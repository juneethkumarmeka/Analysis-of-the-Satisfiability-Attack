module basic_2500_25000_3000_40_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nand U0 (N_0,In_82,In_765);
nor U1 (N_1,In_587,In_1354);
and U2 (N_2,In_2179,In_123);
or U3 (N_3,In_2197,In_2021);
nor U4 (N_4,In_592,In_1819);
and U5 (N_5,In_2267,In_127);
and U6 (N_6,In_1824,In_43);
and U7 (N_7,In_717,In_2441);
or U8 (N_8,In_711,In_1267);
xnor U9 (N_9,In_1784,In_1248);
nor U10 (N_10,In_505,In_2319);
nor U11 (N_11,In_1743,In_2455);
xor U12 (N_12,In_340,In_1995);
nor U13 (N_13,In_1702,In_2271);
and U14 (N_14,In_1509,In_756);
xor U15 (N_15,In_21,In_752);
nor U16 (N_16,In_1302,In_1650);
xnor U17 (N_17,In_1715,In_2272);
or U18 (N_18,In_1393,In_2093);
or U19 (N_19,In_744,In_2183);
or U20 (N_20,In_1944,In_2085);
nor U21 (N_21,In_1659,In_1192);
nand U22 (N_22,In_576,In_1175);
and U23 (N_23,In_512,In_1582);
xor U24 (N_24,In_2376,In_1443);
nor U25 (N_25,In_934,In_166);
xor U26 (N_26,In_821,In_61);
xor U27 (N_27,In_1178,In_282);
xor U28 (N_28,In_295,In_884);
nor U29 (N_29,In_1335,In_2137);
and U30 (N_30,In_2431,In_2445);
xor U31 (N_31,In_1241,In_1775);
nand U32 (N_32,In_213,In_646);
and U33 (N_33,In_984,In_1324);
and U34 (N_34,In_1430,In_1738);
and U35 (N_35,In_2186,In_1841);
or U36 (N_36,In_1952,In_429);
nor U37 (N_37,In_1829,In_411);
and U38 (N_38,In_819,In_2429);
xor U39 (N_39,In_1809,In_815);
nand U40 (N_40,In_1668,In_2022);
or U41 (N_41,In_687,In_1798);
xnor U42 (N_42,In_1135,In_97);
and U43 (N_43,In_300,In_913);
nor U44 (N_44,In_2337,In_1176);
nor U45 (N_45,In_2129,In_2281);
or U46 (N_46,In_113,In_801);
nor U47 (N_47,In_524,In_1867);
or U48 (N_48,In_1918,In_449);
nand U49 (N_49,In_199,In_158);
or U50 (N_50,In_1664,In_1758);
xnor U51 (N_51,In_534,In_255);
nor U52 (N_52,In_1837,In_555);
nand U53 (N_53,In_2471,In_999);
nand U54 (N_54,In_93,In_771);
nor U55 (N_55,In_1202,In_159);
nor U56 (N_56,In_981,In_582);
and U57 (N_57,In_2310,In_1481);
or U58 (N_58,In_50,In_1761);
nand U59 (N_59,In_494,In_693);
nor U60 (N_60,In_1252,In_1941);
nand U61 (N_61,In_948,In_1717);
nor U62 (N_62,In_2472,In_2473);
or U63 (N_63,In_1587,In_1412);
and U64 (N_64,In_691,In_484);
and U65 (N_65,In_1848,In_2059);
or U66 (N_66,In_2460,In_857);
or U67 (N_67,In_457,In_2112);
xor U68 (N_68,In_1359,In_121);
nor U69 (N_69,In_2164,In_925);
and U70 (N_70,In_1682,In_1400);
nand U71 (N_71,In_1705,In_438);
nor U72 (N_72,In_2423,In_883);
and U73 (N_73,In_1862,In_1288);
and U74 (N_74,In_737,In_504);
or U75 (N_75,In_2228,In_2103);
xnor U76 (N_76,In_268,In_877);
or U77 (N_77,In_513,In_2253);
nand U78 (N_78,In_1706,In_1258);
or U79 (N_79,In_788,In_2417);
xor U80 (N_80,In_2362,In_217);
and U81 (N_81,In_1024,In_514);
and U82 (N_82,In_850,In_26);
and U83 (N_83,In_2390,In_361);
xor U84 (N_84,In_810,In_1233);
xnor U85 (N_85,In_1429,In_1933);
nand U86 (N_86,In_720,In_1331);
xnor U87 (N_87,In_1704,In_1234);
and U88 (N_88,In_2291,In_2058);
and U89 (N_89,In_277,In_1467);
xor U90 (N_90,In_214,In_1082);
or U91 (N_91,In_637,In_458);
nor U92 (N_92,In_2344,In_375);
nor U93 (N_93,In_1085,In_1117);
or U94 (N_94,In_2334,In_1218);
nand U95 (N_95,In_1864,In_683);
or U96 (N_96,In_1731,In_702);
and U97 (N_97,In_1576,In_1084);
nand U98 (N_98,In_436,In_254);
nor U99 (N_99,In_498,In_1855);
xor U100 (N_100,In_1732,In_1515);
xnor U101 (N_101,In_951,In_1063);
nand U102 (N_102,In_190,In_986);
and U103 (N_103,In_1080,In_1454);
xor U104 (N_104,In_1247,In_1462);
and U105 (N_105,In_1649,In_1265);
or U106 (N_106,In_152,In_1147);
or U107 (N_107,In_60,In_2213);
xnor U108 (N_108,In_2113,In_526);
nand U109 (N_109,In_1660,In_1527);
and U110 (N_110,In_1860,In_593);
nor U111 (N_111,In_2005,In_615);
nand U112 (N_112,In_732,In_564);
or U113 (N_113,In_1415,In_1012);
and U114 (N_114,In_2225,In_178);
nand U115 (N_115,In_2120,In_2418);
and U116 (N_116,In_349,In_1689);
nand U117 (N_117,In_1273,In_1427);
and U118 (N_118,In_1835,In_1885);
and U119 (N_119,In_2388,In_1710);
nor U120 (N_120,In_599,In_952);
xor U121 (N_121,In_2050,In_1570);
nor U122 (N_122,In_119,In_1103);
xor U123 (N_123,In_1937,In_2410);
nor U124 (N_124,In_1521,In_2248);
xnor U125 (N_125,In_2385,In_1869);
xor U126 (N_126,In_2302,In_729);
nor U127 (N_127,In_1469,In_478);
and U128 (N_128,In_2323,In_1548);
or U129 (N_129,In_380,In_1156);
nor U130 (N_130,In_1368,In_394);
xor U131 (N_131,In_48,In_927);
and U132 (N_132,In_2420,In_2464);
nor U133 (N_133,In_1439,In_929);
nand U134 (N_134,In_16,In_406);
and U135 (N_135,In_1763,In_1399);
nor U136 (N_136,In_56,In_1170);
nand U137 (N_137,In_346,In_2458);
nand U138 (N_138,In_789,In_1380);
and U139 (N_139,In_1264,In_1671);
and U140 (N_140,In_537,In_2081);
xor U141 (N_141,In_1013,In_935);
xnor U142 (N_142,In_1228,In_7);
or U143 (N_143,In_1364,In_1317);
xnor U144 (N_144,In_1046,In_1904);
nand U145 (N_145,In_1594,In_475);
and U146 (N_146,In_1348,In_343);
and U147 (N_147,In_125,In_2140);
nand U148 (N_148,In_1581,In_827);
and U149 (N_149,In_2497,In_1100);
or U150 (N_150,In_2031,In_1930);
nand U151 (N_151,In_654,In_814);
or U152 (N_152,In_2168,In_116);
and U153 (N_153,In_2251,In_303);
or U154 (N_154,In_1795,In_403);
and U155 (N_155,In_1079,In_787);
or U156 (N_156,In_2171,In_2465);
nor U157 (N_157,In_507,In_730);
or U158 (N_158,In_389,In_1994);
nor U159 (N_159,In_2243,In_886);
xor U160 (N_160,In_2208,In_2187);
or U161 (N_161,In_2350,In_226);
and U162 (N_162,In_1459,In_980);
nand U163 (N_163,In_2038,In_973);
nor U164 (N_164,In_1160,In_325);
and U165 (N_165,In_2017,In_1186);
nor U166 (N_166,In_538,In_1398);
nand U167 (N_167,In_1236,In_162);
xor U168 (N_168,In_412,In_1728);
xor U169 (N_169,In_705,In_112);
nand U170 (N_170,In_527,In_2024);
nor U171 (N_171,In_2313,In_1640);
nor U172 (N_172,In_2392,In_578);
xor U173 (N_173,In_597,In_1198);
nor U174 (N_174,In_1676,In_2470);
nor U175 (N_175,In_1433,In_924);
nand U176 (N_176,In_2485,In_841);
or U177 (N_177,In_1998,In_1436);
nor U178 (N_178,In_998,In_1485);
or U179 (N_179,In_1774,In_1711);
nor U180 (N_180,In_1970,In_1655);
or U181 (N_181,In_67,In_292);
or U182 (N_182,In_550,In_760);
nand U183 (N_183,In_1438,In_1628);
nand U184 (N_184,In_1208,In_1183);
and U185 (N_185,In_1,In_910);
xnor U186 (N_186,In_726,In_2249);
xnor U187 (N_187,In_2166,In_695);
and U188 (N_188,In_229,In_1560);
nand U189 (N_189,In_1832,In_14);
and U190 (N_190,In_20,In_305);
or U191 (N_191,In_1406,In_1583);
xnor U192 (N_192,In_2041,In_668);
nand U193 (N_193,In_1982,In_1598);
nor U194 (N_194,In_88,In_2373);
nor U195 (N_195,In_652,In_2034);
nand U196 (N_196,In_182,In_704);
nand U197 (N_197,In_2330,In_2139);
and U198 (N_198,In_2266,In_1672);
nor U199 (N_199,In_1740,In_2071);
nor U200 (N_200,In_501,In_1865);
or U201 (N_201,In_1597,In_1381);
or U202 (N_202,In_710,In_1179);
or U203 (N_203,In_1041,In_803);
or U204 (N_204,In_775,In_692);
or U205 (N_205,In_742,In_1756);
xor U206 (N_206,In_523,In_2199);
nor U207 (N_207,In_1906,In_750);
nand U208 (N_208,In_169,In_1056);
xor U209 (N_209,In_972,In_19);
or U210 (N_210,In_350,In_1644);
nand U211 (N_211,In_2052,In_930);
nand U212 (N_212,In_2459,In_661);
nand U213 (N_213,In_1491,In_189);
and U214 (N_214,In_1356,In_933);
nand U215 (N_215,In_579,In_1677);
xor U216 (N_216,In_2359,In_1159);
and U217 (N_217,In_1118,In_2340);
and U218 (N_218,In_724,In_1440);
nor U219 (N_219,In_263,In_563);
nor U220 (N_220,In_1691,In_3);
nor U221 (N_221,In_1592,In_1000);
or U222 (N_222,In_1185,In_455);
xnor U223 (N_223,In_698,In_792);
nor U224 (N_224,In_1997,In_2185);
or U225 (N_225,In_440,In_804);
nor U226 (N_226,In_1121,In_1723);
xnor U227 (N_227,In_1567,In_1052);
xor U228 (N_228,In_1880,In_1769);
xor U229 (N_229,In_1603,In_84);
xor U230 (N_230,In_674,In_699);
nor U231 (N_231,In_947,In_456);
and U232 (N_232,In_625,In_101);
nand U233 (N_233,In_1311,In_1479);
nand U234 (N_234,In_1981,In_1455);
and U235 (N_235,In_339,In_1210);
nor U236 (N_236,In_1766,In_2076);
nand U237 (N_237,In_596,In_561);
and U238 (N_238,In_1654,In_1757);
nand U239 (N_239,In_1748,In_2073);
nand U240 (N_240,In_535,In_1338);
xor U241 (N_241,In_2082,In_1637);
and U242 (N_242,In_1983,In_1496);
and U243 (N_243,In_1190,In_1653);
and U244 (N_244,In_956,In_1712);
and U245 (N_245,In_805,In_1344);
nand U246 (N_246,In_2428,In_2019);
xnor U247 (N_247,In_1593,In_676);
nor U248 (N_248,In_1600,In_1113);
and U249 (N_249,In_1751,In_1346);
nor U250 (N_250,In_2238,In_1268);
and U251 (N_251,In_74,In_1350);
or U252 (N_252,In_1826,In_2477);
nor U253 (N_253,In_665,In_221);
or U254 (N_254,In_2195,In_1090);
and U255 (N_255,In_2095,In_1441);
nand U256 (N_256,In_2466,In_1701);
nor U257 (N_257,In_892,In_1577);
and U258 (N_258,In_1779,In_1333);
and U259 (N_259,In_1940,In_430);
or U260 (N_260,In_1229,In_212);
nand U261 (N_261,In_660,In_556);
nor U262 (N_262,In_27,In_1822);
nor U263 (N_263,In_586,In_912);
nor U264 (N_264,In_1513,In_1003);
xor U265 (N_265,In_1540,In_868);
nor U266 (N_266,In_5,In_1833);
nor U267 (N_267,In_685,In_1776);
xnor U268 (N_268,In_784,In_2268);
nand U269 (N_269,In_994,In_1942);
nand U270 (N_270,In_1632,In_1029);
nand U271 (N_271,In_181,In_824);
xnor U272 (N_272,In_422,In_2090);
xnor U273 (N_273,In_2210,In_1507);
nor U274 (N_274,In_1352,In_1517);
nor U275 (N_275,In_813,In_2029);
nand U276 (N_276,In_713,In_238);
xor U277 (N_277,In_688,In_1031);
and U278 (N_278,In_1411,In_1726);
nand U279 (N_279,In_1633,In_2496);
nor U280 (N_280,In_271,In_1908);
and U281 (N_281,In_467,In_932);
nor U282 (N_282,In_2227,In_1005);
and U283 (N_283,In_1277,In_383);
nand U284 (N_284,In_274,In_1966);
xor U285 (N_285,In_1887,In_1240);
or U286 (N_286,In_847,In_1017);
or U287 (N_287,In_1999,In_2232);
xnor U288 (N_288,In_552,In_1254);
xor U289 (N_289,In_870,In_366);
or U290 (N_290,In_1503,In_1802);
or U291 (N_291,In_165,In_1066);
and U292 (N_292,In_1518,In_1086);
and U293 (N_293,In_2389,In_1877);
nor U294 (N_294,In_2347,In_1915);
or U295 (N_295,In_37,In_1286);
and U296 (N_296,In_1911,In_2194);
xor U297 (N_297,In_2131,In_1575);
nand U298 (N_298,In_1418,In_989);
nor U299 (N_299,In_1986,In_172);
or U300 (N_300,In_2321,In_2269);
and U301 (N_301,In_1605,In_681);
xor U302 (N_302,In_355,In_1630);
or U303 (N_303,In_1049,In_2259);
nand U304 (N_304,In_1616,In_607);
xor U305 (N_305,In_1670,In_519);
or U306 (N_306,In_2277,In_2457);
xor U307 (N_307,In_2215,In_103);
xnor U308 (N_308,In_269,In_1488);
nand U309 (N_309,In_2386,In_15);
nor U310 (N_310,In_2442,In_2200);
xor U311 (N_311,In_2297,In_2488);
nor U312 (N_312,In_2336,In_2003);
xnor U313 (N_313,In_1935,In_2409);
or U314 (N_314,In_680,In_1604);
or U315 (N_315,In_1285,In_1980);
nor U316 (N_316,In_1355,In_781);
nor U317 (N_317,In_1262,In_915);
and U318 (N_318,In_1667,In_2476);
xnor U319 (N_319,In_1863,In_875);
nor U320 (N_320,In_2155,In_624);
and U321 (N_321,In_584,In_2156);
nor U322 (N_322,In_2008,In_1061);
nor U323 (N_323,In_2494,In_2448);
nor U324 (N_324,In_1133,In_753);
or U325 (N_325,In_1875,In_1501);
or U326 (N_326,In_540,In_1840);
nor U327 (N_327,In_2276,In_2327);
nand U328 (N_328,In_352,In_1790);
xnor U329 (N_329,In_659,In_2088);
and U330 (N_330,In_387,In_1996);
xnor U331 (N_331,In_1688,In_749);
nand U332 (N_332,In_1187,In_1866);
or U333 (N_333,In_942,In_1495);
nand U334 (N_334,In_1168,In_978);
xor U335 (N_335,In_988,In_577);
nor U336 (N_336,In_2127,In_1984);
xor U337 (N_337,In_1016,In_150);
or U338 (N_338,In_823,In_2033);
xor U339 (N_339,In_1416,In_1177);
xnor U340 (N_340,In_2316,In_2468);
xor U341 (N_341,In_2013,In_109);
nor U342 (N_342,In_950,In_1713);
nand U343 (N_343,In_1097,In_1925);
or U344 (N_344,In_469,In_130);
nor U345 (N_345,In_1339,In_1340);
xor U346 (N_346,In_539,In_1145);
nand U347 (N_347,In_2012,In_1098);
or U348 (N_348,In_451,In_1404);
or U349 (N_349,In_920,In_953);
nand U350 (N_350,In_310,In_1217);
nand U351 (N_351,In_1180,In_2001);
nor U352 (N_352,In_746,In_2489);
and U353 (N_353,In_2288,In_2233);
or U354 (N_354,In_1383,In_2105);
nor U355 (N_355,In_32,In_793);
and U356 (N_356,In_1685,In_591);
nor U357 (N_357,In_583,In_156);
and U358 (N_358,In_869,In_1909);
nand U359 (N_359,In_588,In_2252);
or U360 (N_360,In_1902,In_197);
xnor U361 (N_361,In_1326,In_334);
nand U362 (N_362,In_1329,In_1321);
and U363 (N_363,In_1615,In_309);
and U364 (N_364,In_29,In_1621);
and U365 (N_365,In_696,In_1315);
and U366 (N_366,In_606,In_192);
xnor U367 (N_367,In_1992,In_191);
xor U368 (N_368,In_1893,In_376);
and U369 (N_369,In_1261,In_284);
or U370 (N_370,In_1143,In_1303);
and U371 (N_371,In_1754,In_2331);
xor U372 (N_372,In_1222,In_330);
nand U373 (N_373,In_1639,In_2083);
and U374 (N_374,In_2099,In_2175);
nor U375 (N_375,In_671,In_1078);
or U376 (N_376,In_1093,In_293);
xor U377 (N_377,In_1813,In_1461);
nand U378 (N_378,In_1347,In_2294);
nand U379 (N_379,In_1164,In_1225);
nand U380 (N_380,In_1508,In_1746);
nand U381 (N_381,In_2018,In_402);
and U382 (N_382,In_2229,In_2116);
nand U383 (N_383,In_589,In_653);
and U384 (N_384,In_2495,In_890);
nand U385 (N_385,In_2043,In_223);
or U386 (N_386,In_531,In_2256);
or U387 (N_387,In_807,In_2219);
and U388 (N_388,In_2023,In_1945);
xnor U389 (N_389,In_2037,In_997);
nor U390 (N_390,In_517,In_1958);
or U391 (N_391,In_2172,In_1420);
nand U392 (N_392,In_354,In_1679);
nand U393 (N_393,In_2352,In_1382);
nor U394 (N_394,In_2028,In_1808);
or U395 (N_395,In_829,In_2000);
nor U396 (N_396,In_1669,In_686);
xor U397 (N_397,In_1782,In_2318);
nand U398 (N_398,In_1528,In_194);
xnor U399 (N_399,In_2055,In_232);
nand U400 (N_400,In_735,In_1456);
nor U401 (N_401,In_1396,In_1004);
nor U402 (N_402,In_1483,In_766);
xor U403 (N_403,In_2176,In_2221);
nand U404 (N_404,In_2475,In_945);
and U405 (N_405,In_444,In_2415);
nor U406 (N_406,In_1687,In_1112);
xnor U407 (N_407,In_616,In_2380);
and U408 (N_408,In_2371,In_94);
and U409 (N_409,In_610,In_2096);
xnor U410 (N_410,In_1596,In_1988);
or U411 (N_411,In_521,In_1744);
xor U412 (N_412,In_1645,In_278);
nor U413 (N_413,In_969,In_987);
xnor U414 (N_414,In_287,In_1122);
xnor U415 (N_415,In_1614,In_2285);
nor U416 (N_416,In_1874,In_1322);
nor U417 (N_417,In_321,In_393);
xor U418 (N_418,In_64,In_1514);
nor U419 (N_419,In_967,In_1184);
and U420 (N_420,In_522,In_567);
or U421 (N_421,In_1727,In_1349);
nand U422 (N_422,In_80,In_2177);
nor U423 (N_423,In_2400,In_633);
xor U424 (N_424,In_2035,In_891);
nor U425 (N_425,In_2151,In_395);
or U426 (N_426,In_2413,In_2432);
nand U427 (N_427,In_992,In_36);
and U428 (N_428,In_2382,In_1964);
and U429 (N_429,In_888,In_949);
nand U430 (N_430,In_860,In_745);
and U431 (N_431,In_1618,In_1215);
nor U432 (N_432,In_243,In_124);
xnor U433 (N_433,In_432,In_79);
or U434 (N_434,In_427,In_2145);
xor U435 (N_435,In_1408,In_2393);
nand U436 (N_436,In_363,In_357);
nand U437 (N_437,In_2214,In_308);
nand U438 (N_438,In_1846,In_312);
or U439 (N_439,In_1325,In_316);
or U440 (N_440,In_163,In_1033);
xnor U441 (N_441,In_2372,In_1224);
and U442 (N_442,In_8,In_573);
and U443 (N_443,In_1563,In_1094);
or U444 (N_444,In_1536,In_418);
and U445 (N_445,In_2142,In_2286);
xnor U446 (N_446,In_2077,In_1407);
nor U447 (N_447,In_353,In_488);
nand U448 (N_448,In_323,In_1008);
nor U449 (N_449,In_627,In_175);
or U450 (N_450,In_231,In_1607);
nand U451 (N_451,In_799,In_963);
xor U452 (N_452,In_1814,In_1196);
nand U453 (N_453,In_846,In_690);
nor U454 (N_454,In_502,In_1534);
and U455 (N_455,In_2341,In_452);
nand U456 (N_456,In_2306,In_1449);
and U457 (N_457,In_485,In_2170);
xnor U458 (N_458,In_2236,In_1104);
and U459 (N_459,In_1105,In_1213);
and U460 (N_460,In_1316,In_1132);
xor U461 (N_461,In_1070,In_276);
or U462 (N_462,In_1389,In_673);
or U463 (N_463,In_206,In_762);
nand U464 (N_464,In_520,In_544);
or U465 (N_465,In_360,In_2250);
xor U466 (N_466,In_1376,In_533);
nor U467 (N_467,In_441,In_1586);
nor U468 (N_468,In_2365,In_528);
and U469 (N_469,In_10,In_1269);
nand U470 (N_470,In_2182,In_2478);
or U471 (N_471,In_1126,In_768);
xnor U472 (N_472,In_2301,In_1750);
xnor U473 (N_473,In_306,In_1948);
or U474 (N_474,In_1216,In_1551);
and U475 (N_475,In_382,In_2097);
nand U476 (N_476,In_2205,In_714);
nor U477 (N_477,In_1807,In_1367);
xnor U478 (N_478,In_2128,In_1547);
and U479 (N_479,In_2325,In_495);
xor U480 (N_480,In_1162,In_1818);
or U481 (N_481,In_472,In_2079);
and U482 (N_482,In_1073,In_245);
xnor U483 (N_483,In_1535,In_1055);
and U484 (N_484,In_2328,In_408);
and U485 (N_485,In_266,In_2308);
nor U486 (N_486,In_1912,In_2493);
nand U487 (N_487,In_2181,In_1107);
or U488 (N_488,In_828,In_1696);
nand U489 (N_489,In_1419,In_1931);
xor U490 (N_490,In_964,In_1182);
or U491 (N_491,In_2454,In_1036);
xor U492 (N_492,In_725,In_335);
or U493 (N_493,In_1850,In_985);
xor U494 (N_494,In_2235,In_1466);
or U495 (N_495,In_2482,In_2273);
or U496 (N_496,In_1573,In_160);
or U497 (N_497,In_106,In_241);
nand U498 (N_498,In_249,In_1223);
nor U499 (N_499,In_2462,In_58);
or U500 (N_500,In_838,In_2026);
xor U501 (N_501,In_1006,In_2222);
nand U502 (N_502,In_2270,In_2398);
xor U503 (N_503,In_1034,In_837);
nand U504 (N_504,In_52,In_1032);
nor U505 (N_505,In_2346,In_44);
and U506 (N_506,In_1619,In_1313);
nand U507 (N_507,In_2146,In_898);
or U508 (N_508,In_1166,In_405);
nor U509 (N_509,In_1387,In_1805);
xor U510 (N_510,In_235,In_905);
xnor U511 (N_511,In_1881,In_331);
or U512 (N_512,In_1500,In_446);
xnor U513 (N_513,In_859,In_2048);
nand U514 (N_514,In_879,In_1379);
or U515 (N_515,In_701,In_1426);
nand U516 (N_516,In_2204,In_2084);
nand U517 (N_517,In_1658,In_210);
or U518 (N_518,In_1666,In_2074);
nand U519 (N_519,In_1661,In_453);
xnor U520 (N_520,In_1929,In_132);
xor U521 (N_521,In_2191,In_1394);
or U522 (N_522,In_611,In_96);
or U523 (N_523,In_853,In_2122);
nand U524 (N_524,In_634,In_2002);
nor U525 (N_525,In_1845,In_865);
or U526 (N_526,In_2062,In_2007);
xnor U527 (N_527,In_1589,In_222);
xor U528 (N_528,In_1428,In_1295);
xnor U529 (N_529,In_1435,In_2360);
nor U530 (N_530,In_370,In_983);
xor U531 (N_531,In_134,In_2264);
or U532 (N_532,In_940,In_1531);
nor U533 (N_533,In_1559,In_570);
nand U534 (N_534,In_1403,In_1330);
xnor U535 (N_535,In_252,In_2094);
xnor U536 (N_536,In_1519,In_1370);
nor U537 (N_537,In_2339,In_1353);
nand U538 (N_538,In_299,In_251);
nand U539 (N_539,In_1110,In_151);
nand U540 (N_540,In_770,In_1747);
or U541 (N_541,In_2384,In_580);
nand U542 (N_542,In_72,In_54);
nand U543 (N_543,In_198,In_307);
and U544 (N_544,In_2383,In_1762);
xor U545 (N_545,In_1504,In_2421);
xnor U546 (N_546,In_2397,In_2042);
xor U547 (N_547,In_955,In_1889);
or U548 (N_548,In_1623,In_1652);
nand U549 (N_549,In_889,In_1792);
nand U550 (N_550,In_902,In_1384);
xor U551 (N_551,In_2218,In_1884);
nand U552 (N_552,In_1574,In_2154);
xnor U553 (N_553,In_203,In_1657);
or U554 (N_554,In_62,In_1550);
xor U555 (N_555,In_893,In_1291);
nor U556 (N_556,In_1099,In_168);
or U557 (N_557,In_373,In_931);
or U558 (N_558,In_1473,In_81);
nor U559 (N_559,In_809,In_1680);
xnor U560 (N_560,In_842,In_529);
and U561 (N_561,In_220,In_356);
or U562 (N_562,In_620,In_518);
or U563 (N_563,In_1765,In_547);
nor U564 (N_564,In_76,In_1859);
nand U565 (N_565,In_1635,In_1040);
nand U566 (N_566,In_1936,In_1697);
xor U567 (N_567,In_170,In_2387);
nand U568 (N_568,In_2211,In_2064);
nor U569 (N_569,In_854,In_2226);
nor U570 (N_570,In_2299,In_1244);
or U571 (N_571,In_1549,In_908);
nand U572 (N_572,In_397,In_1470);
and U573 (N_573,In_1125,In_55);
and U574 (N_574,In_1625,In_1343);
nor U575 (N_575,In_1725,In_205);
nor U576 (N_576,In_1028,In_290);
nor U577 (N_577,In_1673,In_757);
or U578 (N_578,In_708,In_1457);
xor U579 (N_579,In_911,In_722);
nor U580 (N_580,In_2051,In_1011);
or U581 (N_581,In_542,In_258);
and U582 (N_582,In_230,In_1450);
and U583 (N_583,In_1847,In_872);
and U584 (N_584,In_1502,In_530);
nor U585 (N_585,In_336,In_1719);
and U586 (N_586,In_371,In_1298);
xor U587 (N_587,In_2237,In_1417);
or U588 (N_588,In_463,In_45);
and U589 (N_589,In_1987,In_1764);
and U590 (N_590,In_256,In_1410);
or U591 (N_591,In_2491,In_396);
or U592 (N_592,In_1718,In_715);
xnor U593 (N_593,In_651,In_664);
or U594 (N_594,In_2063,In_1969);
xor U595 (N_595,In_1641,In_1901);
and U596 (N_596,In_1369,In_2463);
xor U597 (N_597,In_2150,In_147);
nand U598 (N_598,In_2449,In_1307);
and U599 (N_599,In_867,In_1195);
nand U600 (N_600,In_234,In_2016);
nor U601 (N_601,In_381,In_35);
or U602 (N_602,In_822,In_1665);
nand U603 (N_603,In_1611,In_2407);
nor U604 (N_604,In_1432,In_2169);
xor U605 (N_605,In_1276,In_1990);
nand U606 (N_606,In_1409,In_1899);
nor U607 (N_607,In_1601,In_979);
or U608 (N_608,In_286,In_2027);
or U609 (N_609,In_1334,In_682);
and U610 (N_610,In_2419,In_92);
or U611 (N_611,In_1283,In_1684);
nor U612 (N_612,In_2114,In_2357);
and U613 (N_613,In_384,In_1448);
and U614 (N_614,In_876,In_2242);
xor U615 (N_615,In_1950,In_684);
or U616 (N_616,In_2298,In_1854);
xnor U617 (N_617,In_129,In_1053);
nand U618 (N_618,In_89,In_1771);
nand U619 (N_619,In_1001,In_608);
nand U620 (N_620,In_95,In_280);
nor U621 (N_621,In_604,In_1043);
xnor U622 (N_622,In_1949,In_49);
nor U623 (N_623,In_2416,In_1836);
xnor U624 (N_624,In_434,In_1249);
and U625 (N_625,In_195,In_2287);
xor U626 (N_626,In_289,In_2098);
nand U627 (N_627,N_119,In_937);
nand U628 (N_628,N_190,In_2424);
xnor U629 (N_629,In_2486,N_489);
nand U630 (N_630,In_1402,In_385);
and U631 (N_631,In_901,N_215);
and U632 (N_632,N_405,In_1245);
nor U633 (N_633,In_24,In_2080);
xnor U634 (N_634,N_184,In_111);
nor U635 (N_635,In_491,In_1760);
and U636 (N_636,In_1562,In_2136);
nand U637 (N_637,N_505,In_1991);
xnor U638 (N_638,In_738,N_612);
and U639 (N_639,N_545,In_509);
xor U640 (N_640,In_1203,In_907);
and U641 (N_641,N_36,In_1968);
or U642 (N_642,N_319,N_459);
xnor U643 (N_643,In_322,In_1900);
xnor U644 (N_644,In_391,In_574);
or U645 (N_645,In_764,N_235);
or U646 (N_646,N_279,N_619);
nand U647 (N_647,In_635,In_1327);
nor U648 (N_648,In_2435,In_786);
xnor U649 (N_649,In_31,N_92);
xnor U650 (N_650,N_9,In_2040);
xor U651 (N_651,In_723,N_604);
xnor U652 (N_652,N_167,In_1868);
xor U653 (N_653,N_504,In_272);
nand U654 (N_654,N_299,N_603);
xor U655 (N_655,In_2123,In_551);
xnor U656 (N_656,In_874,N_611);
or U657 (N_657,N_97,In_239);
nand U658 (N_658,In_1351,N_332);
nor U659 (N_659,In_1972,In_264);
nand U660 (N_660,In_1042,N_82);
and U661 (N_661,In_51,In_1478);
and U662 (N_662,N_418,In_957);
xnor U663 (N_663,In_431,In_1569);
nand U664 (N_664,In_1272,In_1974);
or U665 (N_665,N_188,In_187);
nor U666 (N_666,In_1259,In_2369);
or U667 (N_667,In_763,In_2109);
or U668 (N_668,In_970,In_1674);
or U669 (N_669,N_113,N_433);
and U670 (N_670,N_453,N_352);
nor U671 (N_671,N_227,In_1486);
nor U672 (N_672,In_1894,In_2351);
or U673 (N_673,In_1119,In_137);
and U674 (N_674,In_25,In_1737);
or U675 (N_675,In_1979,In_138);
and U676 (N_676,In_1293,N_272);
and U677 (N_677,In_1511,N_137);
xnor U678 (N_678,N_281,N_91);
nor U679 (N_679,In_663,N_416);
xnor U680 (N_680,In_1212,In_855);
xor U681 (N_681,In_739,In_1921);
nor U682 (N_682,In_941,In_1345);
and U683 (N_683,In_426,N_498);
nand U684 (N_684,In_2216,N_253);
or U685 (N_685,In_808,In_1492);
and U686 (N_686,In_2303,In_2108);
nor U687 (N_687,In_1539,In_2452);
or U688 (N_688,In_1361,In_2147);
or U689 (N_689,N_476,N_597);
nor U690 (N_690,N_39,In_1963);
or U691 (N_691,In_1741,N_134);
and U692 (N_692,N_29,In_69);
nand U693 (N_693,N_528,In_2160);
nand U694 (N_694,In_110,In_2348);
nor U695 (N_695,In_2030,N_24);
or U696 (N_696,In_358,N_491);
or U697 (N_697,In_1363,In_22);
nor U698 (N_698,In_133,In_1067);
xnor U699 (N_699,In_1505,In_34);
xnor U700 (N_700,In_777,In_1136);
or U701 (N_701,In_2133,In_2453);
or U702 (N_702,In_1015,In_594);
nand U703 (N_703,N_204,N_292);
or U704 (N_704,N_359,In_778);
nor U705 (N_705,N_469,N_483);
xor U706 (N_706,N_51,In_291);
or U707 (N_707,In_1220,In_759);
or U708 (N_708,N_187,In_921);
and U709 (N_709,N_307,N_112);
and U710 (N_710,In_1161,N_549);
nand U711 (N_711,N_601,In_1072);
xnor U712 (N_712,In_557,N_270);
nand U713 (N_713,In_1038,In_1266);
xor U714 (N_714,N_74,In_1150);
or U715 (N_715,In_1827,In_302);
and U716 (N_716,In_1445,N_515);
and U717 (N_717,In_1755,In_1544);
nor U718 (N_718,N_560,In_1318);
nor U719 (N_719,In_1799,In_1197);
and U720 (N_720,In_490,N_62);
or U721 (N_721,In_219,N_143);
and U722 (N_722,In_17,N_339);
nand U723 (N_723,N_107,In_1871);
or U724 (N_724,N_42,N_219);
nor U725 (N_725,In_2363,In_2207);
or U726 (N_726,In_174,In_1722);
nand U727 (N_727,In_1768,In_77);
xor U728 (N_728,In_341,N_524);
and U729 (N_729,In_914,In_811);
and U730 (N_730,In_670,In_1852);
and U731 (N_731,In_734,In_1437);
nor U732 (N_732,N_535,In_751);
and U733 (N_733,In_543,In_712);
nand U734 (N_734,In_1898,N_105);
nor U735 (N_735,In_636,In_2364);
nor U736 (N_736,In_208,In_65);
or U737 (N_737,In_2403,In_906);
or U738 (N_738,In_1919,In_1913);
xnor U739 (N_739,N_362,In_640);
nand U740 (N_740,In_975,In_2283);
or U741 (N_741,In_1773,N_141);
or U742 (N_742,In_1643,N_309);
nor U743 (N_743,In_2230,N_344);
or U744 (N_744,In_1844,In_2324);
and U745 (N_745,N_381,N_160);
or U746 (N_746,In_117,In_28);
or U747 (N_747,N_580,In_1377);
nor U748 (N_748,N_199,In_2244);
nor U749 (N_749,In_796,In_1825);
and U750 (N_750,In_1714,In_641);
nand U751 (N_751,In_1171,In_672);
nor U752 (N_752,In_1638,In_1444);
or U753 (N_753,N_413,N_566);
xor U754 (N_754,In_120,In_2006);
nor U755 (N_755,In_18,In_1214);
and U756 (N_756,In_1555,In_740);
xor U757 (N_757,In_1199,N_492);
xnor U758 (N_758,In_2447,In_301);
nand U759 (N_759,In_39,N_77);
nand U760 (N_760,N_325,In_1800);
nand U761 (N_761,In_916,N_590);
nand U762 (N_762,N_320,In_242);
xor U763 (N_763,In_2246,In_483);
nor U764 (N_764,In_1193,In_1853);
xnor U765 (N_765,In_1336,N_126);
or U766 (N_766,N_499,In_2111);
nand U767 (N_767,In_183,In_1453);
nor U768 (N_768,N_130,In_1204);
nand U769 (N_769,N_114,In_1613);
nand U770 (N_770,N_466,In_173);
xor U771 (N_771,N_511,N_19);
or U772 (N_772,In_1786,N_95);
nor U773 (N_773,In_460,N_58);
nand U774 (N_774,N_220,N_437);
or U775 (N_775,In_1525,N_131);
nand U776 (N_776,In_541,N_371);
xor U777 (N_777,In_466,In_1498);
nand U778 (N_778,N_121,In_817);
or U779 (N_779,In_1554,N_496);
nand U780 (N_780,In_2422,In_1116);
or U781 (N_781,In_590,N_506);
nand U782 (N_782,N_264,N_523);
xor U783 (N_783,N_334,N_152);
or U784 (N_784,N_585,In_1320);
nor U785 (N_785,In_2135,In_224);
and U786 (N_786,In_628,In_1910);
xor U787 (N_787,In_612,In_122);
xnor U788 (N_788,In_257,N_522);
or U789 (N_789,In_317,In_840);
or U790 (N_790,N_529,N_103);
or U791 (N_791,N_539,N_395);
xnor U792 (N_792,N_6,N_48);
and U793 (N_793,In_2367,In_562);
or U794 (N_794,In_6,In_2193);
xor U795 (N_795,In_1699,N_425);
nand U796 (N_796,In_1069,N_426);
nand U797 (N_797,In_1044,In_1451);
nor U798 (N_798,N_538,In_897);
and U799 (N_799,N_193,N_596);
or U800 (N_800,In_1882,In_1231);
nand U801 (N_801,In_12,N_370);
nand U802 (N_802,In_2057,N_258);
or U803 (N_803,N_34,In_558);
nand U804 (N_804,In_603,N_100);
xor U805 (N_805,N_449,In_1065);
or U806 (N_806,In_270,In_2241);
xnor U807 (N_807,In_1903,N_558);
and U808 (N_808,N_599,N_290);
nand U809 (N_809,N_398,N_280);
or U810 (N_810,In_454,N_237);
nand U811 (N_811,In_2220,In_1332);
and U812 (N_812,In_873,In_1849);
nor U813 (N_813,In_1695,In_852);
nand U814 (N_814,In_1174,In_2284);
and U815 (N_815,In_2474,In_1310);
nand U816 (N_816,N_254,In_157);
nand U817 (N_817,N_366,In_812);
nand U818 (N_818,N_93,N_348);
and U819 (N_819,In_209,In_525);
nor U820 (N_820,In_177,In_386);
and U821 (N_821,N_620,N_602);
or U822 (N_822,In_1924,N_442);
xor U823 (N_823,In_974,In_1624);
nor U824 (N_824,In_283,In_2192);
nor U825 (N_825,N_456,N_458);
xor U826 (N_826,In_2434,In_2072);
nand U827 (N_827,In_1300,In_423);
nand U828 (N_828,In_848,In_344);
and U829 (N_829,In_1692,In_769);
nand U830 (N_830,N_83,In_1281);
or U831 (N_831,In_1753,In_2437);
and U832 (N_832,In_1083,N_85);
xor U833 (N_833,In_1081,In_894);
nor U834 (N_834,In_631,In_1048);
xor U835 (N_835,In_546,In_1154);
nor U836 (N_836,In_694,In_420);
or U837 (N_837,N_519,In_944);
xor U838 (N_838,N_562,In_1787);
or U839 (N_839,N_229,N_192);
nor U840 (N_840,In_1270,In_1811);
xnor U841 (N_841,In_1690,In_2138);
nor U842 (N_842,In_2209,N_11);
and U843 (N_843,In_1305,In_1130);
or U844 (N_844,In_1626,In_1565);
xnor U845 (N_845,In_9,In_1497);
xor U846 (N_846,In_943,N_159);
and U847 (N_847,N_53,N_401);
xor U848 (N_848,In_2101,In_2345);
and U849 (N_849,In_510,In_748);
nand U850 (N_850,In_831,N_372);
or U851 (N_851,In_959,In_605);
nor U852 (N_852,N_336,N_135);
xor U853 (N_853,In_566,In_1716);
nand U854 (N_854,In_658,N_407);
nor U855 (N_855,In_2356,In_1371);
nor U856 (N_856,N_145,In_131);
and U857 (N_857,In_1405,In_1522);
nand U858 (N_858,In_1308,In_2107);
xnor U859 (N_859,In_2290,In_57);
nand U860 (N_860,In_733,N_308);
xor U861 (N_861,In_1646,In_1250);
and U862 (N_862,N_358,In_2342);
nor U863 (N_863,In_2265,N_615);
and U864 (N_864,In_1778,In_861);
xor U865 (N_865,In_2296,In_23);
or U866 (N_866,In_362,N_500);
nor U867 (N_867,In_1879,In_318);
and U868 (N_868,N_548,N_326);
xor U869 (N_869,N_108,In_2255);
nand U870 (N_870,In_204,N_86);
nand U871 (N_871,In_347,In_1932);
or U872 (N_872,N_559,N_49);
nand U873 (N_873,In_1709,In_2333);
or U874 (N_874,N_123,In_1460);
xnor U875 (N_875,In_1976,In_832);
nor U876 (N_876,In_1791,N_213);
nand U877 (N_877,N_411,In_1817);
or U878 (N_878,In_1951,In_244);
xnor U879 (N_879,In_839,In_1770);
nand U880 (N_880,In_297,N_365);
nor U881 (N_881,N_544,In_677);
nand U882 (N_882,N_387,In_1238);
xnor U883 (N_883,In_1591,In_2282);
or U884 (N_884,N_89,N_570);
and U885 (N_885,In_1357,In_2100);
nand U886 (N_886,In_1752,In_2223);
nand U887 (N_887,In_1595,In_1662);
xnor U888 (N_888,N_179,In_565);
and U889 (N_889,In_1388,In_1678);
and U890 (N_890,In_90,N_110);
or U891 (N_891,In_2295,In_262);
xor U892 (N_892,In_1392,N_587);
and U893 (N_893,In_1922,In_148);
xnor U894 (N_894,In_2061,In_1141);
nor U895 (N_895,In_703,In_1584);
nand U896 (N_896,In_1129,In_1561);
nor U897 (N_897,In_1301,In_2180);
and U898 (N_898,In_783,N_55);
xnor U899 (N_899,N_50,In_878);
or U900 (N_900,N_480,In_2130);
or U901 (N_901,N_195,N_256);
nor U902 (N_902,In_1172,N_534);
xor U903 (N_903,N_269,N_494);
or U904 (N_904,N_59,In_2412);
nand U905 (N_905,In_433,N_317);
xor U906 (N_906,In_2190,N_305);
nor U907 (N_907,In_1794,In_1749);
xor U908 (N_908,In_666,N_233);
nor U909 (N_909,In_2198,In_1961);
nand U910 (N_910,N_10,In_1458);
xor U911 (N_911,N_324,N_331);
xnor U912 (N_912,In_1907,In_553);
xor U913 (N_913,In_864,In_2370);
and U914 (N_914,N_207,In_2010);
xnor U915 (N_915,N_22,N_261);
and U916 (N_916,N_47,In_772);
nand U917 (N_917,In_2396,N_439);
nor U918 (N_918,N_536,In_2158);
and U919 (N_919,N_461,In_2305);
xor U920 (N_920,In_1804,In_100);
or U921 (N_921,In_439,N_424);
and U922 (N_922,In_2425,In_1390);
and U923 (N_923,N_447,In_63);
xor U924 (N_924,In_98,In_961);
or U925 (N_925,In_1721,In_858);
and U926 (N_926,In_1516,In_638);
nor U927 (N_927,In_960,N_474);
xnor U928 (N_928,In_1109,In_2202);
or U929 (N_929,In_1955,In_1447);
and U930 (N_930,In_643,In_754);
nand U931 (N_931,In_516,In_2184);
nand U932 (N_932,In_462,N_115);
or U933 (N_933,In_2404,In_329);
nor U934 (N_934,N_132,N_181);
nand U935 (N_935,In_1279,N_228);
nor U936 (N_936,In_1720,In_2436);
or U937 (N_937,N_383,N_478);
xnor U938 (N_938,In_294,In_946);
and U939 (N_939,N_273,In_1201);
and U940 (N_940,N_482,N_568);
nor U941 (N_941,N_185,In_70);
nor U942 (N_942,In_1360,In_1027);
or U943 (N_943,In_415,In_179);
xnor U944 (N_944,In_71,N_20);
and U945 (N_945,In_497,N_431);
xor U946 (N_946,In_871,In_779);
xnor U947 (N_947,In_1373,N_440);
nor U948 (N_948,N_166,In_962);
nor U949 (N_949,N_212,In_273);
nor U950 (N_950,In_1506,N_87);
xnor U951 (N_951,In_1205,N_313);
and U952 (N_952,In_1167,In_790);
and U953 (N_953,In_421,In_1123);
xnor U954 (N_954,In_794,In_1781);
nand U955 (N_955,In_1480,N_246);
nor U956 (N_956,N_139,In_1928);
and U957 (N_957,In_2315,N_532);
nor U958 (N_958,In_2262,In_1629);
nor U959 (N_959,In_1739,N_162);
nand U960 (N_960,In_320,In_2378);
xor U961 (N_961,In_78,N_406);
and U962 (N_962,In_1856,N_35);
nand U963 (N_963,N_224,N_283);
nand U964 (N_964,In_1953,In_399);
nand U965 (N_965,In_2375,N_127);
and U966 (N_966,In_644,In_1227);
nor U967 (N_967,In_1149,N_443);
or U968 (N_968,In_348,In_87);
xor U969 (N_969,In_171,In_114);
xor U970 (N_970,In_1708,In_1627);
and U971 (N_971,N_520,In_196);
and U972 (N_972,In_1642,In_679);
nand U973 (N_973,In_2163,In_1366);
and U974 (N_974,N_382,In_1188);
xor U975 (N_975,In_1858,N_533);
nor U976 (N_976,N_14,In_164);
nor U977 (N_977,N_584,In_1284);
nor U978 (N_978,In_1058,N_551);
nor U979 (N_979,N_484,N_457);
nor U980 (N_980,In_2430,In_1465);
and U981 (N_981,In_493,In_954);
nor U982 (N_982,N_554,In_1181);
xor U983 (N_983,N_609,N_12);
nand U984 (N_984,In_1489,N_88);
nor U985 (N_985,In_149,In_2);
nand U986 (N_986,In_2143,In_1590);
xnor U987 (N_987,In_459,In_926);
nor U988 (N_988,In_180,In_153);
nand U989 (N_989,In_2408,N_242);
and U990 (N_990,In_73,N_202);
and U991 (N_991,In_1111,In_1108);
and U992 (N_992,N_385,N_189);
or U993 (N_993,In_1051,In_11);
nand U994 (N_994,In_1287,In_996);
nand U995 (N_995,In_379,N_1);
nand U996 (N_996,N_412,N_222);
nand U997 (N_997,In_68,In_1023);
nand U998 (N_998,N_296,N_374);
nor U999 (N_999,N_221,In_1342);
or U1000 (N_1000,In_1742,In_1698);
nor U1001 (N_1001,In_863,In_1905);
nand U1002 (N_1002,In_2086,N_510);
nor U1003 (N_1003,In_2279,In_650);
nor U1004 (N_1004,N_297,In_2092);
and U1005 (N_1005,In_259,N_278);
or U1006 (N_1006,In_1421,In_508);
or U1007 (N_1007,N_378,In_1128);
nand U1008 (N_1008,In_480,In_2068);
nand U1009 (N_1009,In_568,In_656);
nand U1010 (N_1010,In_146,In_834);
xnor U1011 (N_1011,In_1472,N_201);
nor U1012 (N_1012,In_1971,In_2374);
or U1013 (N_1013,In_465,In_1530);
nand U1014 (N_1014,In_601,In_1602);
nor U1015 (N_1015,In_1253,N_621);
xnor U1016 (N_1016,In_845,In_728);
nor U1017 (N_1017,In_900,In_1943);
xnor U1018 (N_1018,In_46,N_565);
nor U1019 (N_1019,N_285,In_572);
nor U1020 (N_1020,N_196,In_2368);
xnor U1021 (N_1021,N_605,In_785);
xor U1022 (N_1022,In_492,N_432);
and U1023 (N_1023,In_409,N_571);
xnor U1024 (N_1024,In_1237,In_1736);
and U1025 (N_1025,In_791,N_479);
xor U1026 (N_1026,N_485,In_136);
or U1027 (N_1027,N_388,In_1985);
nand U1028 (N_1028,In_1803,N_60);
nand U1029 (N_1029,In_2487,In_1612);
nand U1030 (N_1030,In_856,In_1939);
nor U1031 (N_1031,N_303,In_2217);
or U1032 (N_1032,In_1263,In_1965);
nand U1033 (N_1033,N_284,In_365);
and U1034 (N_1034,In_1290,N_206);
nand U1035 (N_1035,N_301,N_214);
nand U1036 (N_1036,N_589,In_104);
or U1037 (N_1037,In_706,In_2104);
xor U1038 (N_1038,In_1579,In_2335);
and U1039 (N_1039,In_2261,In_2377);
xor U1040 (N_1040,In_1442,In_1068);
and U1041 (N_1041,N_396,In_881);
or U1042 (N_1042,N_417,In_825);
xnor U1043 (N_1043,In_202,In_1524);
and U1044 (N_1044,In_1092,In_1337);
and U1045 (N_1045,In_773,In_2047);
and U1046 (N_1046,In_1014,In_767);
or U1047 (N_1047,In_2293,N_473);
or U1048 (N_1048,In_1585,In_1634);
and U1049 (N_1049,In_1144,In_2132);
xnor U1050 (N_1050,In_2115,In_851);
xor U1051 (N_1051,In_1365,In_1401);
and U1052 (N_1052,In_2044,In_899);
nand U1053 (N_1053,N_490,In_1959);
nor U1054 (N_1054,In_1914,In_776);
nor U1055 (N_1055,In_826,N_606);
nand U1056 (N_1056,In_145,N_355);
or U1057 (N_1057,N_488,In_2484);
xnor U1058 (N_1058,In_240,In_2014);
or U1059 (N_1059,In_1271,In_849);
nor U1060 (N_1060,In_142,In_265);
nand U1061 (N_1061,N_150,In_1543);
and U1062 (N_1062,In_1246,In_569);
nand U1063 (N_1063,In_338,N_541);
xnor U1064 (N_1064,In_1686,In_2289);
and U1065 (N_1065,In_1173,In_424);
nand U1066 (N_1066,In_1045,In_2032);
or U1067 (N_1067,N_578,In_675);
nor U1068 (N_1068,In_536,N_226);
nand U1069 (N_1069,In_2174,N_312);
nand U1070 (N_1070,In_369,N_76);
or U1071 (N_1071,In_1493,N_80);
xor U1072 (N_1072,N_438,In_1309);
and U1073 (N_1073,N_0,In_1830);
nand U1074 (N_1074,N_464,In_1475);
nor U1075 (N_1075,In_107,In_218);
nor U1076 (N_1076,In_1636,In_237);
nand U1077 (N_1077,In_2309,In_1648);
xnor U1078 (N_1078,N_30,In_66);
and U1079 (N_1079,In_2203,N_247);
nand U1080 (N_1080,In_1341,In_139);
nor U1081 (N_1081,In_1242,N_477);
or U1082 (N_1082,In_4,In_435);
and U1083 (N_1083,In_2358,In_655);
nand U1084 (N_1084,N_593,N_225);
nor U1085 (N_1085,In_461,N_588);
nand U1086 (N_1086,N_318,In_261);
xnor U1087 (N_1087,In_1206,In_2254);
xnor U1088 (N_1088,N_537,In_797);
or U1089 (N_1089,N_300,N_163);
nand U1090 (N_1090,In_1251,In_982);
nand U1091 (N_1091,In_2499,In_1895);
or U1092 (N_1092,In_1975,N_579);
xor U1093 (N_1093,In_419,N_399);
nor U1094 (N_1094,In_1815,In_820);
and U1095 (N_1095,In_1468,N_350);
or U1096 (N_1096,In_1089,In_621);
or U1097 (N_1097,In_1102,In_1088);
or U1098 (N_1098,In_2015,In_359);
or U1099 (N_1099,N_268,N_321);
nand U1100 (N_1100,N_393,In_1148);
nand U1101 (N_1101,N_521,In_499);
xnor U1102 (N_1102,N_617,N_117);
nand U1103 (N_1103,N_428,N_248);
nor U1104 (N_1104,In_33,In_1883);
or U1105 (N_1105,N_52,N_346);
or U1106 (N_1106,In_410,In_193);
and U1107 (N_1107,In_2426,In_909);
xnor U1108 (N_1108,In_958,N_391);
and U1109 (N_1109,In_1796,N_338);
or U1110 (N_1110,In_1057,N_118);
nand U1111 (N_1111,N_155,In_2165);
xor U1112 (N_1112,N_335,In_741);
and U1113 (N_1113,In_843,In_1037);
nor U1114 (N_1114,In_993,In_1211);
nand U1115 (N_1115,In_2274,N_404);
and U1116 (N_1116,N_41,N_260);
nand U1117 (N_1117,In_1151,N_147);
nand U1118 (N_1118,N_133,In_1730);
xnor U1119 (N_1119,N_44,N_380);
or U1120 (N_1120,N_530,N_68);
xnor U1121 (N_1121,In_1002,In_246);
nand U1122 (N_1122,N_218,N_574);
or U1123 (N_1123,N_63,In_13);
or U1124 (N_1124,In_1810,In_1891);
nor U1125 (N_1125,In_1425,In_2411);
or U1126 (N_1126,N_16,In_118);
nor U1127 (N_1127,In_1610,In_1025);
and U1128 (N_1128,In_1647,In_1050);
nand U1129 (N_1129,In_1675,In_835);
xor U1130 (N_1130,In_342,N_598);
and U1131 (N_1131,In_1523,N_69);
and U1132 (N_1132,N_4,N_54);
nand U1133 (N_1133,In_2110,In_1564);
xnor U1134 (N_1134,In_1512,In_1463);
xnor U1135 (N_1135,In_367,In_176);
nor U1136 (N_1136,In_2054,In_1124);
or U1137 (N_1137,N_231,N_102);
nor U1138 (N_1138,In_2451,N_198);
nor U1139 (N_1139,In_2479,N_168);
nand U1140 (N_1140,In_102,N_509);
nor U1141 (N_1141,In_1312,In_2075);
xnor U1142 (N_1142,In_474,N_450);
nor U1143 (N_1143,In_161,In_40);
nand U1144 (N_1144,In_2300,N_576);
nand U1145 (N_1145,N_333,N_122);
xnor U1146 (N_1146,In_285,In_2091);
nand U1147 (N_1147,N_67,In_228);
or U1148 (N_1148,In_486,N_327);
or U1149 (N_1149,In_2125,In_721);
nor U1150 (N_1150,N_503,N_345);
or U1151 (N_1151,In_425,In_75);
or U1152 (N_1152,In_1131,N_448);
or U1153 (N_1153,In_1838,In_2427);
xnor U1154 (N_1154,In_216,In_1477);
or U1155 (N_1155,N_177,N_194);
and U1156 (N_1156,In_1256,N_573);
or U1157 (N_1157,In_2469,In_345);
and U1158 (N_1158,In_1446,N_614);
nand U1159 (N_1159,N_397,In_1482);
nor U1160 (N_1160,In_2292,N_267);
or U1161 (N_1161,N_341,In_1993);
xnor U1162 (N_1162,In_1385,In_991);
and U1163 (N_1163,In_1064,In_1842);
and U1164 (N_1164,N_197,N_454);
nand U1165 (N_1165,In_1663,N_158);
nand U1166 (N_1166,N_337,In_798);
nand U1167 (N_1167,In_2307,In_816);
xnor U1168 (N_1168,In_1413,In_108);
nor U1169 (N_1169,In_1278,In_313);
and U1170 (N_1170,In_1035,In_1538);
and U1171 (N_1171,In_1568,N_156);
and U1172 (N_1172,In_1872,N_239);
xor U1173 (N_1173,In_1529,In_2304);
nor U1174 (N_1174,In_2070,N_400);
and U1175 (N_1175,N_361,In_2036);
or U1176 (N_1176,N_322,In_2144);
or U1177 (N_1177,N_543,In_2067);
or U1178 (N_1178,N_363,In_2060);
or U1179 (N_1179,In_667,N_569);
or U1180 (N_1180,In_476,In_414);
nor U1181 (N_1181,In_882,N_592);
nor U1182 (N_1182,In_91,N_98);
nand U1183 (N_1183,In_1306,In_2141);
xor U1184 (N_1184,In_619,In_2446);
xnor U1185 (N_1185,In_2153,N_357);
and U1186 (N_1186,In_1707,In_443);
nor U1187 (N_1187,In_1816,In_2467);
and U1188 (N_1188,In_143,In_1510);
or U1189 (N_1189,In_1831,N_471);
xor U1190 (N_1190,N_101,In_885);
nor U1191 (N_1191,In_1734,In_645);
or U1192 (N_1192,In_1978,In_719);
nor U1193 (N_1193,In_1681,In_59);
and U1194 (N_1194,In_662,N_154);
nor U1195 (N_1195,In_326,N_460);
or U1196 (N_1196,N_208,N_186);
or U1197 (N_1197,N_600,N_72);
or U1198 (N_1198,N_15,In_1243);
nor U1199 (N_1199,N_517,In_1414);
nor U1200 (N_1200,In_186,N_21);
xor U1201 (N_1201,In_2379,In_1916);
and U1202 (N_1202,In_500,N_330);
nor U1203 (N_1203,N_81,N_513);
or U1204 (N_1204,N_146,In_758);
xnor U1205 (N_1205,In_1471,In_2196);
and U1206 (N_1206,N_294,N_203);
nor U1207 (N_1207,In_731,N_8);
xor U1208 (N_1208,N_575,In_250);
nand U1209 (N_1209,N_251,In_938);
nand U1210 (N_1210,In_647,In_253);
and U1211 (N_1211,In_281,In_795);
nor U1212 (N_1212,In_140,In_2124);
and U1213 (N_1213,In_2355,In_1059);
or U1214 (N_1214,In_2322,N_28);
and U1215 (N_1215,In_47,In_1431);
nor U1216 (N_1216,N_472,In_1920);
and U1217 (N_1217,N_209,In_1280);
xor U1218 (N_1218,In_1009,In_1372);
xnor U1219 (N_1219,In_2149,In_581);
nand U1220 (N_1220,N_149,N_408);
nand U1221 (N_1221,In_1622,In_1297);
xor U1222 (N_1222,N_314,In_623);
and U1223 (N_1223,In_1155,In_600);
or U1224 (N_1224,In_1537,In_400);
nand U1225 (N_1225,N_169,In_2443);
or U1226 (N_1226,In_2134,N_531);
nor U1227 (N_1227,N_252,N_390);
nor U1228 (N_1228,N_501,In_1464);
xor U1229 (N_1229,In_144,In_1703);
nor U1230 (N_1230,N_266,N_323);
xnor U1231 (N_1231,In_1546,In_1843);
and U1232 (N_1232,N_26,In_207);
or U1233 (N_1233,In_1422,N_43);
nand U1234 (N_1234,In_155,N_125);
nand U1235 (N_1235,In_2314,In_2087);
xnor U1236 (N_1236,In_2157,In_445);
nor U1237 (N_1237,In_1077,In_1021);
xor U1238 (N_1238,N_607,In_1207);
and U1239 (N_1239,N_613,In_1780);
and U1240 (N_1240,In_2414,In_2401);
xor U1241 (N_1241,In_1114,N_557);
or U1242 (N_1242,In_2121,In_2332);
and U1243 (N_1243,In_976,N_245);
xnor U1244 (N_1244,In_1870,In_966);
nand U1245 (N_1245,N_244,In_2320);
or U1246 (N_1246,N_507,In_971);
xor U1247 (N_1247,N_161,In_718);
xnor U1248 (N_1248,In_1886,In_669);
nor U1249 (N_1249,In_1423,In_1018);
xnor U1250 (N_1250,N_263,In_1296);
nor U1251 (N_1251,N_232,N_708);
nor U1252 (N_1252,N_1183,In_1759);
xor U1253 (N_1253,N_384,In_388);
xnor U1254 (N_1254,In_2438,In_939);
xnor U1255 (N_1255,N_928,N_815);
and U1256 (N_1256,N_806,N_655);
nand U1257 (N_1257,N_861,In_560);
nand U1258 (N_1258,N_1227,In_1434);
xor U1259 (N_1259,N_61,N_1236);
or U1260 (N_1260,N_894,In_2405);
nor U1261 (N_1261,In_617,In_154);
or U1262 (N_1262,N_7,N_1234);
nor U1263 (N_1263,In_2326,In_236);
and U1264 (N_1264,N_730,In_1923);
nand U1265 (N_1265,In_1828,N_635);
or U1266 (N_1266,N_1134,N_46);
nand U1267 (N_1267,In_315,N_1242);
nor U1268 (N_1268,N_637,N_937);
and U1269 (N_1269,N_249,N_839);
and U1270 (N_1270,N_701,N_402);
nand U1271 (N_1271,In_515,In_622);
and U1272 (N_1272,In_1299,N_183);
and U1273 (N_1273,N_713,N_784);
and U1274 (N_1274,In_378,N_631);
nand U1275 (N_1275,In_1047,N_610);
xnor U1276 (N_1276,N_1042,In_401);
xor U1277 (N_1277,In_1588,N_809);
xor U1278 (N_1278,In_2004,N_1157);
or U1279 (N_1279,N_658,N_435);
nand U1280 (N_1280,N_1012,N_1002);
xor U1281 (N_1281,N_745,N_756);
and U1282 (N_1282,N_879,In_1319);
nor U1283 (N_1283,N_1057,In_2490);
xnor U1284 (N_1284,In_727,N_866);
xor U1285 (N_1285,N_904,In_928);
nor U1286 (N_1286,N_451,N_851);
xnor U1287 (N_1287,N_1114,N_342);
xnor U1288 (N_1288,N_240,N_1237);
and U1289 (N_1289,In_554,N_75);
xor U1290 (N_1290,N_1080,In_1897);
xor U1291 (N_1291,N_641,In_1729);
and U1292 (N_1292,N_389,N_176);
or U1293 (N_1293,In_1153,N_753);
or U1294 (N_1294,In_1926,N_236);
nand U1295 (N_1295,N_316,N_885);
nor U1296 (N_1296,N_1177,In_1651);
nand U1297 (N_1297,N_487,In_1395);
nand U1298 (N_1298,In_1358,N_709);
and U1299 (N_1299,N_1179,In_1158);
and U1300 (N_1300,N_157,In_1294);
nand U1301 (N_1301,N_1051,N_38);
and U1302 (N_1302,N_785,In_225);
nand U1303 (N_1303,In_1499,N_1142);
and U1304 (N_1304,In_1007,N_174);
nor U1305 (N_1305,In_678,In_904);
xnor U1306 (N_1306,N_1232,N_719);
or U1307 (N_1307,N_802,N_693);
nand U1308 (N_1308,In_1533,In_774);
and U1309 (N_1309,N_1238,N_1054);
xnor U1310 (N_1310,N_1031,In_1375);
nor U1311 (N_1311,N_875,In_2311);
nor U1312 (N_1312,In_1812,N_1219);
and U1313 (N_1313,N_275,In_1275);
nand U1314 (N_1314,N_677,In_2395);
nor U1315 (N_1315,N_271,In_470);
nor U1316 (N_1316,In_1700,In_632);
or U1317 (N_1317,N_165,N_1116);
nor U1318 (N_1318,N_563,N_1035);
or U1319 (N_1319,N_1241,N_564);
and U1320 (N_1320,In_2381,N_369);
and U1321 (N_1321,N_796,N_1158);
or U1322 (N_1322,N_741,N_422);
or U1323 (N_1323,N_778,N_1001);
nor U1324 (N_1324,In_482,In_2450);
nor U1325 (N_1325,N_1082,N_1205);
nor U1326 (N_1326,N_572,In_1973);
nor U1327 (N_1327,In_1541,In_995);
xor U1328 (N_1328,N_973,N_987);
nand U1329 (N_1329,N_1212,N_768);
nor U1330 (N_1330,N_295,In_1552);
or U1331 (N_1331,N_816,N_883);
xnor U1332 (N_1332,N_853,N_1144);
or U1333 (N_1333,N_1137,In_1091);
xor U1334 (N_1334,N_657,N_863);
nor U1335 (N_1335,N_899,N_329);
xor U1336 (N_1336,N_434,In_707);
nor U1337 (N_1337,N_5,N_31);
nand U1338 (N_1338,N_353,N_944);
and U1339 (N_1339,In_1532,N_720);
xnor U1340 (N_1340,In_247,N_948);
nor U1341 (N_1341,N_988,N_732);
and U1342 (N_1342,N_1089,N_516);
and U1343 (N_1343,N_661,N_1162);
or U1344 (N_1344,N_1067,N_1075);
xor U1345 (N_1345,N_1111,In_1946);
and U1346 (N_1346,N_759,N_1211);
xnor U1347 (N_1347,In_489,In_447);
or U1348 (N_1348,In_1797,N_1223);
nand U1349 (N_1349,N_1019,N_737);
nand U1350 (N_1350,In_1960,N_700);
xor U1351 (N_1351,In_1556,In_2498);
nor U1352 (N_1352,N_903,N_116);
xnor U1353 (N_1353,N_967,N_1190);
xor U1354 (N_1354,N_664,N_654);
and U1355 (N_1355,N_25,In_2354);
or U1356 (N_1356,N_905,N_740);
nor U1357 (N_1357,In_437,In_38);
xor U1358 (N_1358,In_288,N_1087);
and U1359 (N_1359,In_716,N_678);
nand U1360 (N_1360,N_1218,In_1127);
and U1361 (N_1361,N_940,N_645);
xor U1362 (N_1362,N_241,N_747);
nand U1363 (N_1363,N_1003,N_874);
nand U1364 (N_1364,N_634,N_648);
xor U1365 (N_1365,In_167,N_871);
and U1366 (N_1366,N_1025,N_675);
or U1367 (N_1367,N_628,N_170);
nor U1368 (N_1368,N_343,N_1086);
nand U1369 (N_1369,N_632,N_429);
xnor U1370 (N_1370,N_764,N_1108);
nand U1371 (N_1371,N_66,N_880);
and U1372 (N_1372,In_1620,N_518);
xnor U1373 (N_1373,In_390,N_182);
nor U1374 (N_1374,In_545,In_1146);
xor U1375 (N_1375,In_1954,N_1167);
xnor U1376 (N_1376,N_1110,In_2148);
and U1377 (N_1377,N_886,In_977);
xor U1378 (N_1378,N_1216,N_1198);
nand U1379 (N_1379,N_1084,N_289);
nand U1380 (N_1380,N_848,N_1121);
nor U1381 (N_1381,N_794,In_1087);
xnor U1382 (N_1382,N_714,N_671);
nand U1383 (N_1383,N_919,N_486);
and U1384 (N_1384,In_1060,In_1362);
xor U1385 (N_1385,N_763,N_981);
nor U1386 (N_1386,In_1219,In_442);
xnor U1387 (N_1387,In_755,In_1967);
nor U1388 (N_1388,In_1397,In_2161);
nor U1389 (N_1389,In_1096,N_890);
xnor U1390 (N_1390,In_1656,In_1823);
and U1391 (N_1391,N_808,In_1232);
nand U1392 (N_1392,N_959,N_1160);
nand U1393 (N_1393,N_1145,In_1917);
xnor U1394 (N_1394,N_787,N_1094);
or U1395 (N_1395,N_835,N_626);
nor U1396 (N_1396,N_703,N_293);
and U1397 (N_1397,In_324,N_742);
xor U1398 (N_1398,N_1127,N_746);
nand U1399 (N_1399,N_757,N_302);
or U1400 (N_1400,N_502,N_445);
xor U1401 (N_1401,N_1154,In_2188);
xnor U1402 (N_1402,N_1182,N_1222);
nor U1403 (N_1403,N_1188,N_111);
nor U1404 (N_1404,N_810,N_814);
or U1405 (N_1405,N_766,N_684);
nand U1406 (N_1406,N_13,N_1024);
nand U1407 (N_1407,In_2189,N_138);
nor U1408 (N_1408,N_1043,N_639);
or U1409 (N_1409,N_1196,N_1053);
nand U1410 (N_1410,N_1018,N_1240);
nor U1411 (N_1411,N_698,N_1150);
and U1412 (N_1412,N_1097,N_1022);
nand U1413 (N_1413,N_1191,N_436);
nand U1414 (N_1414,In_830,In_806);
nand U1415 (N_1415,N_1106,In_296);
nand U1416 (N_1416,N_1030,N_386);
nor U1417 (N_1417,N_931,N_1074);
xor U1418 (N_1418,N_912,N_992);
and U1419 (N_1419,N_913,N_581);
nor U1420 (N_1420,In_141,N_844);
or U1421 (N_1421,In_1255,N_1243);
nand U1422 (N_1422,In_922,N_1090);
and U1423 (N_1423,In_1947,In_267);
nor U1424 (N_1424,N_681,N_1079);
or U1425 (N_1425,N_842,N_769);
or U1426 (N_1426,N_238,In_1209);
nand U1427 (N_1427,N_788,N_749);
or U1428 (N_1428,N_834,N_630);
and U1429 (N_1429,N_1159,In_649);
nand U1430 (N_1430,N_633,N_859);
nor U1431 (N_1431,N_356,N_935);
xnor U1432 (N_1432,N_1209,N_216);
or U1433 (N_1433,N_291,In_1026);
and U1434 (N_1434,N_993,In_1892);
nor U1435 (N_1435,In_2257,N_867);
or U1436 (N_1436,In_1801,N_1247);
nand U1437 (N_1437,N_1153,N_17);
nand U1438 (N_1438,N_567,In_1139);
nor U1439 (N_1439,In_1274,N_983);
and U1440 (N_1440,N_647,N_1005);
nand U1441 (N_1441,N_789,N_104);
nor U1442 (N_1442,N_1015,N_1166);
nor U1443 (N_1443,In_377,N_79);
nor U1444 (N_1444,N_923,N_274);
nor U1445 (N_1445,In_2492,In_1490);
or U1446 (N_1446,N_668,N_864);
xnor U1447 (N_1447,In_2224,N_625);
and U1448 (N_1448,N_423,N_811);
nor U1449 (N_1449,N_462,N_144);
nand U1450 (N_1450,In_1095,N_1220);
nand U1451 (N_1451,In_1292,N_722);
nand U1452 (N_1452,In_1487,N_306);
and U1453 (N_1453,N_1073,In_833);
xnor U1454 (N_1454,N_1164,N_807);
or U1455 (N_1455,In_1861,N_1117);
xor U1456 (N_1456,N_211,N_824);
or U1457 (N_1457,N_629,N_1126);
or U1458 (N_1458,In_1606,N_663);
nand U1459 (N_1459,In_2444,N_27);
nand U1460 (N_1460,In_618,N_743);
nor U1461 (N_1461,N_1136,N_801);
and U1462 (N_1462,N_577,N_985);
nor U1463 (N_1463,N_836,N_837);
nor U1464 (N_1464,N_304,N_415);
and U1465 (N_1465,N_230,N_995);
or U1466 (N_1466,N_1229,N_1007);
xor U1467 (N_1467,In_2025,In_413);
or U1468 (N_1468,In_1572,In_2247);
and U1469 (N_1469,N_1221,N_830);
xnor U1470 (N_1470,N_1058,N_1062);
and U1471 (N_1471,In_2046,N_826);
xor U1472 (N_1472,N_659,N_1101);
nor U1473 (N_1473,In_1793,N_786);
or U1474 (N_1474,N_783,In_2349);
nand U1475 (N_1475,In_2069,N_751);
xnor U1476 (N_1476,N_897,In_2240);
or U1477 (N_1477,N_1113,In_1821);
nor U1478 (N_1478,In_428,N_495);
nor U1479 (N_1479,N_873,In_1878);
nor U1480 (N_1480,N_933,In_374);
nand U1481 (N_1481,In_311,N_727);
and U1482 (N_1482,N_1120,N_1189);
and U1483 (N_1483,N_18,N_591);
nor U1484 (N_1484,In_1806,N_1006);
nand U1485 (N_1485,N_908,In_1386);
nor U1486 (N_1486,In_1163,N_849);
or U1487 (N_1487,N_1204,N_1026);
nor U1488 (N_1488,N_711,In_965);
nor U1489 (N_1489,N_1131,N_679);
or U1490 (N_1490,In_185,N_870);
xor U1491 (N_1491,In_1977,N_367);
and U1492 (N_1492,N_780,N_1152);
and U1493 (N_1493,In_2167,N_1230);
nor U1494 (N_1494,N_898,N_78);
nor U1495 (N_1495,In_614,N_653);
nor U1496 (N_1496,N_696,In_1010);
or U1497 (N_1497,In_1374,N_1207);
nor U1498 (N_1498,In_2329,N_444);
and U1499 (N_1499,N_728,In_2020);
and U1500 (N_1500,N_311,N_234);
xor U1501 (N_1501,In_1323,In_1545);
or U1502 (N_1502,N_843,N_45);
nor U1503 (N_1503,N_468,N_1095);
and U1504 (N_1504,In_1157,N_470);
nand U1505 (N_1505,N_1195,N_896);
and U1506 (N_1506,N_481,N_706);
nand U1507 (N_1507,In_468,In_2178);
xnor U1508 (N_1508,In_42,N_878);
xor U1509 (N_1509,In_642,N_1203);
xor U1510 (N_1510,N_379,N_915);
or U1511 (N_1511,N_1201,N_683);
xnor U1512 (N_1512,N_1200,In_2353);
or U1513 (N_1513,In_1200,N_1235);
nor U1514 (N_1514,In_404,In_260);
nand U1515 (N_1515,In_2280,In_782);
xor U1516 (N_1516,N_669,N_868);
or U1517 (N_1517,N_909,In_2440);
or U1518 (N_1518,N_850,N_889);
nand U1519 (N_1519,In_368,N_858);
or U1520 (N_1520,In_2245,In_2317);
or U1521 (N_1521,N_1050,N_1107);
or U1522 (N_1522,In_917,N_392);
and U1523 (N_1523,In_105,N_1093);
nor U1524 (N_1524,N_1096,N_1004);
and U1525 (N_1525,N_1047,N_642);
nand U1526 (N_1526,In_2089,In_585);
or U1527 (N_1527,In_802,N_739);
or U1528 (N_1528,N_1231,In_1165);
xor U1529 (N_1529,N_555,N_1040);
or U1530 (N_1530,N_1192,In_1484);
or U1531 (N_1531,N_1168,N_962);
xor U1532 (N_1532,In_736,In_2045);
nand U1533 (N_1533,In_1896,N_975);
and U1534 (N_1534,N_1178,N_1105);
xor U1535 (N_1535,N_707,In_1956);
nand U1536 (N_1536,N_65,N_998);
and U1537 (N_1537,N_1070,In_332);
and U1538 (N_1538,N_375,N_882);
nor U1539 (N_1539,In_279,In_1783);
xor U1540 (N_1540,N_724,In_1542);
nand U1541 (N_1541,N_1173,In_275);
nand U1542 (N_1542,N_721,N_968);
or U1543 (N_1543,In_1735,In_392);
xnor U1544 (N_1544,N_800,N_734);
nand U1545 (N_1545,N_795,N_1199);
and U1546 (N_1546,N_761,N_828);
and U1547 (N_1547,In_2212,N_618);
nor U1548 (N_1548,In_398,N_974);
nor U1549 (N_1549,N_1147,In_923);
nor U1550 (N_1550,In_1142,N_803);
xnor U1551 (N_1551,N_1214,N_1175);
or U1552 (N_1552,In_630,N_1194);
nor U1553 (N_1553,N_1029,In_2009);
and U1554 (N_1554,In_1566,N_561);
nand U1555 (N_1555,N_282,N_777);
or U1556 (N_1556,N_1129,In_2011);
and U1557 (N_1557,In_880,N_705);
nand U1558 (N_1558,In_1134,In_481);
nand U1559 (N_1559,In_2066,N_1066);
and U1560 (N_1560,N_148,In_487);
and U1561 (N_1561,In_1733,N_688);
nor U1562 (N_1562,N_2,N_70);
xnor U1563 (N_1563,N_164,N_1083);
nand U1564 (N_1564,N_821,N_1128);
nor U1565 (N_1565,N_1143,N_911);
xor U1566 (N_1566,N_744,N_1009);
or U1567 (N_1567,N_838,N_791);
and U1568 (N_1568,N_178,N_1055);
xor U1569 (N_1569,N_340,N_822);
xnor U1570 (N_1570,In_1189,In_1140);
nand U1571 (N_1571,In_328,In_2078);
xnor U1572 (N_1572,N_1034,In_1075);
xnor U1573 (N_1573,N_527,In_2231);
nand U1574 (N_1574,N_930,N_64);
and U1575 (N_1575,N_627,N_695);
and U1576 (N_1576,N_1100,N_475);
xnor U1577 (N_1577,N_1045,In_417);
or U1578 (N_1578,In_609,N_922);
or U1579 (N_1579,N_941,N_805);
and U1580 (N_1580,In_1239,N_427);
xnor U1581 (N_1581,N_1187,N_1014);
nor U1582 (N_1582,N_368,N_996);
nor U1583 (N_1583,N_1169,N_1068);
or U1584 (N_1584,N_508,N_955);
and U1585 (N_1585,N_616,N_852);
xor U1586 (N_1586,N_1072,N_812);
and U1587 (N_1587,N_550,N_692);
or U1588 (N_1588,N_980,N_907);
or U1589 (N_1589,In_2152,N_1132);
and U1590 (N_1590,N_946,N_1010);
xnor U1591 (N_1591,In_2201,N_455);
and U1592 (N_1592,In_2483,N_430);
xor U1593 (N_1593,N_217,N_969);
and U1594 (N_1594,N_1048,N_594);
or U1595 (N_1595,N_243,In_1789);
nor U1596 (N_1596,N_825,In_2406);
nor U1597 (N_1597,N_622,In_2439);
nand U1598 (N_1598,N_1133,N_666);
xor U1599 (N_1599,In_416,N_1049);
and U1600 (N_1600,In_709,N_965);
or U1601 (N_1601,In_298,N_493);
xnor U1602 (N_1602,In_1235,In_83);
xor U1603 (N_1603,N_1210,N_963);
xnor U1604 (N_1604,N_773,N_799);
nand U1605 (N_1605,N_1081,N_1033);
and U1606 (N_1606,In_2126,N_964);
or U1607 (N_1607,N_638,N_640);
or U1608 (N_1608,N_1246,N_1098);
and U1609 (N_1609,In_184,N_943);
or U1610 (N_1610,In_2263,N_1124);
nor U1611 (N_1611,N_991,N_1011);
and U1612 (N_1612,In_1957,N_1044);
nor U1613 (N_1613,N_644,N_37);
nor U1614 (N_1614,N_797,N_623);
nand U1615 (N_1615,N_142,N_872);
xor U1616 (N_1616,N_465,N_1102);
and U1617 (N_1617,In_1138,N_771);
nor U1618 (N_1618,In_1526,N_662);
nand U1619 (N_1619,N_1059,In_99);
nor U1620 (N_1620,In_1230,N_832);
nor U1621 (N_1621,In_448,N_779);
or U1622 (N_1622,N_920,N_1115);
or U1623 (N_1623,N_1104,In_1137);
nand U1624 (N_1624,In_575,In_896);
nand U1625 (N_1625,In_2162,In_2159);
and U1626 (N_1626,In_648,N_754);
and U1627 (N_1627,N_1118,N_1065);
and U1628 (N_1628,In_1888,N_1000);
nand U1629 (N_1629,In_2049,N_841);
xnor U1630 (N_1630,In_200,N_1109);
nand U1631 (N_1631,N_994,N_23);
or U1632 (N_1632,N_738,N_932);
nand U1633 (N_1633,N_552,N_1088);
nor U1634 (N_1634,N_936,N_715);
and U1635 (N_1635,N_676,N_986);
nand U1636 (N_1636,N_414,In_559);
nand U1637 (N_1637,N_71,In_844);
xnor U1638 (N_1638,N_1017,N_736);
nor U1639 (N_1639,N_942,In_990);
nor U1640 (N_1640,N_525,N_109);
xnor U1641 (N_1641,N_1202,In_918);
or U1642 (N_1642,N_651,N_1226);
nor U1643 (N_1643,In_2394,N_420);
and U1644 (N_1644,In_2278,N_1023);
nor U1645 (N_1645,In_1693,In_571);
and U1646 (N_1646,N_765,N_997);
xor U1647 (N_1647,In_1260,N_1037);
nor U1648 (N_1648,In_1169,N_1174);
xnor U1649 (N_1649,In_479,N_1028);
xor U1650 (N_1650,N_1078,N_1228);
xnor U1651 (N_1651,In_2461,In_1101);
and U1652 (N_1652,In_761,In_364);
and U1653 (N_1653,In_2056,In_1571);
and U1654 (N_1654,N_33,In_85);
nor U1655 (N_1655,N_277,N_151);
nor U1656 (N_1656,In_2260,In_1152);
or U1657 (N_1657,In_511,In_1609);
nor U1658 (N_1658,In_30,N_699);
xnor U1659 (N_1659,N_586,N_288);
or U1660 (N_1660,In_1772,N_646);
or U1661 (N_1661,In_471,N_957);
nand U1662 (N_1662,In_2366,In_549);
nor U1663 (N_1663,N_1125,N_608);
nand U1664 (N_1664,N_1155,N_793);
nand U1665 (N_1665,N_910,In_1062);
or U1666 (N_1666,N_173,N_717);
nand U1667 (N_1667,N_205,N_57);
nor U1668 (N_1668,N_298,In_1553);
nand U1669 (N_1669,N_1061,N_441);
or U1670 (N_1670,N_175,In_1282);
nor U1671 (N_1671,N_286,In_201);
nand U1672 (N_1672,In_2206,In_903);
xnor U1673 (N_1673,N_1008,N_582);
and U1674 (N_1674,In_1106,In_595);
xnor U1675 (N_1675,In_327,In_1328);
nor U1676 (N_1676,N_1180,In_1557);
nor U1677 (N_1677,N_1197,N_1032);
nand U1678 (N_1678,In_2391,N_884);
nand U1679 (N_1679,In_1608,N_360);
nor U1680 (N_1680,N_73,N_990);
nor U1681 (N_1681,N_831,N_956);
or U1682 (N_1682,N_315,N_96);
and U1683 (N_1683,In_818,In_1476);
nand U1684 (N_1684,N_916,In_227);
xnor U1685 (N_1685,In_2106,In_337);
nor U1686 (N_1686,N_40,N_702);
nor U1687 (N_1687,In_450,N_690);
and U1688 (N_1688,N_1172,N_403);
nand U1689 (N_1689,N_971,In_2102);
nor U1690 (N_1690,In_351,In_1054);
and U1691 (N_1691,In_1851,N_583);
or U1692 (N_1692,N_1122,N_902);
nand U1693 (N_1693,N_636,In_1120);
nand U1694 (N_1694,N_804,In_233);
nand U1695 (N_1695,N_817,N_210);
or U1696 (N_1696,N_1186,In_2117);
xnor U1697 (N_1697,N_1016,In_1777);
and U1698 (N_1698,N_925,In_464);
xor U1699 (N_1699,In_372,N_1181);
nand U1700 (N_1700,In_2399,N_553);
nand U1701 (N_1701,In_248,In_1221);
nand U1702 (N_1702,In_1304,In_747);
or U1703 (N_1703,In_1873,N_56);
and U1704 (N_1704,N_497,N_877);
nand U1705 (N_1705,In_2258,In_2118);
and U1706 (N_1706,N_1056,N_798);
or U1707 (N_1707,N_1225,N_180);
nor U1708 (N_1708,N_1064,N_650);
xor U1709 (N_1709,In_2275,N_1239);
nor U1710 (N_1710,N_394,In_1520);
and U1711 (N_1711,N_726,N_84);
or U1712 (N_1712,N_674,N_989);
or U1713 (N_1713,N_823,N_660);
and U1714 (N_1714,N_172,N_961);
nor U1715 (N_1715,In_1839,In_1578);
or U1716 (N_1716,N_128,N_725);
and U1717 (N_1717,N_526,N_1130);
and U1718 (N_1718,N_774,In_532);
and U1719 (N_1719,In_215,N_364);
or U1720 (N_1720,N_847,N_735);
nand U1721 (N_1721,In_2039,In_1631);
nor U1722 (N_1722,N_680,In_1076);
and U1723 (N_1723,N_718,N_1091);
nand U1724 (N_1724,N_949,In_1452);
or U1725 (N_1725,In_613,In_1115);
and U1726 (N_1726,In_1788,N_854);
or U1727 (N_1727,In_1289,N_656);
or U1728 (N_1728,N_755,N_1119);
nand U1729 (N_1729,N_953,In_503);
or U1730 (N_1730,In_211,N_970);
or U1731 (N_1731,In_473,N_1092);
nand U1732 (N_1732,N_540,N_792);
xor U1733 (N_1733,In_919,N_760);
and U1734 (N_1734,N_772,In_1074);
nand U1735 (N_1735,N_347,In_477);
nor U1736 (N_1736,N_276,N_1248);
or U1737 (N_1737,N_750,N_1063);
and U1738 (N_1738,In_1019,N_782);
nor U1739 (N_1739,In_1378,N_865);
or U1740 (N_1740,In_319,N_716);
or U1741 (N_1741,N_1139,N_982);
nand U1742 (N_1742,N_463,In_800);
nand U1743 (N_1743,N_1163,N_901);
or U1744 (N_1744,N_409,N_686);
or U1745 (N_1745,N_856,N_857);
xnor U1746 (N_1746,N_762,N_697);
or U1747 (N_1747,In_1820,N_813);
or U1748 (N_1748,N_1039,N_845);
nand U1749 (N_1749,N_377,N_1020);
or U1750 (N_1750,N_410,N_820);
nand U1751 (N_1751,N_833,N_32);
nand U1752 (N_1752,In_2402,N_643);
and U1753 (N_1753,In_2343,In_2338);
nand U1754 (N_1754,N_895,N_1245);
xnor U1755 (N_1755,In_1617,N_1099);
nand U1756 (N_1756,In_936,N_1071);
and U1757 (N_1757,N_729,N_918);
and U1758 (N_1758,N_1151,N_1077);
nor U1759 (N_1759,N_1036,In_1391);
or U1760 (N_1760,N_1112,N_914);
nor U1761 (N_1761,In_314,In_626);
and U1762 (N_1762,N_351,In_2312);
nor U1763 (N_1763,N_893,N_255);
and U1764 (N_1764,N_287,In_1599);
nor U1765 (N_1765,In_2433,N_976);
xor U1766 (N_1766,N_767,In_697);
nor U1767 (N_1767,N_827,N_1217);
or U1768 (N_1768,In_41,N_1213);
nor U1769 (N_1769,N_1184,In_1938);
and U1770 (N_1770,N_1149,In_598);
nand U1771 (N_1771,N_1170,N_921);
and U1772 (N_1772,In_2456,N_649);
nand U1773 (N_1773,In_2234,N_927);
xor U1774 (N_1774,N_685,In_1494);
and U1775 (N_1775,In_862,N_514);
or U1776 (N_1776,N_257,In_1022);
or U1777 (N_1777,In_866,N_1208);
nor U1778 (N_1778,In_1834,In_2239);
nand U1779 (N_1779,In_86,N_171);
nor U1780 (N_1780,In_700,N_951);
or U1781 (N_1781,N_770,N_1193);
nand U1782 (N_1782,In_1767,In_2065);
nand U1783 (N_1783,In_1558,N_446);
nand U1784 (N_1784,In_629,N_376);
and U1785 (N_1785,In_1030,N_1244);
nand U1786 (N_1786,In_639,N_1076);
nor U1787 (N_1787,N_542,N_556);
and U1788 (N_1788,N_124,In_1745);
nand U1789 (N_1789,N_136,N_819);
nand U1790 (N_1790,N_840,N_250);
nor U1791 (N_1791,N_881,In_1020);
or U1792 (N_1792,N_259,In_304);
xor U1793 (N_1793,In_2481,N_900);
nand U1794 (N_1794,N_977,In_1934);
nor U1795 (N_1795,In_1857,N_512);
nand U1796 (N_1796,N_595,N_546);
nand U1797 (N_1797,In_1424,N_888);
xor U1798 (N_1798,N_776,N_999);
xor U1799 (N_1799,In_1785,N_934);
and U1800 (N_1800,N_140,In_1876);
xor U1801 (N_1801,N_1185,N_1041);
nor U1802 (N_1802,In_496,In_1989);
nor U1803 (N_1803,N_1103,N_748);
nor U1804 (N_1804,N_200,N_467);
nand U1805 (N_1805,N_972,In_1257);
nor U1806 (N_1806,In_1039,In_657);
and U1807 (N_1807,N_1060,In_115);
and U1808 (N_1808,N_818,N_846);
or U1809 (N_1809,In_188,N_1038);
xnor U1810 (N_1810,N_106,N_373);
xor U1811 (N_1811,In_407,In_895);
nand U1812 (N_1812,N_829,N_1046);
and U1813 (N_1813,N_775,In_333);
xnor U1814 (N_1814,N_1123,N_950);
xnor U1815 (N_1815,In_689,N_1146);
nor U1816 (N_1816,N_1140,N_1021);
or U1817 (N_1817,N_328,In_1194);
nand U1818 (N_1818,N_1224,N_652);
or U1819 (N_1819,N_947,N_673);
or U1820 (N_1820,In_53,N_929);
nor U1821 (N_1821,In_1314,N_354);
nand U1822 (N_1822,In_548,In_2173);
or U1823 (N_1823,N_979,N_1052);
xor U1824 (N_1824,N_723,N_667);
and U1825 (N_1825,N_1138,In_1927);
nand U1826 (N_1826,N_1069,In_1580);
xor U1827 (N_1827,N_624,In_2053);
nor U1828 (N_1828,N_1013,In_2480);
or U1829 (N_1829,N_670,N_1135);
and U1830 (N_1830,N_891,In_1191);
nand U1831 (N_1831,N_665,N_120);
and U1832 (N_1832,N_1141,N_694);
or U1833 (N_1833,N_712,N_892);
xor U1834 (N_1834,N_945,N_731);
and U1835 (N_1835,N_3,N_733);
nor U1836 (N_1836,In_1071,N_1027);
or U1837 (N_1837,In_968,N_887);
nand U1838 (N_1838,In_887,N_419);
xnor U1839 (N_1839,N_704,N_855);
xor U1840 (N_1840,In_0,N_262);
and U1841 (N_1841,N_153,In_1474);
nor U1842 (N_1842,N_952,In_1962);
nand U1843 (N_1843,In_743,N_672);
nand U1844 (N_1844,N_758,N_906);
xnor U1845 (N_1845,In_1683,N_752);
and U1846 (N_1846,N_790,N_876);
or U1847 (N_1847,In_1226,N_90);
nor U1848 (N_1848,N_862,N_869);
nand U1849 (N_1849,N_781,N_265);
xor U1850 (N_1850,N_1085,N_978);
nor U1851 (N_1851,N_1233,N_1215);
nor U1852 (N_1852,N_1165,N_939);
nand U1853 (N_1853,N_958,N_938);
nor U1854 (N_1854,In_2361,N_223);
nor U1855 (N_1855,In_1890,N_1161);
or U1856 (N_1856,In_780,N_1249);
nand U1857 (N_1857,N_926,N_710);
or U1858 (N_1858,In_1694,N_687);
and U1859 (N_1859,N_129,N_1156);
nand U1860 (N_1860,N_917,N_984);
xnor U1861 (N_1861,In_836,N_191);
nor U1862 (N_1862,N_860,N_421);
or U1863 (N_1863,N_691,N_547);
nand U1864 (N_1864,N_954,N_452);
and U1865 (N_1865,In_128,N_924);
and U1866 (N_1866,N_1176,In_506);
or U1867 (N_1867,In_126,N_310);
nor U1868 (N_1868,In_2119,N_960);
nor U1869 (N_1869,N_1206,In_135);
xor U1870 (N_1870,N_1171,N_99);
xnor U1871 (N_1871,In_602,N_682);
xnor U1872 (N_1872,N_1148,In_1724);
nand U1873 (N_1873,N_966,N_349);
or U1874 (N_1874,N_689,N_94);
xnor U1875 (N_1875,N_1643,N_1512);
nand U1876 (N_1876,N_1326,N_1274);
nand U1877 (N_1877,N_1854,N_1595);
nor U1878 (N_1878,N_1437,N_1401);
nor U1879 (N_1879,N_1320,N_1608);
nand U1880 (N_1880,N_1728,N_1584);
nor U1881 (N_1881,N_1478,N_1712);
or U1882 (N_1882,N_1353,N_1558);
and U1883 (N_1883,N_1431,N_1604);
or U1884 (N_1884,N_1698,N_1373);
or U1885 (N_1885,N_1511,N_1335);
or U1886 (N_1886,N_1276,N_1283);
and U1887 (N_1887,N_1311,N_1286);
or U1888 (N_1888,N_1535,N_1695);
and U1889 (N_1889,N_1500,N_1497);
xor U1890 (N_1890,N_1328,N_1746);
nor U1891 (N_1891,N_1683,N_1722);
or U1892 (N_1892,N_1570,N_1831);
nand U1893 (N_1893,N_1263,N_1261);
xnor U1894 (N_1894,N_1765,N_1631);
nor U1895 (N_1895,N_1734,N_1813);
nor U1896 (N_1896,N_1563,N_1441);
nor U1897 (N_1897,N_1573,N_1501);
and U1898 (N_1898,N_1634,N_1407);
nand U1899 (N_1899,N_1545,N_1397);
or U1900 (N_1900,N_1541,N_1638);
nand U1901 (N_1901,N_1438,N_1526);
nor U1902 (N_1902,N_1572,N_1823);
xor U1903 (N_1903,N_1816,N_1290);
and U1904 (N_1904,N_1618,N_1783);
nor U1905 (N_1905,N_1537,N_1465);
nand U1906 (N_1906,N_1650,N_1613);
nor U1907 (N_1907,N_1857,N_1384);
nor U1908 (N_1908,N_1296,N_1705);
nand U1909 (N_1909,N_1257,N_1639);
or U1910 (N_1910,N_1798,N_1349);
nand U1911 (N_1911,N_1282,N_1386);
or U1912 (N_1912,N_1351,N_1801);
or U1913 (N_1913,N_1729,N_1778);
nor U1914 (N_1914,N_1389,N_1534);
or U1915 (N_1915,N_1814,N_1488);
nor U1916 (N_1916,N_1250,N_1533);
xnor U1917 (N_1917,N_1499,N_1292);
nor U1918 (N_1918,N_1498,N_1294);
and U1919 (N_1919,N_1319,N_1315);
nand U1920 (N_1920,N_1701,N_1591);
nand U1921 (N_1921,N_1758,N_1521);
xnor U1922 (N_1922,N_1640,N_1606);
nor U1923 (N_1923,N_1792,N_1756);
xnor U1924 (N_1924,N_1428,N_1614);
or U1925 (N_1925,N_1706,N_1797);
xnor U1926 (N_1926,N_1495,N_1254);
or U1927 (N_1927,N_1291,N_1738);
nor U1928 (N_1928,N_1285,N_1770);
xor U1929 (N_1929,N_1364,N_1543);
and U1930 (N_1930,N_1754,N_1416);
nor U1931 (N_1931,N_1777,N_1841);
nand U1932 (N_1932,N_1256,N_1760);
or U1933 (N_1933,N_1630,N_1477);
nand U1934 (N_1934,N_1549,N_1339);
xnor U1935 (N_1935,N_1755,N_1560);
and U1936 (N_1936,N_1779,N_1836);
nor U1937 (N_1937,N_1494,N_1647);
xnor U1938 (N_1938,N_1628,N_1413);
xor U1939 (N_1939,N_1776,N_1480);
nand U1940 (N_1940,N_1767,N_1782);
nand U1941 (N_1941,N_1828,N_1253);
nor U1942 (N_1942,N_1661,N_1696);
nor U1943 (N_1943,N_1289,N_1310);
and U1944 (N_1944,N_1505,N_1751);
or U1945 (N_1945,N_1268,N_1700);
nand U1946 (N_1946,N_1725,N_1307);
and U1947 (N_1947,N_1835,N_1868);
nor U1948 (N_1948,N_1300,N_1626);
xnor U1949 (N_1949,N_1418,N_1405);
and U1950 (N_1950,N_1660,N_1432);
xor U1951 (N_1951,N_1496,N_1623);
nand U1952 (N_1952,N_1516,N_1708);
xnor U1953 (N_1953,N_1561,N_1580);
or U1954 (N_1954,N_1843,N_1436);
and U1955 (N_1955,N_1255,N_1852);
nand U1956 (N_1956,N_1669,N_1596);
nor U1957 (N_1957,N_1601,N_1317);
and U1958 (N_1958,N_1745,N_1404);
and U1959 (N_1959,N_1637,N_1800);
nor U1960 (N_1960,N_1483,N_1342);
nand U1961 (N_1961,N_1636,N_1298);
or U1962 (N_1962,N_1818,N_1527);
nand U1963 (N_1963,N_1301,N_1513);
and U1964 (N_1964,N_1362,N_1517);
and U1965 (N_1965,N_1375,N_1713);
xnor U1966 (N_1966,N_1620,N_1544);
nor U1967 (N_1967,N_1277,N_1665);
xnor U1968 (N_1968,N_1863,N_1808);
or U1969 (N_1969,N_1581,N_1272);
or U1970 (N_1970,N_1279,N_1382);
xor U1971 (N_1971,N_1302,N_1810);
and U1972 (N_1972,N_1491,N_1312);
xnor U1973 (N_1973,N_1592,N_1670);
xnor U1974 (N_1974,N_1262,N_1468);
nand U1975 (N_1975,N_1367,N_1554);
nor U1976 (N_1976,N_1548,N_1588);
nand U1977 (N_1977,N_1391,N_1484);
or U1978 (N_1978,N_1528,N_1809);
nor U1979 (N_1979,N_1786,N_1451);
and U1980 (N_1980,N_1430,N_1486);
nor U1981 (N_1981,N_1550,N_1330);
and U1982 (N_1982,N_1532,N_1733);
nor U1983 (N_1983,N_1392,N_1834);
xnor U1984 (N_1984,N_1470,N_1602);
and U1985 (N_1985,N_1671,N_1506);
nor U1986 (N_1986,N_1799,N_1474);
nor U1987 (N_1987,N_1720,N_1742);
nand U1988 (N_1988,N_1819,N_1444);
or U1989 (N_1989,N_1743,N_1795);
and U1990 (N_1990,N_1771,N_1714);
and U1991 (N_1991,N_1363,N_1802);
nor U1992 (N_1992,N_1749,N_1764);
and U1993 (N_1993,N_1410,N_1514);
nand U1994 (N_1994,N_1675,N_1856);
nand U1995 (N_1995,N_1690,N_1775);
or U1996 (N_1996,N_1615,N_1622);
nor U1997 (N_1997,N_1555,N_1260);
nor U1998 (N_1998,N_1252,N_1653);
xnor U1999 (N_1999,N_1585,N_1370);
xor U2000 (N_2000,N_1414,N_1378);
xor U2001 (N_2001,N_1308,N_1523);
nand U2002 (N_2002,N_1865,N_1387);
and U2003 (N_2003,N_1399,N_1656);
and U2004 (N_2004,N_1377,N_1569);
and U2005 (N_2005,N_1632,N_1763);
xnor U2006 (N_2006,N_1594,N_1425);
xor U2007 (N_2007,N_1462,N_1735);
or U2008 (N_2008,N_1772,N_1693);
xor U2009 (N_2009,N_1603,N_1736);
nor U2010 (N_2010,N_1582,N_1440);
xnor U2011 (N_2011,N_1723,N_1846);
nand U2012 (N_2012,N_1599,N_1519);
xor U2013 (N_2013,N_1361,N_1492);
nor U2014 (N_2014,N_1668,N_1753);
nor U2015 (N_2015,N_1691,N_1458);
nor U2016 (N_2016,N_1536,N_1443);
nand U2017 (N_2017,N_1476,N_1452);
or U2018 (N_2018,N_1464,N_1824);
xnor U2019 (N_2019,N_1385,N_1258);
nor U2020 (N_2020,N_1565,N_1542);
or U2021 (N_2021,N_1578,N_1641);
nor U2022 (N_2022,N_1627,N_1531);
nand U2023 (N_2023,N_1482,N_1791);
or U2024 (N_2024,N_1586,N_1408);
nor U2025 (N_2025,N_1293,N_1461);
and U2026 (N_2026,N_1858,N_1787);
nand U2027 (N_2027,N_1702,N_1270);
and U2028 (N_2028,N_1332,N_1793);
or U2029 (N_2029,N_1420,N_1619);
and U2030 (N_2030,N_1388,N_1336);
and U2031 (N_2031,N_1266,N_1510);
nand U2032 (N_2032,N_1804,N_1768);
and U2033 (N_2033,N_1780,N_1356);
and U2034 (N_2034,N_1340,N_1807);
nor U2035 (N_2035,N_1860,N_1400);
and U2036 (N_2036,N_1822,N_1744);
nand U2037 (N_2037,N_1681,N_1316);
or U2038 (N_2038,N_1844,N_1825);
and U2039 (N_2039,N_1612,N_1659);
xor U2040 (N_2040,N_1562,N_1366);
nor U2041 (N_2041,N_1402,N_1663);
or U2042 (N_2042,N_1333,N_1493);
nand U2043 (N_2043,N_1815,N_1740);
xnor U2044 (N_2044,N_1717,N_1845);
nor U2045 (N_2045,N_1396,N_1520);
xnor U2046 (N_2046,N_1576,N_1394);
or U2047 (N_2047,N_1773,N_1583);
or U2048 (N_2048,N_1721,N_1337);
nand U2049 (N_2049,N_1832,N_1789);
nand U2050 (N_2050,N_1321,N_1314);
or U2051 (N_2051,N_1538,N_1557);
and U2052 (N_2052,N_1442,N_1571);
nor U2053 (N_2053,N_1748,N_1467);
or U2054 (N_2054,N_1371,N_1785);
nor U2055 (N_2055,N_1323,N_1871);
nand U2056 (N_2056,N_1324,N_1463);
and U2057 (N_2057,N_1861,N_1633);
nor U2058 (N_2058,N_1796,N_1654);
or U2059 (N_2059,N_1485,N_1624);
xnor U2060 (N_2060,N_1350,N_1655);
or U2061 (N_2061,N_1426,N_1699);
or U2062 (N_2062,N_1524,N_1649);
nand U2063 (N_2063,N_1446,N_1556);
nor U2064 (N_2064,N_1454,N_1331);
or U2065 (N_2065,N_1611,N_1271);
nand U2066 (N_2066,N_1811,N_1833);
xnor U2067 (N_2067,N_1509,N_1677);
nand U2068 (N_2068,N_1406,N_1475);
nor U2069 (N_2069,N_1295,N_1727);
xnor U2070 (N_2070,N_1817,N_1334);
xnor U2071 (N_2071,N_1692,N_1429);
or U2072 (N_2072,N_1862,N_1433);
nand U2073 (N_2073,N_1642,N_1435);
or U2074 (N_2074,N_1455,N_1372);
nor U2075 (N_2075,N_1354,N_1439);
nor U2076 (N_2076,N_1840,N_1587);
or U2077 (N_2077,N_1415,N_1716);
nand U2078 (N_2078,N_1348,N_1507);
nor U2079 (N_2079,N_1395,N_1445);
or U2080 (N_2080,N_1593,N_1732);
or U2081 (N_2081,N_1322,N_1515);
or U2082 (N_2082,N_1664,N_1551);
nor U2083 (N_2083,N_1769,N_1566);
or U2084 (N_2084,N_1872,N_1502);
and U2085 (N_2085,N_1667,N_1368);
nor U2086 (N_2086,N_1711,N_1518);
or U2087 (N_2087,N_1374,N_1284);
nor U2088 (N_2088,N_1390,N_1674);
nand U2089 (N_2089,N_1423,N_1837);
nor U2090 (N_2090,N_1530,N_1357);
nand U2091 (N_2091,N_1589,N_1522);
and U2092 (N_2092,N_1381,N_1449);
nor U2093 (N_2093,N_1383,N_1473);
nand U2094 (N_2094,N_1305,N_1447);
nor U2095 (N_2095,N_1376,N_1553);
xor U2096 (N_2096,N_1864,N_1605);
xnor U2097 (N_2097,N_1774,N_1345);
or U2098 (N_2098,N_1529,N_1411);
or U2099 (N_2099,N_1848,N_1424);
xor U2100 (N_2100,N_1259,N_1380);
and U2101 (N_2101,N_1409,N_1684);
and U2102 (N_2102,N_1525,N_1412);
and U2103 (N_2103,N_1434,N_1459);
nand U2104 (N_2104,N_1645,N_1471);
nand U2105 (N_2105,N_1597,N_1457);
or U2106 (N_2106,N_1790,N_1873);
nor U2107 (N_2107,N_1874,N_1299);
or U2108 (N_2108,N_1866,N_1629);
xnor U2109 (N_2109,N_1869,N_1278);
xnor U2110 (N_2110,N_1577,N_1621);
nor U2111 (N_2111,N_1564,N_1646);
or U2112 (N_2112,N_1448,N_1269);
xor U2113 (N_2113,N_1829,N_1341);
nor U2114 (N_2114,N_1821,N_1707);
nand U2115 (N_2115,N_1609,N_1697);
xnor U2116 (N_2116,N_1347,N_1710);
xnor U2117 (N_2117,N_1508,N_1304);
nor U2118 (N_2118,N_1847,N_1610);
nand U2119 (N_2119,N_1762,N_1552);
xnor U2120 (N_2120,N_1379,N_1489);
nand U2121 (N_2121,N_1687,N_1781);
or U2122 (N_2122,N_1546,N_1346);
or U2123 (N_2123,N_1369,N_1838);
xor U2124 (N_2124,N_1460,N_1682);
nor U2125 (N_2125,N_1466,N_1427);
xor U2126 (N_2126,N_1867,N_1805);
and U2127 (N_2127,N_1422,N_1303);
nand U2128 (N_2128,N_1694,N_1704);
nor U2129 (N_2129,N_1287,N_1617);
xnor U2130 (N_2130,N_1598,N_1355);
nor U2131 (N_2131,N_1839,N_1718);
nand U2132 (N_2132,N_1715,N_1766);
nor U2133 (N_2133,N_1827,N_1672);
and U2134 (N_2134,N_1559,N_1393);
nor U2135 (N_2135,N_1851,N_1803);
and U2136 (N_2136,N_1306,N_1365);
or U2137 (N_2137,N_1607,N_1421);
or U2138 (N_2138,N_1352,N_1741);
and U2139 (N_2139,N_1281,N_1820);
xor U2140 (N_2140,N_1757,N_1579);
nand U2141 (N_2141,N_1657,N_1686);
nand U2142 (N_2142,N_1726,N_1739);
nor U2143 (N_2143,N_1855,N_1338);
nor U2144 (N_2144,N_1747,N_1275);
and U2145 (N_2145,N_1806,N_1265);
or U2146 (N_2146,N_1842,N_1788);
or U2147 (N_2147,N_1759,N_1719);
and U2148 (N_2148,N_1327,N_1651);
or U2149 (N_2149,N_1264,N_1648);
and U2150 (N_2150,N_1658,N_1644);
nor U2151 (N_2151,N_1625,N_1490);
and U2152 (N_2152,N_1450,N_1547);
nor U2153 (N_2153,N_1329,N_1666);
and U2154 (N_2154,N_1652,N_1360);
xnor U2155 (N_2155,N_1859,N_1456);
xor U2156 (N_2156,N_1812,N_1794);
and U2157 (N_2157,N_1600,N_1403);
xor U2158 (N_2158,N_1419,N_1318);
nor U2159 (N_2159,N_1685,N_1678);
xor U2160 (N_2160,N_1343,N_1730);
and U2161 (N_2161,N_1830,N_1731);
nand U2162 (N_2162,N_1709,N_1679);
nor U2163 (N_2163,N_1761,N_1568);
nand U2164 (N_2164,N_1280,N_1689);
nor U2165 (N_2165,N_1297,N_1481);
xor U2166 (N_2166,N_1662,N_1479);
nor U2167 (N_2167,N_1737,N_1309);
nand U2168 (N_2168,N_1487,N_1574);
and U2169 (N_2169,N_1469,N_1826);
xnor U2170 (N_2170,N_1540,N_1358);
or U2171 (N_2171,N_1359,N_1503);
or U2172 (N_2172,N_1313,N_1251);
nand U2173 (N_2173,N_1344,N_1575);
nor U2174 (N_2174,N_1673,N_1590);
or U2175 (N_2175,N_1273,N_1504);
and U2176 (N_2176,N_1850,N_1567);
nor U2177 (N_2177,N_1688,N_1676);
xor U2178 (N_2178,N_1267,N_1703);
and U2179 (N_2179,N_1453,N_1417);
nand U2180 (N_2180,N_1853,N_1752);
nand U2181 (N_2181,N_1870,N_1724);
nor U2182 (N_2182,N_1398,N_1750);
nor U2183 (N_2183,N_1616,N_1288);
and U2184 (N_2184,N_1635,N_1784);
nand U2185 (N_2185,N_1325,N_1849);
nor U2186 (N_2186,N_1680,N_1472);
nor U2187 (N_2187,N_1539,N_1657);
nor U2188 (N_2188,N_1446,N_1575);
or U2189 (N_2189,N_1488,N_1279);
and U2190 (N_2190,N_1512,N_1628);
xor U2191 (N_2191,N_1581,N_1374);
xnor U2192 (N_2192,N_1449,N_1389);
nor U2193 (N_2193,N_1672,N_1783);
nand U2194 (N_2194,N_1804,N_1252);
nor U2195 (N_2195,N_1388,N_1275);
nand U2196 (N_2196,N_1587,N_1440);
or U2197 (N_2197,N_1775,N_1375);
nand U2198 (N_2198,N_1547,N_1812);
and U2199 (N_2199,N_1527,N_1736);
nand U2200 (N_2200,N_1545,N_1858);
xor U2201 (N_2201,N_1305,N_1310);
xnor U2202 (N_2202,N_1507,N_1772);
nor U2203 (N_2203,N_1853,N_1571);
nand U2204 (N_2204,N_1801,N_1707);
nor U2205 (N_2205,N_1575,N_1612);
nand U2206 (N_2206,N_1685,N_1339);
nor U2207 (N_2207,N_1708,N_1810);
and U2208 (N_2208,N_1320,N_1742);
nor U2209 (N_2209,N_1648,N_1655);
or U2210 (N_2210,N_1453,N_1813);
nor U2211 (N_2211,N_1398,N_1290);
xnor U2212 (N_2212,N_1559,N_1762);
and U2213 (N_2213,N_1648,N_1307);
nand U2214 (N_2214,N_1320,N_1522);
xnor U2215 (N_2215,N_1583,N_1693);
or U2216 (N_2216,N_1616,N_1373);
nand U2217 (N_2217,N_1329,N_1324);
xnor U2218 (N_2218,N_1799,N_1281);
nor U2219 (N_2219,N_1832,N_1753);
or U2220 (N_2220,N_1806,N_1766);
or U2221 (N_2221,N_1464,N_1420);
xnor U2222 (N_2222,N_1860,N_1585);
nor U2223 (N_2223,N_1266,N_1781);
xnor U2224 (N_2224,N_1323,N_1705);
or U2225 (N_2225,N_1864,N_1696);
nor U2226 (N_2226,N_1811,N_1842);
or U2227 (N_2227,N_1255,N_1762);
xnor U2228 (N_2228,N_1652,N_1420);
or U2229 (N_2229,N_1449,N_1742);
and U2230 (N_2230,N_1689,N_1652);
and U2231 (N_2231,N_1672,N_1344);
or U2232 (N_2232,N_1307,N_1813);
xor U2233 (N_2233,N_1266,N_1441);
nand U2234 (N_2234,N_1515,N_1393);
or U2235 (N_2235,N_1710,N_1601);
or U2236 (N_2236,N_1438,N_1588);
xnor U2237 (N_2237,N_1528,N_1537);
and U2238 (N_2238,N_1504,N_1533);
or U2239 (N_2239,N_1345,N_1718);
or U2240 (N_2240,N_1808,N_1414);
and U2241 (N_2241,N_1595,N_1314);
and U2242 (N_2242,N_1443,N_1660);
xor U2243 (N_2243,N_1806,N_1567);
and U2244 (N_2244,N_1508,N_1868);
nor U2245 (N_2245,N_1739,N_1757);
and U2246 (N_2246,N_1716,N_1403);
nand U2247 (N_2247,N_1601,N_1459);
nor U2248 (N_2248,N_1637,N_1703);
nand U2249 (N_2249,N_1274,N_1273);
nor U2250 (N_2250,N_1857,N_1763);
and U2251 (N_2251,N_1487,N_1288);
nand U2252 (N_2252,N_1403,N_1374);
nand U2253 (N_2253,N_1819,N_1541);
xor U2254 (N_2254,N_1520,N_1338);
or U2255 (N_2255,N_1410,N_1449);
nor U2256 (N_2256,N_1437,N_1593);
and U2257 (N_2257,N_1632,N_1257);
nor U2258 (N_2258,N_1379,N_1791);
xnor U2259 (N_2259,N_1853,N_1495);
and U2260 (N_2260,N_1331,N_1846);
xnor U2261 (N_2261,N_1399,N_1512);
and U2262 (N_2262,N_1426,N_1681);
nand U2263 (N_2263,N_1259,N_1554);
nor U2264 (N_2264,N_1429,N_1263);
or U2265 (N_2265,N_1734,N_1729);
nand U2266 (N_2266,N_1735,N_1488);
or U2267 (N_2267,N_1416,N_1575);
xnor U2268 (N_2268,N_1794,N_1786);
xor U2269 (N_2269,N_1393,N_1448);
nor U2270 (N_2270,N_1332,N_1401);
nor U2271 (N_2271,N_1336,N_1311);
nor U2272 (N_2272,N_1776,N_1792);
xor U2273 (N_2273,N_1707,N_1450);
nor U2274 (N_2274,N_1251,N_1258);
xor U2275 (N_2275,N_1689,N_1866);
or U2276 (N_2276,N_1406,N_1527);
xor U2277 (N_2277,N_1463,N_1437);
xor U2278 (N_2278,N_1398,N_1543);
nand U2279 (N_2279,N_1266,N_1515);
nand U2280 (N_2280,N_1501,N_1660);
nor U2281 (N_2281,N_1643,N_1802);
nand U2282 (N_2282,N_1752,N_1410);
and U2283 (N_2283,N_1608,N_1821);
and U2284 (N_2284,N_1857,N_1362);
xor U2285 (N_2285,N_1825,N_1841);
nor U2286 (N_2286,N_1514,N_1447);
nor U2287 (N_2287,N_1443,N_1487);
xnor U2288 (N_2288,N_1726,N_1347);
xor U2289 (N_2289,N_1502,N_1602);
nand U2290 (N_2290,N_1609,N_1631);
and U2291 (N_2291,N_1831,N_1592);
and U2292 (N_2292,N_1613,N_1424);
nand U2293 (N_2293,N_1555,N_1421);
or U2294 (N_2294,N_1461,N_1668);
or U2295 (N_2295,N_1397,N_1322);
or U2296 (N_2296,N_1522,N_1861);
xnor U2297 (N_2297,N_1811,N_1707);
or U2298 (N_2298,N_1677,N_1344);
nor U2299 (N_2299,N_1322,N_1301);
nor U2300 (N_2300,N_1468,N_1744);
nand U2301 (N_2301,N_1606,N_1669);
and U2302 (N_2302,N_1754,N_1773);
nor U2303 (N_2303,N_1811,N_1315);
nand U2304 (N_2304,N_1287,N_1827);
and U2305 (N_2305,N_1337,N_1777);
and U2306 (N_2306,N_1844,N_1659);
nor U2307 (N_2307,N_1452,N_1411);
or U2308 (N_2308,N_1650,N_1671);
and U2309 (N_2309,N_1280,N_1291);
nand U2310 (N_2310,N_1454,N_1321);
nor U2311 (N_2311,N_1406,N_1795);
nor U2312 (N_2312,N_1355,N_1836);
nor U2313 (N_2313,N_1317,N_1261);
xor U2314 (N_2314,N_1485,N_1478);
and U2315 (N_2315,N_1311,N_1738);
xnor U2316 (N_2316,N_1287,N_1575);
and U2317 (N_2317,N_1366,N_1431);
nand U2318 (N_2318,N_1787,N_1278);
xnor U2319 (N_2319,N_1467,N_1347);
or U2320 (N_2320,N_1476,N_1731);
and U2321 (N_2321,N_1763,N_1481);
xor U2322 (N_2322,N_1428,N_1691);
xor U2323 (N_2323,N_1485,N_1554);
xor U2324 (N_2324,N_1662,N_1577);
xnor U2325 (N_2325,N_1716,N_1397);
nor U2326 (N_2326,N_1781,N_1412);
xor U2327 (N_2327,N_1620,N_1538);
and U2328 (N_2328,N_1707,N_1584);
nor U2329 (N_2329,N_1650,N_1494);
and U2330 (N_2330,N_1366,N_1794);
xor U2331 (N_2331,N_1687,N_1577);
nor U2332 (N_2332,N_1772,N_1735);
nor U2333 (N_2333,N_1652,N_1786);
nand U2334 (N_2334,N_1420,N_1485);
nand U2335 (N_2335,N_1372,N_1869);
xnor U2336 (N_2336,N_1642,N_1834);
nand U2337 (N_2337,N_1598,N_1361);
nor U2338 (N_2338,N_1837,N_1612);
nand U2339 (N_2339,N_1443,N_1516);
and U2340 (N_2340,N_1857,N_1593);
or U2341 (N_2341,N_1294,N_1633);
or U2342 (N_2342,N_1284,N_1293);
and U2343 (N_2343,N_1453,N_1427);
xnor U2344 (N_2344,N_1532,N_1456);
nand U2345 (N_2345,N_1563,N_1743);
or U2346 (N_2346,N_1341,N_1527);
xnor U2347 (N_2347,N_1865,N_1662);
nor U2348 (N_2348,N_1812,N_1323);
nor U2349 (N_2349,N_1492,N_1423);
or U2350 (N_2350,N_1843,N_1654);
xor U2351 (N_2351,N_1684,N_1669);
xnor U2352 (N_2352,N_1499,N_1797);
or U2353 (N_2353,N_1825,N_1254);
or U2354 (N_2354,N_1721,N_1674);
nor U2355 (N_2355,N_1296,N_1854);
and U2356 (N_2356,N_1480,N_1803);
and U2357 (N_2357,N_1337,N_1725);
and U2358 (N_2358,N_1589,N_1796);
and U2359 (N_2359,N_1257,N_1762);
nor U2360 (N_2360,N_1727,N_1654);
and U2361 (N_2361,N_1377,N_1458);
or U2362 (N_2362,N_1352,N_1751);
or U2363 (N_2363,N_1511,N_1438);
nor U2364 (N_2364,N_1514,N_1543);
nand U2365 (N_2365,N_1495,N_1658);
nand U2366 (N_2366,N_1843,N_1278);
nor U2367 (N_2367,N_1625,N_1644);
nand U2368 (N_2368,N_1582,N_1335);
xor U2369 (N_2369,N_1447,N_1569);
and U2370 (N_2370,N_1699,N_1544);
or U2371 (N_2371,N_1289,N_1399);
nor U2372 (N_2372,N_1763,N_1337);
and U2373 (N_2373,N_1456,N_1415);
nand U2374 (N_2374,N_1587,N_1781);
xnor U2375 (N_2375,N_1490,N_1580);
xnor U2376 (N_2376,N_1842,N_1531);
and U2377 (N_2377,N_1541,N_1346);
or U2378 (N_2378,N_1339,N_1668);
and U2379 (N_2379,N_1570,N_1658);
and U2380 (N_2380,N_1581,N_1737);
and U2381 (N_2381,N_1497,N_1361);
and U2382 (N_2382,N_1396,N_1515);
xor U2383 (N_2383,N_1653,N_1352);
nand U2384 (N_2384,N_1628,N_1702);
nor U2385 (N_2385,N_1266,N_1762);
or U2386 (N_2386,N_1863,N_1623);
and U2387 (N_2387,N_1580,N_1390);
and U2388 (N_2388,N_1433,N_1719);
or U2389 (N_2389,N_1621,N_1436);
or U2390 (N_2390,N_1263,N_1671);
xnor U2391 (N_2391,N_1263,N_1439);
or U2392 (N_2392,N_1856,N_1290);
xor U2393 (N_2393,N_1807,N_1697);
nor U2394 (N_2394,N_1517,N_1460);
nor U2395 (N_2395,N_1599,N_1369);
or U2396 (N_2396,N_1299,N_1521);
and U2397 (N_2397,N_1812,N_1307);
nand U2398 (N_2398,N_1455,N_1751);
nor U2399 (N_2399,N_1411,N_1282);
nand U2400 (N_2400,N_1381,N_1445);
xnor U2401 (N_2401,N_1566,N_1496);
and U2402 (N_2402,N_1374,N_1517);
and U2403 (N_2403,N_1698,N_1616);
or U2404 (N_2404,N_1319,N_1484);
nand U2405 (N_2405,N_1787,N_1798);
xor U2406 (N_2406,N_1426,N_1548);
or U2407 (N_2407,N_1819,N_1636);
or U2408 (N_2408,N_1620,N_1608);
xor U2409 (N_2409,N_1611,N_1493);
nand U2410 (N_2410,N_1252,N_1352);
nor U2411 (N_2411,N_1525,N_1610);
nor U2412 (N_2412,N_1764,N_1316);
and U2413 (N_2413,N_1369,N_1788);
or U2414 (N_2414,N_1593,N_1300);
xor U2415 (N_2415,N_1789,N_1494);
nand U2416 (N_2416,N_1378,N_1701);
nor U2417 (N_2417,N_1595,N_1643);
and U2418 (N_2418,N_1837,N_1404);
or U2419 (N_2419,N_1742,N_1271);
and U2420 (N_2420,N_1350,N_1613);
nor U2421 (N_2421,N_1722,N_1787);
nor U2422 (N_2422,N_1446,N_1418);
nor U2423 (N_2423,N_1426,N_1408);
or U2424 (N_2424,N_1682,N_1437);
xnor U2425 (N_2425,N_1601,N_1578);
xnor U2426 (N_2426,N_1494,N_1512);
nand U2427 (N_2427,N_1586,N_1671);
nand U2428 (N_2428,N_1720,N_1405);
and U2429 (N_2429,N_1708,N_1842);
nand U2430 (N_2430,N_1403,N_1553);
and U2431 (N_2431,N_1552,N_1291);
and U2432 (N_2432,N_1641,N_1418);
or U2433 (N_2433,N_1821,N_1571);
xor U2434 (N_2434,N_1782,N_1855);
nand U2435 (N_2435,N_1621,N_1858);
nand U2436 (N_2436,N_1448,N_1701);
xor U2437 (N_2437,N_1812,N_1386);
and U2438 (N_2438,N_1715,N_1405);
nand U2439 (N_2439,N_1788,N_1755);
nand U2440 (N_2440,N_1797,N_1565);
xnor U2441 (N_2441,N_1507,N_1754);
xnor U2442 (N_2442,N_1793,N_1715);
nor U2443 (N_2443,N_1442,N_1787);
and U2444 (N_2444,N_1849,N_1766);
xor U2445 (N_2445,N_1576,N_1332);
nand U2446 (N_2446,N_1821,N_1698);
and U2447 (N_2447,N_1376,N_1543);
and U2448 (N_2448,N_1482,N_1734);
or U2449 (N_2449,N_1280,N_1603);
and U2450 (N_2450,N_1705,N_1599);
nand U2451 (N_2451,N_1825,N_1508);
nand U2452 (N_2452,N_1734,N_1750);
nand U2453 (N_2453,N_1339,N_1696);
nand U2454 (N_2454,N_1810,N_1648);
nand U2455 (N_2455,N_1445,N_1751);
nor U2456 (N_2456,N_1822,N_1325);
nor U2457 (N_2457,N_1388,N_1454);
or U2458 (N_2458,N_1479,N_1501);
xor U2459 (N_2459,N_1743,N_1827);
and U2460 (N_2460,N_1537,N_1444);
and U2461 (N_2461,N_1319,N_1491);
nor U2462 (N_2462,N_1686,N_1549);
nand U2463 (N_2463,N_1833,N_1640);
xor U2464 (N_2464,N_1837,N_1858);
xor U2465 (N_2465,N_1580,N_1301);
xor U2466 (N_2466,N_1287,N_1631);
or U2467 (N_2467,N_1596,N_1600);
or U2468 (N_2468,N_1547,N_1509);
xnor U2469 (N_2469,N_1410,N_1684);
xnor U2470 (N_2470,N_1401,N_1496);
and U2471 (N_2471,N_1303,N_1323);
nand U2472 (N_2472,N_1703,N_1771);
or U2473 (N_2473,N_1313,N_1472);
nor U2474 (N_2474,N_1430,N_1267);
nor U2475 (N_2475,N_1272,N_1804);
nor U2476 (N_2476,N_1323,N_1545);
or U2477 (N_2477,N_1625,N_1694);
nand U2478 (N_2478,N_1276,N_1608);
xnor U2479 (N_2479,N_1334,N_1545);
nor U2480 (N_2480,N_1359,N_1573);
nand U2481 (N_2481,N_1325,N_1622);
or U2482 (N_2482,N_1813,N_1800);
or U2483 (N_2483,N_1642,N_1527);
or U2484 (N_2484,N_1840,N_1640);
xor U2485 (N_2485,N_1428,N_1300);
or U2486 (N_2486,N_1444,N_1556);
or U2487 (N_2487,N_1715,N_1768);
nand U2488 (N_2488,N_1371,N_1384);
and U2489 (N_2489,N_1325,N_1396);
nor U2490 (N_2490,N_1590,N_1742);
nand U2491 (N_2491,N_1710,N_1653);
or U2492 (N_2492,N_1567,N_1672);
nand U2493 (N_2493,N_1325,N_1511);
xnor U2494 (N_2494,N_1657,N_1421);
xor U2495 (N_2495,N_1612,N_1862);
nor U2496 (N_2496,N_1612,N_1594);
and U2497 (N_2497,N_1639,N_1697);
xnor U2498 (N_2498,N_1325,N_1856);
and U2499 (N_2499,N_1721,N_1298);
nand U2500 (N_2500,N_2469,N_1931);
nand U2501 (N_2501,N_2455,N_2310);
and U2502 (N_2502,N_1911,N_1992);
or U2503 (N_2503,N_1956,N_2397);
xor U2504 (N_2504,N_1950,N_2157);
nor U2505 (N_2505,N_1924,N_1986);
xnor U2506 (N_2506,N_2279,N_1894);
nor U2507 (N_2507,N_2419,N_2468);
nor U2508 (N_2508,N_2359,N_2206);
and U2509 (N_2509,N_2319,N_2124);
nand U2510 (N_2510,N_1905,N_2480);
xnor U2511 (N_2511,N_2196,N_2345);
nand U2512 (N_2512,N_2172,N_2130);
xnor U2513 (N_2513,N_2213,N_2381);
xnor U2514 (N_2514,N_2485,N_2143);
and U2515 (N_2515,N_2005,N_1975);
xor U2516 (N_2516,N_2446,N_2047);
or U2517 (N_2517,N_2395,N_2431);
or U2518 (N_2518,N_2233,N_2287);
nor U2519 (N_2519,N_2202,N_2475);
nand U2520 (N_2520,N_2409,N_2448);
nand U2521 (N_2521,N_2371,N_2439);
and U2522 (N_2522,N_2356,N_1970);
xor U2523 (N_2523,N_2094,N_2030);
nor U2524 (N_2524,N_2014,N_1916);
and U2525 (N_2525,N_2365,N_2154);
or U2526 (N_2526,N_2236,N_2134);
nor U2527 (N_2527,N_1968,N_2316);
nor U2528 (N_2528,N_2118,N_2248);
or U2529 (N_2529,N_2331,N_2168);
and U2530 (N_2530,N_2243,N_2232);
or U2531 (N_2531,N_1964,N_2360);
and U2532 (N_2532,N_2476,N_1919);
and U2533 (N_2533,N_1935,N_2089);
nand U2534 (N_2534,N_2046,N_2037);
xor U2535 (N_2535,N_2437,N_2065);
xnor U2536 (N_2536,N_2325,N_2499);
nand U2537 (N_2537,N_1980,N_2281);
xnor U2538 (N_2538,N_1988,N_2060);
xnor U2539 (N_2539,N_2497,N_2478);
xnor U2540 (N_2540,N_1929,N_2018);
nor U2541 (N_2541,N_1978,N_2182);
nor U2542 (N_2542,N_2384,N_2408);
nand U2543 (N_2543,N_2225,N_2081);
nand U2544 (N_2544,N_2158,N_1999);
and U2545 (N_2545,N_2457,N_2302);
and U2546 (N_2546,N_1892,N_2488);
xor U2547 (N_2547,N_2412,N_2222);
xor U2548 (N_2548,N_1932,N_1888);
and U2549 (N_2549,N_2283,N_2467);
nand U2550 (N_2550,N_2432,N_2288);
nor U2551 (N_2551,N_2415,N_2038);
nand U2552 (N_2552,N_2271,N_1998);
nor U2553 (N_2553,N_2142,N_2088);
or U2554 (N_2554,N_1943,N_2440);
xor U2555 (N_2555,N_2443,N_2128);
or U2556 (N_2556,N_2436,N_2103);
nor U2557 (N_2557,N_1941,N_2076);
nor U2558 (N_2558,N_2112,N_2194);
xnor U2559 (N_2559,N_2184,N_2390);
and U2560 (N_2560,N_2129,N_2174);
and U2561 (N_2561,N_2035,N_2327);
and U2562 (N_2562,N_2315,N_2460);
and U2563 (N_2563,N_2082,N_2087);
and U2564 (N_2564,N_2256,N_2454);
xnor U2565 (N_2565,N_2337,N_2069);
xor U2566 (N_2566,N_2275,N_2414);
and U2567 (N_2567,N_2246,N_2207);
nand U2568 (N_2568,N_2027,N_2123);
nand U2569 (N_2569,N_2085,N_1966);
nand U2570 (N_2570,N_1938,N_2228);
xor U2571 (N_2571,N_1957,N_2171);
and U2572 (N_2572,N_2219,N_2388);
nand U2573 (N_2573,N_2376,N_2031);
or U2574 (N_2574,N_2297,N_2138);
nor U2575 (N_2575,N_2262,N_2442);
nor U2576 (N_2576,N_2097,N_1948);
nor U2577 (N_2577,N_2276,N_2224);
or U2578 (N_2578,N_2398,N_2355);
xnor U2579 (N_2579,N_2197,N_2402);
and U2580 (N_2580,N_2329,N_2070);
xor U2581 (N_2581,N_2148,N_1936);
nor U2582 (N_2582,N_1912,N_2309);
nand U2583 (N_2583,N_2424,N_2254);
xor U2584 (N_2584,N_2192,N_2349);
xor U2585 (N_2585,N_1944,N_2453);
nand U2586 (N_2586,N_2473,N_1907);
nand U2587 (N_2587,N_2017,N_2020);
xor U2588 (N_2588,N_2176,N_2318);
or U2589 (N_2589,N_2374,N_2111);
nor U2590 (N_2590,N_2472,N_2066);
nand U2591 (N_2591,N_2137,N_2139);
nor U2592 (N_2592,N_2121,N_2255);
xnor U2593 (N_2593,N_2244,N_2106);
and U2594 (N_2594,N_2311,N_2167);
nor U2595 (N_2595,N_1889,N_2152);
nor U2596 (N_2596,N_2144,N_2249);
nand U2597 (N_2597,N_2394,N_2012);
nor U2598 (N_2598,N_2185,N_1979);
xor U2599 (N_2599,N_2377,N_2285);
or U2600 (N_2600,N_2072,N_2362);
nor U2601 (N_2601,N_2320,N_2044);
nor U2602 (N_2602,N_2223,N_2272);
nor U2603 (N_2603,N_2008,N_2486);
nor U2604 (N_2604,N_2164,N_2465);
xor U2605 (N_2605,N_1937,N_2247);
nor U2606 (N_2606,N_2368,N_1977);
and U2607 (N_2607,N_2025,N_2180);
and U2608 (N_2608,N_1883,N_2438);
and U2609 (N_2609,N_2101,N_2253);
or U2610 (N_2610,N_2498,N_2479);
and U2611 (N_2611,N_2383,N_1914);
and U2612 (N_2612,N_2179,N_1906);
xor U2613 (N_2613,N_1878,N_2135);
and U2614 (N_2614,N_2173,N_2334);
and U2615 (N_2615,N_2175,N_2423);
or U2616 (N_2616,N_1927,N_2127);
xor U2617 (N_2617,N_1949,N_2043);
nand U2618 (N_2618,N_2104,N_2265);
nand U2619 (N_2619,N_2369,N_2481);
xor U2620 (N_2620,N_2022,N_2188);
nand U2621 (N_2621,N_2218,N_2096);
nor U2622 (N_2622,N_2002,N_1982);
and U2623 (N_2623,N_2482,N_1960);
nor U2624 (N_2624,N_2463,N_2461);
and U2625 (N_2625,N_2251,N_2338);
xnor U2626 (N_2626,N_2313,N_2039);
or U2627 (N_2627,N_2351,N_2293);
nor U2628 (N_2628,N_1940,N_2492);
nand U2629 (N_2629,N_2308,N_2422);
nand U2630 (N_2630,N_2140,N_1962);
or U2631 (N_2631,N_2161,N_2052);
or U2632 (N_2632,N_1886,N_2100);
nor U2633 (N_2633,N_2084,N_2187);
or U2634 (N_2634,N_2483,N_2322);
nor U2635 (N_2635,N_1947,N_2264);
xnor U2636 (N_2636,N_1922,N_2203);
nand U2637 (N_2637,N_2413,N_2198);
nand U2638 (N_2638,N_2459,N_2263);
nand U2639 (N_2639,N_2462,N_1946);
nor U2640 (N_2640,N_1961,N_2199);
or U2641 (N_2641,N_1995,N_2366);
xor U2642 (N_2642,N_2292,N_2208);
or U2643 (N_2643,N_2056,N_1969);
and U2644 (N_2644,N_2339,N_2058);
and U2645 (N_2645,N_2433,N_2221);
xor U2646 (N_2646,N_2491,N_2274);
nand U2647 (N_2647,N_1879,N_2098);
nand U2648 (N_2648,N_1955,N_2241);
nor U2649 (N_2649,N_1952,N_2163);
or U2650 (N_2650,N_2312,N_2372);
or U2651 (N_2651,N_2450,N_2010);
nor U2652 (N_2652,N_2091,N_2466);
and U2653 (N_2653,N_1959,N_1971);
or U2654 (N_2654,N_2193,N_2386);
xor U2655 (N_2655,N_2231,N_1896);
xor U2656 (N_2656,N_2217,N_2364);
nor U2657 (N_2657,N_2034,N_1910);
and U2658 (N_2658,N_2298,N_2099);
nor U2659 (N_2659,N_1930,N_2400);
nand U2660 (N_2660,N_2132,N_2190);
nor U2661 (N_2661,N_2314,N_2358);
nand U2662 (N_2662,N_1973,N_2237);
and U2663 (N_2663,N_2300,N_1925);
nand U2664 (N_2664,N_2299,N_2280);
and U2665 (N_2665,N_2165,N_2080);
and U2666 (N_2666,N_1920,N_2307);
nor U2667 (N_2667,N_1897,N_2054);
xor U2668 (N_2668,N_2332,N_2363);
and U2669 (N_2669,N_2487,N_1939);
xor U2670 (N_2670,N_2120,N_2107);
nand U2671 (N_2671,N_2278,N_2260);
xor U2672 (N_2672,N_2117,N_2404);
nor U2673 (N_2673,N_2093,N_2456);
nor U2674 (N_2674,N_2258,N_1981);
nand U2675 (N_2675,N_2083,N_1965);
nor U2676 (N_2676,N_2347,N_2162);
nand U2677 (N_2677,N_2346,N_2385);
nor U2678 (N_2678,N_1909,N_1990);
and U2679 (N_2679,N_2133,N_2057);
nor U2680 (N_2680,N_1987,N_2191);
xnor U2681 (N_2681,N_2484,N_2321);
and U2682 (N_2682,N_1885,N_1963);
nand U2683 (N_2683,N_1983,N_2391);
nand U2684 (N_2684,N_2417,N_2382);
xnor U2685 (N_2685,N_2494,N_2477);
nand U2686 (N_2686,N_2426,N_1917);
nand U2687 (N_2687,N_2493,N_2282);
nand U2688 (N_2688,N_2177,N_2421);
nand U2689 (N_2689,N_2048,N_1918);
xor U2690 (N_2690,N_2268,N_2340);
xor U2691 (N_2691,N_2214,N_2013);
xnor U2692 (N_2692,N_2273,N_2040);
xor U2693 (N_2693,N_2301,N_2026);
nor U2694 (N_2694,N_1884,N_2336);
or U2695 (N_2695,N_1903,N_2373);
nor U2696 (N_2696,N_2227,N_2407);
xor U2697 (N_2697,N_2317,N_2335);
or U2698 (N_2698,N_2361,N_2284);
and U2699 (N_2699,N_2250,N_2186);
nand U2700 (N_2700,N_1899,N_2073);
nand U2701 (N_2701,N_2159,N_2141);
nand U2702 (N_2702,N_1900,N_2029);
or U2703 (N_2703,N_2328,N_2153);
xor U2704 (N_2704,N_2016,N_2427);
nand U2705 (N_2705,N_2294,N_1991);
nor U2706 (N_2706,N_2195,N_1984);
xor U2707 (N_2707,N_2036,N_2230);
and U2708 (N_2708,N_2470,N_2201);
nand U2709 (N_2709,N_2090,N_2147);
xor U2710 (N_2710,N_2220,N_1908);
and U2711 (N_2711,N_2053,N_2277);
nand U2712 (N_2712,N_2267,N_1890);
and U2713 (N_2713,N_2049,N_2051);
and U2714 (N_2714,N_2108,N_2126);
nor U2715 (N_2715,N_2032,N_2146);
nor U2716 (N_2716,N_2452,N_1895);
or U2717 (N_2717,N_2403,N_2496);
or U2718 (N_2718,N_2445,N_1934);
xnor U2719 (N_2719,N_2324,N_2149);
and U2720 (N_2720,N_1972,N_1915);
nand U2721 (N_2721,N_1921,N_2114);
xnor U2722 (N_2722,N_2028,N_1875);
nand U2723 (N_2723,N_2155,N_2078);
or U2724 (N_2724,N_2210,N_1913);
and U2725 (N_2725,N_2342,N_2011);
nor U2726 (N_2726,N_2055,N_2489);
or U2727 (N_2727,N_2291,N_2270);
nand U2728 (N_2728,N_2458,N_2102);
nor U2729 (N_2729,N_2357,N_2075);
and U2730 (N_2730,N_2001,N_1898);
and U2731 (N_2731,N_2150,N_2063);
or U2732 (N_2732,N_2405,N_2392);
and U2733 (N_2733,N_2183,N_2068);
or U2734 (N_2734,N_2116,N_2401);
or U2735 (N_2735,N_2399,N_1989);
nand U2736 (N_2736,N_2406,N_2019);
xnor U2737 (N_2737,N_2289,N_2003);
nor U2738 (N_2738,N_2009,N_2136);
or U2739 (N_2739,N_1976,N_2451);
nand U2740 (N_2740,N_2041,N_2259);
xnor U2741 (N_2741,N_1958,N_2326);
nor U2742 (N_2742,N_2434,N_2115);
or U2743 (N_2743,N_2375,N_2189);
or U2744 (N_2744,N_2323,N_2074);
nor U2745 (N_2745,N_2387,N_2023);
nor U2746 (N_2746,N_2435,N_2238);
and U2747 (N_2747,N_2353,N_2425);
or U2748 (N_2748,N_2269,N_1876);
or U2749 (N_2749,N_2064,N_2007);
and U2750 (N_2750,N_1951,N_1933);
and U2751 (N_2751,N_2211,N_2166);
or U2752 (N_2752,N_2092,N_1954);
and U2753 (N_2753,N_2266,N_2042);
nor U2754 (N_2754,N_2416,N_1887);
xor U2755 (N_2755,N_2004,N_2200);
and U2756 (N_2756,N_2204,N_1996);
and U2757 (N_2757,N_1904,N_2113);
nand U2758 (N_2758,N_2086,N_1967);
or U2759 (N_2759,N_2242,N_2050);
or U2760 (N_2760,N_2252,N_2215);
xor U2761 (N_2761,N_2062,N_2370);
nor U2762 (N_2762,N_2354,N_1891);
or U2763 (N_2763,N_2024,N_2061);
xnor U2764 (N_2764,N_2464,N_1997);
xor U2765 (N_2765,N_2333,N_2348);
xnor U2766 (N_2766,N_2109,N_1974);
or U2767 (N_2767,N_2000,N_1926);
or U2768 (N_2768,N_2170,N_1985);
nor U2769 (N_2769,N_2380,N_2067);
xnor U2770 (N_2770,N_2160,N_2430);
and U2771 (N_2771,N_2105,N_2306);
nor U2772 (N_2772,N_2261,N_1923);
or U2773 (N_2773,N_1901,N_2420);
xnor U2774 (N_2774,N_2212,N_2131);
and U2775 (N_2775,N_2235,N_2240);
nand U2776 (N_2776,N_2330,N_2305);
xnor U2777 (N_2777,N_2303,N_1994);
xnor U2778 (N_2778,N_1880,N_2110);
nand U2779 (N_2779,N_2418,N_2156);
xor U2780 (N_2780,N_2033,N_2045);
or U2781 (N_2781,N_2389,N_1928);
and U2782 (N_2782,N_2059,N_2006);
nand U2783 (N_2783,N_2378,N_2344);
nand U2784 (N_2784,N_2145,N_2396);
or U2785 (N_2785,N_2245,N_2447);
and U2786 (N_2786,N_2239,N_2015);
nor U2787 (N_2787,N_2226,N_2471);
and U2788 (N_2788,N_2411,N_2304);
xnor U2789 (N_2789,N_2341,N_2393);
or U2790 (N_2790,N_2444,N_1945);
nand U2791 (N_2791,N_1902,N_2352);
nor U2792 (N_2792,N_2474,N_2169);
nor U2793 (N_2793,N_2125,N_2286);
and U2794 (N_2794,N_2071,N_1877);
nand U2795 (N_2795,N_2449,N_2428);
xor U2796 (N_2796,N_2410,N_1893);
nor U2797 (N_2797,N_2216,N_2379);
xnor U2798 (N_2798,N_1953,N_2021);
and U2799 (N_2799,N_2095,N_1942);
xor U2800 (N_2800,N_2151,N_2077);
or U2801 (N_2801,N_2367,N_2343);
and U2802 (N_2802,N_1993,N_2257);
xnor U2803 (N_2803,N_2350,N_2495);
xnor U2804 (N_2804,N_2122,N_2119);
nand U2805 (N_2805,N_2429,N_2181);
nor U2806 (N_2806,N_2295,N_2296);
and U2807 (N_2807,N_2234,N_1882);
nor U2808 (N_2808,N_2079,N_2178);
nor U2809 (N_2809,N_2290,N_2441);
xor U2810 (N_2810,N_2209,N_2205);
nand U2811 (N_2811,N_2229,N_1881);
xor U2812 (N_2812,N_2490,N_2106);
nor U2813 (N_2813,N_2205,N_1985);
or U2814 (N_2814,N_1928,N_2179);
or U2815 (N_2815,N_2368,N_2397);
xor U2816 (N_2816,N_1971,N_2243);
nand U2817 (N_2817,N_1982,N_2221);
nand U2818 (N_2818,N_2119,N_2261);
and U2819 (N_2819,N_1930,N_2164);
and U2820 (N_2820,N_2187,N_2089);
and U2821 (N_2821,N_2228,N_1961);
and U2822 (N_2822,N_2001,N_2145);
and U2823 (N_2823,N_1952,N_2073);
or U2824 (N_2824,N_1940,N_2482);
nor U2825 (N_2825,N_2055,N_2311);
or U2826 (N_2826,N_2009,N_2377);
and U2827 (N_2827,N_1989,N_2393);
xnor U2828 (N_2828,N_2011,N_2286);
nand U2829 (N_2829,N_2422,N_2419);
or U2830 (N_2830,N_1954,N_2135);
or U2831 (N_2831,N_2021,N_2062);
nor U2832 (N_2832,N_2062,N_2083);
and U2833 (N_2833,N_2368,N_2334);
and U2834 (N_2834,N_2187,N_2459);
nor U2835 (N_2835,N_2477,N_1886);
or U2836 (N_2836,N_2286,N_1881);
or U2837 (N_2837,N_2318,N_2138);
or U2838 (N_2838,N_2216,N_1888);
and U2839 (N_2839,N_2349,N_1958);
and U2840 (N_2840,N_2038,N_2270);
xor U2841 (N_2841,N_2049,N_2181);
nand U2842 (N_2842,N_2257,N_1981);
nor U2843 (N_2843,N_2011,N_1887);
or U2844 (N_2844,N_2321,N_2213);
nor U2845 (N_2845,N_2457,N_1933);
nand U2846 (N_2846,N_1929,N_2214);
nand U2847 (N_2847,N_2287,N_1915);
and U2848 (N_2848,N_2321,N_1950);
or U2849 (N_2849,N_2173,N_1886);
and U2850 (N_2850,N_1951,N_2070);
or U2851 (N_2851,N_2016,N_2041);
and U2852 (N_2852,N_2434,N_2085);
or U2853 (N_2853,N_2180,N_2297);
and U2854 (N_2854,N_2444,N_2183);
nand U2855 (N_2855,N_2188,N_2198);
or U2856 (N_2856,N_2337,N_1883);
nand U2857 (N_2857,N_2232,N_2333);
xor U2858 (N_2858,N_2177,N_2059);
or U2859 (N_2859,N_2149,N_2064);
xnor U2860 (N_2860,N_2318,N_2053);
nor U2861 (N_2861,N_2237,N_1975);
and U2862 (N_2862,N_2477,N_2218);
nor U2863 (N_2863,N_2400,N_2334);
nand U2864 (N_2864,N_2442,N_2114);
and U2865 (N_2865,N_2377,N_2348);
nand U2866 (N_2866,N_1894,N_2119);
nor U2867 (N_2867,N_2347,N_2187);
nor U2868 (N_2868,N_2444,N_2479);
and U2869 (N_2869,N_2422,N_2328);
or U2870 (N_2870,N_2011,N_2007);
xnor U2871 (N_2871,N_2443,N_2101);
xor U2872 (N_2872,N_2317,N_2240);
and U2873 (N_2873,N_2113,N_2259);
nor U2874 (N_2874,N_2003,N_2446);
and U2875 (N_2875,N_2397,N_2205);
nor U2876 (N_2876,N_2142,N_1926);
nand U2877 (N_2877,N_2253,N_1907);
nor U2878 (N_2878,N_2251,N_2442);
or U2879 (N_2879,N_1999,N_2471);
nand U2880 (N_2880,N_2258,N_1965);
nor U2881 (N_2881,N_2019,N_1933);
nand U2882 (N_2882,N_1887,N_2472);
nor U2883 (N_2883,N_2093,N_2415);
xor U2884 (N_2884,N_2481,N_2484);
nor U2885 (N_2885,N_2351,N_2269);
and U2886 (N_2886,N_2460,N_2030);
or U2887 (N_2887,N_2214,N_2153);
nand U2888 (N_2888,N_2124,N_2272);
xor U2889 (N_2889,N_1914,N_2183);
xnor U2890 (N_2890,N_2272,N_2254);
nor U2891 (N_2891,N_2213,N_1884);
nor U2892 (N_2892,N_2068,N_1927);
or U2893 (N_2893,N_2417,N_2327);
xnor U2894 (N_2894,N_2429,N_2239);
xnor U2895 (N_2895,N_2312,N_1884);
or U2896 (N_2896,N_2326,N_2351);
and U2897 (N_2897,N_2172,N_2054);
and U2898 (N_2898,N_1907,N_2155);
nand U2899 (N_2899,N_2106,N_2151);
and U2900 (N_2900,N_2164,N_2120);
nor U2901 (N_2901,N_2420,N_2039);
nand U2902 (N_2902,N_2450,N_2158);
and U2903 (N_2903,N_2203,N_2226);
nor U2904 (N_2904,N_2307,N_2305);
or U2905 (N_2905,N_2070,N_2142);
and U2906 (N_2906,N_2027,N_2395);
nand U2907 (N_2907,N_2204,N_1924);
nor U2908 (N_2908,N_2454,N_2058);
and U2909 (N_2909,N_2045,N_2290);
xnor U2910 (N_2910,N_2099,N_2164);
nor U2911 (N_2911,N_2062,N_2237);
nor U2912 (N_2912,N_2281,N_2085);
xor U2913 (N_2913,N_2048,N_1884);
nand U2914 (N_2914,N_2141,N_2021);
nand U2915 (N_2915,N_1902,N_2291);
xnor U2916 (N_2916,N_2323,N_2247);
nor U2917 (N_2917,N_1909,N_2415);
nor U2918 (N_2918,N_2243,N_2076);
and U2919 (N_2919,N_2318,N_2185);
nand U2920 (N_2920,N_2495,N_2346);
and U2921 (N_2921,N_2170,N_2427);
or U2922 (N_2922,N_1964,N_2486);
and U2923 (N_2923,N_2137,N_1990);
and U2924 (N_2924,N_2320,N_2062);
or U2925 (N_2925,N_2275,N_2091);
or U2926 (N_2926,N_2126,N_2257);
and U2927 (N_2927,N_2427,N_2359);
or U2928 (N_2928,N_2253,N_2285);
nor U2929 (N_2929,N_2344,N_2367);
xor U2930 (N_2930,N_2244,N_2279);
and U2931 (N_2931,N_2318,N_2449);
and U2932 (N_2932,N_2417,N_2464);
xnor U2933 (N_2933,N_1974,N_2230);
nor U2934 (N_2934,N_2465,N_2202);
and U2935 (N_2935,N_1969,N_2478);
or U2936 (N_2936,N_1902,N_2325);
xnor U2937 (N_2937,N_2170,N_2260);
xnor U2938 (N_2938,N_2301,N_2305);
or U2939 (N_2939,N_2397,N_2219);
xor U2940 (N_2940,N_1953,N_1983);
nor U2941 (N_2941,N_2238,N_2232);
nor U2942 (N_2942,N_1952,N_2078);
xnor U2943 (N_2943,N_2010,N_2303);
and U2944 (N_2944,N_2471,N_2036);
nand U2945 (N_2945,N_2054,N_2007);
nand U2946 (N_2946,N_1914,N_2395);
nor U2947 (N_2947,N_2425,N_2288);
nand U2948 (N_2948,N_2285,N_2035);
xnor U2949 (N_2949,N_2235,N_2315);
and U2950 (N_2950,N_1928,N_2263);
nand U2951 (N_2951,N_2186,N_1934);
nor U2952 (N_2952,N_2399,N_2368);
nor U2953 (N_2953,N_2422,N_2396);
nor U2954 (N_2954,N_2017,N_2351);
nand U2955 (N_2955,N_2458,N_2234);
xor U2956 (N_2956,N_2157,N_2380);
nand U2957 (N_2957,N_1914,N_2066);
or U2958 (N_2958,N_2235,N_2052);
or U2959 (N_2959,N_2463,N_2144);
nand U2960 (N_2960,N_2315,N_2257);
nand U2961 (N_2961,N_2421,N_2120);
nand U2962 (N_2962,N_1937,N_2105);
xnor U2963 (N_2963,N_2213,N_2333);
nand U2964 (N_2964,N_2314,N_2433);
and U2965 (N_2965,N_2151,N_1967);
nor U2966 (N_2966,N_2214,N_2448);
xor U2967 (N_2967,N_2341,N_2421);
and U2968 (N_2968,N_2324,N_2201);
nand U2969 (N_2969,N_2042,N_2475);
or U2970 (N_2970,N_1891,N_2213);
nor U2971 (N_2971,N_2249,N_1914);
or U2972 (N_2972,N_2098,N_2314);
nand U2973 (N_2973,N_1962,N_2095);
and U2974 (N_2974,N_2405,N_2095);
or U2975 (N_2975,N_2105,N_2243);
nand U2976 (N_2976,N_2418,N_2351);
nand U2977 (N_2977,N_2190,N_2316);
nor U2978 (N_2978,N_2436,N_2262);
nor U2979 (N_2979,N_2481,N_2436);
nand U2980 (N_2980,N_2059,N_2382);
nor U2981 (N_2981,N_2048,N_2157);
and U2982 (N_2982,N_2058,N_1926);
or U2983 (N_2983,N_2221,N_2362);
nand U2984 (N_2984,N_2237,N_1965);
or U2985 (N_2985,N_2094,N_2328);
nand U2986 (N_2986,N_1985,N_2334);
xor U2987 (N_2987,N_2296,N_2124);
and U2988 (N_2988,N_1897,N_1947);
and U2989 (N_2989,N_1978,N_1928);
nor U2990 (N_2990,N_2355,N_2280);
or U2991 (N_2991,N_2413,N_2158);
xnor U2992 (N_2992,N_2155,N_2081);
nor U2993 (N_2993,N_2116,N_2150);
or U2994 (N_2994,N_2203,N_2094);
and U2995 (N_2995,N_2290,N_2263);
and U2996 (N_2996,N_2001,N_2449);
nand U2997 (N_2997,N_2065,N_2158);
xor U2998 (N_2998,N_2419,N_2054);
or U2999 (N_2999,N_2153,N_2044);
nor U3000 (N_3000,N_2124,N_2267);
or U3001 (N_3001,N_2344,N_2297);
nor U3002 (N_3002,N_2074,N_2082);
xor U3003 (N_3003,N_2172,N_2413);
nor U3004 (N_3004,N_2093,N_2290);
nor U3005 (N_3005,N_2033,N_2347);
or U3006 (N_3006,N_2123,N_2498);
xor U3007 (N_3007,N_2203,N_1985);
or U3008 (N_3008,N_2267,N_2033);
nand U3009 (N_3009,N_2459,N_2377);
xor U3010 (N_3010,N_2331,N_2228);
nor U3011 (N_3011,N_2010,N_2400);
or U3012 (N_3012,N_2075,N_1924);
and U3013 (N_3013,N_1970,N_1961);
or U3014 (N_3014,N_2206,N_2367);
xnor U3015 (N_3015,N_2362,N_2481);
and U3016 (N_3016,N_2388,N_2165);
or U3017 (N_3017,N_1880,N_2125);
nor U3018 (N_3018,N_2262,N_2267);
and U3019 (N_3019,N_1906,N_2414);
or U3020 (N_3020,N_2165,N_2223);
nand U3021 (N_3021,N_2295,N_2024);
nor U3022 (N_3022,N_2047,N_2201);
nor U3023 (N_3023,N_2219,N_1977);
or U3024 (N_3024,N_2084,N_2481);
nor U3025 (N_3025,N_2313,N_2248);
nand U3026 (N_3026,N_2199,N_2142);
or U3027 (N_3027,N_1993,N_2178);
nor U3028 (N_3028,N_2132,N_1937);
nor U3029 (N_3029,N_2205,N_2088);
xor U3030 (N_3030,N_2134,N_2145);
nor U3031 (N_3031,N_1949,N_2158);
or U3032 (N_3032,N_1969,N_2047);
and U3033 (N_3033,N_2027,N_2409);
nor U3034 (N_3034,N_1975,N_2412);
nand U3035 (N_3035,N_1966,N_2282);
nor U3036 (N_3036,N_2072,N_2112);
and U3037 (N_3037,N_2445,N_1940);
nand U3038 (N_3038,N_2190,N_2476);
or U3039 (N_3039,N_2013,N_1904);
nand U3040 (N_3040,N_2282,N_2022);
xnor U3041 (N_3041,N_2450,N_2335);
and U3042 (N_3042,N_2064,N_2316);
xnor U3043 (N_3043,N_1909,N_2222);
nand U3044 (N_3044,N_2049,N_2000);
or U3045 (N_3045,N_2144,N_1926);
xor U3046 (N_3046,N_1937,N_2060);
or U3047 (N_3047,N_1903,N_2070);
nand U3048 (N_3048,N_1978,N_2399);
or U3049 (N_3049,N_1932,N_1886);
nand U3050 (N_3050,N_1992,N_2165);
xnor U3051 (N_3051,N_2233,N_1952);
or U3052 (N_3052,N_2171,N_2161);
xor U3053 (N_3053,N_2304,N_2349);
nor U3054 (N_3054,N_2435,N_2248);
nor U3055 (N_3055,N_1892,N_1941);
nor U3056 (N_3056,N_2007,N_2403);
or U3057 (N_3057,N_2326,N_1986);
xor U3058 (N_3058,N_2207,N_2378);
nand U3059 (N_3059,N_2132,N_2353);
and U3060 (N_3060,N_2479,N_2429);
nand U3061 (N_3061,N_2085,N_2189);
xor U3062 (N_3062,N_1950,N_2267);
xnor U3063 (N_3063,N_2104,N_2102);
and U3064 (N_3064,N_2341,N_2255);
xnor U3065 (N_3065,N_2295,N_1980);
and U3066 (N_3066,N_2291,N_1878);
nand U3067 (N_3067,N_2128,N_2040);
nand U3068 (N_3068,N_2192,N_2329);
nor U3069 (N_3069,N_2270,N_2315);
xnor U3070 (N_3070,N_2153,N_2482);
nand U3071 (N_3071,N_2061,N_2191);
nand U3072 (N_3072,N_1898,N_2136);
or U3073 (N_3073,N_2465,N_2143);
nand U3074 (N_3074,N_2091,N_2049);
nand U3075 (N_3075,N_2322,N_1879);
or U3076 (N_3076,N_2001,N_2485);
nand U3077 (N_3077,N_2207,N_1999);
xnor U3078 (N_3078,N_2080,N_2499);
or U3079 (N_3079,N_2309,N_2335);
and U3080 (N_3080,N_2254,N_2253);
xnor U3081 (N_3081,N_2378,N_2068);
xnor U3082 (N_3082,N_2446,N_2029);
nor U3083 (N_3083,N_2472,N_2088);
or U3084 (N_3084,N_1905,N_2027);
nor U3085 (N_3085,N_2076,N_2330);
xnor U3086 (N_3086,N_2341,N_2072);
nand U3087 (N_3087,N_2092,N_1978);
and U3088 (N_3088,N_2090,N_2279);
and U3089 (N_3089,N_2372,N_1983);
xnor U3090 (N_3090,N_2145,N_1954);
nand U3091 (N_3091,N_2097,N_1978);
nor U3092 (N_3092,N_2143,N_2285);
or U3093 (N_3093,N_2204,N_1958);
xnor U3094 (N_3094,N_2345,N_2123);
or U3095 (N_3095,N_2050,N_2468);
nand U3096 (N_3096,N_2384,N_1883);
and U3097 (N_3097,N_2133,N_2371);
nor U3098 (N_3098,N_2472,N_2416);
or U3099 (N_3099,N_2461,N_2431);
nor U3100 (N_3100,N_2389,N_2171);
nand U3101 (N_3101,N_2050,N_2175);
or U3102 (N_3102,N_2108,N_2059);
or U3103 (N_3103,N_2087,N_2109);
nand U3104 (N_3104,N_2487,N_1964);
xor U3105 (N_3105,N_2024,N_1965);
or U3106 (N_3106,N_2310,N_2438);
xor U3107 (N_3107,N_1994,N_2161);
or U3108 (N_3108,N_2322,N_1995);
xnor U3109 (N_3109,N_2029,N_2480);
or U3110 (N_3110,N_2033,N_2072);
nor U3111 (N_3111,N_2186,N_2036);
nand U3112 (N_3112,N_2236,N_2274);
or U3113 (N_3113,N_1989,N_2061);
xnor U3114 (N_3114,N_2314,N_2089);
and U3115 (N_3115,N_1882,N_2215);
xor U3116 (N_3116,N_2415,N_2375);
nand U3117 (N_3117,N_2389,N_2437);
nor U3118 (N_3118,N_2184,N_2105);
or U3119 (N_3119,N_1985,N_2122);
nand U3120 (N_3120,N_2321,N_2448);
nand U3121 (N_3121,N_2429,N_1929);
nor U3122 (N_3122,N_1921,N_1905);
or U3123 (N_3123,N_2222,N_2430);
nor U3124 (N_3124,N_1997,N_2236);
xor U3125 (N_3125,N_2942,N_2583);
or U3126 (N_3126,N_2878,N_2670);
and U3127 (N_3127,N_2904,N_2982);
xnor U3128 (N_3128,N_3034,N_2764);
xor U3129 (N_3129,N_3094,N_2943);
nor U3130 (N_3130,N_3003,N_2525);
nand U3131 (N_3131,N_3037,N_2926);
or U3132 (N_3132,N_2588,N_2813);
xor U3133 (N_3133,N_3081,N_2681);
nor U3134 (N_3134,N_3087,N_2558);
and U3135 (N_3135,N_2912,N_3031);
or U3136 (N_3136,N_2628,N_2895);
nand U3137 (N_3137,N_2529,N_2799);
or U3138 (N_3138,N_2717,N_3050);
xnor U3139 (N_3139,N_3123,N_2642);
or U3140 (N_3140,N_2719,N_3108);
or U3141 (N_3141,N_2939,N_2809);
xor U3142 (N_3142,N_3106,N_2644);
nor U3143 (N_3143,N_2528,N_2543);
xnor U3144 (N_3144,N_2826,N_2906);
xnor U3145 (N_3145,N_2564,N_2861);
and U3146 (N_3146,N_2533,N_2579);
nand U3147 (N_3147,N_3075,N_2706);
nand U3148 (N_3148,N_2751,N_2936);
nand U3149 (N_3149,N_3090,N_2811);
nor U3150 (N_3150,N_2696,N_2797);
and U3151 (N_3151,N_2546,N_2842);
nor U3152 (N_3152,N_3020,N_2984);
nand U3153 (N_3153,N_2520,N_3112);
nand U3154 (N_3154,N_2871,N_2777);
nand U3155 (N_3155,N_2885,N_2935);
or U3156 (N_3156,N_2674,N_2651);
nand U3157 (N_3157,N_2973,N_2812);
xor U3158 (N_3158,N_3010,N_2837);
nand U3159 (N_3159,N_3122,N_3083);
and U3160 (N_3160,N_3033,N_2580);
and U3161 (N_3161,N_2896,N_2710);
nor U3162 (N_3162,N_2608,N_2945);
and U3163 (N_3163,N_3100,N_2650);
and U3164 (N_3164,N_2881,N_2568);
and U3165 (N_3165,N_2827,N_2793);
xor U3166 (N_3166,N_2841,N_2947);
xor U3167 (N_3167,N_2677,N_2680);
nand U3168 (N_3168,N_2682,N_2541);
or U3169 (N_3169,N_2991,N_2836);
nand U3170 (N_3170,N_2840,N_2995);
xnor U3171 (N_3171,N_2562,N_2603);
nor U3172 (N_3172,N_2846,N_2925);
xor U3173 (N_3173,N_2513,N_2791);
or U3174 (N_3174,N_2767,N_2998);
nor U3175 (N_3175,N_2788,N_2770);
xor U3176 (N_3176,N_3012,N_2910);
and U3177 (N_3177,N_2693,N_2779);
and U3178 (N_3178,N_2699,N_3016);
nand U3179 (N_3179,N_2613,N_2988);
nand U3180 (N_3180,N_2596,N_2989);
nor U3181 (N_3181,N_2610,N_2909);
nand U3182 (N_3182,N_2818,N_2864);
xnor U3183 (N_3183,N_2928,N_3080);
and U3184 (N_3184,N_2934,N_3096);
nand U3185 (N_3185,N_2759,N_3041);
nor U3186 (N_3186,N_2566,N_2614);
and U3187 (N_3187,N_2560,N_2738);
nor U3188 (N_3188,N_2567,N_2940);
and U3189 (N_3189,N_2550,N_2578);
xnor U3190 (N_3190,N_2659,N_3055);
nand U3191 (N_3191,N_2703,N_2866);
nand U3192 (N_3192,N_2741,N_3085);
nor U3193 (N_3193,N_2522,N_2771);
nand U3194 (N_3194,N_3007,N_2730);
nand U3195 (N_3195,N_2966,N_2704);
nand U3196 (N_3196,N_2949,N_2977);
and U3197 (N_3197,N_2675,N_2637);
nor U3198 (N_3198,N_2593,N_2629);
nand U3199 (N_3199,N_2597,N_2729);
and U3200 (N_3200,N_2581,N_3073);
xnor U3201 (N_3201,N_3089,N_2536);
nand U3202 (N_3202,N_2705,N_2669);
nor U3203 (N_3203,N_2551,N_2559);
nand U3204 (N_3204,N_3004,N_2804);
and U3205 (N_3205,N_2586,N_2643);
and U3206 (N_3206,N_2867,N_2946);
nand U3207 (N_3207,N_3098,N_2880);
nor U3208 (N_3208,N_2691,N_2962);
nor U3209 (N_3209,N_2800,N_2532);
or U3210 (N_3210,N_2807,N_3116);
nand U3211 (N_3211,N_2749,N_2666);
and U3212 (N_3212,N_2531,N_2887);
nand U3213 (N_3213,N_3053,N_3078);
xor U3214 (N_3214,N_2623,N_2523);
nand U3215 (N_3215,N_2662,N_3002);
or U3216 (N_3216,N_2868,N_2555);
nor U3217 (N_3217,N_2517,N_2833);
xnor U3218 (N_3218,N_2930,N_2820);
or U3219 (N_3219,N_2734,N_2714);
or U3220 (N_3220,N_2994,N_2582);
xnor U3221 (N_3221,N_3032,N_2755);
xnor U3222 (N_3222,N_2698,N_3088);
and U3223 (N_3223,N_2711,N_2981);
nand U3224 (N_3224,N_2742,N_2944);
and U3225 (N_3225,N_2997,N_2765);
or U3226 (N_3226,N_3074,N_3052);
xnor U3227 (N_3227,N_2636,N_2803);
nand U3228 (N_3228,N_2671,N_3026);
nand U3229 (N_3229,N_3038,N_2592);
or U3230 (N_3230,N_3024,N_2723);
xor U3231 (N_3231,N_2986,N_2908);
or U3232 (N_3232,N_2632,N_2574);
and U3233 (N_3233,N_2883,N_2594);
and U3234 (N_3234,N_2832,N_3095);
nor U3235 (N_3235,N_2585,N_3093);
nand U3236 (N_3236,N_2905,N_2897);
nor U3237 (N_3237,N_2688,N_2778);
nor U3238 (N_3238,N_2924,N_3115);
xnor U3239 (N_3239,N_2515,N_3027);
or U3240 (N_3240,N_2845,N_2960);
or U3241 (N_3241,N_2958,N_2872);
nor U3242 (N_3242,N_2808,N_2859);
or U3243 (N_3243,N_2860,N_2686);
xor U3244 (N_3244,N_2692,N_2544);
nor U3245 (N_3245,N_2587,N_2709);
and U3246 (N_3246,N_2976,N_2873);
nand U3247 (N_3247,N_2911,N_3029);
xnor U3248 (N_3248,N_3048,N_2781);
nor U3249 (N_3249,N_2655,N_2819);
nor U3250 (N_3250,N_2975,N_2985);
nand U3251 (N_3251,N_2921,N_2509);
nand U3252 (N_3252,N_2622,N_2766);
xnor U3253 (N_3253,N_2702,N_3051);
xor U3254 (N_3254,N_2660,N_2679);
or U3255 (N_3255,N_2572,N_2952);
xnor U3256 (N_3256,N_2856,N_2712);
or U3257 (N_3257,N_2862,N_2565);
xnor U3258 (N_3258,N_3014,N_2922);
nand U3259 (N_3259,N_2891,N_2865);
xnor U3260 (N_3260,N_2948,N_2996);
nor U3261 (N_3261,N_3072,N_2801);
nand U3262 (N_3262,N_2663,N_2898);
nor U3263 (N_3263,N_2545,N_2726);
and U3264 (N_3264,N_2701,N_2621);
nor U3265 (N_3265,N_3069,N_2634);
or U3266 (N_3266,N_2538,N_2589);
and U3267 (N_3267,N_3025,N_3111);
or U3268 (N_3268,N_2967,N_2685);
or U3269 (N_3269,N_2516,N_2571);
or U3270 (N_3270,N_2993,N_2715);
or U3271 (N_3271,N_2504,N_2607);
nand U3272 (N_3272,N_3062,N_2831);
xnor U3273 (N_3273,N_2854,N_2968);
and U3274 (N_3274,N_2851,N_2829);
and U3275 (N_3275,N_2810,N_2640);
and U3276 (N_3276,N_2708,N_3077);
xnor U3277 (N_3277,N_2978,N_2920);
nor U3278 (N_3278,N_2821,N_2591);
nand U3279 (N_3279,N_3102,N_2502);
and U3280 (N_3280,N_2773,N_2815);
and U3281 (N_3281,N_2882,N_2556);
xnor U3282 (N_3282,N_2725,N_2697);
and U3283 (N_3283,N_2599,N_2668);
or U3284 (N_3284,N_2760,N_2903);
nor U3285 (N_3285,N_2894,N_3046);
nand U3286 (N_3286,N_2769,N_3120);
xnor U3287 (N_3287,N_2855,N_2507);
xnor U3288 (N_3288,N_2762,N_3104);
xor U3289 (N_3289,N_2774,N_3114);
or U3290 (N_3290,N_2626,N_3045);
or U3291 (N_3291,N_2847,N_3022);
and U3292 (N_3292,N_2990,N_2511);
and U3293 (N_3293,N_2964,N_2519);
xor U3294 (N_3294,N_3121,N_2694);
nand U3295 (N_3295,N_2870,N_3109);
nor U3296 (N_3296,N_2795,N_2913);
nor U3297 (N_3297,N_3008,N_3097);
nand U3298 (N_3298,N_2956,N_2849);
nand U3299 (N_3299,N_2631,N_2652);
nand U3300 (N_3300,N_2600,N_2825);
xnor U3301 (N_3301,N_2877,N_2569);
xor U3302 (N_3302,N_2616,N_2927);
and U3303 (N_3303,N_3068,N_2595);
nand U3304 (N_3304,N_2573,N_3035);
nor U3305 (N_3305,N_3092,N_2684);
nor U3306 (N_3306,N_2915,N_2929);
nand U3307 (N_3307,N_2957,N_3021);
nor U3308 (N_3308,N_3056,N_3001);
and U3309 (N_3309,N_2879,N_2955);
or U3310 (N_3310,N_2888,N_2748);
nor U3311 (N_3311,N_3047,N_2736);
nand U3312 (N_3312,N_2890,N_3061);
nor U3313 (N_3313,N_2501,N_2850);
xnor U3314 (N_3314,N_2733,N_2953);
nand U3315 (N_3315,N_2718,N_2577);
xor U3316 (N_3316,N_2547,N_2941);
nand U3317 (N_3317,N_2602,N_2654);
or U3318 (N_3318,N_2889,N_3000);
nor U3319 (N_3319,N_3076,N_2739);
nor U3320 (N_3320,N_2979,N_2746);
or U3321 (N_3321,N_2763,N_2615);
and U3322 (N_3322,N_3107,N_2822);
nand U3323 (N_3323,N_2852,N_2548);
or U3324 (N_3324,N_2761,N_2690);
or U3325 (N_3325,N_3049,N_2785);
nor U3326 (N_3326,N_2907,N_2969);
nand U3327 (N_3327,N_3067,N_2999);
or U3328 (N_3328,N_2695,N_3036);
nor U3329 (N_3329,N_2796,N_2775);
nor U3330 (N_3330,N_2720,N_3086);
and U3331 (N_3331,N_3013,N_2752);
nand U3332 (N_3332,N_2747,N_2835);
nor U3333 (N_3333,N_2963,N_2639);
or U3334 (N_3334,N_2641,N_3113);
xor U3335 (N_3335,N_2959,N_2892);
and U3336 (N_3336,N_3009,N_2526);
nand U3337 (N_3337,N_2961,N_3124);
and U3338 (N_3338,N_3043,N_2575);
nor U3339 (N_3339,N_2932,N_2500);
or U3340 (N_3340,N_3101,N_2817);
and U3341 (N_3341,N_2784,N_2731);
or U3342 (N_3342,N_2561,N_2974);
and U3343 (N_3343,N_2687,N_2625);
and U3344 (N_3344,N_3054,N_2902);
nor U3345 (N_3345,N_3006,N_2534);
nand U3346 (N_3346,N_2992,N_2553);
or U3347 (N_3347,N_2848,N_2661);
nand U3348 (N_3348,N_3030,N_2798);
xor U3349 (N_3349,N_3018,N_2917);
and U3350 (N_3350,N_2665,N_2965);
nand U3351 (N_3351,N_2554,N_2814);
or U3352 (N_3352,N_2954,N_2950);
xnor U3353 (N_3353,N_3103,N_2689);
or U3354 (N_3354,N_2732,N_2552);
nand U3355 (N_3355,N_2983,N_2790);
nor U3356 (N_3356,N_3017,N_2647);
xor U3357 (N_3357,N_2789,N_2648);
and U3358 (N_3358,N_2753,N_2539);
nand U3359 (N_3359,N_3105,N_2563);
and U3360 (N_3360,N_2970,N_2786);
or U3361 (N_3361,N_2606,N_3011);
and U3362 (N_3362,N_2653,N_2601);
and U3363 (N_3363,N_2524,N_2782);
and U3364 (N_3364,N_3005,N_3015);
or U3365 (N_3365,N_2938,N_2700);
nand U3366 (N_3366,N_2512,N_3082);
or U3367 (N_3367,N_2875,N_2980);
or U3368 (N_3368,N_2619,N_2540);
nand U3369 (N_3369,N_2658,N_2737);
nor U3370 (N_3370,N_2806,N_3058);
and U3371 (N_3371,N_2824,N_3057);
or U3372 (N_3372,N_2792,N_2838);
or U3373 (N_3373,N_2863,N_2618);
xnor U3374 (N_3374,N_2923,N_2527);
nor U3375 (N_3375,N_2627,N_2728);
and U3376 (N_3376,N_2919,N_2816);
nor U3377 (N_3377,N_2743,N_2617);
or U3378 (N_3378,N_2537,N_2542);
xor U3379 (N_3379,N_2722,N_2933);
xnor U3380 (N_3380,N_3019,N_2972);
nand U3381 (N_3381,N_2857,N_2672);
and U3382 (N_3382,N_3064,N_3099);
nor U3383 (N_3383,N_3118,N_2971);
or U3384 (N_3384,N_2900,N_2758);
or U3385 (N_3385,N_2649,N_2508);
and U3386 (N_3386,N_2570,N_2844);
or U3387 (N_3387,N_2505,N_2635);
and U3388 (N_3388,N_2794,N_3042);
and U3389 (N_3389,N_2611,N_2664);
nor U3390 (N_3390,N_2918,N_2805);
nand U3391 (N_3391,N_2744,N_2787);
xnor U3392 (N_3392,N_2514,N_2901);
nor U3393 (N_3393,N_2612,N_2858);
nand U3394 (N_3394,N_2839,N_2853);
nand U3395 (N_3395,N_3059,N_2884);
or U3396 (N_3396,N_2633,N_2506);
and U3397 (N_3397,N_3119,N_2673);
or U3398 (N_3398,N_2780,N_2823);
nand U3399 (N_3399,N_2750,N_2802);
and U3400 (N_3400,N_2638,N_2735);
nor U3401 (N_3401,N_3091,N_2727);
nor U3402 (N_3402,N_2518,N_3066);
xnor U3403 (N_3403,N_2893,N_2745);
or U3404 (N_3404,N_3040,N_3084);
or U3405 (N_3405,N_2828,N_2768);
or U3406 (N_3406,N_2624,N_2724);
nor U3407 (N_3407,N_3071,N_2605);
and U3408 (N_3408,N_2676,N_2886);
or U3409 (N_3409,N_2713,N_2951);
nand U3410 (N_3410,N_2830,N_3044);
or U3411 (N_3411,N_3023,N_2707);
nor U3412 (N_3412,N_2620,N_2874);
or U3413 (N_3413,N_2754,N_2783);
nor U3414 (N_3414,N_2657,N_2584);
or U3415 (N_3415,N_2646,N_2931);
xnor U3416 (N_3416,N_3028,N_2683);
nor U3417 (N_3417,N_3070,N_2609);
nand U3418 (N_3418,N_2776,N_2590);
or U3419 (N_3419,N_3110,N_3039);
nor U3420 (N_3420,N_2521,N_2645);
nor U3421 (N_3421,N_2899,N_2772);
nor U3422 (N_3422,N_2503,N_2667);
nor U3423 (N_3423,N_2914,N_2843);
nor U3424 (N_3424,N_2510,N_2576);
xor U3425 (N_3425,N_2678,N_2721);
xnor U3426 (N_3426,N_3065,N_2604);
nor U3427 (N_3427,N_2535,N_2598);
or U3428 (N_3428,N_2740,N_2630);
nand U3429 (N_3429,N_2656,N_2557);
and U3430 (N_3430,N_2757,N_2987);
nor U3431 (N_3431,N_3063,N_2756);
or U3432 (N_3432,N_2716,N_2834);
xor U3433 (N_3433,N_2530,N_2937);
or U3434 (N_3434,N_2876,N_2916);
nand U3435 (N_3435,N_3079,N_2869);
and U3436 (N_3436,N_3060,N_3117);
nor U3437 (N_3437,N_2549,N_2908);
nand U3438 (N_3438,N_2918,N_2768);
or U3439 (N_3439,N_2731,N_2986);
and U3440 (N_3440,N_3039,N_2950);
xor U3441 (N_3441,N_2870,N_2714);
xnor U3442 (N_3442,N_2647,N_2878);
xnor U3443 (N_3443,N_3105,N_2547);
nand U3444 (N_3444,N_3077,N_2833);
nor U3445 (N_3445,N_3057,N_2879);
nor U3446 (N_3446,N_2820,N_2868);
and U3447 (N_3447,N_2679,N_2777);
nand U3448 (N_3448,N_2795,N_2800);
nand U3449 (N_3449,N_2567,N_2879);
or U3450 (N_3450,N_2544,N_2542);
nor U3451 (N_3451,N_2632,N_2702);
nand U3452 (N_3452,N_2880,N_2658);
nor U3453 (N_3453,N_2944,N_2580);
xnor U3454 (N_3454,N_2511,N_2539);
xor U3455 (N_3455,N_2703,N_2796);
and U3456 (N_3456,N_2686,N_3120);
and U3457 (N_3457,N_2552,N_3048);
nand U3458 (N_3458,N_3063,N_2647);
nor U3459 (N_3459,N_3054,N_2897);
and U3460 (N_3460,N_2743,N_2932);
or U3461 (N_3461,N_2693,N_3035);
and U3462 (N_3462,N_2853,N_3012);
nor U3463 (N_3463,N_2813,N_2771);
nor U3464 (N_3464,N_2512,N_3088);
nand U3465 (N_3465,N_2532,N_2597);
nor U3466 (N_3466,N_2960,N_2844);
nor U3467 (N_3467,N_2614,N_2946);
nand U3468 (N_3468,N_2921,N_2731);
xor U3469 (N_3469,N_2940,N_2504);
and U3470 (N_3470,N_2798,N_2964);
nor U3471 (N_3471,N_2599,N_2802);
nor U3472 (N_3472,N_3121,N_2500);
and U3473 (N_3473,N_2728,N_2629);
and U3474 (N_3474,N_2886,N_2940);
nand U3475 (N_3475,N_2767,N_3081);
and U3476 (N_3476,N_3051,N_3017);
xor U3477 (N_3477,N_2739,N_2636);
nand U3478 (N_3478,N_2646,N_2690);
xor U3479 (N_3479,N_3054,N_2518);
xnor U3480 (N_3480,N_2886,N_2724);
nand U3481 (N_3481,N_3068,N_2943);
nor U3482 (N_3482,N_2797,N_2654);
or U3483 (N_3483,N_2769,N_2632);
nor U3484 (N_3484,N_2747,N_2917);
nor U3485 (N_3485,N_2951,N_3080);
xor U3486 (N_3486,N_2559,N_2792);
or U3487 (N_3487,N_2793,N_2510);
xnor U3488 (N_3488,N_2877,N_2767);
xor U3489 (N_3489,N_3047,N_2766);
and U3490 (N_3490,N_3123,N_2648);
and U3491 (N_3491,N_2898,N_2748);
and U3492 (N_3492,N_3064,N_2933);
nor U3493 (N_3493,N_3068,N_2532);
nor U3494 (N_3494,N_2840,N_2830);
nand U3495 (N_3495,N_2773,N_2605);
nand U3496 (N_3496,N_2822,N_2975);
xnor U3497 (N_3497,N_2883,N_2740);
nand U3498 (N_3498,N_2642,N_3007);
nor U3499 (N_3499,N_2699,N_3027);
nor U3500 (N_3500,N_2606,N_2768);
or U3501 (N_3501,N_2557,N_2870);
xor U3502 (N_3502,N_2769,N_2782);
xnor U3503 (N_3503,N_2759,N_2632);
or U3504 (N_3504,N_2895,N_3101);
and U3505 (N_3505,N_2728,N_2755);
and U3506 (N_3506,N_2542,N_2539);
xor U3507 (N_3507,N_3070,N_2629);
xor U3508 (N_3508,N_2650,N_2520);
nor U3509 (N_3509,N_2548,N_2661);
and U3510 (N_3510,N_2735,N_2850);
nor U3511 (N_3511,N_2681,N_3069);
nand U3512 (N_3512,N_3082,N_2979);
nor U3513 (N_3513,N_3122,N_3110);
xor U3514 (N_3514,N_2859,N_2597);
xor U3515 (N_3515,N_2537,N_2831);
xnor U3516 (N_3516,N_3103,N_2842);
nor U3517 (N_3517,N_2863,N_2543);
nand U3518 (N_3518,N_2657,N_2601);
xor U3519 (N_3519,N_2875,N_2761);
nand U3520 (N_3520,N_2906,N_2521);
or U3521 (N_3521,N_2622,N_2529);
nor U3522 (N_3522,N_2970,N_2869);
and U3523 (N_3523,N_2793,N_2972);
and U3524 (N_3524,N_3058,N_2924);
and U3525 (N_3525,N_2984,N_2702);
xor U3526 (N_3526,N_2582,N_2770);
nand U3527 (N_3527,N_2665,N_2737);
or U3528 (N_3528,N_2627,N_2695);
and U3529 (N_3529,N_2577,N_2768);
nand U3530 (N_3530,N_2992,N_2875);
nand U3531 (N_3531,N_2896,N_3040);
nor U3532 (N_3532,N_2728,N_3091);
nand U3533 (N_3533,N_2709,N_2881);
xor U3534 (N_3534,N_2936,N_3074);
or U3535 (N_3535,N_2718,N_2728);
nand U3536 (N_3536,N_2702,N_3082);
and U3537 (N_3537,N_2869,N_3102);
nor U3538 (N_3538,N_3040,N_2713);
nor U3539 (N_3539,N_2521,N_2552);
nand U3540 (N_3540,N_3066,N_2523);
or U3541 (N_3541,N_2690,N_3022);
xor U3542 (N_3542,N_3021,N_2528);
nand U3543 (N_3543,N_2975,N_2941);
nor U3544 (N_3544,N_2555,N_3116);
and U3545 (N_3545,N_3119,N_2631);
or U3546 (N_3546,N_2986,N_2710);
and U3547 (N_3547,N_2644,N_2548);
xnor U3548 (N_3548,N_2727,N_2835);
and U3549 (N_3549,N_2524,N_2918);
or U3550 (N_3550,N_2720,N_2994);
xor U3551 (N_3551,N_3083,N_2564);
nor U3552 (N_3552,N_2784,N_2734);
and U3553 (N_3553,N_2901,N_2828);
nor U3554 (N_3554,N_2944,N_2745);
nand U3555 (N_3555,N_2858,N_2522);
xor U3556 (N_3556,N_2855,N_2892);
nand U3557 (N_3557,N_2560,N_2987);
nor U3558 (N_3558,N_2875,N_2982);
nor U3559 (N_3559,N_3030,N_2964);
xnor U3560 (N_3560,N_3109,N_2915);
and U3561 (N_3561,N_2598,N_3112);
nand U3562 (N_3562,N_2623,N_3097);
nand U3563 (N_3563,N_3109,N_3030);
or U3564 (N_3564,N_2611,N_2882);
and U3565 (N_3565,N_2889,N_2809);
nand U3566 (N_3566,N_2866,N_3002);
nor U3567 (N_3567,N_2542,N_3119);
nor U3568 (N_3568,N_2986,N_2911);
or U3569 (N_3569,N_2654,N_2986);
nor U3570 (N_3570,N_3081,N_3072);
and U3571 (N_3571,N_2942,N_2995);
or U3572 (N_3572,N_3068,N_2932);
nand U3573 (N_3573,N_2889,N_2801);
xnor U3574 (N_3574,N_2611,N_2539);
nand U3575 (N_3575,N_2888,N_2805);
and U3576 (N_3576,N_3059,N_2952);
xnor U3577 (N_3577,N_2570,N_2910);
xnor U3578 (N_3578,N_2605,N_2655);
and U3579 (N_3579,N_2970,N_2599);
and U3580 (N_3580,N_3072,N_2564);
and U3581 (N_3581,N_2582,N_3018);
nand U3582 (N_3582,N_2643,N_3102);
xnor U3583 (N_3583,N_2746,N_3078);
nor U3584 (N_3584,N_2905,N_3030);
or U3585 (N_3585,N_2584,N_3075);
nand U3586 (N_3586,N_2845,N_3090);
nor U3587 (N_3587,N_3102,N_2530);
or U3588 (N_3588,N_3109,N_2572);
and U3589 (N_3589,N_2887,N_3023);
or U3590 (N_3590,N_2518,N_3021);
or U3591 (N_3591,N_3103,N_2779);
or U3592 (N_3592,N_2946,N_2607);
xor U3593 (N_3593,N_2534,N_2718);
nand U3594 (N_3594,N_2924,N_2601);
and U3595 (N_3595,N_2641,N_2527);
and U3596 (N_3596,N_2543,N_2536);
or U3597 (N_3597,N_2836,N_2841);
or U3598 (N_3598,N_2970,N_2859);
and U3599 (N_3599,N_2597,N_3100);
and U3600 (N_3600,N_2982,N_3108);
nor U3601 (N_3601,N_2711,N_2600);
xor U3602 (N_3602,N_2857,N_3082);
or U3603 (N_3603,N_2721,N_2927);
nand U3604 (N_3604,N_2617,N_2688);
nand U3605 (N_3605,N_3113,N_2913);
nor U3606 (N_3606,N_2975,N_2775);
xor U3607 (N_3607,N_2565,N_2552);
xnor U3608 (N_3608,N_3109,N_2615);
nor U3609 (N_3609,N_2928,N_2814);
nor U3610 (N_3610,N_2618,N_3110);
nand U3611 (N_3611,N_2793,N_2672);
xnor U3612 (N_3612,N_2743,N_2552);
nand U3613 (N_3613,N_2817,N_3022);
xnor U3614 (N_3614,N_2694,N_2838);
and U3615 (N_3615,N_2870,N_2729);
nor U3616 (N_3616,N_2658,N_2595);
and U3617 (N_3617,N_2738,N_2795);
or U3618 (N_3618,N_2863,N_2636);
or U3619 (N_3619,N_2532,N_2836);
and U3620 (N_3620,N_2782,N_2980);
nor U3621 (N_3621,N_2744,N_3061);
and U3622 (N_3622,N_2849,N_2703);
or U3623 (N_3623,N_2581,N_3061);
xnor U3624 (N_3624,N_2596,N_2892);
and U3625 (N_3625,N_2639,N_2992);
and U3626 (N_3626,N_2591,N_2860);
or U3627 (N_3627,N_2522,N_2606);
and U3628 (N_3628,N_3111,N_3007);
nor U3629 (N_3629,N_2797,N_3076);
nand U3630 (N_3630,N_2839,N_2571);
nand U3631 (N_3631,N_3074,N_2911);
or U3632 (N_3632,N_2611,N_2707);
xnor U3633 (N_3633,N_3086,N_2861);
nor U3634 (N_3634,N_2923,N_2604);
nor U3635 (N_3635,N_2571,N_3000);
xor U3636 (N_3636,N_2521,N_2577);
nand U3637 (N_3637,N_2814,N_2908);
nor U3638 (N_3638,N_3093,N_2731);
xnor U3639 (N_3639,N_2711,N_3122);
xor U3640 (N_3640,N_3124,N_2541);
or U3641 (N_3641,N_2685,N_2819);
nor U3642 (N_3642,N_2901,N_2874);
xnor U3643 (N_3643,N_2799,N_2983);
and U3644 (N_3644,N_2679,N_2974);
xor U3645 (N_3645,N_3041,N_2915);
xor U3646 (N_3646,N_2556,N_3051);
and U3647 (N_3647,N_3077,N_3005);
nor U3648 (N_3648,N_2556,N_2723);
and U3649 (N_3649,N_2576,N_2871);
or U3650 (N_3650,N_3044,N_2501);
and U3651 (N_3651,N_2999,N_2505);
xor U3652 (N_3652,N_2646,N_2563);
nor U3653 (N_3653,N_2570,N_2795);
and U3654 (N_3654,N_2938,N_2732);
or U3655 (N_3655,N_2857,N_2977);
xnor U3656 (N_3656,N_2969,N_3081);
and U3657 (N_3657,N_2791,N_2988);
xnor U3658 (N_3658,N_2819,N_2873);
xor U3659 (N_3659,N_2750,N_2579);
xnor U3660 (N_3660,N_2732,N_2672);
and U3661 (N_3661,N_3101,N_2860);
or U3662 (N_3662,N_3044,N_2533);
nor U3663 (N_3663,N_2908,N_2522);
nand U3664 (N_3664,N_2667,N_2525);
nand U3665 (N_3665,N_2778,N_3031);
xnor U3666 (N_3666,N_2800,N_3025);
and U3667 (N_3667,N_2847,N_3095);
nand U3668 (N_3668,N_3082,N_2666);
or U3669 (N_3669,N_2806,N_3109);
and U3670 (N_3670,N_3067,N_2705);
nand U3671 (N_3671,N_2937,N_2794);
xnor U3672 (N_3672,N_2556,N_2532);
nand U3673 (N_3673,N_2633,N_2848);
nand U3674 (N_3674,N_2751,N_2529);
or U3675 (N_3675,N_2571,N_3099);
and U3676 (N_3676,N_3043,N_2628);
nor U3677 (N_3677,N_3072,N_2631);
and U3678 (N_3678,N_2807,N_3086);
xor U3679 (N_3679,N_2582,N_3082);
nand U3680 (N_3680,N_2733,N_2714);
or U3681 (N_3681,N_2948,N_2589);
and U3682 (N_3682,N_2710,N_3077);
nor U3683 (N_3683,N_3022,N_3048);
or U3684 (N_3684,N_3060,N_2855);
nor U3685 (N_3685,N_2979,N_2981);
nand U3686 (N_3686,N_2852,N_2568);
nand U3687 (N_3687,N_3054,N_2728);
or U3688 (N_3688,N_2591,N_2525);
or U3689 (N_3689,N_2664,N_2546);
xnor U3690 (N_3690,N_2910,N_2611);
nand U3691 (N_3691,N_2960,N_2956);
nand U3692 (N_3692,N_2903,N_2578);
nand U3693 (N_3693,N_3000,N_2719);
or U3694 (N_3694,N_2909,N_2852);
nor U3695 (N_3695,N_2801,N_2596);
nand U3696 (N_3696,N_2648,N_2772);
xor U3697 (N_3697,N_2724,N_3056);
or U3698 (N_3698,N_2611,N_3036);
nand U3699 (N_3699,N_2620,N_3109);
xor U3700 (N_3700,N_3104,N_2520);
or U3701 (N_3701,N_2807,N_2540);
and U3702 (N_3702,N_2585,N_2833);
and U3703 (N_3703,N_2523,N_2809);
xor U3704 (N_3704,N_2794,N_2867);
and U3705 (N_3705,N_2864,N_2719);
and U3706 (N_3706,N_2519,N_2656);
nor U3707 (N_3707,N_2681,N_2996);
nand U3708 (N_3708,N_3071,N_2863);
and U3709 (N_3709,N_2641,N_2686);
nand U3710 (N_3710,N_2736,N_2667);
nor U3711 (N_3711,N_2869,N_3095);
nor U3712 (N_3712,N_2678,N_2736);
xor U3713 (N_3713,N_2709,N_2926);
nand U3714 (N_3714,N_2891,N_2974);
nand U3715 (N_3715,N_2970,N_2540);
or U3716 (N_3716,N_2899,N_2587);
nor U3717 (N_3717,N_3105,N_2760);
nand U3718 (N_3718,N_2652,N_2641);
nand U3719 (N_3719,N_2554,N_2804);
nand U3720 (N_3720,N_2626,N_2920);
nor U3721 (N_3721,N_2679,N_2846);
or U3722 (N_3722,N_3099,N_2988);
nor U3723 (N_3723,N_2924,N_2854);
and U3724 (N_3724,N_2913,N_2586);
and U3725 (N_3725,N_2863,N_2667);
xor U3726 (N_3726,N_2926,N_2683);
nor U3727 (N_3727,N_2717,N_3000);
xor U3728 (N_3728,N_3068,N_2691);
nor U3729 (N_3729,N_2761,N_3019);
nand U3730 (N_3730,N_2721,N_2730);
nor U3731 (N_3731,N_3048,N_2950);
xnor U3732 (N_3732,N_2827,N_2930);
nand U3733 (N_3733,N_2515,N_2648);
nor U3734 (N_3734,N_3120,N_2691);
or U3735 (N_3735,N_2660,N_3107);
nand U3736 (N_3736,N_3022,N_2582);
or U3737 (N_3737,N_3091,N_2990);
xor U3738 (N_3738,N_2597,N_3042);
and U3739 (N_3739,N_2507,N_2571);
nor U3740 (N_3740,N_2791,N_2812);
or U3741 (N_3741,N_2541,N_2597);
or U3742 (N_3742,N_2880,N_2731);
or U3743 (N_3743,N_2885,N_2964);
nor U3744 (N_3744,N_2837,N_2826);
xor U3745 (N_3745,N_2607,N_2833);
nand U3746 (N_3746,N_2583,N_2576);
or U3747 (N_3747,N_2983,N_2884);
nor U3748 (N_3748,N_3015,N_2732);
xor U3749 (N_3749,N_2571,N_2982);
nor U3750 (N_3750,N_3354,N_3664);
xor U3751 (N_3751,N_3374,N_3527);
xor U3752 (N_3752,N_3293,N_3360);
nor U3753 (N_3753,N_3684,N_3460);
xnor U3754 (N_3754,N_3333,N_3157);
nand U3755 (N_3755,N_3602,N_3617);
or U3756 (N_3756,N_3309,N_3324);
nand U3757 (N_3757,N_3660,N_3716);
nor U3758 (N_3758,N_3433,N_3364);
nor U3759 (N_3759,N_3181,N_3745);
or U3760 (N_3760,N_3453,N_3539);
nor U3761 (N_3761,N_3462,N_3225);
nand U3762 (N_3762,N_3553,N_3368);
nand U3763 (N_3763,N_3532,N_3277);
nand U3764 (N_3764,N_3696,N_3521);
xnor U3765 (N_3765,N_3214,N_3694);
and U3766 (N_3766,N_3510,N_3281);
and U3767 (N_3767,N_3409,N_3620);
nor U3768 (N_3768,N_3398,N_3383);
xnor U3769 (N_3769,N_3137,N_3549);
nor U3770 (N_3770,N_3247,N_3240);
nand U3771 (N_3771,N_3683,N_3483);
nand U3772 (N_3772,N_3310,N_3722);
nor U3773 (N_3773,N_3266,N_3494);
xor U3774 (N_3774,N_3540,N_3638);
and U3775 (N_3775,N_3252,N_3139);
and U3776 (N_3776,N_3253,N_3315);
nand U3777 (N_3777,N_3296,N_3711);
nand U3778 (N_3778,N_3245,N_3392);
nor U3779 (N_3779,N_3481,N_3352);
and U3780 (N_3780,N_3529,N_3395);
xor U3781 (N_3781,N_3682,N_3704);
and U3782 (N_3782,N_3659,N_3209);
nor U3783 (N_3783,N_3410,N_3326);
or U3784 (N_3784,N_3407,N_3343);
and U3785 (N_3785,N_3730,N_3278);
xor U3786 (N_3786,N_3350,N_3417);
nand U3787 (N_3787,N_3536,N_3457);
xnor U3788 (N_3788,N_3262,N_3236);
nor U3789 (N_3789,N_3256,N_3150);
and U3790 (N_3790,N_3198,N_3743);
or U3791 (N_3791,N_3622,N_3232);
or U3792 (N_3792,N_3675,N_3268);
or U3793 (N_3793,N_3643,N_3386);
xnor U3794 (N_3794,N_3341,N_3126);
nand U3795 (N_3795,N_3448,N_3261);
nand U3796 (N_3796,N_3474,N_3269);
and U3797 (N_3797,N_3738,N_3393);
nand U3798 (N_3798,N_3188,N_3647);
nor U3799 (N_3799,N_3445,N_3479);
nand U3800 (N_3800,N_3165,N_3348);
xnor U3801 (N_3801,N_3312,N_3329);
xnor U3802 (N_3802,N_3400,N_3351);
nand U3803 (N_3803,N_3744,N_3133);
xor U3804 (N_3804,N_3318,N_3687);
nand U3805 (N_3805,N_3446,N_3132);
or U3806 (N_3806,N_3255,N_3185);
nand U3807 (N_3807,N_3636,N_3424);
nor U3808 (N_3808,N_3534,N_3691);
or U3809 (N_3809,N_3606,N_3178);
nor U3810 (N_3810,N_3612,N_3723);
or U3811 (N_3811,N_3740,N_3584);
nor U3812 (N_3812,N_3512,N_3605);
nand U3813 (N_3813,N_3233,N_3273);
nor U3814 (N_3814,N_3451,N_3444);
and U3815 (N_3815,N_3419,N_3594);
xnor U3816 (N_3816,N_3141,N_3624);
or U3817 (N_3817,N_3355,N_3314);
or U3818 (N_3818,N_3183,N_3611);
and U3819 (N_3819,N_3469,N_3306);
and U3820 (N_3820,N_3241,N_3490);
nor U3821 (N_3821,N_3311,N_3561);
and U3822 (N_3822,N_3390,N_3353);
nor U3823 (N_3823,N_3199,N_3712);
nand U3824 (N_3824,N_3248,N_3412);
or U3825 (N_3825,N_3719,N_3697);
or U3826 (N_3826,N_3372,N_3370);
nand U3827 (N_3827,N_3171,N_3283);
xnor U3828 (N_3828,N_3427,N_3747);
xnor U3829 (N_3829,N_3467,N_3206);
nor U3830 (N_3830,N_3470,N_3681);
xor U3831 (N_3831,N_3628,N_3447);
and U3832 (N_3832,N_3369,N_3208);
xnor U3833 (N_3833,N_3486,N_3357);
and U3834 (N_3834,N_3442,N_3610);
nor U3835 (N_3835,N_3559,N_3142);
nand U3836 (N_3836,N_3576,N_3328);
nor U3837 (N_3837,N_3362,N_3303);
nor U3838 (N_3838,N_3587,N_3173);
xnor U3839 (N_3839,N_3519,N_3589);
xnor U3840 (N_3840,N_3601,N_3406);
and U3841 (N_3841,N_3302,N_3503);
xnor U3842 (N_3842,N_3153,N_3569);
nand U3843 (N_3843,N_3389,N_3493);
or U3844 (N_3844,N_3497,N_3147);
or U3845 (N_3845,N_3169,N_3537);
or U3846 (N_3846,N_3555,N_3662);
or U3847 (N_3847,N_3379,N_3699);
nand U3848 (N_3848,N_3193,N_3487);
or U3849 (N_3849,N_3218,N_3518);
nor U3850 (N_3850,N_3706,N_3251);
and U3851 (N_3851,N_3304,N_3471);
nor U3852 (N_3852,N_3524,N_3522);
nand U3853 (N_3853,N_3238,N_3164);
and U3854 (N_3854,N_3346,N_3648);
nor U3855 (N_3855,N_3551,N_3564);
xnor U3856 (N_3856,N_3441,N_3347);
xnor U3857 (N_3857,N_3151,N_3200);
nand U3858 (N_3858,N_3182,N_3590);
nand U3859 (N_3859,N_3621,N_3531);
or U3860 (N_3860,N_3700,N_3645);
or U3861 (N_3861,N_3223,N_3338);
nor U3862 (N_3862,N_3196,N_3274);
or U3863 (N_3863,N_3655,N_3272);
or U3864 (N_3864,N_3415,N_3135);
nor U3865 (N_3865,N_3689,N_3340);
nor U3866 (N_3866,N_3335,N_3159);
xnor U3867 (N_3867,N_3373,N_3168);
xor U3868 (N_3868,N_3154,N_3408);
or U3869 (N_3869,N_3523,N_3160);
xnor U3870 (N_3870,N_3668,N_3653);
nor U3871 (N_3871,N_3657,N_3246);
xnor U3872 (N_3872,N_3425,N_3418);
and U3873 (N_3873,N_3162,N_3686);
nor U3874 (N_3874,N_3525,N_3317);
and U3875 (N_3875,N_3573,N_3466);
xnor U3876 (N_3876,N_3478,N_3290);
or U3877 (N_3877,N_3737,N_3382);
xor U3878 (N_3878,N_3734,N_3205);
nand U3879 (N_3879,N_3320,N_3714);
and U3880 (N_3880,N_3286,N_3579);
or U3881 (N_3881,N_3607,N_3489);
or U3882 (N_3882,N_3739,N_3721);
nand U3883 (N_3883,N_3207,N_3143);
nor U3884 (N_3884,N_3215,N_3468);
or U3885 (N_3885,N_3513,N_3260);
or U3886 (N_3886,N_3705,N_3749);
and U3887 (N_3887,N_3720,N_3161);
nor U3888 (N_3888,N_3365,N_3330);
and U3889 (N_3889,N_3285,N_3498);
nand U3890 (N_3890,N_3725,N_3562);
nor U3891 (N_3891,N_3152,N_3308);
and U3892 (N_3892,N_3685,N_3270);
nor U3893 (N_3893,N_3222,N_3676);
and U3894 (N_3894,N_3204,N_3574);
and U3895 (N_3895,N_3300,N_3595);
nand U3896 (N_3896,N_3736,N_3158);
xnor U3897 (N_3897,N_3414,N_3170);
and U3898 (N_3898,N_3332,N_3615);
nand U3899 (N_3899,N_3630,N_3511);
nand U3900 (N_3900,N_3640,N_3224);
and U3901 (N_3901,N_3291,N_3440);
xnor U3902 (N_3902,N_3432,N_3276);
and U3903 (N_3903,N_3184,N_3550);
xor U3904 (N_3904,N_3526,N_3197);
nand U3905 (N_3905,N_3592,N_3375);
or U3906 (N_3906,N_3136,N_3491);
xor U3907 (N_3907,N_3666,N_3138);
and U3908 (N_3908,N_3288,N_3642);
or U3909 (N_3909,N_3201,N_3456);
and U3910 (N_3910,N_3651,N_3325);
nor U3911 (N_3911,N_3430,N_3639);
and U3912 (N_3912,N_3547,N_3641);
and U3913 (N_3913,N_3267,N_3264);
and U3914 (N_3914,N_3148,N_3342);
and U3915 (N_3915,N_3508,N_3517);
and U3916 (N_3916,N_3577,N_3431);
xor U3917 (N_3917,N_3708,N_3502);
xnor U3918 (N_3918,N_3438,N_3401);
xnor U3919 (N_3919,N_3565,N_3179);
xnor U3920 (N_3920,N_3226,N_3128);
and U3921 (N_3921,N_3604,N_3163);
and U3922 (N_3922,N_3321,N_3724);
nand U3923 (N_3923,N_3598,N_3717);
nand U3924 (N_3924,N_3581,N_3718);
xnor U3925 (N_3925,N_3131,N_3463);
or U3926 (N_3926,N_3495,N_3626);
xnor U3927 (N_3927,N_3403,N_3596);
nand U3928 (N_3928,N_3671,N_3336);
or U3929 (N_3929,N_3216,N_3625);
xor U3930 (N_3930,N_3572,N_3608);
xor U3931 (N_3931,N_3381,N_3242);
xor U3932 (N_3932,N_3220,N_3635);
or U3933 (N_3933,N_3297,N_3501);
or U3934 (N_3934,N_3385,N_3388);
nand U3935 (N_3935,N_3649,N_3287);
and U3936 (N_3936,N_3371,N_3695);
or U3937 (N_3937,N_3437,N_3146);
and U3938 (N_3938,N_3130,N_3500);
or U3939 (N_3939,N_3454,N_3213);
and U3940 (N_3940,N_3480,N_3726);
xor U3941 (N_3941,N_3710,N_3217);
xnor U3942 (N_3942,N_3413,N_3533);
and U3943 (N_3943,N_3542,N_3603);
nand U3944 (N_3944,N_3563,N_3570);
nor U3945 (N_3945,N_3593,N_3709);
and U3946 (N_3946,N_3690,N_3436);
and U3947 (N_3947,N_3679,N_3727);
nand U3948 (N_3948,N_3609,N_3450);
xnor U3949 (N_3949,N_3464,N_3192);
xnor U3950 (N_3950,N_3244,N_3439);
and U3951 (N_3951,N_3212,N_3673);
xor U3952 (N_3952,N_3656,N_3546);
xnor U3953 (N_3953,N_3259,N_3271);
nor U3954 (N_3954,N_3235,N_3391);
and U3955 (N_3955,N_3299,N_3583);
nand U3956 (N_3956,N_3195,N_3482);
xor U3957 (N_3957,N_3384,N_3477);
or U3958 (N_3958,N_3586,N_3472);
nor U3959 (N_3959,N_3399,N_3499);
xnor U3960 (N_3960,N_3249,N_3211);
nor U3961 (N_3961,N_3644,N_3558);
nor U3962 (N_3962,N_3688,N_3254);
xnor U3963 (N_3963,N_3616,N_3396);
or U3964 (N_3964,N_3597,N_3361);
xnor U3965 (N_3965,N_3530,N_3221);
nor U3966 (N_3966,N_3229,N_3337);
or U3967 (N_3967,N_3528,N_3461);
nor U3968 (N_3968,N_3557,N_3514);
and U3969 (N_3969,N_3571,N_3327);
xor U3970 (N_3970,N_3378,N_3515);
nor U3971 (N_3971,N_3632,N_3672);
nand U3972 (N_3972,N_3202,N_3307);
xnor U3973 (N_3973,N_3359,N_3701);
xnor U3974 (N_3974,N_3715,N_3421);
nand U3975 (N_3975,N_3506,N_3358);
nand U3976 (N_3976,N_3728,N_3313);
xor U3977 (N_3977,N_3322,N_3544);
or U3978 (N_3978,N_3543,N_3582);
nor U3979 (N_3979,N_3167,N_3634);
nor U3980 (N_3980,N_3567,N_3652);
xnor U3981 (N_3981,N_3416,N_3674);
and U3982 (N_3982,N_3219,N_3646);
and U3983 (N_3983,N_3692,N_3619);
nor U3984 (N_3984,N_3397,N_3301);
xnor U3985 (N_3985,N_3591,N_3250);
and U3986 (N_3986,N_3339,N_3505);
nand U3987 (N_3987,N_3144,N_3552);
nor U3988 (N_3988,N_3733,N_3742);
nor U3989 (N_3989,N_3134,N_3258);
nor U3990 (N_3990,N_3227,N_3713);
and U3991 (N_3991,N_3560,N_3230);
or U3992 (N_3992,N_3344,N_3585);
and U3993 (N_3993,N_3485,N_3180);
and U3994 (N_3994,N_3488,N_3658);
nor U3995 (N_3995,N_3239,N_3509);
nor U3996 (N_3996,N_3580,N_3746);
nor U3997 (N_3997,N_3669,N_3387);
nor U3998 (N_3998,N_3228,N_3554);
or U3999 (N_3999,N_3145,N_3156);
or U4000 (N_4000,N_3732,N_3190);
nand U4001 (N_4001,N_3556,N_3423);
nor U4002 (N_4002,N_3284,N_3404);
and U4003 (N_4003,N_3535,N_3275);
xnor U4004 (N_4004,N_3588,N_3172);
xor U4005 (N_4005,N_3661,N_3748);
xor U4006 (N_4006,N_3279,N_3599);
xor U4007 (N_4007,N_3678,N_3234);
nor U4008 (N_4008,N_3394,N_3443);
nor U4009 (N_4009,N_3166,N_3367);
nor U4010 (N_4010,N_3475,N_3363);
nor U4011 (N_4011,N_3140,N_3566);
nor U4012 (N_4012,N_3578,N_3422);
and U4013 (N_4013,N_3177,N_3289);
or U4014 (N_4014,N_3376,N_3627);
xor U4015 (N_4015,N_3243,N_3449);
or U4016 (N_4016,N_3623,N_3613);
xor U4017 (N_4017,N_3176,N_3520);
and U4018 (N_4018,N_3575,N_3538);
or U4019 (N_4019,N_3263,N_3316);
and U4020 (N_4020,N_3319,N_3231);
xnor U4021 (N_4021,N_3629,N_3633);
xor U4022 (N_4022,N_3345,N_3476);
nand U4023 (N_4023,N_3465,N_3402);
or U4024 (N_4024,N_3189,N_3237);
xor U4025 (N_4025,N_3420,N_3637);
nand U4026 (N_4026,N_3155,N_3175);
xnor U4027 (N_4027,N_3735,N_3707);
nor U4028 (N_4028,N_3292,N_3366);
or U4029 (N_4029,N_3257,N_3294);
xor U4030 (N_4030,N_3452,N_3129);
and U4031 (N_4031,N_3149,N_3265);
and U4032 (N_4032,N_3295,N_3693);
nor U4033 (N_4033,N_3174,N_3496);
and U4034 (N_4034,N_3654,N_3731);
nor U4035 (N_4035,N_3548,N_3473);
and U4036 (N_4036,N_3282,N_3545);
or U4037 (N_4037,N_3186,N_3323);
xor U4038 (N_4038,N_3677,N_3729);
or U4039 (N_4039,N_3492,N_3614);
or U4040 (N_4040,N_3428,N_3298);
xnor U4041 (N_4041,N_3349,N_3210);
or U4042 (N_4042,N_3680,N_3665);
xor U4043 (N_4043,N_3334,N_3426);
or U4044 (N_4044,N_3663,N_3702);
xor U4045 (N_4045,N_3356,N_3458);
or U4046 (N_4046,N_3568,N_3405);
and U4047 (N_4047,N_3305,N_3127);
xnor U4048 (N_4048,N_3484,N_3631);
xor U4049 (N_4049,N_3667,N_3429);
xnor U4050 (N_4050,N_3411,N_3455);
nor U4051 (N_4051,N_3203,N_3125);
and U4052 (N_4052,N_3741,N_3618);
nand U4053 (N_4053,N_3435,N_3504);
nor U4054 (N_4054,N_3703,N_3670);
and U4055 (N_4055,N_3600,N_3280);
or U4056 (N_4056,N_3541,N_3650);
or U4057 (N_4057,N_3331,N_3459);
xnor U4058 (N_4058,N_3191,N_3434);
or U4059 (N_4059,N_3516,N_3698);
and U4060 (N_4060,N_3194,N_3380);
xnor U4061 (N_4061,N_3507,N_3187);
or U4062 (N_4062,N_3377,N_3148);
nand U4063 (N_4063,N_3126,N_3526);
xor U4064 (N_4064,N_3573,N_3315);
nor U4065 (N_4065,N_3186,N_3212);
and U4066 (N_4066,N_3141,N_3359);
nor U4067 (N_4067,N_3433,N_3220);
nand U4068 (N_4068,N_3152,N_3335);
and U4069 (N_4069,N_3248,N_3488);
xor U4070 (N_4070,N_3304,N_3731);
and U4071 (N_4071,N_3136,N_3389);
nor U4072 (N_4072,N_3743,N_3461);
nor U4073 (N_4073,N_3594,N_3324);
nand U4074 (N_4074,N_3617,N_3648);
or U4075 (N_4075,N_3308,N_3551);
nand U4076 (N_4076,N_3584,N_3665);
and U4077 (N_4077,N_3679,N_3577);
or U4078 (N_4078,N_3583,N_3145);
nand U4079 (N_4079,N_3211,N_3727);
nand U4080 (N_4080,N_3604,N_3627);
xnor U4081 (N_4081,N_3322,N_3377);
and U4082 (N_4082,N_3354,N_3287);
xor U4083 (N_4083,N_3592,N_3593);
or U4084 (N_4084,N_3700,N_3339);
nand U4085 (N_4085,N_3219,N_3356);
nand U4086 (N_4086,N_3503,N_3229);
nand U4087 (N_4087,N_3480,N_3196);
xnor U4088 (N_4088,N_3270,N_3514);
nand U4089 (N_4089,N_3690,N_3552);
nand U4090 (N_4090,N_3586,N_3329);
nor U4091 (N_4091,N_3664,N_3592);
nor U4092 (N_4092,N_3263,N_3264);
and U4093 (N_4093,N_3443,N_3209);
nor U4094 (N_4094,N_3277,N_3643);
and U4095 (N_4095,N_3648,N_3135);
xor U4096 (N_4096,N_3591,N_3630);
and U4097 (N_4097,N_3461,N_3546);
xnor U4098 (N_4098,N_3249,N_3591);
xor U4099 (N_4099,N_3342,N_3219);
xnor U4100 (N_4100,N_3622,N_3611);
and U4101 (N_4101,N_3301,N_3306);
and U4102 (N_4102,N_3155,N_3272);
nor U4103 (N_4103,N_3549,N_3646);
or U4104 (N_4104,N_3541,N_3527);
xnor U4105 (N_4105,N_3401,N_3606);
or U4106 (N_4106,N_3272,N_3177);
nor U4107 (N_4107,N_3728,N_3369);
nand U4108 (N_4108,N_3610,N_3686);
nor U4109 (N_4109,N_3749,N_3427);
or U4110 (N_4110,N_3540,N_3192);
or U4111 (N_4111,N_3665,N_3196);
xnor U4112 (N_4112,N_3379,N_3387);
and U4113 (N_4113,N_3500,N_3370);
or U4114 (N_4114,N_3396,N_3147);
or U4115 (N_4115,N_3307,N_3467);
xor U4116 (N_4116,N_3596,N_3701);
or U4117 (N_4117,N_3457,N_3697);
nor U4118 (N_4118,N_3493,N_3349);
nand U4119 (N_4119,N_3473,N_3630);
xnor U4120 (N_4120,N_3241,N_3141);
or U4121 (N_4121,N_3529,N_3587);
or U4122 (N_4122,N_3226,N_3214);
nand U4123 (N_4123,N_3686,N_3284);
nand U4124 (N_4124,N_3554,N_3157);
xnor U4125 (N_4125,N_3576,N_3131);
xor U4126 (N_4126,N_3381,N_3453);
nor U4127 (N_4127,N_3709,N_3325);
and U4128 (N_4128,N_3339,N_3362);
nand U4129 (N_4129,N_3475,N_3397);
and U4130 (N_4130,N_3449,N_3464);
or U4131 (N_4131,N_3528,N_3436);
xnor U4132 (N_4132,N_3623,N_3603);
xnor U4133 (N_4133,N_3702,N_3673);
nand U4134 (N_4134,N_3476,N_3679);
xnor U4135 (N_4135,N_3717,N_3311);
xor U4136 (N_4136,N_3339,N_3459);
xor U4137 (N_4137,N_3291,N_3342);
xnor U4138 (N_4138,N_3206,N_3496);
xnor U4139 (N_4139,N_3245,N_3510);
or U4140 (N_4140,N_3125,N_3319);
nand U4141 (N_4141,N_3648,N_3618);
or U4142 (N_4142,N_3445,N_3223);
xnor U4143 (N_4143,N_3189,N_3448);
nor U4144 (N_4144,N_3351,N_3354);
and U4145 (N_4145,N_3145,N_3467);
xnor U4146 (N_4146,N_3719,N_3339);
nor U4147 (N_4147,N_3689,N_3490);
xnor U4148 (N_4148,N_3357,N_3533);
xnor U4149 (N_4149,N_3701,N_3232);
nor U4150 (N_4150,N_3575,N_3380);
nor U4151 (N_4151,N_3557,N_3579);
nor U4152 (N_4152,N_3732,N_3677);
nor U4153 (N_4153,N_3414,N_3552);
xor U4154 (N_4154,N_3138,N_3254);
nor U4155 (N_4155,N_3695,N_3498);
and U4156 (N_4156,N_3462,N_3553);
nand U4157 (N_4157,N_3380,N_3348);
and U4158 (N_4158,N_3324,N_3169);
nor U4159 (N_4159,N_3191,N_3375);
nor U4160 (N_4160,N_3536,N_3627);
or U4161 (N_4161,N_3335,N_3285);
nor U4162 (N_4162,N_3349,N_3474);
or U4163 (N_4163,N_3148,N_3417);
or U4164 (N_4164,N_3284,N_3424);
or U4165 (N_4165,N_3594,N_3224);
xnor U4166 (N_4166,N_3445,N_3598);
or U4167 (N_4167,N_3396,N_3152);
nor U4168 (N_4168,N_3732,N_3508);
or U4169 (N_4169,N_3157,N_3397);
xnor U4170 (N_4170,N_3248,N_3413);
xor U4171 (N_4171,N_3281,N_3746);
nand U4172 (N_4172,N_3465,N_3459);
nor U4173 (N_4173,N_3268,N_3516);
or U4174 (N_4174,N_3716,N_3519);
or U4175 (N_4175,N_3597,N_3128);
nand U4176 (N_4176,N_3284,N_3503);
xnor U4177 (N_4177,N_3522,N_3748);
or U4178 (N_4178,N_3372,N_3403);
or U4179 (N_4179,N_3231,N_3698);
nand U4180 (N_4180,N_3609,N_3305);
xnor U4181 (N_4181,N_3714,N_3606);
nor U4182 (N_4182,N_3689,N_3722);
nand U4183 (N_4183,N_3597,N_3166);
nor U4184 (N_4184,N_3536,N_3533);
xnor U4185 (N_4185,N_3622,N_3177);
and U4186 (N_4186,N_3215,N_3385);
or U4187 (N_4187,N_3415,N_3741);
xor U4188 (N_4188,N_3326,N_3472);
nor U4189 (N_4189,N_3208,N_3357);
nor U4190 (N_4190,N_3687,N_3582);
and U4191 (N_4191,N_3576,N_3353);
nand U4192 (N_4192,N_3592,N_3646);
nor U4193 (N_4193,N_3174,N_3628);
or U4194 (N_4194,N_3626,N_3177);
and U4195 (N_4195,N_3342,N_3572);
nand U4196 (N_4196,N_3679,N_3278);
or U4197 (N_4197,N_3243,N_3731);
xnor U4198 (N_4198,N_3598,N_3222);
and U4199 (N_4199,N_3721,N_3232);
nor U4200 (N_4200,N_3343,N_3435);
nor U4201 (N_4201,N_3539,N_3697);
and U4202 (N_4202,N_3432,N_3493);
nand U4203 (N_4203,N_3185,N_3730);
nor U4204 (N_4204,N_3558,N_3379);
nor U4205 (N_4205,N_3603,N_3577);
or U4206 (N_4206,N_3172,N_3508);
xnor U4207 (N_4207,N_3374,N_3252);
and U4208 (N_4208,N_3372,N_3639);
and U4209 (N_4209,N_3335,N_3491);
nor U4210 (N_4210,N_3173,N_3523);
nand U4211 (N_4211,N_3335,N_3299);
or U4212 (N_4212,N_3248,N_3186);
nand U4213 (N_4213,N_3361,N_3621);
xnor U4214 (N_4214,N_3498,N_3734);
or U4215 (N_4215,N_3663,N_3637);
and U4216 (N_4216,N_3453,N_3546);
nor U4217 (N_4217,N_3620,N_3212);
xnor U4218 (N_4218,N_3685,N_3184);
nor U4219 (N_4219,N_3206,N_3332);
nand U4220 (N_4220,N_3712,N_3354);
nand U4221 (N_4221,N_3742,N_3744);
or U4222 (N_4222,N_3330,N_3716);
and U4223 (N_4223,N_3503,N_3613);
nor U4224 (N_4224,N_3749,N_3494);
or U4225 (N_4225,N_3574,N_3450);
nand U4226 (N_4226,N_3586,N_3716);
xnor U4227 (N_4227,N_3578,N_3490);
nor U4228 (N_4228,N_3336,N_3745);
nand U4229 (N_4229,N_3386,N_3146);
xor U4230 (N_4230,N_3615,N_3396);
or U4231 (N_4231,N_3204,N_3187);
nor U4232 (N_4232,N_3254,N_3428);
or U4233 (N_4233,N_3716,N_3748);
xor U4234 (N_4234,N_3505,N_3653);
and U4235 (N_4235,N_3729,N_3165);
xor U4236 (N_4236,N_3432,N_3617);
and U4237 (N_4237,N_3297,N_3172);
nand U4238 (N_4238,N_3618,N_3391);
and U4239 (N_4239,N_3637,N_3584);
or U4240 (N_4240,N_3696,N_3345);
or U4241 (N_4241,N_3616,N_3136);
nand U4242 (N_4242,N_3437,N_3317);
or U4243 (N_4243,N_3323,N_3480);
xor U4244 (N_4244,N_3166,N_3667);
xor U4245 (N_4245,N_3161,N_3245);
or U4246 (N_4246,N_3181,N_3478);
and U4247 (N_4247,N_3592,N_3133);
nand U4248 (N_4248,N_3167,N_3575);
xnor U4249 (N_4249,N_3718,N_3296);
nand U4250 (N_4250,N_3196,N_3669);
and U4251 (N_4251,N_3390,N_3473);
xor U4252 (N_4252,N_3545,N_3638);
nor U4253 (N_4253,N_3167,N_3529);
or U4254 (N_4254,N_3413,N_3726);
or U4255 (N_4255,N_3248,N_3324);
xor U4256 (N_4256,N_3360,N_3501);
xor U4257 (N_4257,N_3150,N_3467);
xnor U4258 (N_4258,N_3565,N_3208);
xor U4259 (N_4259,N_3507,N_3243);
nor U4260 (N_4260,N_3209,N_3257);
nor U4261 (N_4261,N_3673,N_3592);
xnor U4262 (N_4262,N_3310,N_3701);
nor U4263 (N_4263,N_3336,N_3577);
or U4264 (N_4264,N_3417,N_3229);
nand U4265 (N_4265,N_3599,N_3126);
xor U4266 (N_4266,N_3477,N_3484);
and U4267 (N_4267,N_3304,N_3456);
or U4268 (N_4268,N_3226,N_3546);
nor U4269 (N_4269,N_3664,N_3640);
nand U4270 (N_4270,N_3748,N_3343);
nand U4271 (N_4271,N_3745,N_3503);
xnor U4272 (N_4272,N_3331,N_3418);
or U4273 (N_4273,N_3347,N_3683);
xnor U4274 (N_4274,N_3327,N_3260);
and U4275 (N_4275,N_3474,N_3212);
or U4276 (N_4276,N_3603,N_3485);
xnor U4277 (N_4277,N_3405,N_3456);
nor U4278 (N_4278,N_3323,N_3335);
or U4279 (N_4279,N_3517,N_3161);
or U4280 (N_4280,N_3490,N_3239);
nor U4281 (N_4281,N_3157,N_3564);
nand U4282 (N_4282,N_3524,N_3551);
or U4283 (N_4283,N_3734,N_3209);
nand U4284 (N_4284,N_3607,N_3565);
nand U4285 (N_4285,N_3699,N_3378);
and U4286 (N_4286,N_3616,N_3293);
nor U4287 (N_4287,N_3664,N_3179);
and U4288 (N_4288,N_3503,N_3598);
xor U4289 (N_4289,N_3357,N_3187);
nand U4290 (N_4290,N_3695,N_3479);
nand U4291 (N_4291,N_3282,N_3737);
or U4292 (N_4292,N_3474,N_3736);
xor U4293 (N_4293,N_3566,N_3740);
xnor U4294 (N_4294,N_3711,N_3164);
nor U4295 (N_4295,N_3368,N_3633);
nor U4296 (N_4296,N_3231,N_3185);
xor U4297 (N_4297,N_3433,N_3541);
and U4298 (N_4298,N_3264,N_3212);
or U4299 (N_4299,N_3194,N_3435);
or U4300 (N_4300,N_3505,N_3318);
nor U4301 (N_4301,N_3535,N_3487);
nor U4302 (N_4302,N_3691,N_3585);
nor U4303 (N_4303,N_3283,N_3206);
and U4304 (N_4304,N_3707,N_3594);
nand U4305 (N_4305,N_3450,N_3372);
xnor U4306 (N_4306,N_3702,N_3696);
and U4307 (N_4307,N_3734,N_3294);
or U4308 (N_4308,N_3681,N_3472);
and U4309 (N_4309,N_3227,N_3585);
or U4310 (N_4310,N_3247,N_3555);
nor U4311 (N_4311,N_3672,N_3180);
nand U4312 (N_4312,N_3221,N_3719);
nand U4313 (N_4313,N_3194,N_3443);
nor U4314 (N_4314,N_3749,N_3255);
and U4315 (N_4315,N_3229,N_3339);
or U4316 (N_4316,N_3734,N_3335);
and U4317 (N_4317,N_3439,N_3368);
nor U4318 (N_4318,N_3307,N_3522);
and U4319 (N_4319,N_3355,N_3410);
nand U4320 (N_4320,N_3314,N_3437);
nor U4321 (N_4321,N_3640,N_3459);
xnor U4322 (N_4322,N_3585,N_3582);
nand U4323 (N_4323,N_3253,N_3665);
or U4324 (N_4324,N_3385,N_3185);
nand U4325 (N_4325,N_3691,N_3309);
and U4326 (N_4326,N_3408,N_3215);
xor U4327 (N_4327,N_3179,N_3608);
nor U4328 (N_4328,N_3443,N_3273);
xor U4329 (N_4329,N_3704,N_3178);
or U4330 (N_4330,N_3215,N_3503);
nand U4331 (N_4331,N_3343,N_3304);
nor U4332 (N_4332,N_3505,N_3537);
and U4333 (N_4333,N_3453,N_3188);
xor U4334 (N_4334,N_3369,N_3546);
xnor U4335 (N_4335,N_3684,N_3384);
xnor U4336 (N_4336,N_3352,N_3517);
and U4337 (N_4337,N_3640,N_3297);
and U4338 (N_4338,N_3633,N_3208);
nor U4339 (N_4339,N_3615,N_3260);
and U4340 (N_4340,N_3460,N_3425);
xor U4341 (N_4341,N_3391,N_3134);
nand U4342 (N_4342,N_3550,N_3266);
xor U4343 (N_4343,N_3295,N_3618);
nor U4344 (N_4344,N_3717,N_3255);
nand U4345 (N_4345,N_3708,N_3620);
nand U4346 (N_4346,N_3340,N_3550);
or U4347 (N_4347,N_3563,N_3386);
nor U4348 (N_4348,N_3149,N_3493);
nand U4349 (N_4349,N_3318,N_3686);
xnor U4350 (N_4350,N_3440,N_3676);
or U4351 (N_4351,N_3727,N_3616);
and U4352 (N_4352,N_3134,N_3224);
nor U4353 (N_4353,N_3546,N_3673);
or U4354 (N_4354,N_3739,N_3560);
nand U4355 (N_4355,N_3729,N_3307);
nand U4356 (N_4356,N_3718,N_3279);
and U4357 (N_4357,N_3412,N_3506);
nand U4358 (N_4358,N_3517,N_3400);
nand U4359 (N_4359,N_3442,N_3397);
and U4360 (N_4360,N_3511,N_3685);
and U4361 (N_4361,N_3366,N_3686);
nand U4362 (N_4362,N_3464,N_3245);
or U4363 (N_4363,N_3355,N_3345);
and U4364 (N_4364,N_3717,N_3382);
or U4365 (N_4365,N_3366,N_3656);
nand U4366 (N_4366,N_3624,N_3276);
and U4367 (N_4367,N_3319,N_3344);
and U4368 (N_4368,N_3675,N_3695);
or U4369 (N_4369,N_3335,N_3633);
and U4370 (N_4370,N_3174,N_3150);
or U4371 (N_4371,N_3514,N_3699);
xnor U4372 (N_4372,N_3368,N_3146);
or U4373 (N_4373,N_3276,N_3231);
and U4374 (N_4374,N_3184,N_3544);
nand U4375 (N_4375,N_3762,N_4180);
xor U4376 (N_4376,N_4320,N_3901);
xor U4377 (N_4377,N_3957,N_3913);
nor U4378 (N_4378,N_4252,N_4159);
and U4379 (N_4379,N_4280,N_4261);
or U4380 (N_4380,N_3785,N_4076);
nand U4381 (N_4381,N_4006,N_4057);
xnor U4382 (N_4382,N_3969,N_4354);
nor U4383 (N_4383,N_3825,N_3937);
nand U4384 (N_4384,N_4125,N_4153);
nand U4385 (N_4385,N_4060,N_4361);
nor U4386 (N_4386,N_3922,N_4066);
or U4387 (N_4387,N_4337,N_4187);
or U4388 (N_4388,N_4371,N_4161);
and U4389 (N_4389,N_3993,N_3888);
xnor U4390 (N_4390,N_4142,N_4219);
nor U4391 (N_4391,N_4362,N_3874);
or U4392 (N_4392,N_4129,N_4183);
nor U4393 (N_4393,N_3880,N_3926);
nand U4394 (N_4394,N_4214,N_4202);
xnor U4395 (N_4395,N_4245,N_4313);
and U4396 (N_4396,N_3934,N_4020);
or U4397 (N_4397,N_4349,N_3946);
nor U4398 (N_4398,N_4368,N_4072);
nor U4399 (N_4399,N_3989,N_4325);
nand U4400 (N_4400,N_4093,N_4097);
or U4401 (N_4401,N_4206,N_3751);
xnor U4402 (N_4402,N_4208,N_4330);
or U4403 (N_4403,N_4106,N_4373);
and U4404 (N_4404,N_4171,N_3782);
xor U4405 (N_4405,N_3925,N_4001);
nand U4406 (N_4406,N_3803,N_4071);
nand U4407 (N_4407,N_4108,N_4204);
or U4408 (N_4408,N_3871,N_4040);
or U4409 (N_4409,N_4021,N_3793);
xnor U4410 (N_4410,N_3779,N_4136);
nand U4411 (N_4411,N_4063,N_3960);
xor U4412 (N_4412,N_4025,N_4157);
nand U4413 (N_4413,N_4352,N_3933);
and U4414 (N_4414,N_4134,N_4084);
nor U4415 (N_4415,N_4326,N_3919);
nand U4416 (N_4416,N_4017,N_4314);
and U4417 (N_4417,N_3930,N_4168);
nor U4418 (N_4418,N_4177,N_4144);
nand U4419 (N_4419,N_3759,N_4286);
xor U4420 (N_4420,N_4207,N_4217);
xnor U4421 (N_4421,N_3988,N_4185);
nor U4422 (N_4422,N_3850,N_4149);
nor U4423 (N_4423,N_3795,N_4296);
xor U4424 (N_4424,N_3787,N_4317);
xnor U4425 (N_4425,N_4133,N_4227);
nor U4426 (N_4426,N_3774,N_3975);
xnor U4427 (N_4427,N_4119,N_4148);
and U4428 (N_4428,N_4143,N_4090);
and U4429 (N_4429,N_4348,N_4147);
xor U4430 (N_4430,N_4151,N_4290);
nor U4431 (N_4431,N_3833,N_4329);
xnor U4432 (N_4432,N_3861,N_4007);
nand U4433 (N_4433,N_3976,N_4229);
nand U4434 (N_4434,N_3773,N_3921);
or U4435 (N_4435,N_3947,N_3887);
nand U4436 (N_4436,N_3953,N_4141);
nor U4437 (N_4437,N_3906,N_4194);
and U4438 (N_4438,N_3826,N_3829);
nand U4439 (N_4439,N_4221,N_3778);
or U4440 (N_4440,N_3806,N_3883);
nor U4441 (N_4441,N_3894,N_4210);
or U4442 (N_4442,N_3973,N_4268);
and U4443 (N_4443,N_4075,N_4285);
nand U4444 (N_4444,N_4110,N_3903);
xor U4445 (N_4445,N_3941,N_3851);
and U4446 (N_4446,N_4140,N_3893);
or U4447 (N_4447,N_3789,N_4124);
and U4448 (N_4448,N_4045,N_4029);
xnor U4449 (N_4449,N_4074,N_4239);
nor U4450 (N_4450,N_4259,N_4033);
nand U4451 (N_4451,N_4089,N_3996);
and U4452 (N_4452,N_4275,N_4103);
or U4453 (N_4453,N_4253,N_3954);
nand U4454 (N_4454,N_4051,N_3990);
nor U4455 (N_4455,N_3780,N_4172);
nand U4456 (N_4456,N_4297,N_4356);
nor U4457 (N_4457,N_3836,N_3900);
nor U4458 (N_4458,N_4155,N_3827);
or U4459 (N_4459,N_4216,N_4321);
or U4460 (N_4460,N_4096,N_4218);
nor U4461 (N_4461,N_4092,N_4310);
and U4462 (N_4462,N_4228,N_4346);
or U4463 (N_4463,N_3766,N_3809);
and U4464 (N_4464,N_4027,N_4295);
nand U4465 (N_4465,N_4301,N_4241);
nand U4466 (N_4466,N_4294,N_3790);
xor U4467 (N_4467,N_3839,N_3974);
nand U4468 (N_4468,N_4340,N_4240);
xor U4469 (N_4469,N_4236,N_4191);
and U4470 (N_4470,N_3876,N_3799);
xor U4471 (N_4471,N_4199,N_4152);
and U4472 (N_4472,N_4196,N_4101);
nand U4473 (N_4473,N_4350,N_3945);
or U4474 (N_4474,N_3784,N_4169);
xnor U4475 (N_4475,N_4269,N_3964);
and U4476 (N_4476,N_3992,N_4367);
nand U4477 (N_4477,N_3949,N_3943);
xor U4478 (N_4478,N_4137,N_3889);
nor U4479 (N_4479,N_4122,N_4055);
nor U4480 (N_4480,N_4016,N_4192);
nand U4481 (N_4481,N_3791,N_4336);
nand U4482 (N_4482,N_3847,N_4234);
or U4483 (N_4483,N_4095,N_3805);
nor U4484 (N_4484,N_4249,N_4087);
and U4485 (N_4485,N_4083,N_3870);
or U4486 (N_4486,N_4070,N_4111);
and U4487 (N_4487,N_4248,N_3962);
nand U4488 (N_4488,N_3819,N_4156);
xor U4489 (N_4489,N_4267,N_4005);
and U4490 (N_4490,N_3940,N_4260);
nor U4491 (N_4491,N_3882,N_3842);
and U4492 (N_4492,N_3984,N_4195);
nor U4493 (N_4493,N_4044,N_3985);
or U4494 (N_4494,N_4176,N_4053);
nand U4495 (N_4495,N_3936,N_4166);
and U4496 (N_4496,N_4358,N_3886);
or U4497 (N_4497,N_3931,N_3935);
nor U4498 (N_4498,N_4127,N_4131);
and U4499 (N_4499,N_3820,N_4316);
or U4500 (N_4500,N_3783,N_4107);
nor U4501 (N_4501,N_4277,N_3877);
and U4502 (N_4502,N_4279,N_4130);
xnor U4503 (N_4503,N_3797,N_4041);
nand U4504 (N_4504,N_4233,N_4150);
nor U4505 (N_4505,N_4123,N_4292);
or U4506 (N_4506,N_3892,N_4170);
and U4507 (N_4507,N_4372,N_3864);
nand U4508 (N_4508,N_4324,N_4146);
or U4509 (N_4509,N_3927,N_3902);
nor U4510 (N_4510,N_3956,N_4303);
nor U4511 (N_4511,N_3917,N_3952);
xor U4512 (N_4512,N_3757,N_3841);
nand U4513 (N_4513,N_4281,N_3879);
and U4514 (N_4514,N_3763,N_3987);
nand U4515 (N_4515,N_4085,N_3951);
nand U4516 (N_4516,N_4263,N_3760);
and U4517 (N_4517,N_4132,N_3849);
nor U4518 (N_4518,N_3929,N_4175);
or U4519 (N_4519,N_4049,N_4081);
nor U4520 (N_4520,N_4365,N_3948);
or U4521 (N_4521,N_4311,N_4270);
nor U4522 (N_4522,N_3885,N_4312);
nor U4523 (N_4523,N_4154,N_4323);
and U4524 (N_4524,N_4167,N_4193);
and U4525 (N_4525,N_4306,N_4032);
xor U4526 (N_4526,N_4013,N_3875);
xor U4527 (N_4527,N_3979,N_3994);
xor U4528 (N_4528,N_3862,N_4265);
nand U4529 (N_4529,N_4028,N_4264);
xnor U4530 (N_4530,N_3899,N_4205);
or U4531 (N_4531,N_3950,N_4184);
and U4532 (N_4532,N_4360,N_4300);
and U4533 (N_4533,N_4008,N_4220);
nand U4534 (N_4534,N_3852,N_4094);
nand U4535 (N_4535,N_4364,N_3869);
nand U4536 (N_4536,N_4257,N_4067);
nor U4537 (N_4537,N_3752,N_3816);
nand U4538 (N_4538,N_4022,N_4116);
or U4539 (N_4539,N_4222,N_4256);
nand U4540 (N_4540,N_3765,N_4338);
xor U4541 (N_4541,N_3939,N_3968);
xor U4542 (N_4542,N_4363,N_3855);
and U4543 (N_4543,N_4158,N_4226);
nor U4544 (N_4544,N_4047,N_3776);
nand U4545 (N_4545,N_4009,N_4160);
xor U4546 (N_4546,N_4186,N_3831);
or U4547 (N_4547,N_3972,N_3770);
xnor U4548 (N_4548,N_4121,N_3798);
xor U4549 (N_4549,N_3755,N_4298);
nor U4550 (N_4550,N_4283,N_4366);
nor U4551 (N_4551,N_4004,N_4010);
nor U4552 (N_4552,N_4309,N_4225);
and U4553 (N_4553,N_4318,N_3978);
or U4554 (N_4554,N_4117,N_3955);
nor U4555 (N_4555,N_4282,N_4251);
nand U4556 (N_4556,N_4369,N_4339);
nor U4557 (N_4557,N_3853,N_4054);
and U4558 (N_4558,N_3923,N_3928);
and U4559 (N_4559,N_3998,N_4036);
xor U4560 (N_4560,N_4078,N_3966);
nor U4561 (N_4561,N_4198,N_4082);
nor U4562 (N_4562,N_4052,N_3812);
or U4563 (N_4563,N_4333,N_3844);
xnor U4564 (N_4564,N_4299,N_3977);
nand U4565 (N_4565,N_3897,N_4274);
nand U4566 (N_4566,N_3898,N_4182);
nor U4567 (N_4567,N_4014,N_4048);
and U4568 (N_4568,N_3971,N_4258);
or U4569 (N_4569,N_3838,N_3967);
xnor U4570 (N_4570,N_3944,N_4088);
xnor U4571 (N_4571,N_3981,N_3753);
nor U4572 (N_4572,N_4291,N_3801);
nand U4573 (N_4573,N_3970,N_4308);
xor U4574 (N_4574,N_4080,N_4209);
xnor U4575 (N_4575,N_3909,N_3907);
xor U4576 (N_4576,N_3932,N_3811);
xnor U4577 (N_4577,N_3878,N_3961);
xnor U4578 (N_4578,N_4343,N_4328);
xor U4579 (N_4579,N_4068,N_4064);
and U4580 (N_4580,N_4035,N_4197);
or U4581 (N_4581,N_3796,N_4015);
nand U4582 (N_4582,N_4288,N_4293);
and U4583 (N_4583,N_4120,N_4026);
or U4584 (N_4584,N_3915,N_4302);
nor U4585 (N_4585,N_3775,N_4128);
and U4586 (N_4586,N_4138,N_4062);
and U4587 (N_4587,N_3821,N_3808);
or U4588 (N_4588,N_4345,N_3758);
nor U4589 (N_4589,N_3896,N_4342);
xor U4590 (N_4590,N_3788,N_4213);
nand U4591 (N_4591,N_3781,N_4255);
xor U4592 (N_4592,N_4232,N_4109);
nand U4593 (N_4593,N_4099,N_4246);
nand U4594 (N_4594,N_4201,N_4203);
xor U4595 (N_4595,N_3777,N_4019);
or U4596 (N_4596,N_3840,N_3761);
nand U4597 (N_4597,N_4357,N_3817);
or U4598 (N_4598,N_4178,N_4077);
xor U4599 (N_4599,N_3995,N_3828);
nand U4600 (N_4600,N_3980,N_4327);
nand U4601 (N_4601,N_4304,N_3830);
or U4602 (N_4602,N_3848,N_4105);
nor U4603 (N_4603,N_3912,N_4231);
nor U4604 (N_4604,N_4273,N_4250);
or U4605 (N_4605,N_4059,N_4322);
or U4606 (N_4606,N_4031,N_4065);
nor U4607 (N_4607,N_3918,N_3772);
nand U4608 (N_4608,N_4102,N_3911);
nand U4609 (N_4609,N_3910,N_4024);
or U4610 (N_4610,N_4319,N_3916);
nor U4611 (N_4611,N_4100,N_3859);
nor U4612 (N_4612,N_3924,N_3837);
xor U4613 (N_4613,N_3754,N_4242);
and U4614 (N_4614,N_4165,N_4353);
xor U4615 (N_4615,N_3856,N_4179);
nor U4616 (N_4616,N_4262,N_4058);
nor U4617 (N_4617,N_3891,N_3938);
xor U4618 (N_4618,N_3818,N_4139);
xnor U4619 (N_4619,N_3814,N_4023);
and U4620 (N_4620,N_3884,N_4189);
nand U4621 (N_4621,N_4200,N_4069);
or U4622 (N_4622,N_3914,N_3834);
nor U4623 (N_4623,N_3858,N_4287);
xor U4624 (N_4624,N_3804,N_3802);
xor U4625 (N_4625,N_3786,N_4237);
or U4626 (N_4626,N_4098,N_4162);
nand U4627 (N_4627,N_3873,N_3991);
nor U4628 (N_4628,N_4126,N_3835);
nor U4629 (N_4629,N_4223,N_4276);
xor U4630 (N_4630,N_3997,N_3868);
xor U4631 (N_4631,N_3908,N_4284);
and U4632 (N_4632,N_3959,N_4091);
nor U4633 (N_4633,N_4042,N_3792);
or U4634 (N_4634,N_4254,N_4243);
or U4635 (N_4635,N_4012,N_4335);
and U4636 (N_4636,N_4002,N_3942);
nand U4637 (N_4637,N_4039,N_3832);
nand U4638 (N_4638,N_3794,N_4370);
xnor U4639 (N_4639,N_4135,N_4272);
nand U4640 (N_4640,N_4188,N_4000);
xnor U4641 (N_4641,N_4034,N_3843);
nor U4642 (N_4642,N_3958,N_3771);
xnor U4643 (N_4643,N_3920,N_4331);
nor U4644 (N_4644,N_4043,N_3807);
nor U4645 (N_4645,N_4289,N_4315);
xnor U4646 (N_4646,N_4118,N_3860);
or U4647 (N_4647,N_3983,N_3905);
nor U4648 (N_4648,N_4190,N_4215);
or U4649 (N_4649,N_4030,N_4073);
or U4650 (N_4650,N_4011,N_4174);
nand U4651 (N_4651,N_4334,N_4374);
or U4652 (N_4652,N_4163,N_3824);
nand U4653 (N_4653,N_4347,N_4145);
nand U4654 (N_4654,N_3854,N_4341);
xor U4655 (N_4655,N_4113,N_3963);
nand U4656 (N_4656,N_3769,N_4332);
nor U4657 (N_4657,N_3965,N_3756);
nor U4658 (N_4658,N_3764,N_3857);
or U4659 (N_4659,N_4018,N_3865);
or U4660 (N_4660,N_4307,N_3845);
nor U4661 (N_4661,N_4359,N_3904);
xor U4662 (N_4662,N_4244,N_4238);
nand U4663 (N_4663,N_3822,N_3999);
nand U4664 (N_4664,N_4086,N_4181);
nor U4665 (N_4665,N_3846,N_3982);
nand U4666 (N_4666,N_4212,N_4247);
xnor U4667 (N_4667,N_4224,N_3768);
or U4668 (N_4668,N_4211,N_3813);
and U4669 (N_4669,N_3810,N_4056);
or U4670 (N_4670,N_4235,N_3750);
and U4671 (N_4671,N_3800,N_4104);
nor U4672 (N_4672,N_4266,N_3866);
nor U4673 (N_4673,N_4115,N_4305);
xor U4674 (N_4674,N_4173,N_3863);
or U4675 (N_4675,N_3767,N_4164);
or U4676 (N_4676,N_4050,N_4061);
and U4677 (N_4677,N_4112,N_4230);
xor U4678 (N_4678,N_4046,N_4079);
and U4679 (N_4679,N_4355,N_4278);
and U4680 (N_4680,N_3890,N_3867);
and U4681 (N_4681,N_4003,N_4344);
nand U4682 (N_4682,N_4037,N_4271);
xor U4683 (N_4683,N_3986,N_3872);
nand U4684 (N_4684,N_4038,N_3823);
or U4685 (N_4685,N_3881,N_3815);
and U4686 (N_4686,N_4114,N_4351);
and U4687 (N_4687,N_3895,N_4049);
or U4688 (N_4688,N_4315,N_4281);
or U4689 (N_4689,N_4292,N_4333);
or U4690 (N_4690,N_3782,N_3982);
nor U4691 (N_4691,N_4188,N_4192);
and U4692 (N_4692,N_4191,N_4321);
nand U4693 (N_4693,N_4131,N_4138);
and U4694 (N_4694,N_4341,N_4130);
or U4695 (N_4695,N_3787,N_4116);
nor U4696 (N_4696,N_4177,N_4266);
xor U4697 (N_4697,N_4246,N_4232);
or U4698 (N_4698,N_4197,N_4036);
nor U4699 (N_4699,N_3755,N_4108);
xnor U4700 (N_4700,N_4306,N_3784);
and U4701 (N_4701,N_4314,N_4074);
and U4702 (N_4702,N_3974,N_4367);
and U4703 (N_4703,N_3770,N_4059);
xor U4704 (N_4704,N_4114,N_4317);
and U4705 (N_4705,N_3771,N_3950);
nor U4706 (N_4706,N_3961,N_4299);
nand U4707 (N_4707,N_4369,N_4255);
nand U4708 (N_4708,N_4344,N_3902);
and U4709 (N_4709,N_4013,N_4161);
and U4710 (N_4710,N_3829,N_4031);
nor U4711 (N_4711,N_3813,N_4081);
xnor U4712 (N_4712,N_4111,N_4282);
nand U4713 (N_4713,N_3816,N_3977);
and U4714 (N_4714,N_3753,N_3839);
xor U4715 (N_4715,N_3756,N_4270);
and U4716 (N_4716,N_3922,N_4341);
xnor U4717 (N_4717,N_3796,N_3898);
nor U4718 (N_4718,N_4363,N_4115);
and U4719 (N_4719,N_4119,N_4259);
nand U4720 (N_4720,N_4084,N_4313);
and U4721 (N_4721,N_4306,N_3814);
or U4722 (N_4722,N_4188,N_3879);
nand U4723 (N_4723,N_4031,N_3957);
or U4724 (N_4724,N_4300,N_3899);
nand U4725 (N_4725,N_3956,N_3778);
or U4726 (N_4726,N_3770,N_4144);
nand U4727 (N_4727,N_4046,N_4271);
nor U4728 (N_4728,N_4288,N_3808);
nand U4729 (N_4729,N_4268,N_3920);
xnor U4730 (N_4730,N_3952,N_4026);
or U4731 (N_4731,N_4199,N_4291);
xor U4732 (N_4732,N_4203,N_4362);
or U4733 (N_4733,N_3846,N_4275);
xnor U4734 (N_4734,N_4266,N_4150);
xnor U4735 (N_4735,N_3938,N_3988);
nand U4736 (N_4736,N_3884,N_3861);
nand U4737 (N_4737,N_4226,N_3891);
nor U4738 (N_4738,N_3799,N_4224);
or U4739 (N_4739,N_3988,N_4319);
and U4740 (N_4740,N_3866,N_4067);
nor U4741 (N_4741,N_3964,N_4298);
or U4742 (N_4742,N_4049,N_4094);
and U4743 (N_4743,N_3773,N_3815);
or U4744 (N_4744,N_3854,N_3864);
and U4745 (N_4745,N_4307,N_3985);
and U4746 (N_4746,N_4113,N_3929);
or U4747 (N_4747,N_3791,N_3825);
nor U4748 (N_4748,N_4338,N_3759);
nand U4749 (N_4749,N_4366,N_4049);
or U4750 (N_4750,N_4037,N_3756);
and U4751 (N_4751,N_4361,N_3751);
nand U4752 (N_4752,N_4293,N_4122);
nand U4753 (N_4753,N_3820,N_4194);
or U4754 (N_4754,N_4230,N_4315);
nand U4755 (N_4755,N_3854,N_4085);
and U4756 (N_4756,N_4122,N_4017);
or U4757 (N_4757,N_3868,N_3901);
nand U4758 (N_4758,N_4063,N_4211);
or U4759 (N_4759,N_3840,N_3768);
xor U4760 (N_4760,N_4173,N_3875);
nand U4761 (N_4761,N_3941,N_3974);
nand U4762 (N_4762,N_4016,N_3956);
and U4763 (N_4763,N_3828,N_4171);
nor U4764 (N_4764,N_4294,N_3839);
or U4765 (N_4765,N_3983,N_4275);
xor U4766 (N_4766,N_3990,N_3889);
nor U4767 (N_4767,N_3940,N_4078);
nor U4768 (N_4768,N_4143,N_3857);
xor U4769 (N_4769,N_3917,N_4023);
and U4770 (N_4770,N_3792,N_4257);
nor U4771 (N_4771,N_4001,N_4244);
or U4772 (N_4772,N_4355,N_4339);
and U4773 (N_4773,N_3830,N_3846);
and U4774 (N_4774,N_3753,N_3894);
xor U4775 (N_4775,N_4236,N_4241);
or U4776 (N_4776,N_4341,N_3766);
or U4777 (N_4777,N_3852,N_4108);
nor U4778 (N_4778,N_3939,N_4047);
or U4779 (N_4779,N_4206,N_4075);
and U4780 (N_4780,N_3995,N_3867);
nand U4781 (N_4781,N_3956,N_3981);
nand U4782 (N_4782,N_3886,N_4025);
nor U4783 (N_4783,N_4238,N_4098);
and U4784 (N_4784,N_3899,N_4337);
and U4785 (N_4785,N_4339,N_4335);
and U4786 (N_4786,N_4186,N_4326);
xor U4787 (N_4787,N_3880,N_3809);
nand U4788 (N_4788,N_3939,N_4234);
nor U4789 (N_4789,N_4028,N_3865);
xnor U4790 (N_4790,N_3915,N_4322);
or U4791 (N_4791,N_4018,N_3870);
xnor U4792 (N_4792,N_4370,N_4320);
nand U4793 (N_4793,N_3849,N_4001);
xor U4794 (N_4794,N_4332,N_3756);
xor U4795 (N_4795,N_3918,N_3880);
and U4796 (N_4796,N_4175,N_4128);
or U4797 (N_4797,N_4353,N_4067);
or U4798 (N_4798,N_3919,N_3864);
or U4799 (N_4799,N_4019,N_4263);
nand U4800 (N_4800,N_4023,N_4299);
or U4801 (N_4801,N_4312,N_3904);
or U4802 (N_4802,N_3769,N_4154);
nor U4803 (N_4803,N_3793,N_4018);
xor U4804 (N_4804,N_3912,N_3855);
nor U4805 (N_4805,N_3785,N_4011);
nand U4806 (N_4806,N_4170,N_4057);
nand U4807 (N_4807,N_4078,N_3851);
and U4808 (N_4808,N_4213,N_4108);
nor U4809 (N_4809,N_4256,N_3977);
and U4810 (N_4810,N_4298,N_4120);
or U4811 (N_4811,N_3897,N_4055);
xnor U4812 (N_4812,N_4319,N_4316);
nor U4813 (N_4813,N_4366,N_3763);
or U4814 (N_4814,N_4308,N_3910);
nand U4815 (N_4815,N_4030,N_4351);
or U4816 (N_4816,N_4198,N_3864);
or U4817 (N_4817,N_3940,N_3755);
xor U4818 (N_4818,N_3932,N_4343);
nor U4819 (N_4819,N_3834,N_4043);
and U4820 (N_4820,N_4203,N_4113);
nand U4821 (N_4821,N_4017,N_4234);
xor U4822 (N_4822,N_4005,N_3980);
nand U4823 (N_4823,N_4354,N_4036);
or U4824 (N_4824,N_3946,N_4314);
nand U4825 (N_4825,N_4318,N_4226);
xnor U4826 (N_4826,N_4336,N_4302);
and U4827 (N_4827,N_3932,N_4335);
xor U4828 (N_4828,N_3994,N_4249);
nand U4829 (N_4829,N_3832,N_4214);
or U4830 (N_4830,N_3813,N_3910);
nand U4831 (N_4831,N_4085,N_4361);
xnor U4832 (N_4832,N_4097,N_3771);
nand U4833 (N_4833,N_4229,N_4132);
and U4834 (N_4834,N_4283,N_4205);
nor U4835 (N_4835,N_4103,N_4253);
and U4836 (N_4836,N_4018,N_4302);
xor U4837 (N_4837,N_4264,N_4141);
and U4838 (N_4838,N_3903,N_3778);
nor U4839 (N_4839,N_4058,N_4289);
and U4840 (N_4840,N_4039,N_4077);
xnor U4841 (N_4841,N_4142,N_3991);
nor U4842 (N_4842,N_4351,N_4110);
or U4843 (N_4843,N_4177,N_4191);
and U4844 (N_4844,N_3882,N_3967);
xnor U4845 (N_4845,N_4034,N_3999);
xnor U4846 (N_4846,N_3862,N_4197);
nand U4847 (N_4847,N_3955,N_4361);
or U4848 (N_4848,N_4239,N_4261);
nand U4849 (N_4849,N_3952,N_4239);
xor U4850 (N_4850,N_4196,N_4195);
and U4851 (N_4851,N_3958,N_4327);
or U4852 (N_4852,N_4052,N_3806);
and U4853 (N_4853,N_4011,N_3856);
xnor U4854 (N_4854,N_4115,N_3904);
and U4855 (N_4855,N_4280,N_3816);
or U4856 (N_4856,N_4354,N_4060);
nand U4857 (N_4857,N_4030,N_4008);
nor U4858 (N_4858,N_3832,N_4064);
nor U4859 (N_4859,N_4156,N_3806);
nor U4860 (N_4860,N_4092,N_4155);
or U4861 (N_4861,N_3929,N_4292);
nand U4862 (N_4862,N_4247,N_4053);
nand U4863 (N_4863,N_4215,N_3950);
nand U4864 (N_4864,N_3770,N_3878);
and U4865 (N_4865,N_3986,N_4014);
or U4866 (N_4866,N_3820,N_4200);
nand U4867 (N_4867,N_3849,N_4225);
nor U4868 (N_4868,N_4085,N_4109);
xnor U4869 (N_4869,N_4372,N_3794);
or U4870 (N_4870,N_4183,N_4312);
nand U4871 (N_4871,N_4235,N_4033);
and U4872 (N_4872,N_4249,N_4218);
and U4873 (N_4873,N_3799,N_4111);
or U4874 (N_4874,N_3988,N_4042);
nor U4875 (N_4875,N_3948,N_4188);
or U4876 (N_4876,N_4093,N_4265);
and U4877 (N_4877,N_4081,N_4106);
and U4878 (N_4878,N_3980,N_4345);
and U4879 (N_4879,N_4318,N_4107);
nand U4880 (N_4880,N_4042,N_4190);
and U4881 (N_4881,N_4006,N_3759);
or U4882 (N_4882,N_3780,N_4304);
nand U4883 (N_4883,N_3918,N_4010);
nor U4884 (N_4884,N_3856,N_4187);
and U4885 (N_4885,N_3948,N_4090);
xor U4886 (N_4886,N_4203,N_4067);
nand U4887 (N_4887,N_4208,N_4063);
xnor U4888 (N_4888,N_3978,N_4122);
and U4889 (N_4889,N_4325,N_4125);
and U4890 (N_4890,N_3991,N_4064);
and U4891 (N_4891,N_4024,N_4047);
nand U4892 (N_4892,N_4001,N_4199);
nor U4893 (N_4893,N_4257,N_3979);
or U4894 (N_4894,N_4370,N_3817);
nand U4895 (N_4895,N_3864,N_3865);
and U4896 (N_4896,N_3907,N_3775);
nor U4897 (N_4897,N_3982,N_4183);
nand U4898 (N_4898,N_3876,N_4188);
nand U4899 (N_4899,N_4167,N_4040);
nor U4900 (N_4900,N_4296,N_4266);
xnor U4901 (N_4901,N_4359,N_4255);
and U4902 (N_4902,N_4351,N_4054);
nand U4903 (N_4903,N_3798,N_4076);
or U4904 (N_4904,N_3960,N_3814);
xnor U4905 (N_4905,N_4201,N_4018);
nor U4906 (N_4906,N_4173,N_4015);
and U4907 (N_4907,N_3773,N_4201);
or U4908 (N_4908,N_4090,N_4103);
and U4909 (N_4909,N_3928,N_4145);
or U4910 (N_4910,N_4350,N_3813);
nor U4911 (N_4911,N_4113,N_4345);
xnor U4912 (N_4912,N_3953,N_3851);
or U4913 (N_4913,N_3776,N_3808);
xnor U4914 (N_4914,N_3795,N_4027);
or U4915 (N_4915,N_4013,N_4300);
nor U4916 (N_4916,N_3811,N_3788);
and U4917 (N_4917,N_4078,N_4186);
and U4918 (N_4918,N_3798,N_3916);
and U4919 (N_4919,N_3774,N_3895);
and U4920 (N_4920,N_3808,N_3774);
or U4921 (N_4921,N_4181,N_3925);
or U4922 (N_4922,N_3919,N_4246);
or U4923 (N_4923,N_3835,N_3820);
or U4924 (N_4924,N_3808,N_4045);
or U4925 (N_4925,N_4258,N_4226);
xor U4926 (N_4926,N_3994,N_4052);
nor U4927 (N_4927,N_3919,N_4007);
xnor U4928 (N_4928,N_4320,N_4227);
xor U4929 (N_4929,N_3830,N_3928);
or U4930 (N_4930,N_4358,N_4112);
xor U4931 (N_4931,N_3821,N_4206);
or U4932 (N_4932,N_4274,N_3923);
or U4933 (N_4933,N_3801,N_4142);
and U4934 (N_4934,N_4234,N_3924);
nor U4935 (N_4935,N_3853,N_3798);
nand U4936 (N_4936,N_4038,N_4300);
or U4937 (N_4937,N_4003,N_4176);
or U4938 (N_4938,N_3758,N_4048);
nand U4939 (N_4939,N_4213,N_3820);
nor U4940 (N_4940,N_3861,N_3905);
and U4941 (N_4941,N_4171,N_3851);
xnor U4942 (N_4942,N_4067,N_3928);
nor U4943 (N_4943,N_4111,N_4034);
or U4944 (N_4944,N_3761,N_4015);
nor U4945 (N_4945,N_4258,N_3940);
xnor U4946 (N_4946,N_4000,N_4310);
or U4947 (N_4947,N_3848,N_4288);
or U4948 (N_4948,N_4282,N_4181);
and U4949 (N_4949,N_4369,N_4190);
or U4950 (N_4950,N_4205,N_3769);
nand U4951 (N_4951,N_4296,N_3993);
xnor U4952 (N_4952,N_4362,N_4138);
or U4953 (N_4953,N_4155,N_3786);
nor U4954 (N_4954,N_4189,N_3804);
nand U4955 (N_4955,N_4230,N_3992);
xor U4956 (N_4956,N_3913,N_4191);
nor U4957 (N_4957,N_3762,N_3787);
xor U4958 (N_4958,N_4340,N_4308);
nand U4959 (N_4959,N_4252,N_3977);
and U4960 (N_4960,N_4357,N_4016);
nor U4961 (N_4961,N_3920,N_3874);
and U4962 (N_4962,N_3847,N_3914);
nor U4963 (N_4963,N_4190,N_3770);
nand U4964 (N_4964,N_3807,N_4333);
xor U4965 (N_4965,N_4029,N_4048);
nand U4966 (N_4966,N_4311,N_3890);
or U4967 (N_4967,N_4319,N_4158);
nand U4968 (N_4968,N_4216,N_3972);
xor U4969 (N_4969,N_4046,N_3797);
and U4970 (N_4970,N_4261,N_4108);
or U4971 (N_4971,N_4123,N_4039);
nand U4972 (N_4972,N_4184,N_4104);
nand U4973 (N_4973,N_4250,N_4209);
nor U4974 (N_4974,N_4307,N_3812);
and U4975 (N_4975,N_4355,N_4350);
nand U4976 (N_4976,N_4176,N_4144);
and U4977 (N_4977,N_4044,N_3964);
xnor U4978 (N_4978,N_3873,N_4205);
nor U4979 (N_4979,N_4219,N_4178);
xnor U4980 (N_4980,N_4275,N_4360);
xor U4981 (N_4981,N_4343,N_3974);
or U4982 (N_4982,N_3750,N_4118);
or U4983 (N_4983,N_3862,N_3777);
and U4984 (N_4984,N_4062,N_3866);
nand U4985 (N_4985,N_3951,N_4249);
and U4986 (N_4986,N_4060,N_3902);
xnor U4987 (N_4987,N_3921,N_3949);
xnor U4988 (N_4988,N_4057,N_4030);
nand U4989 (N_4989,N_4228,N_4331);
nor U4990 (N_4990,N_3798,N_4012);
nand U4991 (N_4991,N_3902,N_4015);
nand U4992 (N_4992,N_3910,N_4134);
nor U4993 (N_4993,N_3773,N_4369);
nand U4994 (N_4994,N_3892,N_3999);
xor U4995 (N_4995,N_3788,N_3793);
xor U4996 (N_4996,N_4141,N_4302);
and U4997 (N_4997,N_4254,N_4241);
or U4998 (N_4998,N_3884,N_4005);
nor U4999 (N_4999,N_3932,N_4347);
xor U5000 (N_5000,N_4626,N_4987);
and U5001 (N_5001,N_4992,N_4761);
nor U5002 (N_5002,N_4694,N_4946);
or U5003 (N_5003,N_4498,N_4459);
nand U5004 (N_5004,N_4879,N_4656);
xor U5005 (N_5005,N_4468,N_4995);
and U5006 (N_5006,N_4874,N_4377);
nand U5007 (N_5007,N_4617,N_4475);
and U5008 (N_5008,N_4641,N_4764);
or U5009 (N_5009,N_4619,N_4543);
and U5010 (N_5010,N_4984,N_4702);
or U5011 (N_5011,N_4918,N_4881);
or U5012 (N_5012,N_4962,N_4862);
nor U5013 (N_5013,N_4974,N_4418);
or U5014 (N_5014,N_4808,N_4999);
nand U5015 (N_5015,N_4696,N_4826);
nor U5016 (N_5016,N_4965,N_4926);
or U5017 (N_5017,N_4940,N_4513);
xnor U5018 (N_5018,N_4894,N_4506);
or U5019 (N_5019,N_4966,N_4923);
and U5020 (N_5020,N_4857,N_4653);
xnor U5021 (N_5021,N_4781,N_4440);
nor U5022 (N_5022,N_4509,N_4618);
and U5023 (N_5023,N_4804,N_4510);
nor U5024 (N_5024,N_4724,N_4429);
and U5025 (N_5025,N_4603,N_4751);
or U5026 (N_5026,N_4593,N_4929);
nor U5027 (N_5027,N_4456,N_4785);
nor U5028 (N_5028,N_4975,N_4793);
xnor U5029 (N_5029,N_4886,N_4563);
and U5030 (N_5030,N_4730,N_4507);
or U5031 (N_5031,N_4744,N_4909);
nor U5032 (N_5032,N_4531,N_4592);
or U5033 (N_5033,N_4670,N_4508);
nor U5034 (N_5034,N_4994,N_4847);
or U5035 (N_5035,N_4599,N_4578);
nand U5036 (N_5036,N_4411,N_4956);
nor U5037 (N_5037,N_4738,N_4829);
xnor U5038 (N_5038,N_4778,N_4550);
xor U5039 (N_5039,N_4562,N_4587);
nand U5040 (N_5040,N_4579,N_4969);
and U5041 (N_5041,N_4988,N_4824);
and U5042 (N_5042,N_4635,N_4444);
and U5043 (N_5043,N_4941,N_4648);
xor U5044 (N_5044,N_4671,N_4892);
nor U5045 (N_5045,N_4404,N_4771);
nor U5046 (N_5046,N_4750,N_4825);
or U5047 (N_5047,N_4376,N_4476);
nand U5048 (N_5048,N_4414,N_4695);
xor U5049 (N_5049,N_4789,N_4466);
nor U5050 (N_5050,N_4875,N_4767);
nor U5051 (N_5051,N_4640,N_4604);
nor U5052 (N_5052,N_4998,N_4553);
nand U5053 (N_5053,N_4649,N_4853);
xnor U5054 (N_5054,N_4457,N_4484);
nor U5055 (N_5055,N_4814,N_4739);
nor U5056 (N_5056,N_4436,N_4682);
nor U5057 (N_5057,N_4834,N_4405);
nor U5058 (N_5058,N_4445,N_4614);
nand U5059 (N_5059,N_4512,N_4547);
or U5060 (N_5060,N_4548,N_4375);
xor U5061 (N_5061,N_4668,N_4933);
nor U5062 (N_5062,N_4928,N_4759);
and U5063 (N_5063,N_4661,N_4446);
or U5064 (N_5064,N_4514,N_4849);
nand U5065 (N_5065,N_4838,N_4719);
xnor U5066 (N_5066,N_4413,N_4527);
or U5067 (N_5067,N_4938,N_4397);
nor U5068 (N_5068,N_4707,N_4907);
and U5069 (N_5069,N_4708,N_4805);
xnor U5070 (N_5070,N_4625,N_4726);
and U5071 (N_5071,N_4950,N_4557);
and U5072 (N_5072,N_4632,N_4428);
xnor U5073 (N_5073,N_4952,N_4417);
xor U5074 (N_5074,N_4896,N_4817);
nor U5075 (N_5075,N_4379,N_4914);
xor U5076 (N_5076,N_4700,N_4930);
nor U5077 (N_5077,N_4754,N_4423);
xnor U5078 (N_5078,N_4441,N_4678);
and U5079 (N_5079,N_4383,N_4588);
xor U5080 (N_5080,N_4699,N_4891);
and U5081 (N_5081,N_4921,N_4731);
or U5082 (N_5082,N_4747,N_4584);
or U5083 (N_5083,N_4673,N_4679);
nand U5084 (N_5084,N_4692,N_4800);
or U5085 (N_5085,N_4607,N_4981);
or U5086 (N_5086,N_4403,N_4431);
or U5087 (N_5087,N_4585,N_4740);
xnor U5088 (N_5088,N_4898,N_4791);
nor U5089 (N_5089,N_4811,N_4654);
or U5090 (N_5090,N_4645,N_4887);
nand U5091 (N_5091,N_4821,N_4398);
and U5092 (N_5092,N_4608,N_4580);
xnor U5093 (N_5093,N_4684,N_4657);
xor U5094 (N_5094,N_4602,N_4637);
xor U5095 (N_5095,N_4972,N_4442);
nand U5096 (N_5096,N_4903,N_4705);
or U5097 (N_5097,N_4876,N_4421);
nand U5098 (N_5098,N_4452,N_4908);
nand U5099 (N_5099,N_4801,N_4920);
and U5100 (N_5100,N_4480,N_4552);
or U5101 (N_5101,N_4523,N_4772);
or U5102 (N_5102,N_4943,N_4427);
xor U5103 (N_5103,N_4504,N_4683);
and U5104 (N_5104,N_4944,N_4409);
nor U5105 (N_5105,N_4652,N_4776);
and U5106 (N_5106,N_4897,N_4878);
or U5107 (N_5107,N_4471,N_4732);
or U5108 (N_5108,N_4766,N_4674);
and U5109 (N_5109,N_4860,N_4985);
xor U5110 (N_5110,N_4823,N_4917);
xor U5111 (N_5111,N_4520,N_4681);
xnor U5112 (N_5112,N_4386,N_4790);
or U5113 (N_5113,N_4487,N_4991);
or U5114 (N_5114,N_4701,N_4400);
nor U5115 (N_5115,N_4884,N_4447);
nor U5116 (N_5116,N_4852,N_4979);
xor U5117 (N_5117,N_4755,N_4490);
nor U5118 (N_5118,N_4961,N_4639);
nor U5119 (N_5119,N_4560,N_4566);
and U5120 (N_5120,N_4443,N_4752);
or U5121 (N_5121,N_4463,N_4408);
and U5122 (N_5122,N_4983,N_4963);
and U5123 (N_5123,N_4872,N_4746);
or U5124 (N_5124,N_4477,N_4910);
xnor U5125 (N_5125,N_4675,N_4885);
xor U5126 (N_5126,N_4812,N_4720);
xnor U5127 (N_5127,N_4783,N_4378);
and U5128 (N_5128,N_4434,N_4728);
or U5129 (N_5129,N_4802,N_4822);
or U5130 (N_5130,N_4402,N_4807);
nor U5131 (N_5131,N_4798,N_4686);
and U5132 (N_5132,N_4816,N_4380);
and U5133 (N_5133,N_4902,N_4606);
nand U5134 (N_5134,N_4615,N_4664);
or U5135 (N_5135,N_4818,N_4833);
xnor U5136 (N_5136,N_4538,N_4577);
xor U5137 (N_5137,N_4745,N_4757);
or U5138 (N_5138,N_4422,N_4864);
xnor U5139 (N_5139,N_4937,N_4871);
and U5140 (N_5140,N_4688,N_4388);
nand U5141 (N_5141,N_4556,N_4554);
xnor U5142 (N_5142,N_4597,N_4882);
nand U5143 (N_5143,N_4448,N_4387);
nor U5144 (N_5144,N_4742,N_4620);
and U5145 (N_5145,N_4532,N_4623);
nor U5146 (N_5146,N_4646,N_4610);
xnor U5147 (N_5147,N_4458,N_4769);
xnor U5148 (N_5148,N_4787,N_4415);
and U5149 (N_5149,N_4697,N_4954);
nand U5150 (N_5150,N_4890,N_4672);
and U5151 (N_5151,N_4438,N_4912);
nor U5152 (N_5152,N_4989,N_4718);
nor U5153 (N_5153,N_4703,N_4722);
xor U5154 (N_5154,N_4832,N_4780);
or U5155 (N_5155,N_4582,N_4736);
and U5156 (N_5156,N_4714,N_4555);
nand U5157 (N_5157,N_4687,N_4870);
nand U5158 (N_5158,N_4927,N_4502);
and U5159 (N_5159,N_4629,N_4986);
nor U5160 (N_5160,N_4693,N_4919);
xor U5161 (N_5161,N_4549,N_4873);
or U5162 (N_5162,N_4643,N_4899);
or U5163 (N_5163,N_4601,N_4401);
nor U5164 (N_5164,N_4942,N_4454);
and U5165 (N_5165,N_4605,N_4727);
or U5166 (N_5166,N_4779,N_4544);
and U5167 (N_5167,N_4970,N_4916);
nand U5168 (N_5168,N_4644,N_4841);
nand U5169 (N_5169,N_4964,N_4494);
xnor U5170 (N_5170,N_4600,N_4934);
or U5171 (N_5171,N_4830,N_4996);
or U5172 (N_5172,N_4385,N_4689);
xnor U5173 (N_5173,N_4488,N_4535);
or U5174 (N_5174,N_4665,N_4716);
or U5175 (N_5175,N_4658,N_4844);
and U5176 (N_5176,N_4794,N_4416);
and U5177 (N_5177,N_4435,N_4888);
or U5178 (N_5178,N_4541,N_4537);
or U5179 (N_5179,N_4893,N_4889);
nand U5180 (N_5180,N_4638,N_4710);
nor U5181 (N_5181,N_4546,N_4704);
nor U5182 (N_5182,N_4483,N_4472);
and U5183 (N_5183,N_4460,N_4485);
xnor U5184 (N_5184,N_4449,N_4612);
nor U5185 (N_5185,N_4799,N_4721);
or U5186 (N_5186,N_4863,N_4828);
xor U5187 (N_5187,N_4424,N_4997);
nand U5188 (N_5188,N_4925,N_4499);
or U5189 (N_5189,N_4904,N_4384);
or U5190 (N_5190,N_4971,N_4880);
xnor U5191 (N_5191,N_4741,N_4611);
xnor U5192 (N_5192,N_4990,N_4573);
nor U5193 (N_5193,N_4809,N_4810);
xnor U5194 (N_5194,N_4848,N_4394);
xor U5195 (N_5195,N_4945,N_4777);
and U5196 (N_5196,N_4496,N_4539);
and U5197 (N_5197,N_4594,N_4479);
xor U5198 (N_5198,N_4503,N_4806);
xnor U5199 (N_5199,N_4939,N_4486);
xnor U5200 (N_5200,N_4521,N_4450);
or U5201 (N_5201,N_4518,N_4955);
nor U5202 (N_5202,N_4854,N_4391);
xnor U5203 (N_5203,N_4568,N_4725);
or U5204 (N_5204,N_4935,N_4900);
or U5205 (N_5205,N_4712,N_4437);
xor U5206 (N_5206,N_4564,N_4395);
xnor U5207 (N_5207,N_4647,N_4627);
xnor U5208 (N_5208,N_4565,N_4768);
nand U5209 (N_5209,N_4381,N_4760);
xnor U5210 (N_5210,N_4478,N_4856);
nor U5211 (N_5211,N_4973,N_4396);
and U5212 (N_5212,N_4389,N_4851);
xor U5213 (N_5213,N_4784,N_4795);
nand U5214 (N_5214,N_4501,N_4591);
xnor U5215 (N_5215,N_4792,N_4839);
nand U5216 (N_5216,N_4677,N_4574);
or U5217 (N_5217,N_4651,N_4432);
nand U5218 (N_5218,N_4765,N_4932);
and U5219 (N_5219,N_4958,N_4774);
or U5220 (N_5220,N_4978,N_4412);
xnor U5221 (N_5221,N_4390,N_4621);
nand U5222 (N_5222,N_4706,N_4467);
or U5223 (N_5223,N_4551,N_4931);
nand U5224 (N_5224,N_4859,N_4685);
nor U5225 (N_5225,N_4815,N_4559);
or U5226 (N_5226,N_4598,N_4711);
xor U5227 (N_5227,N_4519,N_4426);
and U5228 (N_5228,N_4763,N_4855);
nand U5229 (N_5229,N_4425,N_4906);
or U5230 (N_5230,N_4609,N_4583);
nor U5231 (N_5231,N_4516,N_4676);
or U5232 (N_5232,N_4831,N_4782);
nand U5233 (N_5233,N_4869,N_4515);
nand U5234 (N_5234,N_4877,N_4461);
nor U5235 (N_5235,N_4861,N_4846);
xnor U5236 (N_5236,N_4883,N_4500);
and U5237 (N_5237,N_4419,N_4545);
nor U5238 (N_5238,N_4960,N_4840);
nand U5239 (N_5239,N_4430,N_4663);
and U5240 (N_5240,N_4723,N_4735);
or U5241 (N_5241,N_4756,N_4473);
xnor U5242 (N_5242,N_4481,N_4382);
xor U5243 (N_5243,N_4713,N_4948);
xnor U5244 (N_5244,N_4786,N_4529);
and U5245 (N_5245,N_4775,N_4915);
xnor U5246 (N_5246,N_4843,N_4631);
or U5247 (N_5247,N_4717,N_4406);
or U5248 (N_5248,N_4530,N_4469);
or U5249 (N_5249,N_4850,N_4455);
nand U5250 (N_5250,N_4525,N_4797);
or U5251 (N_5251,N_4526,N_4511);
xor U5252 (N_5252,N_4842,N_4819);
xnor U5253 (N_5253,N_4586,N_4533);
nand U5254 (N_5254,N_4911,N_4570);
or U5255 (N_5255,N_4493,N_4613);
or U5256 (N_5256,N_4392,N_4758);
or U5257 (N_5257,N_4492,N_4953);
nand U5258 (N_5258,N_4462,N_4837);
or U5259 (N_5259,N_4495,N_4616);
nand U5260 (N_5260,N_4836,N_4659);
nand U5261 (N_5261,N_4650,N_4709);
or U5262 (N_5262,N_4749,N_4867);
and U5263 (N_5263,N_4770,N_4451);
or U5264 (N_5264,N_4517,N_4628);
and U5265 (N_5265,N_4420,N_4505);
and U5266 (N_5266,N_4439,N_4596);
or U5267 (N_5267,N_4957,N_4690);
xor U5268 (N_5268,N_4820,N_4866);
xor U5269 (N_5269,N_4977,N_4407);
xor U5270 (N_5270,N_4655,N_4967);
nand U5271 (N_5271,N_4753,N_4715);
nor U5272 (N_5272,N_4922,N_4491);
nand U5273 (N_5273,N_4558,N_4464);
or U5274 (N_5274,N_4976,N_4571);
nor U5275 (N_5275,N_4489,N_4536);
nor U5276 (N_5276,N_4947,N_4729);
xnor U5277 (N_5277,N_4680,N_4575);
xnor U5278 (N_5278,N_4951,N_4773);
or U5279 (N_5279,N_4576,N_4410);
nor U5280 (N_5280,N_4524,N_4636);
xor U5281 (N_5281,N_4788,N_4465);
nand U5282 (N_5282,N_4734,N_4924);
or U5283 (N_5283,N_4803,N_4895);
nand U5284 (N_5284,N_4733,N_4762);
xor U5285 (N_5285,N_4993,N_4968);
xnor U5286 (N_5286,N_4569,N_4737);
xnor U5287 (N_5287,N_4748,N_4865);
and U5288 (N_5288,N_4813,N_4669);
or U5289 (N_5289,N_4622,N_4959);
nor U5290 (N_5290,N_4634,N_4858);
or U5291 (N_5291,N_4642,N_4595);
and U5292 (N_5292,N_4474,N_4590);
or U5293 (N_5293,N_4666,N_4453);
nand U5294 (N_5294,N_4868,N_4581);
xor U5295 (N_5295,N_4572,N_4743);
nor U5296 (N_5296,N_4534,N_4698);
or U5297 (N_5297,N_4691,N_4980);
nand U5298 (N_5298,N_4949,N_4913);
or U5299 (N_5299,N_4522,N_4567);
nor U5300 (N_5300,N_4528,N_4624);
or U5301 (N_5301,N_4630,N_4540);
and U5302 (N_5302,N_4796,N_4433);
xor U5303 (N_5303,N_4835,N_4633);
xor U5304 (N_5304,N_4482,N_4662);
nand U5305 (N_5305,N_4667,N_4399);
and U5306 (N_5306,N_4470,N_4901);
nand U5307 (N_5307,N_4589,N_4497);
or U5308 (N_5308,N_4660,N_4542);
nor U5309 (N_5309,N_4827,N_4393);
nand U5310 (N_5310,N_4905,N_4936);
or U5311 (N_5311,N_4982,N_4561);
or U5312 (N_5312,N_4845,N_4891);
nor U5313 (N_5313,N_4820,N_4977);
xor U5314 (N_5314,N_4635,N_4832);
nand U5315 (N_5315,N_4583,N_4740);
or U5316 (N_5316,N_4793,N_4552);
xor U5317 (N_5317,N_4977,N_4828);
nand U5318 (N_5318,N_4703,N_4729);
and U5319 (N_5319,N_4910,N_4713);
nor U5320 (N_5320,N_4700,N_4947);
xnor U5321 (N_5321,N_4492,N_4728);
or U5322 (N_5322,N_4933,N_4693);
xor U5323 (N_5323,N_4759,N_4662);
or U5324 (N_5324,N_4585,N_4475);
nor U5325 (N_5325,N_4455,N_4746);
or U5326 (N_5326,N_4512,N_4446);
nand U5327 (N_5327,N_4958,N_4832);
nand U5328 (N_5328,N_4862,N_4674);
nand U5329 (N_5329,N_4579,N_4815);
and U5330 (N_5330,N_4418,N_4488);
nor U5331 (N_5331,N_4806,N_4851);
nor U5332 (N_5332,N_4570,N_4902);
and U5333 (N_5333,N_4732,N_4509);
and U5334 (N_5334,N_4901,N_4745);
or U5335 (N_5335,N_4597,N_4453);
and U5336 (N_5336,N_4729,N_4979);
nand U5337 (N_5337,N_4778,N_4981);
xor U5338 (N_5338,N_4517,N_4643);
and U5339 (N_5339,N_4665,N_4521);
xnor U5340 (N_5340,N_4739,N_4391);
or U5341 (N_5341,N_4625,N_4676);
nor U5342 (N_5342,N_4451,N_4631);
nor U5343 (N_5343,N_4628,N_4591);
xor U5344 (N_5344,N_4578,N_4539);
xor U5345 (N_5345,N_4735,N_4675);
xor U5346 (N_5346,N_4846,N_4742);
xnor U5347 (N_5347,N_4607,N_4474);
or U5348 (N_5348,N_4717,N_4884);
xnor U5349 (N_5349,N_4617,N_4552);
nor U5350 (N_5350,N_4685,N_4725);
xnor U5351 (N_5351,N_4979,N_4945);
and U5352 (N_5352,N_4939,N_4383);
or U5353 (N_5353,N_4651,N_4817);
nand U5354 (N_5354,N_4823,N_4964);
xor U5355 (N_5355,N_4545,N_4665);
or U5356 (N_5356,N_4609,N_4671);
and U5357 (N_5357,N_4606,N_4974);
or U5358 (N_5358,N_4508,N_4803);
nor U5359 (N_5359,N_4963,N_4948);
nor U5360 (N_5360,N_4585,N_4951);
xor U5361 (N_5361,N_4445,N_4448);
xnor U5362 (N_5362,N_4746,N_4702);
nand U5363 (N_5363,N_4976,N_4376);
nor U5364 (N_5364,N_4872,N_4815);
and U5365 (N_5365,N_4460,N_4837);
and U5366 (N_5366,N_4983,N_4843);
nor U5367 (N_5367,N_4473,N_4650);
or U5368 (N_5368,N_4458,N_4997);
or U5369 (N_5369,N_4445,N_4592);
nand U5370 (N_5370,N_4494,N_4711);
xnor U5371 (N_5371,N_4954,N_4450);
or U5372 (N_5372,N_4683,N_4858);
or U5373 (N_5373,N_4991,N_4796);
and U5374 (N_5374,N_4449,N_4392);
xnor U5375 (N_5375,N_4431,N_4496);
xor U5376 (N_5376,N_4544,N_4696);
or U5377 (N_5377,N_4680,N_4591);
or U5378 (N_5378,N_4676,N_4956);
nor U5379 (N_5379,N_4952,N_4407);
nor U5380 (N_5380,N_4943,N_4743);
or U5381 (N_5381,N_4383,N_4758);
or U5382 (N_5382,N_4609,N_4780);
or U5383 (N_5383,N_4667,N_4823);
and U5384 (N_5384,N_4478,N_4498);
nand U5385 (N_5385,N_4500,N_4536);
or U5386 (N_5386,N_4967,N_4377);
and U5387 (N_5387,N_4713,N_4788);
xor U5388 (N_5388,N_4510,N_4647);
xor U5389 (N_5389,N_4848,N_4629);
nand U5390 (N_5390,N_4415,N_4510);
nor U5391 (N_5391,N_4588,N_4826);
or U5392 (N_5392,N_4527,N_4600);
or U5393 (N_5393,N_4821,N_4436);
nor U5394 (N_5394,N_4976,N_4840);
xor U5395 (N_5395,N_4852,N_4424);
xor U5396 (N_5396,N_4630,N_4629);
xor U5397 (N_5397,N_4796,N_4609);
or U5398 (N_5398,N_4962,N_4798);
and U5399 (N_5399,N_4916,N_4868);
xnor U5400 (N_5400,N_4625,N_4480);
nand U5401 (N_5401,N_4763,N_4583);
or U5402 (N_5402,N_4559,N_4701);
nand U5403 (N_5403,N_4778,N_4662);
xor U5404 (N_5404,N_4383,N_4473);
xnor U5405 (N_5405,N_4836,N_4789);
nand U5406 (N_5406,N_4990,N_4382);
and U5407 (N_5407,N_4390,N_4733);
xor U5408 (N_5408,N_4430,N_4551);
nor U5409 (N_5409,N_4443,N_4680);
and U5410 (N_5410,N_4472,N_4484);
xor U5411 (N_5411,N_4743,N_4381);
nor U5412 (N_5412,N_4565,N_4716);
xnor U5413 (N_5413,N_4746,N_4696);
and U5414 (N_5414,N_4646,N_4899);
or U5415 (N_5415,N_4574,N_4976);
nand U5416 (N_5416,N_4487,N_4675);
xor U5417 (N_5417,N_4702,N_4887);
and U5418 (N_5418,N_4487,N_4614);
and U5419 (N_5419,N_4813,N_4670);
nor U5420 (N_5420,N_4637,N_4527);
or U5421 (N_5421,N_4826,N_4719);
nand U5422 (N_5422,N_4677,N_4985);
and U5423 (N_5423,N_4712,N_4773);
nand U5424 (N_5424,N_4785,N_4616);
nand U5425 (N_5425,N_4416,N_4508);
or U5426 (N_5426,N_4396,N_4691);
nor U5427 (N_5427,N_4929,N_4719);
and U5428 (N_5428,N_4917,N_4680);
nor U5429 (N_5429,N_4469,N_4731);
and U5430 (N_5430,N_4739,N_4659);
xnor U5431 (N_5431,N_4553,N_4574);
or U5432 (N_5432,N_4636,N_4904);
nor U5433 (N_5433,N_4634,N_4844);
or U5434 (N_5434,N_4855,N_4582);
nor U5435 (N_5435,N_4764,N_4548);
and U5436 (N_5436,N_4470,N_4920);
xor U5437 (N_5437,N_4939,N_4970);
xor U5438 (N_5438,N_4558,N_4436);
nand U5439 (N_5439,N_4502,N_4732);
xnor U5440 (N_5440,N_4922,N_4784);
xor U5441 (N_5441,N_4639,N_4764);
xor U5442 (N_5442,N_4604,N_4671);
xnor U5443 (N_5443,N_4780,N_4872);
xor U5444 (N_5444,N_4667,N_4379);
and U5445 (N_5445,N_4868,N_4481);
xor U5446 (N_5446,N_4981,N_4698);
nor U5447 (N_5447,N_4870,N_4494);
nand U5448 (N_5448,N_4411,N_4853);
nand U5449 (N_5449,N_4717,N_4475);
nand U5450 (N_5450,N_4949,N_4557);
nand U5451 (N_5451,N_4814,N_4625);
nor U5452 (N_5452,N_4704,N_4531);
nand U5453 (N_5453,N_4832,N_4448);
and U5454 (N_5454,N_4647,N_4790);
nor U5455 (N_5455,N_4621,N_4458);
nand U5456 (N_5456,N_4563,N_4902);
nand U5457 (N_5457,N_4751,N_4994);
or U5458 (N_5458,N_4800,N_4941);
nand U5459 (N_5459,N_4472,N_4723);
nand U5460 (N_5460,N_4394,N_4849);
nor U5461 (N_5461,N_4679,N_4726);
or U5462 (N_5462,N_4735,N_4454);
or U5463 (N_5463,N_4856,N_4798);
xnor U5464 (N_5464,N_4810,N_4890);
and U5465 (N_5465,N_4611,N_4567);
nor U5466 (N_5466,N_4778,N_4532);
nor U5467 (N_5467,N_4756,N_4749);
or U5468 (N_5468,N_4965,N_4835);
nand U5469 (N_5469,N_4581,N_4886);
xnor U5470 (N_5470,N_4892,N_4550);
or U5471 (N_5471,N_4391,N_4481);
nand U5472 (N_5472,N_4950,N_4919);
or U5473 (N_5473,N_4432,N_4849);
xor U5474 (N_5474,N_4531,N_4893);
nand U5475 (N_5475,N_4924,N_4565);
xnor U5476 (N_5476,N_4870,N_4578);
nor U5477 (N_5477,N_4507,N_4630);
nor U5478 (N_5478,N_4755,N_4512);
nor U5479 (N_5479,N_4648,N_4695);
and U5480 (N_5480,N_4383,N_4668);
or U5481 (N_5481,N_4827,N_4445);
xnor U5482 (N_5482,N_4784,N_4761);
or U5483 (N_5483,N_4554,N_4718);
xnor U5484 (N_5484,N_4761,N_4703);
nor U5485 (N_5485,N_4916,N_4820);
nor U5486 (N_5486,N_4884,N_4545);
xnor U5487 (N_5487,N_4486,N_4973);
xor U5488 (N_5488,N_4840,N_4503);
nand U5489 (N_5489,N_4901,N_4511);
xor U5490 (N_5490,N_4510,N_4940);
xnor U5491 (N_5491,N_4445,N_4398);
nor U5492 (N_5492,N_4644,N_4886);
nor U5493 (N_5493,N_4455,N_4928);
nand U5494 (N_5494,N_4516,N_4550);
or U5495 (N_5495,N_4922,N_4872);
and U5496 (N_5496,N_4869,N_4762);
and U5497 (N_5497,N_4821,N_4604);
and U5498 (N_5498,N_4971,N_4965);
nand U5499 (N_5499,N_4433,N_4617);
and U5500 (N_5500,N_4755,N_4429);
or U5501 (N_5501,N_4725,N_4535);
or U5502 (N_5502,N_4578,N_4408);
and U5503 (N_5503,N_4725,N_4532);
and U5504 (N_5504,N_4928,N_4446);
nor U5505 (N_5505,N_4863,N_4706);
or U5506 (N_5506,N_4490,N_4679);
xor U5507 (N_5507,N_4789,N_4481);
or U5508 (N_5508,N_4474,N_4765);
nand U5509 (N_5509,N_4379,N_4616);
or U5510 (N_5510,N_4763,N_4460);
nor U5511 (N_5511,N_4868,N_4967);
nor U5512 (N_5512,N_4594,N_4391);
and U5513 (N_5513,N_4537,N_4752);
nor U5514 (N_5514,N_4765,N_4599);
nand U5515 (N_5515,N_4699,N_4560);
nor U5516 (N_5516,N_4977,N_4899);
xnor U5517 (N_5517,N_4580,N_4656);
xnor U5518 (N_5518,N_4760,N_4986);
nor U5519 (N_5519,N_4722,N_4833);
xor U5520 (N_5520,N_4573,N_4541);
xnor U5521 (N_5521,N_4919,N_4443);
nand U5522 (N_5522,N_4863,N_4771);
or U5523 (N_5523,N_4976,N_4450);
nor U5524 (N_5524,N_4632,N_4448);
xnor U5525 (N_5525,N_4469,N_4630);
and U5526 (N_5526,N_4919,N_4497);
nor U5527 (N_5527,N_4901,N_4833);
or U5528 (N_5528,N_4471,N_4939);
or U5529 (N_5529,N_4618,N_4813);
xor U5530 (N_5530,N_4505,N_4842);
and U5531 (N_5531,N_4863,N_4800);
xor U5532 (N_5532,N_4750,N_4842);
or U5533 (N_5533,N_4476,N_4842);
or U5534 (N_5534,N_4469,N_4933);
nand U5535 (N_5535,N_4515,N_4750);
or U5536 (N_5536,N_4402,N_4463);
or U5537 (N_5537,N_4697,N_4904);
and U5538 (N_5538,N_4399,N_4804);
nor U5539 (N_5539,N_4598,N_4635);
nand U5540 (N_5540,N_4763,N_4406);
xor U5541 (N_5541,N_4581,N_4750);
and U5542 (N_5542,N_4426,N_4663);
and U5543 (N_5543,N_4573,N_4477);
nand U5544 (N_5544,N_4478,N_4489);
and U5545 (N_5545,N_4591,N_4963);
nand U5546 (N_5546,N_4505,N_4899);
and U5547 (N_5547,N_4918,N_4759);
and U5548 (N_5548,N_4651,N_4982);
and U5549 (N_5549,N_4517,N_4691);
or U5550 (N_5550,N_4412,N_4956);
nand U5551 (N_5551,N_4801,N_4445);
or U5552 (N_5552,N_4749,N_4909);
and U5553 (N_5553,N_4760,N_4875);
and U5554 (N_5554,N_4498,N_4999);
nand U5555 (N_5555,N_4816,N_4925);
nand U5556 (N_5556,N_4901,N_4966);
xor U5557 (N_5557,N_4676,N_4992);
xor U5558 (N_5558,N_4856,N_4961);
nor U5559 (N_5559,N_4780,N_4830);
nor U5560 (N_5560,N_4815,N_4478);
nand U5561 (N_5561,N_4381,N_4901);
nand U5562 (N_5562,N_4952,N_4896);
nand U5563 (N_5563,N_4556,N_4480);
and U5564 (N_5564,N_4406,N_4798);
or U5565 (N_5565,N_4506,N_4985);
nand U5566 (N_5566,N_4382,N_4688);
nand U5567 (N_5567,N_4472,N_4528);
nand U5568 (N_5568,N_4891,N_4415);
xnor U5569 (N_5569,N_4676,N_4515);
and U5570 (N_5570,N_4823,N_4763);
xnor U5571 (N_5571,N_4956,N_4668);
and U5572 (N_5572,N_4843,N_4799);
or U5573 (N_5573,N_4803,N_4600);
xor U5574 (N_5574,N_4671,N_4785);
or U5575 (N_5575,N_4667,N_4635);
nand U5576 (N_5576,N_4605,N_4909);
nor U5577 (N_5577,N_4792,N_4430);
and U5578 (N_5578,N_4860,N_4552);
nor U5579 (N_5579,N_4608,N_4491);
and U5580 (N_5580,N_4599,N_4823);
or U5581 (N_5581,N_4645,N_4473);
xor U5582 (N_5582,N_4424,N_4376);
or U5583 (N_5583,N_4437,N_4651);
nor U5584 (N_5584,N_4527,N_4547);
xnor U5585 (N_5585,N_4639,N_4648);
xnor U5586 (N_5586,N_4893,N_4632);
nand U5587 (N_5587,N_4442,N_4824);
or U5588 (N_5588,N_4938,N_4407);
and U5589 (N_5589,N_4931,N_4763);
nand U5590 (N_5590,N_4628,N_4477);
or U5591 (N_5591,N_4791,N_4756);
or U5592 (N_5592,N_4468,N_4654);
nand U5593 (N_5593,N_4505,N_4747);
xor U5594 (N_5594,N_4664,N_4473);
xnor U5595 (N_5595,N_4956,N_4777);
and U5596 (N_5596,N_4643,N_4942);
or U5597 (N_5597,N_4439,N_4749);
nor U5598 (N_5598,N_4398,N_4531);
xor U5599 (N_5599,N_4625,N_4895);
and U5600 (N_5600,N_4550,N_4380);
nor U5601 (N_5601,N_4961,N_4716);
nand U5602 (N_5602,N_4761,N_4521);
and U5603 (N_5603,N_4752,N_4665);
or U5604 (N_5604,N_4419,N_4619);
nand U5605 (N_5605,N_4808,N_4878);
nor U5606 (N_5606,N_4995,N_4879);
nor U5607 (N_5607,N_4636,N_4932);
xnor U5608 (N_5608,N_4810,N_4762);
nand U5609 (N_5609,N_4723,N_4965);
nor U5610 (N_5610,N_4716,N_4645);
nand U5611 (N_5611,N_4884,N_4682);
and U5612 (N_5612,N_4501,N_4478);
nor U5613 (N_5613,N_4525,N_4712);
xor U5614 (N_5614,N_4597,N_4948);
or U5615 (N_5615,N_4886,N_4766);
and U5616 (N_5616,N_4733,N_4707);
nand U5617 (N_5617,N_4679,N_4488);
and U5618 (N_5618,N_4606,N_4905);
nand U5619 (N_5619,N_4669,N_4501);
nand U5620 (N_5620,N_4630,N_4602);
nor U5621 (N_5621,N_4824,N_4956);
and U5622 (N_5622,N_4625,N_4569);
and U5623 (N_5623,N_4431,N_4714);
xnor U5624 (N_5624,N_4678,N_4665);
nor U5625 (N_5625,N_5501,N_5307);
and U5626 (N_5626,N_5418,N_5334);
nor U5627 (N_5627,N_5137,N_5443);
nand U5628 (N_5628,N_5188,N_5160);
nor U5629 (N_5629,N_5030,N_5537);
and U5630 (N_5630,N_5166,N_5571);
nand U5631 (N_5631,N_5405,N_5615);
xor U5632 (N_5632,N_5058,N_5108);
or U5633 (N_5633,N_5584,N_5528);
and U5634 (N_5634,N_5050,N_5134);
xnor U5635 (N_5635,N_5277,N_5083);
nand U5636 (N_5636,N_5290,N_5454);
nor U5637 (N_5637,N_5371,N_5172);
nor U5638 (N_5638,N_5230,N_5269);
nor U5639 (N_5639,N_5060,N_5184);
xnor U5640 (N_5640,N_5171,N_5496);
nor U5641 (N_5641,N_5068,N_5211);
xor U5642 (N_5642,N_5154,N_5310);
nor U5643 (N_5643,N_5262,N_5391);
or U5644 (N_5644,N_5516,N_5471);
or U5645 (N_5645,N_5529,N_5389);
or U5646 (N_5646,N_5604,N_5067);
and U5647 (N_5647,N_5512,N_5005);
nor U5648 (N_5648,N_5382,N_5566);
or U5649 (N_5649,N_5077,N_5093);
nor U5650 (N_5650,N_5255,N_5467);
nand U5651 (N_5651,N_5197,N_5619);
or U5652 (N_5652,N_5161,N_5577);
nand U5653 (N_5653,N_5286,N_5463);
or U5654 (N_5654,N_5522,N_5433);
nor U5655 (N_5655,N_5311,N_5003);
nor U5656 (N_5656,N_5147,N_5044);
nand U5657 (N_5657,N_5547,N_5509);
or U5658 (N_5658,N_5556,N_5056);
nor U5659 (N_5659,N_5373,N_5245);
nand U5660 (N_5660,N_5015,N_5029);
nand U5661 (N_5661,N_5458,N_5102);
nor U5662 (N_5662,N_5561,N_5343);
and U5663 (N_5663,N_5295,N_5357);
nand U5664 (N_5664,N_5612,N_5073);
or U5665 (N_5665,N_5287,N_5316);
nor U5666 (N_5666,N_5545,N_5364);
xor U5667 (N_5667,N_5112,N_5497);
or U5668 (N_5668,N_5169,N_5431);
and U5669 (N_5669,N_5106,N_5588);
xor U5670 (N_5670,N_5623,N_5231);
xor U5671 (N_5671,N_5520,N_5317);
or U5672 (N_5672,N_5449,N_5228);
and U5673 (N_5673,N_5369,N_5439);
nand U5674 (N_5674,N_5204,N_5303);
and U5675 (N_5675,N_5012,N_5246);
or U5676 (N_5676,N_5088,N_5020);
nor U5677 (N_5677,N_5089,N_5616);
nand U5678 (N_5678,N_5129,N_5513);
nor U5679 (N_5679,N_5486,N_5218);
nand U5680 (N_5680,N_5333,N_5367);
nand U5681 (N_5681,N_5091,N_5179);
or U5682 (N_5682,N_5283,N_5581);
or U5683 (N_5683,N_5205,N_5385);
or U5684 (N_5684,N_5592,N_5207);
nor U5685 (N_5685,N_5130,N_5387);
xor U5686 (N_5686,N_5265,N_5315);
nor U5687 (N_5687,N_5063,N_5617);
and U5688 (N_5688,N_5535,N_5476);
or U5689 (N_5689,N_5294,N_5007);
nand U5690 (N_5690,N_5576,N_5229);
nand U5691 (N_5691,N_5271,N_5115);
nor U5692 (N_5692,N_5117,N_5244);
xnor U5693 (N_5693,N_5406,N_5506);
nand U5694 (N_5694,N_5248,N_5087);
and U5695 (N_5695,N_5409,N_5014);
or U5696 (N_5696,N_5480,N_5397);
and U5697 (N_5697,N_5527,N_5505);
nand U5698 (N_5698,N_5420,N_5200);
xor U5699 (N_5699,N_5219,N_5238);
nor U5700 (N_5700,N_5173,N_5376);
nand U5701 (N_5701,N_5125,N_5432);
nor U5702 (N_5702,N_5264,N_5233);
or U5703 (N_5703,N_5323,N_5543);
or U5704 (N_5704,N_5350,N_5043);
nor U5705 (N_5705,N_5157,N_5450);
and U5706 (N_5706,N_5455,N_5393);
nand U5707 (N_5707,N_5209,N_5272);
xor U5708 (N_5708,N_5119,N_5567);
or U5709 (N_5709,N_5440,N_5203);
nand U5710 (N_5710,N_5610,N_5568);
nor U5711 (N_5711,N_5275,N_5314);
nor U5712 (N_5712,N_5324,N_5099);
and U5713 (N_5713,N_5423,N_5611);
xor U5714 (N_5714,N_5589,N_5284);
and U5715 (N_5715,N_5402,N_5168);
and U5716 (N_5716,N_5206,N_5319);
xor U5717 (N_5717,N_5195,N_5252);
xor U5718 (N_5718,N_5494,N_5585);
nor U5719 (N_5719,N_5366,N_5349);
and U5720 (N_5720,N_5025,N_5051);
nand U5721 (N_5721,N_5602,N_5356);
nor U5722 (N_5722,N_5113,N_5490);
or U5723 (N_5723,N_5224,N_5379);
or U5724 (N_5724,N_5123,N_5016);
xor U5725 (N_5725,N_5608,N_5540);
nand U5726 (N_5726,N_5097,N_5404);
or U5727 (N_5727,N_5214,N_5081);
and U5728 (N_5728,N_5413,N_5223);
nor U5729 (N_5729,N_5001,N_5066);
nand U5730 (N_5730,N_5282,N_5293);
xnor U5731 (N_5731,N_5309,N_5473);
or U5732 (N_5732,N_5590,N_5410);
and U5733 (N_5733,N_5217,N_5400);
nor U5734 (N_5734,N_5022,N_5041);
xnor U5735 (N_5735,N_5331,N_5110);
nor U5736 (N_5736,N_5359,N_5504);
nor U5737 (N_5737,N_5484,N_5354);
nand U5738 (N_5738,N_5261,N_5442);
and U5739 (N_5739,N_5419,N_5301);
nand U5740 (N_5740,N_5047,N_5388);
and U5741 (N_5741,N_5470,N_5145);
nor U5742 (N_5742,N_5489,N_5575);
nor U5743 (N_5743,N_5268,N_5136);
xnor U5744 (N_5744,N_5362,N_5361);
or U5745 (N_5745,N_5059,N_5139);
and U5746 (N_5746,N_5142,N_5100);
nand U5747 (N_5747,N_5243,N_5411);
nor U5748 (N_5748,N_5553,N_5459);
xor U5749 (N_5749,N_5472,N_5027);
or U5750 (N_5750,N_5594,N_5267);
or U5751 (N_5751,N_5062,N_5614);
xor U5752 (N_5752,N_5580,N_5126);
and U5753 (N_5753,N_5049,N_5181);
xor U5754 (N_5754,N_5398,N_5260);
nor U5755 (N_5755,N_5500,N_5034);
nand U5756 (N_5756,N_5327,N_5563);
xor U5757 (N_5757,N_5372,N_5201);
or U5758 (N_5758,N_5492,N_5511);
xor U5759 (N_5759,N_5336,N_5039);
and U5760 (N_5760,N_5103,N_5053);
nand U5761 (N_5761,N_5457,N_5010);
or U5762 (N_5762,N_5552,N_5558);
nor U5763 (N_5763,N_5539,N_5150);
or U5764 (N_5764,N_5546,N_5464);
and U5765 (N_5765,N_5559,N_5253);
and U5766 (N_5766,N_5624,N_5210);
xnor U5767 (N_5767,N_5312,N_5291);
nand U5768 (N_5768,N_5479,N_5574);
nor U5769 (N_5769,N_5380,N_5105);
and U5770 (N_5770,N_5326,N_5002);
nor U5771 (N_5771,N_5079,N_5085);
and U5772 (N_5772,N_5163,N_5569);
and U5773 (N_5773,N_5011,N_5198);
xor U5774 (N_5774,N_5435,N_5390);
or U5775 (N_5775,N_5075,N_5325);
nand U5776 (N_5776,N_5257,N_5098);
nor U5777 (N_5777,N_5189,N_5318);
nor U5778 (N_5778,N_5055,N_5477);
nand U5779 (N_5779,N_5221,N_5436);
and U5780 (N_5780,N_5370,N_5330);
xnor U5781 (N_5781,N_5313,N_5453);
nand U5782 (N_5782,N_5235,N_5019);
nor U5783 (N_5783,N_5132,N_5140);
or U5784 (N_5784,N_5560,N_5232);
or U5785 (N_5785,N_5178,N_5242);
and U5786 (N_5786,N_5444,N_5536);
nor U5787 (N_5787,N_5266,N_5321);
xnor U5788 (N_5788,N_5076,N_5036);
nand U5789 (N_5789,N_5202,N_5517);
xnor U5790 (N_5790,N_5368,N_5341);
and U5791 (N_5791,N_5375,N_5107);
and U5792 (N_5792,N_5525,N_5414);
nand U5793 (N_5793,N_5095,N_5222);
or U5794 (N_5794,N_5493,N_5488);
nand U5795 (N_5795,N_5342,N_5510);
or U5796 (N_5796,N_5045,N_5279);
xor U5797 (N_5797,N_5226,N_5254);
nor U5798 (N_5798,N_5057,N_5064);
or U5799 (N_5799,N_5399,N_5466);
and U5800 (N_5800,N_5296,N_5305);
nor U5801 (N_5801,N_5482,N_5445);
or U5802 (N_5802,N_5424,N_5052);
or U5803 (N_5803,N_5587,N_5452);
nor U5804 (N_5804,N_5258,N_5236);
and U5805 (N_5805,N_5109,N_5605);
or U5806 (N_5806,N_5141,N_5417);
xnor U5807 (N_5807,N_5143,N_5220);
and U5808 (N_5808,N_5462,N_5237);
nor U5809 (N_5809,N_5550,N_5241);
xnor U5810 (N_5810,N_5618,N_5596);
nor U5811 (N_5811,N_5074,N_5469);
nand U5812 (N_5812,N_5408,N_5329);
nand U5813 (N_5813,N_5167,N_5508);
xor U5814 (N_5814,N_5365,N_5345);
nor U5815 (N_5815,N_5355,N_5092);
or U5816 (N_5816,N_5381,N_5090);
or U5817 (N_5817,N_5101,N_5118);
nor U5818 (N_5818,N_5430,N_5335);
xor U5819 (N_5819,N_5320,N_5447);
and U5820 (N_5820,N_5149,N_5111);
nor U5821 (N_5821,N_5609,N_5152);
or U5822 (N_5822,N_5146,N_5383);
or U5823 (N_5823,N_5082,N_5583);
nor U5824 (N_5824,N_5384,N_5054);
nor U5825 (N_5825,N_5199,N_5557);
xnor U5826 (N_5826,N_5416,N_5292);
nor U5827 (N_5827,N_5347,N_5565);
nor U5828 (N_5828,N_5395,N_5533);
nand U5829 (N_5829,N_5249,N_5374);
or U5830 (N_5830,N_5351,N_5495);
and U5831 (N_5831,N_5170,N_5532);
xnor U5832 (N_5832,N_5280,N_5586);
or U5833 (N_5833,N_5503,N_5593);
nand U5834 (N_5834,N_5518,N_5175);
or U5835 (N_5835,N_5263,N_5606);
xnor U5836 (N_5836,N_5600,N_5270);
and U5837 (N_5837,N_5234,N_5104);
nor U5838 (N_5838,N_5131,N_5620);
nor U5839 (N_5839,N_5256,N_5212);
xnor U5840 (N_5840,N_5162,N_5274);
and U5841 (N_5841,N_5591,N_5185);
nand U5842 (N_5842,N_5250,N_5412);
or U5843 (N_5843,N_5153,N_5128);
nand U5844 (N_5844,N_5124,N_5299);
xnor U5845 (N_5845,N_5438,N_5194);
xnor U5846 (N_5846,N_5156,N_5065);
or U5847 (N_5847,N_5322,N_5048);
and U5848 (N_5848,N_5499,N_5429);
and U5849 (N_5849,N_5281,N_5352);
and U5850 (N_5850,N_5024,N_5071);
and U5851 (N_5851,N_5216,N_5425);
xor U5852 (N_5852,N_5191,N_5507);
xor U5853 (N_5853,N_5300,N_5038);
and U5854 (N_5854,N_5183,N_5122);
and U5855 (N_5855,N_5302,N_5461);
nand U5856 (N_5856,N_5086,N_5538);
nor U5857 (N_5857,N_5564,N_5096);
nand U5858 (N_5858,N_5483,N_5555);
xnor U5859 (N_5859,N_5013,N_5578);
xnor U5860 (N_5860,N_5164,N_5190);
nand U5861 (N_5861,N_5026,N_5622);
nor U5862 (N_5862,N_5475,N_5225);
xor U5863 (N_5863,N_5534,N_5544);
nor U5864 (N_5864,N_5006,N_5017);
or U5865 (N_5865,N_5415,N_5240);
or U5866 (N_5866,N_5363,N_5530);
nand U5867 (N_5867,N_5155,N_5607);
nand U5868 (N_5868,N_5421,N_5531);
or U5869 (N_5869,N_5403,N_5441);
and U5870 (N_5870,N_5394,N_5159);
xnor U5871 (N_5871,N_5448,N_5332);
xnor U5872 (N_5872,N_5148,N_5009);
nor U5873 (N_5873,N_5046,N_5177);
nand U5874 (N_5874,N_5562,N_5514);
or U5875 (N_5875,N_5524,N_5276);
nand U5876 (N_5876,N_5456,N_5042);
nand U5877 (N_5877,N_5072,N_5526);
and U5878 (N_5878,N_5114,N_5460);
nand U5879 (N_5879,N_5033,N_5288);
and U5880 (N_5880,N_5613,N_5008);
nand U5881 (N_5881,N_5032,N_5344);
nor U5882 (N_5882,N_5599,N_5040);
or U5883 (N_5883,N_5396,N_5521);
and U5884 (N_5884,N_5572,N_5478);
or U5885 (N_5885,N_5196,N_5523);
xor U5886 (N_5886,N_5554,N_5061);
nor U5887 (N_5887,N_5289,N_5037);
or U5888 (N_5888,N_5434,N_5428);
xnor U5889 (N_5889,N_5035,N_5069);
or U5890 (N_5890,N_5031,N_5000);
nand U5891 (N_5891,N_5138,N_5601);
and U5892 (N_5892,N_5621,N_5358);
xnor U5893 (N_5893,N_5481,N_5165);
and U5894 (N_5894,N_5144,N_5116);
and U5895 (N_5895,N_5080,N_5273);
or U5896 (N_5896,N_5018,N_5213);
nand U5897 (N_5897,N_5247,N_5192);
nand U5898 (N_5898,N_5541,N_5515);
or U5899 (N_5899,N_5337,N_5377);
or U5900 (N_5900,N_5422,N_5227);
xor U5901 (N_5901,N_5353,N_5004);
or U5902 (N_5902,N_5186,N_5187);
nand U5903 (N_5903,N_5133,N_5151);
nor U5904 (N_5904,N_5519,N_5597);
xnor U5905 (N_5905,N_5339,N_5392);
nor U5906 (N_5906,N_5251,N_5427);
or U5907 (N_5907,N_5570,N_5127);
nand U5908 (N_5908,N_5378,N_5386);
and U5909 (N_5909,N_5468,N_5603);
or U5910 (N_5910,N_5094,N_5306);
or U5911 (N_5911,N_5437,N_5182);
nand U5912 (N_5912,N_5297,N_5135);
nor U5913 (N_5913,N_5278,N_5340);
xnor U5914 (N_5914,N_5465,N_5028);
xnor U5915 (N_5915,N_5239,N_5582);
or U5916 (N_5916,N_5215,N_5120);
nor U5917 (N_5917,N_5078,N_5498);
and U5918 (N_5918,N_5502,N_5551);
and U5919 (N_5919,N_5598,N_5304);
nand U5920 (N_5920,N_5176,N_5348);
and U5921 (N_5921,N_5485,N_5573);
xnor U5922 (N_5922,N_5360,N_5180);
xor U5923 (N_5923,N_5023,N_5021);
or U5924 (N_5924,N_5298,N_5338);
or U5925 (N_5925,N_5346,N_5285);
nand U5926 (N_5926,N_5308,N_5446);
xnor U5927 (N_5927,N_5474,N_5121);
nand U5928 (N_5928,N_5491,N_5174);
nor U5929 (N_5929,N_5426,N_5451);
nand U5930 (N_5930,N_5542,N_5259);
nor U5931 (N_5931,N_5549,N_5548);
nand U5932 (N_5932,N_5193,N_5401);
or U5933 (N_5933,N_5208,N_5328);
nor U5934 (N_5934,N_5158,N_5084);
nor U5935 (N_5935,N_5595,N_5487);
and U5936 (N_5936,N_5579,N_5407);
and U5937 (N_5937,N_5070,N_5227);
nand U5938 (N_5938,N_5043,N_5042);
or U5939 (N_5939,N_5501,N_5279);
or U5940 (N_5940,N_5116,N_5361);
xor U5941 (N_5941,N_5388,N_5336);
nor U5942 (N_5942,N_5393,N_5160);
or U5943 (N_5943,N_5458,N_5568);
xor U5944 (N_5944,N_5563,N_5256);
or U5945 (N_5945,N_5339,N_5527);
nor U5946 (N_5946,N_5175,N_5448);
or U5947 (N_5947,N_5370,N_5534);
nand U5948 (N_5948,N_5564,N_5038);
xor U5949 (N_5949,N_5477,N_5086);
nand U5950 (N_5950,N_5002,N_5518);
nand U5951 (N_5951,N_5496,N_5573);
or U5952 (N_5952,N_5566,N_5325);
or U5953 (N_5953,N_5021,N_5380);
xor U5954 (N_5954,N_5260,N_5330);
xnor U5955 (N_5955,N_5044,N_5509);
nand U5956 (N_5956,N_5444,N_5181);
or U5957 (N_5957,N_5039,N_5567);
nor U5958 (N_5958,N_5497,N_5039);
nor U5959 (N_5959,N_5003,N_5501);
nor U5960 (N_5960,N_5046,N_5529);
and U5961 (N_5961,N_5308,N_5161);
nor U5962 (N_5962,N_5223,N_5480);
xor U5963 (N_5963,N_5360,N_5370);
xnor U5964 (N_5964,N_5143,N_5337);
nor U5965 (N_5965,N_5107,N_5065);
and U5966 (N_5966,N_5180,N_5449);
nand U5967 (N_5967,N_5355,N_5184);
nor U5968 (N_5968,N_5557,N_5611);
xnor U5969 (N_5969,N_5248,N_5322);
or U5970 (N_5970,N_5290,N_5292);
nor U5971 (N_5971,N_5232,N_5205);
nand U5972 (N_5972,N_5018,N_5486);
and U5973 (N_5973,N_5357,N_5213);
nand U5974 (N_5974,N_5151,N_5588);
xnor U5975 (N_5975,N_5487,N_5211);
nor U5976 (N_5976,N_5265,N_5404);
or U5977 (N_5977,N_5599,N_5149);
nor U5978 (N_5978,N_5546,N_5298);
or U5979 (N_5979,N_5610,N_5370);
and U5980 (N_5980,N_5515,N_5413);
and U5981 (N_5981,N_5581,N_5058);
or U5982 (N_5982,N_5406,N_5263);
xor U5983 (N_5983,N_5311,N_5301);
or U5984 (N_5984,N_5365,N_5001);
nand U5985 (N_5985,N_5534,N_5183);
nand U5986 (N_5986,N_5479,N_5409);
nand U5987 (N_5987,N_5196,N_5602);
or U5988 (N_5988,N_5418,N_5003);
or U5989 (N_5989,N_5252,N_5526);
and U5990 (N_5990,N_5515,N_5029);
nand U5991 (N_5991,N_5459,N_5057);
nor U5992 (N_5992,N_5036,N_5451);
or U5993 (N_5993,N_5621,N_5215);
and U5994 (N_5994,N_5273,N_5508);
nand U5995 (N_5995,N_5243,N_5074);
or U5996 (N_5996,N_5528,N_5145);
and U5997 (N_5997,N_5300,N_5433);
xnor U5998 (N_5998,N_5166,N_5264);
or U5999 (N_5999,N_5111,N_5395);
and U6000 (N_6000,N_5040,N_5124);
and U6001 (N_6001,N_5208,N_5081);
nand U6002 (N_6002,N_5193,N_5499);
nor U6003 (N_6003,N_5531,N_5591);
nor U6004 (N_6004,N_5225,N_5030);
xnor U6005 (N_6005,N_5090,N_5412);
nand U6006 (N_6006,N_5038,N_5486);
xor U6007 (N_6007,N_5140,N_5222);
or U6008 (N_6008,N_5426,N_5032);
nor U6009 (N_6009,N_5367,N_5385);
and U6010 (N_6010,N_5582,N_5143);
nand U6011 (N_6011,N_5171,N_5187);
nor U6012 (N_6012,N_5450,N_5311);
xnor U6013 (N_6013,N_5048,N_5209);
xnor U6014 (N_6014,N_5439,N_5428);
nor U6015 (N_6015,N_5330,N_5229);
and U6016 (N_6016,N_5517,N_5578);
xor U6017 (N_6017,N_5033,N_5026);
xor U6018 (N_6018,N_5033,N_5569);
nand U6019 (N_6019,N_5513,N_5392);
xor U6020 (N_6020,N_5358,N_5196);
xnor U6021 (N_6021,N_5114,N_5622);
xor U6022 (N_6022,N_5186,N_5130);
nor U6023 (N_6023,N_5079,N_5328);
or U6024 (N_6024,N_5123,N_5063);
or U6025 (N_6025,N_5483,N_5413);
and U6026 (N_6026,N_5146,N_5347);
or U6027 (N_6027,N_5016,N_5043);
nor U6028 (N_6028,N_5074,N_5049);
or U6029 (N_6029,N_5145,N_5315);
xor U6030 (N_6030,N_5380,N_5446);
nand U6031 (N_6031,N_5546,N_5058);
nor U6032 (N_6032,N_5614,N_5428);
and U6033 (N_6033,N_5300,N_5485);
nand U6034 (N_6034,N_5432,N_5411);
and U6035 (N_6035,N_5313,N_5547);
and U6036 (N_6036,N_5425,N_5540);
xor U6037 (N_6037,N_5221,N_5162);
or U6038 (N_6038,N_5010,N_5306);
nand U6039 (N_6039,N_5144,N_5246);
nor U6040 (N_6040,N_5341,N_5623);
or U6041 (N_6041,N_5172,N_5554);
or U6042 (N_6042,N_5572,N_5140);
and U6043 (N_6043,N_5584,N_5140);
nand U6044 (N_6044,N_5158,N_5185);
and U6045 (N_6045,N_5373,N_5012);
nand U6046 (N_6046,N_5246,N_5457);
and U6047 (N_6047,N_5210,N_5451);
or U6048 (N_6048,N_5114,N_5140);
nand U6049 (N_6049,N_5550,N_5118);
or U6050 (N_6050,N_5160,N_5550);
nand U6051 (N_6051,N_5491,N_5000);
and U6052 (N_6052,N_5340,N_5276);
nand U6053 (N_6053,N_5282,N_5261);
nor U6054 (N_6054,N_5502,N_5206);
nand U6055 (N_6055,N_5358,N_5406);
or U6056 (N_6056,N_5423,N_5001);
xor U6057 (N_6057,N_5193,N_5576);
nor U6058 (N_6058,N_5263,N_5060);
and U6059 (N_6059,N_5158,N_5117);
nor U6060 (N_6060,N_5439,N_5112);
nand U6061 (N_6061,N_5027,N_5552);
or U6062 (N_6062,N_5260,N_5106);
and U6063 (N_6063,N_5326,N_5393);
and U6064 (N_6064,N_5623,N_5237);
nand U6065 (N_6065,N_5215,N_5059);
nand U6066 (N_6066,N_5090,N_5237);
xor U6067 (N_6067,N_5162,N_5571);
nand U6068 (N_6068,N_5022,N_5515);
xor U6069 (N_6069,N_5142,N_5250);
and U6070 (N_6070,N_5044,N_5454);
or U6071 (N_6071,N_5260,N_5137);
or U6072 (N_6072,N_5064,N_5046);
nor U6073 (N_6073,N_5073,N_5591);
and U6074 (N_6074,N_5591,N_5369);
nor U6075 (N_6075,N_5459,N_5275);
and U6076 (N_6076,N_5259,N_5366);
xnor U6077 (N_6077,N_5278,N_5524);
and U6078 (N_6078,N_5213,N_5143);
or U6079 (N_6079,N_5315,N_5113);
nor U6080 (N_6080,N_5530,N_5487);
or U6081 (N_6081,N_5173,N_5331);
or U6082 (N_6082,N_5522,N_5281);
or U6083 (N_6083,N_5094,N_5257);
nor U6084 (N_6084,N_5239,N_5155);
and U6085 (N_6085,N_5178,N_5415);
or U6086 (N_6086,N_5255,N_5233);
or U6087 (N_6087,N_5132,N_5122);
xor U6088 (N_6088,N_5419,N_5256);
xor U6089 (N_6089,N_5115,N_5559);
and U6090 (N_6090,N_5446,N_5273);
or U6091 (N_6091,N_5059,N_5522);
and U6092 (N_6092,N_5088,N_5033);
or U6093 (N_6093,N_5573,N_5025);
xnor U6094 (N_6094,N_5143,N_5094);
nor U6095 (N_6095,N_5501,N_5622);
nand U6096 (N_6096,N_5033,N_5241);
nor U6097 (N_6097,N_5066,N_5412);
nand U6098 (N_6098,N_5047,N_5111);
xor U6099 (N_6099,N_5605,N_5565);
and U6100 (N_6100,N_5049,N_5477);
nor U6101 (N_6101,N_5360,N_5380);
nand U6102 (N_6102,N_5363,N_5383);
or U6103 (N_6103,N_5521,N_5250);
nor U6104 (N_6104,N_5583,N_5540);
or U6105 (N_6105,N_5236,N_5549);
and U6106 (N_6106,N_5223,N_5317);
nand U6107 (N_6107,N_5487,N_5206);
nor U6108 (N_6108,N_5438,N_5178);
and U6109 (N_6109,N_5146,N_5571);
nor U6110 (N_6110,N_5208,N_5498);
and U6111 (N_6111,N_5218,N_5143);
or U6112 (N_6112,N_5510,N_5151);
and U6113 (N_6113,N_5052,N_5351);
xnor U6114 (N_6114,N_5464,N_5354);
or U6115 (N_6115,N_5570,N_5005);
and U6116 (N_6116,N_5088,N_5604);
or U6117 (N_6117,N_5365,N_5049);
nor U6118 (N_6118,N_5112,N_5450);
nor U6119 (N_6119,N_5489,N_5248);
xnor U6120 (N_6120,N_5381,N_5456);
nor U6121 (N_6121,N_5474,N_5074);
nor U6122 (N_6122,N_5256,N_5329);
nor U6123 (N_6123,N_5066,N_5036);
xor U6124 (N_6124,N_5477,N_5179);
or U6125 (N_6125,N_5097,N_5600);
nor U6126 (N_6126,N_5177,N_5424);
and U6127 (N_6127,N_5202,N_5379);
xor U6128 (N_6128,N_5414,N_5558);
nand U6129 (N_6129,N_5012,N_5077);
or U6130 (N_6130,N_5065,N_5180);
or U6131 (N_6131,N_5181,N_5068);
nand U6132 (N_6132,N_5156,N_5119);
nand U6133 (N_6133,N_5197,N_5029);
nand U6134 (N_6134,N_5560,N_5058);
or U6135 (N_6135,N_5030,N_5253);
or U6136 (N_6136,N_5208,N_5284);
or U6137 (N_6137,N_5161,N_5031);
and U6138 (N_6138,N_5048,N_5308);
and U6139 (N_6139,N_5371,N_5151);
or U6140 (N_6140,N_5611,N_5582);
nor U6141 (N_6141,N_5569,N_5115);
nand U6142 (N_6142,N_5549,N_5046);
nand U6143 (N_6143,N_5082,N_5302);
or U6144 (N_6144,N_5211,N_5311);
xnor U6145 (N_6145,N_5044,N_5345);
and U6146 (N_6146,N_5170,N_5312);
nand U6147 (N_6147,N_5070,N_5321);
xor U6148 (N_6148,N_5060,N_5118);
nand U6149 (N_6149,N_5436,N_5147);
xnor U6150 (N_6150,N_5343,N_5012);
xnor U6151 (N_6151,N_5490,N_5007);
nand U6152 (N_6152,N_5022,N_5250);
xor U6153 (N_6153,N_5491,N_5506);
or U6154 (N_6154,N_5357,N_5145);
and U6155 (N_6155,N_5072,N_5374);
nor U6156 (N_6156,N_5537,N_5037);
nor U6157 (N_6157,N_5354,N_5087);
or U6158 (N_6158,N_5618,N_5394);
or U6159 (N_6159,N_5471,N_5517);
and U6160 (N_6160,N_5399,N_5348);
and U6161 (N_6161,N_5172,N_5618);
nor U6162 (N_6162,N_5151,N_5445);
xor U6163 (N_6163,N_5518,N_5424);
nor U6164 (N_6164,N_5607,N_5293);
or U6165 (N_6165,N_5306,N_5312);
nand U6166 (N_6166,N_5247,N_5101);
or U6167 (N_6167,N_5526,N_5091);
and U6168 (N_6168,N_5511,N_5466);
or U6169 (N_6169,N_5531,N_5292);
xor U6170 (N_6170,N_5047,N_5262);
and U6171 (N_6171,N_5248,N_5136);
xnor U6172 (N_6172,N_5131,N_5534);
nor U6173 (N_6173,N_5029,N_5214);
nor U6174 (N_6174,N_5288,N_5579);
or U6175 (N_6175,N_5264,N_5548);
and U6176 (N_6176,N_5396,N_5448);
nand U6177 (N_6177,N_5045,N_5231);
nor U6178 (N_6178,N_5390,N_5049);
nor U6179 (N_6179,N_5420,N_5365);
or U6180 (N_6180,N_5519,N_5527);
or U6181 (N_6181,N_5458,N_5112);
and U6182 (N_6182,N_5372,N_5551);
nand U6183 (N_6183,N_5201,N_5538);
nor U6184 (N_6184,N_5015,N_5023);
nor U6185 (N_6185,N_5534,N_5032);
or U6186 (N_6186,N_5172,N_5583);
nand U6187 (N_6187,N_5468,N_5384);
or U6188 (N_6188,N_5475,N_5288);
and U6189 (N_6189,N_5062,N_5522);
xnor U6190 (N_6190,N_5469,N_5392);
or U6191 (N_6191,N_5599,N_5368);
and U6192 (N_6192,N_5620,N_5504);
and U6193 (N_6193,N_5014,N_5453);
xor U6194 (N_6194,N_5132,N_5106);
nand U6195 (N_6195,N_5320,N_5146);
nand U6196 (N_6196,N_5274,N_5008);
xor U6197 (N_6197,N_5109,N_5021);
nand U6198 (N_6198,N_5416,N_5036);
nand U6199 (N_6199,N_5113,N_5364);
or U6200 (N_6200,N_5205,N_5099);
nand U6201 (N_6201,N_5113,N_5355);
or U6202 (N_6202,N_5122,N_5226);
or U6203 (N_6203,N_5306,N_5036);
xnor U6204 (N_6204,N_5247,N_5196);
and U6205 (N_6205,N_5186,N_5123);
and U6206 (N_6206,N_5546,N_5436);
xor U6207 (N_6207,N_5422,N_5411);
and U6208 (N_6208,N_5260,N_5072);
nand U6209 (N_6209,N_5565,N_5251);
nor U6210 (N_6210,N_5488,N_5051);
nand U6211 (N_6211,N_5231,N_5240);
nand U6212 (N_6212,N_5465,N_5003);
or U6213 (N_6213,N_5593,N_5186);
nand U6214 (N_6214,N_5413,N_5274);
nand U6215 (N_6215,N_5059,N_5500);
nor U6216 (N_6216,N_5255,N_5424);
and U6217 (N_6217,N_5257,N_5292);
and U6218 (N_6218,N_5150,N_5399);
or U6219 (N_6219,N_5507,N_5462);
xnor U6220 (N_6220,N_5230,N_5321);
xor U6221 (N_6221,N_5022,N_5264);
or U6222 (N_6222,N_5098,N_5570);
nand U6223 (N_6223,N_5576,N_5356);
and U6224 (N_6224,N_5421,N_5487);
or U6225 (N_6225,N_5317,N_5213);
or U6226 (N_6226,N_5365,N_5424);
nand U6227 (N_6227,N_5374,N_5385);
and U6228 (N_6228,N_5015,N_5408);
xnor U6229 (N_6229,N_5441,N_5223);
or U6230 (N_6230,N_5035,N_5019);
and U6231 (N_6231,N_5519,N_5120);
or U6232 (N_6232,N_5297,N_5413);
nand U6233 (N_6233,N_5429,N_5307);
nor U6234 (N_6234,N_5624,N_5162);
and U6235 (N_6235,N_5170,N_5259);
xor U6236 (N_6236,N_5326,N_5253);
and U6237 (N_6237,N_5146,N_5250);
nor U6238 (N_6238,N_5425,N_5236);
and U6239 (N_6239,N_5140,N_5139);
nand U6240 (N_6240,N_5512,N_5041);
or U6241 (N_6241,N_5262,N_5213);
xnor U6242 (N_6242,N_5548,N_5531);
nor U6243 (N_6243,N_5021,N_5118);
nor U6244 (N_6244,N_5541,N_5160);
nor U6245 (N_6245,N_5338,N_5030);
or U6246 (N_6246,N_5394,N_5492);
or U6247 (N_6247,N_5057,N_5242);
xor U6248 (N_6248,N_5153,N_5037);
nand U6249 (N_6249,N_5360,N_5620);
or U6250 (N_6250,N_5723,N_5783);
nand U6251 (N_6251,N_6127,N_5876);
nand U6252 (N_6252,N_6024,N_6055);
nand U6253 (N_6253,N_6005,N_6090);
or U6254 (N_6254,N_5934,N_5720);
or U6255 (N_6255,N_5999,N_6152);
nor U6256 (N_6256,N_6056,N_5691);
and U6257 (N_6257,N_6164,N_5705);
nor U6258 (N_6258,N_5696,N_5669);
and U6259 (N_6259,N_6021,N_5891);
and U6260 (N_6260,N_5693,N_5870);
or U6261 (N_6261,N_6242,N_6129);
nor U6262 (N_6262,N_5814,N_5803);
nand U6263 (N_6263,N_6046,N_5730);
and U6264 (N_6264,N_5648,N_5865);
or U6265 (N_6265,N_6113,N_6205);
and U6266 (N_6266,N_6187,N_5958);
and U6267 (N_6267,N_5875,N_6067);
xnor U6268 (N_6268,N_5949,N_5656);
nor U6269 (N_6269,N_6038,N_5627);
xnor U6270 (N_6270,N_5833,N_5796);
xor U6271 (N_6271,N_5973,N_6176);
nor U6272 (N_6272,N_5802,N_5848);
nor U6273 (N_6273,N_5910,N_6248);
or U6274 (N_6274,N_6206,N_6145);
nand U6275 (N_6275,N_6200,N_5962);
and U6276 (N_6276,N_5840,N_5736);
and U6277 (N_6277,N_5662,N_5681);
nor U6278 (N_6278,N_5727,N_5625);
nand U6279 (N_6279,N_6135,N_6173);
and U6280 (N_6280,N_6226,N_5830);
or U6281 (N_6281,N_6149,N_6202);
and U6282 (N_6282,N_6194,N_5647);
xnor U6283 (N_6283,N_5634,N_6209);
nand U6284 (N_6284,N_5700,N_5852);
xor U6285 (N_6285,N_5786,N_5938);
nor U6286 (N_6286,N_5931,N_5685);
nor U6287 (N_6287,N_6210,N_5998);
or U6288 (N_6288,N_5732,N_5823);
xnor U6289 (N_6289,N_6153,N_5714);
nor U6290 (N_6290,N_5837,N_6156);
and U6291 (N_6291,N_6084,N_6217);
nor U6292 (N_6292,N_5925,N_5935);
and U6293 (N_6293,N_5956,N_6207);
or U6294 (N_6294,N_5992,N_6035);
xnor U6295 (N_6295,N_5944,N_5785);
or U6296 (N_6296,N_6018,N_5930);
and U6297 (N_6297,N_5816,N_5942);
xnor U6298 (N_6298,N_5660,N_5645);
nand U6299 (N_6299,N_6114,N_5960);
nor U6300 (N_6300,N_5804,N_6102);
xnor U6301 (N_6301,N_5879,N_5858);
nor U6302 (N_6302,N_6017,N_5948);
xor U6303 (N_6303,N_6077,N_5912);
nor U6304 (N_6304,N_5906,N_6070);
nor U6305 (N_6305,N_5853,N_5997);
nand U6306 (N_6306,N_5911,N_6150);
and U6307 (N_6307,N_5979,N_6010);
and U6308 (N_6308,N_6109,N_5851);
or U6309 (N_6309,N_6057,N_6146);
nand U6310 (N_6310,N_6094,N_5763);
and U6311 (N_6311,N_5943,N_6096);
xnor U6312 (N_6312,N_6000,N_5933);
nand U6313 (N_6313,N_6116,N_6089);
or U6314 (N_6314,N_5985,N_6105);
xnor U6315 (N_6315,N_6174,N_5702);
xnor U6316 (N_6316,N_6110,N_5764);
nand U6317 (N_6317,N_5754,N_5806);
or U6318 (N_6318,N_6155,N_6015);
and U6319 (N_6319,N_5666,N_6030);
xor U6320 (N_6320,N_6120,N_5982);
or U6321 (N_6321,N_5901,N_6119);
nor U6322 (N_6322,N_6062,N_6061);
and U6323 (N_6323,N_5902,N_5756);
or U6324 (N_6324,N_6185,N_6079);
and U6325 (N_6325,N_6126,N_5686);
xnor U6326 (N_6326,N_5922,N_6182);
nand U6327 (N_6327,N_6212,N_6160);
nand U6328 (N_6328,N_5704,N_5955);
and U6329 (N_6329,N_6128,N_6022);
and U6330 (N_6330,N_5805,N_5829);
and U6331 (N_6331,N_5755,N_5710);
nor U6332 (N_6332,N_5977,N_5887);
nor U6333 (N_6333,N_5845,N_6211);
nand U6334 (N_6334,N_6036,N_6052);
nand U6335 (N_6335,N_5978,N_5984);
or U6336 (N_6336,N_5774,N_5672);
nand U6337 (N_6337,N_6159,N_6072);
or U6338 (N_6338,N_5939,N_6189);
and U6339 (N_6339,N_5863,N_6095);
xor U6340 (N_6340,N_6132,N_6112);
nand U6341 (N_6341,N_6231,N_5919);
or U6342 (N_6342,N_5644,N_5684);
nor U6343 (N_6343,N_5855,N_5991);
nor U6344 (N_6344,N_5993,N_5667);
nand U6345 (N_6345,N_5777,N_6196);
xor U6346 (N_6346,N_5807,N_6007);
xor U6347 (N_6347,N_5798,N_6043);
or U6348 (N_6348,N_5972,N_5729);
nand U6349 (N_6349,N_6151,N_5703);
and U6350 (N_6350,N_6118,N_6004);
nor U6351 (N_6351,N_5753,N_5713);
and U6352 (N_6352,N_5904,N_5626);
and U6353 (N_6353,N_5650,N_5743);
nand U6354 (N_6354,N_6106,N_6012);
xor U6355 (N_6355,N_6184,N_5678);
nor U6356 (N_6356,N_5808,N_6040);
xnor U6357 (N_6357,N_5792,N_5834);
nand U6358 (N_6358,N_6177,N_6029);
or U6359 (N_6359,N_5767,N_5746);
nor U6360 (N_6360,N_6097,N_6162);
or U6361 (N_6361,N_5954,N_5752);
nand U6362 (N_6362,N_6082,N_5768);
and U6363 (N_6363,N_5967,N_5668);
or U6364 (N_6364,N_6002,N_5946);
or U6365 (N_6365,N_5969,N_5638);
or U6366 (N_6366,N_5811,N_5940);
or U6367 (N_6367,N_5828,N_5817);
xnor U6368 (N_6368,N_5988,N_5881);
nor U6369 (N_6369,N_6243,N_5689);
or U6370 (N_6370,N_6193,N_5760);
xnor U6371 (N_6371,N_5968,N_5926);
nor U6372 (N_6372,N_5731,N_6093);
nor U6373 (N_6373,N_6224,N_5923);
nor U6374 (N_6374,N_5788,N_6249);
nand U6375 (N_6375,N_5987,N_6221);
or U6376 (N_6376,N_6228,N_5835);
nand U6377 (N_6377,N_5737,N_5894);
nor U6378 (N_6378,N_6181,N_5945);
nor U6379 (N_6379,N_5712,N_5799);
or U6380 (N_6380,N_5758,N_6108);
and U6381 (N_6381,N_5769,N_5709);
nand U6382 (N_6382,N_5741,N_5632);
or U6383 (N_6383,N_5697,N_6215);
nand U6384 (N_6384,N_5809,N_6175);
nand U6385 (N_6385,N_5655,N_5751);
nor U6386 (N_6386,N_5859,N_5963);
nor U6387 (N_6387,N_6183,N_6075);
nand U6388 (N_6388,N_5916,N_6158);
and U6389 (N_6389,N_5950,N_6219);
nand U6390 (N_6390,N_6186,N_6037);
or U6391 (N_6391,N_5747,N_5952);
xnor U6392 (N_6392,N_5694,N_5740);
nand U6393 (N_6393,N_5790,N_6137);
nand U6394 (N_6394,N_5715,N_5953);
xnor U6395 (N_6395,N_5927,N_6016);
nor U6396 (N_6396,N_5765,N_5826);
or U6397 (N_6397,N_6069,N_6134);
nor U6398 (N_6398,N_6147,N_6086);
nor U6399 (N_6399,N_6195,N_5885);
or U6400 (N_6400,N_5818,N_6063);
and U6401 (N_6401,N_6028,N_6227);
nor U6402 (N_6402,N_6085,N_6081);
or U6403 (N_6403,N_5821,N_5961);
nor U6404 (N_6404,N_5815,N_5716);
xnor U6405 (N_6405,N_6078,N_5895);
nor U6406 (N_6406,N_6019,N_6133);
and U6407 (N_6407,N_5976,N_5628);
xnor U6408 (N_6408,N_5890,N_6051);
xnor U6409 (N_6409,N_6073,N_5812);
or U6410 (N_6410,N_5995,N_6060);
nor U6411 (N_6411,N_6168,N_5914);
nor U6412 (N_6412,N_5996,N_5631);
or U6413 (N_6413,N_6032,N_5841);
nand U6414 (N_6414,N_5639,N_6023);
xnor U6415 (N_6415,N_6033,N_6190);
and U6416 (N_6416,N_6115,N_6154);
nand U6417 (N_6417,N_5917,N_6074);
or U6418 (N_6418,N_5793,N_5728);
nor U6419 (N_6419,N_6098,N_6230);
or U6420 (N_6420,N_6009,N_5750);
nand U6421 (N_6421,N_6122,N_5847);
or U6422 (N_6422,N_6218,N_5913);
xor U6423 (N_6423,N_6234,N_6121);
and U6424 (N_6424,N_6001,N_5937);
nor U6425 (N_6425,N_5775,N_5932);
and U6426 (N_6426,N_5918,N_6008);
nand U6427 (N_6427,N_6191,N_5734);
nor U6428 (N_6428,N_5921,N_5849);
xor U6429 (N_6429,N_5800,N_5908);
or U6430 (N_6430,N_5766,N_5983);
xnor U6431 (N_6431,N_5745,N_5905);
and U6432 (N_6432,N_6042,N_6006);
and U6433 (N_6433,N_5838,N_5883);
nor U6434 (N_6434,N_5770,N_6236);
nor U6435 (N_6435,N_6245,N_5653);
nand U6436 (N_6436,N_6104,N_5857);
nor U6437 (N_6437,N_5773,N_6107);
or U6438 (N_6438,N_5629,N_6144);
or U6439 (N_6439,N_5633,N_6179);
or U6440 (N_6440,N_5687,N_5819);
nor U6441 (N_6441,N_5748,N_6223);
or U6442 (N_6442,N_6161,N_6216);
nand U6443 (N_6443,N_5872,N_6229);
xnor U6444 (N_6444,N_6139,N_6166);
and U6445 (N_6445,N_5794,N_5877);
or U6446 (N_6446,N_6165,N_6148);
and U6447 (N_6447,N_5637,N_6238);
xor U6448 (N_6448,N_5959,N_6232);
xor U6449 (N_6449,N_5903,N_6241);
and U6450 (N_6450,N_6064,N_5665);
and U6451 (N_6451,N_5866,N_6197);
nor U6452 (N_6452,N_5749,N_5843);
nor U6453 (N_6453,N_5896,N_5970);
nor U6454 (N_6454,N_5735,N_5780);
xor U6455 (N_6455,N_5630,N_5974);
or U6456 (N_6456,N_6214,N_6050);
nand U6457 (N_6457,N_5782,N_5941);
nor U6458 (N_6458,N_5886,N_6066);
or U6459 (N_6459,N_6235,N_6034);
or U6460 (N_6460,N_5659,N_6013);
nor U6461 (N_6461,N_6140,N_6014);
xor U6462 (N_6462,N_5893,N_5880);
or U6463 (N_6463,N_5836,N_6053);
or U6464 (N_6464,N_5643,N_5784);
nand U6465 (N_6465,N_5928,N_5701);
nor U6466 (N_6466,N_5965,N_6246);
nor U6467 (N_6467,N_5771,N_5688);
and U6468 (N_6468,N_6020,N_5797);
nor U6469 (N_6469,N_5759,N_5680);
nor U6470 (N_6470,N_6171,N_5873);
and U6471 (N_6471,N_5878,N_5658);
or U6472 (N_6472,N_5695,N_5718);
or U6473 (N_6473,N_5677,N_6141);
nand U6474 (N_6474,N_6092,N_5711);
xnor U6475 (N_6475,N_5690,N_6213);
nand U6476 (N_6476,N_5772,N_6172);
or U6477 (N_6477,N_6011,N_6049);
and U6478 (N_6478,N_6198,N_5721);
nand U6479 (N_6479,N_5980,N_5738);
nand U6480 (N_6480,N_5832,N_6103);
xor U6481 (N_6481,N_6239,N_6025);
or U6482 (N_6482,N_5762,N_6054);
xnor U6483 (N_6483,N_5776,N_5692);
nor U6484 (N_6484,N_6045,N_5661);
and U6485 (N_6485,N_5831,N_5884);
nand U6486 (N_6486,N_5882,N_6048);
and U6487 (N_6487,N_5673,N_5820);
or U6488 (N_6488,N_5664,N_5733);
and U6489 (N_6489,N_5654,N_5867);
or U6490 (N_6490,N_5966,N_5708);
nand U6491 (N_6491,N_5844,N_6225);
and U6492 (N_6492,N_6117,N_5856);
and U6493 (N_6493,N_5957,N_5641);
or U6494 (N_6494,N_6136,N_5929);
or U6495 (N_6495,N_5787,N_5850);
nand U6496 (N_6496,N_5719,N_6111);
nand U6497 (N_6497,N_6220,N_5699);
or U6498 (N_6498,N_6076,N_6091);
nor U6499 (N_6499,N_5824,N_5947);
nand U6500 (N_6500,N_5725,N_5924);
or U6501 (N_6501,N_6027,N_6237);
nor U6502 (N_6502,N_5846,N_6240);
and U6503 (N_6503,N_6041,N_6169);
and U6504 (N_6504,N_5936,N_6167);
xor U6505 (N_6505,N_5869,N_6188);
and U6506 (N_6506,N_5892,N_5683);
and U6507 (N_6507,N_5889,N_6031);
and U6508 (N_6508,N_6192,N_6026);
and U6509 (N_6509,N_6100,N_5971);
nor U6510 (N_6510,N_5674,N_5779);
nor U6511 (N_6511,N_6199,N_6059);
nor U6512 (N_6512,N_5860,N_5676);
nor U6513 (N_6513,N_5964,N_5722);
xor U6514 (N_6514,N_5871,N_5757);
xnor U6515 (N_6515,N_5827,N_5717);
nor U6516 (N_6516,N_6071,N_5920);
or U6517 (N_6517,N_5781,N_6222);
xor U6518 (N_6518,N_5868,N_5742);
or U6519 (N_6519,N_5778,N_5795);
or U6520 (N_6520,N_6208,N_6083);
and U6521 (N_6521,N_5675,N_5989);
xor U6522 (N_6522,N_5679,N_6143);
or U6523 (N_6523,N_5789,N_6080);
xnor U6524 (N_6524,N_6138,N_5975);
nand U6525 (N_6525,N_6157,N_6180);
or U6526 (N_6526,N_5862,N_6087);
or U6527 (N_6527,N_5899,N_5986);
and U6528 (N_6528,N_6044,N_6247);
or U6529 (N_6529,N_6123,N_5813);
and U6530 (N_6530,N_6201,N_5642);
xnor U6531 (N_6531,N_5636,N_5898);
nand U6532 (N_6532,N_5909,N_6101);
xor U6533 (N_6533,N_5663,N_6130);
and U6534 (N_6534,N_5897,N_5726);
and U6535 (N_6535,N_5670,N_5649);
nor U6536 (N_6536,N_5900,N_6170);
nand U6537 (N_6537,N_5640,N_5791);
nor U6538 (N_6538,N_6142,N_5915);
or U6539 (N_6539,N_5839,N_5671);
nor U6540 (N_6540,N_5888,N_5761);
nor U6541 (N_6541,N_5854,N_5861);
nor U6542 (N_6542,N_6068,N_6003);
xnor U6543 (N_6543,N_5739,N_6178);
and U6544 (N_6544,N_5842,N_5994);
or U6545 (N_6545,N_6099,N_5724);
and U6546 (N_6546,N_6244,N_6065);
nand U6547 (N_6547,N_5646,N_5907);
or U6548 (N_6548,N_5706,N_6163);
or U6549 (N_6549,N_6039,N_6058);
nand U6550 (N_6550,N_6088,N_6131);
nand U6551 (N_6551,N_6233,N_5635);
nor U6552 (N_6552,N_5801,N_5744);
nor U6553 (N_6553,N_6204,N_5981);
and U6554 (N_6554,N_5651,N_6124);
or U6555 (N_6555,N_5951,N_6125);
nor U6556 (N_6556,N_5990,N_5652);
and U6557 (N_6557,N_5682,N_5825);
xnor U6558 (N_6558,N_6047,N_5810);
and U6559 (N_6559,N_5864,N_6203);
nor U6560 (N_6560,N_5657,N_5707);
nand U6561 (N_6561,N_5698,N_5822);
or U6562 (N_6562,N_5874,N_5764);
nand U6563 (N_6563,N_5744,N_6212);
and U6564 (N_6564,N_5668,N_5697);
or U6565 (N_6565,N_5989,N_5849);
nand U6566 (N_6566,N_6181,N_6036);
nor U6567 (N_6567,N_5829,N_5966);
and U6568 (N_6568,N_6020,N_6147);
nor U6569 (N_6569,N_6220,N_6179);
nand U6570 (N_6570,N_5707,N_5936);
and U6571 (N_6571,N_6095,N_6092);
xor U6572 (N_6572,N_5928,N_5876);
xor U6573 (N_6573,N_5635,N_6111);
or U6574 (N_6574,N_6057,N_6242);
and U6575 (N_6575,N_5983,N_6000);
nor U6576 (N_6576,N_6141,N_6168);
nor U6577 (N_6577,N_6114,N_5910);
or U6578 (N_6578,N_5644,N_5875);
nor U6579 (N_6579,N_6143,N_6057);
nand U6580 (N_6580,N_6091,N_5674);
nor U6581 (N_6581,N_5766,N_6033);
or U6582 (N_6582,N_6246,N_5861);
nand U6583 (N_6583,N_6249,N_5695);
nor U6584 (N_6584,N_5699,N_6232);
nor U6585 (N_6585,N_5839,N_5953);
nor U6586 (N_6586,N_5693,N_5829);
xnor U6587 (N_6587,N_5767,N_6028);
xnor U6588 (N_6588,N_6164,N_5962);
nand U6589 (N_6589,N_6075,N_6220);
and U6590 (N_6590,N_5656,N_5994);
nor U6591 (N_6591,N_5659,N_5822);
and U6592 (N_6592,N_5865,N_6232);
or U6593 (N_6593,N_6194,N_5838);
nand U6594 (N_6594,N_5957,N_6077);
xor U6595 (N_6595,N_6107,N_5650);
nand U6596 (N_6596,N_5945,N_5662);
or U6597 (N_6597,N_6125,N_5726);
or U6598 (N_6598,N_6214,N_6241);
or U6599 (N_6599,N_6090,N_5985);
nand U6600 (N_6600,N_6065,N_6115);
xor U6601 (N_6601,N_6231,N_5790);
or U6602 (N_6602,N_5724,N_6038);
and U6603 (N_6603,N_6194,N_6140);
nor U6604 (N_6604,N_5943,N_5768);
nor U6605 (N_6605,N_6038,N_5771);
nor U6606 (N_6606,N_5899,N_5840);
and U6607 (N_6607,N_5946,N_6052);
nor U6608 (N_6608,N_6232,N_5660);
and U6609 (N_6609,N_6211,N_5756);
xnor U6610 (N_6610,N_6231,N_6196);
xor U6611 (N_6611,N_5818,N_6041);
nor U6612 (N_6612,N_6025,N_5825);
or U6613 (N_6613,N_5834,N_6063);
or U6614 (N_6614,N_6229,N_6140);
nand U6615 (N_6615,N_5858,N_6193);
xor U6616 (N_6616,N_5856,N_6144);
nor U6617 (N_6617,N_5767,N_6096);
nor U6618 (N_6618,N_5981,N_6161);
or U6619 (N_6619,N_5859,N_6205);
nor U6620 (N_6620,N_6135,N_5971);
or U6621 (N_6621,N_5654,N_5703);
and U6622 (N_6622,N_5893,N_5884);
nor U6623 (N_6623,N_6189,N_5800);
and U6624 (N_6624,N_6200,N_5919);
xnor U6625 (N_6625,N_5707,N_5677);
xnor U6626 (N_6626,N_5819,N_5816);
nand U6627 (N_6627,N_5828,N_5629);
or U6628 (N_6628,N_6122,N_6208);
xor U6629 (N_6629,N_6140,N_5892);
xnor U6630 (N_6630,N_6192,N_6246);
and U6631 (N_6631,N_6030,N_6238);
nand U6632 (N_6632,N_6100,N_6187);
and U6633 (N_6633,N_5658,N_6106);
and U6634 (N_6634,N_5889,N_5707);
nor U6635 (N_6635,N_6109,N_5707);
nor U6636 (N_6636,N_5861,N_6011);
xor U6637 (N_6637,N_5926,N_5692);
xnor U6638 (N_6638,N_6040,N_5633);
xor U6639 (N_6639,N_5962,N_6002);
or U6640 (N_6640,N_5655,N_5657);
nand U6641 (N_6641,N_5740,N_5908);
nor U6642 (N_6642,N_5869,N_5732);
or U6643 (N_6643,N_5657,N_5807);
or U6644 (N_6644,N_5634,N_6104);
nand U6645 (N_6645,N_5883,N_5893);
and U6646 (N_6646,N_6202,N_5915);
or U6647 (N_6647,N_5739,N_5755);
or U6648 (N_6648,N_5940,N_6217);
and U6649 (N_6649,N_6113,N_5942);
nand U6650 (N_6650,N_5763,N_6139);
or U6651 (N_6651,N_5896,N_5917);
nor U6652 (N_6652,N_6177,N_5635);
and U6653 (N_6653,N_5660,N_6146);
and U6654 (N_6654,N_5689,N_6246);
and U6655 (N_6655,N_5790,N_5907);
nand U6656 (N_6656,N_5768,N_5712);
and U6657 (N_6657,N_5821,N_5736);
nand U6658 (N_6658,N_5730,N_5701);
or U6659 (N_6659,N_6193,N_6081);
nor U6660 (N_6660,N_5701,N_5947);
xnor U6661 (N_6661,N_5726,N_5712);
and U6662 (N_6662,N_5877,N_6104);
or U6663 (N_6663,N_6200,N_5809);
nor U6664 (N_6664,N_6098,N_5917);
and U6665 (N_6665,N_5718,N_5966);
and U6666 (N_6666,N_6070,N_5640);
nor U6667 (N_6667,N_5925,N_5948);
xor U6668 (N_6668,N_5766,N_6055);
or U6669 (N_6669,N_6202,N_6020);
and U6670 (N_6670,N_5952,N_5742);
or U6671 (N_6671,N_5809,N_6174);
and U6672 (N_6672,N_5788,N_6105);
nand U6673 (N_6673,N_5715,N_6046);
or U6674 (N_6674,N_5709,N_5972);
nand U6675 (N_6675,N_5719,N_6087);
or U6676 (N_6676,N_5975,N_6166);
or U6677 (N_6677,N_5761,N_6010);
and U6678 (N_6678,N_5657,N_5803);
nor U6679 (N_6679,N_5645,N_5869);
nor U6680 (N_6680,N_5802,N_5844);
nor U6681 (N_6681,N_5825,N_6032);
xor U6682 (N_6682,N_6182,N_5778);
or U6683 (N_6683,N_5868,N_6167);
or U6684 (N_6684,N_5727,N_5649);
nor U6685 (N_6685,N_6196,N_5804);
xnor U6686 (N_6686,N_5859,N_6071);
nor U6687 (N_6687,N_5971,N_6112);
nor U6688 (N_6688,N_6068,N_5837);
xor U6689 (N_6689,N_5640,N_6117);
or U6690 (N_6690,N_6086,N_6229);
and U6691 (N_6691,N_5930,N_5906);
and U6692 (N_6692,N_5869,N_6050);
nand U6693 (N_6693,N_5903,N_6187);
nand U6694 (N_6694,N_6039,N_5936);
nand U6695 (N_6695,N_6094,N_5650);
xnor U6696 (N_6696,N_5846,N_5663);
xnor U6697 (N_6697,N_5677,N_5911);
nand U6698 (N_6698,N_5961,N_5776);
and U6699 (N_6699,N_6158,N_6121);
or U6700 (N_6700,N_6188,N_5661);
nor U6701 (N_6701,N_6037,N_6182);
and U6702 (N_6702,N_6241,N_5649);
and U6703 (N_6703,N_6157,N_5860);
or U6704 (N_6704,N_6241,N_6044);
nand U6705 (N_6705,N_6043,N_6004);
xor U6706 (N_6706,N_5918,N_6136);
xor U6707 (N_6707,N_5851,N_5630);
nor U6708 (N_6708,N_5654,N_5798);
or U6709 (N_6709,N_5994,N_5805);
nand U6710 (N_6710,N_6097,N_5712);
or U6711 (N_6711,N_5802,N_5943);
and U6712 (N_6712,N_6218,N_5625);
or U6713 (N_6713,N_5673,N_5941);
nor U6714 (N_6714,N_6190,N_6063);
nor U6715 (N_6715,N_5713,N_5672);
nand U6716 (N_6716,N_6073,N_5659);
and U6717 (N_6717,N_5880,N_6223);
nand U6718 (N_6718,N_5626,N_6128);
and U6719 (N_6719,N_6061,N_5772);
nand U6720 (N_6720,N_5951,N_5851);
and U6721 (N_6721,N_5769,N_5687);
nor U6722 (N_6722,N_6240,N_6122);
and U6723 (N_6723,N_5894,N_5996);
nor U6724 (N_6724,N_5817,N_5683);
or U6725 (N_6725,N_5827,N_6135);
nand U6726 (N_6726,N_6055,N_5913);
nand U6727 (N_6727,N_6210,N_6144);
xor U6728 (N_6728,N_6023,N_6117);
xor U6729 (N_6729,N_5664,N_5679);
and U6730 (N_6730,N_5931,N_5692);
or U6731 (N_6731,N_5968,N_5689);
xor U6732 (N_6732,N_6127,N_5901);
or U6733 (N_6733,N_6058,N_6164);
nand U6734 (N_6734,N_5728,N_5919);
nor U6735 (N_6735,N_5670,N_5919);
or U6736 (N_6736,N_6023,N_5818);
nand U6737 (N_6737,N_5865,N_5988);
nand U6738 (N_6738,N_5859,N_5682);
or U6739 (N_6739,N_5707,N_6194);
or U6740 (N_6740,N_5891,N_5946);
or U6741 (N_6741,N_5796,N_5812);
nor U6742 (N_6742,N_6181,N_6241);
nand U6743 (N_6743,N_5678,N_6187);
nand U6744 (N_6744,N_5964,N_5841);
xnor U6745 (N_6745,N_5871,N_5640);
or U6746 (N_6746,N_5837,N_6170);
and U6747 (N_6747,N_6236,N_6230);
and U6748 (N_6748,N_5921,N_5880);
or U6749 (N_6749,N_5766,N_5850);
nor U6750 (N_6750,N_5884,N_5984);
or U6751 (N_6751,N_5793,N_5736);
nor U6752 (N_6752,N_5806,N_6061);
nor U6753 (N_6753,N_6105,N_6039);
nor U6754 (N_6754,N_6142,N_5774);
nand U6755 (N_6755,N_6129,N_5645);
and U6756 (N_6756,N_6230,N_5739);
xor U6757 (N_6757,N_6051,N_5948);
and U6758 (N_6758,N_6217,N_5784);
xnor U6759 (N_6759,N_6023,N_5672);
nor U6760 (N_6760,N_6196,N_6225);
nand U6761 (N_6761,N_6139,N_5810);
nor U6762 (N_6762,N_6217,N_5797);
nor U6763 (N_6763,N_6037,N_6146);
and U6764 (N_6764,N_5932,N_5804);
and U6765 (N_6765,N_5747,N_6002);
nor U6766 (N_6766,N_5832,N_5865);
or U6767 (N_6767,N_5667,N_6041);
or U6768 (N_6768,N_6118,N_6149);
xor U6769 (N_6769,N_6115,N_5827);
nand U6770 (N_6770,N_6075,N_5652);
nand U6771 (N_6771,N_5830,N_6186);
nor U6772 (N_6772,N_6237,N_5769);
nor U6773 (N_6773,N_6143,N_5983);
and U6774 (N_6774,N_6232,N_6197);
nand U6775 (N_6775,N_6082,N_5685);
or U6776 (N_6776,N_5889,N_5864);
xor U6777 (N_6777,N_6096,N_5868);
or U6778 (N_6778,N_5695,N_5947);
nor U6779 (N_6779,N_6177,N_5906);
nor U6780 (N_6780,N_6179,N_6169);
or U6781 (N_6781,N_6044,N_6210);
or U6782 (N_6782,N_5725,N_5994);
and U6783 (N_6783,N_6193,N_5786);
and U6784 (N_6784,N_5645,N_6168);
xor U6785 (N_6785,N_6040,N_6113);
or U6786 (N_6786,N_5693,N_5733);
nor U6787 (N_6787,N_6037,N_5770);
xor U6788 (N_6788,N_5718,N_5769);
nand U6789 (N_6789,N_5876,N_5819);
nand U6790 (N_6790,N_6221,N_5687);
and U6791 (N_6791,N_6000,N_5673);
nand U6792 (N_6792,N_6136,N_5685);
xnor U6793 (N_6793,N_5768,N_5825);
xnor U6794 (N_6794,N_6082,N_5679);
nor U6795 (N_6795,N_5982,N_5888);
nor U6796 (N_6796,N_5870,N_5710);
nand U6797 (N_6797,N_6036,N_5775);
xor U6798 (N_6798,N_6086,N_5732);
nand U6799 (N_6799,N_5631,N_6019);
xor U6800 (N_6800,N_5634,N_5691);
nand U6801 (N_6801,N_5920,N_5747);
nand U6802 (N_6802,N_5715,N_6114);
or U6803 (N_6803,N_6083,N_5994);
nor U6804 (N_6804,N_5682,N_5766);
xnor U6805 (N_6805,N_6219,N_5974);
or U6806 (N_6806,N_5786,N_6077);
xor U6807 (N_6807,N_6131,N_6243);
xor U6808 (N_6808,N_6193,N_5826);
and U6809 (N_6809,N_6142,N_6014);
or U6810 (N_6810,N_5973,N_5755);
xor U6811 (N_6811,N_5979,N_5995);
nand U6812 (N_6812,N_6006,N_5772);
nand U6813 (N_6813,N_5736,N_6132);
nor U6814 (N_6814,N_6181,N_6040);
nand U6815 (N_6815,N_5679,N_5862);
and U6816 (N_6816,N_5806,N_5640);
or U6817 (N_6817,N_5917,N_6126);
and U6818 (N_6818,N_6056,N_6143);
or U6819 (N_6819,N_6141,N_6032);
nor U6820 (N_6820,N_6077,N_6150);
nand U6821 (N_6821,N_5877,N_5823);
nor U6822 (N_6822,N_6210,N_6134);
nor U6823 (N_6823,N_5626,N_5860);
or U6824 (N_6824,N_5816,N_5727);
or U6825 (N_6825,N_6153,N_5805);
nand U6826 (N_6826,N_5633,N_6171);
or U6827 (N_6827,N_5842,N_6195);
and U6828 (N_6828,N_5849,N_5959);
and U6829 (N_6829,N_6074,N_5818);
nand U6830 (N_6830,N_6126,N_6078);
nor U6831 (N_6831,N_5723,N_5631);
or U6832 (N_6832,N_5721,N_5840);
or U6833 (N_6833,N_5741,N_6067);
nor U6834 (N_6834,N_6249,N_5893);
nor U6835 (N_6835,N_5865,N_5926);
nand U6836 (N_6836,N_5742,N_6112);
nand U6837 (N_6837,N_5628,N_5988);
and U6838 (N_6838,N_5817,N_5908);
or U6839 (N_6839,N_6029,N_5959);
and U6840 (N_6840,N_5911,N_6137);
or U6841 (N_6841,N_6038,N_6170);
nor U6842 (N_6842,N_6165,N_5780);
nor U6843 (N_6843,N_6142,N_6190);
and U6844 (N_6844,N_6164,N_5765);
nand U6845 (N_6845,N_6182,N_5773);
xnor U6846 (N_6846,N_5857,N_5933);
or U6847 (N_6847,N_5854,N_5896);
xor U6848 (N_6848,N_5790,N_5636);
or U6849 (N_6849,N_5702,N_5626);
xnor U6850 (N_6850,N_5688,N_6014);
nand U6851 (N_6851,N_5760,N_5767);
or U6852 (N_6852,N_5996,N_6056);
nor U6853 (N_6853,N_5740,N_5760);
and U6854 (N_6854,N_5654,N_6058);
xnor U6855 (N_6855,N_5729,N_5655);
xor U6856 (N_6856,N_5697,N_5903);
or U6857 (N_6857,N_6043,N_5742);
xnor U6858 (N_6858,N_6005,N_5925);
or U6859 (N_6859,N_6094,N_5775);
or U6860 (N_6860,N_6112,N_5984);
and U6861 (N_6861,N_5984,N_6114);
and U6862 (N_6862,N_5649,N_5860);
xnor U6863 (N_6863,N_6215,N_5682);
or U6864 (N_6864,N_5633,N_6226);
xor U6865 (N_6865,N_6228,N_5805);
xor U6866 (N_6866,N_5648,N_6020);
and U6867 (N_6867,N_5702,N_5766);
xor U6868 (N_6868,N_5780,N_6005);
xnor U6869 (N_6869,N_5635,N_6223);
nor U6870 (N_6870,N_5661,N_5644);
nor U6871 (N_6871,N_5910,N_6125);
or U6872 (N_6872,N_6127,N_6123);
nand U6873 (N_6873,N_6055,N_6089);
and U6874 (N_6874,N_5964,N_5830);
or U6875 (N_6875,N_6619,N_6579);
nand U6876 (N_6876,N_6338,N_6251);
xor U6877 (N_6877,N_6743,N_6637);
xnor U6878 (N_6878,N_6404,N_6826);
nand U6879 (N_6879,N_6312,N_6327);
xnor U6880 (N_6880,N_6700,N_6279);
xor U6881 (N_6881,N_6724,N_6368);
nand U6882 (N_6882,N_6559,N_6446);
nand U6883 (N_6883,N_6361,N_6314);
nor U6884 (N_6884,N_6523,N_6773);
nor U6885 (N_6885,N_6252,N_6692);
or U6886 (N_6886,N_6319,N_6278);
nor U6887 (N_6887,N_6854,N_6767);
or U6888 (N_6888,N_6782,N_6736);
or U6889 (N_6889,N_6483,N_6396);
nand U6890 (N_6890,N_6676,N_6682);
nor U6891 (N_6891,N_6405,N_6495);
nor U6892 (N_6892,N_6778,N_6617);
nor U6893 (N_6893,N_6250,N_6413);
xnor U6894 (N_6894,N_6459,N_6719);
and U6895 (N_6895,N_6273,N_6674);
and U6896 (N_6896,N_6584,N_6397);
and U6897 (N_6897,N_6803,N_6695);
nor U6898 (N_6898,N_6522,N_6355);
xor U6899 (N_6899,N_6783,N_6705);
xor U6900 (N_6900,N_6277,N_6411);
xnor U6901 (N_6901,N_6613,N_6565);
nand U6902 (N_6902,N_6557,N_6722);
and U6903 (N_6903,N_6393,N_6553);
nor U6904 (N_6904,N_6332,N_6640);
xor U6905 (N_6905,N_6482,N_6437);
xor U6906 (N_6906,N_6341,N_6632);
nor U6907 (N_6907,N_6606,N_6721);
nand U6908 (N_6908,N_6690,N_6823);
and U6909 (N_6909,N_6474,N_6763);
or U6910 (N_6910,N_6696,N_6463);
nand U6911 (N_6911,N_6345,N_6321);
xnor U6912 (N_6912,N_6627,N_6386);
and U6913 (N_6913,N_6631,N_6587);
or U6914 (N_6914,N_6264,N_6287);
and U6915 (N_6915,N_6869,N_6518);
nand U6916 (N_6916,N_6745,N_6753);
nor U6917 (N_6917,N_6381,N_6353);
xor U6918 (N_6918,N_6786,N_6612);
nand U6919 (N_6919,N_6816,N_6485);
nor U6920 (N_6920,N_6284,N_6552);
nor U6921 (N_6921,N_6646,N_6357);
nor U6922 (N_6922,N_6817,N_6666);
xnor U6923 (N_6923,N_6863,N_6830);
nor U6924 (N_6924,N_6591,N_6625);
and U6925 (N_6925,N_6293,N_6644);
xor U6926 (N_6926,N_6515,N_6349);
or U6927 (N_6927,N_6257,N_6762);
and U6928 (N_6928,N_6384,N_6311);
nand U6929 (N_6929,N_6813,N_6316);
nand U6930 (N_6930,N_6797,N_6514);
and U6931 (N_6931,N_6756,N_6383);
nor U6932 (N_6932,N_6603,N_6294);
nand U6933 (N_6933,N_6271,N_6575);
nand U6934 (N_6934,N_6549,N_6734);
xor U6935 (N_6935,N_6828,N_6671);
and U6936 (N_6936,N_6716,N_6537);
and U6937 (N_6937,N_6390,N_6687);
xor U6938 (N_6938,N_6595,N_6457);
or U6939 (N_6939,N_6333,N_6852);
or U6940 (N_6940,N_6633,N_6744);
and U6941 (N_6941,N_6620,N_6290);
and U6942 (N_6942,N_6585,N_6313);
nor U6943 (N_6943,N_6471,N_6793);
and U6944 (N_6944,N_6425,N_6706);
or U6945 (N_6945,N_6461,N_6503);
nand U6946 (N_6946,N_6299,N_6592);
or U6947 (N_6947,N_6403,N_6505);
xnor U6948 (N_6948,N_6310,N_6649);
nor U6949 (N_6949,N_6412,N_6426);
nor U6950 (N_6950,N_6328,N_6476);
nor U6951 (N_6951,N_6608,N_6511);
and U6952 (N_6952,N_6547,N_6848);
xnor U6953 (N_6953,N_6697,N_6442);
or U6954 (N_6954,N_6845,N_6540);
nor U6955 (N_6955,N_6406,N_6647);
or U6956 (N_6956,N_6422,N_6473);
nor U6957 (N_6957,N_6401,N_6266);
and U6958 (N_6958,N_6544,N_6868);
nand U6959 (N_6959,N_6610,N_6415);
xnor U6960 (N_6960,N_6851,N_6253);
xnor U6961 (N_6961,N_6770,N_6739);
nand U6962 (N_6962,N_6691,N_6846);
or U6963 (N_6963,N_6533,N_6833);
nand U6964 (N_6964,N_6624,N_6513);
or U6965 (N_6965,N_6410,N_6499);
nor U6966 (N_6966,N_6556,N_6408);
or U6967 (N_6967,N_6811,N_6815);
xnor U6968 (N_6968,N_6254,N_6551);
or U6969 (N_6969,N_6481,N_6870);
xor U6970 (N_6970,N_6267,N_6701);
xnor U6971 (N_6971,N_6433,N_6329);
and U6972 (N_6972,N_6545,N_6789);
or U6973 (N_6973,N_6430,N_6605);
and U6974 (N_6974,N_6360,N_6638);
xnor U6975 (N_6975,N_6356,N_6344);
or U6976 (N_6976,N_6454,N_6806);
nand U6977 (N_6977,N_6458,N_6301);
or U6978 (N_6978,N_6787,N_6658);
or U6979 (N_6979,N_6704,N_6759);
and U6980 (N_6980,N_6414,N_6801);
or U6981 (N_6981,N_6521,N_6867);
nor U6982 (N_6982,N_6827,N_6634);
nor U6983 (N_6983,N_6296,N_6307);
or U6984 (N_6984,N_6643,N_6785);
nor U6985 (N_6985,N_6836,N_6864);
nor U6986 (N_6986,N_6302,N_6661);
xor U6987 (N_6987,N_6470,N_6859);
or U6988 (N_6988,N_6717,N_6711);
or U6989 (N_6989,N_6564,N_6766);
and U6990 (N_6990,N_6378,N_6400);
nand U6991 (N_6991,N_6621,N_6407);
xnor U6992 (N_6992,N_6385,N_6370);
nand U6993 (N_6993,N_6501,N_6727);
or U6994 (N_6994,N_6326,N_6657);
or U6995 (N_6995,N_6256,N_6478);
and U6996 (N_6996,N_6465,N_6375);
and U6997 (N_6997,N_6583,N_6754);
nand U6998 (N_6998,N_6436,N_6519);
and U6999 (N_6999,N_6576,N_6616);
nor U7000 (N_7000,N_6441,N_6315);
xor U7001 (N_7001,N_6512,N_6291);
and U7002 (N_7002,N_6466,N_6298);
or U7003 (N_7003,N_6642,N_6364);
nand U7004 (N_7004,N_6568,N_6418);
nand U7005 (N_7005,N_6784,N_6340);
and U7006 (N_7006,N_6261,N_6856);
xnor U7007 (N_7007,N_6377,N_6731);
and U7008 (N_7008,N_6835,N_6681);
nor U7009 (N_7009,N_6601,N_6765);
xor U7010 (N_7010,N_6652,N_6812);
xor U7011 (N_7011,N_6774,N_6350);
xnor U7012 (N_7012,N_6325,N_6506);
and U7013 (N_7013,N_6358,N_6672);
xor U7014 (N_7014,N_6761,N_6392);
or U7015 (N_7015,N_6680,N_6703);
nor U7016 (N_7016,N_6376,N_6740);
or U7017 (N_7017,N_6309,N_6343);
and U7018 (N_7018,N_6460,N_6710);
xor U7019 (N_7019,N_6464,N_6831);
nor U7020 (N_7020,N_6487,N_6494);
and U7021 (N_7021,N_6819,N_6504);
nand U7022 (N_7022,N_6694,N_6546);
xnor U7023 (N_7023,N_6262,N_6594);
nor U7024 (N_7024,N_6354,N_6741);
and U7025 (N_7025,N_6423,N_6555);
or U7026 (N_7026,N_6873,N_6623);
nor U7027 (N_7027,N_6373,N_6771);
nor U7028 (N_7028,N_6498,N_6853);
nor U7029 (N_7029,N_6489,N_6434);
and U7030 (N_7030,N_6821,N_6604);
or U7031 (N_7031,N_6825,N_6602);
nor U7032 (N_7032,N_6858,N_6500);
nand U7033 (N_7033,N_6820,N_6348);
xor U7034 (N_7034,N_6685,N_6398);
nor U7035 (N_7035,N_6807,N_6342);
nor U7036 (N_7036,N_6574,N_6662);
xnor U7037 (N_7037,N_6752,N_6626);
nand U7038 (N_7038,N_6597,N_6496);
nor U7039 (N_7039,N_6746,N_6804);
and U7040 (N_7040,N_6280,N_6683);
nand U7041 (N_7041,N_6432,N_6805);
and U7042 (N_7042,N_6654,N_6862);
and U7043 (N_7043,N_6281,N_6802);
nand U7044 (N_7044,N_6538,N_6686);
and U7045 (N_7045,N_6269,N_6656);
or U7046 (N_7046,N_6558,N_6331);
or U7047 (N_7047,N_6444,N_6380);
and U7048 (N_7048,N_6794,N_6611);
or U7049 (N_7049,N_6668,N_6490);
or U7050 (N_7050,N_6855,N_6600);
xnor U7051 (N_7051,N_6607,N_6693);
nor U7052 (N_7052,N_6258,N_6352);
nand U7053 (N_7053,N_6834,N_6286);
and U7054 (N_7054,N_6677,N_6292);
xnor U7055 (N_7055,N_6561,N_6359);
and U7056 (N_7056,N_6288,N_6779);
nand U7057 (N_7057,N_6861,N_6289);
nand U7058 (N_7058,N_6275,N_6709);
nand U7059 (N_7059,N_6543,N_6324);
xor U7060 (N_7060,N_6362,N_6502);
and U7061 (N_7061,N_6857,N_6837);
nand U7062 (N_7062,N_6645,N_6394);
xor U7063 (N_7063,N_6492,N_6810);
or U7064 (N_7064,N_6829,N_6443);
and U7065 (N_7065,N_6702,N_6484);
and U7066 (N_7066,N_6548,N_6651);
nor U7067 (N_7067,N_6630,N_6667);
nor U7068 (N_7068,N_6790,N_6566);
or U7069 (N_7069,N_6849,N_6550);
nand U7070 (N_7070,N_6712,N_6757);
nor U7071 (N_7071,N_6416,N_6532);
or U7072 (N_7072,N_6791,N_6578);
or U7073 (N_7073,N_6588,N_6480);
xor U7074 (N_7074,N_6822,N_6402);
or U7075 (N_7075,N_6844,N_6263);
and U7076 (N_7076,N_6509,N_6795);
nand U7077 (N_7077,N_6334,N_6814);
or U7078 (N_7078,N_6641,N_6788);
and U7079 (N_7079,N_6590,N_6516);
xor U7080 (N_7080,N_6429,N_6320);
nand U7081 (N_7081,N_6563,N_6527);
and U7082 (N_7082,N_6776,N_6809);
xor U7083 (N_7083,N_6818,N_6379);
nand U7084 (N_7084,N_6589,N_6367);
xnor U7085 (N_7085,N_6530,N_6768);
nor U7086 (N_7086,N_6421,N_6792);
xnor U7087 (N_7087,N_6477,N_6475);
nor U7088 (N_7088,N_6282,N_6615);
or U7089 (N_7089,N_6308,N_6259);
or U7090 (N_7090,N_6488,N_6554);
xor U7091 (N_7091,N_6562,N_6526);
nor U7092 (N_7092,N_6420,N_6874);
xor U7093 (N_7093,N_6391,N_6469);
nand U7094 (N_7094,N_6387,N_6336);
or U7095 (N_7095,N_6775,N_6268);
and U7096 (N_7096,N_6655,N_6467);
and U7097 (N_7097,N_6593,N_6346);
nand U7098 (N_7098,N_6560,N_6684);
nand U7099 (N_7099,N_6541,N_6614);
nand U7100 (N_7100,N_6586,N_6582);
nor U7101 (N_7101,N_6427,N_6824);
nor U7102 (N_7102,N_6318,N_6440);
xnor U7103 (N_7103,N_6599,N_6742);
or U7104 (N_7104,N_6699,N_6872);
and U7105 (N_7105,N_6339,N_6525);
nand U7106 (N_7106,N_6388,N_6628);
nor U7107 (N_7107,N_6758,N_6842);
xor U7108 (N_7108,N_6839,N_6729);
nor U7109 (N_7109,N_6274,N_6725);
nor U7110 (N_7110,N_6735,N_6520);
nand U7111 (N_7111,N_6718,N_6363);
nand U7112 (N_7112,N_6660,N_6629);
or U7113 (N_7113,N_6351,N_6428);
nor U7114 (N_7114,N_6777,N_6322);
xnor U7115 (N_7115,N_6297,N_6295);
nor U7116 (N_7116,N_6581,N_6799);
nor U7117 (N_7117,N_6452,N_6573);
nor U7118 (N_7118,N_6542,N_6369);
and U7119 (N_7119,N_6409,N_6276);
and U7120 (N_7120,N_6843,N_6664);
xnor U7121 (N_7121,N_6335,N_6838);
and U7122 (N_7122,N_6365,N_6455);
nor U7123 (N_7123,N_6439,N_6860);
nor U7124 (N_7124,N_6708,N_6663);
and U7125 (N_7125,N_6260,N_6323);
or U7126 (N_7126,N_6283,N_6372);
or U7127 (N_7127,N_6737,N_6535);
nand U7128 (N_7128,N_6678,N_6720);
and U7129 (N_7129,N_6781,N_6635);
nand U7130 (N_7130,N_6508,N_6751);
nor U7131 (N_7131,N_6572,N_6749);
and U7132 (N_7132,N_6723,N_6534);
xnor U7133 (N_7133,N_6726,N_6531);
nand U7134 (N_7134,N_6265,N_6389);
and U7135 (N_7135,N_6347,N_6486);
and U7136 (N_7136,N_6650,N_6462);
nand U7137 (N_7137,N_6636,N_6435);
or U7138 (N_7138,N_6445,N_6417);
xnor U7139 (N_7139,N_6732,N_6317);
and U7140 (N_7140,N_6300,N_6303);
and U7141 (N_7141,N_6688,N_6448);
and U7142 (N_7142,N_6728,N_6598);
xor U7143 (N_7143,N_6707,N_6395);
or U7144 (N_7144,N_6528,N_6539);
nand U7145 (N_7145,N_6780,N_6468);
nor U7146 (N_7146,N_6800,N_6639);
or U7147 (N_7147,N_6510,N_6399);
xnor U7148 (N_7148,N_6738,N_6374);
or U7149 (N_7149,N_6330,N_6497);
and U7150 (N_7150,N_6796,N_6456);
nor U7151 (N_7151,N_6733,N_6772);
nand U7152 (N_7152,N_6747,N_6306);
nand U7153 (N_7153,N_6491,N_6865);
nand U7154 (N_7154,N_6272,N_6750);
xnor U7155 (N_7155,N_6648,N_6285);
nor U7156 (N_7156,N_6669,N_6713);
xor U7157 (N_7157,N_6659,N_6507);
and U7158 (N_7158,N_6580,N_6517);
or U7159 (N_7159,N_6755,N_6438);
nor U7160 (N_7160,N_6769,N_6840);
and U7161 (N_7161,N_6596,N_6567);
and U7162 (N_7162,N_6424,N_6764);
xnor U7163 (N_7163,N_6479,N_6670);
or U7164 (N_7164,N_6337,N_6715);
and U7165 (N_7165,N_6451,N_6431);
xor U7166 (N_7166,N_6529,N_6832);
nor U7167 (N_7167,N_6730,N_6665);
nand U7168 (N_7168,N_6371,N_6675);
xnor U7169 (N_7169,N_6571,N_6673);
xnor U7170 (N_7170,N_6305,N_6577);
or U7171 (N_7171,N_6798,N_6453);
and U7172 (N_7172,N_6847,N_6493);
nand U7173 (N_7173,N_6689,N_6866);
or U7174 (N_7174,N_6618,N_6304);
nand U7175 (N_7175,N_6760,N_6841);
nand U7176 (N_7176,N_6472,N_6536);
nor U7177 (N_7177,N_6524,N_6850);
or U7178 (N_7178,N_6714,N_6698);
and U7179 (N_7179,N_6270,N_6609);
and U7180 (N_7180,N_6450,N_6808);
nand U7181 (N_7181,N_6449,N_6569);
nor U7182 (N_7182,N_6447,N_6679);
or U7183 (N_7183,N_6653,N_6382);
or U7184 (N_7184,N_6748,N_6419);
nor U7185 (N_7185,N_6871,N_6255);
nor U7186 (N_7186,N_6570,N_6622);
xor U7187 (N_7187,N_6366,N_6467);
nand U7188 (N_7188,N_6387,N_6493);
nand U7189 (N_7189,N_6823,N_6679);
and U7190 (N_7190,N_6419,N_6547);
and U7191 (N_7191,N_6411,N_6401);
nor U7192 (N_7192,N_6691,N_6779);
nor U7193 (N_7193,N_6576,N_6451);
nand U7194 (N_7194,N_6453,N_6591);
xnor U7195 (N_7195,N_6594,N_6325);
nor U7196 (N_7196,N_6732,N_6812);
xnor U7197 (N_7197,N_6413,N_6700);
nand U7198 (N_7198,N_6476,N_6354);
xor U7199 (N_7199,N_6547,N_6452);
xor U7200 (N_7200,N_6709,N_6638);
nand U7201 (N_7201,N_6856,N_6860);
nand U7202 (N_7202,N_6590,N_6485);
and U7203 (N_7203,N_6823,N_6660);
and U7204 (N_7204,N_6470,N_6665);
and U7205 (N_7205,N_6640,N_6754);
nand U7206 (N_7206,N_6701,N_6358);
or U7207 (N_7207,N_6669,N_6723);
or U7208 (N_7208,N_6684,N_6504);
or U7209 (N_7209,N_6253,N_6648);
xnor U7210 (N_7210,N_6560,N_6625);
nand U7211 (N_7211,N_6617,N_6458);
nor U7212 (N_7212,N_6666,N_6423);
or U7213 (N_7213,N_6714,N_6408);
and U7214 (N_7214,N_6695,N_6571);
or U7215 (N_7215,N_6691,N_6578);
xnor U7216 (N_7216,N_6760,N_6809);
or U7217 (N_7217,N_6554,N_6852);
and U7218 (N_7218,N_6445,N_6605);
nand U7219 (N_7219,N_6403,N_6691);
nor U7220 (N_7220,N_6393,N_6450);
nor U7221 (N_7221,N_6676,N_6689);
xor U7222 (N_7222,N_6582,N_6431);
or U7223 (N_7223,N_6627,N_6366);
or U7224 (N_7224,N_6644,N_6800);
xor U7225 (N_7225,N_6799,N_6292);
xnor U7226 (N_7226,N_6639,N_6680);
and U7227 (N_7227,N_6720,N_6595);
nand U7228 (N_7228,N_6253,N_6754);
and U7229 (N_7229,N_6855,N_6390);
nand U7230 (N_7230,N_6641,N_6379);
or U7231 (N_7231,N_6528,N_6725);
xnor U7232 (N_7232,N_6368,N_6579);
or U7233 (N_7233,N_6397,N_6420);
or U7234 (N_7234,N_6485,N_6384);
and U7235 (N_7235,N_6659,N_6820);
and U7236 (N_7236,N_6457,N_6837);
and U7237 (N_7237,N_6498,N_6627);
nor U7238 (N_7238,N_6319,N_6333);
nand U7239 (N_7239,N_6330,N_6325);
and U7240 (N_7240,N_6461,N_6663);
or U7241 (N_7241,N_6823,N_6257);
xor U7242 (N_7242,N_6282,N_6625);
and U7243 (N_7243,N_6599,N_6740);
nand U7244 (N_7244,N_6560,N_6558);
or U7245 (N_7245,N_6268,N_6528);
and U7246 (N_7246,N_6287,N_6597);
nor U7247 (N_7247,N_6431,N_6433);
and U7248 (N_7248,N_6253,N_6688);
xnor U7249 (N_7249,N_6300,N_6812);
or U7250 (N_7250,N_6661,N_6730);
nand U7251 (N_7251,N_6286,N_6764);
or U7252 (N_7252,N_6813,N_6685);
and U7253 (N_7253,N_6483,N_6848);
or U7254 (N_7254,N_6621,N_6442);
nor U7255 (N_7255,N_6819,N_6834);
or U7256 (N_7256,N_6527,N_6735);
nor U7257 (N_7257,N_6489,N_6545);
or U7258 (N_7258,N_6799,N_6735);
xor U7259 (N_7259,N_6874,N_6283);
nor U7260 (N_7260,N_6757,N_6480);
nor U7261 (N_7261,N_6379,N_6412);
nor U7262 (N_7262,N_6504,N_6591);
xor U7263 (N_7263,N_6534,N_6760);
xnor U7264 (N_7264,N_6382,N_6655);
and U7265 (N_7265,N_6693,N_6481);
and U7266 (N_7266,N_6300,N_6583);
or U7267 (N_7267,N_6740,N_6649);
nand U7268 (N_7268,N_6417,N_6656);
and U7269 (N_7269,N_6380,N_6669);
nand U7270 (N_7270,N_6406,N_6500);
nor U7271 (N_7271,N_6637,N_6374);
or U7272 (N_7272,N_6505,N_6517);
and U7273 (N_7273,N_6386,N_6309);
nand U7274 (N_7274,N_6677,N_6253);
nand U7275 (N_7275,N_6693,N_6568);
xor U7276 (N_7276,N_6311,N_6814);
nor U7277 (N_7277,N_6300,N_6630);
or U7278 (N_7278,N_6413,N_6691);
nand U7279 (N_7279,N_6793,N_6407);
nand U7280 (N_7280,N_6677,N_6784);
or U7281 (N_7281,N_6536,N_6763);
nand U7282 (N_7282,N_6345,N_6645);
nand U7283 (N_7283,N_6360,N_6481);
nand U7284 (N_7284,N_6762,N_6664);
and U7285 (N_7285,N_6694,N_6722);
nand U7286 (N_7286,N_6699,N_6370);
nand U7287 (N_7287,N_6704,N_6412);
nor U7288 (N_7288,N_6302,N_6351);
or U7289 (N_7289,N_6794,N_6582);
or U7290 (N_7290,N_6308,N_6403);
nand U7291 (N_7291,N_6422,N_6653);
nor U7292 (N_7292,N_6704,N_6330);
and U7293 (N_7293,N_6569,N_6555);
and U7294 (N_7294,N_6266,N_6271);
xor U7295 (N_7295,N_6562,N_6753);
nand U7296 (N_7296,N_6836,N_6277);
nand U7297 (N_7297,N_6310,N_6573);
nor U7298 (N_7298,N_6700,N_6409);
or U7299 (N_7299,N_6727,N_6634);
or U7300 (N_7300,N_6775,N_6403);
xor U7301 (N_7301,N_6704,N_6262);
nor U7302 (N_7302,N_6619,N_6486);
or U7303 (N_7303,N_6431,N_6435);
xor U7304 (N_7304,N_6464,N_6434);
and U7305 (N_7305,N_6285,N_6863);
or U7306 (N_7306,N_6393,N_6307);
and U7307 (N_7307,N_6646,N_6664);
nand U7308 (N_7308,N_6856,N_6339);
nor U7309 (N_7309,N_6594,N_6499);
nor U7310 (N_7310,N_6775,N_6479);
and U7311 (N_7311,N_6523,N_6520);
xnor U7312 (N_7312,N_6443,N_6510);
nand U7313 (N_7313,N_6313,N_6636);
nand U7314 (N_7314,N_6526,N_6466);
xnor U7315 (N_7315,N_6592,N_6391);
nor U7316 (N_7316,N_6856,N_6564);
or U7317 (N_7317,N_6759,N_6372);
or U7318 (N_7318,N_6728,N_6356);
xnor U7319 (N_7319,N_6737,N_6655);
nand U7320 (N_7320,N_6751,N_6774);
nand U7321 (N_7321,N_6850,N_6301);
or U7322 (N_7322,N_6287,N_6352);
nand U7323 (N_7323,N_6316,N_6731);
and U7324 (N_7324,N_6806,N_6622);
nor U7325 (N_7325,N_6412,N_6525);
or U7326 (N_7326,N_6828,N_6747);
or U7327 (N_7327,N_6343,N_6375);
nand U7328 (N_7328,N_6343,N_6622);
and U7329 (N_7329,N_6490,N_6777);
and U7330 (N_7330,N_6382,N_6567);
or U7331 (N_7331,N_6298,N_6275);
xnor U7332 (N_7332,N_6739,N_6746);
nand U7333 (N_7333,N_6280,N_6617);
nand U7334 (N_7334,N_6805,N_6327);
nor U7335 (N_7335,N_6667,N_6552);
xnor U7336 (N_7336,N_6755,N_6744);
nor U7337 (N_7337,N_6295,N_6673);
or U7338 (N_7338,N_6867,N_6810);
or U7339 (N_7339,N_6768,N_6467);
nor U7340 (N_7340,N_6664,N_6555);
nand U7341 (N_7341,N_6592,N_6564);
xnor U7342 (N_7342,N_6357,N_6577);
nand U7343 (N_7343,N_6713,N_6686);
nand U7344 (N_7344,N_6758,N_6447);
and U7345 (N_7345,N_6859,N_6266);
nor U7346 (N_7346,N_6552,N_6268);
or U7347 (N_7347,N_6647,N_6748);
xnor U7348 (N_7348,N_6826,N_6855);
xnor U7349 (N_7349,N_6566,N_6779);
xnor U7350 (N_7350,N_6696,N_6554);
nand U7351 (N_7351,N_6724,N_6794);
xnor U7352 (N_7352,N_6484,N_6786);
nand U7353 (N_7353,N_6727,N_6673);
and U7354 (N_7354,N_6486,N_6262);
nand U7355 (N_7355,N_6378,N_6319);
and U7356 (N_7356,N_6536,N_6816);
nor U7357 (N_7357,N_6270,N_6516);
nand U7358 (N_7358,N_6419,N_6388);
xor U7359 (N_7359,N_6470,N_6687);
nand U7360 (N_7360,N_6850,N_6868);
and U7361 (N_7361,N_6588,N_6780);
nand U7362 (N_7362,N_6803,N_6503);
xnor U7363 (N_7363,N_6764,N_6579);
nor U7364 (N_7364,N_6776,N_6483);
or U7365 (N_7365,N_6696,N_6309);
nor U7366 (N_7366,N_6334,N_6620);
or U7367 (N_7367,N_6267,N_6765);
nor U7368 (N_7368,N_6461,N_6662);
and U7369 (N_7369,N_6856,N_6850);
nor U7370 (N_7370,N_6274,N_6682);
nor U7371 (N_7371,N_6469,N_6298);
and U7372 (N_7372,N_6300,N_6304);
or U7373 (N_7373,N_6309,N_6800);
nor U7374 (N_7374,N_6573,N_6411);
and U7375 (N_7375,N_6556,N_6665);
or U7376 (N_7376,N_6417,N_6841);
and U7377 (N_7377,N_6326,N_6757);
and U7378 (N_7378,N_6657,N_6363);
nor U7379 (N_7379,N_6511,N_6325);
nand U7380 (N_7380,N_6430,N_6676);
and U7381 (N_7381,N_6679,N_6740);
nand U7382 (N_7382,N_6846,N_6719);
nand U7383 (N_7383,N_6320,N_6514);
and U7384 (N_7384,N_6749,N_6840);
nor U7385 (N_7385,N_6759,N_6501);
xnor U7386 (N_7386,N_6256,N_6508);
xor U7387 (N_7387,N_6856,N_6293);
xnor U7388 (N_7388,N_6294,N_6811);
xor U7389 (N_7389,N_6669,N_6405);
nor U7390 (N_7390,N_6495,N_6500);
and U7391 (N_7391,N_6568,N_6802);
and U7392 (N_7392,N_6560,N_6495);
nor U7393 (N_7393,N_6318,N_6420);
xor U7394 (N_7394,N_6644,N_6453);
and U7395 (N_7395,N_6851,N_6532);
nand U7396 (N_7396,N_6712,N_6766);
nor U7397 (N_7397,N_6271,N_6470);
nand U7398 (N_7398,N_6673,N_6761);
nor U7399 (N_7399,N_6392,N_6846);
and U7400 (N_7400,N_6836,N_6489);
nor U7401 (N_7401,N_6714,N_6862);
and U7402 (N_7402,N_6532,N_6817);
or U7403 (N_7403,N_6601,N_6820);
nor U7404 (N_7404,N_6839,N_6276);
xnor U7405 (N_7405,N_6757,N_6423);
or U7406 (N_7406,N_6536,N_6353);
and U7407 (N_7407,N_6808,N_6736);
nand U7408 (N_7408,N_6716,N_6327);
nand U7409 (N_7409,N_6779,N_6782);
xnor U7410 (N_7410,N_6596,N_6377);
nand U7411 (N_7411,N_6657,N_6277);
or U7412 (N_7412,N_6449,N_6405);
or U7413 (N_7413,N_6735,N_6339);
or U7414 (N_7414,N_6738,N_6611);
and U7415 (N_7415,N_6387,N_6765);
or U7416 (N_7416,N_6396,N_6385);
or U7417 (N_7417,N_6748,N_6271);
or U7418 (N_7418,N_6680,N_6527);
nand U7419 (N_7419,N_6810,N_6439);
xnor U7420 (N_7420,N_6703,N_6745);
nand U7421 (N_7421,N_6668,N_6505);
or U7422 (N_7422,N_6279,N_6512);
or U7423 (N_7423,N_6292,N_6387);
or U7424 (N_7424,N_6348,N_6308);
xor U7425 (N_7425,N_6569,N_6466);
or U7426 (N_7426,N_6299,N_6799);
nand U7427 (N_7427,N_6744,N_6331);
and U7428 (N_7428,N_6644,N_6404);
or U7429 (N_7429,N_6293,N_6542);
and U7430 (N_7430,N_6769,N_6411);
nand U7431 (N_7431,N_6529,N_6472);
and U7432 (N_7432,N_6436,N_6444);
or U7433 (N_7433,N_6522,N_6509);
nand U7434 (N_7434,N_6457,N_6800);
nand U7435 (N_7435,N_6559,N_6554);
or U7436 (N_7436,N_6650,N_6343);
nand U7437 (N_7437,N_6765,N_6263);
nor U7438 (N_7438,N_6733,N_6301);
nor U7439 (N_7439,N_6394,N_6270);
or U7440 (N_7440,N_6771,N_6564);
nor U7441 (N_7441,N_6417,N_6684);
nor U7442 (N_7442,N_6256,N_6433);
and U7443 (N_7443,N_6443,N_6873);
nor U7444 (N_7444,N_6505,N_6589);
or U7445 (N_7445,N_6683,N_6627);
nor U7446 (N_7446,N_6780,N_6260);
nand U7447 (N_7447,N_6396,N_6290);
nor U7448 (N_7448,N_6482,N_6494);
or U7449 (N_7449,N_6263,N_6557);
nand U7450 (N_7450,N_6521,N_6582);
nor U7451 (N_7451,N_6557,N_6693);
nor U7452 (N_7452,N_6439,N_6710);
nand U7453 (N_7453,N_6292,N_6832);
or U7454 (N_7454,N_6506,N_6825);
nand U7455 (N_7455,N_6763,N_6625);
nand U7456 (N_7456,N_6295,N_6437);
xnor U7457 (N_7457,N_6486,N_6572);
and U7458 (N_7458,N_6679,N_6627);
and U7459 (N_7459,N_6553,N_6512);
nor U7460 (N_7460,N_6359,N_6529);
nor U7461 (N_7461,N_6844,N_6284);
and U7462 (N_7462,N_6578,N_6435);
or U7463 (N_7463,N_6463,N_6666);
and U7464 (N_7464,N_6550,N_6845);
nor U7465 (N_7465,N_6331,N_6484);
or U7466 (N_7466,N_6526,N_6571);
and U7467 (N_7467,N_6874,N_6364);
and U7468 (N_7468,N_6715,N_6642);
nor U7469 (N_7469,N_6548,N_6801);
nand U7470 (N_7470,N_6480,N_6857);
or U7471 (N_7471,N_6378,N_6329);
and U7472 (N_7472,N_6531,N_6656);
xnor U7473 (N_7473,N_6754,N_6730);
nor U7474 (N_7474,N_6780,N_6269);
and U7475 (N_7475,N_6536,N_6874);
nand U7476 (N_7476,N_6730,N_6329);
or U7477 (N_7477,N_6495,N_6328);
nand U7478 (N_7478,N_6431,N_6432);
xor U7479 (N_7479,N_6667,N_6573);
or U7480 (N_7480,N_6811,N_6788);
or U7481 (N_7481,N_6632,N_6785);
nor U7482 (N_7482,N_6488,N_6834);
xnor U7483 (N_7483,N_6376,N_6342);
and U7484 (N_7484,N_6538,N_6560);
or U7485 (N_7485,N_6780,N_6528);
nor U7486 (N_7486,N_6643,N_6268);
nand U7487 (N_7487,N_6409,N_6278);
and U7488 (N_7488,N_6720,N_6514);
or U7489 (N_7489,N_6793,N_6682);
xor U7490 (N_7490,N_6251,N_6319);
nand U7491 (N_7491,N_6415,N_6373);
or U7492 (N_7492,N_6261,N_6646);
xor U7493 (N_7493,N_6710,N_6674);
xor U7494 (N_7494,N_6358,N_6373);
xnor U7495 (N_7495,N_6304,N_6330);
or U7496 (N_7496,N_6266,N_6453);
nand U7497 (N_7497,N_6480,N_6407);
and U7498 (N_7498,N_6445,N_6622);
xnor U7499 (N_7499,N_6281,N_6485);
xor U7500 (N_7500,N_7326,N_6931);
nor U7501 (N_7501,N_6896,N_7417);
nor U7502 (N_7502,N_6945,N_7004);
nand U7503 (N_7503,N_6973,N_6907);
nand U7504 (N_7504,N_7309,N_6943);
or U7505 (N_7505,N_7399,N_7232);
xnor U7506 (N_7506,N_7266,N_7356);
nand U7507 (N_7507,N_7174,N_7291);
nor U7508 (N_7508,N_7261,N_7325);
nand U7509 (N_7509,N_7071,N_6947);
nor U7510 (N_7510,N_7236,N_7223);
nand U7511 (N_7511,N_6909,N_6913);
or U7512 (N_7512,N_7431,N_7407);
xor U7513 (N_7513,N_7051,N_7328);
nand U7514 (N_7514,N_7163,N_7464);
nand U7515 (N_7515,N_7015,N_7436);
nor U7516 (N_7516,N_7005,N_7211);
and U7517 (N_7517,N_7199,N_7140);
nand U7518 (N_7518,N_7082,N_7184);
xnor U7519 (N_7519,N_7432,N_7280);
nor U7520 (N_7520,N_7455,N_7052);
xor U7521 (N_7521,N_7127,N_7076);
xor U7522 (N_7522,N_7305,N_7377);
and U7523 (N_7523,N_7389,N_7249);
or U7524 (N_7524,N_7268,N_7300);
nor U7525 (N_7525,N_7320,N_7347);
nor U7526 (N_7526,N_7074,N_7085);
or U7527 (N_7527,N_7383,N_6929);
and U7528 (N_7528,N_7073,N_7042);
and U7529 (N_7529,N_7272,N_7070);
nand U7530 (N_7530,N_7350,N_7391);
xor U7531 (N_7531,N_7386,N_7486);
nand U7532 (N_7532,N_7296,N_7090);
nor U7533 (N_7533,N_7016,N_7259);
xnor U7534 (N_7534,N_7158,N_7092);
or U7535 (N_7535,N_7164,N_7485);
xnor U7536 (N_7536,N_7478,N_6980);
and U7537 (N_7537,N_7021,N_7243);
or U7538 (N_7538,N_7210,N_7028);
nand U7539 (N_7539,N_7306,N_7061);
or U7540 (N_7540,N_6894,N_6975);
nor U7541 (N_7541,N_6920,N_7418);
xor U7542 (N_7542,N_7014,N_7382);
xor U7543 (N_7543,N_7474,N_7302);
nand U7544 (N_7544,N_7000,N_7240);
xor U7545 (N_7545,N_7394,N_7027);
nor U7546 (N_7546,N_7038,N_7170);
nor U7547 (N_7547,N_7427,N_7238);
or U7548 (N_7548,N_7494,N_7112);
and U7549 (N_7549,N_7186,N_6940);
or U7550 (N_7550,N_7050,N_7117);
nand U7551 (N_7551,N_7343,N_7047);
xnor U7552 (N_7552,N_7145,N_6904);
and U7553 (N_7553,N_7314,N_7321);
xor U7554 (N_7554,N_6983,N_7020);
nor U7555 (N_7555,N_6902,N_7469);
xnor U7556 (N_7556,N_6892,N_7322);
or U7557 (N_7557,N_7088,N_6933);
nand U7558 (N_7558,N_7152,N_7313);
nor U7559 (N_7559,N_6995,N_7330);
nor U7560 (N_7560,N_6887,N_7096);
or U7561 (N_7561,N_7337,N_6890);
nand U7562 (N_7562,N_7196,N_7242);
xnor U7563 (N_7563,N_7404,N_7362);
nor U7564 (N_7564,N_7087,N_7408);
or U7565 (N_7565,N_7026,N_7487);
nor U7566 (N_7566,N_7398,N_7103);
and U7567 (N_7567,N_7176,N_7098);
or U7568 (N_7568,N_7282,N_7034);
and U7569 (N_7569,N_7017,N_7339);
xor U7570 (N_7570,N_7045,N_7284);
nor U7571 (N_7571,N_7361,N_6934);
nand U7572 (N_7572,N_7003,N_6958);
xnor U7573 (N_7573,N_7388,N_7270);
and U7574 (N_7574,N_7493,N_7244);
and U7575 (N_7575,N_7159,N_7497);
and U7576 (N_7576,N_7413,N_7479);
xnor U7577 (N_7577,N_7315,N_7369);
and U7578 (N_7578,N_7414,N_7183);
nand U7579 (N_7579,N_7416,N_7318);
nor U7580 (N_7580,N_7208,N_7205);
nor U7581 (N_7581,N_7009,N_7430);
xor U7582 (N_7582,N_6905,N_6988);
nor U7583 (N_7583,N_7260,N_7068);
nand U7584 (N_7584,N_7466,N_7058);
or U7585 (N_7585,N_7462,N_7125);
or U7586 (N_7586,N_7108,N_7079);
nor U7587 (N_7587,N_6974,N_7379);
xor U7588 (N_7588,N_7372,N_7273);
nor U7589 (N_7589,N_7460,N_7447);
nor U7590 (N_7590,N_6936,N_7024);
nand U7591 (N_7591,N_7498,N_7335);
and U7592 (N_7592,N_7138,N_7143);
and U7593 (N_7593,N_6951,N_7165);
nand U7594 (N_7594,N_7214,N_7317);
xnor U7595 (N_7595,N_7212,N_7064);
xor U7596 (N_7596,N_7329,N_7048);
and U7597 (N_7597,N_7422,N_7075);
or U7598 (N_7598,N_7457,N_7477);
xor U7599 (N_7599,N_6918,N_7336);
or U7600 (N_7600,N_7118,N_7093);
nor U7601 (N_7601,N_7171,N_7482);
xor U7602 (N_7602,N_7195,N_7181);
or U7603 (N_7603,N_7292,N_6901);
nor U7604 (N_7604,N_7278,N_7451);
nor U7605 (N_7605,N_7332,N_7324);
nand U7606 (N_7606,N_7450,N_6898);
nor U7607 (N_7607,N_7147,N_7166);
or U7608 (N_7608,N_7371,N_7080);
nor U7609 (N_7609,N_7380,N_7275);
or U7610 (N_7610,N_7222,N_7049);
nand U7611 (N_7611,N_6993,N_6927);
nor U7612 (N_7612,N_7334,N_7011);
and U7613 (N_7613,N_7409,N_7412);
nor U7614 (N_7614,N_7323,N_7220);
and U7615 (N_7615,N_7423,N_7230);
nand U7616 (N_7616,N_7445,N_7297);
nand U7617 (N_7617,N_6967,N_7002);
nor U7618 (N_7618,N_7354,N_6893);
nor U7619 (N_7619,N_7495,N_7089);
nand U7620 (N_7620,N_6969,N_7472);
xor U7621 (N_7621,N_7031,N_6932);
nand U7622 (N_7622,N_7151,N_7022);
nand U7623 (N_7623,N_7209,N_7131);
nand U7624 (N_7624,N_7149,N_6908);
and U7625 (N_7625,N_7344,N_6957);
xnor U7626 (N_7626,N_7206,N_7218);
or U7627 (N_7627,N_7060,N_7032);
nor U7628 (N_7628,N_7458,N_7374);
or U7629 (N_7629,N_6981,N_7126);
and U7630 (N_7630,N_6895,N_6986);
nor U7631 (N_7631,N_7378,N_7342);
nor U7632 (N_7632,N_7421,N_7191);
or U7633 (N_7633,N_7490,N_7215);
or U7634 (N_7634,N_7440,N_7241);
and U7635 (N_7635,N_7393,N_7100);
and U7636 (N_7636,N_7392,N_7453);
nand U7637 (N_7637,N_6998,N_7109);
nor U7638 (N_7638,N_7056,N_7267);
and U7639 (N_7639,N_6915,N_6930);
xor U7640 (N_7640,N_6991,N_7304);
xnor U7641 (N_7641,N_7426,N_7405);
nand U7642 (N_7642,N_7102,N_6878);
xor U7643 (N_7643,N_7084,N_7247);
or U7644 (N_7644,N_7299,N_7496);
and U7645 (N_7645,N_7072,N_7415);
nand U7646 (N_7646,N_7338,N_7246);
and U7647 (N_7647,N_7256,N_7122);
and U7648 (N_7648,N_6875,N_7144);
xor U7649 (N_7649,N_6886,N_6877);
nor U7650 (N_7650,N_6944,N_7269);
nand U7651 (N_7651,N_7133,N_7274);
and U7652 (N_7652,N_7029,N_7281);
nand U7653 (N_7653,N_7475,N_7465);
nand U7654 (N_7654,N_7177,N_7197);
nor U7655 (N_7655,N_7040,N_6885);
xnor U7656 (N_7656,N_7425,N_7262);
and U7657 (N_7657,N_7258,N_7167);
nand U7658 (N_7658,N_6903,N_7444);
xnor U7659 (N_7659,N_7201,N_7333);
nand U7660 (N_7660,N_7007,N_7289);
or U7661 (N_7661,N_7190,N_7055);
or U7662 (N_7662,N_7437,N_7248);
or U7663 (N_7663,N_6990,N_6964);
and U7664 (N_7664,N_7033,N_6984);
xnor U7665 (N_7665,N_7194,N_7169);
nand U7666 (N_7666,N_7428,N_7341);
xnor U7667 (N_7667,N_7119,N_7067);
xnor U7668 (N_7668,N_7193,N_7271);
xnor U7669 (N_7669,N_7406,N_7010);
and U7670 (N_7670,N_6917,N_7419);
nand U7671 (N_7671,N_6942,N_6914);
nand U7672 (N_7672,N_7233,N_7142);
or U7673 (N_7673,N_7095,N_7429);
xnor U7674 (N_7674,N_7053,N_7018);
and U7675 (N_7675,N_6950,N_6924);
xnor U7676 (N_7676,N_7225,N_6994);
nor U7677 (N_7677,N_6992,N_6926);
nor U7678 (N_7678,N_7039,N_7204);
or U7679 (N_7679,N_6949,N_7463);
and U7680 (N_7680,N_7366,N_7301);
nor U7681 (N_7681,N_6968,N_7285);
and U7682 (N_7682,N_7139,N_7359);
nand U7683 (N_7683,N_6963,N_6966);
and U7684 (N_7684,N_7396,N_7360);
or U7685 (N_7685,N_7065,N_7221);
xor U7686 (N_7686,N_6999,N_7358);
nor U7687 (N_7687,N_7449,N_7006);
nor U7688 (N_7688,N_7349,N_7134);
nor U7689 (N_7689,N_7227,N_7168);
xor U7690 (N_7690,N_7111,N_7254);
or U7691 (N_7691,N_6948,N_7390);
nand U7692 (N_7692,N_7294,N_6977);
xnor U7693 (N_7693,N_7293,N_7381);
xnor U7694 (N_7694,N_7403,N_7251);
xnor U7695 (N_7695,N_7252,N_7121);
nand U7696 (N_7696,N_7120,N_7245);
or U7697 (N_7697,N_7077,N_7387);
nor U7698 (N_7698,N_7008,N_7130);
nand U7699 (N_7699,N_7491,N_7019);
or U7700 (N_7700,N_7373,N_7327);
xor U7701 (N_7701,N_7202,N_7346);
and U7702 (N_7702,N_7172,N_7137);
nand U7703 (N_7703,N_6900,N_7484);
nor U7704 (N_7704,N_7062,N_7146);
and U7705 (N_7705,N_6979,N_7424);
or U7706 (N_7706,N_6939,N_7448);
nor U7707 (N_7707,N_7250,N_6880);
nand U7708 (N_7708,N_7253,N_7030);
xnor U7709 (N_7709,N_7213,N_7298);
or U7710 (N_7710,N_7279,N_7368);
nand U7711 (N_7711,N_7036,N_7277);
or U7712 (N_7712,N_6970,N_7470);
nand U7713 (N_7713,N_6883,N_7043);
or U7714 (N_7714,N_6961,N_7124);
or U7715 (N_7715,N_7364,N_7156);
xor U7716 (N_7716,N_7499,N_6978);
or U7717 (N_7717,N_7441,N_7385);
xor U7718 (N_7718,N_7255,N_7363);
nand U7719 (N_7719,N_7216,N_7400);
xor U7720 (N_7720,N_7001,N_7395);
xor U7721 (N_7721,N_7310,N_7150);
nand U7722 (N_7722,N_7200,N_7483);
nand U7723 (N_7723,N_6911,N_6937);
and U7724 (N_7724,N_7239,N_6925);
and U7725 (N_7725,N_7160,N_7287);
or U7726 (N_7726,N_7207,N_6912);
and U7727 (N_7727,N_7229,N_6960);
and U7728 (N_7728,N_6881,N_7286);
nor U7729 (N_7729,N_7257,N_7037);
or U7730 (N_7730,N_7434,N_6965);
or U7731 (N_7731,N_7288,N_7110);
and U7732 (N_7732,N_7179,N_7459);
nor U7733 (N_7733,N_7066,N_7198);
nor U7734 (N_7734,N_6971,N_7107);
nand U7735 (N_7735,N_7316,N_7471);
or U7736 (N_7736,N_7442,N_7044);
and U7737 (N_7737,N_7263,N_7078);
nor U7738 (N_7738,N_7370,N_7081);
or U7739 (N_7739,N_7148,N_7443);
xor U7740 (N_7740,N_6891,N_7123);
and U7741 (N_7741,N_7135,N_7188);
nand U7742 (N_7742,N_7094,N_7097);
and U7743 (N_7743,N_7203,N_7411);
xor U7744 (N_7744,N_7116,N_7155);
nor U7745 (N_7745,N_7231,N_6935);
xor U7746 (N_7746,N_7153,N_7025);
xnor U7747 (N_7747,N_7136,N_7059);
or U7748 (N_7748,N_7452,N_6959);
or U7749 (N_7749,N_7456,N_7128);
or U7750 (N_7750,N_6952,N_6921);
or U7751 (N_7751,N_6884,N_7086);
xnor U7752 (N_7752,N_6962,N_6996);
and U7753 (N_7753,N_6997,N_7173);
or U7754 (N_7754,N_7105,N_6954);
or U7755 (N_7755,N_7083,N_7224);
or U7756 (N_7756,N_7489,N_7397);
and U7757 (N_7757,N_7446,N_7023);
nor U7758 (N_7758,N_7355,N_7161);
or U7759 (N_7759,N_7467,N_6946);
and U7760 (N_7760,N_7488,N_7132);
or U7761 (N_7761,N_6987,N_6989);
and U7762 (N_7762,N_7013,N_7180);
xnor U7763 (N_7763,N_7384,N_7290);
nor U7764 (N_7764,N_6910,N_7192);
or U7765 (N_7765,N_7219,N_6897);
nor U7766 (N_7766,N_7376,N_6985);
and U7767 (N_7767,N_6879,N_7438);
xor U7768 (N_7768,N_6953,N_7226);
and U7769 (N_7769,N_7115,N_7114);
or U7770 (N_7770,N_6888,N_7420);
xor U7771 (N_7771,N_7473,N_6938);
or U7772 (N_7772,N_7228,N_7357);
or U7773 (N_7773,N_7012,N_7307);
xor U7774 (N_7774,N_7367,N_7154);
nor U7775 (N_7775,N_7454,N_7311);
nor U7776 (N_7776,N_6882,N_7063);
nor U7777 (N_7777,N_7046,N_7480);
nor U7778 (N_7778,N_6922,N_7435);
nor U7779 (N_7779,N_7185,N_7352);
xor U7780 (N_7780,N_7476,N_6955);
nand U7781 (N_7781,N_7433,N_7264);
nand U7782 (N_7782,N_6976,N_7178);
nand U7783 (N_7783,N_6906,N_7401);
and U7784 (N_7784,N_7265,N_7234);
nand U7785 (N_7785,N_7217,N_7351);
and U7786 (N_7786,N_7162,N_7461);
or U7787 (N_7787,N_7402,N_7348);
nor U7788 (N_7788,N_7295,N_6876);
nand U7789 (N_7789,N_6899,N_6916);
nand U7790 (N_7790,N_7091,N_7353);
or U7791 (N_7791,N_7365,N_7069);
xor U7792 (N_7792,N_7340,N_7035);
and U7793 (N_7793,N_6919,N_7175);
xor U7794 (N_7794,N_7345,N_6923);
nor U7795 (N_7795,N_7101,N_7187);
nor U7796 (N_7796,N_7106,N_7057);
and U7797 (N_7797,N_7319,N_7104);
and U7798 (N_7798,N_7235,N_7283);
nor U7799 (N_7799,N_7410,N_6889);
and U7800 (N_7800,N_7331,N_7054);
xnor U7801 (N_7801,N_6982,N_7182);
and U7802 (N_7802,N_7041,N_6972);
nand U7803 (N_7803,N_7312,N_6941);
nor U7804 (N_7804,N_7099,N_7157);
or U7805 (N_7805,N_7113,N_7468);
or U7806 (N_7806,N_7439,N_6928);
xor U7807 (N_7807,N_7189,N_7129);
nor U7808 (N_7808,N_7481,N_7375);
or U7809 (N_7809,N_7303,N_7276);
nand U7810 (N_7810,N_7141,N_7308);
nor U7811 (N_7811,N_6956,N_7237);
and U7812 (N_7812,N_7492,N_7240);
nor U7813 (N_7813,N_7142,N_7014);
nand U7814 (N_7814,N_7177,N_7148);
and U7815 (N_7815,N_7379,N_7131);
nor U7816 (N_7816,N_7204,N_7145);
or U7817 (N_7817,N_6933,N_6907);
and U7818 (N_7818,N_7021,N_7092);
and U7819 (N_7819,N_7425,N_7401);
nor U7820 (N_7820,N_7196,N_7327);
and U7821 (N_7821,N_7069,N_7433);
and U7822 (N_7822,N_7452,N_7141);
nor U7823 (N_7823,N_7103,N_6915);
and U7824 (N_7824,N_7169,N_6916);
nor U7825 (N_7825,N_7210,N_6909);
and U7826 (N_7826,N_7188,N_7086);
nor U7827 (N_7827,N_6945,N_7283);
and U7828 (N_7828,N_7478,N_7411);
nor U7829 (N_7829,N_7239,N_7038);
or U7830 (N_7830,N_7353,N_7060);
nand U7831 (N_7831,N_7307,N_6961);
nor U7832 (N_7832,N_7230,N_7443);
nor U7833 (N_7833,N_7071,N_7385);
nor U7834 (N_7834,N_7251,N_7098);
or U7835 (N_7835,N_7306,N_7262);
or U7836 (N_7836,N_7002,N_7238);
and U7837 (N_7837,N_7101,N_7233);
and U7838 (N_7838,N_7486,N_6942);
nor U7839 (N_7839,N_7018,N_7493);
nor U7840 (N_7840,N_7161,N_6911);
xnor U7841 (N_7841,N_7073,N_7457);
nor U7842 (N_7842,N_7272,N_7047);
and U7843 (N_7843,N_7030,N_7235);
nor U7844 (N_7844,N_7352,N_7411);
and U7845 (N_7845,N_7322,N_7043);
nor U7846 (N_7846,N_7308,N_7422);
nand U7847 (N_7847,N_7342,N_7118);
xnor U7848 (N_7848,N_7367,N_7239);
or U7849 (N_7849,N_6995,N_7301);
nand U7850 (N_7850,N_7406,N_6913);
nand U7851 (N_7851,N_7412,N_7478);
xnor U7852 (N_7852,N_7103,N_7166);
nand U7853 (N_7853,N_7394,N_7024);
or U7854 (N_7854,N_7034,N_7324);
nor U7855 (N_7855,N_7462,N_6883);
or U7856 (N_7856,N_6968,N_7420);
nand U7857 (N_7857,N_7281,N_7363);
or U7858 (N_7858,N_7118,N_7365);
nor U7859 (N_7859,N_7322,N_6907);
and U7860 (N_7860,N_6952,N_7366);
xnor U7861 (N_7861,N_7278,N_6979);
nand U7862 (N_7862,N_6998,N_7298);
or U7863 (N_7863,N_7338,N_7425);
or U7864 (N_7864,N_7279,N_7217);
nor U7865 (N_7865,N_6933,N_6962);
and U7866 (N_7866,N_7375,N_7074);
xnor U7867 (N_7867,N_7018,N_6920);
and U7868 (N_7868,N_7290,N_6887);
and U7869 (N_7869,N_7408,N_7372);
nand U7870 (N_7870,N_6929,N_6908);
or U7871 (N_7871,N_7134,N_7398);
or U7872 (N_7872,N_7082,N_7080);
nand U7873 (N_7873,N_7292,N_6914);
nor U7874 (N_7874,N_7084,N_7471);
nand U7875 (N_7875,N_7360,N_6969);
nand U7876 (N_7876,N_6879,N_7101);
nor U7877 (N_7877,N_7121,N_7135);
nor U7878 (N_7878,N_7194,N_7329);
or U7879 (N_7879,N_7330,N_7486);
nor U7880 (N_7880,N_7490,N_7280);
and U7881 (N_7881,N_7021,N_7489);
and U7882 (N_7882,N_7408,N_7392);
xnor U7883 (N_7883,N_7075,N_7334);
nor U7884 (N_7884,N_7233,N_7126);
nand U7885 (N_7885,N_7128,N_7112);
nor U7886 (N_7886,N_7204,N_7038);
nand U7887 (N_7887,N_7228,N_7389);
and U7888 (N_7888,N_7170,N_7220);
and U7889 (N_7889,N_7365,N_7444);
or U7890 (N_7890,N_6962,N_6886);
xnor U7891 (N_7891,N_7160,N_7064);
nand U7892 (N_7892,N_6968,N_7086);
nor U7893 (N_7893,N_7367,N_7256);
xnor U7894 (N_7894,N_7110,N_7172);
nor U7895 (N_7895,N_7239,N_7121);
nor U7896 (N_7896,N_7380,N_7061);
and U7897 (N_7897,N_7065,N_7495);
or U7898 (N_7898,N_7439,N_7373);
or U7899 (N_7899,N_7350,N_7465);
and U7900 (N_7900,N_7369,N_6939);
and U7901 (N_7901,N_7404,N_7261);
xor U7902 (N_7902,N_6953,N_7295);
nor U7903 (N_7903,N_7395,N_7499);
xor U7904 (N_7904,N_7291,N_7499);
nand U7905 (N_7905,N_7322,N_7011);
xnor U7906 (N_7906,N_7496,N_7141);
nand U7907 (N_7907,N_6915,N_6971);
nor U7908 (N_7908,N_7109,N_6961);
nor U7909 (N_7909,N_7266,N_7454);
nor U7910 (N_7910,N_7460,N_7405);
or U7911 (N_7911,N_7107,N_7159);
nor U7912 (N_7912,N_7360,N_7353);
and U7913 (N_7913,N_7038,N_7485);
and U7914 (N_7914,N_7406,N_6948);
xnor U7915 (N_7915,N_7492,N_7029);
xor U7916 (N_7916,N_7225,N_7172);
nand U7917 (N_7917,N_7436,N_7437);
xor U7918 (N_7918,N_7152,N_7086);
nor U7919 (N_7919,N_6942,N_6947);
xnor U7920 (N_7920,N_7171,N_7299);
or U7921 (N_7921,N_7003,N_6883);
nor U7922 (N_7922,N_7241,N_7234);
and U7923 (N_7923,N_7408,N_7077);
nand U7924 (N_7924,N_7413,N_7045);
xnor U7925 (N_7925,N_7293,N_7023);
nand U7926 (N_7926,N_7444,N_6926);
or U7927 (N_7927,N_6933,N_7373);
nand U7928 (N_7928,N_7149,N_6934);
nor U7929 (N_7929,N_7155,N_7247);
nor U7930 (N_7930,N_6957,N_7051);
or U7931 (N_7931,N_6967,N_7085);
or U7932 (N_7932,N_7141,N_7179);
nand U7933 (N_7933,N_7405,N_7106);
xnor U7934 (N_7934,N_7030,N_7184);
and U7935 (N_7935,N_6927,N_6885);
and U7936 (N_7936,N_6933,N_6884);
nor U7937 (N_7937,N_7392,N_7179);
or U7938 (N_7938,N_7204,N_7205);
or U7939 (N_7939,N_7272,N_7352);
or U7940 (N_7940,N_7147,N_7110);
nand U7941 (N_7941,N_7437,N_7241);
nand U7942 (N_7942,N_7369,N_7389);
xor U7943 (N_7943,N_6990,N_7106);
xnor U7944 (N_7944,N_7089,N_7193);
or U7945 (N_7945,N_7439,N_7428);
nand U7946 (N_7946,N_7439,N_7020);
nand U7947 (N_7947,N_7127,N_7295);
nor U7948 (N_7948,N_7185,N_7378);
nand U7949 (N_7949,N_6937,N_6947);
and U7950 (N_7950,N_7224,N_6878);
or U7951 (N_7951,N_6917,N_7452);
and U7952 (N_7952,N_7475,N_7290);
or U7953 (N_7953,N_7424,N_7128);
and U7954 (N_7954,N_7102,N_7437);
and U7955 (N_7955,N_7312,N_6965);
nor U7956 (N_7956,N_6878,N_7137);
nor U7957 (N_7957,N_7442,N_7226);
or U7958 (N_7958,N_7387,N_7222);
nor U7959 (N_7959,N_6943,N_7148);
nor U7960 (N_7960,N_7117,N_7239);
and U7961 (N_7961,N_6882,N_7104);
xnor U7962 (N_7962,N_7335,N_7198);
xor U7963 (N_7963,N_7223,N_7492);
nor U7964 (N_7964,N_7082,N_7358);
xor U7965 (N_7965,N_7287,N_7490);
nor U7966 (N_7966,N_7134,N_7182);
nor U7967 (N_7967,N_7238,N_7176);
and U7968 (N_7968,N_7150,N_7329);
or U7969 (N_7969,N_7444,N_7069);
nor U7970 (N_7970,N_6960,N_7421);
nor U7971 (N_7971,N_7393,N_7211);
or U7972 (N_7972,N_7444,N_7279);
xor U7973 (N_7973,N_7453,N_7047);
nor U7974 (N_7974,N_7156,N_7193);
or U7975 (N_7975,N_7474,N_7146);
xnor U7976 (N_7976,N_7114,N_7322);
nor U7977 (N_7977,N_7073,N_7425);
or U7978 (N_7978,N_7033,N_7412);
xnor U7979 (N_7979,N_7394,N_7450);
xor U7980 (N_7980,N_7088,N_7230);
nor U7981 (N_7981,N_7348,N_7084);
nor U7982 (N_7982,N_6943,N_6935);
xnor U7983 (N_7983,N_6955,N_7096);
and U7984 (N_7984,N_7285,N_7014);
nor U7985 (N_7985,N_7262,N_7310);
and U7986 (N_7986,N_7431,N_7357);
or U7987 (N_7987,N_7366,N_7201);
nor U7988 (N_7988,N_7317,N_7245);
or U7989 (N_7989,N_7353,N_7026);
xor U7990 (N_7990,N_7473,N_7421);
xnor U7991 (N_7991,N_6899,N_7496);
nor U7992 (N_7992,N_7388,N_7246);
or U7993 (N_7993,N_7104,N_7192);
nor U7994 (N_7994,N_6962,N_7176);
or U7995 (N_7995,N_7204,N_7301);
xor U7996 (N_7996,N_7075,N_7357);
and U7997 (N_7997,N_7114,N_6884);
or U7998 (N_7998,N_7158,N_7265);
nor U7999 (N_7999,N_7062,N_6958);
or U8000 (N_8000,N_7410,N_7477);
and U8001 (N_8001,N_6913,N_7492);
nand U8002 (N_8002,N_7159,N_7327);
nor U8003 (N_8003,N_7322,N_6940);
nor U8004 (N_8004,N_7049,N_7458);
xnor U8005 (N_8005,N_6923,N_7400);
nor U8006 (N_8006,N_7360,N_7085);
xor U8007 (N_8007,N_7288,N_7318);
and U8008 (N_8008,N_6974,N_7133);
nand U8009 (N_8009,N_7318,N_7296);
nand U8010 (N_8010,N_7199,N_7466);
and U8011 (N_8011,N_7069,N_7041);
or U8012 (N_8012,N_6954,N_7211);
nand U8013 (N_8013,N_7439,N_6889);
nor U8014 (N_8014,N_6991,N_7272);
nor U8015 (N_8015,N_7036,N_6998);
nand U8016 (N_8016,N_7394,N_7050);
and U8017 (N_8017,N_7157,N_7431);
nand U8018 (N_8018,N_7368,N_7481);
and U8019 (N_8019,N_7418,N_7267);
and U8020 (N_8020,N_7235,N_6914);
and U8021 (N_8021,N_7061,N_7430);
or U8022 (N_8022,N_7093,N_7270);
xor U8023 (N_8023,N_7157,N_7266);
nand U8024 (N_8024,N_7283,N_7418);
nand U8025 (N_8025,N_7417,N_7225);
nor U8026 (N_8026,N_7478,N_7402);
and U8027 (N_8027,N_7489,N_7061);
nand U8028 (N_8028,N_7056,N_7035);
and U8029 (N_8029,N_6989,N_7093);
and U8030 (N_8030,N_7155,N_7443);
and U8031 (N_8031,N_7385,N_7329);
xnor U8032 (N_8032,N_6978,N_6969);
nor U8033 (N_8033,N_7078,N_7444);
nor U8034 (N_8034,N_7323,N_7151);
nor U8035 (N_8035,N_7400,N_7329);
nor U8036 (N_8036,N_7483,N_7268);
nand U8037 (N_8037,N_7440,N_7286);
xor U8038 (N_8038,N_7024,N_7045);
or U8039 (N_8039,N_7234,N_7133);
nand U8040 (N_8040,N_7431,N_6992);
nand U8041 (N_8041,N_7241,N_7154);
nor U8042 (N_8042,N_7026,N_6994);
xnor U8043 (N_8043,N_7247,N_7442);
nor U8044 (N_8044,N_7174,N_7439);
and U8045 (N_8045,N_6970,N_7338);
and U8046 (N_8046,N_7499,N_7366);
or U8047 (N_8047,N_7200,N_7017);
xor U8048 (N_8048,N_7048,N_7119);
or U8049 (N_8049,N_6934,N_7131);
and U8050 (N_8050,N_7160,N_7241);
xor U8051 (N_8051,N_7303,N_6993);
and U8052 (N_8052,N_7185,N_7196);
nand U8053 (N_8053,N_7267,N_7283);
and U8054 (N_8054,N_7058,N_7103);
or U8055 (N_8055,N_6905,N_7329);
nor U8056 (N_8056,N_7496,N_7125);
nor U8057 (N_8057,N_7373,N_7064);
and U8058 (N_8058,N_6896,N_7208);
xnor U8059 (N_8059,N_7321,N_7179);
and U8060 (N_8060,N_7479,N_7296);
and U8061 (N_8061,N_7443,N_6881);
or U8062 (N_8062,N_7348,N_6945);
nor U8063 (N_8063,N_7027,N_6999);
and U8064 (N_8064,N_7408,N_7044);
nand U8065 (N_8065,N_6914,N_7349);
nand U8066 (N_8066,N_7013,N_7302);
nand U8067 (N_8067,N_7035,N_7176);
or U8068 (N_8068,N_7242,N_7324);
nor U8069 (N_8069,N_7138,N_7027);
nor U8070 (N_8070,N_7425,N_6877);
nand U8071 (N_8071,N_7042,N_7248);
nor U8072 (N_8072,N_7312,N_6931);
or U8073 (N_8073,N_7198,N_7011);
or U8074 (N_8074,N_7122,N_7251);
or U8075 (N_8075,N_7368,N_7157);
and U8076 (N_8076,N_7268,N_6960);
and U8077 (N_8077,N_7369,N_7186);
or U8078 (N_8078,N_7445,N_7417);
nand U8079 (N_8079,N_7417,N_7034);
or U8080 (N_8080,N_7482,N_7256);
nand U8081 (N_8081,N_6962,N_7439);
xnor U8082 (N_8082,N_7425,N_7491);
xnor U8083 (N_8083,N_7471,N_6953);
nand U8084 (N_8084,N_7493,N_7479);
nor U8085 (N_8085,N_7308,N_7441);
nor U8086 (N_8086,N_7051,N_6995);
xor U8087 (N_8087,N_7409,N_7281);
xor U8088 (N_8088,N_7061,N_6992);
nand U8089 (N_8089,N_6956,N_6974);
xor U8090 (N_8090,N_7359,N_7173);
nor U8091 (N_8091,N_7074,N_7202);
xor U8092 (N_8092,N_6981,N_7111);
and U8093 (N_8093,N_7095,N_7200);
and U8094 (N_8094,N_7430,N_7341);
and U8095 (N_8095,N_7422,N_7167);
nand U8096 (N_8096,N_7098,N_7220);
and U8097 (N_8097,N_6960,N_7013);
and U8098 (N_8098,N_7321,N_7436);
nand U8099 (N_8099,N_7479,N_7285);
nor U8100 (N_8100,N_6958,N_6909);
or U8101 (N_8101,N_7484,N_7380);
or U8102 (N_8102,N_7245,N_7248);
xnor U8103 (N_8103,N_7172,N_7469);
and U8104 (N_8104,N_7110,N_7186);
and U8105 (N_8105,N_7311,N_7446);
xnor U8106 (N_8106,N_6963,N_7110);
xor U8107 (N_8107,N_7340,N_7162);
nand U8108 (N_8108,N_7144,N_7127);
xnor U8109 (N_8109,N_6944,N_7396);
and U8110 (N_8110,N_7134,N_7095);
xor U8111 (N_8111,N_7043,N_7027);
or U8112 (N_8112,N_6953,N_7029);
nand U8113 (N_8113,N_6972,N_6947);
nor U8114 (N_8114,N_7025,N_7126);
xnor U8115 (N_8115,N_6949,N_6976);
or U8116 (N_8116,N_7001,N_7414);
or U8117 (N_8117,N_6936,N_7239);
nor U8118 (N_8118,N_7181,N_7095);
or U8119 (N_8119,N_7225,N_7128);
xor U8120 (N_8120,N_7147,N_7171);
nor U8121 (N_8121,N_7142,N_7073);
nand U8122 (N_8122,N_7330,N_7180);
nand U8123 (N_8123,N_7445,N_7423);
or U8124 (N_8124,N_6926,N_7023);
or U8125 (N_8125,N_8029,N_7505);
and U8126 (N_8126,N_7867,N_7745);
nand U8127 (N_8127,N_8002,N_7592);
xor U8128 (N_8128,N_7872,N_7934);
nor U8129 (N_8129,N_7859,N_7705);
and U8130 (N_8130,N_7643,N_7656);
nor U8131 (N_8131,N_8115,N_7980);
nor U8132 (N_8132,N_7988,N_8045);
nor U8133 (N_8133,N_7681,N_7997);
xnor U8134 (N_8134,N_7968,N_7612);
nor U8135 (N_8135,N_7858,N_7640);
nor U8136 (N_8136,N_7668,N_8123);
xor U8137 (N_8137,N_7521,N_7690);
or U8138 (N_8138,N_7911,N_7599);
or U8139 (N_8139,N_7834,N_7930);
nand U8140 (N_8140,N_7605,N_8052);
nand U8141 (N_8141,N_7927,N_7685);
nor U8142 (N_8142,N_7562,N_7869);
or U8143 (N_8143,N_8094,N_8116);
and U8144 (N_8144,N_7670,N_7862);
nand U8145 (N_8145,N_7851,N_7765);
nand U8146 (N_8146,N_7866,N_7757);
or U8147 (N_8147,N_8012,N_8032);
xor U8148 (N_8148,N_8005,N_7642);
or U8149 (N_8149,N_7926,N_7766);
or U8150 (N_8150,N_7913,N_7828);
nand U8151 (N_8151,N_7616,N_7707);
xor U8152 (N_8152,N_7792,N_7751);
nand U8153 (N_8153,N_7929,N_8073);
and U8154 (N_8154,N_7966,N_7735);
nor U8155 (N_8155,N_7641,N_8118);
nor U8156 (N_8156,N_7910,N_7830);
nor U8157 (N_8157,N_8086,N_7512);
nor U8158 (N_8158,N_7931,N_7507);
nor U8159 (N_8159,N_7701,N_8081);
and U8160 (N_8160,N_8063,N_7710);
and U8161 (N_8161,N_7838,N_7879);
nor U8162 (N_8162,N_8098,N_7763);
xnor U8163 (N_8163,N_7993,N_7970);
nor U8164 (N_8164,N_8004,N_8117);
nor U8165 (N_8165,N_8064,N_7938);
nand U8166 (N_8166,N_7882,N_8077);
or U8167 (N_8167,N_7808,N_7714);
xor U8168 (N_8168,N_7983,N_7753);
nor U8169 (N_8169,N_8107,N_7853);
nor U8170 (N_8170,N_7939,N_8104);
or U8171 (N_8171,N_7564,N_7604);
nor U8172 (N_8172,N_7624,N_7613);
nand U8173 (N_8173,N_7919,N_7550);
nor U8174 (N_8174,N_7947,N_7885);
nor U8175 (N_8175,N_7807,N_7504);
xnor U8176 (N_8176,N_7796,N_8022);
or U8177 (N_8177,N_7734,N_7536);
nor U8178 (N_8178,N_7845,N_7533);
xnor U8179 (N_8179,N_8120,N_7769);
nand U8180 (N_8180,N_7799,N_7894);
xnor U8181 (N_8181,N_7991,N_7633);
or U8182 (N_8182,N_7958,N_7703);
nor U8183 (N_8183,N_8001,N_7779);
nor U8184 (N_8184,N_7918,N_7595);
nor U8185 (N_8185,N_7875,N_7951);
nor U8186 (N_8186,N_7777,N_7678);
and U8187 (N_8187,N_7606,N_7709);
nand U8188 (N_8188,N_7530,N_8097);
nand U8189 (N_8189,N_7547,N_7649);
nand U8190 (N_8190,N_7909,N_7551);
nand U8191 (N_8191,N_7596,N_8071);
or U8192 (N_8192,N_7684,N_8099);
or U8193 (N_8193,N_7713,N_8056);
or U8194 (N_8194,N_8042,N_7806);
and U8195 (N_8195,N_7812,N_7933);
nor U8196 (N_8196,N_8011,N_7733);
xnor U8197 (N_8197,N_8016,N_7586);
xnor U8198 (N_8198,N_7590,N_7514);
xor U8199 (N_8199,N_7750,N_7657);
nand U8200 (N_8200,N_7601,N_7591);
nor U8201 (N_8201,N_7546,N_7863);
xor U8202 (N_8202,N_7767,N_7925);
nand U8203 (N_8203,N_7669,N_7688);
nand U8204 (N_8204,N_7961,N_7627);
nor U8205 (N_8205,N_7956,N_7946);
or U8206 (N_8206,N_7732,N_8083);
or U8207 (N_8207,N_7542,N_8106);
or U8208 (N_8208,N_7888,N_7996);
and U8209 (N_8209,N_8088,N_7865);
and U8210 (N_8210,N_7602,N_7520);
xnor U8211 (N_8211,N_7600,N_7772);
and U8212 (N_8212,N_7936,N_7902);
nor U8213 (N_8213,N_7771,N_7538);
nor U8214 (N_8214,N_8044,N_7708);
xnor U8215 (N_8215,N_7664,N_7691);
xnor U8216 (N_8216,N_7809,N_7724);
xor U8217 (N_8217,N_7746,N_7680);
xor U8218 (N_8218,N_7963,N_7857);
xnor U8219 (N_8219,N_8096,N_7923);
and U8220 (N_8220,N_7575,N_7658);
nor U8221 (N_8221,N_7972,N_7741);
xor U8222 (N_8222,N_7572,N_7976);
and U8223 (N_8223,N_7556,N_7854);
xor U8224 (N_8224,N_8006,N_7916);
nand U8225 (N_8225,N_7742,N_7775);
nand U8226 (N_8226,N_7646,N_7846);
nor U8227 (N_8227,N_8110,N_7560);
nand U8228 (N_8228,N_7700,N_7903);
or U8229 (N_8229,N_7768,N_7841);
nor U8230 (N_8230,N_7573,N_7842);
and U8231 (N_8231,N_8100,N_7905);
nand U8232 (N_8232,N_7644,N_7529);
nor U8233 (N_8233,N_7557,N_7881);
xor U8234 (N_8234,N_7873,N_7503);
and U8235 (N_8235,N_7712,N_8112);
xor U8236 (N_8236,N_7860,N_7890);
xnor U8237 (N_8237,N_7623,N_7886);
and U8238 (N_8238,N_7543,N_7937);
xor U8239 (N_8239,N_7718,N_8050);
and U8240 (N_8240,N_7528,N_7728);
and U8241 (N_8241,N_7810,N_8075);
nor U8242 (N_8242,N_7719,N_7813);
nor U8243 (N_8243,N_7539,N_7797);
nor U8244 (N_8244,N_7566,N_8010);
and U8245 (N_8245,N_7762,N_7588);
xor U8246 (N_8246,N_7548,N_7897);
nor U8247 (N_8247,N_8019,N_7935);
nand U8248 (N_8248,N_7944,N_7725);
and U8249 (N_8249,N_8007,N_7655);
and U8250 (N_8250,N_7698,N_7518);
nand U8251 (N_8251,N_7949,N_8122);
nand U8252 (N_8252,N_7662,N_7508);
and U8253 (N_8253,N_7686,N_7693);
and U8254 (N_8254,N_7626,N_8092);
and U8255 (N_8255,N_8066,N_7598);
nor U8256 (N_8256,N_7695,N_7738);
xnor U8257 (N_8257,N_7977,N_7790);
or U8258 (N_8258,N_7821,N_7515);
nand U8259 (N_8259,N_7585,N_7801);
and U8260 (N_8260,N_7984,N_7583);
xnor U8261 (N_8261,N_8062,N_7831);
and U8262 (N_8262,N_7803,N_8085);
nor U8263 (N_8263,N_7786,N_7893);
xor U8264 (N_8264,N_8111,N_7755);
or U8265 (N_8265,N_7877,N_8095);
or U8266 (N_8266,N_8072,N_8082);
or U8267 (N_8267,N_7697,N_7511);
nor U8268 (N_8268,N_7534,N_7904);
xor U8269 (N_8269,N_7816,N_7773);
nand U8270 (N_8270,N_7565,N_7593);
xnor U8271 (N_8271,N_8058,N_7694);
xor U8272 (N_8272,N_7739,N_8008);
or U8273 (N_8273,N_7513,N_7780);
and U8274 (N_8274,N_7761,N_7558);
or U8275 (N_8275,N_7615,N_7722);
xnor U8276 (N_8276,N_7782,N_7822);
and U8277 (N_8277,N_8039,N_8087);
and U8278 (N_8278,N_7985,N_7617);
xnor U8279 (N_8279,N_7594,N_7577);
xnor U8280 (N_8280,N_7990,N_8105);
or U8281 (N_8281,N_7764,N_7844);
nand U8282 (N_8282,N_7884,N_8003);
or U8283 (N_8283,N_7638,N_7667);
and U8284 (N_8284,N_7524,N_7544);
nor U8285 (N_8285,N_8074,N_8035);
nor U8286 (N_8286,N_7715,N_8047);
xor U8287 (N_8287,N_7908,N_7915);
or U8288 (N_8288,N_7829,N_7942);
nand U8289 (N_8289,N_7648,N_8114);
or U8290 (N_8290,N_7843,N_7945);
xnor U8291 (N_8291,N_7981,N_7948);
nor U8292 (N_8292,N_7721,N_7836);
and U8293 (N_8293,N_7620,N_7653);
or U8294 (N_8294,N_7986,N_7517);
and U8295 (N_8295,N_7943,N_7759);
nor U8296 (N_8296,N_8014,N_7537);
nand U8297 (N_8297,N_7749,N_7509);
or U8298 (N_8298,N_7621,N_7540);
and U8299 (N_8299,N_7832,N_7614);
nor U8300 (N_8300,N_7630,N_7785);
xor U8301 (N_8301,N_7635,N_7979);
and U8302 (N_8302,N_8000,N_7969);
xnor U8303 (N_8303,N_7964,N_7849);
or U8304 (N_8304,N_7576,N_7898);
and U8305 (N_8305,N_7663,N_8015);
nor U8306 (N_8306,N_7567,N_8018);
nor U8307 (N_8307,N_7580,N_7752);
nor U8308 (N_8308,N_8060,N_7597);
or U8309 (N_8309,N_8051,N_7848);
nand U8310 (N_8310,N_7650,N_7696);
or U8311 (N_8311,N_7629,N_7502);
or U8312 (N_8312,N_7868,N_7870);
xor U8313 (N_8313,N_7794,N_7744);
or U8314 (N_8314,N_8067,N_7525);
or U8315 (N_8315,N_7609,N_7727);
nand U8316 (N_8316,N_7535,N_7571);
or U8317 (N_8317,N_7819,N_7864);
nor U8318 (N_8318,N_7804,N_8069);
nand U8319 (N_8319,N_7631,N_7561);
or U8320 (N_8320,N_7820,N_7555);
or U8321 (N_8321,N_8053,N_7527);
xnor U8322 (N_8322,N_7673,N_7895);
or U8323 (N_8323,N_8038,N_8026);
nand U8324 (N_8324,N_7754,N_7523);
nor U8325 (N_8325,N_7774,N_7999);
or U8326 (N_8326,N_7954,N_7639);
and U8327 (N_8327,N_7559,N_7675);
xor U8328 (N_8328,N_7652,N_8048);
nor U8329 (N_8329,N_7871,N_7815);
nor U8330 (N_8330,N_7682,N_7574);
xnor U8331 (N_8331,N_7516,N_7920);
nor U8332 (N_8332,N_7581,N_7798);
nand U8333 (N_8333,N_8084,N_7940);
nand U8334 (N_8334,N_7553,N_7619);
nor U8335 (N_8335,N_7628,N_8080);
nor U8336 (N_8336,N_8030,N_7827);
or U8337 (N_8337,N_7730,N_7967);
and U8338 (N_8338,N_7634,N_7998);
nor U8339 (N_8339,N_8090,N_7907);
and U8340 (N_8340,N_7955,N_7659);
nand U8341 (N_8341,N_7510,N_8049);
nor U8342 (N_8342,N_7784,N_7729);
nor U8343 (N_8343,N_7717,N_8013);
xnor U8344 (N_8344,N_8057,N_8070);
xnor U8345 (N_8345,N_8079,N_7971);
nor U8346 (N_8346,N_7906,N_7924);
xnor U8347 (N_8347,N_7687,N_7587);
xor U8348 (N_8348,N_7824,N_7519);
nor U8349 (N_8349,N_8043,N_8102);
nand U8350 (N_8350,N_7672,N_8119);
nand U8351 (N_8351,N_7541,N_7770);
and U8352 (N_8352,N_7787,N_7526);
xnor U8353 (N_8353,N_7552,N_7950);
or U8354 (N_8354,N_8027,N_7778);
and U8355 (N_8355,N_7665,N_8041);
xor U8356 (N_8356,N_7975,N_7711);
nand U8357 (N_8357,N_7800,N_7569);
nor U8358 (N_8358,N_7758,N_7720);
or U8359 (N_8359,N_7532,N_7833);
or U8360 (N_8360,N_8121,N_7899);
nand U8361 (N_8361,N_7837,N_7953);
or U8362 (N_8362,N_8009,N_7699);
or U8363 (N_8363,N_7660,N_8113);
and U8364 (N_8364,N_7531,N_7878);
xnor U8365 (N_8365,N_8020,N_8031);
or U8366 (N_8366,N_7666,N_7932);
or U8367 (N_8367,N_7570,N_7716);
nand U8368 (N_8368,N_8033,N_8124);
xor U8369 (N_8369,N_7995,N_7989);
and U8370 (N_8370,N_7625,N_7723);
nor U8371 (N_8371,N_7802,N_8046);
nand U8372 (N_8372,N_7982,N_7579);
nor U8373 (N_8373,N_7994,N_8078);
or U8374 (N_8374,N_7793,N_7689);
and U8375 (N_8375,N_7957,N_7637);
nand U8376 (N_8376,N_7611,N_7776);
nand U8377 (N_8377,N_7651,N_7789);
or U8378 (N_8378,N_7880,N_7737);
and U8379 (N_8379,N_7607,N_7545);
and U8380 (N_8380,N_7760,N_7563);
and U8381 (N_8381,N_8024,N_7568);
xnor U8382 (N_8382,N_7679,N_8017);
or U8383 (N_8383,N_7900,N_8101);
and U8384 (N_8384,N_7965,N_8021);
nand U8385 (N_8385,N_7952,N_8028);
nand U8386 (N_8386,N_8055,N_7676);
and U8387 (N_8387,N_7582,N_7636);
nand U8388 (N_8388,N_7856,N_7781);
and U8389 (N_8389,N_7839,N_8040);
xor U8390 (N_8390,N_7960,N_7610);
or U8391 (N_8391,N_7941,N_7921);
and U8392 (N_8392,N_7726,N_7855);
nor U8393 (N_8393,N_8068,N_7817);
nor U8394 (N_8394,N_7811,N_8034);
and U8395 (N_8395,N_7840,N_7818);
and U8396 (N_8396,N_7835,N_7874);
nor U8397 (N_8397,N_7795,N_7522);
or U8398 (N_8398,N_7743,N_7974);
or U8399 (N_8399,N_7683,N_8065);
nand U8400 (N_8400,N_7825,N_7740);
or U8401 (N_8401,N_8025,N_7692);
nand U8402 (N_8402,N_7992,N_7674);
and U8403 (N_8403,N_7671,N_7661);
or U8404 (N_8404,N_7645,N_7584);
xnor U8405 (N_8405,N_8061,N_7883);
nand U8406 (N_8406,N_7962,N_7747);
or U8407 (N_8407,N_7706,N_7677);
xnor U8408 (N_8408,N_7861,N_7731);
and U8409 (N_8409,N_8059,N_7736);
nand U8410 (N_8410,N_7632,N_8054);
nor U8411 (N_8411,N_8076,N_8023);
or U8412 (N_8412,N_7914,N_7876);
and U8413 (N_8413,N_7654,N_7917);
nor U8414 (N_8414,N_7501,N_7702);
and U8415 (N_8415,N_7896,N_7887);
and U8416 (N_8416,N_7889,N_7901);
xnor U8417 (N_8417,N_7850,N_8109);
nor U8418 (N_8418,N_7622,N_8089);
xor U8419 (N_8419,N_7892,N_7618);
xnor U8420 (N_8420,N_7788,N_7928);
and U8421 (N_8421,N_7814,N_7891);
xnor U8422 (N_8422,N_8093,N_8103);
nor U8423 (N_8423,N_8091,N_7978);
or U8424 (N_8424,N_7554,N_7647);
or U8425 (N_8425,N_7847,N_8108);
xor U8426 (N_8426,N_7756,N_7589);
or U8427 (N_8427,N_8036,N_7748);
and U8428 (N_8428,N_7959,N_7912);
or U8429 (N_8429,N_7987,N_8037);
or U8430 (N_8430,N_7506,N_7922);
or U8431 (N_8431,N_7500,N_7973);
and U8432 (N_8432,N_7852,N_7826);
xnor U8433 (N_8433,N_7549,N_7791);
or U8434 (N_8434,N_7608,N_7783);
and U8435 (N_8435,N_7578,N_7603);
xnor U8436 (N_8436,N_7805,N_7704);
nor U8437 (N_8437,N_7823,N_8039);
nor U8438 (N_8438,N_7530,N_8114);
and U8439 (N_8439,N_7887,N_8016);
nand U8440 (N_8440,N_7524,N_7522);
nor U8441 (N_8441,N_7600,N_8032);
and U8442 (N_8442,N_7647,N_7572);
nor U8443 (N_8443,N_7876,N_7709);
nor U8444 (N_8444,N_8076,N_7520);
and U8445 (N_8445,N_7976,N_7748);
nand U8446 (N_8446,N_7811,N_7816);
and U8447 (N_8447,N_7746,N_8056);
nand U8448 (N_8448,N_8108,N_7891);
nand U8449 (N_8449,N_7819,N_7640);
or U8450 (N_8450,N_7650,N_7990);
nor U8451 (N_8451,N_7978,N_7726);
nor U8452 (N_8452,N_7791,N_7748);
nand U8453 (N_8453,N_7521,N_7750);
nor U8454 (N_8454,N_7669,N_7598);
nor U8455 (N_8455,N_7897,N_7577);
or U8456 (N_8456,N_7529,N_7770);
or U8457 (N_8457,N_8039,N_7772);
and U8458 (N_8458,N_7632,N_8002);
nand U8459 (N_8459,N_7854,N_7677);
and U8460 (N_8460,N_7613,N_7799);
and U8461 (N_8461,N_7741,N_8071);
and U8462 (N_8462,N_8077,N_8048);
and U8463 (N_8463,N_7582,N_7940);
or U8464 (N_8464,N_8015,N_8114);
xor U8465 (N_8465,N_7717,N_7910);
and U8466 (N_8466,N_8106,N_8087);
nor U8467 (N_8467,N_8071,N_7603);
xor U8468 (N_8468,N_7575,N_8077);
or U8469 (N_8469,N_7828,N_7850);
nor U8470 (N_8470,N_7891,N_8028);
nand U8471 (N_8471,N_7505,N_7803);
and U8472 (N_8472,N_7982,N_7907);
nor U8473 (N_8473,N_7941,N_7859);
and U8474 (N_8474,N_7719,N_8063);
and U8475 (N_8475,N_7588,N_7853);
nand U8476 (N_8476,N_8110,N_7821);
and U8477 (N_8477,N_7673,N_7788);
and U8478 (N_8478,N_7802,N_8107);
nor U8479 (N_8479,N_7605,N_7710);
nor U8480 (N_8480,N_7508,N_7782);
and U8481 (N_8481,N_7630,N_8062);
nand U8482 (N_8482,N_7593,N_7748);
xnor U8483 (N_8483,N_7776,N_7521);
xnor U8484 (N_8484,N_7847,N_7867);
xnor U8485 (N_8485,N_8009,N_7644);
nand U8486 (N_8486,N_7944,N_7560);
and U8487 (N_8487,N_8064,N_7773);
nand U8488 (N_8488,N_7655,N_7888);
or U8489 (N_8489,N_7672,N_7721);
xor U8490 (N_8490,N_8075,N_7946);
or U8491 (N_8491,N_7520,N_7816);
or U8492 (N_8492,N_7516,N_7865);
nand U8493 (N_8493,N_7884,N_8022);
nand U8494 (N_8494,N_7994,N_7739);
or U8495 (N_8495,N_8117,N_7709);
or U8496 (N_8496,N_7892,N_7639);
nor U8497 (N_8497,N_7933,N_8120);
or U8498 (N_8498,N_7893,N_8066);
or U8499 (N_8499,N_7830,N_8102);
or U8500 (N_8500,N_8065,N_7898);
nor U8501 (N_8501,N_8055,N_7677);
or U8502 (N_8502,N_8018,N_7559);
nor U8503 (N_8503,N_8071,N_7554);
xnor U8504 (N_8504,N_7628,N_7908);
nand U8505 (N_8505,N_7812,N_7702);
and U8506 (N_8506,N_8052,N_7505);
nand U8507 (N_8507,N_7847,N_7707);
xor U8508 (N_8508,N_7826,N_7962);
nor U8509 (N_8509,N_7909,N_8054);
and U8510 (N_8510,N_8033,N_7590);
nand U8511 (N_8511,N_7738,N_7698);
nand U8512 (N_8512,N_7843,N_7846);
nand U8513 (N_8513,N_8087,N_7958);
nor U8514 (N_8514,N_7647,N_7932);
nor U8515 (N_8515,N_8052,N_7633);
or U8516 (N_8516,N_7673,N_7718);
nor U8517 (N_8517,N_7739,N_7605);
nand U8518 (N_8518,N_7532,N_7989);
and U8519 (N_8519,N_7500,N_7744);
xor U8520 (N_8520,N_8016,N_7935);
and U8521 (N_8521,N_7698,N_7506);
nor U8522 (N_8522,N_7560,N_7671);
xor U8523 (N_8523,N_8005,N_7910);
and U8524 (N_8524,N_7654,N_7797);
xnor U8525 (N_8525,N_7750,N_7733);
and U8526 (N_8526,N_7919,N_7673);
xnor U8527 (N_8527,N_7567,N_7970);
and U8528 (N_8528,N_8019,N_7945);
or U8529 (N_8529,N_7505,N_8122);
nor U8530 (N_8530,N_8032,N_8109);
nor U8531 (N_8531,N_8087,N_7995);
and U8532 (N_8532,N_8040,N_7601);
nor U8533 (N_8533,N_8006,N_7813);
and U8534 (N_8534,N_7504,N_7928);
and U8535 (N_8535,N_7516,N_7518);
xor U8536 (N_8536,N_7837,N_7705);
nor U8537 (N_8537,N_7889,N_7676);
nor U8538 (N_8538,N_7754,N_7554);
or U8539 (N_8539,N_7860,N_7743);
and U8540 (N_8540,N_7883,N_7884);
nand U8541 (N_8541,N_7647,N_8080);
or U8542 (N_8542,N_7911,N_7904);
xnor U8543 (N_8543,N_7568,N_8022);
xor U8544 (N_8544,N_7904,N_7957);
nand U8545 (N_8545,N_7892,N_8064);
nor U8546 (N_8546,N_7508,N_7999);
xor U8547 (N_8547,N_7780,N_7708);
xnor U8548 (N_8548,N_7617,N_7766);
nand U8549 (N_8549,N_7521,N_8065);
or U8550 (N_8550,N_8060,N_8087);
nor U8551 (N_8551,N_7726,N_8001);
and U8552 (N_8552,N_7632,N_7761);
xnor U8553 (N_8553,N_7507,N_7551);
xor U8554 (N_8554,N_7969,N_7691);
or U8555 (N_8555,N_7704,N_8054);
and U8556 (N_8556,N_7568,N_7825);
nor U8557 (N_8557,N_7510,N_7920);
xnor U8558 (N_8558,N_7826,N_8010);
xor U8559 (N_8559,N_7768,N_7759);
nor U8560 (N_8560,N_7745,N_7968);
nand U8561 (N_8561,N_7614,N_7751);
nand U8562 (N_8562,N_7747,N_7663);
and U8563 (N_8563,N_8028,N_7552);
nor U8564 (N_8564,N_7899,N_8085);
nand U8565 (N_8565,N_7800,N_7734);
or U8566 (N_8566,N_8079,N_7926);
xnor U8567 (N_8567,N_7652,N_8028);
and U8568 (N_8568,N_8009,N_7930);
nor U8569 (N_8569,N_7715,N_7613);
nand U8570 (N_8570,N_7777,N_7654);
nor U8571 (N_8571,N_7938,N_7578);
nand U8572 (N_8572,N_7668,N_7954);
nand U8573 (N_8573,N_8073,N_7627);
and U8574 (N_8574,N_8056,N_8111);
nand U8575 (N_8575,N_8031,N_7949);
and U8576 (N_8576,N_7997,N_7525);
or U8577 (N_8577,N_7678,N_7614);
xor U8578 (N_8578,N_7784,N_7669);
nand U8579 (N_8579,N_7787,N_7936);
xor U8580 (N_8580,N_7633,N_7892);
or U8581 (N_8581,N_7513,N_7979);
nand U8582 (N_8582,N_7687,N_7595);
nor U8583 (N_8583,N_8051,N_7911);
or U8584 (N_8584,N_7515,N_7872);
xnor U8585 (N_8585,N_7777,N_8003);
or U8586 (N_8586,N_7935,N_7784);
or U8587 (N_8587,N_7849,N_7917);
nor U8588 (N_8588,N_8034,N_7724);
nor U8589 (N_8589,N_8047,N_7546);
or U8590 (N_8590,N_7929,N_7725);
or U8591 (N_8591,N_7785,N_7744);
nand U8592 (N_8592,N_7924,N_8046);
or U8593 (N_8593,N_8109,N_7838);
xor U8594 (N_8594,N_7971,N_8083);
nor U8595 (N_8595,N_7573,N_8022);
xor U8596 (N_8596,N_7817,N_8092);
or U8597 (N_8597,N_7863,N_7853);
or U8598 (N_8598,N_7605,N_7654);
or U8599 (N_8599,N_8074,N_7799);
nand U8600 (N_8600,N_7822,N_8026);
xor U8601 (N_8601,N_8011,N_8031);
or U8602 (N_8602,N_7989,N_7522);
and U8603 (N_8603,N_7715,N_7977);
nand U8604 (N_8604,N_8034,N_7956);
nor U8605 (N_8605,N_8090,N_7978);
or U8606 (N_8606,N_7987,N_7685);
nand U8607 (N_8607,N_7599,N_7954);
xor U8608 (N_8608,N_7724,N_8089);
or U8609 (N_8609,N_7661,N_7697);
and U8610 (N_8610,N_7542,N_7609);
nand U8611 (N_8611,N_7724,N_8045);
nor U8612 (N_8612,N_7982,N_7753);
xor U8613 (N_8613,N_7880,N_7885);
or U8614 (N_8614,N_7781,N_7577);
nor U8615 (N_8615,N_7512,N_7734);
and U8616 (N_8616,N_7845,N_7968);
nand U8617 (N_8617,N_7842,N_7630);
xnor U8618 (N_8618,N_7857,N_7577);
or U8619 (N_8619,N_7702,N_7881);
and U8620 (N_8620,N_8052,N_8012);
or U8621 (N_8621,N_7800,N_8078);
nand U8622 (N_8622,N_8030,N_7851);
nor U8623 (N_8623,N_7853,N_7919);
and U8624 (N_8624,N_7741,N_7721);
nand U8625 (N_8625,N_7812,N_7755);
nand U8626 (N_8626,N_7795,N_7569);
nand U8627 (N_8627,N_7746,N_7500);
xnor U8628 (N_8628,N_8068,N_7500);
xnor U8629 (N_8629,N_7720,N_7914);
nand U8630 (N_8630,N_7921,N_7958);
nor U8631 (N_8631,N_8101,N_7990);
xor U8632 (N_8632,N_7892,N_7985);
xnor U8633 (N_8633,N_7717,N_7658);
and U8634 (N_8634,N_7923,N_7642);
or U8635 (N_8635,N_7605,N_7854);
nand U8636 (N_8636,N_7674,N_7881);
nand U8637 (N_8637,N_7685,N_7749);
nor U8638 (N_8638,N_7869,N_7956);
or U8639 (N_8639,N_7539,N_7529);
xor U8640 (N_8640,N_8064,N_7605);
and U8641 (N_8641,N_7554,N_8065);
nor U8642 (N_8642,N_7528,N_7775);
nand U8643 (N_8643,N_7841,N_7853);
xnor U8644 (N_8644,N_7511,N_7732);
xnor U8645 (N_8645,N_7504,N_7898);
xor U8646 (N_8646,N_7725,N_7503);
xor U8647 (N_8647,N_7580,N_7704);
nand U8648 (N_8648,N_7865,N_8018);
nor U8649 (N_8649,N_7816,N_7718);
nand U8650 (N_8650,N_8111,N_7665);
nand U8651 (N_8651,N_7786,N_7914);
nor U8652 (N_8652,N_7828,N_7899);
or U8653 (N_8653,N_7528,N_7552);
nor U8654 (N_8654,N_8072,N_7552);
or U8655 (N_8655,N_7560,N_7759);
or U8656 (N_8656,N_8029,N_7622);
or U8657 (N_8657,N_7699,N_7563);
xnor U8658 (N_8658,N_7763,N_8108);
nand U8659 (N_8659,N_7895,N_7668);
or U8660 (N_8660,N_8112,N_8015);
xor U8661 (N_8661,N_7837,N_7635);
nand U8662 (N_8662,N_8031,N_7946);
and U8663 (N_8663,N_7755,N_7805);
and U8664 (N_8664,N_7938,N_7908);
nor U8665 (N_8665,N_7714,N_7512);
xor U8666 (N_8666,N_7891,N_7914);
and U8667 (N_8667,N_7856,N_7708);
or U8668 (N_8668,N_7892,N_7969);
xor U8669 (N_8669,N_7724,N_7563);
and U8670 (N_8670,N_8089,N_8054);
xnor U8671 (N_8671,N_7699,N_8050);
and U8672 (N_8672,N_7856,N_7565);
and U8673 (N_8673,N_7712,N_7938);
or U8674 (N_8674,N_7955,N_7581);
and U8675 (N_8675,N_7501,N_7863);
xnor U8676 (N_8676,N_7881,N_7825);
xor U8677 (N_8677,N_7595,N_8019);
xor U8678 (N_8678,N_7609,N_7830);
xnor U8679 (N_8679,N_8072,N_7992);
nor U8680 (N_8680,N_7977,N_7975);
xnor U8681 (N_8681,N_7776,N_7949);
xnor U8682 (N_8682,N_8038,N_7738);
nor U8683 (N_8683,N_7510,N_7650);
and U8684 (N_8684,N_8084,N_7675);
xor U8685 (N_8685,N_7985,N_7980);
nor U8686 (N_8686,N_7847,N_7632);
and U8687 (N_8687,N_7743,N_7792);
and U8688 (N_8688,N_8109,N_7662);
xor U8689 (N_8689,N_7928,N_7828);
or U8690 (N_8690,N_7621,N_7894);
xnor U8691 (N_8691,N_7708,N_7694);
and U8692 (N_8692,N_7917,N_8007);
nor U8693 (N_8693,N_7578,N_8089);
nand U8694 (N_8694,N_7946,N_7521);
nor U8695 (N_8695,N_7684,N_8118);
nor U8696 (N_8696,N_7961,N_7573);
or U8697 (N_8697,N_7699,N_8052);
xor U8698 (N_8698,N_7599,N_7692);
nand U8699 (N_8699,N_8046,N_7973);
xnor U8700 (N_8700,N_7903,N_8118);
nand U8701 (N_8701,N_7740,N_7990);
and U8702 (N_8702,N_7597,N_7936);
and U8703 (N_8703,N_8033,N_7524);
or U8704 (N_8704,N_7938,N_7534);
xnor U8705 (N_8705,N_7881,N_7929);
and U8706 (N_8706,N_7981,N_8117);
nor U8707 (N_8707,N_7657,N_7985);
nor U8708 (N_8708,N_7864,N_8031);
or U8709 (N_8709,N_7867,N_8109);
nor U8710 (N_8710,N_7765,N_7863);
and U8711 (N_8711,N_7708,N_7696);
nor U8712 (N_8712,N_7909,N_8117);
or U8713 (N_8713,N_8118,N_7955);
nor U8714 (N_8714,N_7569,N_7639);
nor U8715 (N_8715,N_7993,N_7650);
xnor U8716 (N_8716,N_7999,N_7606);
nor U8717 (N_8717,N_7589,N_8096);
nand U8718 (N_8718,N_8059,N_8050);
and U8719 (N_8719,N_7726,N_7559);
nor U8720 (N_8720,N_8119,N_7725);
nand U8721 (N_8721,N_7886,N_7593);
and U8722 (N_8722,N_7593,N_7982);
nand U8723 (N_8723,N_7524,N_7825);
xnor U8724 (N_8724,N_7826,N_7690);
xor U8725 (N_8725,N_7626,N_7584);
nor U8726 (N_8726,N_7824,N_8021);
xor U8727 (N_8727,N_8043,N_7539);
nand U8728 (N_8728,N_7844,N_7574);
or U8729 (N_8729,N_7666,N_7942);
xnor U8730 (N_8730,N_7567,N_7730);
nor U8731 (N_8731,N_7598,N_7746);
and U8732 (N_8732,N_7680,N_7606);
nand U8733 (N_8733,N_7908,N_8111);
nand U8734 (N_8734,N_8051,N_7975);
and U8735 (N_8735,N_8009,N_7606);
xnor U8736 (N_8736,N_7857,N_8018);
nand U8737 (N_8737,N_7884,N_7673);
nand U8738 (N_8738,N_8121,N_7956);
or U8739 (N_8739,N_7866,N_7669);
xor U8740 (N_8740,N_7887,N_7739);
nor U8741 (N_8741,N_7936,N_7964);
nand U8742 (N_8742,N_7582,N_7953);
or U8743 (N_8743,N_8027,N_8029);
xor U8744 (N_8744,N_8020,N_8099);
nor U8745 (N_8745,N_7936,N_7577);
nand U8746 (N_8746,N_7860,N_7586);
nand U8747 (N_8747,N_8044,N_7728);
or U8748 (N_8748,N_7752,N_7641);
or U8749 (N_8749,N_7596,N_7953);
nand U8750 (N_8750,N_8729,N_8213);
xor U8751 (N_8751,N_8377,N_8706);
nand U8752 (N_8752,N_8385,N_8402);
xnor U8753 (N_8753,N_8637,N_8351);
nor U8754 (N_8754,N_8310,N_8180);
xor U8755 (N_8755,N_8391,N_8575);
xnor U8756 (N_8756,N_8307,N_8683);
and U8757 (N_8757,N_8531,N_8263);
nand U8758 (N_8758,N_8185,N_8295);
xnor U8759 (N_8759,N_8326,N_8138);
nor U8760 (N_8760,N_8261,N_8126);
xnor U8761 (N_8761,N_8444,N_8223);
and U8762 (N_8762,N_8217,N_8211);
and U8763 (N_8763,N_8166,N_8409);
xor U8764 (N_8764,N_8288,N_8182);
or U8765 (N_8765,N_8155,N_8458);
nor U8766 (N_8766,N_8141,N_8748);
or U8767 (N_8767,N_8610,N_8544);
xnor U8768 (N_8768,N_8227,N_8538);
and U8769 (N_8769,N_8313,N_8499);
xnor U8770 (N_8770,N_8417,N_8736);
or U8771 (N_8771,N_8718,N_8202);
nand U8772 (N_8772,N_8507,N_8215);
xor U8773 (N_8773,N_8557,N_8521);
and U8774 (N_8774,N_8431,N_8560);
and U8775 (N_8775,N_8262,N_8194);
nor U8776 (N_8776,N_8308,N_8614);
nand U8777 (N_8777,N_8206,N_8594);
nand U8778 (N_8778,N_8135,N_8269);
nand U8779 (N_8779,N_8635,N_8707);
xor U8780 (N_8780,N_8519,N_8245);
xor U8781 (N_8781,N_8636,N_8484);
and U8782 (N_8782,N_8148,N_8320);
nor U8783 (N_8783,N_8568,N_8670);
nand U8784 (N_8784,N_8451,N_8655);
nor U8785 (N_8785,N_8429,N_8410);
or U8786 (N_8786,N_8586,N_8401);
xor U8787 (N_8787,N_8724,N_8510);
and U8788 (N_8788,N_8495,N_8475);
xnor U8789 (N_8789,N_8192,N_8183);
nor U8790 (N_8790,N_8381,N_8622);
nand U8791 (N_8791,N_8321,N_8243);
xnor U8792 (N_8792,N_8570,N_8149);
nand U8793 (N_8793,N_8527,N_8144);
nand U8794 (N_8794,N_8201,N_8668);
nor U8795 (N_8795,N_8592,N_8450);
and U8796 (N_8796,N_8547,N_8246);
xor U8797 (N_8797,N_8546,N_8745);
and U8798 (N_8798,N_8616,N_8386);
nand U8799 (N_8799,N_8419,N_8690);
nor U8800 (N_8800,N_8593,N_8222);
or U8801 (N_8801,N_8688,N_8405);
or U8802 (N_8802,N_8198,N_8604);
nor U8803 (N_8803,N_8699,N_8721);
xnor U8804 (N_8804,N_8168,N_8464);
xor U8805 (N_8805,N_8530,N_8711);
and U8806 (N_8806,N_8717,N_8383);
and U8807 (N_8807,N_8642,N_8139);
nand U8808 (N_8808,N_8504,N_8657);
nor U8809 (N_8809,N_8150,N_8145);
and U8810 (N_8810,N_8459,N_8669);
or U8811 (N_8811,N_8129,N_8533);
xor U8812 (N_8812,N_8463,N_8329);
xnor U8813 (N_8813,N_8481,N_8333);
nor U8814 (N_8814,N_8188,N_8249);
nor U8815 (N_8815,N_8382,N_8306);
or U8816 (N_8816,N_8432,N_8633);
and U8817 (N_8817,N_8700,N_8467);
xnor U8818 (N_8818,N_8389,N_8644);
nor U8819 (N_8819,N_8453,N_8500);
or U8820 (N_8820,N_8485,N_8366);
nand U8821 (N_8821,N_8457,N_8371);
xor U8822 (N_8822,N_8181,N_8653);
or U8823 (N_8823,N_8302,N_8415);
or U8824 (N_8824,N_8733,N_8572);
and U8825 (N_8825,N_8131,N_8638);
nand U8826 (N_8826,N_8392,N_8318);
or U8827 (N_8827,N_8742,N_8259);
nor U8828 (N_8828,N_8523,N_8403);
and U8829 (N_8829,N_8679,N_8618);
and U8830 (N_8830,N_8501,N_8399);
xnor U8831 (N_8831,N_8734,N_8137);
or U8832 (N_8832,N_8551,N_8577);
or U8833 (N_8833,N_8713,N_8229);
or U8834 (N_8834,N_8210,N_8502);
and U8835 (N_8835,N_8353,N_8579);
nand U8836 (N_8836,N_8589,N_8542);
and U8837 (N_8837,N_8199,N_8257);
nor U8838 (N_8838,N_8341,N_8271);
nor U8839 (N_8839,N_8611,N_8230);
xor U8840 (N_8840,N_8225,N_8516);
or U8841 (N_8841,N_8446,N_8541);
or U8842 (N_8842,N_8413,N_8605);
and U8843 (N_8843,N_8489,N_8665);
or U8844 (N_8844,N_8440,N_8556);
or U8845 (N_8845,N_8497,N_8619);
or U8846 (N_8846,N_8553,N_8704);
nor U8847 (N_8847,N_8494,N_8651);
and U8848 (N_8848,N_8473,N_8612);
nor U8849 (N_8849,N_8449,N_8294);
nor U8850 (N_8850,N_8498,N_8411);
nor U8851 (N_8851,N_8387,N_8634);
xnor U8852 (N_8852,N_8581,N_8408);
nand U8853 (N_8853,N_8646,N_8241);
nor U8854 (N_8854,N_8443,N_8599);
nand U8855 (N_8855,N_8208,N_8357);
nor U8856 (N_8856,N_8393,N_8349);
and U8857 (N_8857,N_8514,N_8746);
nor U8858 (N_8858,N_8284,N_8375);
xor U8859 (N_8859,N_8370,N_8445);
and U8860 (N_8860,N_8532,N_8674);
nand U8861 (N_8861,N_8332,N_8477);
and U8862 (N_8862,N_8480,N_8520);
and U8863 (N_8863,N_8508,N_8396);
nand U8864 (N_8864,N_8133,N_8434);
or U8865 (N_8865,N_8348,N_8325);
xnor U8866 (N_8866,N_8379,N_8278);
xnor U8867 (N_8867,N_8735,N_8731);
and U8868 (N_8868,N_8256,N_8394);
nand U8869 (N_8869,N_8142,N_8338);
nand U8870 (N_8870,N_8174,N_8276);
or U8871 (N_8871,N_8555,N_8491);
xor U8872 (N_8872,N_8407,N_8730);
nand U8873 (N_8873,N_8462,N_8558);
nand U8874 (N_8874,N_8291,N_8191);
xnor U8875 (N_8875,N_8146,N_8441);
nand U8876 (N_8876,N_8672,N_8661);
and U8877 (N_8877,N_8265,N_8696);
nor U8878 (N_8878,N_8219,N_8388);
and U8879 (N_8879,N_8378,N_8728);
xnor U8880 (N_8880,N_8512,N_8316);
nor U8881 (N_8881,N_8554,N_8630);
nand U8882 (N_8882,N_8285,N_8304);
xor U8883 (N_8883,N_8430,N_8582);
nor U8884 (N_8884,N_8452,N_8334);
or U8885 (N_8885,N_8648,N_8597);
or U8886 (N_8886,N_8226,N_8303);
and U8887 (N_8887,N_8352,N_8539);
or U8888 (N_8888,N_8177,N_8479);
xnor U8889 (N_8889,N_8345,N_8741);
and U8890 (N_8890,N_8682,N_8626);
or U8891 (N_8891,N_8628,N_8448);
xor U8892 (N_8892,N_8234,N_8273);
and U8893 (N_8893,N_8160,N_8471);
or U8894 (N_8894,N_8296,N_8496);
xnor U8895 (N_8895,N_8505,N_8654);
nand U8896 (N_8896,N_8412,N_8190);
nand U8897 (N_8897,N_8373,N_8209);
nor U8898 (N_8898,N_8606,N_8487);
nor U8899 (N_8899,N_8425,N_8687);
xor U8900 (N_8900,N_8297,N_8216);
nand U8901 (N_8901,N_8358,N_8641);
and U8902 (N_8902,N_8565,N_8561);
and U8903 (N_8903,N_8134,N_8167);
nand U8904 (N_8904,N_8660,N_8433);
and U8905 (N_8905,N_8712,N_8438);
xor U8906 (N_8906,N_8609,N_8571);
or U8907 (N_8907,N_8197,N_8737);
xnor U8908 (N_8908,N_8725,N_8543);
nand U8909 (N_8909,N_8398,N_8684);
and U8910 (N_8910,N_8406,N_8685);
and U8911 (N_8911,N_8580,N_8478);
xnor U8912 (N_8912,N_8221,N_8524);
nor U8913 (N_8913,N_8613,N_8299);
xor U8914 (N_8914,N_8242,N_8354);
nand U8915 (N_8915,N_8355,N_8550);
nor U8916 (N_8916,N_8342,N_8239);
nand U8917 (N_8917,N_8298,N_8418);
xor U8918 (N_8918,N_8335,N_8372);
and U8919 (N_8919,N_8359,N_8629);
xor U8920 (N_8920,N_8689,N_8511);
nand U8921 (N_8921,N_8702,N_8474);
or U8922 (N_8922,N_8603,N_8281);
or U8923 (N_8923,N_8492,N_8136);
nor U8924 (N_8924,N_8339,N_8164);
or U8925 (N_8925,N_8694,N_8368);
and U8926 (N_8926,N_8356,N_8178);
or U8927 (N_8927,N_8266,N_8526);
xor U8928 (N_8928,N_8300,N_8466);
nor U8929 (N_8929,N_8255,N_8749);
nand U8930 (N_8930,N_8390,N_8627);
and U8931 (N_8931,N_8395,N_8469);
nor U8932 (N_8932,N_8143,N_8203);
nand U8933 (N_8933,N_8301,N_8513);
or U8934 (N_8934,N_8360,N_8666);
and U8935 (N_8935,N_8250,N_8678);
and U8936 (N_8936,N_8293,N_8331);
nand U8937 (N_8937,N_8574,N_8639);
nand U8938 (N_8938,N_8218,N_8722);
nand U8939 (N_8939,N_8309,N_8647);
and U8940 (N_8940,N_8552,N_8624);
and U8941 (N_8941,N_8283,N_8128);
xor U8942 (N_8942,N_8472,N_8376);
or U8943 (N_8943,N_8562,N_8156);
nand U8944 (N_8944,N_8343,N_8184);
nor U8945 (N_8945,N_8251,N_8548);
xnor U8946 (N_8946,N_8732,N_8365);
nor U8947 (N_8947,N_8344,N_8468);
or U8948 (N_8948,N_8328,N_8607);
nand U8949 (N_8949,N_8436,N_8153);
or U8950 (N_8950,N_8154,N_8253);
and U8951 (N_8951,N_8187,N_8525);
nand U8952 (N_8952,N_8274,N_8454);
nand U8953 (N_8953,N_8695,N_8374);
nor U8954 (N_8954,N_8640,N_8567);
or U8955 (N_8955,N_8244,N_8286);
nor U8956 (N_8956,N_8709,N_8439);
and U8957 (N_8957,N_8305,N_8214);
xor U8958 (N_8958,N_8127,N_8327);
nor U8959 (N_8959,N_8204,N_8125);
xor U8960 (N_8960,N_8692,N_8727);
nand U8961 (N_8961,N_8726,N_8130);
and U8962 (N_8962,N_8236,N_8559);
xnor U8963 (N_8963,N_8632,N_8189);
and U8964 (N_8964,N_8673,N_8282);
nor U8965 (N_8965,N_8465,N_8659);
and U8966 (N_8966,N_8311,N_8631);
xnor U8967 (N_8967,N_8602,N_8535);
nand U8968 (N_8968,N_8165,N_8264);
nand U8969 (N_8969,N_8260,N_8205);
nor U8970 (N_8970,N_8158,N_8503);
xnor U8971 (N_8971,N_8416,N_8254);
nand U8972 (N_8972,N_8258,N_8220);
xnor U8973 (N_8973,N_8233,N_8228);
xnor U8974 (N_8974,N_8147,N_8171);
nor U8975 (N_8975,N_8705,N_8545);
nor U8976 (N_8976,N_8346,N_8159);
and U8977 (N_8977,N_8714,N_8677);
or U8978 (N_8978,N_8140,N_8238);
nand U8979 (N_8979,N_8330,N_8384);
nand U8980 (N_8980,N_8287,N_8460);
xor U8981 (N_8981,N_8461,N_8176);
nand U8982 (N_8982,N_8723,N_8361);
or U8983 (N_8983,N_8540,N_8625);
and U8984 (N_8984,N_8566,N_8186);
xnor U8985 (N_8985,N_8277,N_8280);
nand U8986 (N_8986,N_8470,N_8601);
or U8987 (N_8987,N_8400,N_8595);
and U8988 (N_8988,N_8650,N_8515);
and U8989 (N_8989,N_8195,N_8573);
and U8990 (N_8990,N_8738,N_8369);
and U8991 (N_8991,N_8350,N_8179);
nand U8992 (N_8992,N_8697,N_8322);
xnor U8993 (N_8993,N_8317,N_8314);
xor U8994 (N_8994,N_8663,N_8272);
or U8995 (N_8995,N_8658,N_8193);
xnor U8996 (N_8996,N_8172,N_8275);
xnor U8997 (N_8997,N_8578,N_8643);
xor U8998 (N_8998,N_8151,N_8740);
nor U8999 (N_8999,N_8232,N_8456);
or U9000 (N_9000,N_8426,N_8267);
and U9001 (N_9001,N_8623,N_8224);
nand U9002 (N_9002,N_8427,N_8157);
or U9003 (N_9003,N_8701,N_8173);
or U9004 (N_9004,N_8170,N_8739);
nand U9005 (N_9005,N_8437,N_8591);
or U9006 (N_9006,N_8621,N_8681);
nor U9007 (N_9007,N_8667,N_8482);
or U9008 (N_9008,N_8200,N_8315);
or U9009 (N_9009,N_8420,N_8649);
or U9010 (N_9010,N_8656,N_8488);
xnor U9011 (N_9011,N_8537,N_8506);
nor U9012 (N_9012,N_8596,N_8585);
xor U9013 (N_9013,N_8652,N_8719);
nand U9014 (N_9014,N_8671,N_8620);
or U9015 (N_9015,N_8698,N_8340);
and U9016 (N_9016,N_8587,N_8645);
nor U9017 (N_9017,N_8536,N_8231);
and U9018 (N_9018,N_8336,N_8615);
and U9019 (N_9019,N_8528,N_8583);
nand U9020 (N_9020,N_8319,N_8292);
and U9021 (N_9021,N_8397,N_8703);
or U9022 (N_9022,N_8509,N_8132);
xor U9023 (N_9023,N_8240,N_8161);
nand U9024 (N_9024,N_8691,N_8347);
or U9025 (N_9025,N_8600,N_8212);
and U9026 (N_9026,N_8686,N_8435);
xor U9027 (N_9027,N_8743,N_8337);
xnor U9028 (N_9028,N_8708,N_8608);
nand U9029 (N_9029,N_8680,N_8442);
and U9030 (N_9030,N_8693,N_8720);
and U9031 (N_9031,N_8324,N_8493);
and U9032 (N_9032,N_8569,N_8422);
xnor U9033 (N_9033,N_8529,N_8428);
or U9034 (N_9034,N_8175,N_8270);
nand U9035 (N_9035,N_8414,N_8380);
and U9036 (N_9036,N_8404,N_8424);
xnor U9037 (N_9037,N_8747,N_8196);
nor U9038 (N_9038,N_8664,N_8364);
nor U9039 (N_9039,N_8744,N_8447);
nor U9040 (N_9040,N_8710,N_8563);
nand U9041 (N_9041,N_8522,N_8675);
xnor U9042 (N_9042,N_8549,N_8676);
and U9043 (N_9043,N_8248,N_8367);
or U9044 (N_9044,N_8716,N_8163);
nand U9045 (N_9045,N_8169,N_8584);
nor U9046 (N_9046,N_8476,N_8455);
or U9047 (N_9047,N_8312,N_8421);
and U9048 (N_9048,N_8590,N_8207);
and U9049 (N_9049,N_8252,N_8662);
nor U9050 (N_9050,N_8237,N_8423);
and U9051 (N_9051,N_8715,N_8363);
and U9052 (N_9052,N_8247,N_8598);
xnor U9053 (N_9053,N_8617,N_8576);
xnor U9054 (N_9054,N_8534,N_8268);
nor U9055 (N_9055,N_8564,N_8362);
or U9056 (N_9056,N_8323,N_8483);
or U9057 (N_9057,N_8290,N_8235);
or U9058 (N_9058,N_8588,N_8152);
nor U9059 (N_9059,N_8518,N_8279);
xor U9060 (N_9060,N_8490,N_8162);
nand U9061 (N_9061,N_8486,N_8517);
and U9062 (N_9062,N_8289,N_8578);
or U9063 (N_9063,N_8578,N_8642);
nand U9064 (N_9064,N_8699,N_8467);
xor U9065 (N_9065,N_8703,N_8732);
or U9066 (N_9066,N_8398,N_8390);
and U9067 (N_9067,N_8438,N_8717);
and U9068 (N_9068,N_8733,N_8620);
and U9069 (N_9069,N_8189,N_8206);
nand U9070 (N_9070,N_8230,N_8686);
and U9071 (N_9071,N_8707,N_8308);
xnor U9072 (N_9072,N_8594,N_8586);
nand U9073 (N_9073,N_8378,N_8207);
nand U9074 (N_9074,N_8561,N_8465);
and U9075 (N_9075,N_8304,N_8373);
nand U9076 (N_9076,N_8181,N_8312);
and U9077 (N_9077,N_8508,N_8491);
nand U9078 (N_9078,N_8407,N_8306);
or U9079 (N_9079,N_8145,N_8436);
nand U9080 (N_9080,N_8173,N_8606);
xor U9081 (N_9081,N_8409,N_8485);
nand U9082 (N_9082,N_8449,N_8747);
and U9083 (N_9083,N_8160,N_8163);
or U9084 (N_9084,N_8704,N_8686);
nor U9085 (N_9085,N_8586,N_8168);
nor U9086 (N_9086,N_8665,N_8422);
or U9087 (N_9087,N_8452,N_8568);
xor U9088 (N_9088,N_8159,N_8355);
xor U9089 (N_9089,N_8312,N_8557);
and U9090 (N_9090,N_8494,N_8254);
and U9091 (N_9091,N_8462,N_8445);
xor U9092 (N_9092,N_8408,N_8310);
or U9093 (N_9093,N_8137,N_8302);
xor U9094 (N_9094,N_8640,N_8418);
nor U9095 (N_9095,N_8569,N_8566);
xnor U9096 (N_9096,N_8608,N_8300);
or U9097 (N_9097,N_8351,N_8544);
and U9098 (N_9098,N_8657,N_8737);
nor U9099 (N_9099,N_8186,N_8401);
nor U9100 (N_9100,N_8487,N_8400);
and U9101 (N_9101,N_8718,N_8343);
nand U9102 (N_9102,N_8147,N_8179);
xnor U9103 (N_9103,N_8490,N_8463);
xnor U9104 (N_9104,N_8455,N_8553);
xnor U9105 (N_9105,N_8336,N_8144);
xnor U9106 (N_9106,N_8551,N_8700);
and U9107 (N_9107,N_8433,N_8420);
and U9108 (N_9108,N_8282,N_8240);
nor U9109 (N_9109,N_8279,N_8673);
xnor U9110 (N_9110,N_8643,N_8211);
nor U9111 (N_9111,N_8531,N_8738);
nor U9112 (N_9112,N_8540,N_8595);
xor U9113 (N_9113,N_8572,N_8549);
nor U9114 (N_9114,N_8344,N_8127);
or U9115 (N_9115,N_8367,N_8363);
xnor U9116 (N_9116,N_8172,N_8154);
nand U9117 (N_9117,N_8248,N_8207);
xor U9118 (N_9118,N_8284,N_8506);
nor U9119 (N_9119,N_8548,N_8458);
and U9120 (N_9120,N_8581,N_8612);
and U9121 (N_9121,N_8136,N_8482);
nor U9122 (N_9122,N_8514,N_8650);
or U9123 (N_9123,N_8233,N_8731);
xnor U9124 (N_9124,N_8262,N_8435);
nor U9125 (N_9125,N_8330,N_8262);
nand U9126 (N_9126,N_8296,N_8641);
nand U9127 (N_9127,N_8354,N_8513);
xnor U9128 (N_9128,N_8143,N_8542);
nor U9129 (N_9129,N_8174,N_8402);
or U9130 (N_9130,N_8701,N_8146);
nor U9131 (N_9131,N_8685,N_8330);
and U9132 (N_9132,N_8736,N_8217);
nand U9133 (N_9133,N_8476,N_8556);
and U9134 (N_9134,N_8319,N_8131);
nor U9135 (N_9135,N_8428,N_8384);
and U9136 (N_9136,N_8250,N_8235);
xnor U9137 (N_9137,N_8482,N_8452);
nand U9138 (N_9138,N_8281,N_8540);
nand U9139 (N_9139,N_8382,N_8363);
and U9140 (N_9140,N_8146,N_8627);
nor U9141 (N_9141,N_8734,N_8351);
nand U9142 (N_9142,N_8398,N_8357);
xnor U9143 (N_9143,N_8645,N_8339);
and U9144 (N_9144,N_8148,N_8180);
and U9145 (N_9145,N_8653,N_8428);
nand U9146 (N_9146,N_8660,N_8633);
xnor U9147 (N_9147,N_8722,N_8681);
nand U9148 (N_9148,N_8620,N_8628);
xor U9149 (N_9149,N_8547,N_8204);
nand U9150 (N_9150,N_8355,N_8518);
and U9151 (N_9151,N_8712,N_8548);
and U9152 (N_9152,N_8138,N_8161);
nand U9153 (N_9153,N_8506,N_8249);
or U9154 (N_9154,N_8265,N_8360);
and U9155 (N_9155,N_8170,N_8714);
xor U9156 (N_9156,N_8659,N_8419);
nand U9157 (N_9157,N_8632,N_8262);
nand U9158 (N_9158,N_8402,N_8593);
xor U9159 (N_9159,N_8507,N_8486);
and U9160 (N_9160,N_8721,N_8341);
nor U9161 (N_9161,N_8366,N_8658);
xor U9162 (N_9162,N_8349,N_8684);
and U9163 (N_9163,N_8387,N_8199);
or U9164 (N_9164,N_8230,N_8291);
nor U9165 (N_9165,N_8322,N_8288);
and U9166 (N_9166,N_8282,N_8359);
xor U9167 (N_9167,N_8234,N_8329);
xnor U9168 (N_9168,N_8263,N_8250);
nand U9169 (N_9169,N_8419,N_8233);
nand U9170 (N_9170,N_8326,N_8424);
or U9171 (N_9171,N_8299,N_8602);
xor U9172 (N_9172,N_8606,N_8458);
or U9173 (N_9173,N_8416,N_8313);
and U9174 (N_9174,N_8331,N_8192);
nand U9175 (N_9175,N_8241,N_8676);
xnor U9176 (N_9176,N_8221,N_8466);
nand U9177 (N_9177,N_8361,N_8472);
and U9178 (N_9178,N_8533,N_8645);
or U9179 (N_9179,N_8555,N_8134);
nor U9180 (N_9180,N_8599,N_8171);
and U9181 (N_9181,N_8463,N_8368);
nor U9182 (N_9182,N_8247,N_8384);
nand U9183 (N_9183,N_8627,N_8258);
and U9184 (N_9184,N_8636,N_8585);
or U9185 (N_9185,N_8350,N_8383);
nor U9186 (N_9186,N_8282,N_8659);
nand U9187 (N_9187,N_8302,N_8665);
nand U9188 (N_9188,N_8194,N_8594);
xor U9189 (N_9189,N_8133,N_8630);
nand U9190 (N_9190,N_8241,N_8400);
nand U9191 (N_9191,N_8703,N_8731);
or U9192 (N_9192,N_8665,N_8721);
or U9193 (N_9193,N_8311,N_8255);
xnor U9194 (N_9194,N_8450,N_8594);
xnor U9195 (N_9195,N_8665,N_8611);
xor U9196 (N_9196,N_8718,N_8171);
and U9197 (N_9197,N_8617,N_8280);
xor U9198 (N_9198,N_8384,N_8546);
and U9199 (N_9199,N_8457,N_8332);
and U9200 (N_9200,N_8151,N_8278);
and U9201 (N_9201,N_8414,N_8306);
xor U9202 (N_9202,N_8493,N_8606);
or U9203 (N_9203,N_8246,N_8406);
xor U9204 (N_9204,N_8453,N_8257);
xnor U9205 (N_9205,N_8373,N_8324);
or U9206 (N_9206,N_8384,N_8252);
nand U9207 (N_9207,N_8213,N_8426);
xor U9208 (N_9208,N_8363,N_8279);
and U9209 (N_9209,N_8465,N_8266);
xor U9210 (N_9210,N_8737,N_8620);
and U9211 (N_9211,N_8128,N_8749);
nand U9212 (N_9212,N_8363,N_8310);
nor U9213 (N_9213,N_8161,N_8198);
xor U9214 (N_9214,N_8175,N_8441);
xnor U9215 (N_9215,N_8179,N_8682);
nor U9216 (N_9216,N_8377,N_8306);
or U9217 (N_9217,N_8241,N_8478);
and U9218 (N_9218,N_8691,N_8336);
nor U9219 (N_9219,N_8292,N_8320);
or U9220 (N_9220,N_8230,N_8600);
nor U9221 (N_9221,N_8165,N_8705);
nor U9222 (N_9222,N_8130,N_8236);
xnor U9223 (N_9223,N_8539,N_8383);
xnor U9224 (N_9224,N_8514,N_8491);
and U9225 (N_9225,N_8424,N_8510);
nand U9226 (N_9226,N_8721,N_8560);
nor U9227 (N_9227,N_8389,N_8721);
or U9228 (N_9228,N_8473,N_8500);
xor U9229 (N_9229,N_8195,N_8677);
or U9230 (N_9230,N_8185,N_8407);
and U9231 (N_9231,N_8131,N_8327);
nor U9232 (N_9232,N_8139,N_8280);
nand U9233 (N_9233,N_8159,N_8651);
and U9234 (N_9234,N_8331,N_8256);
nor U9235 (N_9235,N_8288,N_8443);
nand U9236 (N_9236,N_8557,N_8512);
or U9237 (N_9237,N_8749,N_8721);
or U9238 (N_9238,N_8488,N_8164);
nor U9239 (N_9239,N_8150,N_8277);
and U9240 (N_9240,N_8400,N_8510);
and U9241 (N_9241,N_8239,N_8611);
xnor U9242 (N_9242,N_8574,N_8618);
and U9243 (N_9243,N_8391,N_8397);
or U9244 (N_9244,N_8540,N_8660);
nor U9245 (N_9245,N_8254,N_8367);
nor U9246 (N_9246,N_8447,N_8642);
xor U9247 (N_9247,N_8540,N_8175);
nor U9248 (N_9248,N_8349,N_8749);
nor U9249 (N_9249,N_8234,N_8316);
nor U9250 (N_9250,N_8636,N_8384);
xnor U9251 (N_9251,N_8524,N_8626);
nor U9252 (N_9252,N_8175,N_8559);
and U9253 (N_9253,N_8566,N_8458);
and U9254 (N_9254,N_8700,N_8430);
nor U9255 (N_9255,N_8591,N_8693);
and U9256 (N_9256,N_8161,N_8322);
or U9257 (N_9257,N_8726,N_8135);
or U9258 (N_9258,N_8579,N_8277);
or U9259 (N_9259,N_8451,N_8471);
nand U9260 (N_9260,N_8165,N_8748);
nor U9261 (N_9261,N_8658,N_8323);
nand U9262 (N_9262,N_8549,N_8405);
nand U9263 (N_9263,N_8567,N_8555);
or U9264 (N_9264,N_8231,N_8511);
nand U9265 (N_9265,N_8349,N_8310);
nand U9266 (N_9266,N_8379,N_8481);
nand U9267 (N_9267,N_8526,N_8713);
or U9268 (N_9268,N_8324,N_8184);
xor U9269 (N_9269,N_8747,N_8315);
nor U9270 (N_9270,N_8510,N_8246);
nand U9271 (N_9271,N_8270,N_8199);
nand U9272 (N_9272,N_8664,N_8208);
nor U9273 (N_9273,N_8733,N_8448);
xnor U9274 (N_9274,N_8301,N_8377);
and U9275 (N_9275,N_8299,N_8201);
nand U9276 (N_9276,N_8293,N_8554);
xnor U9277 (N_9277,N_8428,N_8406);
or U9278 (N_9278,N_8366,N_8460);
nor U9279 (N_9279,N_8232,N_8538);
nor U9280 (N_9280,N_8539,N_8597);
and U9281 (N_9281,N_8377,N_8249);
nor U9282 (N_9282,N_8729,N_8410);
nand U9283 (N_9283,N_8742,N_8129);
or U9284 (N_9284,N_8685,N_8332);
or U9285 (N_9285,N_8358,N_8325);
nand U9286 (N_9286,N_8618,N_8266);
or U9287 (N_9287,N_8445,N_8461);
and U9288 (N_9288,N_8508,N_8445);
nand U9289 (N_9289,N_8529,N_8354);
and U9290 (N_9290,N_8343,N_8706);
xnor U9291 (N_9291,N_8360,N_8459);
or U9292 (N_9292,N_8565,N_8571);
or U9293 (N_9293,N_8622,N_8273);
nand U9294 (N_9294,N_8434,N_8473);
or U9295 (N_9295,N_8137,N_8727);
nand U9296 (N_9296,N_8136,N_8303);
nor U9297 (N_9297,N_8253,N_8690);
nand U9298 (N_9298,N_8381,N_8723);
xor U9299 (N_9299,N_8476,N_8572);
or U9300 (N_9300,N_8535,N_8154);
and U9301 (N_9301,N_8137,N_8149);
and U9302 (N_9302,N_8343,N_8685);
and U9303 (N_9303,N_8518,N_8471);
or U9304 (N_9304,N_8622,N_8490);
and U9305 (N_9305,N_8615,N_8675);
xor U9306 (N_9306,N_8587,N_8265);
nor U9307 (N_9307,N_8379,N_8602);
or U9308 (N_9308,N_8233,N_8562);
nor U9309 (N_9309,N_8593,N_8632);
nor U9310 (N_9310,N_8234,N_8514);
and U9311 (N_9311,N_8724,N_8294);
or U9312 (N_9312,N_8547,N_8157);
and U9313 (N_9313,N_8636,N_8563);
and U9314 (N_9314,N_8335,N_8296);
or U9315 (N_9315,N_8304,N_8138);
xor U9316 (N_9316,N_8582,N_8480);
nand U9317 (N_9317,N_8265,N_8223);
nor U9318 (N_9318,N_8131,N_8602);
xnor U9319 (N_9319,N_8707,N_8244);
or U9320 (N_9320,N_8282,N_8459);
or U9321 (N_9321,N_8683,N_8514);
xor U9322 (N_9322,N_8669,N_8615);
and U9323 (N_9323,N_8667,N_8320);
nand U9324 (N_9324,N_8691,N_8359);
and U9325 (N_9325,N_8468,N_8573);
nand U9326 (N_9326,N_8149,N_8283);
nor U9327 (N_9327,N_8269,N_8597);
nor U9328 (N_9328,N_8506,N_8195);
nor U9329 (N_9329,N_8147,N_8735);
nand U9330 (N_9330,N_8371,N_8217);
xnor U9331 (N_9331,N_8398,N_8737);
or U9332 (N_9332,N_8199,N_8390);
nor U9333 (N_9333,N_8240,N_8574);
nor U9334 (N_9334,N_8603,N_8645);
xnor U9335 (N_9335,N_8137,N_8146);
nand U9336 (N_9336,N_8551,N_8261);
xnor U9337 (N_9337,N_8599,N_8553);
nor U9338 (N_9338,N_8212,N_8485);
and U9339 (N_9339,N_8396,N_8385);
nand U9340 (N_9340,N_8177,N_8303);
nor U9341 (N_9341,N_8385,N_8725);
nand U9342 (N_9342,N_8602,N_8289);
nand U9343 (N_9343,N_8140,N_8244);
xor U9344 (N_9344,N_8196,N_8525);
and U9345 (N_9345,N_8158,N_8741);
nor U9346 (N_9346,N_8455,N_8190);
nor U9347 (N_9347,N_8580,N_8482);
or U9348 (N_9348,N_8338,N_8552);
and U9349 (N_9349,N_8244,N_8648);
and U9350 (N_9350,N_8698,N_8191);
nand U9351 (N_9351,N_8307,N_8141);
nand U9352 (N_9352,N_8434,N_8629);
nand U9353 (N_9353,N_8586,N_8746);
or U9354 (N_9354,N_8520,N_8217);
or U9355 (N_9355,N_8419,N_8559);
nor U9356 (N_9356,N_8630,N_8583);
nor U9357 (N_9357,N_8233,N_8387);
xor U9358 (N_9358,N_8275,N_8600);
and U9359 (N_9359,N_8421,N_8266);
xnor U9360 (N_9360,N_8151,N_8279);
xnor U9361 (N_9361,N_8498,N_8748);
or U9362 (N_9362,N_8487,N_8717);
and U9363 (N_9363,N_8376,N_8633);
nand U9364 (N_9364,N_8262,N_8506);
and U9365 (N_9365,N_8596,N_8376);
or U9366 (N_9366,N_8367,N_8298);
xnor U9367 (N_9367,N_8416,N_8519);
or U9368 (N_9368,N_8705,N_8500);
and U9369 (N_9369,N_8218,N_8195);
nand U9370 (N_9370,N_8709,N_8487);
or U9371 (N_9371,N_8552,N_8176);
nand U9372 (N_9372,N_8731,N_8397);
or U9373 (N_9373,N_8368,N_8286);
nor U9374 (N_9374,N_8181,N_8532);
xnor U9375 (N_9375,N_9255,N_9177);
nand U9376 (N_9376,N_8775,N_9339);
and U9377 (N_9377,N_9211,N_9149);
or U9378 (N_9378,N_9090,N_9155);
nor U9379 (N_9379,N_9374,N_9007);
or U9380 (N_9380,N_9049,N_8780);
or U9381 (N_9381,N_8788,N_9027);
nor U9382 (N_9382,N_8808,N_8774);
nor U9383 (N_9383,N_8932,N_9205);
or U9384 (N_9384,N_8823,N_8786);
and U9385 (N_9385,N_9171,N_9253);
nor U9386 (N_9386,N_9278,N_9256);
nor U9387 (N_9387,N_9033,N_9099);
and U9388 (N_9388,N_8977,N_9113);
nor U9389 (N_9389,N_9103,N_8996);
xor U9390 (N_9390,N_8900,N_9055);
nand U9391 (N_9391,N_8989,N_8763);
nor U9392 (N_9392,N_9137,N_8857);
and U9393 (N_9393,N_9236,N_9292);
nand U9394 (N_9394,N_8965,N_8968);
and U9395 (N_9395,N_9296,N_9015);
nor U9396 (N_9396,N_9119,N_9367);
nor U9397 (N_9397,N_8874,N_9096);
and U9398 (N_9398,N_8807,N_9012);
nor U9399 (N_9399,N_9220,N_9248);
nand U9400 (N_9400,N_9262,N_8952);
nand U9401 (N_9401,N_9228,N_8962);
and U9402 (N_9402,N_9309,N_9330);
nand U9403 (N_9403,N_9305,N_9216);
or U9404 (N_9404,N_9125,N_9023);
nor U9405 (N_9405,N_8751,N_9226);
or U9406 (N_9406,N_9025,N_9131);
and U9407 (N_9407,N_8850,N_8862);
nand U9408 (N_9408,N_9053,N_8908);
or U9409 (N_9409,N_8803,N_9293);
xor U9410 (N_9410,N_8997,N_8809);
xnor U9411 (N_9411,N_9089,N_9298);
xor U9412 (N_9412,N_9288,N_9347);
nand U9413 (N_9413,N_9279,N_9129);
xor U9414 (N_9414,N_8990,N_8776);
or U9415 (N_9415,N_8949,N_8929);
xnor U9416 (N_9416,N_9212,N_9084);
and U9417 (N_9417,N_9344,N_8921);
nand U9418 (N_9418,N_8914,N_8777);
nand U9419 (N_9419,N_8766,N_8873);
or U9420 (N_9420,N_9206,N_9195);
xor U9421 (N_9421,N_9136,N_9366);
or U9422 (N_9422,N_9071,N_9139);
and U9423 (N_9423,N_9218,N_9277);
nand U9424 (N_9424,N_9038,N_8846);
or U9425 (N_9425,N_9289,N_8887);
nand U9426 (N_9426,N_9264,N_8866);
and U9427 (N_9427,N_9043,N_9303);
nor U9428 (N_9428,N_8794,N_9187);
nand U9429 (N_9429,N_9168,N_8833);
and U9430 (N_9430,N_9140,N_8799);
nand U9431 (N_9431,N_9359,N_9350);
and U9432 (N_9432,N_9234,N_9317);
nor U9433 (N_9433,N_8938,N_8993);
nand U9434 (N_9434,N_9276,N_8934);
or U9435 (N_9435,N_8769,N_9146);
xor U9436 (N_9436,N_8843,N_8975);
xnor U9437 (N_9437,N_9108,N_8950);
and U9438 (N_9438,N_9267,N_8883);
and U9439 (N_9439,N_9176,N_9325);
nand U9440 (N_9440,N_9243,N_8859);
xor U9441 (N_9441,N_9313,N_9324);
xor U9442 (N_9442,N_9338,N_9078);
nor U9443 (N_9443,N_9065,N_9247);
xor U9444 (N_9444,N_8773,N_9068);
nor U9445 (N_9445,N_9002,N_8836);
nor U9446 (N_9446,N_8798,N_8813);
or U9447 (N_9447,N_9127,N_8838);
or U9448 (N_9448,N_9196,N_9105);
nand U9449 (N_9449,N_8964,N_9057);
and U9450 (N_9450,N_9286,N_8957);
xor U9451 (N_9451,N_9353,N_9351);
nor U9452 (N_9452,N_9284,N_8853);
nand U9453 (N_9453,N_8827,N_9174);
and U9454 (N_9454,N_8854,N_9118);
nand U9455 (N_9455,N_8924,N_9100);
xnor U9456 (N_9456,N_9230,N_8753);
xnor U9457 (N_9457,N_9148,N_8919);
xor U9458 (N_9458,N_8871,N_9249);
nor U9459 (N_9459,N_8872,N_8868);
xor U9460 (N_9460,N_9362,N_9063);
nand U9461 (N_9461,N_8875,N_9151);
or U9462 (N_9462,N_8917,N_9335);
and U9463 (N_9463,N_9192,N_8999);
or U9464 (N_9464,N_9181,N_9029);
or U9465 (N_9465,N_9275,N_9164);
xnor U9466 (N_9466,N_9101,N_8907);
nand U9467 (N_9467,N_8909,N_9020);
or U9468 (N_9468,N_8876,N_8778);
nand U9469 (N_9469,N_9001,N_9154);
xor U9470 (N_9470,N_8985,N_9165);
nor U9471 (N_9471,N_9021,N_9036);
nand U9472 (N_9472,N_8994,N_8987);
and U9473 (N_9473,N_9287,N_9348);
xor U9474 (N_9474,N_9083,N_9087);
nand U9475 (N_9475,N_9209,N_8764);
and U9476 (N_9476,N_8953,N_9133);
nor U9477 (N_9477,N_8841,N_8955);
and U9478 (N_9478,N_9032,N_8946);
or U9479 (N_9479,N_9183,N_9039);
or U9480 (N_9480,N_9056,N_9024);
and U9481 (N_9481,N_9132,N_9217);
and U9482 (N_9482,N_9144,N_9368);
or U9483 (N_9483,N_9156,N_9184);
or U9484 (N_9484,N_8792,N_8954);
or U9485 (N_9485,N_8933,N_9157);
nand U9486 (N_9486,N_8886,N_8937);
nand U9487 (N_9487,N_8967,N_9357);
nor U9488 (N_9488,N_8811,N_8761);
and U9489 (N_9489,N_8752,N_9016);
or U9490 (N_9490,N_8852,N_9030);
nor U9491 (N_9491,N_9169,N_9308);
nand U9492 (N_9492,N_8963,N_8756);
nor U9493 (N_9493,N_9369,N_9372);
xnor U9494 (N_9494,N_9221,N_8970);
and U9495 (N_9495,N_9019,N_9079);
nor U9496 (N_9496,N_8771,N_9048);
or U9497 (N_9497,N_9214,N_9088);
nand U9498 (N_9498,N_9361,N_8787);
and U9499 (N_9499,N_8842,N_9327);
or U9500 (N_9500,N_9290,N_9210);
xor U9501 (N_9501,N_9259,N_8982);
nand U9502 (N_9502,N_9091,N_8926);
nor U9503 (N_9503,N_9081,N_8762);
xor U9504 (N_9504,N_8884,N_9269);
or U9505 (N_9505,N_8925,N_9035);
or U9506 (N_9506,N_9252,N_9198);
nand U9507 (N_9507,N_9005,N_9258);
nor U9508 (N_9508,N_9110,N_9340);
and U9509 (N_9509,N_8856,N_8782);
and U9510 (N_9510,N_8895,N_9158);
and U9511 (N_9511,N_9336,N_9180);
xnor U9512 (N_9512,N_9354,N_8943);
nor U9513 (N_9513,N_8897,N_9190);
and U9514 (N_9514,N_9143,N_9349);
and U9515 (N_9515,N_8892,N_8837);
or U9516 (N_9516,N_9345,N_8801);
nand U9517 (N_9517,N_8972,N_9297);
xor U9518 (N_9518,N_8861,N_9343);
or U9519 (N_9519,N_9213,N_9251);
and U9520 (N_9520,N_9166,N_9054);
xnor U9521 (N_9521,N_9026,N_8941);
xor U9522 (N_9522,N_9014,N_8911);
xor U9523 (N_9523,N_8991,N_8898);
nor U9524 (N_9524,N_8863,N_9172);
nand U9525 (N_9525,N_9215,N_8793);
nand U9526 (N_9526,N_9283,N_8881);
or U9527 (N_9527,N_8885,N_8758);
or U9528 (N_9528,N_9334,N_9315);
nor U9529 (N_9529,N_9152,N_8961);
and U9530 (N_9530,N_9041,N_8848);
nor U9531 (N_9531,N_9320,N_8855);
nand U9532 (N_9532,N_8849,N_9203);
xnor U9533 (N_9533,N_9145,N_8916);
and U9534 (N_9534,N_9060,N_9082);
xnor U9535 (N_9535,N_8870,N_8928);
xnor U9536 (N_9536,N_9042,N_8992);
nand U9537 (N_9537,N_8800,N_9009);
or U9538 (N_9538,N_9075,N_9322);
xnor U9539 (N_9539,N_8858,N_9207);
or U9540 (N_9540,N_9365,N_8879);
nor U9541 (N_9541,N_9161,N_8750);
or U9542 (N_9542,N_8789,N_8810);
or U9543 (N_9543,N_9363,N_8893);
or U9544 (N_9544,N_8821,N_8903);
xor U9545 (N_9545,N_8828,N_8783);
xnor U9546 (N_9546,N_8944,N_9202);
xor U9547 (N_9547,N_9044,N_9333);
or U9548 (N_9548,N_9018,N_9273);
nand U9549 (N_9549,N_9291,N_9186);
and U9550 (N_9550,N_8817,N_8832);
or U9551 (N_9551,N_9245,N_8816);
nor U9552 (N_9552,N_8978,N_9128);
xnor U9553 (N_9553,N_8939,N_8940);
nor U9554 (N_9554,N_9329,N_8819);
nand U9555 (N_9555,N_9229,N_8820);
or U9556 (N_9556,N_9170,N_9022);
and U9557 (N_9557,N_8865,N_9310);
or U9558 (N_9558,N_9240,N_8971);
nand U9559 (N_9559,N_8945,N_9233);
nand U9560 (N_9560,N_8878,N_9059);
or U9561 (N_9561,N_9270,N_9073);
and U9562 (N_9562,N_8935,N_8896);
nor U9563 (N_9563,N_9062,N_9077);
xnor U9564 (N_9564,N_9097,N_9070);
nor U9565 (N_9565,N_9052,N_9311);
and U9566 (N_9566,N_8923,N_9342);
nand U9567 (N_9567,N_9178,N_8797);
and U9568 (N_9568,N_8905,N_9112);
nor U9569 (N_9569,N_9163,N_9098);
and U9570 (N_9570,N_9093,N_9352);
or U9571 (N_9571,N_9318,N_9111);
or U9572 (N_9572,N_9130,N_8845);
nor U9573 (N_9573,N_8806,N_8980);
or U9574 (N_9574,N_9355,N_8770);
xnor U9575 (N_9575,N_9314,N_8976);
nor U9576 (N_9576,N_9280,N_8768);
nand U9577 (N_9577,N_9373,N_9199);
nand U9578 (N_9578,N_9179,N_9326);
nor U9579 (N_9579,N_9306,N_8966);
or U9580 (N_9580,N_8785,N_9069);
nand U9581 (N_9581,N_9147,N_8959);
xor U9582 (N_9582,N_8796,N_8894);
nand U9583 (N_9583,N_9197,N_9235);
and U9584 (N_9584,N_8784,N_9159);
nor U9585 (N_9585,N_9225,N_8890);
nand U9586 (N_9586,N_9200,N_8981);
or U9587 (N_9587,N_8830,N_8882);
xnor U9588 (N_9588,N_9321,N_9358);
and U9589 (N_9589,N_9061,N_9246);
nor U9590 (N_9590,N_9086,N_9281);
and U9591 (N_9591,N_8973,N_9028);
xnor U9592 (N_9592,N_9301,N_8984);
or U9593 (N_9593,N_8825,N_9201);
and U9594 (N_9594,N_9360,N_9328);
nor U9595 (N_9595,N_9319,N_8767);
nor U9596 (N_9596,N_8927,N_9141);
and U9597 (N_9597,N_8891,N_8983);
xnor U9598 (N_9598,N_9064,N_8974);
or U9599 (N_9599,N_9004,N_8986);
nor U9600 (N_9600,N_9307,N_8931);
and U9601 (N_9601,N_9121,N_9185);
or U9602 (N_9602,N_8835,N_9371);
nor U9603 (N_9603,N_8851,N_8951);
nand U9604 (N_9604,N_8826,N_8888);
and U9605 (N_9605,N_9045,N_9266);
nand U9606 (N_9606,N_9223,N_9260);
nor U9607 (N_9607,N_8791,N_8757);
xnor U9608 (N_9608,N_8805,N_9006);
nand U9609 (N_9609,N_9150,N_8912);
or U9610 (N_9610,N_9116,N_9067);
and U9611 (N_9611,N_9117,N_9126);
or U9612 (N_9612,N_9316,N_8979);
nor U9613 (N_9613,N_8901,N_9302);
nor U9614 (N_9614,N_9191,N_8899);
nand U9615 (N_9615,N_9104,N_9194);
nor U9616 (N_9616,N_9250,N_9346);
xnor U9617 (N_9617,N_8824,N_9135);
or U9618 (N_9618,N_8904,N_8867);
or U9619 (N_9619,N_8902,N_9051);
and U9620 (N_9620,N_9046,N_9323);
nand U9621 (N_9621,N_8814,N_8918);
or U9622 (N_9622,N_9162,N_9254);
or U9623 (N_9623,N_9175,N_8880);
nand U9624 (N_9624,N_9265,N_9094);
and U9625 (N_9625,N_9189,N_8995);
and U9626 (N_9626,N_9072,N_9300);
and U9627 (N_9627,N_9034,N_8812);
nand U9628 (N_9628,N_8834,N_8958);
and U9629 (N_9629,N_9173,N_9010);
and U9630 (N_9630,N_9241,N_9050);
nand U9631 (N_9631,N_8831,N_9124);
xor U9632 (N_9632,N_8818,N_9120);
xor U9633 (N_9633,N_9232,N_8942);
and U9634 (N_9634,N_9058,N_9364);
xnor U9635 (N_9635,N_8781,N_9341);
xnor U9636 (N_9636,N_9263,N_8998);
xnor U9637 (N_9637,N_9080,N_8802);
and U9638 (N_9638,N_8765,N_8956);
or U9639 (N_9639,N_9193,N_8815);
nor U9640 (N_9640,N_9295,N_8906);
nor U9641 (N_9641,N_9011,N_9047);
nand U9642 (N_9642,N_8847,N_9031);
and U9643 (N_9643,N_9224,N_8947);
or U9644 (N_9644,N_9003,N_9182);
xor U9645 (N_9645,N_9160,N_8844);
xnor U9646 (N_9646,N_8795,N_9092);
and U9647 (N_9647,N_9037,N_8829);
xnor U9648 (N_9648,N_8864,N_9008);
nor U9649 (N_9649,N_8930,N_9123);
and U9650 (N_9650,N_8860,N_8869);
nor U9651 (N_9651,N_9017,N_8913);
nor U9652 (N_9652,N_8910,N_9331);
and U9653 (N_9653,N_9257,N_9134);
and U9654 (N_9654,N_9013,N_8760);
nor U9655 (N_9655,N_9095,N_9102);
and U9656 (N_9656,N_9337,N_8969);
and U9657 (N_9657,N_9294,N_9268);
or U9658 (N_9658,N_9107,N_8922);
and U9659 (N_9659,N_9271,N_9237);
nor U9660 (N_9660,N_9142,N_9312);
and U9661 (N_9661,N_8822,N_9261);
nor U9662 (N_9662,N_9285,N_9085);
nand U9663 (N_9663,N_9122,N_9282);
xor U9664 (N_9664,N_8915,N_9356);
or U9665 (N_9665,N_8755,N_9167);
nand U9666 (N_9666,N_9138,N_8759);
nor U9667 (N_9667,N_9074,N_9106);
xnor U9668 (N_9668,N_9114,N_8804);
nor U9669 (N_9669,N_9238,N_9040);
or U9670 (N_9670,N_8948,N_9332);
and U9671 (N_9671,N_9219,N_8960);
or U9672 (N_9672,N_9370,N_8772);
and U9673 (N_9673,N_9231,N_8779);
nor U9674 (N_9674,N_9239,N_9076);
and U9675 (N_9675,N_9272,N_8790);
xor U9676 (N_9676,N_9109,N_9227);
nor U9677 (N_9677,N_8754,N_8840);
nand U9678 (N_9678,N_9208,N_9000);
nor U9679 (N_9679,N_9066,N_9274);
and U9680 (N_9680,N_8839,N_9115);
xor U9681 (N_9681,N_8920,N_9153);
nor U9682 (N_9682,N_8877,N_9242);
nor U9683 (N_9683,N_9222,N_9304);
nand U9684 (N_9684,N_8889,N_8988);
nor U9685 (N_9685,N_9244,N_9204);
or U9686 (N_9686,N_9188,N_9299);
xnor U9687 (N_9687,N_8936,N_8872);
nor U9688 (N_9688,N_8956,N_9255);
nor U9689 (N_9689,N_9287,N_9009);
nor U9690 (N_9690,N_8882,N_9122);
and U9691 (N_9691,N_8924,N_9200);
nor U9692 (N_9692,N_8859,N_9158);
or U9693 (N_9693,N_8765,N_9193);
or U9694 (N_9694,N_8852,N_9034);
nand U9695 (N_9695,N_8816,N_9163);
xnor U9696 (N_9696,N_9362,N_9223);
or U9697 (N_9697,N_9262,N_8752);
nand U9698 (N_9698,N_8917,N_8887);
nand U9699 (N_9699,N_8811,N_9233);
nor U9700 (N_9700,N_9202,N_9048);
or U9701 (N_9701,N_8993,N_8815);
nor U9702 (N_9702,N_9166,N_8775);
xor U9703 (N_9703,N_9016,N_9268);
or U9704 (N_9704,N_9338,N_8969);
nor U9705 (N_9705,N_9235,N_9246);
and U9706 (N_9706,N_8783,N_9014);
nand U9707 (N_9707,N_9063,N_9316);
xnor U9708 (N_9708,N_8815,N_9314);
or U9709 (N_9709,N_9312,N_9072);
nand U9710 (N_9710,N_8770,N_9333);
xor U9711 (N_9711,N_8940,N_9373);
and U9712 (N_9712,N_8984,N_9224);
or U9713 (N_9713,N_9165,N_8972);
or U9714 (N_9714,N_8992,N_9157);
xnor U9715 (N_9715,N_8840,N_9371);
and U9716 (N_9716,N_8938,N_8914);
and U9717 (N_9717,N_9053,N_9222);
xor U9718 (N_9718,N_8851,N_9214);
or U9719 (N_9719,N_9004,N_9347);
nand U9720 (N_9720,N_8814,N_8902);
xor U9721 (N_9721,N_8951,N_8927);
nor U9722 (N_9722,N_8793,N_9224);
xnor U9723 (N_9723,N_9160,N_9172);
or U9724 (N_9724,N_8767,N_9230);
nand U9725 (N_9725,N_9024,N_9369);
and U9726 (N_9726,N_9178,N_9151);
or U9727 (N_9727,N_9141,N_8844);
nor U9728 (N_9728,N_9341,N_8864);
or U9729 (N_9729,N_8863,N_8840);
xnor U9730 (N_9730,N_8783,N_9335);
or U9731 (N_9731,N_8996,N_9224);
or U9732 (N_9732,N_8957,N_9347);
nor U9733 (N_9733,N_8890,N_9003);
nand U9734 (N_9734,N_9184,N_8966);
xor U9735 (N_9735,N_9079,N_9358);
and U9736 (N_9736,N_9155,N_9232);
nand U9737 (N_9737,N_8859,N_8880);
nor U9738 (N_9738,N_8958,N_8760);
xor U9739 (N_9739,N_9186,N_8800);
nand U9740 (N_9740,N_8818,N_8881);
xnor U9741 (N_9741,N_9220,N_9333);
xor U9742 (N_9742,N_9308,N_9044);
or U9743 (N_9743,N_9210,N_8784);
xnor U9744 (N_9744,N_8860,N_9001);
nand U9745 (N_9745,N_9203,N_9224);
nand U9746 (N_9746,N_8768,N_8945);
nand U9747 (N_9747,N_8829,N_8853);
nor U9748 (N_9748,N_9269,N_8905);
nand U9749 (N_9749,N_8935,N_9220);
nand U9750 (N_9750,N_9362,N_8821);
nand U9751 (N_9751,N_9045,N_8845);
nor U9752 (N_9752,N_9000,N_8766);
or U9753 (N_9753,N_9330,N_8867);
xor U9754 (N_9754,N_9058,N_9147);
nor U9755 (N_9755,N_8940,N_8929);
and U9756 (N_9756,N_9190,N_9030);
xnor U9757 (N_9757,N_8849,N_8929);
and U9758 (N_9758,N_9087,N_9243);
and U9759 (N_9759,N_8925,N_9295);
nor U9760 (N_9760,N_8806,N_9051);
nor U9761 (N_9761,N_9053,N_8846);
or U9762 (N_9762,N_8976,N_9096);
or U9763 (N_9763,N_8811,N_9173);
and U9764 (N_9764,N_9365,N_8812);
nand U9765 (N_9765,N_8923,N_9184);
or U9766 (N_9766,N_9057,N_9180);
nor U9767 (N_9767,N_9233,N_8891);
nor U9768 (N_9768,N_8805,N_9029);
nand U9769 (N_9769,N_8998,N_9325);
and U9770 (N_9770,N_9003,N_9297);
nand U9771 (N_9771,N_8971,N_9294);
nor U9772 (N_9772,N_8898,N_9207);
nand U9773 (N_9773,N_9229,N_9258);
nand U9774 (N_9774,N_9300,N_9080);
nand U9775 (N_9775,N_8891,N_9046);
or U9776 (N_9776,N_8850,N_9300);
and U9777 (N_9777,N_9132,N_8839);
or U9778 (N_9778,N_8765,N_9369);
xor U9779 (N_9779,N_8998,N_9372);
and U9780 (N_9780,N_9367,N_9253);
nand U9781 (N_9781,N_8876,N_9063);
nand U9782 (N_9782,N_8971,N_9119);
and U9783 (N_9783,N_8760,N_8916);
nor U9784 (N_9784,N_8824,N_8961);
nand U9785 (N_9785,N_9182,N_9248);
or U9786 (N_9786,N_9328,N_9226);
or U9787 (N_9787,N_9035,N_9230);
nand U9788 (N_9788,N_8838,N_8980);
nor U9789 (N_9789,N_9068,N_8793);
xnor U9790 (N_9790,N_8928,N_9126);
or U9791 (N_9791,N_9272,N_8781);
xor U9792 (N_9792,N_9352,N_8859);
or U9793 (N_9793,N_9211,N_9340);
or U9794 (N_9794,N_9336,N_9333);
nand U9795 (N_9795,N_9361,N_8891);
and U9796 (N_9796,N_9214,N_8792);
and U9797 (N_9797,N_8804,N_8755);
nor U9798 (N_9798,N_8973,N_9164);
nor U9799 (N_9799,N_9335,N_8761);
nor U9800 (N_9800,N_9052,N_8819);
nand U9801 (N_9801,N_8826,N_8753);
nand U9802 (N_9802,N_8804,N_9367);
or U9803 (N_9803,N_8880,N_9194);
xor U9804 (N_9804,N_9149,N_9355);
or U9805 (N_9805,N_9020,N_8919);
and U9806 (N_9806,N_9123,N_8845);
xor U9807 (N_9807,N_8987,N_9212);
nor U9808 (N_9808,N_9212,N_9056);
nor U9809 (N_9809,N_9360,N_9195);
xnor U9810 (N_9810,N_8995,N_8880);
nand U9811 (N_9811,N_9076,N_8949);
xor U9812 (N_9812,N_9300,N_8841);
nor U9813 (N_9813,N_8753,N_8861);
or U9814 (N_9814,N_9261,N_9159);
xor U9815 (N_9815,N_8899,N_8818);
xnor U9816 (N_9816,N_9214,N_9322);
and U9817 (N_9817,N_9356,N_9023);
or U9818 (N_9818,N_9147,N_8800);
nor U9819 (N_9819,N_8871,N_9266);
nand U9820 (N_9820,N_8783,N_8924);
or U9821 (N_9821,N_8834,N_8937);
and U9822 (N_9822,N_8800,N_9096);
nor U9823 (N_9823,N_9320,N_9135);
nand U9824 (N_9824,N_9255,N_9226);
xnor U9825 (N_9825,N_9030,N_9047);
and U9826 (N_9826,N_9247,N_8773);
and U9827 (N_9827,N_8793,N_9210);
nand U9828 (N_9828,N_9047,N_9291);
and U9829 (N_9829,N_9036,N_8751);
xnor U9830 (N_9830,N_9066,N_9008);
xor U9831 (N_9831,N_9159,N_9265);
or U9832 (N_9832,N_9298,N_8991);
nor U9833 (N_9833,N_9318,N_8778);
nor U9834 (N_9834,N_8846,N_9082);
or U9835 (N_9835,N_8901,N_8831);
or U9836 (N_9836,N_8906,N_9271);
nor U9837 (N_9837,N_9125,N_8873);
xor U9838 (N_9838,N_8956,N_9322);
nand U9839 (N_9839,N_9288,N_9301);
or U9840 (N_9840,N_9215,N_9117);
xnor U9841 (N_9841,N_9168,N_9053);
and U9842 (N_9842,N_8918,N_9118);
nor U9843 (N_9843,N_8871,N_9160);
nand U9844 (N_9844,N_9353,N_9361);
nand U9845 (N_9845,N_9310,N_8992);
nor U9846 (N_9846,N_8951,N_9009);
nand U9847 (N_9847,N_9368,N_9347);
or U9848 (N_9848,N_9153,N_9130);
xor U9849 (N_9849,N_9060,N_9085);
xor U9850 (N_9850,N_9106,N_8779);
or U9851 (N_9851,N_9001,N_9200);
or U9852 (N_9852,N_8918,N_9299);
and U9853 (N_9853,N_8780,N_8992);
or U9854 (N_9854,N_9163,N_9037);
nor U9855 (N_9855,N_9042,N_9000);
nand U9856 (N_9856,N_9003,N_8856);
and U9857 (N_9857,N_9028,N_9184);
nor U9858 (N_9858,N_8766,N_9075);
nand U9859 (N_9859,N_8942,N_8968);
nor U9860 (N_9860,N_8848,N_9178);
nand U9861 (N_9861,N_8831,N_9148);
and U9862 (N_9862,N_9368,N_9095);
nand U9863 (N_9863,N_9088,N_8902);
nor U9864 (N_9864,N_9348,N_9000);
nand U9865 (N_9865,N_8982,N_8926);
or U9866 (N_9866,N_9126,N_9234);
or U9867 (N_9867,N_9336,N_9030);
and U9868 (N_9868,N_8776,N_9255);
or U9869 (N_9869,N_8806,N_8994);
nor U9870 (N_9870,N_8842,N_9323);
nand U9871 (N_9871,N_9226,N_9238);
and U9872 (N_9872,N_8818,N_9224);
nand U9873 (N_9873,N_9056,N_9224);
xor U9874 (N_9874,N_8849,N_9020);
nand U9875 (N_9875,N_9116,N_9261);
xor U9876 (N_9876,N_8911,N_9314);
and U9877 (N_9877,N_8973,N_9229);
nand U9878 (N_9878,N_8898,N_8974);
nor U9879 (N_9879,N_9154,N_8937);
nor U9880 (N_9880,N_9274,N_8963);
nor U9881 (N_9881,N_9164,N_8911);
or U9882 (N_9882,N_9012,N_8873);
nor U9883 (N_9883,N_9175,N_9314);
nor U9884 (N_9884,N_9234,N_8945);
xor U9885 (N_9885,N_8760,N_9253);
or U9886 (N_9886,N_9368,N_9342);
or U9887 (N_9887,N_9235,N_9093);
nor U9888 (N_9888,N_8843,N_9160);
nor U9889 (N_9889,N_9230,N_9353);
nor U9890 (N_9890,N_9159,N_9319);
and U9891 (N_9891,N_9111,N_8803);
nand U9892 (N_9892,N_8804,N_8853);
nand U9893 (N_9893,N_9024,N_9222);
or U9894 (N_9894,N_8884,N_8933);
xor U9895 (N_9895,N_9103,N_9069);
or U9896 (N_9896,N_8913,N_9156);
nand U9897 (N_9897,N_9318,N_9369);
nor U9898 (N_9898,N_8822,N_9228);
nand U9899 (N_9899,N_9278,N_9312);
nand U9900 (N_9900,N_8829,N_9202);
or U9901 (N_9901,N_8989,N_8924);
or U9902 (N_9902,N_9157,N_9247);
or U9903 (N_9903,N_9326,N_9268);
and U9904 (N_9904,N_9204,N_9346);
xor U9905 (N_9905,N_9338,N_9320);
and U9906 (N_9906,N_9164,N_9154);
nor U9907 (N_9907,N_8798,N_9288);
or U9908 (N_9908,N_9128,N_8862);
xnor U9909 (N_9909,N_9318,N_9133);
or U9910 (N_9910,N_9254,N_9248);
nand U9911 (N_9911,N_9150,N_8992);
xnor U9912 (N_9912,N_8779,N_9304);
and U9913 (N_9913,N_8899,N_9167);
or U9914 (N_9914,N_8829,N_8851);
nor U9915 (N_9915,N_9277,N_9088);
and U9916 (N_9916,N_9111,N_9303);
nand U9917 (N_9917,N_8957,N_9322);
nor U9918 (N_9918,N_9369,N_9085);
nand U9919 (N_9919,N_9339,N_9151);
nand U9920 (N_9920,N_8924,N_9106);
nand U9921 (N_9921,N_8789,N_9370);
or U9922 (N_9922,N_9234,N_9131);
or U9923 (N_9923,N_9029,N_8762);
and U9924 (N_9924,N_9058,N_8875);
and U9925 (N_9925,N_9152,N_8839);
nand U9926 (N_9926,N_9074,N_8791);
nand U9927 (N_9927,N_9316,N_8901);
nor U9928 (N_9928,N_9009,N_9023);
nor U9929 (N_9929,N_9246,N_9202);
xor U9930 (N_9930,N_9052,N_9069);
nand U9931 (N_9931,N_8802,N_9099);
nand U9932 (N_9932,N_9034,N_9164);
or U9933 (N_9933,N_8855,N_9105);
nand U9934 (N_9934,N_8761,N_9156);
xnor U9935 (N_9935,N_9320,N_8945);
xnor U9936 (N_9936,N_8796,N_8942);
nor U9937 (N_9937,N_9183,N_9116);
and U9938 (N_9938,N_9064,N_8967);
and U9939 (N_9939,N_9313,N_9065);
xnor U9940 (N_9940,N_9304,N_9276);
or U9941 (N_9941,N_9024,N_9110);
nand U9942 (N_9942,N_9289,N_9007);
nand U9943 (N_9943,N_9355,N_9322);
nor U9944 (N_9944,N_9011,N_9126);
nor U9945 (N_9945,N_8757,N_9070);
or U9946 (N_9946,N_8835,N_9257);
nand U9947 (N_9947,N_9060,N_8994);
or U9948 (N_9948,N_9090,N_9133);
nand U9949 (N_9949,N_9198,N_9184);
and U9950 (N_9950,N_8775,N_9357);
nand U9951 (N_9951,N_9335,N_8874);
or U9952 (N_9952,N_9325,N_9324);
nor U9953 (N_9953,N_8930,N_9275);
nand U9954 (N_9954,N_8942,N_9071);
xor U9955 (N_9955,N_9348,N_9088);
or U9956 (N_9956,N_8770,N_9064);
or U9957 (N_9957,N_9095,N_9338);
xor U9958 (N_9958,N_9131,N_8993);
nor U9959 (N_9959,N_9020,N_8841);
and U9960 (N_9960,N_9105,N_8772);
nor U9961 (N_9961,N_8966,N_9049);
and U9962 (N_9962,N_8964,N_8762);
and U9963 (N_9963,N_9039,N_9365);
nor U9964 (N_9964,N_8763,N_9357);
and U9965 (N_9965,N_9004,N_8996);
and U9966 (N_9966,N_9256,N_8782);
and U9967 (N_9967,N_9249,N_8780);
nor U9968 (N_9968,N_9098,N_9286);
and U9969 (N_9969,N_9230,N_8852);
or U9970 (N_9970,N_8947,N_9327);
nand U9971 (N_9971,N_9128,N_9247);
nand U9972 (N_9972,N_9059,N_8906);
nand U9973 (N_9973,N_8956,N_8943);
nand U9974 (N_9974,N_8761,N_9081);
or U9975 (N_9975,N_9165,N_8871);
or U9976 (N_9976,N_9049,N_8789);
or U9977 (N_9977,N_8904,N_9046);
nand U9978 (N_9978,N_9059,N_9034);
and U9979 (N_9979,N_9266,N_9215);
nor U9980 (N_9980,N_8942,N_8905);
or U9981 (N_9981,N_9297,N_9051);
xor U9982 (N_9982,N_9174,N_8991);
xnor U9983 (N_9983,N_8812,N_9173);
xnor U9984 (N_9984,N_8834,N_9231);
or U9985 (N_9985,N_9244,N_9336);
or U9986 (N_9986,N_8809,N_8778);
xnor U9987 (N_9987,N_8798,N_8820);
or U9988 (N_9988,N_9280,N_9251);
nor U9989 (N_9989,N_8949,N_9163);
or U9990 (N_9990,N_9007,N_9136);
and U9991 (N_9991,N_8899,N_9227);
nor U9992 (N_9992,N_9016,N_9290);
nor U9993 (N_9993,N_9304,N_9005);
nor U9994 (N_9994,N_8934,N_9320);
xnor U9995 (N_9995,N_9347,N_9033);
or U9996 (N_9996,N_9142,N_9297);
nor U9997 (N_9997,N_8890,N_9220);
nand U9998 (N_9998,N_9018,N_8983);
nor U9999 (N_9999,N_8863,N_8926);
xnor U10000 (N_10000,N_9971,N_9675);
or U10001 (N_10001,N_9855,N_9583);
nand U10002 (N_10002,N_9790,N_9611);
xor U10003 (N_10003,N_9875,N_9740);
or U10004 (N_10004,N_9757,N_9990);
nor U10005 (N_10005,N_9625,N_9500);
xor U10006 (N_10006,N_9390,N_9963);
xor U10007 (N_10007,N_9932,N_9408);
or U10008 (N_10008,N_9524,N_9737);
xnor U10009 (N_10009,N_9923,N_9848);
nor U10010 (N_10010,N_9989,N_9957);
or U10011 (N_10011,N_9938,N_9707);
xor U10012 (N_10012,N_9872,N_9378);
or U10013 (N_10013,N_9942,N_9433);
nor U10014 (N_10014,N_9947,N_9847);
and U10015 (N_10015,N_9561,N_9973);
nor U10016 (N_10016,N_9577,N_9443);
or U10017 (N_10017,N_9764,N_9775);
xnor U10018 (N_10018,N_9385,N_9685);
and U10019 (N_10019,N_9455,N_9566);
xor U10020 (N_10020,N_9567,N_9656);
nor U10021 (N_10021,N_9734,N_9442);
and U10022 (N_10022,N_9575,N_9763);
and U10023 (N_10023,N_9826,N_9642);
xnor U10024 (N_10024,N_9890,N_9979);
nor U10025 (N_10025,N_9594,N_9823);
xnor U10026 (N_10026,N_9440,N_9687);
nand U10027 (N_10027,N_9520,N_9405);
nand U10028 (N_10028,N_9754,N_9411);
nor U10029 (N_10029,N_9840,N_9976);
nand U10030 (N_10030,N_9878,N_9821);
and U10031 (N_10031,N_9673,N_9589);
nand U10032 (N_10032,N_9515,N_9811);
or U10033 (N_10033,N_9869,N_9670);
nand U10034 (N_10034,N_9743,N_9574);
nand U10035 (N_10035,N_9531,N_9784);
or U10036 (N_10036,N_9972,N_9491);
or U10037 (N_10037,N_9857,N_9404);
nor U10038 (N_10038,N_9450,N_9424);
nor U10039 (N_10039,N_9783,N_9586);
nand U10040 (N_10040,N_9560,N_9530);
nor U10041 (N_10041,N_9839,N_9709);
nor U10042 (N_10042,N_9981,N_9744);
and U10043 (N_10043,N_9850,N_9987);
and U10044 (N_10044,N_9765,N_9624);
nor U10045 (N_10045,N_9471,N_9711);
xor U10046 (N_10046,N_9845,N_9527);
xor U10047 (N_10047,N_9650,N_9836);
nor U10048 (N_10048,N_9633,N_9526);
nor U10049 (N_10049,N_9948,N_9389);
and U10050 (N_10050,N_9517,N_9806);
and U10051 (N_10051,N_9539,N_9638);
and U10052 (N_10052,N_9729,N_9851);
and U10053 (N_10053,N_9809,N_9564);
xnor U10054 (N_10054,N_9508,N_9608);
xor U10055 (N_10055,N_9759,N_9829);
or U10056 (N_10056,N_9718,N_9620);
nand U10057 (N_10057,N_9710,N_9944);
or U10058 (N_10058,N_9464,N_9580);
and U10059 (N_10059,N_9984,N_9745);
and U10060 (N_10060,N_9644,N_9476);
xor U10061 (N_10061,N_9936,N_9735);
or U10062 (N_10062,N_9792,N_9406);
nand U10063 (N_10063,N_9495,N_9590);
nand U10064 (N_10064,N_9645,N_9513);
or U10065 (N_10065,N_9488,N_9447);
xor U10066 (N_10066,N_9769,N_9696);
nand U10067 (N_10067,N_9893,N_9615);
or U10068 (N_10068,N_9982,N_9804);
xor U10069 (N_10069,N_9714,N_9381);
nand U10070 (N_10070,N_9983,N_9396);
nand U10071 (N_10071,N_9647,N_9886);
or U10072 (N_10072,N_9756,N_9668);
nand U10073 (N_10073,N_9658,N_9761);
and U10074 (N_10074,N_9665,N_9475);
or U10075 (N_10075,N_9572,N_9771);
xor U10076 (N_10076,N_9410,N_9593);
xnor U10077 (N_10077,N_9607,N_9723);
nor U10078 (N_10078,N_9628,N_9437);
or U10079 (N_10079,N_9777,N_9767);
or U10080 (N_10080,N_9430,N_9487);
xnor U10081 (N_10081,N_9698,N_9810);
nor U10082 (N_10082,N_9486,N_9701);
and U10083 (N_10083,N_9964,N_9807);
nand U10084 (N_10084,N_9525,N_9591);
and U10085 (N_10085,N_9399,N_9879);
and U10086 (N_10086,N_9678,N_9796);
xnor U10087 (N_10087,N_9930,N_9721);
nand U10088 (N_10088,N_9789,N_9425);
or U10089 (N_10089,N_9570,N_9417);
and U10090 (N_10090,N_9444,N_9968);
or U10091 (N_10091,N_9470,N_9835);
nand U10092 (N_10092,N_9724,N_9421);
nor U10093 (N_10093,N_9733,N_9728);
or U10094 (N_10094,N_9479,N_9797);
nor U10095 (N_10095,N_9774,N_9720);
and U10096 (N_10096,N_9474,N_9603);
nor U10097 (N_10097,N_9816,N_9629);
or U10098 (N_10098,N_9993,N_9705);
xnor U10099 (N_10099,N_9866,N_9694);
nor U10100 (N_10100,N_9492,N_9716);
xnor U10101 (N_10101,N_9379,N_9827);
and U10102 (N_10102,N_9817,N_9686);
or U10103 (N_10103,N_9802,N_9945);
and U10104 (N_10104,N_9906,N_9894);
nand U10105 (N_10105,N_9951,N_9913);
nand U10106 (N_10106,N_9920,N_9387);
or U10107 (N_10107,N_9898,N_9482);
and U10108 (N_10108,N_9785,N_9897);
nor U10109 (N_10109,N_9534,N_9940);
or U10110 (N_10110,N_9565,N_9929);
and U10111 (N_10111,N_9553,N_9375);
nor U10112 (N_10112,N_9556,N_9978);
nand U10113 (N_10113,N_9516,N_9618);
xor U10114 (N_10114,N_9787,N_9856);
nand U10115 (N_10115,N_9991,N_9895);
nand U10116 (N_10116,N_9900,N_9616);
nand U10117 (N_10117,N_9742,N_9518);
xnor U10118 (N_10118,N_9697,N_9880);
nand U10119 (N_10119,N_9545,N_9926);
and U10120 (N_10120,N_9581,N_9794);
nand U10121 (N_10121,N_9786,N_9782);
xnor U10122 (N_10122,N_9521,N_9960);
nand U10123 (N_10123,N_9676,N_9966);
or U10124 (N_10124,N_9388,N_9382);
nor U10125 (N_10125,N_9852,N_9457);
and U10126 (N_10126,N_9919,N_9507);
and U10127 (N_10127,N_9666,N_9392);
and U10128 (N_10128,N_9631,N_9477);
xor U10129 (N_10129,N_9671,N_9576);
and U10130 (N_10130,N_9397,N_9755);
nand U10131 (N_10131,N_9415,N_9768);
nor U10132 (N_10132,N_9465,N_9533);
and U10133 (N_10133,N_9717,N_9496);
nor U10134 (N_10134,N_9512,N_9610);
xor U10135 (N_10135,N_9652,N_9837);
and U10136 (N_10136,N_9509,N_9612);
or U10137 (N_10137,N_9695,N_9925);
or U10138 (N_10138,N_9414,N_9883);
or U10139 (N_10139,N_9677,N_9497);
nor U10140 (N_10140,N_9587,N_9458);
nand U10141 (N_10141,N_9597,N_9498);
nor U10142 (N_10142,N_9478,N_9937);
nand U10143 (N_10143,N_9598,N_9461);
nand U10144 (N_10144,N_9877,N_9861);
or U10145 (N_10145,N_9600,N_9849);
or U10146 (N_10146,N_9803,N_9649);
or U10147 (N_10147,N_9599,N_9452);
nand U10148 (N_10148,N_9451,N_9941);
and U10149 (N_10149,N_9651,N_9967);
and U10150 (N_10150,N_9918,N_9928);
or U10151 (N_10151,N_9641,N_9445);
xnor U10152 (N_10152,N_9502,N_9888);
and U10153 (N_10153,N_9772,N_9820);
xnor U10154 (N_10154,N_9506,N_9870);
nor U10155 (N_10155,N_9791,N_9899);
xnor U10156 (N_10156,N_9722,N_9884);
nand U10157 (N_10157,N_9688,N_9532);
nand U10158 (N_10158,N_9431,N_9760);
nand U10159 (N_10159,N_9965,N_9632);
nand U10160 (N_10160,N_9674,N_9682);
and U10161 (N_10161,N_9758,N_9838);
nand U10162 (N_10162,N_9619,N_9874);
nor U10163 (N_10163,N_9604,N_9501);
or U10164 (N_10164,N_9902,N_9778);
nor U10165 (N_10165,N_9505,N_9690);
and U10166 (N_10166,N_9739,N_9639);
and U10167 (N_10167,N_9751,N_9995);
xnor U10168 (N_10168,N_9814,N_9562);
nand U10169 (N_10169,N_9749,N_9988);
nand U10170 (N_10170,N_9766,N_9727);
or U10171 (N_10171,N_9958,N_9536);
and U10172 (N_10172,N_9626,N_9891);
nor U10173 (N_10173,N_9860,N_9640);
and U10174 (N_10174,N_9681,N_9833);
xor U10175 (N_10175,N_9726,N_9691);
and U10176 (N_10176,N_9595,N_9912);
nand U10177 (N_10177,N_9386,N_9384);
nor U10178 (N_10178,N_9655,N_9904);
or U10179 (N_10179,N_9917,N_9887);
nor U10180 (N_10180,N_9395,N_9956);
nor U10181 (N_10181,N_9914,N_9435);
and U10182 (N_10182,N_9842,N_9403);
nor U10183 (N_10183,N_9980,N_9801);
and U10184 (N_10184,N_9997,N_9438);
xnor U10185 (N_10185,N_9601,N_9376);
xnor U10186 (N_10186,N_9499,N_9402);
or U10187 (N_10187,N_9547,N_9962);
xor U10188 (N_10188,N_9793,N_9511);
or U10189 (N_10189,N_9746,N_9393);
xor U10190 (N_10190,N_9578,N_9684);
nand U10191 (N_10191,N_9909,N_9819);
nor U10192 (N_10192,N_9831,N_9954);
nand U10193 (N_10193,N_9892,N_9523);
nand U10194 (N_10194,N_9552,N_9571);
nor U10195 (N_10195,N_9462,N_9416);
xor U10196 (N_10196,N_9996,N_9911);
nor U10197 (N_10197,N_9868,N_9975);
and U10198 (N_10198,N_9579,N_9854);
nand U10199 (N_10199,N_9514,N_9466);
nor U10200 (N_10200,N_9605,N_9994);
nor U10201 (N_10201,N_9830,N_9961);
nor U10202 (N_10202,N_9770,N_9529);
nor U10203 (N_10203,N_9776,N_9692);
xor U10204 (N_10204,N_9485,N_9584);
nor U10205 (N_10205,N_9537,N_9448);
nor U10206 (N_10206,N_9931,N_9859);
xor U10207 (N_10207,N_9672,N_9568);
xor U10208 (N_10208,N_9921,N_9955);
or U10209 (N_10209,N_9704,N_9489);
and U10210 (N_10210,N_9992,N_9467);
xnor U10211 (N_10211,N_9689,N_9683);
xor U10212 (N_10212,N_9834,N_9569);
or U10213 (N_10213,N_9881,N_9910);
nor U10214 (N_10214,N_9419,N_9781);
nor U10215 (N_10215,N_9719,N_9977);
xnor U10216 (N_10216,N_9473,N_9544);
nand U10217 (N_10217,N_9730,N_9805);
nor U10218 (N_10218,N_9627,N_9563);
nand U10219 (N_10219,N_9661,N_9551);
nor U10220 (N_10220,N_9637,N_9420);
and U10221 (N_10221,N_9708,N_9548);
xnor U10222 (N_10222,N_9472,N_9907);
nor U10223 (N_10223,N_9469,N_9858);
nor U10224 (N_10224,N_9428,N_9985);
xor U10225 (N_10225,N_9915,N_9922);
or U10226 (N_10226,N_9454,N_9933);
nor U10227 (N_10227,N_9622,N_9494);
and U10228 (N_10228,N_9646,N_9519);
or U10229 (N_10229,N_9795,N_9453);
or U10230 (N_10230,N_9950,N_9818);
and U10231 (N_10231,N_9703,N_9480);
xor U10232 (N_10232,N_9449,N_9542);
or U10233 (N_10233,N_9680,N_9813);
or U10234 (N_10234,N_9828,N_9939);
nor U10235 (N_10235,N_9762,N_9844);
or U10236 (N_10236,N_9779,N_9377);
or U10237 (N_10237,N_9463,N_9602);
and U10238 (N_10238,N_9538,N_9934);
xnor U10239 (N_10239,N_9853,N_9460);
nor U10240 (N_10240,N_9959,N_9434);
nor U10241 (N_10241,N_9409,N_9715);
nor U10242 (N_10242,N_9617,N_9660);
nand U10243 (N_10243,N_9662,N_9400);
nor U10244 (N_10244,N_9750,N_9484);
and U10245 (N_10245,N_9557,N_9391);
xor U10246 (N_10246,N_9481,N_9422);
nand U10247 (N_10247,N_9394,N_9825);
nand U10248 (N_10248,N_9873,N_9446);
or U10249 (N_10249,N_9712,N_9490);
nand U10250 (N_10250,N_9780,N_9528);
nor U10251 (N_10251,N_9613,N_9654);
and U10252 (N_10252,N_9383,N_9582);
nand U10253 (N_10253,N_9558,N_9441);
and U10254 (N_10254,N_9423,N_9664);
or U10255 (N_10255,N_9946,N_9832);
or U10256 (N_10256,N_9636,N_9550);
xor U10257 (N_10257,N_9864,N_9401);
and U10258 (N_10258,N_9555,N_9535);
xnor U10259 (N_10259,N_9432,N_9667);
or U10260 (N_10260,N_9439,N_9653);
nand U10261 (N_10261,N_9741,N_9876);
nor U10262 (N_10262,N_9596,N_9752);
nand U10263 (N_10263,N_9812,N_9679);
nor U10264 (N_10264,N_9846,N_9953);
xor U10265 (N_10265,N_9483,N_9952);
nor U10266 (N_10266,N_9540,N_9503);
nor U10267 (N_10267,N_9738,N_9554);
and U10268 (N_10268,N_9706,N_9871);
nand U10269 (N_10269,N_9634,N_9903);
nand U10270 (N_10270,N_9585,N_9669);
and U10271 (N_10271,N_9429,N_9663);
or U10272 (N_10272,N_9841,N_9459);
and U10273 (N_10273,N_9700,N_9969);
xor U10274 (N_10274,N_9693,N_9736);
nor U10275 (N_10275,N_9541,N_9808);
xor U10276 (N_10276,N_9456,N_9882);
nor U10277 (N_10277,N_9549,N_9799);
nand U10278 (N_10278,N_9588,N_9510);
nor U10279 (N_10279,N_9732,N_9824);
nand U10280 (N_10280,N_9643,N_9748);
nand U10281 (N_10281,N_9407,N_9935);
and U10282 (N_10282,N_9788,N_9623);
or U10283 (N_10283,N_9635,N_9747);
xnor U10284 (N_10284,N_9606,N_9998);
xnor U10285 (N_10285,N_9468,N_9949);
and U10286 (N_10286,N_9800,N_9822);
nand U10287 (N_10287,N_9657,N_9798);
and U10288 (N_10288,N_9885,N_9699);
nand U10289 (N_10289,N_9504,N_9862);
xor U10290 (N_10290,N_9867,N_9927);
and U10291 (N_10291,N_9573,N_9999);
nor U10292 (N_10292,N_9986,N_9621);
or U10293 (N_10293,N_9413,N_9543);
xor U10294 (N_10294,N_9559,N_9916);
xor U10295 (N_10295,N_9943,N_9731);
xor U10296 (N_10296,N_9426,N_9924);
and U10297 (N_10297,N_9773,N_9713);
nor U10298 (N_10298,N_9865,N_9974);
nand U10299 (N_10299,N_9702,N_9380);
nand U10300 (N_10300,N_9863,N_9493);
and U10301 (N_10301,N_9427,N_9436);
xnor U10302 (N_10302,N_9648,N_9630);
or U10303 (N_10303,N_9889,N_9609);
or U10304 (N_10304,N_9908,N_9614);
nor U10305 (N_10305,N_9901,N_9592);
nor U10306 (N_10306,N_9725,N_9546);
or U10307 (N_10307,N_9418,N_9522);
nor U10308 (N_10308,N_9896,N_9815);
or U10309 (N_10309,N_9970,N_9843);
or U10310 (N_10310,N_9412,N_9398);
xor U10311 (N_10311,N_9753,N_9659);
and U10312 (N_10312,N_9905,N_9851);
nor U10313 (N_10313,N_9423,N_9807);
nor U10314 (N_10314,N_9898,N_9451);
nand U10315 (N_10315,N_9566,N_9531);
xor U10316 (N_10316,N_9863,N_9922);
or U10317 (N_10317,N_9404,N_9435);
xnor U10318 (N_10318,N_9956,N_9412);
and U10319 (N_10319,N_9959,N_9847);
and U10320 (N_10320,N_9846,N_9393);
nor U10321 (N_10321,N_9889,N_9872);
nand U10322 (N_10322,N_9792,N_9428);
nand U10323 (N_10323,N_9736,N_9401);
nand U10324 (N_10324,N_9923,N_9862);
nor U10325 (N_10325,N_9850,N_9908);
nand U10326 (N_10326,N_9937,N_9380);
nor U10327 (N_10327,N_9940,N_9540);
xor U10328 (N_10328,N_9974,N_9501);
and U10329 (N_10329,N_9548,N_9436);
or U10330 (N_10330,N_9958,N_9849);
and U10331 (N_10331,N_9933,N_9667);
xnor U10332 (N_10332,N_9647,N_9573);
or U10333 (N_10333,N_9821,N_9706);
nand U10334 (N_10334,N_9477,N_9937);
nand U10335 (N_10335,N_9876,N_9773);
xnor U10336 (N_10336,N_9466,N_9547);
nand U10337 (N_10337,N_9697,N_9490);
xnor U10338 (N_10338,N_9628,N_9646);
xnor U10339 (N_10339,N_9520,N_9396);
nand U10340 (N_10340,N_9458,N_9377);
nor U10341 (N_10341,N_9724,N_9696);
nor U10342 (N_10342,N_9531,N_9927);
nor U10343 (N_10343,N_9772,N_9589);
nor U10344 (N_10344,N_9918,N_9652);
or U10345 (N_10345,N_9971,N_9842);
or U10346 (N_10346,N_9651,N_9741);
xnor U10347 (N_10347,N_9966,N_9445);
or U10348 (N_10348,N_9823,N_9980);
or U10349 (N_10349,N_9723,N_9960);
nand U10350 (N_10350,N_9573,N_9902);
nand U10351 (N_10351,N_9522,N_9991);
xnor U10352 (N_10352,N_9564,N_9949);
nor U10353 (N_10353,N_9941,N_9968);
nand U10354 (N_10354,N_9992,N_9460);
nand U10355 (N_10355,N_9577,N_9642);
or U10356 (N_10356,N_9858,N_9866);
xor U10357 (N_10357,N_9989,N_9703);
or U10358 (N_10358,N_9800,N_9949);
xor U10359 (N_10359,N_9389,N_9418);
nand U10360 (N_10360,N_9385,N_9607);
or U10361 (N_10361,N_9710,N_9784);
nand U10362 (N_10362,N_9727,N_9683);
and U10363 (N_10363,N_9840,N_9381);
nor U10364 (N_10364,N_9618,N_9686);
and U10365 (N_10365,N_9748,N_9792);
and U10366 (N_10366,N_9544,N_9619);
xnor U10367 (N_10367,N_9772,N_9828);
nor U10368 (N_10368,N_9729,N_9516);
and U10369 (N_10369,N_9619,N_9975);
nand U10370 (N_10370,N_9729,N_9823);
and U10371 (N_10371,N_9919,N_9570);
or U10372 (N_10372,N_9864,N_9487);
or U10373 (N_10373,N_9691,N_9817);
nor U10374 (N_10374,N_9496,N_9536);
nand U10375 (N_10375,N_9902,N_9943);
xor U10376 (N_10376,N_9568,N_9972);
and U10377 (N_10377,N_9846,N_9986);
nand U10378 (N_10378,N_9736,N_9628);
nor U10379 (N_10379,N_9526,N_9878);
xor U10380 (N_10380,N_9495,N_9777);
nor U10381 (N_10381,N_9719,N_9829);
nor U10382 (N_10382,N_9737,N_9888);
and U10383 (N_10383,N_9502,N_9868);
xor U10384 (N_10384,N_9653,N_9818);
or U10385 (N_10385,N_9465,N_9513);
nand U10386 (N_10386,N_9524,N_9379);
nand U10387 (N_10387,N_9651,N_9765);
and U10388 (N_10388,N_9625,N_9907);
nor U10389 (N_10389,N_9856,N_9633);
xor U10390 (N_10390,N_9779,N_9443);
nand U10391 (N_10391,N_9630,N_9598);
xor U10392 (N_10392,N_9419,N_9384);
nand U10393 (N_10393,N_9462,N_9414);
and U10394 (N_10394,N_9656,N_9752);
xnor U10395 (N_10395,N_9785,N_9859);
and U10396 (N_10396,N_9944,N_9504);
nor U10397 (N_10397,N_9995,N_9730);
or U10398 (N_10398,N_9744,N_9507);
or U10399 (N_10399,N_9607,N_9490);
nor U10400 (N_10400,N_9875,N_9727);
or U10401 (N_10401,N_9558,N_9818);
nor U10402 (N_10402,N_9476,N_9953);
and U10403 (N_10403,N_9961,N_9833);
and U10404 (N_10404,N_9831,N_9728);
and U10405 (N_10405,N_9665,N_9963);
and U10406 (N_10406,N_9553,N_9737);
nor U10407 (N_10407,N_9872,N_9780);
xor U10408 (N_10408,N_9480,N_9410);
xnor U10409 (N_10409,N_9992,N_9500);
or U10410 (N_10410,N_9616,N_9651);
nand U10411 (N_10411,N_9725,N_9711);
or U10412 (N_10412,N_9678,N_9605);
xnor U10413 (N_10413,N_9477,N_9786);
or U10414 (N_10414,N_9538,N_9897);
xor U10415 (N_10415,N_9729,N_9535);
nand U10416 (N_10416,N_9627,N_9512);
and U10417 (N_10417,N_9885,N_9478);
nor U10418 (N_10418,N_9454,N_9555);
and U10419 (N_10419,N_9938,N_9479);
or U10420 (N_10420,N_9773,N_9730);
and U10421 (N_10421,N_9746,N_9969);
nor U10422 (N_10422,N_9453,N_9963);
nand U10423 (N_10423,N_9775,N_9487);
nand U10424 (N_10424,N_9853,N_9991);
or U10425 (N_10425,N_9378,N_9969);
or U10426 (N_10426,N_9722,N_9378);
and U10427 (N_10427,N_9427,N_9623);
and U10428 (N_10428,N_9812,N_9819);
nor U10429 (N_10429,N_9678,N_9824);
xor U10430 (N_10430,N_9733,N_9392);
xnor U10431 (N_10431,N_9496,N_9805);
and U10432 (N_10432,N_9472,N_9791);
nand U10433 (N_10433,N_9539,N_9621);
and U10434 (N_10434,N_9900,N_9928);
nor U10435 (N_10435,N_9836,N_9877);
nor U10436 (N_10436,N_9882,N_9590);
and U10437 (N_10437,N_9612,N_9564);
xor U10438 (N_10438,N_9914,N_9813);
nand U10439 (N_10439,N_9736,N_9629);
nor U10440 (N_10440,N_9880,N_9656);
and U10441 (N_10441,N_9469,N_9568);
or U10442 (N_10442,N_9478,N_9815);
xnor U10443 (N_10443,N_9590,N_9681);
xor U10444 (N_10444,N_9893,N_9452);
and U10445 (N_10445,N_9858,N_9558);
xnor U10446 (N_10446,N_9649,N_9492);
nand U10447 (N_10447,N_9419,N_9463);
nand U10448 (N_10448,N_9659,N_9399);
nand U10449 (N_10449,N_9778,N_9515);
nor U10450 (N_10450,N_9964,N_9967);
and U10451 (N_10451,N_9665,N_9889);
nor U10452 (N_10452,N_9993,N_9470);
or U10453 (N_10453,N_9683,N_9404);
nand U10454 (N_10454,N_9394,N_9490);
nor U10455 (N_10455,N_9836,N_9922);
and U10456 (N_10456,N_9678,N_9519);
and U10457 (N_10457,N_9855,N_9784);
xnor U10458 (N_10458,N_9576,N_9739);
nand U10459 (N_10459,N_9396,N_9681);
or U10460 (N_10460,N_9905,N_9979);
and U10461 (N_10461,N_9557,N_9773);
or U10462 (N_10462,N_9906,N_9768);
and U10463 (N_10463,N_9696,N_9718);
nand U10464 (N_10464,N_9760,N_9905);
or U10465 (N_10465,N_9919,N_9800);
xnor U10466 (N_10466,N_9816,N_9489);
nand U10467 (N_10467,N_9882,N_9938);
or U10468 (N_10468,N_9931,N_9612);
nor U10469 (N_10469,N_9479,N_9545);
nand U10470 (N_10470,N_9609,N_9627);
nor U10471 (N_10471,N_9457,N_9923);
nor U10472 (N_10472,N_9921,N_9722);
and U10473 (N_10473,N_9713,N_9792);
nor U10474 (N_10474,N_9541,N_9639);
and U10475 (N_10475,N_9482,N_9417);
and U10476 (N_10476,N_9442,N_9497);
and U10477 (N_10477,N_9770,N_9932);
xnor U10478 (N_10478,N_9911,N_9975);
and U10479 (N_10479,N_9520,N_9956);
and U10480 (N_10480,N_9866,N_9624);
or U10481 (N_10481,N_9389,N_9611);
and U10482 (N_10482,N_9999,N_9887);
or U10483 (N_10483,N_9736,N_9969);
and U10484 (N_10484,N_9859,N_9866);
xor U10485 (N_10485,N_9847,N_9777);
or U10486 (N_10486,N_9503,N_9505);
nor U10487 (N_10487,N_9940,N_9429);
nor U10488 (N_10488,N_9482,N_9689);
or U10489 (N_10489,N_9707,N_9583);
xor U10490 (N_10490,N_9818,N_9964);
and U10491 (N_10491,N_9883,N_9493);
xnor U10492 (N_10492,N_9823,N_9723);
nand U10493 (N_10493,N_9443,N_9974);
xnor U10494 (N_10494,N_9447,N_9990);
xnor U10495 (N_10495,N_9702,N_9591);
nand U10496 (N_10496,N_9725,N_9672);
or U10497 (N_10497,N_9723,N_9842);
xor U10498 (N_10498,N_9547,N_9943);
or U10499 (N_10499,N_9408,N_9607);
xor U10500 (N_10500,N_9854,N_9404);
and U10501 (N_10501,N_9828,N_9782);
nor U10502 (N_10502,N_9481,N_9644);
and U10503 (N_10503,N_9861,N_9808);
xnor U10504 (N_10504,N_9896,N_9902);
nor U10505 (N_10505,N_9514,N_9735);
nor U10506 (N_10506,N_9706,N_9995);
and U10507 (N_10507,N_9883,N_9505);
or U10508 (N_10508,N_9652,N_9494);
or U10509 (N_10509,N_9772,N_9767);
nor U10510 (N_10510,N_9452,N_9555);
or U10511 (N_10511,N_9590,N_9619);
nor U10512 (N_10512,N_9546,N_9507);
and U10513 (N_10513,N_9844,N_9701);
or U10514 (N_10514,N_9803,N_9675);
xor U10515 (N_10515,N_9994,N_9408);
nor U10516 (N_10516,N_9622,N_9384);
and U10517 (N_10517,N_9810,N_9605);
and U10518 (N_10518,N_9519,N_9942);
or U10519 (N_10519,N_9439,N_9921);
nand U10520 (N_10520,N_9481,N_9483);
nor U10521 (N_10521,N_9512,N_9402);
nand U10522 (N_10522,N_9674,N_9807);
and U10523 (N_10523,N_9893,N_9681);
nand U10524 (N_10524,N_9972,N_9978);
nor U10525 (N_10525,N_9580,N_9811);
nand U10526 (N_10526,N_9543,N_9810);
and U10527 (N_10527,N_9847,N_9477);
xor U10528 (N_10528,N_9996,N_9406);
nand U10529 (N_10529,N_9822,N_9556);
xor U10530 (N_10530,N_9411,N_9628);
xnor U10531 (N_10531,N_9575,N_9999);
xnor U10532 (N_10532,N_9548,N_9617);
nand U10533 (N_10533,N_9800,N_9763);
nand U10534 (N_10534,N_9594,N_9945);
or U10535 (N_10535,N_9970,N_9727);
or U10536 (N_10536,N_9439,N_9786);
and U10537 (N_10537,N_9417,N_9762);
and U10538 (N_10538,N_9586,N_9902);
xor U10539 (N_10539,N_9642,N_9757);
nand U10540 (N_10540,N_9665,N_9980);
or U10541 (N_10541,N_9618,N_9651);
or U10542 (N_10542,N_9883,N_9800);
nand U10543 (N_10543,N_9878,N_9684);
or U10544 (N_10544,N_9789,N_9850);
nor U10545 (N_10545,N_9702,N_9870);
nand U10546 (N_10546,N_9671,N_9533);
xor U10547 (N_10547,N_9561,N_9654);
nand U10548 (N_10548,N_9441,N_9950);
nor U10549 (N_10549,N_9558,N_9761);
xor U10550 (N_10550,N_9453,N_9657);
and U10551 (N_10551,N_9691,N_9916);
or U10552 (N_10552,N_9870,N_9849);
and U10553 (N_10553,N_9949,N_9822);
nand U10554 (N_10554,N_9968,N_9456);
nor U10555 (N_10555,N_9455,N_9868);
and U10556 (N_10556,N_9445,N_9464);
xor U10557 (N_10557,N_9931,N_9734);
xor U10558 (N_10558,N_9711,N_9475);
nand U10559 (N_10559,N_9839,N_9934);
and U10560 (N_10560,N_9504,N_9984);
xor U10561 (N_10561,N_9823,N_9915);
or U10562 (N_10562,N_9391,N_9737);
nor U10563 (N_10563,N_9914,N_9608);
nor U10564 (N_10564,N_9845,N_9492);
nand U10565 (N_10565,N_9630,N_9572);
nor U10566 (N_10566,N_9705,N_9711);
or U10567 (N_10567,N_9759,N_9945);
nand U10568 (N_10568,N_9507,N_9435);
nand U10569 (N_10569,N_9886,N_9930);
nor U10570 (N_10570,N_9554,N_9536);
and U10571 (N_10571,N_9973,N_9992);
and U10572 (N_10572,N_9820,N_9791);
and U10573 (N_10573,N_9968,N_9950);
xnor U10574 (N_10574,N_9788,N_9565);
and U10575 (N_10575,N_9785,N_9421);
nand U10576 (N_10576,N_9865,N_9986);
nand U10577 (N_10577,N_9494,N_9426);
xor U10578 (N_10578,N_9614,N_9541);
nor U10579 (N_10579,N_9717,N_9997);
nor U10580 (N_10580,N_9589,N_9379);
nand U10581 (N_10581,N_9757,N_9770);
nor U10582 (N_10582,N_9979,N_9767);
nor U10583 (N_10583,N_9900,N_9479);
and U10584 (N_10584,N_9933,N_9416);
and U10585 (N_10585,N_9546,N_9537);
nor U10586 (N_10586,N_9403,N_9646);
and U10587 (N_10587,N_9788,N_9625);
or U10588 (N_10588,N_9769,N_9998);
and U10589 (N_10589,N_9960,N_9773);
nor U10590 (N_10590,N_9958,N_9845);
and U10591 (N_10591,N_9434,N_9505);
xor U10592 (N_10592,N_9478,N_9796);
nor U10593 (N_10593,N_9864,N_9415);
and U10594 (N_10594,N_9637,N_9959);
and U10595 (N_10595,N_9435,N_9471);
or U10596 (N_10596,N_9535,N_9476);
and U10597 (N_10597,N_9415,N_9888);
nand U10598 (N_10598,N_9620,N_9632);
xnor U10599 (N_10599,N_9581,N_9467);
and U10600 (N_10600,N_9556,N_9537);
xor U10601 (N_10601,N_9447,N_9411);
nand U10602 (N_10602,N_9918,N_9412);
nor U10603 (N_10603,N_9885,N_9653);
and U10604 (N_10604,N_9790,N_9806);
and U10605 (N_10605,N_9670,N_9388);
nand U10606 (N_10606,N_9859,N_9842);
or U10607 (N_10607,N_9912,N_9964);
or U10608 (N_10608,N_9585,N_9947);
nor U10609 (N_10609,N_9779,N_9651);
or U10610 (N_10610,N_9486,N_9995);
xor U10611 (N_10611,N_9772,N_9628);
xnor U10612 (N_10612,N_9954,N_9447);
nor U10613 (N_10613,N_9914,N_9689);
or U10614 (N_10614,N_9815,N_9526);
xor U10615 (N_10615,N_9676,N_9385);
and U10616 (N_10616,N_9647,N_9890);
nor U10617 (N_10617,N_9716,N_9532);
or U10618 (N_10618,N_9638,N_9399);
nand U10619 (N_10619,N_9868,N_9412);
or U10620 (N_10620,N_9488,N_9821);
nor U10621 (N_10621,N_9556,N_9761);
nor U10622 (N_10622,N_9857,N_9378);
xnor U10623 (N_10623,N_9781,N_9888);
nor U10624 (N_10624,N_9468,N_9925);
xnor U10625 (N_10625,N_10321,N_10294);
nor U10626 (N_10626,N_10156,N_10582);
and U10627 (N_10627,N_10237,N_10167);
nand U10628 (N_10628,N_10388,N_10064);
nand U10629 (N_10629,N_10576,N_10322);
nand U10630 (N_10630,N_10245,N_10508);
and U10631 (N_10631,N_10136,N_10225);
and U10632 (N_10632,N_10111,N_10144);
or U10633 (N_10633,N_10300,N_10212);
nand U10634 (N_10634,N_10303,N_10356);
nor U10635 (N_10635,N_10468,N_10330);
nand U10636 (N_10636,N_10423,N_10395);
or U10637 (N_10637,N_10045,N_10147);
xnor U10638 (N_10638,N_10620,N_10062);
and U10639 (N_10639,N_10096,N_10295);
or U10640 (N_10640,N_10099,N_10509);
and U10641 (N_10641,N_10074,N_10059);
and U10642 (N_10642,N_10493,N_10569);
and U10643 (N_10643,N_10396,N_10187);
and U10644 (N_10644,N_10198,N_10407);
or U10645 (N_10645,N_10548,N_10063);
nor U10646 (N_10646,N_10276,N_10171);
or U10647 (N_10647,N_10526,N_10514);
nor U10648 (N_10648,N_10179,N_10476);
xnor U10649 (N_10649,N_10484,N_10457);
nand U10650 (N_10650,N_10140,N_10465);
and U10651 (N_10651,N_10551,N_10302);
xor U10652 (N_10652,N_10405,N_10478);
nand U10653 (N_10653,N_10490,N_10265);
nand U10654 (N_10654,N_10286,N_10350);
nor U10655 (N_10655,N_10539,N_10338);
or U10656 (N_10656,N_10267,N_10596);
or U10657 (N_10657,N_10052,N_10558);
nor U10658 (N_10658,N_10239,N_10009);
and U10659 (N_10659,N_10556,N_10614);
nand U10660 (N_10660,N_10107,N_10199);
or U10661 (N_10661,N_10318,N_10464);
and U10662 (N_10662,N_10126,N_10222);
xnor U10663 (N_10663,N_10005,N_10116);
nand U10664 (N_10664,N_10605,N_10621);
nor U10665 (N_10665,N_10220,N_10599);
nand U10666 (N_10666,N_10354,N_10501);
and U10667 (N_10667,N_10002,N_10175);
nand U10668 (N_10668,N_10349,N_10149);
xor U10669 (N_10669,N_10240,N_10264);
or U10670 (N_10670,N_10304,N_10432);
and U10671 (N_10671,N_10439,N_10309);
nand U10672 (N_10672,N_10194,N_10134);
or U10673 (N_10673,N_10298,N_10458);
or U10674 (N_10674,N_10269,N_10177);
or U10675 (N_10675,N_10412,N_10431);
xnor U10676 (N_10676,N_10219,N_10221);
and U10677 (N_10677,N_10447,N_10244);
or U10678 (N_10678,N_10437,N_10340);
or U10679 (N_10679,N_10320,N_10095);
and U10680 (N_10680,N_10131,N_10335);
and U10681 (N_10681,N_10544,N_10342);
nand U10682 (N_10682,N_10402,N_10281);
nor U10683 (N_10683,N_10319,N_10532);
nor U10684 (N_10684,N_10311,N_10477);
nor U10685 (N_10685,N_10504,N_10624);
or U10686 (N_10686,N_10085,N_10553);
and U10687 (N_10687,N_10380,N_10475);
nor U10688 (N_10688,N_10176,N_10128);
nor U10689 (N_10689,N_10157,N_10251);
nor U10690 (N_10690,N_10016,N_10248);
xor U10691 (N_10691,N_10538,N_10077);
or U10692 (N_10692,N_10056,N_10589);
nor U10693 (N_10693,N_10399,N_10060);
xnor U10694 (N_10694,N_10270,N_10293);
and U10695 (N_10695,N_10272,N_10352);
xor U10696 (N_10696,N_10084,N_10141);
xor U10697 (N_10697,N_10263,N_10332);
nor U10698 (N_10698,N_10604,N_10507);
xor U10699 (N_10699,N_10215,N_10491);
and U10700 (N_10700,N_10425,N_10463);
nor U10701 (N_10701,N_10414,N_10154);
and U10702 (N_10702,N_10571,N_10090);
nand U10703 (N_10703,N_10190,N_10500);
nand U10704 (N_10704,N_10257,N_10210);
nor U10705 (N_10705,N_10075,N_10474);
and U10706 (N_10706,N_10573,N_10071);
or U10707 (N_10707,N_10602,N_10334);
or U10708 (N_10708,N_10313,N_10622);
or U10709 (N_10709,N_10361,N_10527);
and U10710 (N_10710,N_10051,N_10003);
or U10711 (N_10711,N_10242,N_10470);
nand U10712 (N_10712,N_10578,N_10201);
and U10713 (N_10713,N_10254,N_10381);
nand U10714 (N_10714,N_10452,N_10205);
nor U10715 (N_10715,N_10284,N_10502);
nand U10716 (N_10716,N_10410,N_10442);
nor U10717 (N_10717,N_10089,N_10329);
and U10718 (N_10718,N_10387,N_10482);
nor U10719 (N_10719,N_10486,N_10427);
or U10720 (N_10720,N_10574,N_10555);
xor U10721 (N_10721,N_10181,N_10013);
or U10722 (N_10722,N_10278,N_10531);
xnor U10723 (N_10723,N_10554,N_10441);
and U10724 (N_10724,N_10367,N_10103);
and U10725 (N_10725,N_10042,N_10448);
or U10726 (N_10726,N_10068,N_10364);
xnor U10727 (N_10727,N_10080,N_10580);
xor U10728 (N_10728,N_10515,N_10454);
or U10729 (N_10729,N_10250,N_10236);
and U10730 (N_10730,N_10218,N_10228);
nand U10731 (N_10731,N_10344,N_10216);
and U10732 (N_10732,N_10044,N_10362);
nor U10733 (N_10733,N_10192,N_10168);
xor U10734 (N_10734,N_10200,N_10496);
xnor U10735 (N_10735,N_10472,N_10301);
xnor U10736 (N_10736,N_10041,N_10160);
xor U10737 (N_10737,N_10413,N_10565);
nand U10738 (N_10738,N_10460,N_10488);
and U10739 (N_10739,N_10162,N_10266);
nor U10740 (N_10740,N_10253,N_10235);
and U10741 (N_10741,N_10004,N_10389);
nor U10742 (N_10742,N_10393,N_10489);
xor U10743 (N_10743,N_10053,N_10241);
or U10744 (N_10744,N_10196,N_10048);
or U10745 (N_10745,N_10542,N_10503);
nand U10746 (N_10746,N_10082,N_10261);
nand U10747 (N_10747,N_10007,N_10050);
xnor U10748 (N_10748,N_10383,N_10310);
nor U10749 (N_10749,N_10583,N_10069);
and U10750 (N_10750,N_10469,N_10424);
xnor U10751 (N_10751,N_10451,N_10481);
nor U10752 (N_10752,N_10015,N_10588);
xor U10753 (N_10753,N_10043,N_10203);
xor U10754 (N_10754,N_10487,N_10365);
xor U10755 (N_10755,N_10535,N_10592);
and U10756 (N_10756,N_10204,N_10260);
nand U10757 (N_10757,N_10453,N_10135);
nor U10758 (N_10758,N_10230,N_10390);
and U10759 (N_10759,N_10234,N_10331);
xnor U10760 (N_10760,N_10594,N_10185);
nor U10761 (N_10761,N_10382,N_10581);
nand U10762 (N_10762,N_10000,N_10081);
nor U10763 (N_10763,N_10597,N_10540);
nor U10764 (N_10764,N_10434,N_10151);
and U10765 (N_10765,N_10512,N_10110);
xnor U10766 (N_10766,N_10546,N_10567);
nand U10767 (N_10767,N_10568,N_10559);
nor U10768 (N_10768,N_10288,N_10392);
and U10769 (N_10769,N_10169,N_10208);
nand U10770 (N_10770,N_10557,N_10146);
nand U10771 (N_10771,N_10530,N_10566);
nor U10772 (N_10772,N_10223,N_10207);
nor U10773 (N_10773,N_10249,N_10355);
and U10774 (N_10774,N_10017,N_10353);
nor U10775 (N_10775,N_10229,N_10455);
and U10776 (N_10776,N_10022,N_10271);
or U10777 (N_10777,N_10426,N_10188);
and U10778 (N_10778,N_10613,N_10109);
nand U10779 (N_10779,N_10522,N_10511);
and U10780 (N_10780,N_10438,N_10255);
nor U10781 (N_10781,N_10243,N_10485);
nand U10782 (N_10782,N_10498,N_10608);
and U10783 (N_10783,N_10384,N_10397);
xor U10784 (N_10784,N_10366,N_10586);
nand U10785 (N_10785,N_10623,N_10195);
nor U10786 (N_10786,N_10315,N_10280);
nor U10787 (N_10787,N_10363,N_10445);
nand U10788 (N_10788,N_10379,N_10088);
xnor U10789 (N_10789,N_10585,N_10520);
and U10790 (N_10790,N_10391,N_10214);
or U10791 (N_10791,N_10117,N_10370);
xnor U10792 (N_10792,N_10070,N_10411);
xor U10793 (N_10793,N_10600,N_10341);
nand U10794 (N_10794,N_10180,N_10087);
and U10795 (N_10795,N_10152,N_10609);
or U10796 (N_10796,N_10430,N_10505);
xnor U10797 (N_10797,N_10415,N_10227);
nor U10798 (N_10798,N_10590,N_10078);
nor U10799 (N_10799,N_10516,N_10076);
nand U10800 (N_10800,N_10521,N_10118);
xor U10801 (N_10801,N_10037,N_10183);
nor U10802 (N_10802,N_10419,N_10114);
nand U10803 (N_10803,N_10357,N_10466);
or U10804 (N_10804,N_10209,N_10549);
xnor U10805 (N_10805,N_10579,N_10404);
nor U10806 (N_10806,N_10065,N_10150);
and U10807 (N_10807,N_10433,N_10036);
and U10808 (N_10808,N_10057,N_10417);
and U10809 (N_10809,N_10400,N_10137);
and U10810 (N_10810,N_10058,N_10011);
and U10811 (N_10811,N_10471,N_10495);
xnor U10812 (N_10812,N_10348,N_10273);
or U10813 (N_10813,N_10497,N_10038);
xnor U10814 (N_10814,N_10106,N_10232);
or U10815 (N_10815,N_10347,N_10577);
nand U10816 (N_10816,N_10186,N_10224);
xnor U10817 (N_10817,N_10494,N_10610);
nor U10818 (N_10818,N_10023,N_10299);
and U10819 (N_10819,N_10473,N_10336);
or U10820 (N_10820,N_10086,N_10525);
or U10821 (N_10821,N_10001,N_10155);
and U10822 (N_10822,N_10429,N_10305);
nor U10823 (N_10823,N_10373,N_10256);
and U10824 (N_10824,N_10115,N_10285);
nand U10825 (N_10825,N_10105,N_10572);
xor U10826 (N_10826,N_10359,N_10523);
and U10827 (N_10827,N_10297,N_10378);
xnor U10828 (N_10828,N_10345,N_10132);
and U10829 (N_10829,N_10158,N_10587);
xnor U10830 (N_10830,N_10025,N_10534);
nand U10831 (N_10831,N_10591,N_10039);
xnor U10832 (N_10832,N_10593,N_10125);
nor U10833 (N_10833,N_10283,N_10275);
and U10834 (N_10834,N_10462,N_10282);
nor U10835 (N_10835,N_10461,N_10337);
nor U10836 (N_10836,N_10121,N_10279);
or U10837 (N_10837,N_10563,N_10124);
and U10838 (N_10838,N_10010,N_10166);
and U10839 (N_10839,N_10371,N_10324);
xor U10840 (N_10840,N_10130,N_10161);
and U10841 (N_10841,N_10312,N_10385);
and U10842 (N_10842,N_10327,N_10524);
xnor U10843 (N_10843,N_10346,N_10323);
xnor U10844 (N_10844,N_10550,N_10211);
nand U10845 (N_10845,N_10032,N_10376);
and U10846 (N_10846,N_10450,N_10499);
nor U10847 (N_10847,N_10061,N_10422);
nand U10848 (N_10848,N_10326,N_10193);
or U10849 (N_10849,N_10091,N_10047);
xor U10850 (N_10850,N_10416,N_10449);
or U10851 (N_10851,N_10307,N_10617);
and U10852 (N_10852,N_10164,N_10226);
xor U10853 (N_10853,N_10612,N_10231);
and U10854 (N_10854,N_10174,N_10092);
xor U10855 (N_10855,N_10619,N_10163);
nor U10856 (N_10856,N_10142,N_10428);
or U10857 (N_10857,N_10197,N_10533);
xnor U10858 (N_10858,N_10277,N_10072);
nor U10859 (N_10859,N_10238,N_10459);
nand U10860 (N_10860,N_10360,N_10456);
and U10861 (N_10861,N_10306,N_10386);
or U10862 (N_10862,N_10601,N_10394);
and U10863 (N_10863,N_10570,N_10561);
or U10864 (N_10864,N_10153,N_10054);
xnor U10865 (N_10865,N_10444,N_10374);
or U10866 (N_10866,N_10541,N_10552);
nand U10867 (N_10867,N_10406,N_10104);
or U10868 (N_10868,N_10372,N_10420);
nand U10869 (N_10869,N_10020,N_10006);
xnor U10870 (N_10870,N_10079,N_10202);
nor U10871 (N_10871,N_10100,N_10049);
nor U10872 (N_10872,N_10316,N_10518);
nand U10873 (N_10873,N_10409,N_10102);
nor U10874 (N_10874,N_10246,N_10019);
xnor U10875 (N_10875,N_10519,N_10435);
nand U10876 (N_10876,N_10119,N_10480);
nand U10877 (N_10877,N_10517,N_10606);
xnor U10878 (N_10878,N_10217,N_10268);
nor U10879 (N_10879,N_10401,N_10206);
xnor U10880 (N_10880,N_10618,N_10012);
xnor U10881 (N_10881,N_10607,N_10536);
nor U10882 (N_10882,N_10028,N_10528);
and U10883 (N_10883,N_10339,N_10446);
nor U10884 (N_10884,N_10259,N_10008);
xnor U10885 (N_10885,N_10421,N_10014);
nand U10886 (N_10886,N_10513,N_10408);
nor U10887 (N_10887,N_10184,N_10040);
and U10888 (N_10888,N_10398,N_10024);
nor U10889 (N_10889,N_10584,N_10545);
and U10890 (N_10890,N_10467,N_10560);
nor U10891 (N_10891,N_10443,N_10120);
xnor U10892 (N_10892,N_10289,N_10314);
nand U10893 (N_10893,N_10066,N_10030);
and U10894 (N_10894,N_10479,N_10325);
and U10895 (N_10895,N_10287,N_10138);
nand U10896 (N_10896,N_10213,N_10375);
and U10897 (N_10897,N_10133,N_10369);
and U10898 (N_10898,N_10317,N_10093);
nor U10899 (N_10899,N_10543,N_10252);
and U10900 (N_10900,N_10575,N_10182);
xor U10901 (N_10901,N_10094,N_10562);
or U10902 (N_10902,N_10127,N_10296);
and U10903 (N_10903,N_10035,N_10510);
nor U10904 (N_10904,N_10148,N_10178);
nand U10905 (N_10905,N_10483,N_10122);
or U10906 (N_10906,N_10189,N_10595);
and U10907 (N_10907,N_10159,N_10027);
or U10908 (N_10908,N_10247,N_10172);
nor U10909 (N_10909,N_10191,N_10615);
nor U10910 (N_10910,N_10073,N_10258);
xnor U10911 (N_10911,N_10537,N_10112);
xnor U10912 (N_10912,N_10129,N_10291);
nor U10913 (N_10913,N_10021,N_10274);
xnor U10914 (N_10914,N_10143,N_10083);
xnor U10915 (N_10915,N_10603,N_10018);
xor U10916 (N_10916,N_10165,N_10611);
or U10917 (N_10917,N_10598,N_10173);
or U10918 (N_10918,N_10098,N_10292);
xnor U10919 (N_10919,N_10055,N_10377);
nand U10920 (N_10920,N_10139,N_10113);
xor U10921 (N_10921,N_10108,N_10262);
or U10922 (N_10922,N_10031,N_10403);
nand U10923 (N_10923,N_10233,N_10351);
nor U10924 (N_10924,N_10529,N_10067);
xor U10925 (N_10925,N_10046,N_10616);
nor U10926 (N_10926,N_10123,N_10170);
xor U10927 (N_10927,N_10358,N_10436);
xnor U10928 (N_10928,N_10029,N_10101);
nand U10929 (N_10929,N_10308,N_10492);
xnor U10930 (N_10930,N_10034,N_10145);
or U10931 (N_10931,N_10418,N_10440);
or U10932 (N_10932,N_10290,N_10506);
or U10933 (N_10933,N_10328,N_10026);
and U10934 (N_10934,N_10368,N_10333);
nor U10935 (N_10935,N_10564,N_10033);
or U10936 (N_10936,N_10343,N_10097);
or U10937 (N_10937,N_10547,N_10503);
nor U10938 (N_10938,N_10277,N_10100);
or U10939 (N_10939,N_10606,N_10335);
xor U10940 (N_10940,N_10466,N_10012);
nor U10941 (N_10941,N_10312,N_10623);
nand U10942 (N_10942,N_10098,N_10263);
nand U10943 (N_10943,N_10488,N_10570);
nor U10944 (N_10944,N_10376,N_10284);
and U10945 (N_10945,N_10000,N_10235);
xor U10946 (N_10946,N_10222,N_10277);
xnor U10947 (N_10947,N_10188,N_10153);
nor U10948 (N_10948,N_10006,N_10356);
nor U10949 (N_10949,N_10259,N_10183);
and U10950 (N_10950,N_10097,N_10492);
nor U10951 (N_10951,N_10534,N_10278);
nand U10952 (N_10952,N_10017,N_10540);
nor U10953 (N_10953,N_10037,N_10056);
and U10954 (N_10954,N_10579,N_10609);
nor U10955 (N_10955,N_10277,N_10009);
and U10956 (N_10956,N_10182,N_10075);
and U10957 (N_10957,N_10184,N_10377);
nand U10958 (N_10958,N_10033,N_10129);
and U10959 (N_10959,N_10026,N_10117);
nand U10960 (N_10960,N_10340,N_10551);
and U10961 (N_10961,N_10592,N_10438);
nor U10962 (N_10962,N_10543,N_10006);
xnor U10963 (N_10963,N_10093,N_10139);
or U10964 (N_10964,N_10127,N_10267);
nand U10965 (N_10965,N_10322,N_10512);
or U10966 (N_10966,N_10600,N_10283);
nand U10967 (N_10967,N_10097,N_10179);
xnor U10968 (N_10968,N_10550,N_10158);
nor U10969 (N_10969,N_10372,N_10336);
nand U10970 (N_10970,N_10423,N_10188);
nor U10971 (N_10971,N_10014,N_10457);
xnor U10972 (N_10972,N_10533,N_10353);
or U10973 (N_10973,N_10572,N_10169);
xor U10974 (N_10974,N_10172,N_10344);
or U10975 (N_10975,N_10104,N_10102);
xnor U10976 (N_10976,N_10339,N_10146);
and U10977 (N_10977,N_10010,N_10576);
nor U10978 (N_10978,N_10392,N_10284);
xnor U10979 (N_10979,N_10521,N_10405);
xnor U10980 (N_10980,N_10122,N_10518);
nor U10981 (N_10981,N_10520,N_10521);
nor U10982 (N_10982,N_10237,N_10078);
nor U10983 (N_10983,N_10163,N_10495);
nor U10984 (N_10984,N_10234,N_10600);
or U10985 (N_10985,N_10282,N_10034);
nand U10986 (N_10986,N_10421,N_10520);
xor U10987 (N_10987,N_10305,N_10470);
and U10988 (N_10988,N_10107,N_10604);
nor U10989 (N_10989,N_10194,N_10580);
nand U10990 (N_10990,N_10525,N_10523);
nor U10991 (N_10991,N_10053,N_10609);
or U10992 (N_10992,N_10401,N_10242);
xnor U10993 (N_10993,N_10364,N_10345);
and U10994 (N_10994,N_10300,N_10192);
nand U10995 (N_10995,N_10202,N_10104);
or U10996 (N_10996,N_10177,N_10133);
nand U10997 (N_10997,N_10019,N_10535);
or U10998 (N_10998,N_10519,N_10596);
nand U10999 (N_10999,N_10328,N_10374);
and U11000 (N_11000,N_10520,N_10532);
nor U11001 (N_11001,N_10100,N_10290);
xor U11002 (N_11002,N_10094,N_10006);
nor U11003 (N_11003,N_10443,N_10617);
and U11004 (N_11004,N_10201,N_10565);
nor U11005 (N_11005,N_10527,N_10389);
nand U11006 (N_11006,N_10176,N_10149);
or U11007 (N_11007,N_10618,N_10361);
and U11008 (N_11008,N_10000,N_10337);
xor U11009 (N_11009,N_10463,N_10135);
and U11010 (N_11010,N_10044,N_10479);
or U11011 (N_11011,N_10199,N_10022);
xnor U11012 (N_11012,N_10222,N_10391);
or U11013 (N_11013,N_10464,N_10123);
or U11014 (N_11014,N_10544,N_10372);
or U11015 (N_11015,N_10085,N_10135);
nor U11016 (N_11016,N_10424,N_10475);
or U11017 (N_11017,N_10498,N_10501);
or U11018 (N_11018,N_10051,N_10322);
and U11019 (N_11019,N_10557,N_10018);
xnor U11020 (N_11020,N_10419,N_10498);
nand U11021 (N_11021,N_10571,N_10392);
xnor U11022 (N_11022,N_10296,N_10563);
and U11023 (N_11023,N_10342,N_10231);
and U11024 (N_11024,N_10585,N_10608);
or U11025 (N_11025,N_10308,N_10083);
xnor U11026 (N_11026,N_10331,N_10562);
nand U11027 (N_11027,N_10195,N_10279);
nor U11028 (N_11028,N_10274,N_10251);
nor U11029 (N_11029,N_10030,N_10323);
or U11030 (N_11030,N_10358,N_10621);
or U11031 (N_11031,N_10574,N_10175);
and U11032 (N_11032,N_10358,N_10078);
nand U11033 (N_11033,N_10027,N_10019);
nor U11034 (N_11034,N_10373,N_10526);
nor U11035 (N_11035,N_10403,N_10231);
nand U11036 (N_11036,N_10061,N_10582);
or U11037 (N_11037,N_10071,N_10242);
nand U11038 (N_11038,N_10015,N_10238);
and U11039 (N_11039,N_10173,N_10193);
nor U11040 (N_11040,N_10534,N_10603);
nand U11041 (N_11041,N_10391,N_10102);
xor U11042 (N_11042,N_10532,N_10359);
and U11043 (N_11043,N_10311,N_10476);
xor U11044 (N_11044,N_10030,N_10306);
nand U11045 (N_11045,N_10355,N_10443);
xor U11046 (N_11046,N_10383,N_10374);
xor U11047 (N_11047,N_10496,N_10423);
or U11048 (N_11048,N_10381,N_10505);
nor U11049 (N_11049,N_10110,N_10484);
and U11050 (N_11050,N_10267,N_10450);
xnor U11051 (N_11051,N_10572,N_10167);
nand U11052 (N_11052,N_10259,N_10509);
nand U11053 (N_11053,N_10039,N_10076);
nor U11054 (N_11054,N_10120,N_10335);
or U11055 (N_11055,N_10071,N_10000);
nor U11056 (N_11056,N_10240,N_10169);
and U11057 (N_11057,N_10374,N_10099);
and U11058 (N_11058,N_10219,N_10471);
xor U11059 (N_11059,N_10141,N_10525);
and U11060 (N_11060,N_10611,N_10510);
and U11061 (N_11061,N_10516,N_10066);
and U11062 (N_11062,N_10573,N_10532);
nor U11063 (N_11063,N_10606,N_10014);
xor U11064 (N_11064,N_10356,N_10529);
xnor U11065 (N_11065,N_10196,N_10197);
and U11066 (N_11066,N_10282,N_10373);
xor U11067 (N_11067,N_10210,N_10003);
and U11068 (N_11068,N_10469,N_10123);
xnor U11069 (N_11069,N_10344,N_10099);
nor U11070 (N_11070,N_10552,N_10407);
xor U11071 (N_11071,N_10529,N_10176);
or U11072 (N_11072,N_10274,N_10120);
or U11073 (N_11073,N_10588,N_10119);
or U11074 (N_11074,N_10413,N_10576);
nor U11075 (N_11075,N_10139,N_10273);
or U11076 (N_11076,N_10166,N_10518);
and U11077 (N_11077,N_10449,N_10419);
nor U11078 (N_11078,N_10334,N_10109);
xor U11079 (N_11079,N_10582,N_10470);
nand U11080 (N_11080,N_10116,N_10372);
nor U11081 (N_11081,N_10087,N_10352);
xor U11082 (N_11082,N_10266,N_10567);
and U11083 (N_11083,N_10002,N_10048);
nor U11084 (N_11084,N_10177,N_10066);
nand U11085 (N_11085,N_10333,N_10409);
nand U11086 (N_11086,N_10575,N_10201);
nand U11087 (N_11087,N_10312,N_10115);
xor U11088 (N_11088,N_10170,N_10087);
nor U11089 (N_11089,N_10409,N_10506);
and U11090 (N_11090,N_10575,N_10047);
nand U11091 (N_11091,N_10245,N_10124);
xor U11092 (N_11092,N_10243,N_10378);
nand U11093 (N_11093,N_10413,N_10551);
nor U11094 (N_11094,N_10247,N_10162);
and U11095 (N_11095,N_10186,N_10537);
and U11096 (N_11096,N_10551,N_10396);
xnor U11097 (N_11097,N_10277,N_10328);
xnor U11098 (N_11098,N_10265,N_10050);
nand U11099 (N_11099,N_10400,N_10559);
xor U11100 (N_11100,N_10617,N_10453);
nand U11101 (N_11101,N_10367,N_10033);
xor U11102 (N_11102,N_10082,N_10518);
nand U11103 (N_11103,N_10323,N_10131);
and U11104 (N_11104,N_10366,N_10463);
or U11105 (N_11105,N_10401,N_10365);
or U11106 (N_11106,N_10349,N_10497);
and U11107 (N_11107,N_10070,N_10375);
or U11108 (N_11108,N_10331,N_10279);
and U11109 (N_11109,N_10179,N_10143);
xor U11110 (N_11110,N_10514,N_10370);
nor U11111 (N_11111,N_10143,N_10359);
nor U11112 (N_11112,N_10167,N_10563);
or U11113 (N_11113,N_10418,N_10317);
xnor U11114 (N_11114,N_10250,N_10237);
nor U11115 (N_11115,N_10582,N_10446);
and U11116 (N_11116,N_10091,N_10290);
nand U11117 (N_11117,N_10521,N_10477);
nor U11118 (N_11118,N_10162,N_10084);
nand U11119 (N_11119,N_10549,N_10286);
nor U11120 (N_11120,N_10218,N_10240);
nand U11121 (N_11121,N_10440,N_10355);
xor U11122 (N_11122,N_10083,N_10330);
or U11123 (N_11123,N_10607,N_10187);
nand U11124 (N_11124,N_10395,N_10212);
nor U11125 (N_11125,N_10518,N_10431);
and U11126 (N_11126,N_10317,N_10354);
xnor U11127 (N_11127,N_10206,N_10611);
nor U11128 (N_11128,N_10127,N_10383);
nor U11129 (N_11129,N_10101,N_10057);
or U11130 (N_11130,N_10162,N_10068);
or U11131 (N_11131,N_10253,N_10128);
nor U11132 (N_11132,N_10623,N_10345);
xor U11133 (N_11133,N_10268,N_10210);
nand U11134 (N_11134,N_10329,N_10073);
nor U11135 (N_11135,N_10591,N_10523);
and U11136 (N_11136,N_10048,N_10428);
and U11137 (N_11137,N_10356,N_10313);
and U11138 (N_11138,N_10233,N_10544);
and U11139 (N_11139,N_10347,N_10196);
xor U11140 (N_11140,N_10083,N_10168);
xnor U11141 (N_11141,N_10092,N_10183);
xor U11142 (N_11142,N_10181,N_10269);
and U11143 (N_11143,N_10491,N_10356);
and U11144 (N_11144,N_10137,N_10024);
and U11145 (N_11145,N_10101,N_10530);
nand U11146 (N_11146,N_10469,N_10543);
or U11147 (N_11147,N_10545,N_10247);
nand U11148 (N_11148,N_10424,N_10385);
or U11149 (N_11149,N_10409,N_10028);
xor U11150 (N_11150,N_10481,N_10316);
and U11151 (N_11151,N_10519,N_10567);
and U11152 (N_11152,N_10591,N_10621);
or U11153 (N_11153,N_10614,N_10451);
nand U11154 (N_11154,N_10219,N_10399);
or U11155 (N_11155,N_10332,N_10250);
nor U11156 (N_11156,N_10540,N_10579);
or U11157 (N_11157,N_10074,N_10176);
xor U11158 (N_11158,N_10074,N_10542);
xnor U11159 (N_11159,N_10349,N_10449);
nor U11160 (N_11160,N_10056,N_10104);
and U11161 (N_11161,N_10602,N_10532);
nor U11162 (N_11162,N_10325,N_10424);
nor U11163 (N_11163,N_10277,N_10187);
xor U11164 (N_11164,N_10208,N_10621);
xor U11165 (N_11165,N_10413,N_10143);
and U11166 (N_11166,N_10097,N_10000);
nand U11167 (N_11167,N_10437,N_10529);
or U11168 (N_11168,N_10619,N_10518);
xor U11169 (N_11169,N_10465,N_10199);
xor U11170 (N_11170,N_10245,N_10597);
and U11171 (N_11171,N_10447,N_10298);
nor U11172 (N_11172,N_10309,N_10145);
and U11173 (N_11173,N_10604,N_10480);
nand U11174 (N_11174,N_10549,N_10217);
xor U11175 (N_11175,N_10254,N_10317);
and U11176 (N_11176,N_10088,N_10383);
and U11177 (N_11177,N_10447,N_10605);
nand U11178 (N_11178,N_10306,N_10511);
and U11179 (N_11179,N_10455,N_10212);
xnor U11180 (N_11180,N_10508,N_10339);
xor U11181 (N_11181,N_10488,N_10196);
nand U11182 (N_11182,N_10473,N_10268);
and U11183 (N_11183,N_10305,N_10476);
nor U11184 (N_11184,N_10303,N_10255);
nand U11185 (N_11185,N_10303,N_10364);
and U11186 (N_11186,N_10081,N_10153);
nand U11187 (N_11187,N_10439,N_10097);
nor U11188 (N_11188,N_10134,N_10305);
xnor U11189 (N_11189,N_10532,N_10154);
xnor U11190 (N_11190,N_10203,N_10210);
or U11191 (N_11191,N_10598,N_10365);
and U11192 (N_11192,N_10015,N_10080);
nand U11193 (N_11193,N_10621,N_10276);
or U11194 (N_11194,N_10352,N_10586);
xor U11195 (N_11195,N_10415,N_10314);
and U11196 (N_11196,N_10023,N_10194);
nand U11197 (N_11197,N_10476,N_10068);
nand U11198 (N_11198,N_10186,N_10519);
and U11199 (N_11199,N_10050,N_10222);
xnor U11200 (N_11200,N_10338,N_10055);
nand U11201 (N_11201,N_10010,N_10330);
and U11202 (N_11202,N_10561,N_10461);
nor U11203 (N_11203,N_10406,N_10145);
xor U11204 (N_11204,N_10357,N_10365);
nand U11205 (N_11205,N_10439,N_10184);
or U11206 (N_11206,N_10326,N_10054);
and U11207 (N_11207,N_10602,N_10530);
nand U11208 (N_11208,N_10517,N_10051);
or U11209 (N_11209,N_10332,N_10198);
and U11210 (N_11210,N_10100,N_10163);
xnor U11211 (N_11211,N_10236,N_10177);
and U11212 (N_11212,N_10429,N_10307);
nor U11213 (N_11213,N_10350,N_10278);
nor U11214 (N_11214,N_10347,N_10497);
or U11215 (N_11215,N_10579,N_10523);
or U11216 (N_11216,N_10514,N_10473);
and U11217 (N_11217,N_10203,N_10372);
nor U11218 (N_11218,N_10176,N_10416);
or U11219 (N_11219,N_10171,N_10614);
or U11220 (N_11220,N_10419,N_10128);
nor U11221 (N_11221,N_10238,N_10380);
nor U11222 (N_11222,N_10615,N_10416);
nor U11223 (N_11223,N_10179,N_10019);
xor U11224 (N_11224,N_10374,N_10586);
or U11225 (N_11225,N_10136,N_10537);
or U11226 (N_11226,N_10581,N_10178);
or U11227 (N_11227,N_10366,N_10018);
xor U11228 (N_11228,N_10275,N_10338);
nor U11229 (N_11229,N_10268,N_10495);
nor U11230 (N_11230,N_10237,N_10383);
nand U11231 (N_11231,N_10016,N_10290);
or U11232 (N_11232,N_10269,N_10502);
nor U11233 (N_11233,N_10099,N_10316);
or U11234 (N_11234,N_10213,N_10138);
nand U11235 (N_11235,N_10573,N_10109);
nor U11236 (N_11236,N_10218,N_10152);
nand U11237 (N_11237,N_10039,N_10586);
nor U11238 (N_11238,N_10219,N_10558);
nand U11239 (N_11239,N_10053,N_10085);
xnor U11240 (N_11240,N_10206,N_10338);
and U11241 (N_11241,N_10496,N_10326);
nor U11242 (N_11242,N_10429,N_10031);
and U11243 (N_11243,N_10102,N_10051);
nand U11244 (N_11244,N_10555,N_10237);
nand U11245 (N_11245,N_10022,N_10437);
xnor U11246 (N_11246,N_10455,N_10043);
nand U11247 (N_11247,N_10198,N_10278);
xor U11248 (N_11248,N_10546,N_10376);
nand U11249 (N_11249,N_10496,N_10555);
xnor U11250 (N_11250,N_11175,N_11132);
xnor U11251 (N_11251,N_11188,N_11172);
and U11252 (N_11252,N_10641,N_11189);
or U11253 (N_11253,N_10947,N_11160);
nor U11254 (N_11254,N_11021,N_10969);
xor U11255 (N_11255,N_10653,N_10640);
xnor U11256 (N_11256,N_10973,N_11112);
nor U11257 (N_11257,N_11141,N_10975);
nand U11258 (N_11258,N_11084,N_11232);
and U11259 (N_11259,N_10815,N_11098);
nor U11260 (N_11260,N_11181,N_11031);
xnor U11261 (N_11261,N_11209,N_11137);
and U11262 (N_11262,N_11065,N_11004);
or U11263 (N_11263,N_11022,N_10883);
and U11264 (N_11264,N_10962,N_10761);
nand U11265 (N_11265,N_11239,N_11122);
nor U11266 (N_11266,N_10944,N_10771);
nand U11267 (N_11267,N_10943,N_10999);
or U11268 (N_11268,N_11086,N_11238);
nand U11269 (N_11269,N_10749,N_10825);
and U11270 (N_11270,N_10680,N_10797);
or U11271 (N_11271,N_11087,N_11214);
xnor U11272 (N_11272,N_11040,N_11143);
nand U11273 (N_11273,N_10778,N_11201);
nand U11274 (N_11274,N_10991,N_10723);
nand U11275 (N_11275,N_10908,N_10632);
nand U11276 (N_11276,N_10775,N_10644);
nor U11277 (N_11277,N_10781,N_11124);
xnor U11278 (N_11278,N_10869,N_10732);
nand U11279 (N_11279,N_10626,N_11186);
nand U11280 (N_11280,N_10746,N_10774);
nand U11281 (N_11281,N_11231,N_10839);
or U11282 (N_11282,N_10966,N_11217);
nor U11283 (N_11283,N_10655,N_11013);
or U11284 (N_11284,N_11035,N_10683);
nand U11285 (N_11285,N_11233,N_10638);
or U11286 (N_11286,N_11116,N_11042);
nor U11287 (N_11287,N_11223,N_10634);
and U11288 (N_11288,N_11166,N_11151);
nor U11289 (N_11289,N_10990,N_10919);
or U11290 (N_11290,N_10950,N_10836);
or U11291 (N_11291,N_10851,N_11082);
nand U11292 (N_11292,N_11154,N_10870);
nand U11293 (N_11293,N_10901,N_10806);
xnor U11294 (N_11294,N_10629,N_10691);
nand U11295 (N_11295,N_11121,N_10789);
xnor U11296 (N_11296,N_11144,N_10956);
nor U11297 (N_11297,N_11003,N_10730);
nand U11298 (N_11298,N_10959,N_10736);
or U11299 (N_11299,N_10881,N_11218);
or U11300 (N_11300,N_10960,N_10935);
and U11301 (N_11301,N_10756,N_11049);
nor U11302 (N_11302,N_10809,N_10831);
nand U11303 (N_11303,N_11044,N_10742);
and U11304 (N_11304,N_11246,N_10646);
nand U11305 (N_11305,N_10793,N_10660);
or U11306 (N_11306,N_11227,N_10647);
or U11307 (N_11307,N_10910,N_11178);
or U11308 (N_11308,N_10829,N_10695);
nand U11309 (N_11309,N_10710,N_11016);
nor U11310 (N_11310,N_11046,N_10738);
xnor U11311 (N_11311,N_10874,N_10783);
or U11312 (N_11312,N_10631,N_10984);
or U11313 (N_11313,N_10740,N_10992);
nand U11314 (N_11314,N_11200,N_11052);
nand U11315 (N_11315,N_11133,N_11105);
or U11316 (N_11316,N_10859,N_10835);
and U11317 (N_11317,N_10843,N_10721);
or U11318 (N_11318,N_10711,N_10807);
xor U11319 (N_11319,N_10639,N_10968);
nor U11320 (N_11320,N_11029,N_10997);
nand U11321 (N_11321,N_10860,N_10864);
nand U11322 (N_11322,N_11208,N_10800);
nor U11323 (N_11323,N_11069,N_10817);
nor U11324 (N_11324,N_11169,N_11017);
or U11325 (N_11325,N_11102,N_11094);
xor U11326 (N_11326,N_10987,N_10755);
xor U11327 (N_11327,N_11131,N_10924);
xor U11328 (N_11328,N_11176,N_10834);
xor U11329 (N_11329,N_10718,N_10934);
and U11330 (N_11330,N_11006,N_10830);
or U11331 (N_11331,N_11005,N_10914);
nor U11332 (N_11332,N_10767,N_10709);
nor U11333 (N_11333,N_10678,N_11202);
nor U11334 (N_11334,N_10694,N_11236);
nor U11335 (N_11335,N_11047,N_10798);
nand U11336 (N_11336,N_11015,N_10760);
or U11337 (N_11337,N_10823,N_10844);
nand U11338 (N_11338,N_10982,N_11184);
or U11339 (N_11339,N_10974,N_10887);
nor U11340 (N_11340,N_10878,N_11114);
or U11341 (N_11341,N_11010,N_11159);
nor U11342 (N_11342,N_11039,N_10762);
nand U11343 (N_11343,N_11030,N_10895);
nand U11344 (N_11344,N_10983,N_10790);
xnor U11345 (N_11345,N_10970,N_10673);
nor U11346 (N_11346,N_10648,N_10805);
xnor U11347 (N_11347,N_10770,N_10977);
or U11348 (N_11348,N_10784,N_10656);
or U11349 (N_11349,N_10957,N_10666);
nand U11350 (N_11350,N_11061,N_10757);
or U11351 (N_11351,N_10929,N_11092);
and U11352 (N_11352,N_10669,N_10667);
or U11353 (N_11353,N_11228,N_10759);
nand U11354 (N_11354,N_10838,N_11135);
xnor U11355 (N_11355,N_10722,N_10628);
nand U11356 (N_11356,N_10980,N_10681);
and U11357 (N_11357,N_11157,N_11148);
and U11358 (N_11358,N_10802,N_10668);
or U11359 (N_11359,N_11206,N_10854);
nor U11360 (N_11360,N_11070,N_11099);
nand U11361 (N_11361,N_10703,N_11075);
nor U11362 (N_11362,N_10720,N_10677);
or U11363 (N_11363,N_10689,N_10692);
or U11364 (N_11364,N_11090,N_11230);
nand U11365 (N_11365,N_11113,N_10922);
xor U11366 (N_11366,N_11054,N_10712);
or U11367 (N_11367,N_11242,N_11192);
nand U11368 (N_11368,N_11180,N_10735);
nand U11369 (N_11369,N_10855,N_10727);
and U11370 (N_11370,N_10985,N_11191);
and U11371 (N_11371,N_10650,N_11025);
nor U11372 (N_11372,N_11018,N_11179);
xnor U11373 (N_11373,N_10857,N_10989);
and U11374 (N_11374,N_10937,N_10779);
nand U11375 (N_11375,N_10745,N_10821);
xnor U11376 (N_11376,N_11243,N_11038);
and U11377 (N_11377,N_10981,N_10911);
nand U11378 (N_11378,N_10785,N_10662);
nor U11379 (N_11379,N_10682,N_10765);
and U11380 (N_11380,N_10876,N_10946);
nor U11381 (N_11381,N_11118,N_10868);
xor U11382 (N_11382,N_10717,N_11109);
nand U11383 (N_11383,N_10896,N_11168);
nand U11384 (N_11384,N_10842,N_10953);
or U11385 (N_11385,N_10875,N_11211);
or U11386 (N_11386,N_10900,N_10636);
xor U11387 (N_11387,N_10769,N_10810);
or U11388 (N_11388,N_11150,N_11164);
xnor U11389 (N_11389,N_11080,N_10951);
and U11390 (N_11390,N_11119,N_11177);
or U11391 (N_11391,N_10766,N_11245);
xor U11392 (N_11392,N_11207,N_10697);
nand U11393 (N_11393,N_11055,N_11123);
nand U11394 (N_11394,N_10884,N_10867);
and U11395 (N_11395,N_11183,N_10933);
xor U11396 (N_11396,N_10816,N_11111);
nand U11397 (N_11397,N_10863,N_10643);
nand U11398 (N_11398,N_10812,N_10897);
nand U11399 (N_11399,N_11012,N_10993);
nor U11400 (N_11400,N_10871,N_10845);
or U11401 (N_11401,N_10941,N_10702);
or U11402 (N_11402,N_10915,N_10688);
xnor U11403 (N_11403,N_11063,N_11064);
nand U11404 (N_11404,N_10903,N_11174);
xor U11405 (N_11405,N_10995,N_10671);
xnor U11406 (N_11406,N_10724,N_11117);
nand U11407 (N_11407,N_11210,N_10964);
nand U11408 (N_11408,N_10741,N_10729);
and U11409 (N_11409,N_11036,N_10967);
xnor U11410 (N_11410,N_10872,N_10719);
xnor U11411 (N_11411,N_11222,N_11002);
nand U11412 (N_11412,N_10961,N_11104);
or U11413 (N_11413,N_11107,N_10936);
xnor U11414 (N_11414,N_10913,N_11156);
and U11415 (N_11415,N_10909,N_10885);
xnor U11416 (N_11416,N_11163,N_10866);
xor U11417 (N_11417,N_10856,N_10725);
and U11418 (N_11418,N_11028,N_10891);
or U11419 (N_11419,N_11126,N_10700);
nand U11420 (N_11420,N_10888,N_10906);
nand U11421 (N_11421,N_10728,N_10748);
xnor U11422 (N_11422,N_10803,N_10898);
xnor U11423 (N_11423,N_11155,N_11045);
and U11424 (N_11424,N_10926,N_11173);
or U11425 (N_11425,N_11101,N_10776);
nor U11426 (N_11426,N_10925,N_10786);
nand U11427 (N_11427,N_11129,N_10998);
nand U11428 (N_11428,N_10690,N_10832);
and U11429 (N_11429,N_10743,N_10826);
and U11430 (N_11430,N_11139,N_10706);
and U11431 (N_11431,N_10813,N_10963);
and U11432 (N_11432,N_10696,N_11062);
xor U11433 (N_11433,N_10847,N_10679);
nor U11434 (N_11434,N_11023,N_11158);
or U11435 (N_11435,N_10750,N_11162);
or U11436 (N_11436,N_11234,N_11091);
xnor U11437 (N_11437,N_11056,N_11127);
and U11438 (N_11438,N_11165,N_11068);
and U11439 (N_11439,N_11224,N_10972);
nor U11440 (N_11440,N_10685,N_10971);
nand U11441 (N_11441,N_11130,N_10945);
or U11442 (N_11442,N_10822,N_10658);
xor U11443 (N_11443,N_10905,N_10930);
or U11444 (N_11444,N_11134,N_10958);
nand U11445 (N_11445,N_11235,N_10733);
xnor U11446 (N_11446,N_11247,N_11226);
nor U11447 (N_11447,N_11215,N_10955);
nor U11448 (N_11448,N_11203,N_10726);
xor U11449 (N_11449,N_11145,N_10704);
or U11450 (N_11450,N_10670,N_11220);
or U11451 (N_11451,N_10853,N_10996);
and U11452 (N_11452,N_10894,N_11198);
nand U11453 (N_11453,N_11152,N_10799);
or U11454 (N_11454,N_10652,N_10976);
nand U11455 (N_11455,N_10986,N_11147);
or U11456 (N_11456,N_11050,N_10751);
or U11457 (N_11457,N_10753,N_11237);
xor U11458 (N_11458,N_10848,N_10841);
and U11459 (N_11459,N_10828,N_10676);
or U11460 (N_11460,N_10931,N_11219);
nor U11461 (N_11461,N_11033,N_11193);
or U11462 (N_11462,N_10824,N_10877);
and U11463 (N_11463,N_11019,N_10674);
or U11464 (N_11464,N_10782,N_11161);
or U11465 (N_11465,N_10928,N_10837);
nand U11466 (N_11466,N_10890,N_11043);
xnor U11467 (N_11467,N_10893,N_11110);
nand U11468 (N_11468,N_10664,N_10788);
and U11469 (N_11469,N_11059,N_10633);
or U11470 (N_11470,N_10715,N_11108);
and U11471 (N_11471,N_10818,N_11205);
nand U11472 (N_11472,N_10965,N_10949);
and U11473 (N_11473,N_11244,N_11120);
and U11474 (N_11474,N_10792,N_10820);
nand U11475 (N_11475,N_11057,N_10846);
nand U11476 (N_11476,N_11204,N_10791);
nand U11477 (N_11477,N_10850,N_10713);
and U11478 (N_11478,N_11053,N_10747);
nor U11479 (N_11479,N_10952,N_10659);
nor U11480 (N_11480,N_10708,N_10737);
and U11481 (N_11481,N_11027,N_10739);
and U11482 (N_11482,N_10892,N_11249);
and U11483 (N_11483,N_11195,N_10651);
and U11484 (N_11484,N_10663,N_11149);
xor U11485 (N_11485,N_11194,N_10627);
nand U11486 (N_11486,N_11100,N_10804);
and U11487 (N_11487,N_10777,N_11066);
xor U11488 (N_11488,N_11115,N_10787);
nor U11489 (N_11489,N_11196,N_10714);
and U11490 (N_11490,N_10716,N_11095);
nor U11491 (N_11491,N_10862,N_11128);
xor U11492 (N_11492,N_10904,N_11071);
or U11493 (N_11493,N_11081,N_11026);
nor U11494 (N_11494,N_11140,N_10827);
and U11495 (N_11495,N_10923,N_10882);
nor U11496 (N_11496,N_11001,N_11197);
nand U11497 (N_11497,N_10907,N_10686);
xor U11498 (N_11498,N_10918,N_10625);
or U11499 (N_11499,N_10858,N_11007);
nand U11500 (N_11500,N_10795,N_10927);
nor U11501 (N_11501,N_11009,N_10879);
or U11502 (N_11502,N_10796,N_11020);
nand U11503 (N_11503,N_11138,N_11058);
and U11504 (N_11504,N_11088,N_10661);
or U11505 (N_11505,N_11212,N_10773);
and U11506 (N_11506,N_11248,N_11032);
xnor U11507 (N_11507,N_10917,N_11067);
xor U11508 (N_11508,N_10978,N_11125);
or U11509 (N_11509,N_10657,N_11034);
or U11510 (N_11510,N_11216,N_11079);
nor U11511 (N_11511,N_10654,N_10701);
nand U11512 (N_11512,N_11011,N_10988);
xor U11513 (N_11513,N_10687,N_10649);
nand U11514 (N_11514,N_11083,N_11089);
or U11515 (N_11515,N_11146,N_11170);
or U11516 (N_11516,N_10705,N_10635);
and U11517 (N_11517,N_11213,N_10840);
nand U11518 (N_11518,N_10794,N_10642);
nor U11519 (N_11519,N_10675,N_11225);
nand U11520 (N_11520,N_10880,N_10852);
nor U11521 (N_11521,N_10698,N_11190);
nor U11522 (N_11522,N_10684,N_11153);
nor U11523 (N_11523,N_10693,N_11097);
nor U11524 (N_11524,N_11037,N_10912);
nor U11525 (N_11525,N_10932,N_10754);
nor U11526 (N_11526,N_11187,N_10630);
nand U11527 (N_11527,N_11048,N_10899);
nor U11528 (N_11528,N_10731,N_11008);
nand U11529 (N_11529,N_10758,N_10744);
xnor U11530 (N_11530,N_10886,N_11077);
or U11531 (N_11531,N_11072,N_11093);
or U11532 (N_11532,N_11024,N_10921);
and U11533 (N_11533,N_10994,N_10699);
and U11534 (N_11534,N_11060,N_10920);
nor U11535 (N_11535,N_11041,N_10889);
and U11536 (N_11536,N_11076,N_10811);
nor U11537 (N_11537,N_10801,N_10849);
xnor U11538 (N_11538,N_11106,N_10954);
nand U11539 (N_11539,N_10752,N_10764);
xnor U11540 (N_11540,N_11103,N_10707);
xor U11541 (N_11541,N_10763,N_11229);
nand U11542 (N_11542,N_11171,N_10772);
nor U11543 (N_11543,N_11085,N_10861);
xnor U11544 (N_11544,N_10819,N_10808);
and U11545 (N_11545,N_11014,N_10939);
xor U11546 (N_11546,N_10948,N_11185);
nand U11547 (N_11547,N_10873,N_10665);
or U11548 (N_11548,N_10768,N_11096);
nand U11549 (N_11549,N_10916,N_10672);
nor U11550 (N_11550,N_10780,N_10979);
or U11551 (N_11551,N_10940,N_10645);
xor U11552 (N_11552,N_11000,N_11078);
nor U11553 (N_11553,N_11051,N_11142);
or U11554 (N_11554,N_11240,N_11221);
and U11555 (N_11555,N_10865,N_10938);
nor U11556 (N_11556,N_10637,N_11241);
nand U11557 (N_11557,N_10734,N_10833);
nand U11558 (N_11558,N_11073,N_11136);
nand U11559 (N_11559,N_10942,N_10902);
xor U11560 (N_11560,N_11199,N_11074);
xnor U11561 (N_11561,N_11182,N_10814);
nor U11562 (N_11562,N_11167,N_10956);
nand U11563 (N_11563,N_11128,N_11056);
nor U11564 (N_11564,N_10702,N_11054);
and U11565 (N_11565,N_11037,N_10631);
nor U11566 (N_11566,N_10807,N_10901);
or U11567 (N_11567,N_10769,N_10871);
nor U11568 (N_11568,N_10731,N_11218);
nand U11569 (N_11569,N_10655,N_10901);
xnor U11570 (N_11570,N_10733,N_11218);
or U11571 (N_11571,N_10723,N_10992);
nor U11572 (N_11572,N_10890,N_10960);
and U11573 (N_11573,N_11053,N_11092);
nor U11574 (N_11574,N_10811,N_10863);
nand U11575 (N_11575,N_11190,N_11006);
and U11576 (N_11576,N_11182,N_11242);
or U11577 (N_11577,N_11059,N_11206);
xnor U11578 (N_11578,N_10800,N_10888);
nor U11579 (N_11579,N_11076,N_10886);
xnor U11580 (N_11580,N_11171,N_11097);
nor U11581 (N_11581,N_10917,N_10925);
or U11582 (N_11582,N_10708,N_10735);
nand U11583 (N_11583,N_11220,N_10785);
and U11584 (N_11584,N_11098,N_11121);
or U11585 (N_11585,N_11200,N_10843);
nor U11586 (N_11586,N_11097,N_10944);
nand U11587 (N_11587,N_10825,N_10634);
nor U11588 (N_11588,N_11238,N_11200);
nor U11589 (N_11589,N_11115,N_10688);
nand U11590 (N_11590,N_11215,N_11031);
nor U11591 (N_11591,N_10890,N_10917);
xor U11592 (N_11592,N_10987,N_11199);
nand U11593 (N_11593,N_10709,N_10919);
and U11594 (N_11594,N_10944,N_10762);
or U11595 (N_11595,N_10930,N_10950);
and U11596 (N_11596,N_10881,N_10791);
and U11597 (N_11597,N_11152,N_10822);
xnor U11598 (N_11598,N_10820,N_11038);
or U11599 (N_11599,N_11244,N_10912);
nand U11600 (N_11600,N_10745,N_10913);
xnor U11601 (N_11601,N_10937,N_10829);
nand U11602 (N_11602,N_11025,N_10701);
xor U11603 (N_11603,N_11208,N_11010);
xnor U11604 (N_11604,N_11248,N_11200);
and U11605 (N_11605,N_10724,N_11047);
nand U11606 (N_11606,N_10851,N_11240);
xor U11607 (N_11607,N_11210,N_10998);
xnor U11608 (N_11608,N_10677,N_10674);
xnor U11609 (N_11609,N_10988,N_11145);
nor U11610 (N_11610,N_11157,N_11115);
xor U11611 (N_11611,N_10990,N_10793);
nand U11612 (N_11612,N_11051,N_11132);
nor U11613 (N_11613,N_10901,N_11225);
nand U11614 (N_11614,N_11166,N_11135);
and U11615 (N_11615,N_11141,N_10629);
xnor U11616 (N_11616,N_11187,N_11183);
nor U11617 (N_11617,N_10852,N_10865);
nand U11618 (N_11618,N_10739,N_11121);
or U11619 (N_11619,N_10728,N_11219);
nand U11620 (N_11620,N_11077,N_10629);
and U11621 (N_11621,N_10803,N_10987);
or U11622 (N_11622,N_10821,N_11007);
xnor U11623 (N_11623,N_10976,N_11120);
or U11624 (N_11624,N_10951,N_11064);
xor U11625 (N_11625,N_11043,N_11133);
xor U11626 (N_11626,N_11227,N_10812);
nor U11627 (N_11627,N_10832,N_10850);
and U11628 (N_11628,N_11134,N_10816);
xnor U11629 (N_11629,N_11082,N_10803);
and U11630 (N_11630,N_11169,N_11116);
nor U11631 (N_11631,N_10907,N_11016);
or U11632 (N_11632,N_11213,N_10822);
nand U11633 (N_11633,N_10764,N_10920);
nand U11634 (N_11634,N_11080,N_11021);
xor U11635 (N_11635,N_10646,N_11239);
nand U11636 (N_11636,N_10714,N_11045);
and U11637 (N_11637,N_11105,N_10892);
nand U11638 (N_11638,N_10923,N_11036);
nor U11639 (N_11639,N_10886,N_11135);
nor U11640 (N_11640,N_10967,N_11066);
xnor U11641 (N_11641,N_10792,N_10905);
nand U11642 (N_11642,N_10753,N_11151);
nand U11643 (N_11643,N_10702,N_10746);
nand U11644 (N_11644,N_10873,N_10907);
nand U11645 (N_11645,N_10957,N_10719);
nand U11646 (N_11646,N_10976,N_10874);
or U11647 (N_11647,N_11181,N_10926);
nor U11648 (N_11648,N_11206,N_10739);
nand U11649 (N_11649,N_10735,N_11111);
or U11650 (N_11650,N_11079,N_10750);
nand U11651 (N_11651,N_10803,N_10760);
and U11652 (N_11652,N_10818,N_11249);
and U11653 (N_11653,N_10808,N_10644);
and U11654 (N_11654,N_10661,N_11190);
nor U11655 (N_11655,N_11053,N_10625);
and U11656 (N_11656,N_11048,N_11184);
nor U11657 (N_11657,N_10682,N_11051);
nor U11658 (N_11658,N_10634,N_10937);
xnor U11659 (N_11659,N_10724,N_10855);
nor U11660 (N_11660,N_10698,N_10776);
and U11661 (N_11661,N_11049,N_10993);
nand U11662 (N_11662,N_10986,N_11138);
nor U11663 (N_11663,N_11094,N_11166);
xor U11664 (N_11664,N_11015,N_11081);
xnor U11665 (N_11665,N_10784,N_10964);
or U11666 (N_11666,N_10874,N_10890);
and U11667 (N_11667,N_11031,N_11052);
nand U11668 (N_11668,N_10672,N_11128);
nand U11669 (N_11669,N_10863,N_10806);
xor U11670 (N_11670,N_10955,N_10798);
and U11671 (N_11671,N_10841,N_11114);
nand U11672 (N_11672,N_11032,N_10811);
nand U11673 (N_11673,N_11162,N_11017);
or U11674 (N_11674,N_11030,N_10965);
xnor U11675 (N_11675,N_11225,N_11169);
nand U11676 (N_11676,N_11145,N_10636);
or U11677 (N_11677,N_11092,N_10676);
and U11678 (N_11678,N_10841,N_11248);
nor U11679 (N_11679,N_10997,N_10708);
or U11680 (N_11680,N_10664,N_10800);
nand U11681 (N_11681,N_10790,N_11103);
xor U11682 (N_11682,N_11243,N_11234);
nand U11683 (N_11683,N_11022,N_10816);
and U11684 (N_11684,N_11247,N_10674);
nand U11685 (N_11685,N_11147,N_10940);
xor U11686 (N_11686,N_10872,N_10942);
nor U11687 (N_11687,N_11177,N_11042);
nand U11688 (N_11688,N_10835,N_11205);
xor U11689 (N_11689,N_11183,N_10930);
xnor U11690 (N_11690,N_10905,N_11097);
and U11691 (N_11691,N_11179,N_11052);
nand U11692 (N_11692,N_10829,N_10946);
nand U11693 (N_11693,N_10684,N_10988);
and U11694 (N_11694,N_11241,N_11118);
and U11695 (N_11695,N_10868,N_10867);
and U11696 (N_11696,N_11004,N_10747);
or U11697 (N_11697,N_10912,N_10724);
nor U11698 (N_11698,N_10791,N_10866);
xor U11699 (N_11699,N_10939,N_11183);
nor U11700 (N_11700,N_11017,N_11035);
xor U11701 (N_11701,N_11200,N_11002);
nor U11702 (N_11702,N_10743,N_10849);
nand U11703 (N_11703,N_10806,N_10703);
nor U11704 (N_11704,N_11158,N_10758);
or U11705 (N_11705,N_10958,N_11220);
nor U11706 (N_11706,N_11112,N_11098);
xnor U11707 (N_11707,N_11170,N_11139);
and U11708 (N_11708,N_10651,N_11194);
xnor U11709 (N_11709,N_11164,N_10693);
or U11710 (N_11710,N_10638,N_11147);
or U11711 (N_11711,N_10672,N_10733);
nand U11712 (N_11712,N_11128,N_11133);
or U11713 (N_11713,N_10649,N_11073);
nor U11714 (N_11714,N_10845,N_11029);
xor U11715 (N_11715,N_11087,N_10917);
and U11716 (N_11716,N_11230,N_10930);
and U11717 (N_11717,N_10887,N_10909);
nand U11718 (N_11718,N_11088,N_10781);
nor U11719 (N_11719,N_11232,N_10901);
nor U11720 (N_11720,N_10650,N_10813);
or U11721 (N_11721,N_11233,N_10735);
or U11722 (N_11722,N_10783,N_11109);
and U11723 (N_11723,N_10985,N_11095);
xor U11724 (N_11724,N_10870,N_10970);
or U11725 (N_11725,N_11080,N_11172);
or U11726 (N_11726,N_10804,N_11123);
and U11727 (N_11727,N_10646,N_10867);
xnor U11728 (N_11728,N_10987,N_11054);
nand U11729 (N_11729,N_10882,N_11069);
or U11730 (N_11730,N_10950,N_10676);
nand U11731 (N_11731,N_11235,N_11020);
and U11732 (N_11732,N_11195,N_10636);
and U11733 (N_11733,N_10894,N_10939);
or U11734 (N_11734,N_11173,N_11004);
nand U11735 (N_11735,N_10909,N_11200);
xnor U11736 (N_11736,N_10943,N_10919);
nor U11737 (N_11737,N_10779,N_10644);
xnor U11738 (N_11738,N_10743,N_11162);
nor U11739 (N_11739,N_11022,N_10771);
xnor U11740 (N_11740,N_10756,N_11094);
nor U11741 (N_11741,N_10790,N_10748);
nor U11742 (N_11742,N_11199,N_10928);
nand U11743 (N_11743,N_10679,N_10835);
nor U11744 (N_11744,N_11215,N_10809);
nand U11745 (N_11745,N_11010,N_11045);
and U11746 (N_11746,N_10995,N_11108);
nand U11747 (N_11747,N_10746,N_11214);
xor U11748 (N_11748,N_10885,N_10851);
and U11749 (N_11749,N_11132,N_11109);
nand U11750 (N_11750,N_10647,N_10758);
xor U11751 (N_11751,N_11028,N_10822);
nand U11752 (N_11752,N_10833,N_10717);
and U11753 (N_11753,N_11003,N_10734);
and U11754 (N_11754,N_10889,N_10703);
xor U11755 (N_11755,N_10746,N_11194);
or U11756 (N_11756,N_11112,N_11123);
nor U11757 (N_11757,N_10833,N_10825);
nand U11758 (N_11758,N_10891,N_11202);
nand U11759 (N_11759,N_11172,N_10897);
xnor U11760 (N_11760,N_10887,N_10627);
and U11761 (N_11761,N_10863,N_10683);
xor U11762 (N_11762,N_11129,N_11147);
nor U11763 (N_11763,N_10702,N_11068);
and U11764 (N_11764,N_10908,N_10950);
nor U11765 (N_11765,N_11174,N_10653);
and U11766 (N_11766,N_11102,N_11083);
xnor U11767 (N_11767,N_10669,N_11155);
nand U11768 (N_11768,N_10804,N_11136);
nand U11769 (N_11769,N_10810,N_10794);
or U11770 (N_11770,N_10717,N_10918);
or U11771 (N_11771,N_10732,N_11045);
or U11772 (N_11772,N_11164,N_10761);
xnor U11773 (N_11773,N_11249,N_11181);
xor U11774 (N_11774,N_10786,N_10695);
xnor U11775 (N_11775,N_11062,N_10722);
xnor U11776 (N_11776,N_10969,N_11022);
nor U11777 (N_11777,N_10667,N_11238);
xor U11778 (N_11778,N_11064,N_11062);
nand U11779 (N_11779,N_10763,N_10808);
or U11780 (N_11780,N_11218,N_10754);
and U11781 (N_11781,N_11066,N_11094);
and U11782 (N_11782,N_10859,N_11178);
or U11783 (N_11783,N_11223,N_10657);
nor U11784 (N_11784,N_11239,N_11107);
and U11785 (N_11785,N_11216,N_10689);
and U11786 (N_11786,N_10880,N_11086);
nor U11787 (N_11787,N_11207,N_11239);
nor U11788 (N_11788,N_11173,N_11169);
nand U11789 (N_11789,N_11120,N_10647);
nor U11790 (N_11790,N_10639,N_10849);
and U11791 (N_11791,N_10684,N_10810);
or U11792 (N_11792,N_11147,N_11203);
nor U11793 (N_11793,N_11104,N_10634);
nor U11794 (N_11794,N_10883,N_10970);
and U11795 (N_11795,N_10902,N_11021);
nor U11796 (N_11796,N_10917,N_11222);
xnor U11797 (N_11797,N_10950,N_10778);
nor U11798 (N_11798,N_10850,N_11146);
nand U11799 (N_11799,N_10835,N_10805);
or U11800 (N_11800,N_10927,N_10742);
and U11801 (N_11801,N_10792,N_10824);
and U11802 (N_11802,N_10970,N_10990);
and U11803 (N_11803,N_11160,N_11064);
and U11804 (N_11804,N_11201,N_11114);
nand U11805 (N_11805,N_10830,N_10802);
nor U11806 (N_11806,N_10716,N_10987);
nand U11807 (N_11807,N_10941,N_10780);
nor U11808 (N_11808,N_10680,N_10852);
and U11809 (N_11809,N_11203,N_10661);
or U11810 (N_11810,N_11005,N_10898);
nor U11811 (N_11811,N_10641,N_11077);
nor U11812 (N_11812,N_10639,N_11103);
xnor U11813 (N_11813,N_11180,N_10872);
nand U11814 (N_11814,N_10815,N_10886);
nand U11815 (N_11815,N_10986,N_11000);
or U11816 (N_11816,N_11065,N_10800);
and U11817 (N_11817,N_10696,N_10861);
xnor U11818 (N_11818,N_11053,N_11190);
or U11819 (N_11819,N_11046,N_10779);
xor U11820 (N_11820,N_10810,N_10888);
nor U11821 (N_11821,N_11115,N_11184);
and U11822 (N_11822,N_10824,N_10915);
nand U11823 (N_11823,N_11211,N_10696);
or U11824 (N_11824,N_11027,N_10899);
or U11825 (N_11825,N_11099,N_10833);
xor U11826 (N_11826,N_11143,N_11230);
nor U11827 (N_11827,N_10902,N_11079);
nand U11828 (N_11828,N_11103,N_10889);
nand U11829 (N_11829,N_11131,N_10792);
nand U11830 (N_11830,N_11072,N_10774);
xor U11831 (N_11831,N_10820,N_10797);
and U11832 (N_11832,N_10837,N_11012);
and U11833 (N_11833,N_11225,N_11239);
nand U11834 (N_11834,N_11054,N_11001);
nor U11835 (N_11835,N_11115,N_11113);
nand U11836 (N_11836,N_10696,N_11213);
xor U11837 (N_11837,N_11249,N_10766);
nor U11838 (N_11838,N_11123,N_11108);
nand U11839 (N_11839,N_10670,N_11154);
xnor U11840 (N_11840,N_10705,N_11051);
xor U11841 (N_11841,N_10659,N_11247);
and U11842 (N_11842,N_10809,N_11213);
or U11843 (N_11843,N_10639,N_10796);
nor U11844 (N_11844,N_11227,N_11147);
and U11845 (N_11845,N_10637,N_10671);
xor U11846 (N_11846,N_11132,N_10626);
nor U11847 (N_11847,N_10763,N_10737);
nor U11848 (N_11848,N_10697,N_10948);
or U11849 (N_11849,N_10667,N_11181);
or U11850 (N_11850,N_11148,N_10704);
or U11851 (N_11851,N_11045,N_11077);
nand U11852 (N_11852,N_10894,N_11029);
and U11853 (N_11853,N_10713,N_10652);
or U11854 (N_11854,N_10751,N_10917);
and U11855 (N_11855,N_11239,N_10742);
xor U11856 (N_11856,N_10884,N_11022);
and U11857 (N_11857,N_10936,N_10867);
and U11858 (N_11858,N_11141,N_11093);
or U11859 (N_11859,N_10929,N_11167);
nor U11860 (N_11860,N_10738,N_11017);
nor U11861 (N_11861,N_11233,N_10799);
or U11862 (N_11862,N_11157,N_10696);
and U11863 (N_11863,N_10725,N_10694);
xnor U11864 (N_11864,N_10850,N_10658);
xnor U11865 (N_11865,N_10875,N_10773);
nand U11866 (N_11866,N_10873,N_10949);
or U11867 (N_11867,N_10916,N_10976);
and U11868 (N_11868,N_10802,N_10873);
nor U11869 (N_11869,N_11152,N_10870);
xor U11870 (N_11870,N_10730,N_11156);
nand U11871 (N_11871,N_10712,N_10667);
or U11872 (N_11872,N_10894,N_11192);
and U11873 (N_11873,N_10888,N_10728);
nand U11874 (N_11874,N_10911,N_10900);
nand U11875 (N_11875,N_11774,N_11653);
nor U11876 (N_11876,N_11632,N_11331);
and U11877 (N_11877,N_11669,N_11451);
or U11878 (N_11878,N_11666,N_11856);
nand U11879 (N_11879,N_11701,N_11499);
and U11880 (N_11880,N_11668,N_11271);
xor U11881 (N_11881,N_11692,N_11556);
nand U11882 (N_11882,N_11438,N_11413);
nor U11883 (N_11883,N_11498,N_11627);
xor U11884 (N_11884,N_11317,N_11487);
nand U11885 (N_11885,N_11850,N_11562);
xnor U11886 (N_11886,N_11426,N_11848);
nand U11887 (N_11887,N_11332,N_11358);
or U11888 (N_11888,N_11546,N_11353);
or U11889 (N_11889,N_11571,N_11625);
nor U11890 (N_11890,N_11281,N_11691);
xor U11891 (N_11891,N_11743,N_11443);
nand U11892 (N_11892,N_11769,N_11832);
nor U11893 (N_11893,N_11650,N_11536);
or U11894 (N_11894,N_11693,N_11541);
nor U11895 (N_11895,N_11420,N_11697);
nand U11896 (N_11896,N_11570,N_11335);
and U11897 (N_11897,N_11720,N_11297);
nand U11898 (N_11898,N_11385,N_11591);
xor U11899 (N_11899,N_11865,N_11261);
nand U11900 (N_11900,N_11314,N_11767);
nand U11901 (N_11901,N_11548,N_11471);
nand U11902 (N_11902,N_11860,N_11700);
xor U11903 (N_11903,N_11847,N_11797);
or U11904 (N_11904,N_11791,N_11495);
and U11905 (N_11905,N_11586,N_11383);
nand U11906 (N_11906,N_11394,N_11783);
and U11907 (N_11907,N_11798,N_11690);
and U11908 (N_11908,N_11753,N_11581);
and U11909 (N_11909,N_11679,N_11654);
xnor U11910 (N_11910,N_11522,N_11736);
or U11911 (N_11911,N_11852,N_11544);
nand U11912 (N_11912,N_11773,N_11606);
xnor U11913 (N_11913,N_11651,N_11366);
and U11914 (N_11914,N_11369,N_11657);
nor U11915 (N_11915,N_11491,N_11806);
or U11916 (N_11916,N_11826,N_11871);
nor U11917 (N_11917,N_11766,N_11842);
xor U11918 (N_11918,N_11260,N_11592);
nand U11919 (N_11919,N_11755,N_11255);
or U11920 (N_11920,N_11685,N_11279);
nand U11921 (N_11921,N_11409,N_11702);
xnor U11922 (N_11922,N_11731,N_11275);
and U11923 (N_11923,N_11772,N_11288);
nor U11924 (N_11924,N_11602,N_11867);
or U11925 (N_11925,N_11721,N_11362);
nor U11926 (N_11926,N_11551,N_11858);
nand U11927 (N_11927,N_11628,N_11757);
nor U11928 (N_11928,N_11648,N_11728);
xor U11929 (N_11929,N_11818,N_11284);
xor U11930 (N_11930,N_11449,N_11620);
nor U11931 (N_11931,N_11518,N_11354);
nand U11932 (N_11932,N_11272,N_11251);
and U11933 (N_11933,N_11589,N_11843);
xnor U11934 (N_11934,N_11543,N_11454);
or U11935 (N_11935,N_11550,N_11419);
xor U11936 (N_11936,N_11578,N_11390);
nand U11937 (N_11937,N_11684,N_11304);
and U11938 (N_11938,N_11453,N_11500);
or U11939 (N_11939,N_11738,N_11593);
nand U11940 (N_11940,N_11294,N_11545);
xor U11941 (N_11941,N_11370,N_11457);
and U11942 (N_11942,N_11841,N_11611);
and U11943 (N_11943,N_11638,N_11286);
and U11944 (N_11944,N_11483,N_11553);
nor U11945 (N_11945,N_11373,N_11431);
xor U11946 (N_11946,N_11756,N_11801);
nand U11947 (N_11947,N_11463,N_11316);
xor U11948 (N_11948,N_11762,N_11315);
nand U11949 (N_11949,N_11482,N_11812);
or U11950 (N_11950,N_11754,N_11566);
nor U11951 (N_11951,N_11568,N_11530);
nor U11952 (N_11952,N_11792,N_11485);
and U11953 (N_11953,N_11819,N_11367);
nor U11954 (N_11954,N_11633,N_11861);
and U11955 (N_11955,N_11790,N_11557);
xnor U11956 (N_11956,N_11296,N_11706);
and U11957 (N_11957,N_11722,N_11647);
or U11958 (N_11958,N_11595,N_11799);
nor U11959 (N_11959,N_11254,N_11795);
xnor U11960 (N_11960,N_11868,N_11696);
nand U11961 (N_11961,N_11352,N_11376);
nor U11962 (N_11962,N_11382,N_11405);
xnor U11963 (N_11963,N_11282,N_11854);
or U11964 (N_11964,N_11660,N_11285);
and U11965 (N_11965,N_11273,N_11779);
xnor U11966 (N_11966,N_11310,N_11688);
nor U11967 (N_11967,N_11613,N_11555);
and U11968 (N_11968,N_11448,N_11505);
nor U11969 (N_11969,N_11302,N_11450);
nand U11970 (N_11970,N_11817,N_11857);
and U11971 (N_11971,N_11403,N_11597);
and U11972 (N_11972,N_11293,N_11547);
nand U11973 (N_11973,N_11590,N_11326);
and U11974 (N_11974,N_11308,N_11624);
xnor U11975 (N_11975,N_11765,N_11723);
xnor U11976 (N_11976,N_11838,N_11318);
nand U11977 (N_11977,N_11674,N_11612);
xor U11978 (N_11978,N_11807,N_11621);
xor U11979 (N_11979,N_11513,N_11337);
nor U11980 (N_11980,N_11733,N_11363);
and U11981 (N_11981,N_11422,N_11712);
nor U11982 (N_11982,N_11676,N_11836);
or U11983 (N_11983,N_11575,N_11710);
nand U11984 (N_11984,N_11360,N_11425);
nor U11985 (N_11985,N_11835,N_11565);
and U11986 (N_11986,N_11440,N_11444);
nor U11987 (N_11987,N_11349,N_11257);
nand U11988 (N_11988,N_11672,N_11834);
nand U11989 (N_11989,N_11325,N_11312);
or U11990 (N_11990,N_11408,N_11637);
nand U11991 (N_11991,N_11645,N_11291);
nor U11992 (N_11992,N_11262,N_11404);
xnor U11993 (N_11993,N_11782,N_11713);
nor U11994 (N_11994,N_11474,N_11564);
and U11995 (N_11995,N_11378,N_11446);
nor U11996 (N_11996,N_11516,N_11537);
nand U11997 (N_11997,N_11872,N_11377);
and U11998 (N_11998,N_11828,N_11560);
nand U11999 (N_11999,N_11705,N_11699);
xor U12000 (N_12000,N_11667,N_11748);
nand U12001 (N_12001,N_11810,N_11734);
or U12002 (N_12002,N_11531,N_11829);
nand U12003 (N_12003,N_11781,N_11504);
nand U12004 (N_12004,N_11458,N_11300);
nand U12005 (N_12005,N_11489,N_11439);
xnor U12006 (N_12006,N_11689,N_11729);
nand U12007 (N_12007,N_11533,N_11343);
nor U12008 (N_12008,N_11618,N_11269);
xnor U12009 (N_12009,N_11365,N_11601);
and U12010 (N_12010,N_11703,N_11567);
nand U12011 (N_12011,N_11608,N_11759);
xor U12012 (N_12012,N_11374,N_11777);
nor U12013 (N_12013,N_11780,N_11472);
or U12014 (N_12014,N_11649,N_11789);
xor U12015 (N_12015,N_11816,N_11421);
and U12016 (N_12016,N_11484,N_11341);
or U12017 (N_12017,N_11375,N_11423);
nand U12018 (N_12018,N_11574,N_11855);
nand U12019 (N_12019,N_11460,N_11350);
nor U12020 (N_12020,N_11686,N_11704);
nand U12021 (N_12021,N_11747,N_11481);
or U12022 (N_12022,N_11609,N_11348);
nor U12023 (N_12023,N_11724,N_11256);
xnor U12024 (N_12024,N_11815,N_11813);
and U12025 (N_12025,N_11506,N_11603);
nand U12026 (N_12026,N_11406,N_11596);
nor U12027 (N_12027,N_11735,N_11321);
xnor U12028 (N_12028,N_11739,N_11727);
and U12029 (N_12029,N_11695,N_11726);
or U12030 (N_12030,N_11267,N_11455);
or U12031 (N_12031,N_11535,N_11324);
nor U12032 (N_12032,N_11344,N_11824);
and U12033 (N_12033,N_11558,N_11322);
nor U12034 (N_12034,N_11298,N_11336);
or U12035 (N_12035,N_11418,N_11540);
and U12036 (N_12036,N_11682,N_11776);
nor U12037 (N_12037,N_11263,N_11845);
and U12038 (N_12038,N_11497,N_11496);
nand U12039 (N_12039,N_11626,N_11554);
nor U12040 (N_12040,N_11414,N_11866);
or U12041 (N_12041,N_11640,N_11561);
and U12042 (N_12042,N_11342,N_11644);
and U12043 (N_12043,N_11604,N_11831);
or U12044 (N_12044,N_11507,N_11830);
nor U12045 (N_12045,N_11741,N_11347);
nor U12046 (N_12046,N_11641,N_11587);
or U12047 (N_12047,N_11737,N_11687);
nand U12048 (N_12048,N_11796,N_11771);
and U12049 (N_12049,N_11268,N_11786);
or U12050 (N_12050,N_11465,N_11396);
and U12051 (N_12051,N_11785,N_11718);
or U12052 (N_12052,N_11614,N_11844);
or U12053 (N_12053,N_11663,N_11610);
xor U12054 (N_12054,N_11675,N_11368);
and U12055 (N_12055,N_11576,N_11313);
xor U12056 (N_12056,N_11278,N_11708);
nor U12057 (N_12057,N_11768,N_11473);
and U12058 (N_12058,N_11399,N_11673);
and U12059 (N_12059,N_11311,N_11873);
xnor U12060 (N_12060,N_11745,N_11433);
nor U12061 (N_12061,N_11664,N_11569);
and U12062 (N_12062,N_11820,N_11821);
or U12063 (N_12063,N_11508,N_11631);
and U12064 (N_12064,N_11635,N_11655);
and U12065 (N_12065,N_11351,N_11274);
nand U12066 (N_12066,N_11636,N_11289);
nand U12067 (N_12067,N_11447,N_11659);
nor U12068 (N_12068,N_11276,N_11392);
and U12069 (N_12069,N_11441,N_11870);
and U12070 (N_12070,N_11502,N_11853);
and U12071 (N_12071,N_11469,N_11400);
and U12072 (N_12072,N_11266,N_11577);
xnor U12073 (N_12073,N_11709,N_11778);
nand U12074 (N_12074,N_11599,N_11563);
and U12075 (N_12075,N_11521,N_11719);
nand U12076 (N_12076,N_11717,N_11730);
nor U12077 (N_12077,N_11520,N_11467);
xnor U12078 (N_12078,N_11805,N_11452);
nand U12079 (N_12079,N_11761,N_11386);
nand U12080 (N_12080,N_11387,N_11456);
nand U12081 (N_12081,N_11427,N_11411);
and U12082 (N_12082,N_11542,N_11580);
nor U12083 (N_12083,N_11346,N_11477);
nor U12084 (N_12084,N_11364,N_11320);
and U12085 (N_12085,N_11671,N_11760);
or U12086 (N_12086,N_11519,N_11391);
or U12087 (N_12087,N_11534,N_11490);
and U12088 (N_12088,N_11355,N_11616);
or U12089 (N_12089,N_11714,N_11598);
or U12090 (N_12090,N_11804,N_11784);
nor U12091 (N_12091,N_11379,N_11430);
xor U12092 (N_12092,N_11306,N_11680);
and U12093 (N_12093,N_11800,N_11607);
nand U12094 (N_12094,N_11814,N_11793);
nor U12095 (N_12095,N_11594,N_11512);
and U12096 (N_12096,N_11582,N_11742);
or U12097 (N_12097,N_11407,N_11840);
and U12098 (N_12098,N_11389,N_11361);
nand U12099 (N_12099,N_11359,N_11523);
or U12100 (N_12100,N_11334,N_11656);
or U12101 (N_12101,N_11333,N_11851);
and U12102 (N_12102,N_11356,N_11479);
nand U12103 (N_12103,N_11429,N_11770);
xnor U12104 (N_12104,N_11401,N_11579);
and U12105 (N_12105,N_11639,N_11573);
nand U12106 (N_12106,N_11694,N_11707);
nor U12107 (N_12107,N_11476,N_11677);
and U12108 (N_12108,N_11559,N_11827);
xor U12109 (N_12109,N_11811,N_11417);
or U12110 (N_12110,N_11524,N_11265);
xor U12111 (N_12111,N_11464,N_11652);
nand U12112 (N_12112,N_11292,N_11380);
nor U12113 (N_12113,N_11287,N_11746);
nand U12114 (N_12114,N_11301,N_11461);
xor U12115 (N_12115,N_11445,N_11340);
nand U12116 (N_12116,N_11809,N_11280);
xor U12117 (N_12117,N_11290,N_11462);
and U12118 (N_12118,N_11517,N_11357);
and U12119 (N_12119,N_11678,N_11509);
and U12120 (N_12120,N_11393,N_11309);
or U12121 (N_12121,N_11410,N_11526);
and U12122 (N_12122,N_11338,N_11750);
nor U12123 (N_12123,N_11527,N_11492);
xor U12124 (N_12124,N_11584,N_11862);
and U12125 (N_12125,N_11665,N_11511);
nor U12126 (N_12126,N_11681,N_11869);
xnor U12127 (N_12127,N_11822,N_11588);
or U12128 (N_12128,N_11528,N_11859);
nor U12129 (N_12129,N_11670,N_11823);
or U12130 (N_12130,N_11395,N_11788);
or U12131 (N_12131,N_11258,N_11758);
or U12132 (N_12132,N_11299,N_11549);
or U12133 (N_12133,N_11252,N_11615);
xnor U12134 (N_12134,N_11864,N_11794);
nor U12135 (N_12135,N_11442,N_11397);
nand U12136 (N_12136,N_11839,N_11605);
nor U12137 (N_12137,N_11643,N_11388);
and U12138 (N_12138,N_11330,N_11398);
or U12139 (N_12139,N_11833,N_11529);
and U12140 (N_12140,N_11466,N_11307);
or U12141 (N_12141,N_11539,N_11583);
nand U12142 (N_12142,N_11416,N_11328);
xor U12143 (N_12143,N_11501,N_11740);
nor U12144 (N_12144,N_11253,N_11837);
nand U12145 (N_12145,N_11323,N_11424);
xor U12146 (N_12146,N_11402,N_11488);
nand U12147 (N_12147,N_11270,N_11436);
or U12148 (N_12148,N_11849,N_11428);
nand U12149 (N_12149,N_11622,N_11259);
nor U12150 (N_12150,N_11277,N_11803);
and U12151 (N_12151,N_11658,N_11585);
and U12152 (N_12152,N_11538,N_11478);
nor U12153 (N_12153,N_11732,N_11415);
xor U12154 (N_12154,N_11480,N_11634);
nor U12155 (N_12155,N_11283,N_11874);
and U12156 (N_12156,N_11381,N_11475);
nand U12157 (N_12157,N_11305,N_11808);
nor U12158 (N_12158,N_11372,N_11763);
and U12159 (N_12159,N_11617,N_11646);
xnor U12160 (N_12160,N_11510,N_11503);
nand U12161 (N_12161,N_11327,N_11846);
nor U12162 (N_12162,N_11339,N_11752);
nor U12163 (N_12163,N_11494,N_11572);
xnor U12164 (N_12164,N_11514,N_11384);
nand U12165 (N_12165,N_11345,N_11802);
nand U12166 (N_12166,N_11532,N_11515);
or U12167 (N_12167,N_11600,N_11437);
or U12168 (N_12168,N_11764,N_11434);
xor U12169 (N_12169,N_11715,N_11459);
and U12170 (N_12170,N_11319,N_11744);
or U12171 (N_12171,N_11725,N_11825);
nor U12172 (N_12172,N_11642,N_11412);
xor U12173 (N_12173,N_11329,N_11468);
and U12174 (N_12174,N_11751,N_11432);
nand U12175 (N_12175,N_11629,N_11661);
xnor U12176 (N_12176,N_11863,N_11698);
or U12177 (N_12177,N_11371,N_11525);
and U12178 (N_12178,N_11630,N_11749);
and U12179 (N_12179,N_11683,N_11552);
or U12180 (N_12180,N_11470,N_11486);
xor U12181 (N_12181,N_11787,N_11493);
nand U12182 (N_12182,N_11303,N_11264);
or U12183 (N_12183,N_11435,N_11619);
xnor U12184 (N_12184,N_11250,N_11711);
nand U12185 (N_12185,N_11775,N_11623);
xnor U12186 (N_12186,N_11295,N_11716);
nand U12187 (N_12187,N_11662,N_11795);
and U12188 (N_12188,N_11775,N_11536);
nand U12189 (N_12189,N_11645,N_11838);
and U12190 (N_12190,N_11479,N_11288);
nor U12191 (N_12191,N_11281,N_11851);
nor U12192 (N_12192,N_11393,N_11376);
nor U12193 (N_12193,N_11725,N_11684);
xnor U12194 (N_12194,N_11426,N_11646);
or U12195 (N_12195,N_11440,N_11760);
nor U12196 (N_12196,N_11681,N_11318);
or U12197 (N_12197,N_11460,N_11411);
or U12198 (N_12198,N_11607,N_11483);
nand U12199 (N_12199,N_11530,N_11368);
nand U12200 (N_12200,N_11382,N_11397);
nand U12201 (N_12201,N_11760,N_11583);
or U12202 (N_12202,N_11697,N_11402);
xor U12203 (N_12203,N_11856,N_11607);
nor U12204 (N_12204,N_11270,N_11556);
xor U12205 (N_12205,N_11333,N_11682);
nand U12206 (N_12206,N_11680,N_11422);
nand U12207 (N_12207,N_11581,N_11874);
nor U12208 (N_12208,N_11658,N_11508);
or U12209 (N_12209,N_11433,N_11760);
nor U12210 (N_12210,N_11648,N_11839);
nor U12211 (N_12211,N_11363,N_11868);
xor U12212 (N_12212,N_11566,N_11604);
nand U12213 (N_12213,N_11562,N_11639);
nand U12214 (N_12214,N_11261,N_11821);
or U12215 (N_12215,N_11550,N_11608);
nand U12216 (N_12216,N_11676,N_11682);
and U12217 (N_12217,N_11713,N_11686);
nand U12218 (N_12218,N_11786,N_11668);
nand U12219 (N_12219,N_11381,N_11862);
and U12220 (N_12220,N_11610,N_11542);
nor U12221 (N_12221,N_11300,N_11688);
nand U12222 (N_12222,N_11289,N_11255);
nand U12223 (N_12223,N_11714,N_11251);
xor U12224 (N_12224,N_11402,N_11506);
or U12225 (N_12225,N_11690,N_11844);
nor U12226 (N_12226,N_11441,N_11487);
and U12227 (N_12227,N_11352,N_11548);
nand U12228 (N_12228,N_11687,N_11705);
and U12229 (N_12229,N_11408,N_11318);
nand U12230 (N_12230,N_11436,N_11757);
xnor U12231 (N_12231,N_11809,N_11271);
or U12232 (N_12232,N_11284,N_11697);
xnor U12233 (N_12233,N_11284,N_11782);
xor U12234 (N_12234,N_11688,N_11835);
nor U12235 (N_12235,N_11767,N_11519);
nand U12236 (N_12236,N_11624,N_11806);
xnor U12237 (N_12237,N_11390,N_11682);
nand U12238 (N_12238,N_11611,N_11550);
or U12239 (N_12239,N_11588,N_11720);
nor U12240 (N_12240,N_11397,N_11455);
xor U12241 (N_12241,N_11698,N_11491);
nand U12242 (N_12242,N_11262,N_11453);
or U12243 (N_12243,N_11862,N_11750);
xor U12244 (N_12244,N_11370,N_11437);
nor U12245 (N_12245,N_11530,N_11493);
nor U12246 (N_12246,N_11472,N_11504);
nand U12247 (N_12247,N_11597,N_11315);
xor U12248 (N_12248,N_11659,N_11837);
or U12249 (N_12249,N_11446,N_11300);
nand U12250 (N_12250,N_11675,N_11700);
nor U12251 (N_12251,N_11707,N_11383);
nand U12252 (N_12252,N_11782,N_11526);
and U12253 (N_12253,N_11453,N_11553);
and U12254 (N_12254,N_11659,N_11375);
nand U12255 (N_12255,N_11521,N_11683);
xnor U12256 (N_12256,N_11683,N_11842);
and U12257 (N_12257,N_11274,N_11485);
nor U12258 (N_12258,N_11761,N_11414);
or U12259 (N_12259,N_11399,N_11450);
and U12260 (N_12260,N_11855,N_11313);
nor U12261 (N_12261,N_11578,N_11558);
xnor U12262 (N_12262,N_11397,N_11453);
nand U12263 (N_12263,N_11859,N_11564);
nor U12264 (N_12264,N_11580,N_11771);
xor U12265 (N_12265,N_11373,N_11850);
or U12266 (N_12266,N_11820,N_11340);
and U12267 (N_12267,N_11628,N_11817);
nand U12268 (N_12268,N_11407,N_11602);
xor U12269 (N_12269,N_11422,N_11520);
xnor U12270 (N_12270,N_11274,N_11278);
or U12271 (N_12271,N_11644,N_11592);
xor U12272 (N_12272,N_11492,N_11514);
nor U12273 (N_12273,N_11307,N_11689);
nand U12274 (N_12274,N_11641,N_11784);
xor U12275 (N_12275,N_11414,N_11292);
or U12276 (N_12276,N_11770,N_11833);
nor U12277 (N_12277,N_11730,N_11800);
nor U12278 (N_12278,N_11671,N_11629);
and U12279 (N_12279,N_11761,N_11603);
nor U12280 (N_12280,N_11504,N_11536);
nor U12281 (N_12281,N_11252,N_11639);
nor U12282 (N_12282,N_11360,N_11719);
nand U12283 (N_12283,N_11597,N_11685);
nand U12284 (N_12284,N_11403,N_11674);
and U12285 (N_12285,N_11481,N_11864);
or U12286 (N_12286,N_11669,N_11711);
and U12287 (N_12287,N_11701,N_11521);
xnor U12288 (N_12288,N_11606,N_11463);
nand U12289 (N_12289,N_11603,N_11451);
nor U12290 (N_12290,N_11539,N_11402);
or U12291 (N_12291,N_11783,N_11856);
nand U12292 (N_12292,N_11340,N_11794);
xor U12293 (N_12293,N_11296,N_11721);
and U12294 (N_12294,N_11452,N_11857);
xnor U12295 (N_12295,N_11342,N_11620);
nor U12296 (N_12296,N_11681,N_11576);
nor U12297 (N_12297,N_11493,N_11460);
nor U12298 (N_12298,N_11257,N_11796);
nand U12299 (N_12299,N_11337,N_11364);
or U12300 (N_12300,N_11558,N_11526);
xor U12301 (N_12301,N_11754,N_11687);
xnor U12302 (N_12302,N_11515,N_11276);
or U12303 (N_12303,N_11570,N_11775);
nor U12304 (N_12304,N_11650,N_11443);
and U12305 (N_12305,N_11644,N_11772);
nor U12306 (N_12306,N_11803,N_11751);
and U12307 (N_12307,N_11651,N_11629);
nand U12308 (N_12308,N_11499,N_11330);
nand U12309 (N_12309,N_11469,N_11423);
or U12310 (N_12310,N_11713,N_11568);
nor U12311 (N_12311,N_11513,N_11306);
or U12312 (N_12312,N_11771,N_11424);
xor U12313 (N_12313,N_11552,N_11606);
xnor U12314 (N_12314,N_11810,N_11807);
nor U12315 (N_12315,N_11774,N_11717);
or U12316 (N_12316,N_11872,N_11600);
nand U12317 (N_12317,N_11494,N_11770);
nor U12318 (N_12318,N_11633,N_11464);
and U12319 (N_12319,N_11349,N_11393);
or U12320 (N_12320,N_11777,N_11688);
xnor U12321 (N_12321,N_11577,N_11824);
or U12322 (N_12322,N_11323,N_11664);
nor U12323 (N_12323,N_11275,N_11411);
nand U12324 (N_12324,N_11332,N_11359);
nand U12325 (N_12325,N_11816,N_11297);
xnor U12326 (N_12326,N_11294,N_11734);
xor U12327 (N_12327,N_11637,N_11336);
nor U12328 (N_12328,N_11743,N_11641);
nor U12329 (N_12329,N_11355,N_11468);
and U12330 (N_12330,N_11839,N_11419);
or U12331 (N_12331,N_11602,N_11752);
xnor U12332 (N_12332,N_11607,N_11641);
and U12333 (N_12333,N_11355,N_11441);
xor U12334 (N_12334,N_11726,N_11510);
or U12335 (N_12335,N_11841,N_11363);
nor U12336 (N_12336,N_11330,N_11636);
nor U12337 (N_12337,N_11774,N_11694);
nand U12338 (N_12338,N_11273,N_11427);
or U12339 (N_12339,N_11788,N_11817);
and U12340 (N_12340,N_11625,N_11641);
and U12341 (N_12341,N_11709,N_11297);
nor U12342 (N_12342,N_11367,N_11458);
nand U12343 (N_12343,N_11600,N_11664);
or U12344 (N_12344,N_11865,N_11552);
and U12345 (N_12345,N_11818,N_11304);
nand U12346 (N_12346,N_11646,N_11412);
nor U12347 (N_12347,N_11365,N_11546);
xor U12348 (N_12348,N_11353,N_11795);
xnor U12349 (N_12349,N_11618,N_11363);
xor U12350 (N_12350,N_11783,N_11768);
nor U12351 (N_12351,N_11441,N_11395);
nor U12352 (N_12352,N_11347,N_11825);
nand U12353 (N_12353,N_11826,N_11383);
xnor U12354 (N_12354,N_11445,N_11733);
nor U12355 (N_12355,N_11290,N_11528);
or U12356 (N_12356,N_11604,N_11549);
xnor U12357 (N_12357,N_11575,N_11873);
xor U12358 (N_12358,N_11351,N_11435);
nor U12359 (N_12359,N_11694,N_11523);
nand U12360 (N_12360,N_11316,N_11346);
xnor U12361 (N_12361,N_11867,N_11587);
xor U12362 (N_12362,N_11270,N_11551);
xnor U12363 (N_12363,N_11545,N_11714);
nor U12364 (N_12364,N_11661,N_11529);
nor U12365 (N_12365,N_11379,N_11538);
nand U12366 (N_12366,N_11859,N_11505);
nor U12367 (N_12367,N_11724,N_11494);
xnor U12368 (N_12368,N_11567,N_11276);
and U12369 (N_12369,N_11309,N_11281);
nand U12370 (N_12370,N_11479,N_11675);
or U12371 (N_12371,N_11614,N_11831);
or U12372 (N_12372,N_11620,N_11396);
xnor U12373 (N_12373,N_11474,N_11395);
xnor U12374 (N_12374,N_11532,N_11712);
nor U12375 (N_12375,N_11330,N_11622);
or U12376 (N_12376,N_11312,N_11620);
or U12377 (N_12377,N_11700,N_11390);
and U12378 (N_12378,N_11692,N_11622);
and U12379 (N_12379,N_11585,N_11375);
and U12380 (N_12380,N_11695,N_11472);
nor U12381 (N_12381,N_11397,N_11678);
and U12382 (N_12382,N_11493,N_11531);
xor U12383 (N_12383,N_11608,N_11421);
nor U12384 (N_12384,N_11668,N_11530);
or U12385 (N_12385,N_11809,N_11326);
or U12386 (N_12386,N_11712,N_11873);
and U12387 (N_12387,N_11719,N_11354);
and U12388 (N_12388,N_11667,N_11458);
and U12389 (N_12389,N_11700,N_11624);
nor U12390 (N_12390,N_11419,N_11596);
nor U12391 (N_12391,N_11523,N_11559);
or U12392 (N_12392,N_11477,N_11267);
and U12393 (N_12393,N_11709,N_11419);
or U12394 (N_12394,N_11271,N_11854);
and U12395 (N_12395,N_11476,N_11595);
and U12396 (N_12396,N_11560,N_11548);
and U12397 (N_12397,N_11867,N_11670);
xor U12398 (N_12398,N_11795,N_11464);
and U12399 (N_12399,N_11489,N_11568);
nand U12400 (N_12400,N_11363,N_11470);
nor U12401 (N_12401,N_11579,N_11833);
or U12402 (N_12402,N_11509,N_11609);
xnor U12403 (N_12403,N_11383,N_11615);
nor U12404 (N_12404,N_11349,N_11734);
and U12405 (N_12405,N_11770,N_11459);
or U12406 (N_12406,N_11794,N_11631);
nor U12407 (N_12407,N_11547,N_11307);
and U12408 (N_12408,N_11799,N_11536);
or U12409 (N_12409,N_11544,N_11632);
xor U12410 (N_12410,N_11819,N_11716);
xnor U12411 (N_12411,N_11266,N_11755);
or U12412 (N_12412,N_11608,N_11691);
or U12413 (N_12413,N_11522,N_11462);
or U12414 (N_12414,N_11592,N_11252);
nand U12415 (N_12415,N_11568,N_11838);
nand U12416 (N_12416,N_11260,N_11375);
or U12417 (N_12417,N_11495,N_11291);
or U12418 (N_12418,N_11630,N_11653);
or U12419 (N_12419,N_11622,N_11588);
nand U12420 (N_12420,N_11415,N_11712);
and U12421 (N_12421,N_11612,N_11386);
xor U12422 (N_12422,N_11648,N_11403);
or U12423 (N_12423,N_11635,N_11367);
xor U12424 (N_12424,N_11774,N_11589);
nand U12425 (N_12425,N_11675,N_11392);
nand U12426 (N_12426,N_11714,N_11485);
and U12427 (N_12427,N_11800,N_11344);
and U12428 (N_12428,N_11313,N_11662);
xnor U12429 (N_12429,N_11491,N_11294);
or U12430 (N_12430,N_11483,N_11511);
nand U12431 (N_12431,N_11266,N_11414);
and U12432 (N_12432,N_11338,N_11425);
and U12433 (N_12433,N_11260,N_11373);
xnor U12434 (N_12434,N_11446,N_11265);
and U12435 (N_12435,N_11593,N_11530);
nor U12436 (N_12436,N_11540,N_11819);
nand U12437 (N_12437,N_11503,N_11343);
nor U12438 (N_12438,N_11513,N_11417);
or U12439 (N_12439,N_11390,N_11395);
or U12440 (N_12440,N_11689,N_11401);
and U12441 (N_12441,N_11695,N_11377);
nor U12442 (N_12442,N_11823,N_11727);
and U12443 (N_12443,N_11590,N_11806);
nor U12444 (N_12444,N_11469,N_11429);
or U12445 (N_12445,N_11416,N_11740);
and U12446 (N_12446,N_11416,N_11779);
xnor U12447 (N_12447,N_11512,N_11631);
xnor U12448 (N_12448,N_11468,N_11843);
xor U12449 (N_12449,N_11490,N_11765);
and U12450 (N_12450,N_11725,N_11740);
nor U12451 (N_12451,N_11397,N_11345);
and U12452 (N_12452,N_11337,N_11696);
nor U12453 (N_12453,N_11678,N_11630);
nand U12454 (N_12454,N_11758,N_11574);
xnor U12455 (N_12455,N_11395,N_11415);
nand U12456 (N_12456,N_11621,N_11761);
and U12457 (N_12457,N_11473,N_11343);
nand U12458 (N_12458,N_11307,N_11729);
or U12459 (N_12459,N_11849,N_11266);
or U12460 (N_12460,N_11463,N_11770);
nor U12461 (N_12461,N_11465,N_11838);
xnor U12462 (N_12462,N_11532,N_11802);
xor U12463 (N_12463,N_11738,N_11555);
or U12464 (N_12464,N_11471,N_11815);
and U12465 (N_12465,N_11824,N_11331);
nor U12466 (N_12466,N_11853,N_11551);
nand U12467 (N_12467,N_11806,N_11275);
or U12468 (N_12468,N_11643,N_11332);
nor U12469 (N_12469,N_11346,N_11465);
or U12470 (N_12470,N_11799,N_11593);
nor U12471 (N_12471,N_11784,N_11625);
xor U12472 (N_12472,N_11745,N_11653);
xor U12473 (N_12473,N_11702,N_11729);
or U12474 (N_12474,N_11511,N_11296);
nand U12475 (N_12475,N_11855,N_11674);
nand U12476 (N_12476,N_11618,N_11619);
and U12477 (N_12477,N_11675,N_11845);
xnor U12478 (N_12478,N_11254,N_11502);
nor U12479 (N_12479,N_11252,N_11531);
nand U12480 (N_12480,N_11580,N_11484);
xor U12481 (N_12481,N_11870,N_11358);
or U12482 (N_12482,N_11776,N_11309);
nand U12483 (N_12483,N_11356,N_11749);
and U12484 (N_12484,N_11574,N_11612);
nand U12485 (N_12485,N_11622,N_11343);
or U12486 (N_12486,N_11420,N_11832);
nor U12487 (N_12487,N_11355,N_11720);
xor U12488 (N_12488,N_11641,N_11498);
xnor U12489 (N_12489,N_11254,N_11264);
nor U12490 (N_12490,N_11282,N_11830);
or U12491 (N_12491,N_11855,N_11730);
nor U12492 (N_12492,N_11714,N_11681);
or U12493 (N_12493,N_11497,N_11767);
and U12494 (N_12494,N_11393,N_11837);
nand U12495 (N_12495,N_11466,N_11753);
and U12496 (N_12496,N_11847,N_11665);
and U12497 (N_12497,N_11345,N_11858);
nand U12498 (N_12498,N_11439,N_11366);
and U12499 (N_12499,N_11672,N_11275);
or U12500 (N_12500,N_12067,N_12253);
nand U12501 (N_12501,N_12061,N_12396);
or U12502 (N_12502,N_12459,N_11902);
and U12503 (N_12503,N_11979,N_12335);
and U12504 (N_12504,N_11926,N_12123);
xor U12505 (N_12505,N_12117,N_12444);
xor U12506 (N_12506,N_12007,N_12467);
nor U12507 (N_12507,N_12348,N_12005);
or U12508 (N_12508,N_12199,N_12343);
xnor U12509 (N_12509,N_11890,N_12355);
nand U12510 (N_12510,N_12351,N_11962);
nand U12511 (N_12511,N_12428,N_11950);
or U12512 (N_12512,N_11984,N_12200);
nand U12513 (N_12513,N_12080,N_12224);
or U12514 (N_12514,N_12051,N_11992);
and U12515 (N_12515,N_12213,N_12304);
nor U12516 (N_12516,N_12106,N_11918);
nand U12517 (N_12517,N_12104,N_12497);
nand U12518 (N_12518,N_12038,N_12074);
nand U12519 (N_12519,N_12491,N_12205);
nor U12520 (N_12520,N_11999,N_11996);
nand U12521 (N_12521,N_12210,N_12391);
or U12522 (N_12522,N_12327,N_12345);
nand U12523 (N_12523,N_11885,N_12385);
xnor U12524 (N_12524,N_11877,N_12220);
or U12525 (N_12525,N_12232,N_12119);
nand U12526 (N_12526,N_12115,N_12093);
nand U12527 (N_12527,N_12401,N_12369);
or U12528 (N_12528,N_12047,N_12181);
or U12529 (N_12529,N_12379,N_12053);
or U12530 (N_12530,N_12322,N_12145);
xnor U12531 (N_12531,N_12308,N_12399);
or U12532 (N_12532,N_12163,N_12154);
nor U12533 (N_12533,N_12045,N_12483);
and U12534 (N_12534,N_12350,N_12419);
xor U12535 (N_12535,N_12009,N_12493);
nor U12536 (N_12536,N_12344,N_12073);
nor U12537 (N_12537,N_12250,N_12226);
nand U12538 (N_12538,N_12398,N_12132);
nand U12539 (N_12539,N_12171,N_11947);
nand U12540 (N_12540,N_11881,N_12457);
and U12541 (N_12541,N_12228,N_12394);
and U12542 (N_12542,N_11923,N_11980);
nor U12543 (N_12543,N_12258,N_12020);
or U12544 (N_12544,N_12179,N_11987);
nor U12545 (N_12545,N_12184,N_12138);
or U12546 (N_12546,N_11944,N_11989);
xor U12547 (N_12547,N_12278,N_12384);
nand U12548 (N_12548,N_12230,N_11888);
xnor U12549 (N_12549,N_12447,N_12361);
nand U12550 (N_12550,N_12421,N_12412);
or U12551 (N_12551,N_12298,N_12388);
xnor U12552 (N_12552,N_11879,N_12353);
and U12553 (N_12553,N_12075,N_11978);
and U12554 (N_12554,N_11912,N_11922);
or U12555 (N_12555,N_12206,N_12452);
xor U12556 (N_12556,N_12269,N_12069);
or U12557 (N_12557,N_12393,N_11955);
nand U12558 (N_12558,N_12267,N_12078);
or U12559 (N_12559,N_12328,N_12368);
xor U12560 (N_12560,N_12266,N_12141);
xnor U12561 (N_12561,N_12499,N_12144);
nand U12562 (N_12562,N_12019,N_12221);
and U12563 (N_12563,N_12071,N_12188);
or U12564 (N_12564,N_12131,N_12116);
or U12565 (N_12565,N_12498,N_12279);
and U12566 (N_12566,N_12111,N_12418);
nand U12567 (N_12567,N_12032,N_12317);
or U12568 (N_12568,N_12281,N_12100);
or U12569 (N_12569,N_12041,N_12357);
and U12570 (N_12570,N_12150,N_12195);
and U12571 (N_12571,N_11986,N_12110);
nand U12572 (N_12572,N_11908,N_12052);
or U12573 (N_12573,N_12187,N_11892);
xnor U12574 (N_12574,N_12089,N_12270);
and U12575 (N_12575,N_12063,N_12326);
or U12576 (N_12576,N_12347,N_12022);
nor U12577 (N_12577,N_12470,N_12462);
nor U12578 (N_12578,N_11905,N_12120);
nand U12579 (N_12579,N_12072,N_11993);
nor U12580 (N_12580,N_11981,N_12157);
and U12581 (N_12581,N_12377,N_12215);
nand U12582 (N_12582,N_12092,N_12122);
nor U12583 (N_12583,N_12336,N_12128);
xor U12584 (N_12584,N_12370,N_11973);
nand U12585 (N_12585,N_12318,N_12284);
nand U12586 (N_12586,N_12170,N_12433);
xor U12587 (N_12587,N_12243,N_12028);
xnor U12588 (N_12588,N_12314,N_12241);
xnor U12589 (N_12589,N_11891,N_12341);
nor U12590 (N_12590,N_12222,N_12360);
nor U12591 (N_12591,N_11900,N_12012);
and U12592 (N_12592,N_12313,N_12404);
nor U12593 (N_12593,N_12136,N_12422);
xor U12594 (N_12594,N_11896,N_11974);
nor U12595 (N_12595,N_12425,N_12091);
and U12596 (N_12596,N_12358,N_11954);
and U12597 (N_12597,N_11901,N_11972);
and U12598 (N_12598,N_12137,N_12485);
and U12599 (N_12599,N_12246,N_12437);
nor U12600 (N_12600,N_11941,N_12134);
and U12601 (N_12601,N_12302,N_12242);
and U12602 (N_12602,N_12449,N_11924);
and U12603 (N_12603,N_12133,N_12159);
nand U12604 (N_12604,N_11878,N_11969);
xor U12605 (N_12605,N_11991,N_12446);
nor U12606 (N_12606,N_12000,N_12265);
nand U12607 (N_12607,N_12477,N_12306);
or U12608 (N_12608,N_12407,N_12310);
nand U12609 (N_12609,N_12008,N_12097);
nand U12610 (N_12610,N_12465,N_12056);
xor U12611 (N_12611,N_11988,N_12489);
nand U12612 (N_12612,N_12453,N_12408);
or U12613 (N_12613,N_12135,N_12436);
or U12614 (N_12614,N_12011,N_12216);
xor U12615 (N_12615,N_11958,N_12186);
and U12616 (N_12616,N_12088,N_12321);
xor U12617 (N_12617,N_12229,N_12395);
or U12618 (N_12618,N_12147,N_12148);
xnor U12619 (N_12619,N_12027,N_12440);
xor U12620 (N_12620,N_11968,N_11935);
and U12621 (N_12621,N_12176,N_12429);
or U12622 (N_12622,N_12125,N_12160);
xor U12623 (N_12623,N_12264,N_12451);
nand U12624 (N_12624,N_12225,N_11917);
or U12625 (N_12625,N_12083,N_12413);
nand U12626 (N_12626,N_11966,N_12285);
nor U12627 (N_12627,N_11889,N_12001);
xor U12628 (N_12628,N_12139,N_12113);
or U12629 (N_12629,N_12261,N_12098);
nor U12630 (N_12630,N_11975,N_12496);
nand U12631 (N_12631,N_12185,N_12202);
nand U12632 (N_12632,N_12417,N_12247);
xor U12633 (N_12633,N_12030,N_12256);
and U12634 (N_12634,N_12077,N_12441);
or U12635 (N_12635,N_11951,N_12323);
nor U12636 (N_12636,N_12479,N_12332);
and U12637 (N_12637,N_12237,N_12356);
nand U12638 (N_12638,N_12240,N_12114);
xor U12639 (N_12639,N_12108,N_12082);
and U12640 (N_12640,N_12183,N_12055);
xor U12641 (N_12641,N_12272,N_12456);
xor U12642 (N_12642,N_12227,N_12464);
xnor U12643 (N_12643,N_12442,N_12448);
or U12644 (N_12644,N_12168,N_11931);
xnor U12645 (N_12645,N_11976,N_12178);
nor U12646 (N_12646,N_12014,N_12434);
xor U12647 (N_12647,N_12214,N_11990);
xor U12648 (N_12648,N_12024,N_12129);
nand U12649 (N_12649,N_11894,N_12312);
or U12650 (N_12650,N_11956,N_12432);
and U12651 (N_12651,N_12295,N_12219);
nand U12652 (N_12652,N_11934,N_12198);
xnor U12653 (N_12653,N_12372,N_12424);
nor U12654 (N_12654,N_12268,N_12153);
nand U12655 (N_12655,N_12300,N_12263);
and U12656 (N_12656,N_11898,N_12040);
and U12657 (N_12657,N_12380,N_12244);
nand U12658 (N_12658,N_11884,N_11961);
or U12659 (N_12659,N_12165,N_12469);
and U12660 (N_12660,N_11940,N_11964);
and U12661 (N_12661,N_12487,N_11959);
and U12662 (N_12662,N_12233,N_12478);
xor U12663 (N_12663,N_12172,N_12340);
nor U12664 (N_12664,N_12017,N_11893);
or U12665 (N_12665,N_11919,N_11977);
nand U12666 (N_12666,N_12271,N_12021);
and U12667 (N_12667,N_12494,N_11909);
xnor U12668 (N_12668,N_12495,N_12420);
and U12669 (N_12669,N_12238,N_12048);
and U12670 (N_12670,N_12293,N_12324);
nand U12671 (N_12671,N_12463,N_12189);
xor U12672 (N_12672,N_12414,N_12085);
nor U12673 (N_12673,N_12068,N_12239);
or U12674 (N_12674,N_11998,N_11921);
nand U12675 (N_12675,N_12410,N_12212);
nand U12676 (N_12676,N_11882,N_11939);
or U12677 (N_12677,N_11895,N_12130);
xnor U12678 (N_12678,N_12337,N_12297);
or U12679 (N_12679,N_12066,N_11965);
nor U12680 (N_12680,N_12445,N_12392);
and U12681 (N_12681,N_12015,N_12288);
nand U12682 (N_12682,N_12018,N_12010);
nor U12683 (N_12683,N_12415,N_12315);
xor U12684 (N_12684,N_12059,N_11929);
nand U12685 (N_12685,N_12174,N_12107);
and U12686 (N_12686,N_11906,N_12329);
xnor U12687 (N_12687,N_12466,N_12177);
xor U12688 (N_12688,N_12127,N_12034);
and U12689 (N_12689,N_12164,N_11948);
nor U12690 (N_12690,N_12458,N_11903);
xnor U12691 (N_12691,N_11949,N_12109);
or U12692 (N_12692,N_12362,N_12101);
or U12693 (N_12693,N_12480,N_12096);
and U12694 (N_12694,N_11995,N_12382);
xor U12695 (N_12695,N_12389,N_12249);
xnor U12696 (N_12696,N_12076,N_12488);
and U12697 (N_12697,N_12367,N_12140);
nand U12698 (N_12698,N_12474,N_12305);
nand U12699 (N_12699,N_12276,N_12283);
nor U12700 (N_12700,N_12484,N_12460);
nor U12701 (N_12701,N_12065,N_11887);
nand U12702 (N_12702,N_12402,N_12042);
nand U12703 (N_12703,N_12058,N_12173);
nand U12704 (N_12704,N_12426,N_11911);
nand U12705 (N_12705,N_12403,N_12245);
or U12706 (N_12706,N_11963,N_12405);
nand U12707 (N_12707,N_12430,N_12259);
nand U12708 (N_12708,N_12359,N_11937);
xor U12709 (N_12709,N_12274,N_12231);
xnor U12710 (N_12710,N_12217,N_12255);
or U12711 (N_12711,N_12029,N_12036);
and U12712 (N_12712,N_12390,N_12049);
and U12713 (N_12713,N_11910,N_11883);
xor U12714 (N_12714,N_12475,N_12280);
nor U12715 (N_12715,N_12381,N_11957);
and U12716 (N_12716,N_12349,N_12218);
nand U12717 (N_12717,N_12476,N_12364);
nand U12718 (N_12718,N_12025,N_12124);
or U12719 (N_12719,N_11876,N_12481);
or U12720 (N_12720,N_12490,N_11936);
xnor U12721 (N_12721,N_12169,N_12375);
nand U12722 (N_12722,N_12152,N_12383);
nand U12723 (N_12723,N_12211,N_12333);
or U12724 (N_12724,N_11942,N_12050);
or U12725 (N_12725,N_12090,N_12182);
nand U12726 (N_12726,N_12035,N_12316);
nand U12727 (N_12727,N_12190,N_12363);
and U12728 (N_12728,N_12473,N_12033);
nand U12729 (N_12729,N_12064,N_12095);
nor U12730 (N_12730,N_12112,N_12287);
xnor U12731 (N_12731,N_12286,N_12006);
nor U12732 (N_12732,N_12037,N_11927);
and U12733 (N_12733,N_12234,N_12290);
and U12734 (N_12734,N_11945,N_12443);
xor U12735 (N_12735,N_12235,N_11897);
nand U12736 (N_12736,N_12207,N_12303);
nand U12737 (N_12737,N_11953,N_12439);
nor U12738 (N_12738,N_12292,N_12197);
nand U12739 (N_12739,N_11930,N_12406);
or U12740 (N_12740,N_12400,N_12026);
and U12741 (N_12741,N_12167,N_12282);
and U12742 (N_12742,N_11913,N_12468);
and U12743 (N_12743,N_12455,N_12378);
and U12744 (N_12744,N_12325,N_12454);
or U12745 (N_12745,N_12423,N_12252);
nor U12746 (N_12746,N_12193,N_12338);
xor U12747 (N_12747,N_12309,N_12311);
or U12748 (N_12748,N_12334,N_12411);
and U12749 (N_12749,N_12373,N_12166);
and U12750 (N_12750,N_12438,N_11983);
xor U12751 (N_12751,N_12260,N_12158);
or U12752 (N_12752,N_12492,N_12149);
or U12753 (N_12753,N_12427,N_11938);
nor U12754 (N_12754,N_12203,N_12275);
nand U12755 (N_12755,N_12201,N_12194);
nor U12756 (N_12756,N_12002,N_11971);
nand U12757 (N_12757,N_12376,N_11933);
or U12758 (N_12758,N_12482,N_12081);
nand U12759 (N_12759,N_12086,N_12277);
nor U12760 (N_12760,N_12013,N_12191);
nor U12761 (N_12761,N_11920,N_11960);
nor U12762 (N_12762,N_12208,N_12435);
nor U12763 (N_12763,N_12156,N_12461);
xnor U12764 (N_12764,N_12057,N_12043);
nand U12765 (N_12765,N_11946,N_12342);
and U12766 (N_12766,N_12084,N_12118);
nor U12767 (N_12767,N_12121,N_12196);
nor U12768 (N_12768,N_12162,N_12431);
xnor U12769 (N_12769,N_12307,N_12161);
or U12770 (N_12770,N_12262,N_12102);
or U12771 (N_12771,N_12054,N_12352);
nand U12772 (N_12772,N_11997,N_12039);
nand U12773 (N_12773,N_11967,N_12155);
and U12774 (N_12774,N_12103,N_12004);
or U12775 (N_12775,N_12371,N_12320);
or U12776 (N_12776,N_12254,N_12331);
nor U12777 (N_12777,N_11925,N_12319);
xor U12778 (N_12778,N_12099,N_12248);
nand U12779 (N_12779,N_12472,N_12062);
nand U12780 (N_12780,N_11943,N_11928);
and U12781 (N_12781,N_12471,N_12209);
nand U12782 (N_12782,N_12236,N_11994);
xnor U12783 (N_12783,N_11970,N_11952);
nand U12784 (N_12784,N_12079,N_12204);
nand U12785 (N_12785,N_12023,N_12450);
or U12786 (N_12786,N_11904,N_11915);
xor U12787 (N_12787,N_12105,N_12126);
and U12788 (N_12788,N_12301,N_12346);
nor U12789 (N_12789,N_12142,N_12289);
or U12790 (N_12790,N_12486,N_12044);
nand U12791 (N_12791,N_12192,N_12087);
xor U12792 (N_12792,N_11916,N_12273);
or U12793 (N_12793,N_12299,N_12257);
and U12794 (N_12794,N_12016,N_12151);
nor U12795 (N_12795,N_11914,N_12060);
xor U12796 (N_12796,N_11985,N_12416);
or U12797 (N_12797,N_12143,N_11880);
nor U12798 (N_12798,N_12387,N_12223);
xnor U12799 (N_12799,N_12365,N_12386);
nand U12800 (N_12800,N_12180,N_12354);
or U12801 (N_12801,N_12339,N_11932);
or U12802 (N_12802,N_11899,N_12330);
nor U12803 (N_12803,N_11875,N_12070);
xor U12804 (N_12804,N_12251,N_11886);
nand U12805 (N_12805,N_12003,N_12146);
and U12806 (N_12806,N_12291,N_12366);
nor U12807 (N_12807,N_11907,N_12094);
nor U12808 (N_12808,N_12175,N_12294);
xnor U12809 (N_12809,N_12031,N_12046);
or U12810 (N_12810,N_12374,N_11982);
nor U12811 (N_12811,N_12296,N_12409);
or U12812 (N_12812,N_12397,N_12358);
nand U12813 (N_12813,N_12264,N_11946);
xor U12814 (N_12814,N_12328,N_12237);
and U12815 (N_12815,N_11972,N_12013);
nand U12816 (N_12816,N_11893,N_12426);
and U12817 (N_12817,N_12359,N_12029);
xor U12818 (N_12818,N_11909,N_12430);
nor U12819 (N_12819,N_12437,N_12333);
xnor U12820 (N_12820,N_12493,N_12413);
nor U12821 (N_12821,N_12083,N_12038);
xnor U12822 (N_12822,N_11945,N_12290);
nor U12823 (N_12823,N_12359,N_12377);
nor U12824 (N_12824,N_12482,N_11986);
nor U12825 (N_12825,N_12350,N_12171);
nand U12826 (N_12826,N_11938,N_12196);
or U12827 (N_12827,N_12424,N_12483);
nand U12828 (N_12828,N_11990,N_12036);
xor U12829 (N_12829,N_12493,N_12377);
nor U12830 (N_12830,N_11937,N_11916);
or U12831 (N_12831,N_12079,N_12101);
xnor U12832 (N_12832,N_11936,N_11887);
xor U12833 (N_12833,N_11917,N_12209);
nor U12834 (N_12834,N_12270,N_11962);
nor U12835 (N_12835,N_11884,N_12293);
nand U12836 (N_12836,N_11956,N_11882);
and U12837 (N_12837,N_12475,N_12095);
xor U12838 (N_12838,N_12140,N_11974);
nand U12839 (N_12839,N_12358,N_12010);
and U12840 (N_12840,N_12069,N_12459);
and U12841 (N_12841,N_12490,N_12018);
or U12842 (N_12842,N_11895,N_12314);
xnor U12843 (N_12843,N_12348,N_11988);
nor U12844 (N_12844,N_12392,N_11904);
or U12845 (N_12845,N_12409,N_12168);
and U12846 (N_12846,N_12296,N_12445);
nor U12847 (N_12847,N_12137,N_12352);
and U12848 (N_12848,N_12373,N_11911);
and U12849 (N_12849,N_12016,N_12152);
nor U12850 (N_12850,N_12438,N_12116);
or U12851 (N_12851,N_12020,N_12040);
nand U12852 (N_12852,N_12377,N_12389);
xnor U12853 (N_12853,N_12130,N_12236);
or U12854 (N_12854,N_11975,N_11979);
nor U12855 (N_12855,N_12022,N_12316);
nor U12856 (N_12856,N_12057,N_11890);
xor U12857 (N_12857,N_12428,N_12242);
or U12858 (N_12858,N_12204,N_12307);
nor U12859 (N_12859,N_12263,N_12071);
or U12860 (N_12860,N_11994,N_11909);
xnor U12861 (N_12861,N_11881,N_11882);
xnor U12862 (N_12862,N_11901,N_12201);
and U12863 (N_12863,N_12020,N_12048);
xor U12864 (N_12864,N_12109,N_12409);
or U12865 (N_12865,N_12222,N_12096);
and U12866 (N_12866,N_12243,N_12168);
nand U12867 (N_12867,N_12251,N_12160);
or U12868 (N_12868,N_12070,N_12316);
and U12869 (N_12869,N_12103,N_12210);
nand U12870 (N_12870,N_11979,N_12074);
nor U12871 (N_12871,N_11898,N_12239);
or U12872 (N_12872,N_12383,N_12340);
or U12873 (N_12873,N_12468,N_12212);
nand U12874 (N_12874,N_11907,N_12417);
nor U12875 (N_12875,N_12194,N_12427);
and U12876 (N_12876,N_11943,N_12059);
and U12877 (N_12877,N_12115,N_11921);
or U12878 (N_12878,N_12270,N_12070);
or U12879 (N_12879,N_12062,N_12449);
nor U12880 (N_12880,N_11953,N_11936);
or U12881 (N_12881,N_12469,N_12036);
xnor U12882 (N_12882,N_12217,N_12365);
nor U12883 (N_12883,N_12277,N_12168);
or U12884 (N_12884,N_12362,N_12042);
xnor U12885 (N_12885,N_12465,N_12249);
or U12886 (N_12886,N_11966,N_12283);
or U12887 (N_12887,N_11993,N_12116);
or U12888 (N_12888,N_12496,N_12058);
or U12889 (N_12889,N_12062,N_12073);
xor U12890 (N_12890,N_11980,N_12140);
nor U12891 (N_12891,N_11883,N_12439);
xnor U12892 (N_12892,N_12274,N_12005);
or U12893 (N_12893,N_12443,N_12375);
nand U12894 (N_12894,N_11887,N_11954);
and U12895 (N_12895,N_12312,N_12250);
or U12896 (N_12896,N_12499,N_12454);
or U12897 (N_12897,N_12458,N_12181);
and U12898 (N_12898,N_12314,N_11902);
and U12899 (N_12899,N_11912,N_12232);
or U12900 (N_12900,N_12123,N_12004);
or U12901 (N_12901,N_12033,N_12482);
nand U12902 (N_12902,N_12419,N_12477);
and U12903 (N_12903,N_12361,N_12188);
xor U12904 (N_12904,N_12363,N_12468);
nand U12905 (N_12905,N_12267,N_12486);
xnor U12906 (N_12906,N_11908,N_12381);
xor U12907 (N_12907,N_12103,N_12347);
nor U12908 (N_12908,N_12164,N_12072);
and U12909 (N_12909,N_12032,N_12279);
and U12910 (N_12910,N_12478,N_12168);
and U12911 (N_12911,N_12424,N_12446);
and U12912 (N_12912,N_12354,N_11897);
or U12913 (N_12913,N_11906,N_11982);
nand U12914 (N_12914,N_12236,N_12157);
nand U12915 (N_12915,N_11933,N_12335);
nor U12916 (N_12916,N_12386,N_12387);
or U12917 (N_12917,N_12329,N_12236);
xnor U12918 (N_12918,N_12217,N_12472);
or U12919 (N_12919,N_12315,N_11978);
or U12920 (N_12920,N_12124,N_12203);
xor U12921 (N_12921,N_11921,N_12441);
nor U12922 (N_12922,N_12380,N_12450);
xnor U12923 (N_12923,N_11980,N_12094);
or U12924 (N_12924,N_12390,N_12202);
nand U12925 (N_12925,N_12307,N_12387);
xor U12926 (N_12926,N_12198,N_12033);
xnor U12927 (N_12927,N_12459,N_11903);
nand U12928 (N_12928,N_11906,N_11976);
nand U12929 (N_12929,N_12173,N_12105);
or U12930 (N_12930,N_12472,N_12380);
and U12931 (N_12931,N_12325,N_12420);
or U12932 (N_12932,N_12028,N_12001);
or U12933 (N_12933,N_11939,N_12010);
nor U12934 (N_12934,N_12466,N_12082);
or U12935 (N_12935,N_12094,N_11902);
nand U12936 (N_12936,N_12234,N_12424);
nand U12937 (N_12937,N_12425,N_11973);
xnor U12938 (N_12938,N_12058,N_11897);
nand U12939 (N_12939,N_12380,N_11908);
and U12940 (N_12940,N_11954,N_12498);
nor U12941 (N_12941,N_12210,N_12279);
or U12942 (N_12942,N_11952,N_11950);
and U12943 (N_12943,N_12239,N_11917);
nand U12944 (N_12944,N_12052,N_12222);
and U12945 (N_12945,N_12175,N_11898);
nor U12946 (N_12946,N_11976,N_12403);
xnor U12947 (N_12947,N_12035,N_11979);
and U12948 (N_12948,N_12143,N_12292);
xor U12949 (N_12949,N_12079,N_12487);
or U12950 (N_12950,N_12458,N_12363);
nand U12951 (N_12951,N_11897,N_12057);
nand U12952 (N_12952,N_12021,N_12285);
xor U12953 (N_12953,N_11992,N_12285);
or U12954 (N_12954,N_12176,N_11887);
nor U12955 (N_12955,N_12030,N_12136);
xnor U12956 (N_12956,N_12434,N_11902);
nand U12957 (N_12957,N_11899,N_12403);
and U12958 (N_12958,N_12362,N_12114);
nor U12959 (N_12959,N_12156,N_12339);
xnor U12960 (N_12960,N_12096,N_12092);
or U12961 (N_12961,N_12342,N_12298);
xor U12962 (N_12962,N_12388,N_12471);
or U12963 (N_12963,N_12341,N_12194);
nand U12964 (N_12964,N_12101,N_12210);
nand U12965 (N_12965,N_11964,N_12208);
nor U12966 (N_12966,N_12197,N_11899);
and U12967 (N_12967,N_12217,N_11988);
nand U12968 (N_12968,N_12331,N_12224);
xor U12969 (N_12969,N_12196,N_12428);
and U12970 (N_12970,N_12491,N_12055);
or U12971 (N_12971,N_12362,N_12408);
or U12972 (N_12972,N_12289,N_11905);
xor U12973 (N_12973,N_12157,N_12097);
and U12974 (N_12974,N_12163,N_12133);
and U12975 (N_12975,N_11910,N_12474);
and U12976 (N_12976,N_12263,N_12436);
nor U12977 (N_12977,N_12455,N_12388);
or U12978 (N_12978,N_12388,N_12189);
nor U12979 (N_12979,N_12006,N_12315);
nor U12980 (N_12980,N_12467,N_12102);
and U12981 (N_12981,N_12021,N_11875);
nor U12982 (N_12982,N_11900,N_12202);
nand U12983 (N_12983,N_12293,N_12411);
nand U12984 (N_12984,N_12251,N_12123);
xor U12985 (N_12985,N_12206,N_12040);
or U12986 (N_12986,N_12337,N_12376);
xor U12987 (N_12987,N_12230,N_12404);
nor U12988 (N_12988,N_11906,N_12233);
and U12989 (N_12989,N_12238,N_12439);
nor U12990 (N_12990,N_12466,N_11886);
or U12991 (N_12991,N_12319,N_11894);
nand U12992 (N_12992,N_12494,N_12166);
nor U12993 (N_12993,N_11957,N_11923);
nand U12994 (N_12994,N_12127,N_12411);
xnor U12995 (N_12995,N_12373,N_11912);
or U12996 (N_12996,N_12379,N_12123);
or U12997 (N_12997,N_12406,N_12442);
or U12998 (N_12998,N_12197,N_12282);
and U12999 (N_12999,N_11896,N_12220);
or U13000 (N_13000,N_12497,N_12371);
nor U13001 (N_13001,N_11963,N_12428);
xnor U13002 (N_13002,N_11932,N_12366);
xnor U13003 (N_13003,N_12364,N_12261);
xor U13004 (N_13004,N_12234,N_12199);
nand U13005 (N_13005,N_12321,N_12044);
nand U13006 (N_13006,N_12369,N_12024);
nand U13007 (N_13007,N_12258,N_11991);
xor U13008 (N_13008,N_11995,N_12105);
or U13009 (N_13009,N_11901,N_12078);
and U13010 (N_13010,N_12260,N_12234);
nand U13011 (N_13011,N_12372,N_12488);
nand U13012 (N_13012,N_11971,N_12187);
xnor U13013 (N_13013,N_12019,N_12183);
or U13014 (N_13014,N_11875,N_12421);
nand U13015 (N_13015,N_12194,N_12020);
and U13016 (N_13016,N_11910,N_12362);
nor U13017 (N_13017,N_12047,N_12201);
or U13018 (N_13018,N_12323,N_12472);
nor U13019 (N_13019,N_12436,N_11944);
and U13020 (N_13020,N_12329,N_12428);
and U13021 (N_13021,N_12477,N_12400);
nor U13022 (N_13022,N_12497,N_11894);
and U13023 (N_13023,N_12293,N_12371);
nand U13024 (N_13024,N_12468,N_12204);
xor U13025 (N_13025,N_12189,N_11900);
nor U13026 (N_13026,N_12470,N_11924);
or U13027 (N_13027,N_12218,N_12432);
nor U13028 (N_13028,N_12295,N_12442);
xnor U13029 (N_13029,N_12088,N_11940);
and U13030 (N_13030,N_11985,N_12499);
or U13031 (N_13031,N_12433,N_12200);
and U13032 (N_13032,N_12250,N_12496);
or U13033 (N_13033,N_12251,N_12158);
xnor U13034 (N_13034,N_12331,N_12386);
nand U13035 (N_13035,N_12088,N_12465);
nand U13036 (N_13036,N_12475,N_12344);
xor U13037 (N_13037,N_12166,N_12298);
nand U13038 (N_13038,N_11978,N_12190);
nand U13039 (N_13039,N_12038,N_12164);
or U13040 (N_13040,N_12449,N_11887);
or U13041 (N_13041,N_12081,N_12462);
nand U13042 (N_13042,N_12026,N_12322);
and U13043 (N_13043,N_11979,N_12150);
xor U13044 (N_13044,N_12260,N_12164);
nand U13045 (N_13045,N_12407,N_12475);
xor U13046 (N_13046,N_12227,N_12171);
or U13047 (N_13047,N_12140,N_12195);
and U13048 (N_13048,N_12113,N_11876);
nand U13049 (N_13049,N_12238,N_12450);
nor U13050 (N_13050,N_12462,N_12172);
and U13051 (N_13051,N_12427,N_12005);
or U13052 (N_13052,N_12279,N_12406);
nand U13053 (N_13053,N_12238,N_12392);
xnor U13054 (N_13054,N_12031,N_12342);
or U13055 (N_13055,N_11984,N_12181);
and U13056 (N_13056,N_12414,N_12112);
xnor U13057 (N_13057,N_12448,N_12189);
xor U13058 (N_13058,N_12091,N_12154);
xnor U13059 (N_13059,N_12466,N_12005);
nor U13060 (N_13060,N_12264,N_12340);
nand U13061 (N_13061,N_12041,N_12249);
xor U13062 (N_13062,N_11954,N_12116);
xnor U13063 (N_13063,N_12234,N_11966);
xnor U13064 (N_13064,N_12267,N_12274);
nand U13065 (N_13065,N_12475,N_12220);
nand U13066 (N_13066,N_12242,N_12008);
or U13067 (N_13067,N_12027,N_11992);
nand U13068 (N_13068,N_12007,N_12091);
nand U13069 (N_13069,N_12481,N_12296);
xor U13070 (N_13070,N_12203,N_11956);
or U13071 (N_13071,N_12472,N_12143);
xor U13072 (N_13072,N_12138,N_12260);
xnor U13073 (N_13073,N_12052,N_12448);
xor U13074 (N_13074,N_12061,N_12385);
or U13075 (N_13075,N_12451,N_12434);
xor U13076 (N_13076,N_11970,N_12003);
xor U13077 (N_13077,N_12256,N_11926);
xnor U13078 (N_13078,N_12441,N_12406);
and U13079 (N_13079,N_12014,N_12012);
xnor U13080 (N_13080,N_11902,N_12276);
or U13081 (N_13081,N_12320,N_12195);
or U13082 (N_13082,N_12278,N_12498);
nor U13083 (N_13083,N_12312,N_12029);
or U13084 (N_13084,N_12179,N_11968);
xor U13085 (N_13085,N_11978,N_11989);
nand U13086 (N_13086,N_11881,N_12261);
and U13087 (N_13087,N_11989,N_12455);
xor U13088 (N_13088,N_12246,N_11944);
nor U13089 (N_13089,N_12268,N_12345);
nor U13090 (N_13090,N_12086,N_12178);
and U13091 (N_13091,N_12124,N_12007);
and U13092 (N_13092,N_12488,N_12349);
or U13093 (N_13093,N_12487,N_12494);
or U13094 (N_13094,N_12410,N_12114);
xnor U13095 (N_13095,N_11884,N_12164);
xor U13096 (N_13096,N_12495,N_12295);
xnor U13097 (N_13097,N_12148,N_12408);
xor U13098 (N_13098,N_12444,N_12201);
or U13099 (N_13099,N_11892,N_12013);
and U13100 (N_13100,N_12004,N_12115);
and U13101 (N_13101,N_12381,N_12318);
and U13102 (N_13102,N_12256,N_12141);
nor U13103 (N_13103,N_12372,N_11915);
and U13104 (N_13104,N_12088,N_11962);
nor U13105 (N_13105,N_12135,N_11880);
nand U13106 (N_13106,N_11903,N_11985);
xnor U13107 (N_13107,N_12459,N_12017);
xnor U13108 (N_13108,N_12390,N_12322);
nor U13109 (N_13109,N_11972,N_11990);
or U13110 (N_13110,N_12271,N_12432);
nor U13111 (N_13111,N_12283,N_12167);
xnor U13112 (N_13112,N_12136,N_12216);
and U13113 (N_13113,N_12331,N_12323);
nand U13114 (N_13114,N_12160,N_12202);
or U13115 (N_13115,N_12113,N_12389);
xor U13116 (N_13116,N_12264,N_12089);
and U13117 (N_13117,N_11913,N_12253);
or U13118 (N_13118,N_12210,N_12360);
nand U13119 (N_13119,N_12348,N_11987);
nor U13120 (N_13120,N_12286,N_12335);
nand U13121 (N_13121,N_12304,N_12081);
or U13122 (N_13122,N_11880,N_11877);
nand U13123 (N_13123,N_12202,N_12067);
nand U13124 (N_13124,N_12226,N_12351);
xor U13125 (N_13125,N_12700,N_13017);
nand U13126 (N_13126,N_12989,N_12679);
or U13127 (N_13127,N_13102,N_12835);
xnor U13128 (N_13128,N_12721,N_12939);
nand U13129 (N_13129,N_12588,N_12547);
nand U13130 (N_13130,N_12572,N_12836);
xor U13131 (N_13131,N_12732,N_12957);
nor U13132 (N_13132,N_12845,N_12581);
and U13133 (N_13133,N_13006,N_12508);
nand U13134 (N_13134,N_13019,N_12841);
or U13135 (N_13135,N_13112,N_12675);
nand U13136 (N_13136,N_12544,N_12551);
and U13137 (N_13137,N_12652,N_12931);
nor U13138 (N_13138,N_13034,N_12698);
or U13139 (N_13139,N_13098,N_12659);
xnor U13140 (N_13140,N_12871,N_12828);
or U13141 (N_13141,N_13042,N_12999);
nor U13142 (N_13142,N_12580,N_13046);
xor U13143 (N_13143,N_13050,N_12833);
nor U13144 (N_13144,N_12952,N_12537);
xnor U13145 (N_13145,N_13108,N_12578);
nor U13146 (N_13146,N_12896,N_12759);
nor U13147 (N_13147,N_12583,N_12812);
nor U13148 (N_13148,N_12861,N_12628);
xnor U13149 (N_13149,N_12716,N_12942);
or U13150 (N_13150,N_13103,N_12656);
xnor U13151 (N_13151,N_13057,N_12921);
or U13152 (N_13152,N_13079,N_12631);
xnor U13153 (N_13153,N_12596,N_12762);
nand U13154 (N_13154,N_12662,N_12976);
nor U13155 (N_13155,N_12653,N_12515);
or U13156 (N_13156,N_12829,N_12963);
xnor U13157 (N_13157,N_12938,N_12809);
nand U13158 (N_13158,N_12726,N_12985);
or U13159 (N_13159,N_12814,N_12830);
nand U13160 (N_13160,N_13047,N_12786);
xor U13161 (N_13161,N_12876,N_13059);
or U13162 (N_13162,N_12710,N_12774);
and U13163 (N_13163,N_12758,N_12579);
or U13164 (N_13164,N_12901,N_12624);
and U13165 (N_13165,N_12980,N_12586);
nand U13166 (N_13166,N_12816,N_12600);
and U13167 (N_13167,N_12849,N_12855);
xnor U13168 (N_13168,N_13029,N_13093);
or U13169 (N_13169,N_12571,N_13099);
nand U13170 (N_13170,N_12977,N_12740);
xnor U13171 (N_13171,N_13066,N_12927);
xnor U13172 (N_13172,N_12920,N_12949);
nand U13173 (N_13173,N_12868,N_12639);
nor U13174 (N_13174,N_12561,N_12872);
xnor U13175 (N_13175,N_12516,N_12840);
nand U13176 (N_13176,N_12533,N_12661);
or U13177 (N_13177,N_12574,N_13115);
and U13178 (N_13178,N_12608,N_12904);
or U13179 (N_13179,N_12994,N_12900);
xor U13180 (N_13180,N_12644,N_12617);
nor U13181 (N_13181,N_12875,N_12787);
nor U13182 (N_13182,N_13088,N_12567);
and U13183 (N_13183,N_13001,N_12687);
nor U13184 (N_13184,N_12711,N_12688);
and U13185 (N_13185,N_12650,N_12613);
nand U13186 (N_13186,N_12693,N_12540);
or U13187 (N_13187,N_12893,N_12757);
nor U13188 (N_13188,N_12919,N_13061);
xor U13189 (N_13189,N_12504,N_12665);
xor U13190 (N_13190,N_12727,N_12903);
nor U13191 (N_13191,N_12674,N_13003);
xor U13192 (N_13192,N_12983,N_12995);
xnor U13193 (N_13193,N_13082,N_12546);
or U13194 (N_13194,N_12704,N_12801);
nor U13195 (N_13195,N_12843,N_13005);
or U13196 (N_13196,N_12557,N_12792);
xnor U13197 (N_13197,N_12569,N_12592);
or U13198 (N_13198,N_12930,N_12634);
and U13199 (N_13199,N_12556,N_12852);
xor U13200 (N_13200,N_13122,N_12510);
nor U13201 (N_13201,N_12768,N_12509);
xor U13202 (N_13202,N_12753,N_12971);
and U13203 (N_13203,N_13055,N_12582);
or U13204 (N_13204,N_12691,N_12606);
nor U13205 (N_13205,N_12568,N_12718);
and U13206 (N_13206,N_12746,N_12857);
or U13207 (N_13207,N_12605,N_12851);
nand U13208 (N_13208,N_12584,N_12941);
or U13209 (N_13209,N_12793,N_12791);
and U13210 (N_13210,N_12666,N_12623);
and U13211 (N_13211,N_12587,N_12784);
nand U13212 (N_13212,N_12678,N_13014);
and U13213 (N_13213,N_12979,N_12991);
or U13214 (N_13214,N_12724,N_12689);
xnor U13215 (N_13215,N_13117,N_12535);
or U13216 (N_13216,N_13012,N_12695);
nand U13217 (N_13217,N_12684,N_12632);
and U13218 (N_13218,N_12987,N_12880);
or U13219 (N_13219,N_13013,N_12839);
nor U13220 (N_13220,N_13036,N_12621);
and U13221 (N_13221,N_13077,N_12682);
nand U13222 (N_13222,N_12506,N_12668);
xor U13223 (N_13223,N_12525,N_12501);
or U13224 (N_13224,N_12545,N_12646);
xnor U13225 (N_13225,N_12573,N_12869);
xnor U13226 (N_13226,N_12602,N_12697);
and U13227 (N_13227,N_12813,N_12673);
xor U13228 (N_13228,N_12672,N_12860);
and U13229 (N_13229,N_12625,N_12519);
nand U13230 (N_13230,N_12731,N_13053);
xnor U13231 (N_13231,N_12645,N_12954);
and U13232 (N_13232,N_12680,N_12748);
nor U13233 (N_13233,N_12785,N_13097);
nor U13234 (N_13234,N_12790,N_13056);
nand U13235 (N_13235,N_13107,N_13062);
nand U13236 (N_13236,N_12637,N_12648);
nor U13237 (N_13237,N_12733,N_12570);
and U13238 (N_13238,N_12970,N_12946);
nor U13239 (N_13239,N_12948,N_12803);
nor U13240 (N_13240,N_12928,N_13040);
nor U13241 (N_13241,N_12912,N_12603);
nor U13242 (N_13242,N_12619,N_12781);
and U13243 (N_13243,N_12523,N_12526);
nand U13244 (N_13244,N_13045,N_12993);
nand U13245 (N_13245,N_12873,N_12734);
nand U13246 (N_13246,N_13052,N_13124);
xor U13247 (N_13247,N_12595,N_13025);
and U13248 (N_13248,N_13054,N_12788);
nand U13249 (N_13249,N_12522,N_12914);
xor U13250 (N_13250,N_13026,N_13049);
and U13251 (N_13251,N_12910,N_12658);
nor U13252 (N_13252,N_12969,N_12959);
nand U13253 (N_13253,N_12685,N_13120);
and U13254 (N_13254,N_12549,N_13101);
nand U13255 (N_13255,N_12530,N_12520);
nor U13256 (N_13256,N_12922,N_12647);
and U13257 (N_13257,N_12874,N_12690);
nor U13258 (N_13258,N_12925,N_12892);
or U13259 (N_13259,N_13007,N_12708);
and U13260 (N_13260,N_13072,N_12565);
nand U13261 (N_13261,N_12692,N_13116);
and U13262 (N_13262,N_12918,N_12854);
nand U13263 (N_13263,N_12823,N_12771);
nand U13264 (N_13264,N_13118,N_13091);
or U13265 (N_13265,N_13113,N_12769);
nor U13266 (N_13266,N_12597,N_13011);
nand U13267 (N_13267,N_12736,N_12507);
or U13268 (N_13268,N_12550,N_12681);
or U13269 (N_13269,N_13092,N_12907);
nand U13270 (N_13270,N_12825,N_12890);
nor U13271 (N_13271,N_12958,N_12780);
nor U13272 (N_13272,N_12953,N_13078);
or U13273 (N_13273,N_12538,N_12911);
xor U13274 (N_13274,N_13090,N_12915);
nor U13275 (N_13275,N_12749,N_12966);
or U13276 (N_13276,N_13123,N_12935);
or U13277 (N_13277,N_13105,N_12933);
and U13278 (N_13278,N_12782,N_13028);
xor U13279 (N_13279,N_12737,N_12752);
or U13280 (N_13280,N_12834,N_13031);
nand U13281 (N_13281,N_13044,N_13018);
or U13282 (N_13282,N_12601,N_13027);
nand U13283 (N_13283,N_12539,N_12616);
xor U13284 (N_13284,N_12811,N_12778);
xor U13285 (N_13285,N_13051,N_12548);
or U13286 (N_13286,N_12763,N_13089);
and U13287 (N_13287,N_13104,N_12642);
and U13288 (N_13288,N_12973,N_12831);
and U13289 (N_13289,N_12651,N_12889);
and U13290 (N_13290,N_12730,N_13084);
nand U13291 (N_13291,N_12968,N_12870);
or U13292 (N_13292,N_12905,N_12945);
xor U13293 (N_13293,N_13073,N_12967);
or U13294 (N_13294,N_12775,N_13020);
nand U13295 (N_13295,N_12513,N_13037);
nand U13296 (N_13296,N_12745,N_13109);
nand U13297 (N_13297,N_13075,N_12858);
or U13298 (N_13298,N_12575,N_13015);
nor U13299 (N_13299,N_12978,N_12951);
and U13300 (N_13300,N_12611,N_12883);
or U13301 (N_13301,N_13085,N_13043);
nor U13302 (N_13302,N_13087,N_12837);
nand U13303 (N_13303,N_13048,N_12885);
and U13304 (N_13304,N_12932,N_12898);
or U13305 (N_13305,N_12936,N_13094);
and U13306 (N_13306,N_13121,N_12773);
xor U13307 (N_13307,N_12856,N_12879);
nand U13308 (N_13308,N_12822,N_12853);
or U13309 (N_13309,N_13068,N_12997);
nor U13310 (N_13310,N_12529,N_12554);
nor U13311 (N_13311,N_12820,N_12585);
nand U13312 (N_13312,N_12747,N_12514);
and U13313 (N_13313,N_12709,N_12947);
nand U13314 (N_13314,N_12622,N_12598);
nand U13315 (N_13315,N_12988,N_12660);
nand U13316 (N_13316,N_12566,N_13038);
or U13317 (N_13317,N_13076,N_12810);
nor U13318 (N_13318,N_12795,N_12772);
xor U13319 (N_13319,N_12975,N_12909);
xor U13320 (N_13320,N_12886,N_12738);
nor U13321 (N_13321,N_12728,N_12511);
nor U13322 (N_13322,N_12913,N_12850);
nand U13323 (N_13323,N_13041,N_13096);
xor U13324 (N_13324,N_12589,N_12821);
or U13325 (N_13325,N_12524,N_12641);
or U13326 (N_13326,N_12751,N_12766);
xnor U13327 (N_13327,N_12804,N_12884);
nand U13328 (N_13328,N_13111,N_13106);
xor U13329 (N_13329,N_12703,N_12649);
or U13330 (N_13330,N_12517,N_12714);
nor U13331 (N_13331,N_12654,N_12760);
xor U13332 (N_13332,N_13058,N_12705);
and U13333 (N_13333,N_12640,N_12729);
nand U13334 (N_13334,N_12723,N_12630);
and U13335 (N_13335,N_12541,N_12962);
and U13336 (N_13336,N_12577,N_13070);
nand U13337 (N_13337,N_12827,N_12609);
nor U13338 (N_13338,N_13010,N_12844);
nor U13339 (N_13339,N_12564,N_12767);
or U13340 (N_13340,N_12859,N_12940);
nand U13341 (N_13341,N_12990,N_12532);
nand U13342 (N_13342,N_12750,N_13000);
xor U13343 (N_13343,N_13064,N_12981);
and U13344 (N_13344,N_12902,N_13114);
nor U13345 (N_13345,N_12965,N_12826);
nor U13346 (N_13346,N_12802,N_12770);
nor U13347 (N_13347,N_12563,N_12505);
nor U13348 (N_13348,N_12614,N_12742);
or U13349 (N_13349,N_12629,N_12846);
nand U13350 (N_13350,N_12618,N_13008);
or U13351 (N_13351,N_13100,N_12776);
or U13352 (N_13352,N_12719,N_12518);
xor U13353 (N_13353,N_12842,N_12699);
xor U13354 (N_13354,N_12677,N_12916);
nor U13355 (N_13355,N_12754,N_12725);
nand U13356 (N_13356,N_12756,N_12819);
and U13357 (N_13357,N_12635,N_13086);
or U13358 (N_13358,N_12862,N_12713);
nand U13359 (N_13359,N_12865,N_12996);
and U13360 (N_13360,N_12552,N_13030);
and U13361 (N_13361,N_12937,N_12739);
nor U13362 (N_13362,N_12906,N_12735);
or U13363 (N_13363,N_12599,N_12923);
and U13364 (N_13364,N_12663,N_12534);
or U13365 (N_13365,N_12838,N_12832);
and U13366 (N_13366,N_12972,N_12657);
xnor U13367 (N_13367,N_12669,N_12798);
or U13368 (N_13368,N_12615,N_12512);
nand U13369 (N_13369,N_12559,N_12655);
nand U13370 (N_13370,N_12591,N_12960);
or U13371 (N_13371,N_12926,N_12562);
nor U13372 (N_13372,N_12761,N_12717);
nor U13373 (N_13373,N_12878,N_12531);
and U13374 (N_13374,N_12604,N_12779);
or U13375 (N_13375,N_12882,N_12897);
xor U13376 (N_13376,N_12807,N_12636);
xor U13377 (N_13377,N_12743,N_12908);
or U13378 (N_13378,N_12887,N_12722);
xnor U13379 (N_13379,N_13110,N_12593);
nor U13380 (N_13380,N_12917,N_12929);
nand U13381 (N_13381,N_13063,N_12744);
nor U13382 (N_13382,N_12638,N_12943);
nor U13383 (N_13383,N_12824,N_12694);
nand U13384 (N_13384,N_12720,N_12696);
xnor U13385 (N_13385,N_13083,N_12702);
and U13386 (N_13386,N_12986,N_12671);
or U13387 (N_13387,N_13002,N_12502);
nand U13388 (N_13388,N_12500,N_12964);
nor U13389 (N_13389,N_12796,N_12982);
xor U13390 (N_13390,N_12899,N_12560);
xnor U13391 (N_13391,N_12764,N_12818);
nand U13392 (N_13392,N_12806,N_12894);
nand U13393 (N_13393,N_12895,N_12794);
nand U13394 (N_13394,N_12633,N_12706);
or U13395 (N_13395,N_12542,N_12797);
xor U13396 (N_13396,N_12799,N_12558);
nand U13397 (N_13397,N_12555,N_12715);
nor U13398 (N_13398,N_12594,N_12888);
and U13399 (N_13399,N_12643,N_12686);
nand U13400 (N_13400,N_12701,N_12956);
and U13401 (N_13401,N_13119,N_12664);
xor U13402 (N_13402,N_13033,N_12961);
and U13403 (N_13403,N_12815,N_13035);
or U13404 (N_13404,N_12998,N_12881);
and U13405 (N_13405,N_12864,N_12805);
xnor U13406 (N_13406,N_12707,N_12863);
or U13407 (N_13407,N_12950,N_12610);
nand U13408 (N_13408,N_12627,N_12777);
and U13409 (N_13409,N_12808,N_13081);
xnor U13410 (N_13410,N_13009,N_13021);
or U13411 (N_13411,N_12576,N_12848);
xnor U13412 (N_13412,N_12866,N_13067);
nand U13413 (N_13413,N_13095,N_12924);
xnor U13414 (N_13414,N_12607,N_13069);
nand U13415 (N_13415,N_13004,N_12800);
xnor U13416 (N_13416,N_12528,N_12620);
or U13417 (N_13417,N_12667,N_12543);
xor U13418 (N_13418,N_12553,N_12984);
and U13419 (N_13419,N_12934,N_13060);
or U13420 (N_13420,N_13071,N_12741);
and U13421 (N_13421,N_12536,N_12765);
xor U13422 (N_13422,N_12683,N_12527);
xor U13423 (N_13423,N_13074,N_12676);
nand U13424 (N_13424,N_12712,N_12755);
nand U13425 (N_13425,N_12944,N_12817);
and U13426 (N_13426,N_13080,N_12867);
nand U13427 (N_13427,N_12612,N_13032);
and U13428 (N_13428,N_12847,N_12521);
nand U13429 (N_13429,N_13023,N_13024);
nor U13430 (N_13430,N_12974,N_13016);
and U13431 (N_13431,N_12891,N_12590);
nor U13432 (N_13432,N_12789,N_12955);
xor U13433 (N_13433,N_12783,N_13022);
xnor U13434 (N_13434,N_13065,N_13039);
nor U13435 (N_13435,N_12670,N_12626);
or U13436 (N_13436,N_12503,N_12877);
xor U13437 (N_13437,N_12992,N_12902);
xnor U13438 (N_13438,N_13070,N_12822);
nor U13439 (N_13439,N_12759,N_12680);
or U13440 (N_13440,N_13010,N_12947);
xor U13441 (N_13441,N_12977,N_12562);
nand U13442 (N_13442,N_12668,N_13070);
nand U13443 (N_13443,N_12844,N_12927);
nand U13444 (N_13444,N_12599,N_12958);
and U13445 (N_13445,N_12657,N_13107);
nand U13446 (N_13446,N_12806,N_12940);
and U13447 (N_13447,N_12528,N_13116);
and U13448 (N_13448,N_12624,N_13003);
nor U13449 (N_13449,N_13038,N_12690);
nand U13450 (N_13450,N_13111,N_12530);
xnor U13451 (N_13451,N_12515,N_12770);
nand U13452 (N_13452,N_12763,N_12992);
and U13453 (N_13453,N_12830,N_12701);
xor U13454 (N_13454,N_12827,N_12929);
nor U13455 (N_13455,N_12519,N_12602);
nand U13456 (N_13456,N_12672,N_12728);
nand U13457 (N_13457,N_12896,N_12714);
and U13458 (N_13458,N_12550,N_12820);
or U13459 (N_13459,N_12597,N_12992);
xnor U13460 (N_13460,N_12539,N_12675);
or U13461 (N_13461,N_12521,N_12913);
or U13462 (N_13462,N_12552,N_13073);
or U13463 (N_13463,N_12968,N_12559);
or U13464 (N_13464,N_12517,N_12695);
and U13465 (N_13465,N_12571,N_12781);
nor U13466 (N_13466,N_12872,N_12834);
nor U13467 (N_13467,N_12785,N_12634);
and U13468 (N_13468,N_12940,N_12977);
nor U13469 (N_13469,N_12783,N_12583);
and U13470 (N_13470,N_12576,N_12514);
xnor U13471 (N_13471,N_12758,N_12666);
xnor U13472 (N_13472,N_12687,N_12957);
nand U13473 (N_13473,N_13038,N_12796);
or U13474 (N_13474,N_12595,N_12764);
or U13475 (N_13475,N_12816,N_13030);
xor U13476 (N_13476,N_12751,N_12708);
nor U13477 (N_13477,N_12721,N_13001);
or U13478 (N_13478,N_12739,N_12911);
and U13479 (N_13479,N_13104,N_13049);
or U13480 (N_13480,N_12872,N_12505);
or U13481 (N_13481,N_12540,N_12568);
nor U13482 (N_13482,N_12980,N_12899);
xor U13483 (N_13483,N_12654,N_12882);
nor U13484 (N_13484,N_12500,N_12738);
xnor U13485 (N_13485,N_13024,N_12918);
nand U13486 (N_13486,N_12541,N_12544);
xnor U13487 (N_13487,N_13075,N_12523);
nor U13488 (N_13488,N_12826,N_13042);
nand U13489 (N_13489,N_13123,N_12891);
xnor U13490 (N_13490,N_12905,N_12944);
and U13491 (N_13491,N_12754,N_13014);
nand U13492 (N_13492,N_12873,N_12738);
and U13493 (N_13493,N_12535,N_12996);
xnor U13494 (N_13494,N_12864,N_13074);
xnor U13495 (N_13495,N_12551,N_12801);
nor U13496 (N_13496,N_13124,N_12670);
nor U13497 (N_13497,N_12768,N_12857);
or U13498 (N_13498,N_12840,N_12783);
nor U13499 (N_13499,N_12755,N_12590);
nand U13500 (N_13500,N_12854,N_13102);
and U13501 (N_13501,N_12785,N_12728);
nor U13502 (N_13502,N_12627,N_12902);
nand U13503 (N_13503,N_12789,N_12885);
or U13504 (N_13504,N_12769,N_12781);
xor U13505 (N_13505,N_12663,N_12693);
xnor U13506 (N_13506,N_12563,N_12893);
nor U13507 (N_13507,N_12743,N_12725);
xnor U13508 (N_13508,N_13054,N_12748);
and U13509 (N_13509,N_12699,N_12876);
and U13510 (N_13510,N_13068,N_12785);
or U13511 (N_13511,N_12866,N_12534);
nand U13512 (N_13512,N_12737,N_12592);
or U13513 (N_13513,N_12978,N_12972);
or U13514 (N_13514,N_12850,N_12513);
and U13515 (N_13515,N_12768,N_12508);
xnor U13516 (N_13516,N_12968,N_12546);
xnor U13517 (N_13517,N_13069,N_12533);
or U13518 (N_13518,N_12639,N_13096);
or U13519 (N_13519,N_12770,N_12540);
nor U13520 (N_13520,N_12933,N_12567);
or U13521 (N_13521,N_12790,N_12846);
nor U13522 (N_13522,N_12806,N_12814);
xnor U13523 (N_13523,N_13088,N_12562);
or U13524 (N_13524,N_13035,N_12932);
nor U13525 (N_13525,N_12896,N_12546);
xor U13526 (N_13526,N_12956,N_12677);
and U13527 (N_13527,N_12698,N_13007);
nand U13528 (N_13528,N_12983,N_12724);
and U13529 (N_13529,N_12783,N_12805);
nor U13530 (N_13530,N_12554,N_12949);
xnor U13531 (N_13531,N_12802,N_12920);
and U13532 (N_13532,N_12929,N_12742);
nand U13533 (N_13533,N_12824,N_12888);
xor U13534 (N_13534,N_13105,N_12781);
or U13535 (N_13535,N_12789,N_12957);
nand U13536 (N_13536,N_12757,N_12902);
nor U13537 (N_13537,N_13046,N_12602);
nor U13538 (N_13538,N_12882,N_13044);
xor U13539 (N_13539,N_12555,N_12823);
xor U13540 (N_13540,N_12567,N_12534);
or U13541 (N_13541,N_12507,N_12583);
or U13542 (N_13542,N_13075,N_12958);
or U13543 (N_13543,N_13007,N_12760);
nand U13544 (N_13544,N_12820,N_13009);
or U13545 (N_13545,N_12904,N_12870);
or U13546 (N_13546,N_12864,N_12510);
and U13547 (N_13547,N_12676,N_13122);
or U13548 (N_13548,N_12715,N_13010);
xnor U13549 (N_13549,N_12984,N_13013);
xnor U13550 (N_13550,N_12588,N_12535);
or U13551 (N_13551,N_12653,N_12911);
or U13552 (N_13552,N_12563,N_12796);
nand U13553 (N_13553,N_12801,N_12783);
nor U13554 (N_13554,N_12735,N_13089);
nand U13555 (N_13555,N_12817,N_12933);
xnor U13556 (N_13556,N_12713,N_12518);
nor U13557 (N_13557,N_12628,N_12741);
or U13558 (N_13558,N_13006,N_12674);
nand U13559 (N_13559,N_13005,N_12768);
nor U13560 (N_13560,N_12556,N_12648);
nand U13561 (N_13561,N_12873,N_12984);
or U13562 (N_13562,N_12792,N_12791);
xor U13563 (N_13563,N_13003,N_12857);
or U13564 (N_13564,N_13122,N_13006);
xnor U13565 (N_13565,N_12798,N_12536);
or U13566 (N_13566,N_12701,N_12975);
nor U13567 (N_13567,N_13025,N_12565);
and U13568 (N_13568,N_12850,N_12687);
nand U13569 (N_13569,N_12780,N_13102);
or U13570 (N_13570,N_12881,N_12752);
nand U13571 (N_13571,N_12651,N_12602);
or U13572 (N_13572,N_12958,N_12914);
nor U13573 (N_13573,N_12628,N_12700);
and U13574 (N_13574,N_12982,N_12680);
and U13575 (N_13575,N_12521,N_12758);
nor U13576 (N_13576,N_13037,N_13114);
nor U13577 (N_13577,N_12755,N_12919);
nand U13578 (N_13578,N_12969,N_12851);
nor U13579 (N_13579,N_12970,N_12675);
nor U13580 (N_13580,N_12548,N_12702);
xnor U13581 (N_13581,N_12786,N_12767);
xnor U13582 (N_13582,N_12664,N_12662);
nor U13583 (N_13583,N_12807,N_12514);
xor U13584 (N_13584,N_12675,N_13118);
nand U13585 (N_13585,N_12852,N_12550);
nor U13586 (N_13586,N_13092,N_12819);
xor U13587 (N_13587,N_12785,N_13116);
nand U13588 (N_13588,N_13111,N_12865);
nand U13589 (N_13589,N_13097,N_12690);
or U13590 (N_13590,N_13002,N_12686);
or U13591 (N_13591,N_12747,N_12643);
nor U13592 (N_13592,N_12861,N_12857);
or U13593 (N_13593,N_12759,N_13098);
and U13594 (N_13594,N_12935,N_12654);
or U13595 (N_13595,N_12631,N_13026);
and U13596 (N_13596,N_12687,N_12880);
and U13597 (N_13597,N_12635,N_13063);
or U13598 (N_13598,N_13043,N_12935);
nand U13599 (N_13599,N_12824,N_13065);
or U13600 (N_13600,N_12750,N_12856);
nor U13601 (N_13601,N_13082,N_13051);
xor U13602 (N_13602,N_12952,N_12644);
and U13603 (N_13603,N_12932,N_12755);
or U13604 (N_13604,N_12503,N_13119);
or U13605 (N_13605,N_12536,N_12736);
xor U13606 (N_13606,N_13005,N_12950);
and U13607 (N_13607,N_12562,N_12655);
and U13608 (N_13608,N_12791,N_12703);
and U13609 (N_13609,N_12586,N_12516);
nor U13610 (N_13610,N_13065,N_13068);
nand U13611 (N_13611,N_12938,N_12528);
or U13612 (N_13612,N_12697,N_12574);
nor U13613 (N_13613,N_12652,N_12674);
or U13614 (N_13614,N_12785,N_13051);
nor U13615 (N_13615,N_13099,N_12605);
nor U13616 (N_13616,N_12805,N_12964);
or U13617 (N_13617,N_13070,N_12651);
and U13618 (N_13618,N_12990,N_12860);
or U13619 (N_13619,N_12550,N_12710);
xor U13620 (N_13620,N_13116,N_12831);
or U13621 (N_13621,N_13023,N_12680);
nor U13622 (N_13622,N_12790,N_13067);
xnor U13623 (N_13623,N_12782,N_12697);
nor U13624 (N_13624,N_12507,N_12604);
and U13625 (N_13625,N_12807,N_12720);
or U13626 (N_13626,N_12677,N_12689);
and U13627 (N_13627,N_12753,N_12591);
xnor U13628 (N_13628,N_13026,N_12645);
nand U13629 (N_13629,N_13071,N_12665);
nand U13630 (N_13630,N_12570,N_13065);
nor U13631 (N_13631,N_12504,N_13099);
and U13632 (N_13632,N_12859,N_12842);
nand U13633 (N_13633,N_12537,N_12784);
and U13634 (N_13634,N_12517,N_12532);
xor U13635 (N_13635,N_12801,N_12711);
and U13636 (N_13636,N_12841,N_12726);
and U13637 (N_13637,N_12984,N_12535);
xor U13638 (N_13638,N_12870,N_12614);
xor U13639 (N_13639,N_12638,N_13018);
and U13640 (N_13640,N_13009,N_12704);
or U13641 (N_13641,N_12926,N_12875);
xor U13642 (N_13642,N_12861,N_12902);
nand U13643 (N_13643,N_12874,N_13086);
nand U13644 (N_13644,N_13069,N_12635);
nand U13645 (N_13645,N_12650,N_12563);
and U13646 (N_13646,N_12705,N_12972);
nor U13647 (N_13647,N_12941,N_12614);
or U13648 (N_13648,N_12697,N_13095);
and U13649 (N_13649,N_12513,N_12799);
and U13650 (N_13650,N_12869,N_12585);
and U13651 (N_13651,N_12967,N_12706);
and U13652 (N_13652,N_13104,N_12731);
and U13653 (N_13653,N_12898,N_12960);
or U13654 (N_13654,N_12897,N_12837);
xnor U13655 (N_13655,N_12757,N_12908);
xnor U13656 (N_13656,N_12787,N_12881);
or U13657 (N_13657,N_12686,N_13066);
nor U13658 (N_13658,N_12649,N_13007);
nor U13659 (N_13659,N_12755,N_12510);
and U13660 (N_13660,N_12533,N_12804);
xnor U13661 (N_13661,N_12995,N_13106);
xnor U13662 (N_13662,N_12671,N_12652);
nand U13663 (N_13663,N_12605,N_12806);
and U13664 (N_13664,N_12675,N_12595);
and U13665 (N_13665,N_12858,N_12559);
or U13666 (N_13666,N_13101,N_12898);
or U13667 (N_13667,N_13109,N_12589);
or U13668 (N_13668,N_12614,N_13031);
nor U13669 (N_13669,N_12698,N_12526);
xnor U13670 (N_13670,N_13073,N_12853);
or U13671 (N_13671,N_13038,N_12960);
xor U13672 (N_13672,N_12764,N_12786);
xor U13673 (N_13673,N_12843,N_12875);
and U13674 (N_13674,N_13084,N_12928);
nor U13675 (N_13675,N_12820,N_12743);
nor U13676 (N_13676,N_12564,N_12738);
nor U13677 (N_13677,N_12879,N_12983);
or U13678 (N_13678,N_12559,N_12944);
nand U13679 (N_13679,N_12787,N_12524);
xnor U13680 (N_13680,N_12595,N_12894);
nor U13681 (N_13681,N_12561,N_12625);
and U13682 (N_13682,N_12663,N_13060);
nor U13683 (N_13683,N_13102,N_12572);
nor U13684 (N_13684,N_12743,N_12602);
xor U13685 (N_13685,N_13020,N_13098);
nand U13686 (N_13686,N_12655,N_12781);
and U13687 (N_13687,N_12646,N_12803);
nor U13688 (N_13688,N_13008,N_12921);
nor U13689 (N_13689,N_13014,N_13031);
xnor U13690 (N_13690,N_12850,N_12669);
and U13691 (N_13691,N_13058,N_12739);
nor U13692 (N_13692,N_12592,N_12973);
and U13693 (N_13693,N_12977,N_12998);
nor U13694 (N_13694,N_12830,N_12720);
nand U13695 (N_13695,N_12552,N_13120);
nor U13696 (N_13696,N_12999,N_12815);
nand U13697 (N_13697,N_13006,N_12990);
xor U13698 (N_13698,N_12608,N_12968);
and U13699 (N_13699,N_12560,N_12781);
nand U13700 (N_13700,N_12531,N_12826);
or U13701 (N_13701,N_12888,N_12870);
and U13702 (N_13702,N_13071,N_12633);
nand U13703 (N_13703,N_13033,N_12789);
nand U13704 (N_13704,N_12548,N_12977);
xor U13705 (N_13705,N_12867,N_12603);
or U13706 (N_13706,N_13014,N_12616);
nand U13707 (N_13707,N_12834,N_12505);
and U13708 (N_13708,N_12665,N_12620);
or U13709 (N_13709,N_12677,N_12554);
or U13710 (N_13710,N_13024,N_13070);
xnor U13711 (N_13711,N_12749,N_12708);
and U13712 (N_13712,N_12598,N_12679);
and U13713 (N_13713,N_12834,N_13063);
nor U13714 (N_13714,N_12669,N_12694);
or U13715 (N_13715,N_12886,N_12935);
and U13716 (N_13716,N_12851,N_12761);
xor U13717 (N_13717,N_12510,N_12842);
nand U13718 (N_13718,N_12728,N_12637);
xor U13719 (N_13719,N_12500,N_12675);
nor U13720 (N_13720,N_13069,N_12544);
nand U13721 (N_13721,N_12560,N_12518);
nand U13722 (N_13722,N_12582,N_12990);
xnor U13723 (N_13723,N_12886,N_13062);
xnor U13724 (N_13724,N_13111,N_12742);
nor U13725 (N_13725,N_12953,N_12928);
or U13726 (N_13726,N_12500,N_12887);
xnor U13727 (N_13727,N_12572,N_12681);
nand U13728 (N_13728,N_12983,N_13106);
nor U13729 (N_13729,N_12679,N_12906);
nor U13730 (N_13730,N_12856,N_12596);
and U13731 (N_13731,N_12663,N_12905);
nand U13732 (N_13732,N_12772,N_12925);
nor U13733 (N_13733,N_12749,N_13108);
nor U13734 (N_13734,N_12700,N_13052);
nor U13735 (N_13735,N_13063,N_12764);
or U13736 (N_13736,N_12828,N_12861);
nor U13737 (N_13737,N_12815,N_12597);
xnor U13738 (N_13738,N_13072,N_13071);
xor U13739 (N_13739,N_13084,N_12966);
nand U13740 (N_13740,N_13052,N_12543);
nand U13741 (N_13741,N_12978,N_12599);
nand U13742 (N_13742,N_12519,N_12803);
or U13743 (N_13743,N_12610,N_13057);
nor U13744 (N_13744,N_12659,N_12894);
nand U13745 (N_13745,N_12872,N_12624);
and U13746 (N_13746,N_12710,N_12828);
nand U13747 (N_13747,N_12585,N_12738);
nor U13748 (N_13748,N_13061,N_12751);
nor U13749 (N_13749,N_12701,N_13031);
nand U13750 (N_13750,N_13705,N_13246);
and U13751 (N_13751,N_13180,N_13307);
and U13752 (N_13752,N_13135,N_13494);
xnor U13753 (N_13753,N_13143,N_13410);
or U13754 (N_13754,N_13161,N_13546);
xor U13755 (N_13755,N_13679,N_13181);
or U13756 (N_13756,N_13346,N_13305);
nor U13757 (N_13757,N_13235,N_13518);
or U13758 (N_13758,N_13170,N_13262);
nor U13759 (N_13759,N_13236,N_13298);
xnor U13760 (N_13760,N_13209,N_13684);
nor U13761 (N_13761,N_13535,N_13357);
xor U13762 (N_13762,N_13444,N_13403);
nand U13763 (N_13763,N_13664,N_13304);
or U13764 (N_13764,N_13147,N_13282);
nor U13765 (N_13765,N_13211,N_13730);
or U13766 (N_13766,N_13738,N_13476);
and U13767 (N_13767,N_13436,N_13416);
xor U13768 (N_13768,N_13432,N_13640);
xor U13769 (N_13769,N_13643,N_13258);
nor U13770 (N_13770,N_13712,N_13396);
nor U13771 (N_13771,N_13573,N_13361);
nand U13772 (N_13772,N_13478,N_13302);
nand U13773 (N_13773,N_13136,N_13187);
or U13774 (N_13774,N_13690,N_13253);
or U13775 (N_13775,N_13454,N_13184);
or U13776 (N_13776,N_13356,N_13353);
nand U13777 (N_13777,N_13537,N_13744);
nor U13778 (N_13778,N_13565,N_13313);
nor U13779 (N_13779,N_13425,N_13237);
xnor U13780 (N_13780,N_13188,N_13580);
nand U13781 (N_13781,N_13477,N_13658);
xor U13782 (N_13782,N_13651,N_13501);
nand U13783 (N_13783,N_13192,N_13467);
nand U13784 (N_13784,N_13491,N_13201);
xor U13785 (N_13785,N_13665,N_13322);
nor U13786 (N_13786,N_13391,N_13232);
and U13787 (N_13787,N_13171,N_13626);
xnor U13788 (N_13788,N_13141,N_13153);
or U13789 (N_13789,N_13214,N_13610);
nor U13790 (N_13790,N_13614,N_13321);
nor U13791 (N_13791,N_13548,N_13320);
nor U13792 (N_13792,N_13554,N_13149);
nand U13793 (N_13793,N_13281,N_13492);
nand U13794 (N_13794,N_13578,N_13677);
nand U13795 (N_13795,N_13166,N_13725);
xnor U13796 (N_13796,N_13452,N_13287);
and U13797 (N_13797,N_13351,N_13566);
or U13798 (N_13798,N_13631,N_13680);
xor U13799 (N_13799,N_13504,N_13230);
xor U13800 (N_13800,N_13132,N_13398);
or U13801 (N_13801,N_13222,N_13486);
and U13802 (N_13802,N_13389,N_13433);
or U13803 (N_13803,N_13303,N_13524);
xor U13804 (N_13804,N_13649,N_13641);
nand U13805 (N_13805,N_13700,N_13577);
and U13806 (N_13806,N_13148,N_13646);
xor U13807 (N_13807,N_13688,N_13526);
xnor U13808 (N_13808,N_13194,N_13458);
and U13809 (N_13809,N_13370,N_13190);
or U13810 (N_13810,N_13411,N_13508);
and U13811 (N_13811,N_13707,N_13460);
or U13812 (N_13812,N_13251,N_13638);
nand U13813 (N_13813,N_13393,N_13428);
nor U13814 (N_13814,N_13423,N_13159);
or U13815 (N_13815,N_13715,N_13269);
and U13816 (N_13816,N_13395,N_13582);
and U13817 (N_13817,N_13341,N_13365);
nor U13818 (N_13818,N_13552,N_13364);
xnor U13819 (N_13819,N_13203,N_13556);
nand U13820 (N_13820,N_13593,N_13613);
nor U13821 (N_13821,N_13719,N_13709);
nor U13822 (N_13822,N_13291,N_13366);
and U13823 (N_13823,N_13496,N_13420);
or U13824 (N_13824,N_13345,N_13482);
and U13825 (N_13825,N_13157,N_13331);
and U13826 (N_13826,N_13511,N_13602);
xnor U13827 (N_13827,N_13134,N_13290);
and U13828 (N_13828,N_13256,N_13284);
nand U13829 (N_13829,N_13318,N_13129);
xnor U13830 (N_13830,N_13668,N_13481);
xnor U13831 (N_13831,N_13238,N_13131);
nand U13832 (N_13832,N_13430,N_13301);
and U13833 (N_13833,N_13446,N_13337);
xnor U13834 (N_13834,N_13274,N_13294);
and U13835 (N_13835,N_13673,N_13563);
nor U13836 (N_13836,N_13158,N_13348);
nand U13837 (N_13837,N_13419,N_13133);
or U13838 (N_13838,N_13463,N_13590);
xor U13839 (N_13839,N_13193,N_13650);
or U13840 (N_13840,N_13470,N_13245);
and U13841 (N_13841,N_13404,N_13354);
or U13842 (N_13842,N_13160,N_13126);
nor U13843 (N_13843,N_13344,N_13599);
and U13844 (N_13844,N_13571,N_13451);
and U13845 (N_13845,N_13666,N_13178);
nand U13846 (N_13846,N_13234,N_13384);
nand U13847 (N_13847,N_13621,N_13415);
nand U13848 (N_13848,N_13182,N_13579);
or U13849 (N_13849,N_13311,N_13721);
nand U13850 (N_13850,N_13377,N_13739);
nor U13851 (N_13851,N_13561,N_13567);
nor U13852 (N_13852,N_13695,N_13408);
nand U13853 (N_13853,N_13375,N_13340);
and U13854 (N_13854,N_13600,N_13551);
or U13855 (N_13855,N_13264,N_13630);
and U13856 (N_13856,N_13442,N_13441);
xor U13857 (N_13857,N_13516,N_13227);
or U13858 (N_13858,N_13314,N_13701);
xnor U13859 (N_13859,N_13588,N_13474);
or U13860 (N_13860,N_13150,N_13286);
and U13861 (N_13861,N_13713,N_13468);
and U13862 (N_13862,N_13620,N_13402);
and U13863 (N_13863,N_13603,N_13597);
nand U13864 (N_13864,N_13417,N_13449);
nor U13865 (N_13865,N_13622,N_13268);
xor U13866 (N_13866,N_13542,N_13525);
nand U13867 (N_13867,N_13270,N_13689);
and U13868 (N_13868,N_13198,N_13362);
nand U13869 (N_13869,N_13448,N_13392);
nand U13870 (N_13870,N_13239,N_13595);
nand U13871 (N_13871,N_13657,N_13257);
nand U13872 (N_13872,N_13529,N_13670);
nor U13873 (N_13873,N_13197,N_13685);
nand U13874 (N_13874,N_13745,N_13386);
nor U13875 (N_13875,N_13249,N_13706);
or U13876 (N_13876,N_13173,N_13407);
nor U13877 (N_13877,N_13475,N_13659);
xor U13878 (N_13878,N_13255,N_13718);
xor U13879 (N_13879,N_13555,N_13473);
xor U13880 (N_13880,N_13729,N_13265);
and U13881 (N_13881,N_13698,N_13285);
and U13882 (N_13882,N_13326,N_13628);
nand U13883 (N_13883,N_13376,N_13466);
nand U13884 (N_13884,N_13213,N_13488);
or U13885 (N_13885,N_13592,N_13374);
xnor U13886 (N_13886,N_13371,N_13687);
nor U13887 (N_13887,N_13300,N_13164);
nand U13888 (N_13888,N_13342,N_13619);
xnor U13889 (N_13889,N_13560,N_13229);
and U13890 (N_13890,N_13639,N_13167);
or U13891 (N_13891,N_13584,N_13517);
and U13892 (N_13892,N_13733,N_13272);
nand U13893 (N_13893,N_13426,N_13278);
nor U13894 (N_13894,N_13704,N_13710);
or U13895 (N_13895,N_13748,N_13325);
xor U13896 (N_13896,N_13316,N_13210);
nor U13897 (N_13897,N_13692,N_13216);
xor U13898 (N_13898,N_13708,N_13330);
or U13899 (N_13899,N_13735,N_13324);
nor U13900 (N_13900,N_13312,N_13437);
and U13901 (N_13901,N_13233,N_13155);
or U13902 (N_13902,N_13645,N_13472);
xnor U13903 (N_13903,N_13438,N_13280);
or U13904 (N_13904,N_13485,N_13703);
xnor U13905 (N_13905,N_13443,N_13728);
and U13906 (N_13906,N_13623,N_13399);
or U13907 (N_13907,N_13177,N_13225);
xnor U13908 (N_13908,N_13431,N_13352);
nor U13909 (N_13909,N_13202,N_13562);
xnor U13910 (N_13910,N_13372,N_13461);
xor U13911 (N_13911,N_13292,N_13223);
xnor U13912 (N_13912,N_13369,N_13539);
and U13913 (N_13913,N_13746,N_13576);
or U13914 (N_13914,N_13279,N_13145);
or U13915 (N_13915,N_13315,N_13457);
or U13916 (N_13916,N_13534,N_13724);
xor U13917 (N_13917,N_13734,N_13359);
and U13918 (N_13918,N_13711,N_13598);
or U13919 (N_13919,N_13137,N_13189);
xnor U13920 (N_13920,N_13163,N_13140);
xnor U13921 (N_13921,N_13484,N_13221);
xnor U13922 (N_13922,N_13642,N_13168);
and U13923 (N_13923,N_13297,N_13632);
nor U13924 (N_13924,N_13263,N_13726);
and U13925 (N_13925,N_13678,N_13334);
xnor U13926 (N_13926,N_13306,N_13544);
or U13927 (N_13927,N_13681,N_13413);
or U13928 (N_13928,N_13569,N_13655);
xor U13929 (N_13929,N_13741,N_13401);
nand U13930 (N_13930,N_13559,N_13434);
nor U13931 (N_13931,N_13204,N_13379);
nor U13932 (N_13932,N_13347,N_13414);
or U13933 (N_13933,N_13199,N_13328);
nand U13934 (N_13934,N_13549,N_13327);
nand U13935 (N_13935,N_13633,N_13697);
nand U13936 (N_13936,N_13217,N_13388);
nor U13937 (N_13937,N_13228,N_13195);
and U13938 (N_13938,N_13627,N_13509);
or U13939 (N_13939,N_13656,N_13382);
xnor U13940 (N_13940,N_13489,N_13545);
and U13941 (N_13941,N_13506,N_13499);
nand U13942 (N_13942,N_13742,N_13186);
nand U13943 (N_13943,N_13200,N_13536);
and U13944 (N_13944,N_13275,N_13661);
and U13945 (N_13945,N_13338,N_13654);
nand U13946 (N_13946,N_13543,N_13412);
nand U13947 (N_13947,N_13378,N_13462);
xor U13948 (N_13948,N_13702,N_13455);
or U13949 (N_13949,N_13521,N_13266);
or U13950 (N_13950,N_13634,N_13226);
and U13951 (N_13951,N_13146,N_13144);
xnor U13952 (N_13952,N_13717,N_13747);
nand U13953 (N_13953,N_13653,N_13243);
nand U13954 (N_13954,N_13261,N_13125);
nand U13955 (N_13955,N_13605,N_13250);
nand U13956 (N_13956,N_13663,N_13127);
nand U13957 (N_13957,N_13191,N_13240);
nand U13958 (N_13958,N_13740,N_13514);
nand U13959 (N_13959,N_13683,N_13604);
and U13960 (N_13960,N_13349,N_13682);
nand U13961 (N_13961,N_13154,N_13541);
nand U13962 (N_13962,N_13637,N_13616);
or U13963 (N_13963,N_13723,N_13676);
or U13964 (N_13964,N_13380,N_13570);
and U13965 (N_13965,N_13358,N_13368);
nand U13966 (N_13966,N_13727,N_13456);
or U13967 (N_13967,N_13130,N_13714);
or U13968 (N_13968,N_13618,N_13424);
nor U13969 (N_13969,N_13299,N_13156);
xor U13970 (N_13970,N_13520,N_13479);
xnor U13971 (N_13971,N_13471,N_13336);
xnor U13972 (N_13972,N_13502,N_13736);
xnor U13973 (N_13973,N_13553,N_13505);
nor U13974 (N_13974,N_13531,N_13343);
nor U13975 (N_13975,N_13271,N_13667);
xor U13976 (N_13976,N_13293,N_13220);
xnor U13977 (N_13977,N_13648,N_13587);
and U13978 (N_13978,N_13422,N_13179);
and U13979 (N_13979,N_13558,N_13208);
xor U13980 (N_13980,N_13737,N_13174);
xnor U13981 (N_13981,N_13288,N_13215);
or U13982 (N_13982,N_13405,N_13421);
nand U13983 (N_13983,N_13607,N_13267);
or U13984 (N_13984,N_13406,N_13205);
nor U13985 (N_13985,N_13572,N_13373);
nand U13986 (N_13986,N_13276,N_13512);
nor U13987 (N_13987,N_13550,N_13498);
xnor U13988 (N_13988,N_13691,N_13241);
xnor U13989 (N_13989,N_13367,N_13453);
nand U13990 (N_13990,N_13409,N_13629);
nor U13991 (N_13991,N_13647,N_13252);
nor U13992 (N_13992,N_13445,N_13360);
nor U13993 (N_13993,N_13615,N_13635);
or U13994 (N_13994,N_13254,N_13500);
nand U13995 (N_13995,N_13277,N_13686);
and U13996 (N_13996,N_13447,N_13557);
xnor U13997 (N_13997,N_13259,N_13696);
xor U13998 (N_13998,N_13400,N_13247);
and U13999 (N_13999,N_13185,N_13295);
nor U14000 (N_14000,N_13152,N_13139);
nand U14001 (N_14001,N_13749,N_13601);
nand U14002 (N_14002,N_13142,N_13465);
and U14003 (N_14003,N_13716,N_13669);
nand U14004 (N_14004,N_13439,N_13527);
and U14005 (N_14005,N_13617,N_13283);
nor U14006 (N_14006,N_13339,N_13574);
or U14007 (N_14007,N_13260,N_13625);
and U14008 (N_14008,N_13538,N_13497);
nand U14009 (N_14009,N_13459,N_13212);
and U14010 (N_14010,N_13586,N_13672);
or U14011 (N_14011,N_13591,N_13381);
xor U14012 (N_14012,N_13699,N_13487);
and U14013 (N_14013,N_13530,N_13532);
and U14014 (N_14014,N_13289,N_13169);
xor U14015 (N_14015,N_13503,N_13510);
or U14016 (N_14016,N_13540,N_13429);
nor U14017 (N_14017,N_13507,N_13317);
nor U14018 (N_14018,N_13493,N_13469);
nand U14019 (N_14019,N_13693,N_13490);
xnor U14020 (N_14020,N_13652,N_13231);
nand U14021 (N_14021,N_13172,N_13450);
nor U14022 (N_14022,N_13583,N_13218);
or U14023 (N_14023,N_13310,N_13611);
nand U14024 (N_14024,N_13547,N_13660);
nand U14025 (N_14025,N_13513,N_13722);
xnor U14026 (N_14026,N_13355,N_13694);
nand U14027 (N_14027,N_13319,N_13162);
xnor U14028 (N_14028,N_13196,N_13418);
or U14029 (N_14029,N_13464,N_13427);
nor U14030 (N_14030,N_13363,N_13397);
and U14031 (N_14031,N_13440,N_13176);
xor U14032 (N_14032,N_13515,N_13206);
or U14033 (N_14033,N_13522,N_13383);
and U14034 (N_14034,N_13596,N_13350);
nor U14035 (N_14035,N_13732,N_13675);
nand U14036 (N_14036,N_13219,N_13606);
nand U14037 (N_14037,N_13662,N_13308);
or U14038 (N_14038,N_13575,N_13731);
nor U14039 (N_14039,N_13242,N_13483);
nor U14040 (N_14040,N_13296,N_13612);
nand U14041 (N_14041,N_13323,N_13720);
and U14042 (N_14042,N_13394,N_13671);
nor U14043 (N_14043,N_13495,N_13175);
nand U14044 (N_14044,N_13151,N_13387);
nor U14045 (N_14045,N_13568,N_13435);
or U14046 (N_14046,N_13224,N_13309);
and U14047 (N_14047,N_13585,N_13743);
or U14048 (N_14048,N_13138,N_13528);
or U14049 (N_14049,N_13523,N_13332);
or U14050 (N_14050,N_13589,N_13165);
nand U14051 (N_14051,N_13248,N_13183);
and U14052 (N_14052,N_13644,N_13594);
and U14053 (N_14053,N_13608,N_13390);
xor U14054 (N_14054,N_13624,N_13128);
nand U14055 (N_14055,N_13564,N_13533);
and U14056 (N_14056,N_13581,N_13207);
xor U14057 (N_14057,N_13636,N_13333);
or U14058 (N_14058,N_13674,N_13519);
or U14059 (N_14059,N_13329,N_13244);
and U14060 (N_14060,N_13385,N_13480);
xnor U14061 (N_14061,N_13335,N_13273);
nor U14062 (N_14062,N_13609,N_13545);
xnor U14063 (N_14063,N_13437,N_13491);
nand U14064 (N_14064,N_13317,N_13182);
nand U14065 (N_14065,N_13510,N_13423);
and U14066 (N_14066,N_13653,N_13619);
nand U14067 (N_14067,N_13628,N_13645);
or U14068 (N_14068,N_13160,N_13437);
nand U14069 (N_14069,N_13325,N_13152);
or U14070 (N_14070,N_13434,N_13143);
xnor U14071 (N_14071,N_13449,N_13547);
nand U14072 (N_14072,N_13144,N_13356);
xnor U14073 (N_14073,N_13647,N_13340);
or U14074 (N_14074,N_13136,N_13416);
xor U14075 (N_14075,N_13674,N_13345);
nand U14076 (N_14076,N_13351,N_13272);
nand U14077 (N_14077,N_13630,N_13130);
nand U14078 (N_14078,N_13166,N_13330);
xor U14079 (N_14079,N_13275,N_13419);
nor U14080 (N_14080,N_13479,N_13593);
nand U14081 (N_14081,N_13745,N_13143);
and U14082 (N_14082,N_13315,N_13663);
xor U14083 (N_14083,N_13406,N_13633);
nand U14084 (N_14084,N_13502,N_13711);
xor U14085 (N_14085,N_13357,N_13611);
xor U14086 (N_14086,N_13590,N_13250);
xor U14087 (N_14087,N_13689,N_13208);
and U14088 (N_14088,N_13557,N_13201);
and U14089 (N_14089,N_13632,N_13616);
nor U14090 (N_14090,N_13667,N_13167);
nor U14091 (N_14091,N_13589,N_13659);
nand U14092 (N_14092,N_13563,N_13383);
nor U14093 (N_14093,N_13489,N_13716);
nor U14094 (N_14094,N_13208,N_13244);
and U14095 (N_14095,N_13329,N_13235);
xor U14096 (N_14096,N_13344,N_13593);
nor U14097 (N_14097,N_13150,N_13530);
xor U14098 (N_14098,N_13480,N_13174);
nor U14099 (N_14099,N_13680,N_13217);
and U14100 (N_14100,N_13330,N_13319);
and U14101 (N_14101,N_13697,N_13598);
nor U14102 (N_14102,N_13626,N_13340);
nor U14103 (N_14103,N_13206,N_13356);
and U14104 (N_14104,N_13172,N_13625);
nor U14105 (N_14105,N_13563,N_13267);
nand U14106 (N_14106,N_13160,N_13609);
and U14107 (N_14107,N_13403,N_13212);
xor U14108 (N_14108,N_13333,N_13472);
nor U14109 (N_14109,N_13478,N_13181);
nor U14110 (N_14110,N_13687,N_13519);
nor U14111 (N_14111,N_13211,N_13726);
and U14112 (N_14112,N_13147,N_13702);
nor U14113 (N_14113,N_13294,N_13629);
or U14114 (N_14114,N_13296,N_13433);
nor U14115 (N_14115,N_13421,N_13509);
xor U14116 (N_14116,N_13409,N_13459);
or U14117 (N_14117,N_13697,N_13708);
nand U14118 (N_14118,N_13603,N_13653);
nand U14119 (N_14119,N_13698,N_13547);
or U14120 (N_14120,N_13246,N_13321);
xor U14121 (N_14121,N_13207,N_13206);
nand U14122 (N_14122,N_13701,N_13725);
and U14123 (N_14123,N_13450,N_13238);
nand U14124 (N_14124,N_13313,N_13590);
or U14125 (N_14125,N_13223,N_13631);
or U14126 (N_14126,N_13126,N_13573);
and U14127 (N_14127,N_13510,N_13617);
xor U14128 (N_14128,N_13178,N_13272);
and U14129 (N_14129,N_13199,N_13387);
nor U14130 (N_14130,N_13726,N_13486);
and U14131 (N_14131,N_13496,N_13421);
nor U14132 (N_14132,N_13210,N_13441);
nor U14133 (N_14133,N_13430,N_13307);
nand U14134 (N_14134,N_13636,N_13159);
and U14135 (N_14135,N_13140,N_13372);
nor U14136 (N_14136,N_13403,N_13143);
nand U14137 (N_14137,N_13589,N_13573);
nor U14138 (N_14138,N_13595,N_13628);
nand U14139 (N_14139,N_13443,N_13434);
xnor U14140 (N_14140,N_13361,N_13666);
or U14141 (N_14141,N_13310,N_13271);
nor U14142 (N_14142,N_13425,N_13359);
nor U14143 (N_14143,N_13460,N_13375);
nand U14144 (N_14144,N_13350,N_13255);
and U14145 (N_14145,N_13147,N_13546);
nand U14146 (N_14146,N_13501,N_13174);
and U14147 (N_14147,N_13709,N_13515);
xnor U14148 (N_14148,N_13388,N_13140);
xor U14149 (N_14149,N_13586,N_13227);
nand U14150 (N_14150,N_13148,N_13723);
or U14151 (N_14151,N_13599,N_13384);
nor U14152 (N_14152,N_13209,N_13680);
or U14153 (N_14153,N_13737,N_13396);
and U14154 (N_14154,N_13232,N_13649);
nor U14155 (N_14155,N_13420,N_13158);
nor U14156 (N_14156,N_13508,N_13178);
xnor U14157 (N_14157,N_13499,N_13192);
xnor U14158 (N_14158,N_13469,N_13734);
or U14159 (N_14159,N_13515,N_13613);
nand U14160 (N_14160,N_13280,N_13585);
xor U14161 (N_14161,N_13431,N_13550);
xor U14162 (N_14162,N_13730,N_13167);
nand U14163 (N_14163,N_13485,N_13158);
or U14164 (N_14164,N_13735,N_13219);
xor U14165 (N_14165,N_13275,N_13285);
xnor U14166 (N_14166,N_13348,N_13537);
nand U14167 (N_14167,N_13561,N_13651);
nand U14168 (N_14168,N_13454,N_13251);
and U14169 (N_14169,N_13238,N_13213);
nand U14170 (N_14170,N_13596,N_13697);
xnor U14171 (N_14171,N_13710,N_13392);
and U14172 (N_14172,N_13439,N_13683);
xnor U14173 (N_14173,N_13142,N_13256);
or U14174 (N_14174,N_13130,N_13306);
nand U14175 (N_14175,N_13657,N_13401);
or U14176 (N_14176,N_13661,N_13151);
xor U14177 (N_14177,N_13501,N_13719);
and U14178 (N_14178,N_13591,N_13438);
and U14179 (N_14179,N_13471,N_13579);
or U14180 (N_14180,N_13472,N_13730);
or U14181 (N_14181,N_13330,N_13583);
nor U14182 (N_14182,N_13135,N_13225);
nor U14183 (N_14183,N_13299,N_13378);
nand U14184 (N_14184,N_13349,N_13275);
or U14185 (N_14185,N_13160,N_13643);
and U14186 (N_14186,N_13536,N_13145);
nand U14187 (N_14187,N_13470,N_13486);
and U14188 (N_14188,N_13134,N_13321);
nand U14189 (N_14189,N_13219,N_13285);
nor U14190 (N_14190,N_13642,N_13575);
xor U14191 (N_14191,N_13223,N_13303);
and U14192 (N_14192,N_13178,N_13304);
or U14193 (N_14193,N_13212,N_13719);
xnor U14194 (N_14194,N_13171,N_13554);
nor U14195 (N_14195,N_13365,N_13348);
or U14196 (N_14196,N_13234,N_13405);
xor U14197 (N_14197,N_13232,N_13193);
nor U14198 (N_14198,N_13233,N_13681);
nand U14199 (N_14199,N_13543,N_13743);
and U14200 (N_14200,N_13280,N_13482);
or U14201 (N_14201,N_13724,N_13428);
and U14202 (N_14202,N_13564,N_13171);
nor U14203 (N_14203,N_13201,N_13623);
or U14204 (N_14204,N_13697,N_13728);
nor U14205 (N_14205,N_13242,N_13206);
or U14206 (N_14206,N_13540,N_13681);
or U14207 (N_14207,N_13684,N_13519);
and U14208 (N_14208,N_13198,N_13736);
or U14209 (N_14209,N_13560,N_13417);
xor U14210 (N_14210,N_13233,N_13706);
and U14211 (N_14211,N_13469,N_13145);
nor U14212 (N_14212,N_13181,N_13702);
and U14213 (N_14213,N_13505,N_13384);
and U14214 (N_14214,N_13389,N_13352);
nor U14215 (N_14215,N_13480,N_13642);
xor U14216 (N_14216,N_13634,N_13174);
nand U14217 (N_14217,N_13617,N_13425);
xor U14218 (N_14218,N_13266,N_13734);
or U14219 (N_14219,N_13296,N_13393);
xor U14220 (N_14220,N_13660,N_13329);
nor U14221 (N_14221,N_13652,N_13604);
or U14222 (N_14222,N_13688,N_13708);
nand U14223 (N_14223,N_13193,N_13558);
or U14224 (N_14224,N_13577,N_13242);
xnor U14225 (N_14225,N_13331,N_13250);
xor U14226 (N_14226,N_13490,N_13485);
xnor U14227 (N_14227,N_13701,N_13627);
xnor U14228 (N_14228,N_13738,N_13348);
or U14229 (N_14229,N_13299,N_13398);
or U14230 (N_14230,N_13554,N_13129);
and U14231 (N_14231,N_13200,N_13412);
nor U14232 (N_14232,N_13262,N_13421);
nand U14233 (N_14233,N_13228,N_13210);
nor U14234 (N_14234,N_13305,N_13463);
xor U14235 (N_14235,N_13314,N_13641);
and U14236 (N_14236,N_13681,N_13299);
nand U14237 (N_14237,N_13553,N_13265);
and U14238 (N_14238,N_13652,N_13659);
nand U14239 (N_14239,N_13396,N_13157);
nand U14240 (N_14240,N_13231,N_13637);
nand U14241 (N_14241,N_13181,N_13294);
or U14242 (N_14242,N_13472,N_13225);
and U14243 (N_14243,N_13228,N_13702);
nor U14244 (N_14244,N_13578,N_13575);
nor U14245 (N_14245,N_13503,N_13515);
nand U14246 (N_14246,N_13350,N_13338);
nor U14247 (N_14247,N_13473,N_13564);
and U14248 (N_14248,N_13306,N_13479);
and U14249 (N_14249,N_13464,N_13461);
and U14250 (N_14250,N_13600,N_13578);
xor U14251 (N_14251,N_13556,N_13559);
nand U14252 (N_14252,N_13698,N_13591);
xnor U14253 (N_14253,N_13260,N_13502);
xnor U14254 (N_14254,N_13698,N_13595);
xnor U14255 (N_14255,N_13126,N_13623);
and U14256 (N_14256,N_13513,N_13354);
and U14257 (N_14257,N_13504,N_13666);
or U14258 (N_14258,N_13687,N_13679);
nand U14259 (N_14259,N_13275,N_13200);
xor U14260 (N_14260,N_13634,N_13430);
nand U14261 (N_14261,N_13415,N_13617);
nand U14262 (N_14262,N_13621,N_13270);
or U14263 (N_14263,N_13681,N_13716);
xnor U14264 (N_14264,N_13640,N_13161);
nor U14265 (N_14265,N_13251,N_13579);
and U14266 (N_14266,N_13412,N_13403);
or U14267 (N_14267,N_13135,N_13600);
nor U14268 (N_14268,N_13195,N_13643);
nand U14269 (N_14269,N_13664,N_13589);
nand U14270 (N_14270,N_13374,N_13190);
or U14271 (N_14271,N_13696,N_13323);
xnor U14272 (N_14272,N_13135,N_13547);
xor U14273 (N_14273,N_13489,N_13699);
nor U14274 (N_14274,N_13711,N_13562);
nand U14275 (N_14275,N_13331,N_13284);
and U14276 (N_14276,N_13545,N_13166);
nor U14277 (N_14277,N_13323,N_13211);
nor U14278 (N_14278,N_13179,N_13339);
nor U14279 (N_14279,N_13479,N_13365);
xor U14280 (N_14280,N_13150,N_13747);
or U14281 (N_14281,N_13631,N_13399);
and U14282 (N_14282,N_13453,N_13395);
xnor U14283 (N_14283,N_13447,N_13128);
nor U14284 (N_14284,N_13456,N_13564);
xnor U14285 (N_14285,N_13561,N_13716);
nand U14286 (N_14286,N_13483,N_13727);
xor U14287 (N_14287,N_13183,N_13735);
xnor U14288 (N_14288,N_13669,N_13665);
nor U14289 (N_14289,N_13330,N_13189);
and U14290 (N_14290,N_13126,N_13248);
nand U14291 (N_14291,N_13744,N_13432);
nand U14292 (N_14292,N_13402,N_13644);
nor U14293 (N_14293,N_13471,N_13406);
nor U14294 (N_14294,N_13459,N_13429);
nor U14295 (N_14295,N_13369,N_13433);
nand U14296 (N_14296,N_13231,N_13223);
or U14297 (N_14297,N_13406,N_13288);
and U14298 (N_14298,N_13577,N_13456);
nor U14299 (N_14299,N_13612,N_13489);
nor U14300 (N_14300,N_13714,N_13267);
xnor U14301 (N_14301,N_13667,N_13528);
or U14302 (N_14302,N_13684,N_13463);
nor U14303 (N_14303,N_13613,N_13550);
or U14304 (N_14304,N_13235,N_13569);
nand U14305 (N_14305,N_13565,N_13397);
or U14306 (N_14306,N_13585,N_13377);
and U14307 (N_14307,N_13144,N_13208);
nand U14308 (N_14308,N_13551,N_13689);
nor U14309 (N_14309,N_13637,N_13265);
and U14310 (N_14310,N_13520,N_13313);
or U14311 (N_14311,N_13597,N_13561);
nand U14312 (N_14312,N_13213,N_13500);
and U14313 (N_14313,N_13513,N_13252);
xor U14314 (N_14314,N_13193,N_13457);
xor U14315 (N_14315,N_13585,N_13457);
and U14316 (N_14316,N_13678,N_13587);
nor U14317 (N_14317,N_13678,N_13542);
nor U14318 (N_14318,N_13663,N_13541);
xnor U14319 (N_14319,N_13606,N_13411);
and U14320 (N_14320,N_13534,N_13354);
and U14321 (N_14321,N_13620,N_13718);
nor U14322 (N_14322,N_13354,N_13392);
nor U14323 (N_14323,N_13431,N_13594);
and U14324 (N_14324,N_13455,N_13378);
nand U14325 (N_14325,N_13438,N_13286);
or U14326 (N_14326,N_13304,N_13541);
nor U14327 (N_14327,N_13403,N_13593);
and U14328 (N_14328,N_13627,N_13260);
nand U14329 (N_14329,N_13440,N_13499);
nand U14330 (N_14330,N_13175,N_13240);
or U14331 (N_14331,N_13269,N_13516);
nor U14332 (N_14332,N_13553,N_13539);
and U14333 (N_14333,N_13294,N_13345);
nand U14334 (N_14334,N_13658,N_13183);
nor U14335 (N_14335,N_13530,N_13307);
xor U14336 (N_14336,N_13553,N_13475);
or U14337 (N_14337,N_13611,N_13176);
or U14338 (N_14338,N_13697,N_13699);
nand U14339 (N_14339,N_13361,N_13209);
or U14340 (N_14340,N_13191,N_13417);
or U14341 (N_14341,N_13741,N_13180);
nand U14342 (N_14342,N_13671,N_13469);
nor U14343 (N_14343,N_13359,N_13575);
xor U14344 (N_14344,N_13432,N_13334);
nand U14345 (N_14345,N_13216,N_13194);
nand U14346 (N_14346,N_13356,N_13264);
nor U14347 (N_14347,N_13352,N_13726);
nor U14348 (N_14348,N_13234,N_13497);
or U14349 (N_14349,N_13704,N_13676);
xnor U14350 (N_14350,N_13262,N_13232);
xor U14351 (N_14351,N_13382,N_13664);
xor U14352 (N_14352,N_13284,N_13678);
and U14353 (N_14353,N_13359,N_13303);
or U14354 (N_14354,N_13711,N_13621);
xor U14355 (N_14355,N_13650,N_13303);
and U14356 (N_14356,N_13137,N_13734);
and U14357 (N_14357,N_13580,N_13545);
nand U14358 (N_14358,N_13655,N_13310);
xor U14359 (N_14359,N_13330,N_13474);
and U14360 (N_14360,N_13650,N_13301);
nand U14361 (N_14361,N_13211,N_13144);
xor U14362 (N_14362,N_13677,N_13169);
nor U14363 (N_14363,N_13599,N_13666);
nand U14364 (N_14364,N_13611,N_13649);
and U14365 (N_14365,N_13719,N_13253);
nand U14366 (N_14366,N_13523,N_13127);
xnor U14367 (N_14367,N_13420,N_13276);
nor U14368 (N_14368,N_13663,N_13358);
or U14369 (N_14369,N_13551,N_13666);
nand U14370 (N_14370,N_13342,N_13195);
nand U14371 (N_14371,N_13154,N_13634);
and U14372 (N_14372,N_13515,N_13184);
nand U14373 (N_14373,N_13309,N_13265);
and U14374 (N_14374,N_13129,N_13357);
nor U14375 (N_14375,N_14276,N_13760);
nor U14376 (N_14376,N_14113,N_13796);
or U14377 (N_14377,N_14190,N_13765);
nor U14378 (N_14378,N_13787,N_13935);
nor U14379 (N_14379,N_13945,N_13984);
nand U14380 (N_14380,N_14289,N_14092);
nand U14381 (N_14381,N_14286,N_13978);
or U14382 (N_14382,N_13847,N_14258);
xor U14383 (N_14383,N_14325,N_14212);
nor U14384 (N_14384,N_14341,N_14326);
and U14385 (N_14385,N_14089,N_14226);
nand U14386 (N_14386,N_13975,N_14310);
and U14387 (N_14387,N_14315,N_14227);
nand U14388 (N_14388,N_13986,N_14231);
nand U14389 (N_14389,N_14008,N_13805);
and U14390 (N_14390,N_14120,N_14003);
nor U14391 (N_14391,N_14211,N_14216);
nor U14392 (N_14392,N_14112,N_13777);
and U14393 (N_14393,N_13970,N_13839);
nor U14394 (N_14394,N_13902,N_14246);
and U14395 (N_14395,N_13816,N_14207);
and U14396 (N_14396,N_13886,N_14343);
nand U14397 (N_14397,N_14232,N_14305);
nand U14398 (N_14398,N_14183,N_14168);
or U14399 (N_14399,N_13987,N_14235);
nor U14400 (N_14400,N_13904,N_14050);
nand U14401 (N_14401,N_14031,N_13927);
nand U14402 (N_14402,N_14060,N_14123);
or U14403 (N_14403,N_14108,N_14063);
nor U14404 (N_14404,N_14057,N_14161);
nand U14405 (N_14405,N_13890,N_13813);
or U14406 (N_14406,N_14138,N_14115);
or U14407 (N_14407,N_14275,N_14155);
nor U14408 (N_14408,N_14223,N_14094);
and U14409 (N_14409,N_13939,N_14082);
nor U14410 (N_14410,N_14051,N_13963);
or U14411 (N_14411,N_14015,N_14293);
xnor U14412 (N_14412,N_13782,N_14011);
xnor U14413 (N_14413,N_14323,N_13942);
xor U14414 (N_14414,N_14032,N_13922);
and U14415 (N_14415,N_13947,N_14164);
or U14416 (N_14416,N_14070,N_14300);
nand U14417 (N_14417,N_14002,N_14218);
xnor U14418 (N_14418,N_14023,N_13926);
nor U14419 (N_14419,N_13916,N_13982);
xor U14420 (N_14420,N_14364,N_13844);
and U14421 (N_14421,N_13775,N_14171);
nand U14422 (N_14422,N_14154,N_13812);
xnor U14423 (N_14423,N_14283,N_13780);
nor U14424 (N_14424,N_13951,N_14318);
nand U14425 (N_14425,N_14121,N_13857);
nand U14426 (N_14426,N_13856,N_13894);
xor U14427 (N_14427,N_14345,N_13799);
xnor U14428 (N_14428,N_14087,N_14206);
nor U14429 (N_14429,N_13818,N_13759);
and U14430 (N_14430,N_14105,N_14312);
xnor U14431 (N_14431,N_13983,N_14137);
or U14432 (N_14432,N_13924,N_14109);
or U14433 (N_14433,N_13852,N_14146);
or U14434 (N_14434,N_13851,N_14142);
or U14435 (N_14435,N_14198,N_13993);
or U14436 (N_14436,N_14321,N_13838);
nand U14437 (N_14437,N_14119,N_13898);
nand U14438 (N_14438,N_13825,N_13815);
xor U14439 (N_14439,N_14254,N_13908);
or U14440 (N_14440,N_14176,N_14238);
or U14441 (N_14441,N_14337,N_14157);
xor U14442 (N_14442,N_14030,N_13944);
nand U14443 (N_14443,N_13881,N_13776);
nor U14444 (N_14444,N_14044,N_14361);
or U14445 (N_14445,N_14222,N_13961);
and U14446 (N_14446,N_13871,N_13814);
nor U14447 (N_14447,N_14065,N_14225);
and U14448 (N_14448,N_13974,N_13959);
and U14449 (N_14449,N_13784,N_13912);
and U14450 (N_14450,N_14111,N_13899);
xor U14451 (N_14451,N_14193,N_13973);
and U14452 (N_14452,N_13964,N_14165);
or U14453 (N_14453,N_14219,N_14340);
xor U14454 (N_14454,N_14103,N_13948);
nand U14455 (N_14455,N_14072,N_14230);
xnor U14456 (N_14456,N_14097,N_13958);
or U14457 (N_14457,N_13845,N_14224);
nor U14458 (N_14458,N_14195,N_14314);
and U14459 (N_14459,N_13761,N_14149);
or U14460 (N_14460,N_13867,N_13907);
and U14461 (N_14461,N_13891,N_14124);
nor U14462 (N_14462,N_14181,N_13833);
nand U14463 (N_14463,N_14253,N_13981);
and U14464 (N_14464,N_14369,N_14255);
xor U14465 (N_14465,N_14152,N_14324);
xnor U14466 (N_14466,N_14180,N_14129);
and U14467 (N_14467,N_14288,N_13909);
xor U14468 (N_14468,N_14203,N_14153);
xnor U14469 (N_14469,N_13929,N_14029);
nand U14470 (N_14470,N_14292,N_14042);
and U14471 (N_14471,N_13794,N_13795);
and U14472 (N_14472,N_13992,N_14160);
or U14473 (N_14473,N_14143,N_13769);
and U14474 (N_14474,N_14177,N_13877);
or U14475 (N_14475,N_14052,N_13883);
and U14476 (N_14476,N_13789,N_14248);
xor U14477 (N_14477,N_14173,N_14294);
and U14478 (N_14478,N_14162,N_14067);
or U14479 (N_14479,N_14304,N_14132);
nand U14480 (N_14480,N_14273,N_14004);
xnor U14481 (N_14481,N_13868,N_14217);
nand U14482 (N_14482,N_13837,N_13917);
nand U14483 (N_14483,N_14045,N_13788);
and U14484 (N_14484,N_14297,N_13785);
xnor U14485 (N_14485,N_14352,N_14351);
xnor U14486 (N_14486,N_14236,N_13893);
nand U14487 (N_14487,N_13937,N_13905);
or U14488 (N_14488,N_14291,N_13832);
xnor U14489 (N_14489,N_13864,N_14259);
nor U14490 (N_14490,N_13800,N_13870);
and U14491 (N_14491,N_13878,N_14266);
and U14492 (N_14492,N_13820,N_14139);
nor U14493 (N_14493,N_14041,N_14018);
or U14494 (N_14494,N_14281,N_14038);
or U14495 (N_14495,N_14362,N_14090);
or U14496 (N_14496,N_14241,N_14338);
and U14497 (N_14497,N_13807,N_14141);
nor U14498 (N_14498,N_14037,N_14339);
nand U14499 (N_14499,N_14064,N_14167);
or U14500 (N_14500,N_14010,N_14301);
nor U14501 (N_14501,N_13873,N_14194);
nor U14502 (N_14502,N_14075,N_13758);
or U14503 (N_14503,N_14012,N_14163);
nand U14504 (N_14504,N_13779,N_14006);
nor U14505 (N_14505,N_14200,N_14117);
or U14506 (N_14506,N_14184,N_13919);
nor U14507 (N_14507,N_13941,N_14130);
nor U14508 (N_14508,N_14335,N_13778);
nand U14509 (N_14509,N_13849,N_14122);
nand U14510 (N_14510,N_14019,N_14332);
nand U14511 (N_14511,N_14001,N_13914);
and U14512 (N_14512,N_13854,N_14144);
xor U14513 (N_14513,N_13766,N_14192);
nand U14514 (N_14514,N_13876,N_13827);
or U14515 (N_14515,N_13888,N_14069);
and U14516 (N_14516,N_13753,N_14363);
or U14517 (N_14517,N_14150,N_13985);
nor U14518 (N_14518,N_13930,N_14210);
xor U14519 (N_14519,N_13892,N_13921);
or U14520 (N_14520,N_14342,N_13969);
and U14521 (N_14521,N_13841,N_14213);
nor U14522 (N_14522,N_13882,N_14368);
nand U14523 (N_14523,N_14147,N_14020);
and U14524 (N_14524,N_14280,N_13910);
and U14525 (N_14525,N_14228,N_13853);
xnor U14526 (N_14526,N_14178,N_14056);
and U14527 (N_14527,N_13806,N_13804);
and U14528 (N_14528,N_13936,N_13762);
nor U14529 (N_14529,N_14265,N_13829);
xor U14530 (N_14530,N_14360,N_14093);
nand U14531 (N_14531,N_14202,N_13858);
and U14532 (N_14532,N_14262,N_14270);
and U14533 (N_14533,N_14017,N_13798);
or U14534 (N_14534,N_13925,N_14073);
and U14535 (N_14535,N_13931,N_14214);
nor U14536 (N_14536,N_14024,N_14048);
nand U14537 (N_14537,N_14188,N_13783);
nor U14538 (N_14538,N_14347,N_14196);
or U14539 (N_14539,N_14096,N_14025);
nor U14540 (N_14540,N_14009,N_13950);
or U14541 (N_14541,N_14327,N_14336);
nand U14542 (N_14542,N_13932,N_14085);
nor U14543 (N_14543,N_14302,N_14296);
and U14544 (N_14544,N_13906,N_13770);
and U14545 (N_14545,N_13808,N_13980);
xor U14546 (N_14546,N_14243,N_13880);
and U14547 (N_14547,N_13957,N_14014);
xnor U14548 (N_14548,N_14058,N_14267);
or U14549 (N_14549,N_14088,N_14035);
or U14550 (N_14550,N_14140,N_14328);
nor U14551 (N_14551,N_14016,N_14229);
or U14552 (N_14552,N_13962,N_13866);
nor U14553 (N_14553,N_13928,N_14174);
and U14554 (N_14554,N_14319,N_13819);
or U14555 (N_14555,N_14242,N_13771);
and U14556 (N_14556,N_13911,N_13822);
nor U14557 (N_14557,N_14099,N_14299);
xnor U14558 (N_14558,N_14322,N_14274);
nor U14559 (N_14559,N_14106,N_13920);
nand U14560 (N_14560,N_14354,N_14040);
xor U14561 (N_14561,N_14145,N_14127);
or U14562 (N_14562,N_14049,N_14366);
nor U14563 (N_14563,N_14128,N_14077);
nand U14564 (N_14564,N_13817,N_14131);
nor U14565 (N_14565,N_14239,N_14237);
or U14566 (N_14566,N_14197,N_13843);
or U14567 (N_14567,N_14187,N_14007);
nor U14568 (N_14568,N_13767,N_14205);
nand U14569 (N_14569,N_13752,N_14148);
and U14570 (N_14570,N_14027,N_14133);
xor U14571 (N_14571,N_13952,N_13850);
xor U14572 (N_14572,N_14334,N_14320);
xnor U14573 (N_14573,N_14136,N_13934);
or U14574 (N_14574,N_13996,N_14272);
nor U14575 (N_14575,N_13913,N_14028);
xor U14576 (N_14576,N_13938,N_13979);
xor U14577 (N_14577,N_13810,N_13768);
nor U14578 (N_14578,N_14250,N_14329);
nor U14579 (N_14579,N_14185,N_14126);
xnor U14580 (N_14580,N_14370,N_13802);
or U14581 (N_14581,N_13988,N_14282);
nand U14582 (N_14582,N_14344,N_13887);
nor U14583 (N_14583,N_14373,N_14251);
xnor U14584 (N_14584,N_14348,N_13828);
or U14585 (N_14585,N_14220,N_14083);
and U14586 (N_14586,N_14252,N_13903);
or U14587 (N_14587,N_13772,N_13790);
or U14588 (N_14588,N_13956,N_14054);
and U14589 (N_14589,N_13823,N_13781);
nand U14590 (N_14590,N_14079,N_13791);
and U14591 (N_14591,N_13757,N_14022);
nand U14592 (N_14592,N_14257,N_13995);
and U14593 (N_14593,N_13879,N_14278);
nor U14594 (N_14594,N_14039,N_14084);
nor U14595 (N_14595,N_13896,N_14268);
nor U14596 (N_14596,N_14234,N_14261);
nand U14597 (N_14597,N_14201,N_14316);
xnor U14598 (N_14598,N_14175,N_13989);
and U14599 (N_14599,N_13859,N_14271);
nand U14600 (N_14600,N_13889,N_14371);
and U14601 (N_14601,N_14365,N_14172);
and U14602 (N_14602,N_14215,N_14086);
nor U14603 (N_14603,N_13809,N_13863);
nor U14604 (N_14604,N_14306,N_14313);
and U14605 (N_14605,N_14374,N_14247);
xor U14606 (N_14606,N_14071,N_13834);
and U14607 (N_14607,N_13940,N_14043);
xnor U14608 (N_14608,N_13786,N_14118);
nand U14609 (N_14609,N_14331,N_14182);
nand U14610 (N_14610,N_14298,N_13865);
xnor U14611 (N_14611,N_14100,N_13860);
nand U14612 (N_14612,N_13835,N_13764);
nand U14613 (N_14613,N_14053,N_14284);
or U14614 (N_14614,N_14279,N_14066);
xor U14615 (N_14615,N_13971,N_13830);
nand U14616 (N_14616,N_13793,N_14036);
xor U14617 (N_14617,N_13756,N_13831);
or U14618 (N_14618,N_14159,N_13994);
or U14619 (N_14619,N_13965,N_14134);
xor U14620 (N_14620,N_14191,N_14204);
and U14621 (N_14621,N_14104,N_14333);
nand U14622 (N_14622,N_14151,N_14367);
or U14623 (N_14623,N_13897,N_14156);
nor U14624 (N_14624,N_14353,N_13869);
xor U14625 (N_14625,N_14372,N_14356);
nand U14626 (N_14626,N_14033,N_13842);
xnor U14627 (N_14627,N_14055,N_14021);
xnor U14628 (N_14628,N_14078,N_13773);
nand U14629 (N_14629,N_13977,N_14260);
and U14630 (N_14630,N_13923,N_13763);
or U14631 (N_14631,N_13955,N_14080);
xor U14632 (N_14632,N_14026,N_13953);
or U14633 (N_14633,N_13821,N_13885);
or U14634 (N_14634,N_14287,N_14034);
and U14635 (N_14635,N_14199,N_13751);
or U14636 (N_14636,N_13990,N_13933);
xor U14637 (N_14637,N_13874,N_13755);
nor U14638 (N_14638,N_14308,N_13855);
or U14639 (N_14639,N_14269,N_14303);
xor U14640 (N_14640,N_14076,N_13901);
xor U14641 (N_14641,N_14061,N_13918);
or U14642 (N_14642,N_13895,N_13915);
nand U14643 (N_14643,N_14098,N_13861);
or U14644 (N_14644,N_14135,N_14062);
xor U14645 (N_14645,N_13797,N_14166);
or U14646 (N_14646,N_14114,N_13872);
or U14647 (N_14647,N_13875,N_14233);
nand U14648 (N_14648,N_14101,N_14189);
or U14649 (N_14649,N_14209,N_14221);
nor U14650 (N_14650,N_13972,N_13954);
nand U14651 (N_14651,N_14047,N_13998);
nor U14652 (N_14652,N_13750,N_13824);
nand U14653 (N_14653,N_14081,N_14091);
or U14654 (N_14654,N_13946,N_13884);
and U14655 (N_14655,N_13801,N_14095);
and U14656 (N_14656,N_14158,N_14330);
or U14657 (N_14657,N_13966,N_14240);
and U14658 (N_14658,N_14102,N_14295);
and U14659 (N_14659,N_13997,N_14359);
or U14660 (N_14660,N_13968,N_14170);
and U14661 (N_14661,N_14307,N_14046);
and U14662 (N_14662,N_13976,N_13949);
nor U14663 (N_14663,N_14059,N_14311);
nor U14664 (N_14664,N_13754,N_13803);
xor U14665 (N_14665,N_14116,N_13811);
and U14666 (N_14666,N_14256,N_13999);
xor U14667 (N_14667,N_14358,N_14355);
or U14668 (N_14668,N_14277,N_13991);
xor U14669 (N_14669,N_14350,N_14346);
and U14670 (N_14670,N_13967,N_14208);
nand U14671 (N_14671,N_14074,N_13836);
xor U14672 (N_14672,N_14245,N_14349);
nor U14673 (N_14673,N_14264,N_14179);
or U14674 (N_14674,N_14357,N_13862);
nand U14675 (N_14675,N_14186,N_13943);
nor U14676 (N_14676,N_13900,N_14068);
nor U14677 (N_14677,N_14244,N_14005);
nand U14678 (N_14678,N_14263,N_13792);
nor U14679 (N_14679,N_14107,N_14110);
or U14680 (N_14680,N_14309,N_13960);
xnor U14681 (N_14681,N_13840,N_13774);
xnor U14682 (N_14682,N_14285,N_13848);
nand U14683 (N_14683,N_14013,N_14249);
xnor U14684 (N_14684,N_14000,N_14169);
xnor U14685 (N_14685,N_13826,N_13846);
xor U14686 (N_14686,N_14290,N_14125);
nand U14687 (N_14687,N_14317,N_13980);
nor U14688 (N_14688,N_14057,N_14160);
or U14689 (N_14689,N_13861,N_14190);
nor U14690 (N_14690,N_14286,N_14290);
nand U14691 (N_14691,N_13800,N_14235);
nand U14692 (N_14692,N_14323,N_14129);
or U14693 (N_14693,N_13791,N_14074);
xor U14694 (N_14694,N_13964,N_14362);
xor U14695 (N_14695,N_14142,N_14309);
and U14696 (N_14696,N_14018,N_14017);
and U14697 (N_14697,N_14089,N_14309);
or U14698 (N_14698,N_14097,N_13855);
nand U14699 (N_14699,N_13962,N_13857);
and U14700 (N_14700,N_14171,N_14188);
xor U14701 (N_14701,N_13870,N_13772);
nor U14702 (N_14702,N_14019,N_14034);
nand U14703 (N_14703,N_14164,N_13934);
or U14704 (N_14704,N_14263,N_14116);
nor U14705 (N_14705,N_13961,N_14208);
nor U14706 (N_14706,N_13914,N_13868);
or U14707 (N_14707,N_14012,N_14263);
nand U14708 (N_14708,N_14072,N_14145);
nor U14709 (N_14709,N_13836,N_14179);
xor U14710 (N_14710,N_14329,N_14290);
nor U14711 (N_14711,N_13941,N_14172);
nor U14712 (N_14712,N_14370,N_14037);
nor U14713 (N_14713,N_14365,N_14201);
or U14714 (N_14714,N_14130,N_13849);
nor U14715 (N_14715,N_14142,N_14102);
and U14716 (N_14716,N_13800,N_14091);
or U14717 (N_14717,N_13942,N_13897);
or U14718 (N_14718,N_14000,N_14289);
nand U14719 (N_14719,N_13771,N_13778);
or U14720 (N_14720,N_14236,N_13936);
or U14721 (N_14721,N_14093,N_13809);
nand U14722 (N_14722,N_13856,N_13970);
and U14723 (N_14723,N_14228,N_14188);
and U14724 (N_14724,N_14067,N_14010);
nand U14725 (N_14725,N_13842,N_14195);
nand U14726 (N_14726,N_14115,N_14274);
nor U14727 (N_14727,N_13806,N_14356);
or U14728 (N_14728,N_14066,N_13847);
nor U14729 (N_14729,N_14143,N_13924);
nand U14730 (N_14730,N_14341,N_13865);
or U14731 (N_14731,N_13813,N_13894);
nor U14732 (N_14732,N_14322,N_14230);
and U14733 (N_14733,N_14179,N_14334);
nand U14734 (N_14734,N_14054,N_14347);
nor U14735 (N_14735,N_14176,N_13964);
nor U14736 (N_14736,N_14185,N_14267);
nor U14737 (N_14737,N_14122,N_13970);
nand U14738 (N_14738,N_13836,N_13847);
nor U14739 (N_14739,N_14295,N_14335);
nor U14740 (N_14740,N_14154,N_14366);
nand U14741 (N_14741,N_14283,N_14032);
and U14742 (N_14742,N_14071,N_14350);
or U14743 (N_14743,N_14115,N_13881);
nor U14744 (N_14744,N_13845,N_14120);
nor U14745 (N_14745,N_14138,N_13897);
nand U14746 (N_14746,N_13985,N_14162);
nor U14747 (N_14747,N_14053,N_13838);
and U14748 (N_14748,N_13994,N_14082);
xnor U14749 (N_14749,N_14265,N_14230);
and U14750 (N_14750,N_14172,N_14031);
nor U14751 (N_14751,N_14246,N_14315);
or U14752 (N_14752,N_14006,N_13888);
xor U14753 (N_14753,N_13780,N_14264);
nor U14754 (N_14754,N_14306,N_14368);
nand U14755 (N_14755,N_14303,N_14244);
nor U14756 (N_14756,N_14193,N_14283);
or U14757 (N_14757,N_14319,N_13960);
nor U14758 (N_14758,N_13862,N_14341);
nand U14759 (N_14759,N_13974,N_13834);
xor U14760 (N_14760,N_13890,N_13896);
and U14761 (N_14761,N_13909,N_13991);
nand U14762 (N_14762,N_14254,N_13808);
xnor U14763 (N_14763,N_13782,N_13827);
xnor U14764 (N_14764,N_14089,N_14373);
xnor U14765 (N_14765,N_13969,N_13944);
nand U14766 (N_14766,N_13805,N_14150);
nand U14767 (N_14767,N_14269,N_13771);
or U14768 (N_14768,N_14315,N_14169);
nor U14769 (N_14769,N_14225,N_14192);
and U14770 (N_14770,N_13782,N_13778);
nor U14771 (N_14771,N_13974,N_14203);
and U14772 (N_14772,N_14206,N_13919);
and U14773 (N_14773,N_14172,N_14167);
xnor U14774 (N_14774,N_13790,N_13814);
or U14775 (N_14775,N_13963,N_13985);
nor U14776 (N_14776,N_13924,N_14249);
and U14777 (N_14777,N_14054,N_14312);
or U14778 (N_14778,N_14181,N_13938);
and U14779 (N_14779,N_13760,N_13955);
and U14780 (N_14780,N_13873,N_13946);
or U14781 (N_14781,N_13897,N_13936);
or U14782 (N_14782,N_14152,N_14343);
and U14783 (N_14783,N_14112,N_14256);
nand U14784 (N_14784,N_14074,N_14269);
nor U14785 (N_14785,N_14263,N_14152);
xor U14786 (N_14786,N_14026,N_14250);
nand U14787 (N_14787,N_13974,N_14158);
xnor U14788 (N_14788,N_13768,N_14296);
nor U14789 (N_14789,N_13786,N_13792);
nand U14790 (N_14790,N_13765,N_14162);
and U14791 (N_14791,N_13831,N_13982);
nand U14792 (N_14792,N_14185,N_13778);
and U14793 (N_14793,N_13854,N_14074);
or U14794 (N_14794,N_14004,N_14216);
xor U14795 (N_14795,N_14045,N_13956);
xnor U14796 (N_14796,N_14253,N_14168);
and U14797 (N_14797,N_13794,N_13900);
nand U14798 (N_14798,N_13778,N_14208);
and U14799 (N_14799,N_14183,N_13897);
or U14800 (N_14800,N_14158,N_14309);
xnor U14801 (N_14801,N_13942,N_14209);
and U14802 (N_14802,N_14062,N_13804);
nor U14803 (N_14803,N_13802,N_14249);
nor U14804 (N_14804,N_14234,N_13791);
xnor U14805 (N_14805,N_14134,N_14350);
and U14806 (N_14806,N_14045,N_13924);
and U14807 (N_14807,N_13859,N_14335);
nor U14808 (N_14808,N_13919,N_13854);
or U14809 (N_14809,N_14068,N_13809);
nor U14810 (N_14810,N_14207,N_14235);
or U14811 (N_14811,N_13759,N_13761);
nand U14812 (N_14812,N_14172,N_13940);
nor U14813 (N_14813,N_14161,N_14203);
nor U14814 (N_14814,N_14007,N_13837);
and U14815 (N_14815,N_14134,N_14001);
and U14816 (N_14816,N_14332,N_13788);
and U14817 (N_14817,N_13903,N_14042);
nand U14818 (N_14818,N_14224,N_14236);
or U14819 (N_14819,N_13822,N_13851);
or U14820 (N_14820,N_13920,N_14320);
nor U14821 (N_14821,N_14202,N_13949);
xnor U14822 (N_14822,N_14118,N_14135);
nor U14823 (N_14823,N_13984,N_13918);
xnor U14824 (N_14824,N_13930,N_14313);
xnor U14825 (N_14825,N_13770,N_14153);
xnor U14826 (N_14826,N_14237,N_14304);
nand U14827 (N_14827,N_14153,N_13905);
nand U14828 (N_14828,N_14018,N_13865);
nand U14829 (N_14829,N_13942,N_13992);
or U14830 (N_14830,N_14080,N_13949);
or U14831 (N_14831,N_14086,N_13996);
nor U14832 (N_14832,N_13788,N_14022);
xnor U14833 (N_14833,N_14137,N_14277);
nand U14834 (N_14834,N_14267,N_13930);
nand U14835 (N_14835,N_14227,N_13927);
xnor U14836 (N_14836,N_13831,N_13896);
or U14837 (N_14837,N_14255,N_13884);
nand U14838 (N_14838,N_14187,N_14297);
or U14839 (N_14839,N_14316,N_13997);
nor U14840 (N_14840,N_14080,N_14251);
xnor U14841 (N_14841,N_13789,N_13940);
and U14842 (N_14842,N_13885,N_14050);
or U14843 (N_14843,N_14293,N_13959);
and U14844 (N_14844,N_13757,N_14236);
nor U14845 (N_14845,N_14316,N_13898);
nor U14846 (N_14846,N_13950,N_13924);
xor U14847 (N_14847,N_14343,N_14211);
or U14848 (N_14848,N_14054,N_14285);
nor U14849 (N_14849,N_14268,N_14148);
nor U14850 (N_14850,N_14369,N_14266);
and U14851 (N_14851,N_14370,N_13902);
nor U14852 (N_14852,N_14023,N_13815);
xor U14853 (N_14853,N_13964,N_13853);
nand U14854 (N_14854,N_14351,N_13855);
nand U14855 (N_14855,N_14362,N_14085);
or U14856 (N_14856,N_14365,N_13847);
and U14857 (N_14857,N_14081,N_14134);
nor U14858 (N_14858,N_13759,N_13993);
nand U14859 (N_14859,N_14319,N_13921);
xor U14860 (N_14860,N_13783,N_13897);
nand U14861 (N_14861,N_13922,N_14145);
and U14862 (N_14862,N_13820,N_13848);
nor U14863 (N_14863,N_13926,N_13945);
nand U14864 (N_14864,N_14069,N_13775);
and U14865 (N_14865,N_14218,N_14154);
xnor U14866 (N_14866,N_14267,N_14150);
xor U14867 (N_14867,N_13805,N_13888);
and U14868 (N_14868,N_14220,N_14306);
or U14869 (N_14869,N_13990,N_14158);
nor U14870 (N_14870,N_14248,N_14076);
or U14871 (N_14871,N_13774,N_14053);
nand U14872 (N_14872,N_13850,N_13972);
nand U14873 (N_14873,N_14074,N_13786);
and U14874 (N_14874,N_14048,N_14135);
nand U14875 (N_14875,N_14268,N_14009);
nand U14876 (N_14876,N_13885,N_13881);
nor U14877 (N_14877,N_13906,N_14134);
and U14878 (N_14878,N_13947,N_14211);
or U14879 (N_14879,N_14340,N_14290);
nand U14880 (N_14880,N_14247,N_14177);
nand U14881 (N_14881,N_13804,N_14217);
and U14882 (N_14882,N_13845,N_14081);
or U14883 (N_14883,N_13955,N_13861);
or U14884 (N_14884,N_13878,N_13898);
or U14885 (N_14885,N_13763,N_13838);
and U14886 (N_14886,N_13937,N_14177);
nand U14887 (N_14887,N_14219,N_13935);
nor U14888 (N_14888,N_13775,N_13944);
nand U14889 (N_14889,N_14180,N_13929);
and U14890 (N_14890,N_14112,N_14062);
nand U14891 (N_14891,N_13861,N_13991);
and U14892 (N_14892,N_14104,N_13993);
nor U14893 (N_14893,N_14341,N_14241);
nor U14894 (N_14894,N_14263,N_13751);
nand U14895 (N_14895,N_14337,N_14076);
and U14896 (N_14896,N_14306,N_13948);
xor U14897 (N_14897,N_14052,N_14092);
nor U14898 (N_14898,N_14041,N_14190);
xnor U14899 (N_14899,N_13991,N_14248);
or U14900 (N_14900,N_14039,N_14234);
xnor U14901 (N_14901,N_13756,N_14065);
and U14902 (N_14902,N_13962,N_13995);
and U14903 (N_14903,N_14093,N_13898);
nor U14904 (N_14904,N_14018,N_14266);
nor U14905 (N_14905,N_13977,N_14234);
or U14906 (N_14906,N_14029,N_13962);
or U14907 (N_14907,N_14127,N_14097);
and U14908 (N_14908,N_13951,N_14203);
nor U14909 (N_14909,N_14132,N_14202);
nor U14910 (N_14910,N_13956,N_13780);
nand U14911 (N_14911,N_14241,N_14292);
xor U14912 (N_14912,N_14301,N_13881);
nor U14913 (N_14913,N_13881,N_14233);
nor U14914 (N_14914,N_13879,N_14354);
and U14915 (N_14915,N_14130,N_13881);
nor U14916 (N_14916,N_14091,N_14051);
xnor U14917 (N_14917,N_14064,N_13750);
xnor U14918 (N_14918,N_14195,N_13755);
or U14919 (N_14919,N_14105,N_14177);
or U14920 (N_14920,N_14015,N_13859);
and U14921 (N_14921,N_13960,N_13967);
or U14922 (N_14922,N_14186,N_14330);
or U14923 (N_14923,N_14352,N_13934);
or U14924 (N_14924,N_14368,N_14335);
xor U14925 (N_14925,N_14058,N_14170);
or U14926 (N_14926,N_14175,N_13754);
and U14927 (N_14927,N_13775,N_13870);
nor U14928 (N_14928,N_14176,N_14091);
nand U14929 (N_14929,N_14031,N_14320);
nand U14930 (N_14930,N_13887,N_13755);
or U14931 (N_14931,N_13945,N_13767);
nor U14932 (N_14932,N_13779,N_13778);
and U14933 (N_14933,N_13758,N_14094);
xor U14934 (N_14934,N_14056,N_13946);
and U14935 (N_14935,N_13922,N_13796);
and U14936 (N_14936,N_14044,N_13909);
or U14937 (N_14937,N_13803,N_14232);
nand U14938 (N_14938,N_14249,N_13925);
and U14939 (N_14939,N_14052,N_14286);
xnor U14940 (N_14940,N_13798,N_14179);
and U14941 (N_14941,N_13801,N_14248);
nor U14942 (N_14942,N_14173,N_13967);
or U14943 (N_14943,N_13983,N_14217);
and U14944 (N_14944,N_14045,N_13965);
nor U14945 (N_14945,N_14300,N_13877);
xnor U14946 (N_14946,N_13956,N_14210);
nand U14947 (N_14947,N_13890,N_13832);
nand U14948 (N_14948,N_13908,N_13999);
nand U14949 (N_14949,N_14210,N_13834);
nor U14950 (N_14950,N_13776,N_14209);
nor U14951 (N_14951,N_13972,N_13951);
and U14952 (N_14952,N_14149,N_13785);
or U14953 (N_14953,N_14371,N_13774);
and U14954 (N_14954,N_14098,N_14257);
nand U14955 (N_14955,N_14059,N_14222);
nor U14956 (N_14956,N_14126,N_13816);
nand U14957 (N_14957,N_13866,N_14024);
xnor U14958 (N_14958,N_13980,N_14040);
nor U14959 (N_14959,N_14337,N_13760);
xor U14960 (N_14960,N_13870,N_14097);
nand U14961 (N_14961,N_14060,N_13928);
nor U14962 (N_14962,N_13988,N_14347);
nand U14963 (N_14963,N_13837,N_13998);
and U14964 (N_14964,N_13804,N_14251);
xor U14965 (N_14965,N_14140,N_14366);
nand U14966 (N_14966,N_14332,N_14299);
nor U14967 (N_14967,N_13809,N_14138);
xor U14968 (N_14968,N_13884,N_14122);
and U14969 (N_14969,N_14054,N_13791);
and U14970 (N_14970,N_14090,N_13872);
and U14971 (N_14971,N_13909,N_14238);
nand U14972 (N_14972,N_14266,N_14343);
nand U14973 (N_14973,N_14359,N_14164);
or U14974 (N_14974,N_14109,N_14139);
or U14975 (N_14975,N_14012,N_13854);
and U14976 (N_14976,N_13833,N_14287);
xor U14977 (N_14977,N_14102,N_14286);
and U14978 (N_14978,N_14337,N_14281);
nor U14979 (N_14979,N_14221,N_14126);
xnor U14980 (N_14980,N_13995,N_14213);
nor U14981 (N_14981,N_14038,N_14123);
xor U14982 (N_14982,N_14259,N_13819);
and U14983 (N_14983,N_14145,N_14133);
or U14984 (N_14984,N_14144,N_14211);
nor U14985 (N_14985,N_14226,N_14330);
nor U14986 (N_14986,N_14046,N_14176);
and U14987 (N_14987,N_14126,N_13896);
nand U14988 (N_14988,N_14066,N_14244);
or U14989 (N_14989,N_14053,N_13928);
nand U14990 (N_14990,N_14320,N_14141);
and U14991 (N_14991,N_13828,N_13820);
or U14992 (N_14992,N_14127,N_14013);
nand U14993 (N_14993,N_14350,N_14295);
and U14994 (N_14994,N_13754,N_14139);
and U14995 (N_14995,N_14016,N_14038);
nand U14996 (N_14996,N_13980,N_14077);
nand U14997 (N_14997,N_14190,N_14312);
xnor U14998 (N_14998,N_14222,N_14211);
or U14999 (N_14999,N_13923,N_13792);
or U15000 (N_15000,N_14546,N_14583);
nand U15001 (N_15001,N_14396,N_14525);
and U15002 (N_15002,N_14906,N_14764);
nor U15003 (N_15003,N_14547,N_14873);
nand U15004 (N_15004,N_14725,N_14457);
and U15005 (N_15005,N_14612,N_14759);
xnor U15006 (N_15006,N_14375,N_14474);
and U15007 (N_15007,N_14624,N_14951);
and U15008 (N_15008,N_14463,N_14862);
and U15009 (N_15009,N_14614,N_14544);
nor U15010 (N_15010,N_14813,N_14393);
or U15011 (N_15011,N_14839,N_14826);
and U15012 (N_15012,N_14406,N_14424);
xor U15013 (N_15013,N_14833,N_14732);
xnor U15014 (N_15014,N_14617,N_14863);
nand U15015 (N_15015,N_14635,N_14967);
and U15016 (N_15016,N_14729,N_14886);
or U15017 (N_15017,N_14961,N_14670);
or U15018 (N_15018,N_14545,N_14709);
and U15019 (N_15019,N_14652,N_14927);
nand U15020 (N_15020,N_14739,N_14777);
nor U15021 (N_15021,N_14956,N_14508);
or U15022 (N_15022,N_14467,N_14609);
nand U15023 (N_15023,N_14390,N_14840);
or U15024 (N_15024,N_14660,N_14828);
nand U15025 (N_15025,N_14963,N_14619);
nand U15026 (N_15026,N_14388,N_14563);
xor U15027 (N_15027,N_14398,N_14613);
and U15028 (N_15028,N_14662,N_14626);
or U15029 (N_15029,N_14402,N_14628);
nor U15030 (N_15030,N_14451,N_14608);
or U15031 (N_15031,N_14941,N_14819);
and U15032 (N_15032,N_14940,N_14384);
xor U15033 (N_15033,N_14431,N_14722);
nor U15034 (N_15034,N_14610,N_14554);
nor U15035 (N_15035,N_14853,N_14841);
or U15036 (N_15036,N_14576,N_14925);
nand U15037 (N_15037,N_14380,N_14797);
xor U15038 (N_15038,N_14671,N_14493);
and U15039 (N_15039,N_14781,N_14439);
xor U15040 (N_15040,N_14791,N_14646);
nor U15041 (N_15041,N_14399,N_14557);
xnor U15042 (N_15042,N_14414,N_14538);
xor U15043 (N_15043,N_14426,N_14513);
nand U15044 (N_15044,N_14938,N_14550);
nand U15045 (N_15045,N_14654,N_14498);
nor U15046 (N_15046,N_14539,N_14857);
or U15047 (N_15047,N_14893,N_14549);
and U15048 (N_15048,N_14464,N_14778);
or U15049 (N_15049,N_14425,N_14438);
and U15050 (N_15050,N_14981,N_14490);
xnor U15051 (N_15051,N_14977,N_14383);
and U15052 (N_15052,N_14885,N_14703);
nand U15053 (N_15053,N_14410,N_14912);
and U15054 (N_15054,N_14803,N_14907);
nor U15055 (N_15055,N_14387,N_14872);
and U15056 (N_15056,N_14731,N_14452);
or U15057 (N_15057,N_14959,N_14392);
xor U15058 (N_15058,N_14611,N_14903);
or U15059 (N_15059,N_14753,N_14623);
and U15060 (N_15060,N_14672,N_14681);
xnor U15061 (N_15061,N_14700,N_14409);
nand U15062 (N_15062,N_14687,N_14586);
nand U15063 (N_15063,N_14567,N_14765);
nand U15064 (N_15064,N_14802,N_14405);
nor U15065 (N_15065,N_14458,N_14790);
nand U15066 (N_15066,N_14939,N_14536);
and U15067 (N_15067,N_14541,N_14752);
nor U15068 (N_15068,N_14879,N_14480);
nor U15069 (N_15069,N_14589,N_14994);
or U15070 (N_15070,N_14894,N_14779);
nor U15071 (N_15071,N_14835,N_14943);
or U15072 (N_15072,N_14898,N_14966);
or U15073 (N_15073,N_14740,N_14920);
xor U15074 (N_15074,N_14533,N_14641);
or U15075 (N_15075,N_14642,N_14553);
nor U15076 (N_15076,N_14761,N_14984);
xnor U15077 (N_15077,N_14607,N_14528);
and U15078 (N_15078,N_14572,N_14858);
xnor U15079 (N_15079,N_14808,N_14511);
nor U15080 (N_15080,N_14686,N_14957);
xor U15081 (N_15081,N_14798,N_14677);
nor U15082 (N_15082,N_14876,N_14823);
and U15083 (N_15083,N_14568,N_14408);
or U15084 (N_15084,N_14401,N_14807);
xor U15085 (N_15085,N_14794,N_14986);
xor U15086 (N_15086,N_14762,N_14389);
and U15087 (N_15087,N_14809,N_14908);
or U15088 (N_15088,N_14673,N_14806);
nand U15089 (N_15089,N_14397,N_14514);
or U15090 (N_15090,N_14877,N_14810);
nor U15091 (N_15091,N_14747,N_14697);
or U15092 (N_15092,N_14944,N_14844);
nand U15093 (N_15093,N_14995,N_14974);
nor U15094 (N_15094,N_14701,N_14475);
and U15095 (N_15095,N_14690,N_14379);
or U15096 (N_15096,N_14655,N_14648);
xor U15097 (N_15097,N_14429,N_14897);
nor U15098 (N_15098,N_14805,N_14849);
or U15099 (N_15099,N_14910,N_14597);
nor U15100 (N_15100,N_14588,N_14931);
nor U15101 (N_15101,N_14666,N_14960);
or U15102 (N_15102,N_14587,N_14584);
or U15103 (N_15103,N_14901,N_14712);
xnor U15104 (N_15104,N_14921,N_14481);
or U15105 (N_15105,N_14830,N_14933);
nand U15106 (N_15106,N_14815,N_14675);
or U15107 (N_15107,N_14705,N_14904);
nor U15108 (N_15108,N_14645,N_14721);
xnor U15109 (N_15109,N_14579,N_14510);
or U15110 (N_15110,N_14564,N_14825);
and U15111 (N_15111,N_14971,N_14770);
and U15112 (N_15112,N_14887,N_14743);
xor U15113 (N_15113,N_14469,N_14638);
nor U15114 (N_15114,N_14512,N_14559);
nor U15115 (N_15115,N_14945,N_14804);
and U15116 (N_15116,N_14500,N_14683);
nor U15117 (N_15117,N_14676,N_14569);
xor U15118 (N_15118,N_14627,N_14892);
and U15119 (N_15119,N_14750,N_14767);
xor U15120 (N_15120,N_14888,N_14834);
and U15121 (N_15121,N_14706,N_14485);
xnor U15122 (N_15122,N_14965,N_14860);
and U15123 (N_15123,N_14420,N_14922);
or U15124 (N_15124,N_14713,N_14923);
nor U15125 (N_15125,N_14914,N_14870);
nor U15126 (N_15126,N_14621,N_14932);
xor U15127 (N_15127,N_14783,N_14400);
nand U15128 (N_15128,N_14869,N_14952);
or U15129 (N_15129,N_14565,N_14726);
or U15130 (N_15130,N_14404,N_14385);
nand U15131 (N_15131,N_14518,N_14978);
nand U15132 (N_15132,N_14968,N_14822);
and U15133 (N_15133,N_14575,N_14606);
xnor U15134 (N_15134,N_14598,N_14501);
nor U15135 (N_15135,N_14854,N_14975);
xnor U15136 (N_15136,N_14454,N_14386);
and U15137 (N_15137,N_14622,N_14896);
and U15138 (N_15138,N_14407,N_14827);
nor U15139 (N_15139,N_14989,N_14976);
or U15140 (N_15140,N_14856,N_14911);
or U15141 (N_15141,N_14625,N_14682);
and U15142 (N_15142,N_14878,N_14678);
or U15143 (N_15143,N_14382,N_14616);
xor U15144 (N_15144,N_14580,N_14434);
nor U15145 (N_15145,N_14883,N_14499);
xnor U15146 (N_15146,N_14708,N_14766);
nand U15147 (N_15147,N_14774,N_14378);
nand U15148 (N_15148,N_14446,N_14585);
nand U15149 (N_15149,N_14688,N_14506);
and U15150 (N_15150,N_14685,N_14692);
xor U15151 (N_15151,N_14937,N_14942);
nand U15152 (N_15152,N_14442,N_14736);
or U15153 (N_15153,N_14799,N_14930);
xor U15154 (N_15154,N_14691,N_14737);
or U15155 (N_15155,N_14988,N_14573);
nor U15156 (N_15156,N_14814,N_14466);
or U15157 (N_15157,N_14430,N_14522);
or U15158 (N_15158,N_14704,N_14891);
nand U15159 (N_15159,N_14647,N_14482);
or U15160 (N_15160,N_14763,N_14667);
or U15161 (N_15161,N_14768,N_14643);
xnor U15162 (N_15162,N_14899,N_14832);
nor U15163 (N_15163,N_14459,N_14479);
nand U15164 (N_15164,N_14594,N_14601);
and U15165 (N_15165,N_14644,N_14950);
nor U15166 (N_15166,N_14465,N_14542);
nor U15167 (N_15167,N_14758,N_14754);
and U15168 (N_15168,N_14502,N_14818);
and U15169 (N_15169,N_14633,N_14448);
nor U15170 (N_15170,N_14720,N_14497);
xnor U15171 (N_15171,N_14560,N_14570);
xnor U15172 (N_15172,N_14926,N_14668);
or U15173 (N_15173,N_14900,N_14577);
nor U15174 (N_15174,N_14574,N_14450);
nor U15175 (N_15175,N_14377,N_14787);
or U15176 (N_15176,N_14916,N_14884);
xor U15177 (N_15177,N_14817,N_14483);
xor U15178 (N_15178,N_14918,N_14848);
or U15179 (N_15179,N_14786,N_14650);
or U15180 (N_15180,N_14821,N_14669);
nand U15181 (N_15181,N_14537,N_14503);
xor U15182 (N_15182,N_14531,N_14412);
nor U15183 (N_15183,N_14949,N_14868);
and U15184 (N_15184,N_14842,N_14615);
and U15185 (N_15185,N_14491,N_14435);
and U15186 (N_15186,N_14634,N_14394);
xor U15187 (N_15187,N_14551,N_14505);
xnor U15188 (N_15188,N_14707,N_14432);
and U15189 (N_15189,N_14526,N_14521);
nor U15190 (N_15190,N_14756,N_14422);
or U15191 (N_15191,N_14784,N_14954);
nand U15192 (N_15192,N_14717,N_14581);
or U15193 (N_15193,N_14970,N_14694);
nor U15194 (N_15194,N_14630,N_14590);
nand U15195 (N_15195,N_14780,N_14487);
xor U15196 (N_15196,N_14534,N_14795);
or U15197 (N_15197,N_14443,N_14693);
xor U15198 (N_15198,N_14947,N_14516);
and U15199 (N_15199,N_14846,N_14865);
and U15200 (N_15200,N_14769,N_14741);
and U15201 (N_15201,N_14733,N_14855);
nand U15202 (N_15202,N_14782,N_14785);
and U15203 (N_15203,N_14562,N_14788);
nor U15204 (N_15204,N_14411,N_14556);
and U15205 (N_15205,N_14462,N_14983);
or U15206 (N_15206,N_14689,N_14376);
nand U15207 (N_15207,N_14603,N_14757);
xor U15208 (N_15208,N_14702,N_14811);
or U15209 (N_15209,N_14934,N_14674);
and U15210 (N_15210,N_14760,N_14504);
nand U15211 (N_15211,N_14776,N_14596);
nand U15212 (N_15212,N_14591,N_14793);
or U15213 (N_15213,N_14851,N_14419);
and U15214 (N_15214,N_14812,N_14484);
nand U15215 (N_15215,N_14843,N_14629);
and U15216 (N_15216,N_14875,N_14695);
nand U15217 (N_15217,N_14656,N_14958);
xnor U15218 (N_15218,N_14418,N_14992);
or U15219 (N_15219,N_14964,N_14699);
nand U15220 (N_15220,N_14471,N_14486);
nand U15221 (N_15221,N_14456,N_14595);
nand U15222 (N_15222,N_14998,N_14973);
nand U15223 (N_15223,N_14987,N_14980);
or U15224 (N_15224,N_14792,N_14716);
nor U15225 (N_15225,N_14519,N_14663);
xor U15226 (N_15226,N_14664,N_14836);
and U15227 (N_15227,N_14800,N_14403);
and U15228 (N_15228,N_14838,N_14867);
nor U15229 (N_15229,N_14472,N_14924);
or U15230 (N_15230,N_14520,N_14651);
or U15231 (N_15231,N_14558,N_14935);
nand U15232 (N_15232,N_14755,N_14847);
nand U15233 (N_15233,N_14751,N_14515);
xnor U15234 (N_15234,N_14665,N_14509);
xnor U15235 (N_15235,N_14730,N_14715);
and U15236 (N_15236,N_14602,N_14972);
nand U15237 (N_15237,N_14566,N_14571);
nand U15238 (N_15238,N_14734,N_14928);
or U15239 (N_15239,N_14495,N_14746);
or U15240 (N_15240,N_14936,N_14946);
and U15241 (N_15241,N_14837,N_14582);
nand U15242 (N_15242,N_14468,N_14969);
nor U15243 (N_15243,N_14993,N_14748);
and U15244 (N_15244,N_14489,N_14861);
and U15245 (N_15245,N_14527,N_14631);
xor U15246 (N_15246,N_14962,N_14473);
and U15247 (N_15247,N_14447,N_14789);
xor U15248 (N_15248,N_14529,N_14824);
and U15249 (N_15249,N_14874,N_14455);
nand U15250 (N_15250,N_14738,N_14773);
or U15251 (N_15251,N_14649,N_14902);
nand U15252 (N_15252,N_14492,N_14801);
nand U15253 (N_15253,N_14684,N_14679);
nor U15254 (N_15254,N_14530,N_14535);
and U15255 (N_15255,N_14478,N_14919);
nand U15256 (N_15256,N_14997,N_14561);
xor U15257 (N_15257,N_14578,N_14996);
xnor U15258 (N_15258,N_14657,N_14552);
and U15259 (N_15259,N_14735,N_14831);
nand U15260 (N_15260,N_14600,N_14415);
and U15261 (N_15261,N_14453,N_14852);
and U15262 (N_15262,N_14727,N_14433);
xor U15263 (N_15263,N_14909,N_14953);
nor U15264 (N_15264,N_14895,N_14444);
and U15265 (N_15265,N_14391,N_14723);
xor U15266 (N_15266,N_14477,N_14890);
and U15267 (N_15267,N_14620,N_14659);
or U15268 (N_15268,N_14658,N_14437);
xnor U15269 (N_15269,N_14653,N_14999);
xnor U15270 (N_15270,N_14711,N_14985);
xor U15271 (N_15271,N_14881,N_14540);
xor U15272 (N_15272,N_14775,N_14982);
nor U15273 (N_15273,N_14604,N_14742);
nand U15274 (N_15274,N_14524,N_14772);
nand U15275 (N_15275,N_14460,N_14593);
nor U15276 (N_15276,N_14859,N_14661);
xor U15277 (N_15277,N_14905,N_14543);
nand U15278 (N_15278,N_14476,N_14488);
nor U15279 (N_15279,N_14850,N_14990);
nand U15280 (N_15280,N_14441,N_14866);
or U15281 (N_15281,N_14915,N_14436);
and U15282 (N_15282,N_14423,N_14421);
and U15283 (N_15283,N_14427,N_14745);
nand U15284 (N_15284,N_14882,N_14449);
and U15285 (N_15285,N_14955,N_14929);
nor U15286 (N_15286,N_14820,N_14771);
nand U15287 (N_15287,N_14880,N_14718);
nand U15288 (N_15288,N_14416,N_14637);
nor U15289 (N_15289,N_14461,N_14991);
and U15290 (N_15290,N_14719,N_14639);
nor U15291 (N_15291,N_14381,N_14698);
nand U15292 (N_15292,N_14710,N_14829);
or U15293 (N_15293,N_14889,N_14948);
xor U15294 (N_15294,N_14496,N_14523);
nand U15295 (N_15295,N_14395,N_14440);
nor U15296 (N_15296,N_14796,N_14696);
and U15297 (N_15297,N_14605,N_14494);
and U15298 (N_15298,N_14680,N_14871);
nand U15299 (N_15299,N_14816,N_14636);
and U15300 (N_15300,N_14979,N_14917);
nor U15301 (N_15301,N_14618,N_14470);
or U15302 (N_15302,N_14728,N_14913);
xnor U15303 (N_15303,N_14864,N_14413);
or U15304 (N_15304,N_14749,N_14632);
and U15305 (N_15305,N_14555,N_14417);
nor U15306 (N_15306,N_14532,N_14714);
and U15307 (N_15307,N_14592,N_14744);
nor U15308 (N_15308,N_14845,N_14640);
or U15309 (N_15309,N_14724,N_14507);
or U15310 (N_15310,N_14428,N_14548);
xnor U15311 (N_15311,N_14445,N_14599);
nor U15312 (N_15312,N_14517,N_14612);
and U15313 (N_15313,N_14504,N_14399);
xnor U15314 (N_15314,N_14846,N_14911);
nand U15315 (N_15315,N_14563,N_14967);
nand U15316 (N_15316,N_14949,N_14642);
and U15317 (N_15317,N_14579,N_14926);
or U15318 (N_15318,N_14956,N_14531);
and U15319 (N_15319,N_14640,N_14995);
nand U15320 (N_15320,N_14782,N_14863);
nand U15321 (N_15321,N_14698,N_14595);
nand U15322 (N_15322,N_14809,N_14522);
xnor U15323 (N_15323,N_14711,N_14950);
xnor U15324 (N_15324,N_14721,N_14608);
nand U15325 (N_15325,N_14582,N_14633);
and U15326 (N_15326,N_14669,N_14436);
nor U15327 (N_15327,N_14454,N_14467);
nand U15328 (N_15328,N_14428,N_14740);
and U15329 (N_15329,N_14587,N_14778);
xnor U15330 (N_15330,N_14971,N_14637);
nor U15331 (N_15331,N_14930,N_14596);
and U15332 (N_15332,N_14561,N_14764);
nor U15333 (N_15333,N_14738,N_14457);
or U15334 (N_15334,N_14865,N_14610);
or U15335 (N_15335,N_14864,N_14427);
xnor U15336 (N_15336,N_14689,N_14781);
nand U15337 (N_15337,N_14640,N_14769);
xnor U15338 (N_15338,N_14840,N_14538);
or U15339 (N_15339,N_14989,N_14851);
nor U15340 (N_15340,N_14944,N_14733);
and U15341 (N_15341,N_14615,N_14576);
or U15342 (N_15342,N_14685,N_14442);
nand U15343 (N_15343,N_14809,N_14467);
nor U15344 (N_15344,N_14496,N_14452);
nand U15345 (N_15345,N_14689,N_14582);
nand U15346 (N_15346,N_14524,N_14568);
xnor U15347 (N_15347,N_14685,N_14606);
nor U15348 (N_15348,N_14427,N_14858);
nor U15349 (N_15349,N_14468,N_14668);
or U15350 (N_15350,N_14499,N_14916);
or U15351 (N_15351,N_14411,N_14985);
xnor U15352 (N_15352,N_14735,N_14659);
nor U15353 (N_15353,N_14687,N_14670);
and U15354 (N_15354,N_14648,N_14669);
xnor U15355 (N_15355,N_14378,N_14992);
xor U15356 (N_15356,N_14972,N_14769);
nand U15357 (N_15357,N_14617,N_14382);
and U15358 (N_15358,N_14847,N_14454);
xnor U15359 (N_15359,N_14588,N_14799);
nor U15360 (N_15360,N_14762,N_14597);
or U15361 (N_15361,N_14912,N_14691);
nor U15362 (N_15362,N_14802,N_14822);
nand U15363 (N_15363,N_14400,N_14912);
xor U15364 (N_15364,N_14633,N_14966);
xor U15365 (N_15365,N_14465,N_14658);
nor U15366 (N_15366,N_14394,N_14392);
nor U15367 (N_15367,N_14566,N_14525);
nor U15368 (N_15368,N_14437,N_14420);
nor U15369 (N_15369,N_14759,N_14989);
xor U15370 (N_15370,N_14906,N_14392);
and U15371 (N_15371,N_14797,N_14648);
and U15372 (N_15372,N_14733,N_14909);
nand U15373 (N_15373,N_14855,N_14585);
nand U15374 (N_15374,N_14575,N_14905);
xnor U15375 (N_15375,N_14994,N_14859);
and U15376 (N_15376,N_14754,N_14395);
xor U15377 (N_15377,N_14731,N_14386);
or U15378 (N_15378,N_14633,N_14450);
and U15379 (N_15379,N_14881,N_14454);
nand U15380 (N_15380,N_14619,N_14669);
nor U15381 (N_15381,N_14508,N_14898);
xor U15382 (N_15382,N_14737,N_14950);
and U15383 (N_15383,N_14677,N_14581);
and U15384 (N_15384,N_14643,N_14787);
or U15385 (N_15385,N_14466,N_14756);
xor U15386 (N_15386,N_14523,N_14891);
nor U15387 (N_15387,N_14567,N_14595);
nor U15388 (N_15388,N_14746,N_14955);
nor U15389 (N_15389,N_14916,N_14812);
or U15390 (N_15390,N_14482,N_14499);
and U15391 (N_15391,N_14720,N_14877);
nor U15392 (N_15392,N_14834,N_14816);
or U15393 (N_15393,N_14703,N_14790);
nand U15394 (N_15394,N_14937,N_14705);
nor U15395 (N_15395,N_14784,N_14671);
or U15396 (N_15396,N_14517,N_14450);
and U15397 (N_15397,N_14590,N_14515);
or U15398 (N_15398,N_14628,N_14413);
xnor U15399 (N_15399,N_14916,N_14647);
nor U15400 (N_15400,N_14433,N_14934);
xor U15401 (N_15401,N_14431,N_14698);
or U15402 (N_15402,N_14838,N_14752);
and U15403 (N_15403,N_14755,N_14619);
xor U15404 (N_15404,N_14548,N_14583);
or U15405 (N_15405,N_14717,N_14723);
nor U15406 (N_15406,N_14589,N_14938);
and U15407 (N_15407,N_14527,N_14810);
nor U15408 (N_15408,N_14803,N_14825);
or U15409 (N_15409,N_14834,N_14956);
and U15410 (N_15410,N_14647,N_14673);
or U15411 (N_15411,N_14942,N_14667);
nor U15412 (N_15412,N_14912,N_14380);
and U15413 (N_15413,N_14669,N_14839);
nor U15414 (N_15414,N_14752,N_14420);
and U15415 (N_15415,N_14822,N_14832);
or U15416 (N_15416,N_14658,N_14972);
xor U15417 (N_15417,N_14827,N_14495);
xnor U15418 (N_15418,N_14389,N_14556);
and U15419 (N_15419,N_14764,N_14496);
or U15420 (N_15420,N_14646,N_14918);
nor U15421 (N_15421,N_14587,N_14745);
nor U15422 (N_15422,N_14651,N_14476);
nor U15423 (N_15423,N_14661,N_14887);
xnor U15424 (N_15424,N_14584,N_14888);
or U15425 (N_15425,N_14610,N_14416);
and U15426 (N_15426,N_14652,N_14498);
or U15427 (N_15427,N_14806,N_14432);
xnor U15428 (N_15428,N_14914,N_14436);
nor U15429 (N_15429,N_14619,N_14404);
nand U15430 (N_15430,N_14850,N_14584);
or U15431 (N_15431,N_14669,N_14970);
nand U15432 (N_15432,N_14769,N_14920);
xnor U15433 (N_15433,N_14814,N_14737);
or U15434 (N_15434,N_14503,N_14887);
and U15435 (N_15435,N_14933,N_14432);
and U15436 (N_15436,N_14845,N_14992);
nand U15437 (N_15437,N_14889,N_14579);
nor U15438 (N_15438,N_14642,N_14518);
and U15439 (N_15439,N_14877,N_14739);
nand U15440 (N_15440,N_14577,N_14601);
and U15441 (N_15441,N_14759,N_14413);
nand U15442 (N_15442,N_14723,N_14729);
nand U15443 (N_15443,N_14963,N_14876);
nand U15444 (N_15444,N_14893,N_14712);
nor U15445 (N_15445,N_14442,N_14892);
xnor U15446 (N_15446,N_14878,N_14384);
nor U15447 (N_15447,N_14915,N_14761);
nand U15448 (N_15448,N_14921,N_14552);
xor U15449 (N_15449,N_14941,N_14676);
nand U15450 (N_15450,N_14749,N_14742);
xor U15451 (N_15451,N_14684,N_14743);
and U15452 (N_15452,N_14921,N_14635);
or U15453 (N_15453,N_14380,N_14614);
nor U15454 (N_15454,N_14982,N_14585);
and U15455 (N_15455,N_14683,N_14384);
nor U15456 (N_15456,N_14965,N_14696);
and U15457 (N_15457,N_14728,N_14784);
nor U15458 (N_15458,N_14636,N_14896);
nor U15459 (N_15459,N_14566,N_14808);
nand U15460 (N_15460,N_14907,N_14743);
nand U15461 (N_15461,N_14651,N_14690);
nand U15462 (N_15462,N_14535,N_14767);
nor U15463 (N_15463,N_14836,N_14834);
nor U15464 (N_15464,N_14473,N_14664);
xor U15465 (N_15465,N_14735,N_14997);
nor U15466 (N_15466,N_14714,N_14906);
xnor U15467 (N_15467,N_14803,N_14719);
and U15468 (N_15468,N_14732,N_14971);
xnor U15469 (N_15469,N_14694,N_14721);
and U15470 (N_15470,N_14994,N_14601);
nand U15471 (N_15471,N_14525,N_14556);
xnor U15472 (N_15472,N_14912,N_14442);
nand U15473 (N_15473,N_14697,N_14760);
xnor U15474 (N_15474,N_14492,N_14529);
or U15475 (N_15475,N_14588,N_14972);
and U15476 (N_15476,N_14744,N_14726);
xnor U15477 (N_15477,N_14532,N_14508);
and U15478 (N_15478,N_14862,N_14731);
or U15479 (N_15479,N_14793,N_14986);
xnor U15480 (N_15480,N_14857,N_14898);
nand U15481 (N_15481,N_14602,N_14505);
nand U15482 (N_15482,N_14583,N_14409);
and U15483 (N_15483,N_14965,N_14381);
nor U15484 (N_15484,N_14829,N_14861);
and U15485 (N_15485,N_14776,N_14420);
nand U15486 (N_15486,N_14851,N_14832);
or U15487 (N_15487,N_14666,N_14651);
or U15488 (N_15488,N_14424,N_14774);
and U15489 (N_15489,N_14494,N_14527);
nand U15490 (N_15490,N_14387,N_14802);
nand U15491 (N_15491,N_14803,N_14380);
or U15492 (N_15492,N_14736,N_14403);
nand U15493 (N_15493,N_14975,N_14602);
nand U15494 (N_15494,N_14462,N_14832);
xnor U15495 (N_15495,N_14699,N_14954);
nor U15496 (N_15496,N_14515,N_14596);
or U15497 (N_15497,N_14695,N_14652);
nand U15498 (N_15498,N_14538,N_14406);
and U15499 (N_15499,N_14704,N_14476);
xor U15500 (N_15500,N_14449,N_14522);
xor U15501 (N_15501,N_14884,N_14430);
or U15502 (N_15502,N_14911,N_14725);
nor U15503 (N_15503,N_14587,N_14917);
xor U15504 (N_15504,N_14584,N_14615);
and U15505 (N_15505,N_14545,N_14963);
nand U15506 (N_15506,N_14833,N_14404);
nand U15507 (N_15507,N_14919,N_14847);
or U15508 (N_15508,N_14572,N_14710);
nand U15509 (N_15509,N_14678,N_14561);
xnor U15510 (N_15510,N_14517,N_14754);
xnor U15511 (N_15511,N_14598,N_14619);
or U15512 (N_15512,N_14510,N_14690);
or U15513 (N_15513,N_14676,N_14977);
xor U15514 (N_15514,N_14863,N_14940);
or U15515 (N_15515,N_14884,N_14676);
nor U15516 (N_15516,N_14636,N_14906);
or U15517 (N_15517,N_14797,N_14864);
nand U15518 (N_15518,N_14912,N_14430);
nand U15519 (N_15519,N_14545,N_14671);
xnor U15520 (N_15520,N_14376,N_14431);
nand U15521 (N_15521,N_14769,N_14735);
nand U15522 (N_15522,N_14551,N_14504);
nor U15523 (N_15523,N_14981,N_14425);
and U15524 (N_15524,N_14751,N_14631);
nor U15525 (N_15525,N_14535,N_14757);
or U15526 (N_15526,N_14675,N_14700);
xor U15527 (N_15527,N_14983,N_14870);
nor U15528 (N_15528,N_14603,N_14520);
nand U15529 (N_15529,N_14794,N_14719);
nand U15530 (N_15530,N_14386,N_14861);
nand U15531 (N_15531,N_14548,N_14837);
nor U15532 (N_15532,N_14438,N_14448);
or U15533 (N_15533,N_14605,N_14453);
xnor U15534 (N_15534,N_14518,N_14780);
nor U15535 (N_15535,N_14725,N_14625);
and U15536 (N_15536,N_14413,N_14515);
nor U15537 (N_15537,N_14929,N_14571);
xor U15538 (N_15538,N_14765,N_14785);
nor U15539 (N_15539,N_14516,N_14798);
and U15540 (N_15540,N_14439,N_14389);
nand U15541 (N_15541,N_14750,N_14789);
nor U15542 (N_15542,N_14830,N_14785);
nor U15543 (N_15543,N_14472,N_14804);
and U15544 (N_15544,N_14947,N_14424);
xnor U15545 (N_15545,N_14510,N_14875);
and U15546 (N_15546,N_14769,N_14895);
nand U15547 (N_15547,N_14990,N_14648);
or U15548 (N_15548,N_14711,N_14545);
xor U15549 (N_15549,N_14680,N_14497);
nor U15550 (N_15550,N_14846,N_14612);
nand U15551 (N_15551,N_14828,N_14832);
nor U15552 (N_15552,N_14981,N_14831);
nor U15553 (N_15553,N_14558,N_14978);
nor U15554 (N_15554,N_14390,N_14868);
xor U15555 (N_15555,N_14588,N_14600);
nor U15556 (N_15556,N_14766,N_14513);
or U15557 (N_15557,N_14934,N_14769);
or U15558 (N_15558,N_14945,N_14808);
or U15559 (N_15559,N_14398,N_14816);
or U15560 (N_15560,N_14437,N_14920);
nand U15561 (N_15561,N_14658,N_14747);
or U15562 (N_15562,N_14591,N_14828);
nand U15563 (N_15563,N_14485,N_14956);
nand U15564 (N_15564,N_14635,N_14800);
or U15565 (N_15565,N_14606,N_14637);
nor U15566 (N_15566,N_14919,N_14548);
and U15567 (N_15567,N_14424,N_14934);
or U15568 (N_15568,N_14487,N_14388);
xor U15569 (N_15569,N_14710,N_14904);
nand U15570 (N_15570,N_14959,N_14673);
nand U15571 (N_15571,N_14956,N_14991);
nand U15572 (N_15572,N_14380,N_14549);
or U15573 (N_15573,N_14785,N_14412);
or U15574 (N_15574,N_14582,N_14898);
nand U15575 (N_15575,N_14778,N_14996);
nor U15576 (N_15576,N_14430,N_14474);
xnor U15577 (N_15577,N_14445,N_14548);
xor U15578 (N_15578,N_14760,N_14935);
nand U15579 (N_15579,N_14901,N_14670);
nand U15580 (N_15580,N_14621,N_14716);
and U15581 (N_15581,N_14978,N_14748);
or U15582 (N_15582,N_14590,N_14979);
and U15583 (N_15583,N_14422,N_14955);
and U15584 (N_15584,N_14850,N_14601);
xor U15585 (N_15585,N_14534,N_14916);
or U15586 (N_15586,N_14735,N_14961);
nand U15587 (N_15587,N_14532,N_14967);
or U15588 (N_15588,N_14732,N_14825);
nor U15589 (N_15589,N_14507,N_14495);
and U15590 (N_15590,N_14413,N_14921);
and U15591 (N_15591,N_14451,N_14679);
or U15592 (N_15592,N_14820,N_14783);
nand U15593 (N_15593,N_14656,N_14463);
or U15594 (N_15594,N_14846,N_14994);
or U15595 (N_15595,N_14822,N_14787);
nand U15596 (N_15596,N_14958,N_14565);
or U15597 (N_15597,N_14782,N_14589);
nand U15598 (N_15598,N_14751,N_14665);
xnor U15599 (N_15599,N_14796,N_14701);
nand U15600 (N_15600,N_14383,N_14957);
xnor U15601 (N_15601,N_14387,N_14843);
xor U15602 (N_15602,N_14485,N_14620);
nand U15603 (N_15603,N_14431,N_14785);
nor U15604 (N_15604,N_14484,N_14730);
and U15605 (N_15605,N_14883,N_14994);
xnor U15606 (N_15606,N_14740,N_14742);
or U15607 (N_15607,N_14428,N_14451);
or U15608 (N_15608,N_14944,N_14429);
and U15609 (N_15609,N_14999,N_14694);
nand U15610 (N_15610,N_14481,N_14967);
nor U15611 (N_15611,N_14748,N_14399);
xor U15612 (N_15612,N_14734,N_14956);
nor U15613 (N_15613,N_14450,N_14683);
or U15614 (N_15614,N_14513,N_14800);
nand U15615 (N_15615,N_14752,N_14453);
and U15616 (N_15616,N_14979,N_14789);
nor U15617 (N_15617,N_14750,N_14738);
nand U15618 (N_15618,N_14543,N_14493);
or U15619 (N_15619,N_14429,N_14398);
xor U15620 (N_15620,N_14522,N_14406);
nand U15621 (N_15621,N_14477,N_14483);
xor U15622 (N_15622,N_14413,N_14896);
or U15623 (N_15623,N_14783,N_14447);
nor U15624 (N_15624,N_14694,N_14409);
nand U15625 (N_15625,N_15316,N_15073);
nand U15626 (N_15626,N_15515,N_15580);
xor U15627 (N_15627,N_15415,N_15134);
nand U15628 (N_15628,N_15300,N_15216);
or U15629 (N_15629,N_15416,N_15195);
nor U15630 (N_15630,N_15425,N_15505);
nand U15631 (N_15631,N_15143,N_15520);
nand U15632 (N_15632,N_15503,N_15160);
xor U15633 (N_15633,N_15056,N_15349);
nand U15634 (N_15634,N_15547,N_15156);
and U15635 (N_15635,N_15394,N_15271);
nand U15636 (N_15636,N_15240,N_15550);
or U15637 (N_15637,N_15612,N_15613);
nand U15638 (N_15638,N_15051,N_15152);
nand U15639 (N_15639,N_15578,N_15048);
nand U15640 (N_15640,N_15212,N_15010);
nand U15641 (N_15641,N_15042,N_15269);
or U15642 (N_15642,N_15275,N_15486);
or U15643 (N_15643,N_15317,N_15280);
or U15644 (N_15644,N_15003,N_15245);
xnor U15645 (N_15645,N_15226,N_15514);
and U15646 (N_15646,N_15436,N_15465);
nand U15647 (N_15647,N_15287,N_15090);
or U15648 (N_15648,N_15379,N_15462);
xnor U15649 (N_15649,N_15584,N_15421);
or U15650 (N_15650,N_15137,N_15603);
or U15651 (N_15651,N_15086,N_15323);
and U15652 (N_15652,N_15359,N_15201);
or U15653 (N_15653,N_15501,N_15313);
xor U15654 (N_15654,N_15293,N_15267);
or U15655 (N_15655,N_15609,N_15083);
xnor U15656 (N_15656,N_15062,N_15527);
and U15657 (N_15657,N_15571,N_15423);
nand U15658 (N_15658,N_15412,N_15213);
nand U15659 (N_15659,N_15124,N_15464);
or U15660 (N_15660,N_15344,N_15182);
or U15661 (N_15661,N_15385,N_15035);
or U15662 (N_15662,N_15327,N_15573);
nor U15663 (N_15663,N_15373,N_15176);
and U15664 (N_15664,N_15184,N_15457);
and U15665 (N_15665,N_15006,N_15542);
xnor U15666 (N_15666,N_15288,N_15526);
or U15667 (N_15667,N_15286,N_15130);
xnor U15668 (N_15668,N_15538,N_15189);
nor U15669 (N_15669,N_15570,N_15388);
nand U15670 (N_15670,N_15235,N_15561);
xnor U15671 (N_15671,N_15282,N_15377);
nand U15672 (N_15672,N_15046,N_15264);
nand U15673 (N_15673,N_15432,N_15548);
and U15674 (N_15674,N_15471,N_15504);
nor U15675 (N_15675,N_15311,N_15133);
xnor U15676 (N_15676,N_15304,N_15424);
and U15677 (N_15677,N_15025,N_15370);
xnor U15678 (N_15678,N_15446,N_15175);
or U15679 (N_15679,N_15163,N_15050);
or U15680 (N_15680,N_15326,N_15484);
nor U15681 (N_15681,N_15162,N_15539);
xor U15682 (N_15682,N_15509,N_15097);
nor U15683 (N_15683,N_15441,N_15599);
nor U15684 (N_15684,N_15249,N_15399);
nand U15685 (N_15685,N_15418,N_15618);
nor U15686 (N_15686,N_15071,N_15445);
nand U15687 (N_15687,N_15200,N_15408);
xnor U15688 (N_15688,N_15365,N_15467);
nand U15689 (N_15689,N_15207,N_15497);
and U15690 (N_15690,N_15104,N_15531);
nand U15691 (N_15691,N_15159,N_15543);
or U15692 (N_15692,N_15145,N_15289);
xor U15693 (N_15693,N_15219,N_15146);
xor U15694 (N_15694,N_15202,N_15103);
nand U15695 (N_15695,N_15227,N_15502);
xnor U15696 (N_15696,N_15248,N_15382);
nand U15697 (N_15697,N_15440,N_15234);
xor U15698 (N_15698,N_15591,N_15558);
and U15699 (N_15699,N_15252,N_15498);
or U15700 (N_15700,N_15028,N_15259);
and U15701 (N_15701,N_15582,N_15572);
nand U15702 (N_15702,N_15125,N_15278);
nand U15703 (N_15703,N_15400,N_15040);
xnor U15704 (N_15704,N_15358,N_15563);
and U15705 (N_15705,N_15560,N_15161);
xor U15706 (N_15706,N_15192,N_15238);
xnor U15707 (N_15707,N_15037,N_15528);
and U15708 (N_15708,N_15458,N_15617);
nand U15709 (N_15709,N_15138,N_15169);
or U15710 (N_15710,N_15517,N_15545);
and U15711 (N_15711,N_15622,N_15452);
nor U15712 (N_15712,N_15310,N_15453);
or U15713 (N_15713,N_15360,N_15448);
xor U15714 (N_15714,N_15144,N_15142);
or U15715 (N_15715,N_15002,N_15291);
nand U15716 (N_15716,N_15565,N_15211);
xor U15717 (N_15717,N_15055,N_15390);
and U15718 (N_15718,N_15020,N_15410);
nand U15719 (N_15719,N_15017,N_15540);
nand U15720 (N_15720,N_15567,N_15129);
or U15721 (N_15721,N_15038,N_15203);
and U15722 (N_15722,N_15149,N_15397);
xnor U15723 (N_15723,N_15244,N_15199);
or U15724 (N_15724,N_15292,N_15487);
xnor U15725 (N_15725,N_15091,N_15566);
and U15726 (N_15726,N_15583,N_15209);
nand U15727 (N_15727,N_15180,N_15556);
nand U15728 (N_15728,N_15336,N_15296);
and U15729 (N_15729,N_15481,N_15620);
or U15730 (N_15730,N_15237,N_15615);
and U15731 (N_15731,N_15574,N_15380);
nand U15732 (N_15732,N_15546,N_15529);
xor U15733 (N_15733,N_15034,N_15014);
nor U15734 (N_15734,N_15466,N_15215);
or U15735 (N_15735,N_15343,N_15404);
or U15736 (N_15736,N_15030,N_15590);
nor U15737 (N_15737,N_15396,N_15364);
nand U15738 (N_15738,N_15141,N_15032);
and U15739 (N_15739,N_15549,N_15621);
nand U15740 (N_15740,N_15513,N_15460);
nand U15741 (N_15741,N_15554,N_15284);
nand U15742 (N_15742,N_15575,N_15011);
xnor U15743 (N_15743,N_15229,N_15600);
nor U15744 (N_15744,N_15070,N_15270);
xnor U15745 (N_15745,N_15409,N_15601);
and U15746 (N_15746,N_15496,N_15510);
and U15747 (N_15747,N_15345,N_15322);
nand U15748 (N_15748,N_15290,N_15076);
and U15749 (N_15749,N_15263,N_15589);
nand U15750 (N_15750,N_15241,N_15395);
and U15751 (N_15751,N_15031,N_15350);
nor U15752 (N_15752,N_15158,N_15111);
xnor U15753 (N_15753,N_15593,N_15472);
nand U15754 (N_15754,N_15494,N_15431);
xor U15755 (N_15755,N_15063,N_15206);
or U15756 (N_15756,N_15614,N_15177);
nor U15757 (N_15757,N_15398,N_15616);
or U15758 (N_15758,N_15340,N_15255);
nand U15759 (N_15759,N_15151,N_15450);
nand U15760 (N_15760,N_15007,N_15272);
xor U15761 (N_15761,N_15131,N_15419);
and U15762 (N_15762,N_15171,N_15555);
or U15763 (N_15763,N_15164,N_15039);
and U15764 (N_15764,N_15389,N_15027);
xnor U15765 (N_15765,N_15420,N_15516);
and U15766 (N_15766,N_15059,N_15427);
and U15767 (N_15767,N_15198,N_15321);
or U15768 (N_15768,N_15606,N_15455);
or U15769 (N_15769,N_15181,N_15607);
xnor U15770 (N_15770,N_15536,N_15602);
and U15771 (N_15771,N_15208,N_15266);
xnor U15772 (N_15772,N_15491,N_15384);
xor U15773 (N_15773,N_15518,N_15507);
nand U15774 (N_15774,N_15081,N_15052);
and U15775 (N_15775,N_15231,N_15594);
nor U15776 (N_15776,N_15474,N_15387);
xnor U15777 (N_15777,N_15069,N_15298);
and U15778 (N_15778,N_15033,N_15595);
xor U15779 (N_15779,N_15470,N_15115);
nand U15780 (N_15780,N_15089,N_15147);
and U15781 (N_15781,N_15347,N_15619);
nor U15782 (N_15782,N_15224,N_15068);
nand U15783 (N_15783,N_15114,N_15085);
nand U15784 (N_15784,N_15155,N_15302);
xnor U15785 (N_15785,N_15375,N_15523);
and U15786 (N_15786,N_15093,N_15413);
or U15787 (N_15787,N_15443,N_15499);
or U15788 (N_15788,N_15016,N_15154);
and U15789 (N_15789,N_15108,N_15495);
or U15790 (N_15790,N_15333,N_15305);
and U15791 (N_15791,N_15009,N_15066);
xnor U15792 (N_15792,N_15294,N_15407);
nor U15793 (N_15793,N_15019,N_15352);
and U15794 (N_15794,N_15537,N_15274);
or U15795 (N_15795,N_15449,N_15511);
nand U15796 (N_15796,N_15329,N_15045);
nand U15797 (N_15797,N_15354,N_15193);
nand U15798 (N_15798,N_15429,N_15488);
and U15799 (N_15799,N_15053,N_15475);
nand U15800 (N_15800,N_15469,N_15544);
nor U15801 (N_15801,N_15074,N_15139);
nor U15802 (N_15802,N_15353,N_15306);
and U15803 (N_15803,N_15276,N_15119);
xnor U15804 (N_15804,N_15338,N_15218);
or U15805 (N_15805,N_15087,N_15341);
and U15806 (N_15806,N_15433,N_15004);
or U15807 (N_15807,N_15188,N_15592);
nor U15808 (N_15808,N_15109,N_15230);
and U15809 (N_15809,N_15301,N_15000);
or U15810 (N_15810,N_15233,N_15330);
and U15811 (N_15811,N_15172,N_15604);
xnor U15812 (N_15812,N_15092,N_15026);
and U15813 (N_15813,N_15493,N_15043);
nand U15814 (N_15814,N_15477,N_15369);
xnor U15815 (N_15815,N_15082,N_15307);
and U15816 (N_15816,N_15223,N_15439);
and U15817 (N_15817,N_15075,N_15150);
xor U15818 (N_15818,N_15437,N_15557);
nand U15819 (N_15819,N_15552,N_15283);
and U15820 (N_15820,N_15442,N_15403);
xnor U15821 (N_15821,N_15113,N_15140);
or U15822 (N_15822,N_15148,N_15568);
or U15823 (N_15823,N_15112,N_15444);
nand U15824 (N_15824,N_15366,N_15088);
nand U15825 (N_15825,N_15170,N_15118);
xor U15826 (N_15826,N_15553,N_15247);
xor U15827 (N_15827,N_15179,N_15157);
nor U15828 (N_15828,N_15361,N_15058);
and U15829 (N_15829,N_15374,N_15610);
and U15830 (N_15830,N_15253,N_15183);
and U15831 (N_15831,N_15588,N_15220);
and U15832 (N_15832,N_15428,N_15079);
nor U15833 (N_15833,N_15232,N_15015);
or U15834 (N_15834,N_15239,N_15204);
xnor U15835 (N_15835,N_15562,N_15222);
nor U15836 (N_15836,N_15049,N_15101);
nand U15837 (N_15837,N_15054,N_15100);
nand U15838 (N_15838,N_15228,N_15411);
nand U15839 (N_15839,N_15587,N_15367);
xor U15840 (N_15840,N_15022,N_15559);
nor U15841 (N_15841,N_15351,N_15297);
xor U15842 (N_15842,N_15386,N_15196);
nand U15843 (N_15843,N_15459,N_15107);
nor U15844 (N_15844,N_15479,N_15257);
or U15845 (N_15845,N_15047,N_15067);
xor U15846 (N_15846,N_15197,N_15094);
or U15847 (N_15847,N_15483,N_15564);
and U15848 (N_15848,N_15106,N_15057);
xor U15849 (N_15849,N_15476,N_15569);
nor U15850 (N_15850,N_15210,N_15318);
xor U15851 (N_15851,N_15256,N_15029);
nor U15852 (N_15852,N_15173,N_15324);
nor U15853 (N_15853,N_15013,N_15008);
nand U15854 (N_15854,N_15530,N_15331);
or U15855 (N_15855,N_15246,N_15187);
xor U15856 (N_15856,N_15191,N_15576);
nor U15857 (N_15857,N_15402,N_15277);
nand U15858 (N_15858,N_15102,N_15328);
nor U15859 (N_15859,N_15339,N_15356);
xnor U15860 (N_15860,N_15371,N_15186);
nand U15861 (N_15861,N_15036,N_15185);
nor U15862 (N_15862,N_15392,N_15041);
or U15863 (N_15863,N_15126,N_15312);
and U15864 (N_15864,N_15174,N_15096);
nand U15865 (N_15865,N_15468,N_15018);
or U15866 (N_15866,N_15205,N_15167);
or U15867 (N_15867,N_15372,N_15078);
or U15868 (N_15868,N_15451,N_15190);
and U15869 (N_15869,N_15273,N_15251);
xor U15870 (N_15870,N_15586,N_15116);
nor U15871 (N_15871,N_15363,N_15378);
nand U15872 (N_15872,N_15262,N_15426);
nor U15873 (N_15873,N_15524,N_15492);
xnor U15874 (N_15874,N_15065,N_15585);
or U15875 (N_15875,N_15095,N_15105);
nand U15876 (N_15876,N_15295,N_15362);
and U15877 (N_15877,N_15532,N_15221);
nor U15878 (N_15878,N_15012,N_15368);
and U15879 (N_15879,N_15447,N_15414);
nor U15880 (N_15880,N_15577,N_15463);
or U15881 (N_15881,N_15454,N_15393);
nor U15882 (N_15882,N_15506,N_15005);
and U15883 (N_15883,N_15456,N_15519);
nor U15884 (N_15884,N_15348,N_15383);
nor U15885 (N_15885,N_15250,N_15332);
nor U15886 (N_15886,N_15072,N_15422);
or U15887 (N_15887,N_15099,N_15334);
or U15888 (N_15888,N_15279,N_15521);
nand U15889 (N_15889,N_15533,N_15024);
and U15890 (N_15890,N_15417,N_15254);
and U15891 (N_15891,N_15060,N_15551);
and U15892 (N_15892,N_15315,N_15461);
or U15893 (N_15893,N_15534,N_15123);
xnor U15894 (N_15894,N_15136,N_15243);
and U15895 (N_15895,N_15061,N_15605);
xnor U15896 (N_15896,N_15473,N_15608);
and U15897 (N_15897,N_15303,N_15522);
and U15898 (N_15898,N_15512,N_15117);
nor U15899 (N_15899,N_15597,N_15342);
or U15900 (N_15900,N_15611,N_15077);
or U15901 (N_15901,N_15541,N_15281);
nand U15902 (N_15902,N_15581,N_15023);
or U15903 (N_15903,N_15261,N_15128);
nand U15904 (N_15904,N_15355,N_15135);
and U15905 (N_15905,N_15535,N_15225);
or U15906 (N_15906,N_15381,N_15320);
nor U15907 (N_15907,N_15120,N_15098);
nor U15908 (N_15908,N_15508,N_15110);
and U15909 (N_15909,N_15265,N_15480);
xnor U15910 (N_15910,N_15064,N_15335);
nor U15911 (N_15911,N_15319,N_15485);
or U15912 (N_15912,N_15435,N_15122);
and U15913 (N_15913,N_15478,N_15127);
and U15914 (N_15914,N_15214,N_15121);
xnor U15915 (N_15915,N_15268,N_15482);
or U15916 (N_15916,N_15260,N_15242);
xor U15917 (N_15917,N_15500,N_15525);
and U15918 (N_15918,N_15217,N_15337);
nor U15919 (N_15919,N_15598,N_15044);
and U15920 (N_15920,N_15596,N_15258);
nor U15921 (N_15921,N_15401,N_15236);
or U15922 (N_15922,N_15376,N_15132);
nor U15923 (N_15923,N_15406,N_15490);
or U15924 (N_15924,N_15391,N_15579);
nand U15925 (N_15925,N_15084,N_15325);
nand U15926 (N_15926,N_15489,N_15194);
nand U15927 (N_15927,N_15623,N_15405);
or U15928 (N_15928,N_15178,N_15001);
and U15929 (N_15929,N_15314,N_15309);
nor U15930 (N_15930,N_15080,N_15168);
nand U15931 (N_15931,N_15285,N_15430);
and U15932 (N_15932,N_15308,N_15021);
xor U15933 (N_15933,N_15346,N_15166);
xor U15934 (N_15934,N_15153,N_15357);
nand U15935 (N_15935,N_15299,N_15165);
nand U15936 (N_15936,N_15434,N_15624);
and U15937 (N_15937,N_15438,N_15223);
or U15938 (N_15938,N_15075,N_15194);
xor U15939 (N_15939,N_15323,N_15595);
or U15940 (N_15940,N_15612,N_15221);
and U15941 (N_15941,N_15563,N_15309);
xnor U15942 (N_15942,N_15026,N_15397);
nand U15943 (N_15943,N_15301,N_15478);
and U15944 (N_15944,N_15549,N_15019);
nand U15945 (N_15945,N_15269,N_15544);
nor U15946 (N_15946,N_15029,N_15284);
xnor U15947 (N_15947,N_15565,N_15532);
and U15948 (N_15948,N_15030,N_15293);
or U15949 (N_15949,N_15338,N_15256);
or U15950 (N_15950,N_15486,N_15212);
or U15951 (N_15951,N_15355,N_15040);
and U15952 (N_15952,N_15514,N_15517);
or U15953 (N_15953,N_15216,N_15232);
nor U15954 (N_15954,N_15098,N_15252);
xnor U15955 (N_15955,N_15584,N_15099);
xnor U15956 (N_15956,N_15099,N_15484);
xor U15957 (N_15957,N_15080,N_15216);
nor U15958 (N_15958,N_15085,N_15176);
and U15959 (N_15959,N_15427,N_15565);
nor U15960 (N_15960,N_15257,N_15169);
nand U15961 (N_15961,N_15564,N_15470);
and U15962 (N_15962,N_15329,N_15175);
nand U15963 (N_15963,N_15279,N_15592);
xor U15964 (N_15964,N_15441,N_15197);
or U15965 (N_15965,N_15129,N_15078);
nand U15966 (N_15966,N_15536,N_15106);
and U15967 (N_15967,N_15121,N_15522);
nor U15968 (N_15968,N_15021,N_15384);
nor U15969 (N_15969,N_15212,N_15232);
nor U15970 (N_15970,N_15478,N_15416);
and U15971 (N_15971,N_15303,N_15558);
xor U15972 (N_15972,N_15477,N_15065);
nand U15973 (N_15973,N_15230,N_15573);
and U15974 (N_15974,N_15332,N_15026);
or U15975 (N_15975,N_15515,N_15218);
and U15976 (N_15976,N_15470,N_15212);
xor U15977 (N_15977,N_15234,N_15532);
xor U15978 (N_15978,N_15093,N_15362);
or U15979 (N_15979,N_15482,N_15109);
nor U15980 (N_15980,N_15410,N_15268);
nand U15981 (N_15981,N_15550,N_15527);
nand U15982 (N_15982,N_15039,N_15001);
nor U15983 (N_15983,N_15513,N_15541);
nand U15984 (N_15984,N_15045,N_15130);
xor U15985 (N_15985,N_15418,N_15044);
or U15986 (N_15986,N_15047,N_15307);
xor U15987 (N_15987,N_15396,N_15146);
nor U15988 (N_15988,N_15539,N_15554);
and U15989 (N_15989,N_15268,N_15557);
or U15990 (N_15990,N_15087,N_15296);
and U15991 (N_15991,N_15516,N_15621);
and U15992 (N_15992,N_15562,N_15124);
nor U15993 (N_15993,N_15550,N_15579);
nand U15994 (N_15994,N_15399,N_15041);
and U15995 (N_15995,N_15568,N_15278);
nor U15996 (N_15996,N_15569,N_15275);
xnor U15997 (N_15997,N_15350,N_15063);
xnor U15998 (N_15998,N_15129,N_15450);
xor U15999 (N_15999,N_15097,N_15281);
nand U16000 (N_16000,N_15346,N_15111);
or U16001 (N_16001,N_15035,N_15614);
and U16002 (N_16002,N_15560,N_15573);
or U16003 (N_16003,N_15544,N_15120);
nor U16004 (N_16004,N_15074,N_15070);
nand U16005 (N_16005,N_15585,N_15214);
and U16006 (N_16006,N_15085,N_15116);
or U16007 (N_16007,N_15085,N_15243);
nor U16008 (N_16008,N_15563,N_15295);
nor U16009 (N_16009,N_15146,N_15267);
nor U16010 (N_16010,N_15136,N_15011);
or U16011 (N_16011,N_15384,N_15420);
nor U16012 (N_16012,N_15615,N_15441);
nor U16013 (N_16013,N_15440,N_15443);
nor U16014 (N_16014,N_15329,N_15272);
or U16015 (N_16015,N_15410,N_15480);
or U16016 (N_16016,N_15009,N_15535);
nor U16017 (N_16017,N_15482,N_15210);
nor U16018 (N_16018,N_15096,N_15245);
nand U16019 (N_16019,N_15204,N_15099);
nor U16020 (N_16020,N_15399,N_15272);
nor U16021 (N_16021,N_15119,N_15107);
nand U16022 (N_16022,N_15300,N_15353);
and U16023 (N_16023,N_15183,N_15048);
xnor U16024 (N_16024,N_15401,N_15050);
nor U16025 (N_16025,N_15375,N_15252);
nand U16026 (N_16026,N_15217,N_15293);
and U16027 (N_16027,N_15322,N_15021);
nand U16028 (N_16028,N_15528,N_15597);
or U16029 (N_16029,N_15003,N_15347);
and U16030 (N_16030,N_15571,N_15371);
xor U16031 (N_16031,N_15096,N_15081);
nor U16032 (N_16032,N_15132,N_15048);
xnor U16033 (N_16033,N_15538,N_15373);
nor U16034 (N_16034,N_15280,N_15113);
xor U16035 (N_16035,N_15343,N_15069);
or U16036 (N_16036,N_15162,N_15038);
and U16037 (N_16037,N_15122,N_15093);
nand U16038 (N_16038,N_15406,N_15561);
and U16039 (N_16039,N_15059,N_15206);
xnor U16040 (N_16040,N_15459,N_15043);
nand U16041 (N_16041,N_15510,N_15146);
nand U16042 (N_16042,N_15379,N_15593);
xor U16043 (N_16043,N_15276,N_15287);
xnor U16044 (N_16044,N_15196,N_15395);
or U16045 (N_16045,N_15356,N_15374);
xnor U16046 (N_16046,N_15128,N_15072);
and U16047 (N_16047,N_15345,N_15030);
xor U16048 (N_16048,N_15151,N_15389);
nand U16049 (N_16049,N_15614,N_15365);
xnor U16050 (N_16050,N_15585,N_15030);
xnor U16051 (N_16051,N_15528,N_15277);
xnor U16052 (N_16052,N_15030,N_15358);
nand U16053 (N_16053,N_15098,N_15609);
nor U16054 (N_16054,N_15603,N_15294);
nor U16055 (N_16055,N_15074,N_15078);
xor U16056 (N_16056,N_15134,N_15126);
xnor U16057 (N_16057,N_15231,N_15511);
and U16058 (N_16058,N_15065,N_15511);
nand U16059 (N_16059,N_15614,N_15245);
nor U16060 (N_16060,N_15590,N_15519);
nor U16061 (N_16061,N_15312,N_15584);
and U16062 (N_16062,N_15059,N_15218);
and U16063 (N_16063,N_15165,N_15002);
or U16064 (N_16064,N_15622,N_15521);
and U16065 (N_16065,N_15005,N_15401);
nand U16066 (N_16066,N_15507,N_15145);
nor U16067 (N_16067,N_15323,N_15503);
nor U16068 (N_16068,N_15401,N_15519);
nand U16069 (N_16069,N_15480,N_15315);
xor U16070 (N_16070,N_15033,N_15241);
nor U16071 (N_16071,N_15114,N_15279);
nand U16072 (N_16072,N_15084,N_15441);
and U16073 (N_16073,N_15022,N_15210);
xor U16074 (N_16074,N_15268,N_15020);
nor U16075 (N_16075,N_15280,N_15619);
nor U16076 (N_16076,N_15183,N_15197);
nor U16077 (N_16077,N_15198,N_15318);
or U16078 (N_16078,N_15084,N_15013);
nand U16079 (N_16079,N_15354,N_15559);
or U16080 (N_16080,N_15503,N_15174);
and U16081 (N_16081,N_15382,N_15247);
or U16082 (N_16082,N_15335,N_15137);
nand U16083 (N_16083,N_15252,N_15289);
and U16084 (N_16084,N_15496,N_15564);
xnor U16085 (N_16085,N_15102,N_15341);
xor U16086 (N_16086,N_15476,N_15103);
nor U16087 (N_16087,N_15439,N_15157);
xor U16088 (N_16088,N_15620,N_15245);
and U16089 (N_16089,N_15404,N_15318);
and U16090 (N_16090,N_15355,N_15127);
xnor U16091 (N_16091,N_15328,N_15375);
or U16092 (N_16092,N_15375,N_15096);
or U16093 (N_16093,N_15583,N_15140);
and U16094 (N_16094,N_15123,N_15154);
and U16095 (N_16095,N_15448,N_15610);
and U16096 (N_16096,N_15514,N_15606);
or U16097 (N_16097,N_15200,N_15208);
or U16098 (N_16098,N_15392,N_15528);
and U16099 (N_16099,N_15269,N_15343);
nand U16100 (N_16100,N_15439,N_15516);
or U16101 (N_16101,N_15474,N_15226);
nor U16102 (N_16102,N_15151,N_15583);
nor U16103 (N_16103,N_15520,N_15150);
nand U16104 (N_16104,N_15616,N_15109);
or U16105 (N_16105,N_15442,N_15581);
and U16106 (N_16106,N_15344,N_15170);
and U16107 (N_16107,N_15281,N_15577);
and U16108 (N_16108,N_15295,N_15364);
nand U16109 (N_16109,N_15496,N_15331);
and U16110 (N_16110,N_15360,N_15598);
xor U16111 (N_16111,N_15257,N_15533);
or U16112 (N_16112,N_15553,N_15338);
nand U16113 (N_16113,N_15216,N_15118);
or U16114 (N_16114,N_15434,N_15047);
or U16115 (N_16115,N_15422,N_15164);
nor U16116 (N_16116,N_15489,N_15315);
nor U16117 (N_16117,N_15235,N_15166);
or U16118 (N_16118,N_15043,N_15172);
nand U16119 (N_16119,N_15431,N_15112);
or U16120 (N_16120,N_15473,N_15567);
and U16121 (N_16121,N_15620,N_15314);
or U16122 (N_16122,N_15301,N_15615);
nand U16123 (N_16123,N_15164,N_15043);
nor U16124 (N_16124,N_15004,N_15607);
nor U16125 (N_16125,N_15451,N_15410);
xnor U16126 (N_16126,N_15260,N_15482);
and U16127 (N_16127,N_15155,N_15576);
nor U16128 (N_16128,N_15157,N_15543);
xor U16129 (N_16129,N_15329,N_15243);
and U16130 (N_16130,N_15051,N_15484);
nand U16131 (N_16131,N_15189,N_15168);
nor U16132 (N_16132,N_15129,N_15063);
nand U16133 (N_16133,N_15423,N_15446);
or U16134 (N_16134,N_15119,N_15290);
xor U16135 (N_16135,N_15215,N_15136);
or U16136 (N_16136,N_15286,N_15214);
xor U16137 (N_16137,N_15134,N_15214);
and U16138 (N_16138,N_15521,N_15266);
nor U16139 (N_16139,N_15586,N_15045);
or U16140 (N_16140,N_15109,N_15457);
nand U16141 (N_16141,N_15517,N_15533);
or U16142 (N_16142,N_15064,N_15084);
nor U16143 (N_16143,N_15494,N_15425);
or U16144 (N_16144,N_15584,N_15131);
or U16145 (N_16145,N_15478,N_15586);
xor U16146 (N_16146,N_15459,N_15083);
nor U16147 (N_16147,N_15465,N_15332);
or U16148 (N_16148,N_15192,N_15353);
xor U16149 (N_16149,N_15167,N_15411);
nor U16150 (N_16150,N_15375,N_15168);
nor U16151 (N_16151,N_15332,N_15329);
or U16152 (N_16152,N_15303,N_15370);
nor U16153 (N_16153,N_15339,N_15017);
nor U16154 (N_16154,N_15028,N_15218);
xor U16155 (N_16155,N_15129,N_15552);
nand U16156 (N_16156,N_15256,N_15604);
xnor U16157 (N_16157,N_15263,N_15573);
or U16158 (N_16158,N_15522,N_15375);
nor U16159 (N_16159,N_15611,N_15064);
or U16160 (N_16160,N_15186,N_15278);
and U16161 (N_16161,N_15219,N_15366);
nand U16162 (N_16162,N_15110,N_15396);
nor U16163 (N_16163,N_15159,N_15173);
nor U16164 (N_16164,N_15339,N_15066);
nor U16165 (N_16165,N_15402,N_15131);
and U16166 (N_16166,N_15328,N_15516);
nor U16167 (N_16167,N_15597,N_15411);
or U16168 (N_16168,N_15215,N_15256);
nand U16169 (N_16169,N_15415,N_15025);
nand U16170 (N_16170,N_15173,N_15571);
xor U16171 (N_16171,N_15466,N_15147);
nor U16172 (N_16172,N_15365,N_15606);
nor U16173 (N_16173,N_15252,N_15204);
nor U16174 (N_16174,N_15300,N_15596);
or U16175 (N_16175,N_15581,N_15584);
and U16176 (N_16176,N_15390,N_15313);
nor U16177 (N_16177,N_15060,N_15321);
nand U16178 (N_16178,N_15468,N_15033);
nand U16179 (N_16179,N_15532,N_15217);
or U16180 (N_16180,N_15359,N_15145);
nor U16181 (N_16181,N_15411,N_15059);
nor U16182 (N_16182,N_15213,N_15441);
and U16183 (N_16183,N_15285,N_15515);
xor U16184 (N_16184,N_15016,N_15082);
or U16185 (N_16185,N_15451,N_15179);
nand U16186 (N_16186,N_15457,N_15426);
nand U16187 (N_16187,N_15602,N_15026);
xor U16188 (N_16188,N_15315,N_15211);
nor U16189 (N_16189,N_15495,N_15270);
and U16190 (N_16190,N_15211,N_15531);
or U16191 (N_16191,N_15620,N_15156);
xnor U16192 (N_16192,N_15072,N_15020);
or U16193 (N_16193,N_15071,N_15443);
nand U16194 (N_16194,N_15270,N_15408);
or U16195 (N_16195,N_15202,N_15573);
nor U16196 (N_16196,N_15090,N_15283);
nor U16197 (N_16197,N_15052,N_15162);
nor U16198 (N_16198,N_15371,N_15450);
nand U16199 (N_16199,N_15564,N_15527);
and U16200 (N_16200,N_15071,N_15592);
xor U16201 (N_16201,N_15136,N_15439);
or U16202 (N_16202,N_15495,N_15461);
nor U16203 (N_16203,N_15016,N_15227);
xor U16204 (N_16204,N_15281,N_15422);
xor U16205 (N_16205,N_15039,N_15050);
nor U16206 (N_16206,N_15144,N_15038);
or U16207 (N_16207,N_15439,N_15597);
or U16208 (N_16208,N_15274,N_15221);
or U16209 (N_16209,N_15026,N_15550);
nor U16210 (N_16210,N_15436,N_15532);
and U16211 (N_16211,N_15265,N_15162);
and U16212 (N_16212,N_15092,N_15170);
and U16213 (N_16213,N_15298,N_15074);
and U16214 (N_16214,N_15014,N_15096);
nor U16215 (N_16215,N_15004,N_15448);
nand U16216 (N_16216,N_15249,N_15186);
or U16217 (N_16217,N_15341,N_15582);
and U16218 (N_16218,N_15463,N_15039);
and U16219 (N_16219,N_15350,N_15065);
or U16220 (N_16220,N_15317,N_15234);
nor U16221 (N_16221,N_15013,N_15003);
xor U16222 (N_16222,N_15208,N_15141);
nor U16223 (N_16223,N_15492,N_15410);
nor U16224 (N_16224,N_15064,N_15429);
nand U16225 (N_16225,N_15254,N_15439);
or U16226 (N_16226,N_15560,N_15185);
or U16227 (N_16227,N_15622,N_15548);
and U16228 (N_16228,N_15434,N_15238);
and U16229 (N_16229,N_15305,N_15113);
nand U16230 (N_16230,N_15189,N_15503);
nor U16231 (N_16231,N_15338,N_15491);
nor U16232 (N_16232,N_15138,N_15413);
or U16233 (N_16233,N_15225,N_15464);
or U16234 (N_16234,N_15154,N_15614);
or U16235 (N_16235,N_15231,N_15347);
nor U16236 (N_16236,N_15497,N_15581);
nor U16237 (N_16237,N_15250,N_15148);
or U16238 (N_16238,N_15548,N_15583);
nor U16239 (N_16239,N_15362,N_15228);
nor U16240 (N_16240,N_15227,N_15545);
or U16241 (N_16241,N_15394,N_15007);
or U16242 (N_16242,N_15158,N_15268);
nand U16243 (N_16243,N_15561,N_15216);
and U16244 (N_16244,N_15108,N_15178);
nand U16245 (N_16245,N_15539,N_15575);
xnor U16246 (N_16246,N_15169,N_15436);
xnor U16247 (N_16247,N_15097,N_15334);
and U16248 (N_16248,N_15116,N_15172);
or U16249 (N_16249,N_15126,N_15552);
nand U16250 (N_16250,N_15914,N_15672);
xnor U16251 (N_16251,N_15905,N_16101);
xnor U16252 (N_16252,N_16200,N_15920);
nand U16253 (N_16253,N_16193,N_15719);
xor U16254 (N_16254,N_15828,N_16174);
nand U16255 (N_16255,N_15701,N_16197);
nand U16256 (N_16256,N_16219,N_15922);
and U16257 (N_16257,N_16068,N_16236);
and U16258 (N_16258,N_16071,N_16194);
and U16259 (N_16259,N_16038,N_16110);
xnor U16260 (N_16260,N_15885,N_15637);
xnor U16261 (N_16261,N_15663,N_15945);
or U16262 (N_16262,N_16098,N_16074);
and U16263 (N_16263,N_15711,N_15951);
nand U16264 (N_16264,N_15941,N_15875);
nand U16265 (N_16265,N_15819,N_16225);
xor U16266 (N_16266,N_16120,N_15915);
nor U16267 (N_16267,N_15666,N_15759);
nor U16268 (N_16268,N_15659,N_15751);
nand U16269 (N_16269,N_15859,N_16094);
nor U16270 (N_16270,N_15849,N_15928);
xnor U16271 (N_16271,N_15833,N_16083);
nor U16272 (N_16272,N_15767,N_15886);
nand U16273 (N_16273,N_16076,N_15668);
and U16274 (N_16274,N_15664,N_15726);
nor U16275 (N_16275,N_15873,N_15808);
or U16276 (N_16276,N_15946,N_15647);
nand U16277 (N_16277,N_15916,N_15682);
and U16278 (N_16278,N_15702,N_15684);
or U16279 (N_16279,N_15827,N_15938);
xor U16280 (N_16280,N_16012,N_16000);
nor U16281 (N_16281,N_15626,N_15636);
nand U16282 (N_16282,N_15776,N_16018);
xnor U16283 (N_16283,N_16141,N_15689);
xor U16284 (N_16284,N_15734,N_15692);
nor U16285 (N_16285,N_15925,N_15822);
and U16286 (N_16286,N_16165,N_15867);
nand U16287 (N_16287,N_15694,N_15820);
and U16288 (N_16288,N_16234,N_16053);
xor U16289 (N_16289,N_16213,N_16228);
nand U16290 (N_16290,N_15932,N_15796);
xnor U16291 (N_16291,N_15688,N_16080);
or U16292 (N_16292,N_15840,N_16001);
nand U16293 (N_16293,N_15816,N_16026);
nand U16294 (N_16294,N_15812,N_16181);
xor U16295 (N_16295,N_15721,N_16161);
or U16296 (N_16296,N_15780,N_16077);
and U16297 (N_16297,N_15940,N_16099);
or U16298 (N_16298,N_15802,N_15844);
or U16299 (N_16299,N_15720,N_15893);
and U16300 (N_16300,N_16243,N_15884);
nand U16301 (N_16301,N_15912,N_15927);
xnor U16302 (N_16302,N_16007,N_15674);
xnor U16303 (N_16303,N_15696,N_16072);
and U16304 (N_16304,N_15864,N_15671);
nand U16305 (N_16305,N_15649,N_15628);
nor U16306 (N_16306,N_15980,N_16056);
or U16307 (N_16307,N_16132,N_15657);
or U16308 (N_16308,N_15866,N_16180);
and U16309 (N_16309,N_15846,N_15960);
nand U16310 (N_16310,N_15662,N_15740);
and U16311 (N_16311,N_16017,N_16048);
or U16312 (N_16312,N_15797,N_15937);
or U16313 (N_16313,N_15970,N_16221);
and U16314 (N_16314,N_15803,N_16081);
nor U16315 (N_16315,N_15641,N_15775);
xor U16316 (N_16316,N_16037,N_15973);
xnor U16317 (N_16317,N_16058,N_15708);
and U16318 (N_16318,N_16168,N_15838);
nand U16319 (N_16319,N_15790,N_15826);
xor U16320 (N_16320,N_15817,N_15997);
xnor U16321 (N_16321,N_16237,N_15986);
and U16322 (N_16322,N_16104,N_15648);
or U16323 (N_16323,N_15761,N_16060);
nand U16324 (N_16324,N_16059,N_16023);
nand U16325 (N_16325,N_15800,N_16019);
nor U16326 (N_16326,N_16136,N_16046);
nand U16327 (N_16327,N_15995,N_16041);
xnor U16328 (N_16328,N_16008,N_16126);
nor U16329 (N_16329,N_16129,N_15839);
and U16330 (N_16330,N_15673,N_16108);
or U16331 (N_16331,N_16172,N_15752);
and U16332 (N_16332,N_15789,N_15918);
nand U16333 (N_16333,N_16179,N_16182);
nor U16334 (N_16334,N_15877,N_16201);
and U16335 (N_16335,N_15677,N_16118);
nor U16336 (N_16336,N_15934,N_16152);
and U16337 (N_16337,N_15627,N_16128);
xnor U16338 (N_16338,N_15923,N_16249);
nor U16339 (N_16339,N_16208,N_16044);
xnor U16340 (N_16340,N_15658,N_15656);
and U16341 (N_16341,N_15795,N_15785);
or U16342 (N_16342,N_15758,N_15793);
xnor U16343 (N_16343,N_15948,N_16163);
xor U16344 (N_16344,N_15836,N_15978);
xnor U16345 (N_16345,N_15907,N_16186);
and U16346 (N_16346,N_15896,N_15917);
and U16347 (N_16347,N_15814,N_15869);
nand U16348 (N_16348,N_16214,N_15999);
xnor U16349 (N_16349,N_16184,N_16138);
nand U16350 (N_16350,N_15742,N_16220);
nand U16351 (N_16351,N_16177,N_15850);
nand U16352 (N_16352,N_16215,N_16052);
xor U16353 (N_16353,N_15756,N_16016);
nor U16354 (N_16354,N_15676,N_15732);
xor U16355 (N_16355,N_16004,N_15853);
or U16356 (N_16356,N_16027,N_15772);
nor U16357 (N_16357,N_16209,N_15961);
nor U16358 (N_16358,N_16010,N_16106);
and U16359 (N_16359,N_16231,N_16040);
or U16360 (N_16360,N_15746,N_15863);
nor U16361 (N_16361,N_15955,N_16051);
nand U16362 (N_16362,N_15757,N_16034);
nand U16363 (N_16363,N_15868,N_16121);
xnor U16364 (N_16364,N_15716,N_16005);
and U16365 (N_16365,N_15977,N_16109);
or U16366 (N_16366,N_16245,N_15901);
nand U16367 (N_16367,N_16217,N_15679);
nor U16368 (N_16368,N_15965,N_15991);
nand U16369 (N_16369,N_15747,N_15798);
or U16370 (N_16370,N_16167,N_16227);
nor U16371 (N_16371,N_16155,N_15810);
nor U16372 (N_16372,N_15754,N_15992);
nor U16373 (N_16373,N_15723,N_15971);
and U16374 (N_16374,N_15931,N_15930);
nor U16375 (N_16375,N_15944,N_15736);
and U16376 (N_16376,N_15703,N_15653);
xor U16377 (N_16377,N_15942,N_16205);
xor U16378 (N_16378,N_15890,N_16084);
and U16379 (N_16379,N_16154,N_16095);
and U16380 (N_16380,N_16247,N_15635);
or U16381 (N_16381,N_16123,N_15963);
or U16382 (N_16382,N_15897,N_15686);
xor U16383 (N_16383,N_16229,N_16192);
nor U16384 (N_16384,N_15646,N_16156);
nor U16385 (N_16385,N_15749,N_15981);
or U16386 (N_16386,N_15783,N_15782);
and U16387 (N_16387,N_16146,N_16173);
and U16388 (N_16388,N_16047,N_15821);
nand U16389 (N_16389,N_16031,N_16160);
and U16390 (N_16390,N_15809,N_16055);
or U16391 (N_16391,N_15744,N_15625);
or U16392 (N_16392,N_16238,N_16142);
nor U16393 (N_16393,N_15862,N_16024);
and U16394 (N_16394,N_16149,N_16157);
or U16395 (N_16395,N_15962,N_15794);
nand U16396 (N_16396,N_15640,N_16067);
nand U16397 (N_16397,N_15698,N_16100);
or U16398 (N_16398,N_15832,N_16233);
and U16399 (N_16399,N_15988,N_15874);
xor U16400 (N_16400,N_15678,N_15706);
xor U16401 (N_16401,N_16096,N_15730);
nor U16402 (N_16402,N_15745,N_16097);
nand U16403 (N_16403,N_16039,N_15910);
xnor U16404 (N_16404,N_15713,N_15987);
or U16405 (N_16405,N_15704,N_15829);
xnor U16406 (N_16406,N_16033,N_15781);
nand U16407 (N_16407,N_15709,N_15633);
or U16408 (N_16408,N_16013,N_16196);
or U16409 (N_16409,N_16043,N_16158);
or U16410 (N_16410,N_15825,N_15926);
nor U16411 (N_16411,N_15911,N_16078);
nor U16412 (N_16412,N_15788,N_15909);
nand U16413 (N_16413,N_16062,N_15630);
or U16414 (N_16414,N_16117,N_15860);
nand U16415 (N_16415,N_15984,N_16011);
xor U16416 (N_16416,N_16119,N_15900);
and U16417 (N_16417,N_15714,N_15919);
nor U16418 (N_16418,N_15876,N_16075);
xnor U16419 (N_16419,N_16144,N_16103);
nand U16420 (N_16420,N_16107,N_16206);
nor U16421 (N_16421,N_16150,N_15771);
nand U16422 (N_16422,N_15936,N_15690);
xnor U16423 (N_16423,N_15887,N_16178);
nand U16424 (N_16424,N_16171,N_15697);
and U16425 (N_16425,N_15717,N_16065);
and U16426 (N_16426,N_15718,N_15939);
xnor U16427 (N_16427,N_15950,N_16223);
or U16428 (N_16428,N_16187,N_15787);
and U16429 (N_16429,N_15733,N_15729);
or U16430 (N_16430,N_16042,N_16089);
and U16431 (N_16431,N_16242,N_16151);
nor U16432 (N_16432,N_15969,N_15766);
nor U16433 (N_16433,N_15791,N_16122);
nand U16434 (N_16434,N_15765,N_15731);
nor U16435 (N_16435,N_15768,N_16112);
nor U16436 (N_16436,N_16162,N_16087);
xnor U16437 (N_16437,N_15854,N_16057);
or U16438 (N_16438,N_15952,N_16091);
or U16439 (N_16439,N_16199,N_15975);
nand U16440 (N_16440,N_15959,N_15786);
nor U16441 (N_16441,N_15638,N_15737);
nor U16442 (N_16442,N_15865,N_15888);
nand U16443 (N_16443,N_16022,N_15705);
and U16444 (N_16444,N_15958,N_15892);
and U16445 (N_16445,N_16079,N_15906);
nand U16446 (N_16446,N_16226,N_16222);
nor U16447 (N_16447,N_16085,N_15779);
xor U16448 (N_16448,N_15848,N_16015);
xnor U16449 (N_16449,N_15835,N_15903);
nor U16450 (N_16450,N_16239,N_15799);
and U16451 (N_16451,N_16183,N_15943);
nand U16452 (N_16452,N_16166,N_15968);
or U16453 (N_16453,N_16248,N_16086);
and U16454 (N_16454,N_15871,N_15727);
nand U16455 (N_16455,N_15990,N_16202);
nand U16456 (N_16456,N_15957,N_15629);
and U16457 (N_16457,N_15974,N_16131);
and U16458 (N_16458,N_15989,N_16020);
xor U16459 (N_16459,N_15985,N_15748);
xor U16460 (N_16460,N_16069,N_15660);
nor U16461 (N_16461,N_16064,N_15728);
xor U16462 (N_16462,N_15895,N_15841);
nor U16463 (N_16463,N_15883,N_16232);
nand U16464 (N_16464,N_16207,N_15699);
nand U16465 (N_16465,N_15966,N_16216);
nand U16466 (N_16466,N_15880,N_15675);
or U16467 (N_16467,N_15760,N_16133);
and U16468 (N_16468,N_16045,N_16203);
xor U16469 (N_16469,N_15845,N_16090);
nor U16470 (N_16470,N_15847,N_15954);
and U16471 (N_16471,N_16025,N_16190);
nor U16472 (N_16472,N_16240,N_15643);
nand U16473 (N_16473,N_16139,N_15651);
nor U16474 (N_16474,N_16164,N_15993);
or U16475 (N_16475,N_16115,N_15687);
and U16476 (N_16476,N_15665,N_15956);
and U16477 (N_16477,N_15824,N_16127);
nor U16478 (N_16478,N_15891,N_16088);
xor U16479 (N_16479,N_15654,N_15724);
nand U16480 (N_16480,N_15639,N_16073);
or U16481 (N_16481,N_16125,N_15998);
xor U16482 (N_16482,N_15680,N_16169);
nand U16483 (N_16483,N_15889,N_16049);
nand U16484 (N_16484,N_15933,N_16145);
and U16485 (N_16485,N_16218,N_16054);
nor U16486 (N_16486,N_16134,N_15715);
nor U16487 (N_16487,N_15964,N_15842);
and U16488 (N_16488,N_16003,N_16082);
or U16489 (N_16489,N_16148,N_15878);
nor U16490 (N_16490,N_15750,N_15818);
nor U16491 (N_16491,N_15685,N_16140);
xor U16492 (N_16492,N_15764,N_15655);
and U16493 (N_16493,N_16130,N_16006);
nor U16494 (N_16494,N_15904,N_15792);
or U16495 (N_16495,N_16030,N_15778);
and U16496 (N_16496,N_15642,N_15898);
or U16497 (N_16497,N_16021,N_15650);
nand U16498 (N_16498,N_16009,N_16189);
nor U16499 (N_16499,N_15852,N_15773);
xnor U16500 (N_16500,N_15661,N_15857);
xnor U16501 (N_16501,N_15881,N_16241);
nor U16502 (N_16502,N_15953,N_15631);
or U16503 (N_16503,N_16092,N_15929);
nand U16504 (N_16504,N_15879,N_15804);
nand U16505 (N_16505,N_16188,N_16135);
nand U16506 (N_16506,N_15924,N_16093);
or U16507 (N_16507,N_16246,N_16070);
nand U16508 (N_16508,N_15632,N_15935);
nand U16509 (N_16509,N_16210,N_15801);
and U16510 (N_16510,N_16111,N_16224);
or U16511 (N_16511,N_15972,N_16143);
nand U16512 (N_16512,N_15741,N_15681);
nor U16513 (N_16513,N_15806,N_15902);
nor U16514 (N_16514,N_15851,N_16170);
or U16515 (N_16515,N_15967,N_16147);
nand U16516 (N_16516,N_15645,N_15979);
or U16517 (N_16517,N_16198,N_15710);
xnor U16518 (N_16518,N_15976,N_16124);
and U16519 (N_16519,N_16114,N_15834);
xor U16520 (N_16520,N_15996,N_15815);
nand U16521 (N_16521,N_15994,N_15693);
nand U16522 (N_16522,N_15743,N_15813);
xnor U16523 (N_16523,N_15805,N_16235);
xnor U16524 (N_16524,N_16185,N_15669);
xor U16525 (N_16525,N_16061,N_15739);
and U16526 (N_16526,N_15921,N_15843);
and U16527 (N_16527,N_16212,N_15683);
or U16528 (N_16528,N_16113,N_15823);
and U16529 (N_16529,N_15763,N_15770);
and U16530 (N_16530,N_16195,N_16204);
xnor U16531 (N_16531,N_16211,N_15753);
nand U16532 (N_16532,N_15700,N_15725);
xnor U16533 (N_16533,N_16014,N_15652);
xnor U16534 (N_16534,N_15735,N_16002);
nand U16535 (N_16535,N_15882,N_15769);
nor U16536 (N_16536,N_15811,N_15670);
and U16537 (N_16537,N_16050,N_15830);
or U16538 (N_16538,N_15872,N_15738);
nor U16539 (N_16539,N_15762,N_15712);
nand U16540 (N_16540,N_15722,N_15691);
nor U16541 (N_16541,N_15908,N_16028);
or U16542 (N_16542,N_15983,N_15837);
nand U16543 (N_16543,N_16029,N_16102);
xor U16544 (N_16544,N_15870,N_16153);
or U16545 (N_16545,N_16066,N_15707);
nand U16546 (N_16546,N_15634,N_15755);
and U16547 (N_16547,N_16176,N_16159);
nand U16548 (N_16548,N_15856,N_16036);
and U16549 (N_16549,N_15855,N_15947);
or U16550 (N_16550,N_16137,N_15807);
nand U16551 (N_16551,N_15894,N_15858);
and U16552 (N_16552,N_16105,N_15949);
or U16553 (N_16553,N_16244,N_15913);
xor U16554 (N_16554,N_16032,N_15831);
nor U16555 (N_16555,N_15784,N_16035);
or U16556 (N_16556,N_16230,N_15667);
or U16557 (N_16557,N_15644,N_16063);
or U16558 (N_16558,N_15774,N_15695);
and U16559 (N_16559,N_15861,N_15899);
nand U16560 (N_16560,N_16175,N_16191);
nor U16561 (N_16561,N_15982,N_15777);
nor U16562 (N_16562,N_16116,N_16071);
nand U16563 (N_16563,N_15861,N_15973);
and U16564 (N_16564,N_16113,N_15782);
or U16565 (N_16565,N_15675,N_15698);
xnor U16566 (N_16566,N_15669,N_16017);
nor U16567 (N_16567,N_15743,N_15699);
xor U16568 (N_16568,N_15815,N_15831);
or U16569 (N_16569,N_15650,N_15819);
nand U16570 (N_16570,N_16183,N_15886);
nand U16571 (N_16571,N_15749,N_16231);
and U16572 (N_16572,N_15861,N_15784);
nand U16573 (N_16573,N_15632,N_15808);
and U16574 (N_16574,N_15795,N_16166);
or U16575 (N_16575,N_16099,N_15895);
or U16576 (N_16576,N_15691,N_15719);
nand U16577 (N_16577,N_16094,N_16200);
or U16578 (N_16578,N_16054,N_15975);
or U16579 (N_16579,N_15782,N_15720);
and U16580 (N_16580,N_15941,N_15879);
nand U16581 (N_16581,N_16012,N_15643);
and U16582 (N_16582,N_16154,N_15737);
or U16583 (N_16583,N_16066,N_16006);
or U16584 (N_16584,N_16152,N_16190);
xnor U16585 (N_16585,N_15683,N_15871);
nor U16586 (N_16586,N_15850,N_15971);
or U16587 (N_16587,N_16080,N_15685);
xnor U16588 (N_16588,N_16082,N_16066);
nand U16589 (N_16589,N_16165,N_16139);
and U16590 (N_16590,N_15677,N_16248);
or U16591 (N_16591,N_16014,N_15897);
and U16592 (N_16592,N_15774,N_15643);
or U16593 (N_16593,N_15649,N_16169);
and U16594 (N_16594,N_15964,N_16244);
or U16595 (N_16595,N_16235,N_16131);
nor U16596 (N_16596,N_16030,N_15699);
and U16597 (N_16597,N_15702,N_16185);
xnor U16598 (N_16598,N_15941,N_15981);
nand U16599 (N_16599,N_15804,N_16037);
nor U16600 (N_16600,N_15917,N_15711);
nand U16601 (N_16601,N_16012,N_15725);
and U16602 (N_16602,N_15760,N_16182);
and U16603 (N_16603,N_15946,N_16235);
and U16604 (N_16604,N_15874,N_15786);
or U16605 (N_16605,N_16151,N_16055);
or U16606 (N_16606,N_15824,N_15961);
xor U16607 (N_16607,N_16181,N_15731);
xnor U16608 (N_16608,N_15756,N_15674);
or U16609 (N_16609,N_16081,N_16064);
nor U16610 (N_16610,N_16199,N_15820);
xor U16611 (N_16611,N_15664,N_15817);
nor U16612 (N_16612,N_16072,N_15736);
xnor U16613 (N_16613,N_16073,N_15954);
nor U16614 (N_16614,N_15944,N_15959);
or U16615 (N_16615,N_16199,N_15694);
nor U16616 (N_16616,N_16136,N_15632);
nand U16617 (N_16617,N_16179,N_15885);
and U16618 (N_16618,N_15634,N_16198);
nor U16619 (N_16619,N_15813,N_15763);
or U16620 (N_16620,N_16070,N_15854);
nand U16621 (N_16621,N_15771,N_15625);
or U16622 (N_16622,N_15999,N_15681);
xor U16623 (N_16623,N_16205,N_16246);
nor U16624 (N_16624,N_16072,N_15872);
or U16625 (N_16625,N_15818,N_15925);
or U16626 (N_16626,N_15656,N_15976);
nor U16627 (N_16627,N_16119,N_16183);
nand U16628 (N_16628,N_15808,N_15734);
nand U16629 (N_16629,N_16190,N_15649);
and U16630 (N_16630,N_15860,N_16053);
nor U16631 (N_16631,N_15794,N_16136);
nor U16632 (N_16632,N_15958,N_16231);
and U16633 (N_16633,N_15906,N_16095);
or U16634 (N_16634,N_15758,N_16049);
xor U16635 (N_16635,N_16103,N_15944);
nor U16636 (N_16636,N_16176,N_15971);
nand U16637 (N_16637,N_16156,N_16205);
nor U16638 (N_16638,N_15660,N_15664);
nor U16639 (N_16639,N_16137,N_15846);
or U16640 (N_16640,N_15845,N_15856);
xor U16641 (N_16641,N_15914,N_16202);
and U16642 (N_16642,N_16113,N_15655);
and U16643 (N_16643,N_16054,N_16141);
nand U16644 (N_16644,N_16059,N_15863);
nand U16645 (N_16645,N_15827,N_15886);
nand U16646 (N_16646,N_16072,N_15821);
nor U16647 (N_16647,N_15720,N_15894);
and U16648 (N_16648,N_16225,N_15887);
and U16649 (N_16649,N_16017,N_16050);
nor U16650 (N_16650,N_16241,N_15951);
or U16651 (N_16651,N_16097,N_16185);
nand U16652 (N_16652,N_16217,N_16229);
nor U16653 (N_16653,N_16097,N_15968);
xor U16654 (N_16654,N_16163,N_15857);
xor U16655 (N_16655,N_15730,N_15806);
nand U16656 (N_16656,N_15890,N_15876);
nand U16657 (N_16657,N_15679,N_15671);
nor U16658 (N_16658,N_15808,N_15822);
or U16659 (N_16659,N_15730,N_16017);
xor U16660 (N_16660,N_15789,N_16192);
nand U16661 (N_16661,N_15899,N_15660);
nor U16662 (N_16662,N_15645,N_15773);
xnor U16663 (N_16663,N_15698,N_16233);
or U16664 (N_16664,N_16188,N_16067);
and U16665 (N_16665,N_15757,N_15906);
and U16666 (N_16666,N_15840,N_15723);
nand U16667 (N_16667,N_15961,N_15759);
or U16668 (N_16668,N_15799,N_16104);
nand U16669 (N_16669,N_15643,N_16088);
or U16670 (N_16670,N_15832,N_15711);
xnor U16671 (N_16671,N_15848,N_15717);
xor U16672 (N_16672,N_16074,N_16081);
or U16673 (N_16673,N_15917,N_16181);
and U16674 (N_16674,N_15626,N_16094);
xor U16675 (N_16675,N_16072,N_15752);
nor U16676 (N_16676,N_16070,N_15879);
xnor U16677 (N_16677,N_15787,N_15922);
nand U16678 (N_16678,N_16097,N_16035);
or U16679 (N_16679,N_15905,N_16191);
nor U16680 (N_16680,N_15655,N_15646);
or U16681 (N_16681,N_15632,N_15799);
nor U16682 (N_16682,N_15872,N_15910);
nand U16683 (N_16683,N_15952,N_16185);
and U16684 (N_16684,N_15937,N_15812);
nand U16685 (N_16685,N_16123,N_15809);
nand U16686 (N_16686,N_15810,N_15961);
xor U16687 (N_16687,N_16119,N_16230);
nand U16688 (N_16688,N_16123,N_15820);
xnor U16689 (N_16689,N_15772,N_15988);
nand U16690 (N_16690,N_15727,N_16246);
nor U16691 (N_16691,N_15892,N_15837);
or U16692 (N_16692,N_15785,N_15673);
xor U16693 (N_16693,N_15897,N_16210);
and U16694 (N_16694,N_16218,N_15737);
nor U16695 (N_16695,N_15782,N_16178);
or U16696 (N_16696,N_15794,N_16209);
nand U16697 (N_16697,N_16006,N_16093);
nand U16698 (N_16698,N_16009,N_15625);
nand U16699 (N_16699,N_15767,N_15644);
xor U16700 (N_16700,N_16209,N_16150);
xor U16701 (N_16701,N_15810,N_16242);
or U16702 (N_16702,N_16027,N_16108);
and U16703 (N_16703,N_15842,N_15836);
xnor U16704 (N_16704,N_16207,N_15907);
xor U16705 (N_16705,N_15765,N_16176);
and U16706 (N_16706,N_16048,N_16060);
xnor U16707 (N_16707,N_16230,N_15815);
nand U16708 (N_16708,N_16234,N_15917);
nand U16709 (N_16709,N_15983,N_15834);
or U16710 (N_16710,N_15983,N_15955);
or U16711 (N_16711,N_16017,N_15784);
nand U16712 (N_16712,N_15849,N_15895);
xnor U16713 (N_16713,N_15627,N_15936);
xor U16714 (N_16714,N_16203,N_15650);
nor U16715 (N_16715,N_15738,N_16189);
nand U16716 (N_16716,N_15983,N_15704);
xnor U16717 (N_16717,N_16216,N_15858);
and U16718 (N_16718,N_15738,N_15664);
and U16719 (N_16719,N_16240,N_16201);
nor U16720 (N_16720,N_16179,N_16082);
nor U16721 (N_16721,N_15987,N_16102);
nand U16722 (N_16722,N_15756,N_16020);
xnor U16723 (N_16723,N_16187,N_15713);
nor U16724 (N_16724,N_15801,N_15870);
xor U16725 (N_16725,N_16049,N_16022);
nor U16726 (N_16726,N_15636,N_16116);
xor U16727 (N_16727,N_15862,N_16080);
xor U16728 (N_16728,N_16028,N_16056);
xor U16729 (N_16729,N_15888,N_15802);
or U16730 (N_16730,N_15744,N_16010);
or U16731 (N_16731,N_15836,N_15718);
xor U16732 (N_16732,N_15754,N_16227);
xor U16733 (N_16733,N_15824,N_15653);
or U16734 (N_16734,N_15923,N_15658);
and U16735 (N_16735,N_15842,N_15924);
and U16736 (N_16736,N_16108,N_16174);
or U16737 (N_16737,N_15681,N_15627);
and U16738 (N_16738,N_16036,N_16186);
nor U16739 (N_16739,N_16172,N_16097);
xnor U16740 (N_16740,N_15691,N_16082);
and U16741 (N_16741,N_15932,N_15713);
nand U16742 (N_16742,N_15659,N_15954);
xor U16743 (N_16743,N_15668,N_15746);
or U16744 (N_16744,N_16244,N_15732);
nand U16745 (N_16745,N_15911,N_16161);
nand U16746 (N_16746,N_16219,N_16159);
nand U16747 (N_16747,N_15908,N_15885);
xor U16748 (N_16748,N_16073,N_16178);
and U16749 (N_16749,N_16045,N_15740);
and U16750 (N_16750,N_16213,N_15900);
xnor U16751 (N_16751,N_15732,N_15716);
nand U16752 (N_16752,N_16074,N_15793);
xor U16753 (N_16753,N_15995,N_15642);
nor U16754 (N_16754,N_15751,N_15738);
and U16755 (N_16755,N_15933,N_16169);
or U16756 (N_16756,N_16188,N_16230);
xnor U16757 (N_16757,N_16087,N_16153);
or U16758 (N_16758,N_15920,N_16001);
or U16759 (N_16759,N_16139,N_16075);
nor U16760 (N_16760,N_15730,N_15913);
or U16761 (N_16761,N_15836,N_15972);
xor U16762 (N_16762,N_15985,N_16009);
nand U16763 (N_16763,N_16025,N_15857);
or U16764 (N_16764,N_16194,N_16049);
and U16765 (N_16765,N_16005,N_15860);
nand U16766 (N_16766,N_15969,N_16031);
nand U16767 (N_16767,N_15861,N_16118);
nand U16768 (N_16768,N_15759,N_15936);
and U16769 (N_16769,N_15647,N_15715);
and U16770 (N_16770,N_16148,N_15688);
nor U16771 (N_16771,N_16169,N_16220);
or U16772 (N_16772,N_15850,N_16113);
nand U16773 (N_16773,N_15941,N_16164);
or U16774 (N_16774,N_16165,N_15965);
nand U16775 (N_16775,N_15989,N_16002);
nand U16776 (N_16776,N_15781,N_15963);
nor U16777 (N_16777,N_16134,N_15855);
nor U16778 (N_16778,N_16039,N_16211);
nor U16779 (N_16779,N_15872,N_15948);
and U16780 (N_16780,N_15689,N_15915);
and U16781 (N_16781,N_15970,N_16045);
nand U16782 (N_16782,N_15956,N_15916);
and U16783 (N_16783,N_16028,N_16230);
and U16784 (N_16784,N_16224,N_15996);
nand U16785 (N_16785,N_16086,N_16110);
xnor U16786 (N_16786,N_15903,N_16021);
nor U16787 (N_16787,N_15876,N_16157);
nand U16788 (N_16788,N_15784,N_16098);
and U16789 (N_16789,N_15849,N_15634);
nor U16790 (N_16790,N_15858,N_15767);
nor U16791 (N_16791,N_15796,N_15940);
nor U16792 (N_16792,N_15749,N_15791);
xnor U16793 (N_16793,N_16204,N_16205);
nand U16794 (N_16794,N_15770,N_15629);
nor U16795 (N_16795,N_15959,N_15968);
or U16796 (N_16796,N_15625,N_16137);
nand U16797 (N_16797,N_15711,N_15886);
nand U16798 (N_16798,N_16180,N_15744);
or U16799 (N_16799,N_16195,N_15922);
nand U16800 (N_16800,N_16081,N_15855);
nor U16801 (N_16801,N_16082,N_16114);
nand U16802 (N_16802,N_15673,N_16006);
xnor U16803 (N_16803,N_15781,N_15821);
nor U16804 (N_16804,N_15737,N_16075);
nand U16805 (N_16805,N_16025,N_16077);
or U16806 (N_16806,N_16056,N_16123);
nor U16807 (N_16807,N_16249,N_16163);
and U16808 (N_16808,N_15920,N_16051);
nand U16809 (N_16809,N_16159,N_15921);
xor U16810 (N_16810,N_15959,N_16231);
and U16811 (N_16811,N_15744,N_15844);
nand U16812 (N_16812,N_15859,N_16060);
and U16813 (N_16813,N_15793,N_15839);
nor U16814 (N_16814,N_16042,N_15874);
xnor U16815 (N_16815,N_16058,N_16025);
and U16816 (N_16816,N_15908,N_15836);
or U16817 (N_16817,N_15637,N_15962);
nand U16818 (N_16818,N_16187,N_15936);
and U16819 (N_16819,N_15891,N_15812);
xor U16820 (N_16820,N_15723,N_15976);
xor U16821 (N_16821,N_15824,N_15810);
xor U16822 (N_16822,N_15664,N_15890);
or U16823 (N_16823,N_16005,N_15986);
nand U16824 (N_16824,N_15768,N_15653);
and U16825 (N_16825,N_16177,N_16104);
nor U16826 (N_16826,N_15637,N_16248);
xnor U16827 (N_16827,N_16102,N_16139);
or U16828 (N_16828,N_15765,N_16112);
or U16829 (N_16829,N_15929,N_15999);
or U16830 (N_16830,N_16075,N_16245);
nand U16831 (N_16831,N_16175,N_16142);
or U16832 (N_16832,N_15962,N_16234);
or U16833 (N_16833,N_16032,N_15676);
and U16834 (N_16834,N_16103,N_15907);
or U16835 (N_16835,N_16206,N_15692);
and U16836 (N_16836,N_15684,N_16042);
xor U16837 (N_16837,N_15657,N_16050);
nand U16838 (N_16838,N_15788,N_15875);
xnor U16839 (N_16839,N_15806,N_16164);
xnor U16840 (N_16840,N_16148,N_16135);
xor U16841 (N_16841,N_16202,N_15950);
nor U16842 (N_16842,N_15871,N_15732);
xnor U16843 (N_16843,N_16181,N_16081);
and U16844 (N_16844,N_16212,N_15759);
xnor U16845 (N_16845,N_15804,N_16224);
or U16846 (N_16846,N_16049,N_15815);
nand U16847 (N_16847,N_15756,N_15981);
xor U16848 (N_16848,N_16192,N_15911);
and U16849 (N_16849,N_16147,N_15803);
xnor U16850 (N_16850,N_16029,N_15701);
xor U16851 (N_16851,N_16138,N_15849);
or U16852 (N_16852,N_16087,N_15655);
and U16853 (N_16853,N_16207,N_16124);
or U16854 (N_16854,N_16156,N_15640);
or U16855 (N_16855,N_16034,N_16047);
nand U16856 (N_16856,N_15641,N_15634);
xor U16857 (N_16857,N_16082,N_16192);
or U16858 (N_16858,N_15844,N_16092);
nand U16859 (N_16859,N_15987,N_16122);
and U16860 (N_16860,N_16028,N_15757);
and U16861 (N_16861,N_16094,N_16089);
and U16862 (N_16862,N_16025,N_16196);
and U16863 (N_16863,N_15735,N_15977);
or U16864 (N_16864,N_16232,N_16071);
or U16865 (N_16865,N_15700,N_15971);
nor U16866 (N_16866,N_15877,N_16109);
and U16867 (N_16867,N_16066,N_15852);
and U16868 (N_16868,N_16049,N_15635);
nor U16869 (N_16869,N_15711,N_15726);
and U16870 (N_16870,N_16116,N_16011);
and U16871 (N_16871,N_16002,N_15830);
or U16872 (N_16872,N_16151,N_16006);
xnor U16873 (N_16873,N_15749,N_15637);
and U16874 (N_16874,N_16018,N_15654);
nor U16875 (N_16875,N_16262,N_16849);
nand U16876 (N_16876,N_16792,N_16752);
and U16877 (N_16877,N_16345,N_16523);
nor U16878 (N_16878,N_16534,N_16348);
and U16879 (N_16879,N_16399,N_16826);
nor U16880 (N_16880,N_16822,N_16647);
nor U16881 (N_16881,N_16786,N_16535);
nand U16882 (N_16882,N_16868,N_16467);
nand U16883 (N_16883,N_16758,N_16430);
and U16884 (N_16884,N_16625,N_16725);
xnor U16885 (N_16885,N_16410,N_16843);
xnor U16886 (N_16886,N_16714,N_16325);
or U16887 (N_16887,N_16276,N_16766);
nand U16888 (N_16888,N_16602,N_16655);
nand U16889 (N_16889,N_16729,N_16308);
nor U16890 (N_16890,N_16596,N_16356);
or U16891 (N_16891,N_16414,N_16802);
nand U16892 (N_16892,N_16420,N_16586);
nor U16893 (N_16893,N_16608,N_16854);
and U16894 (N_16894,N_16491,N_16691);
xnor U16895 (N_16895,N_16605,N_16690);
nor U16896 (N_16896,N_16524,N_16657);
nor U16897 (N_16897,N_16400,N_16260);
nor U16898 (N_16898,N_16372,N_16552);
nand U16899 (N_16899,N_16342,N_16483);
xor U16900 (N_16900,N_16417,N_16263);
nand U16901 (N_16901,N_16307,N_16486);
nand U16902 (N_16902,N_16277,N_16546);
xnor U16903 (N_16903,N_16561,N_16509);
xnor U16904 (N_16904,N_16869,N_16795);
nor U16905 (N_16905,N_16812,N_16823);
nand U16906 (N_16906,N_16303,N_16451);
nand U16907 (N_16907,N_16753,N_16265);
nand U16908 (N_16908,N_16848,N_16540);
or U16909 (N_16909,N_16668,N_16858);
nor U16910 (N_16910,N_16692,N_16353);
nor U16911 (N_16911,N_16615,N_16403);
or U16912 (N_16912,N_16306,N_16512);
nand U16913 (N_16913,N_16489,N_16374);
or U16914 (N_16914,N_16623,N_16801);
or U16915 (N_16915,N_16847,N_16257);
xor U16916 (N_16916,N_16418,N_16548);
or U16917 (N_16917,N_16867,N_16677);
or U16918 (N_16918,N_16779,N_16568);
nand U16919 (N_16919,N_16631,N_16819);
or U16920 (N_16920,N_16354,N_16783);
or U16921 (N_16921,N_16375,N_16538);
nand U16922 (N_16922,N_16532,N_16737);
nand U16923 (N_16923,N_16385,N_16748);
xnor U16924 (N_16924,N_16699,N_16793);
and U16925 (N_16925,N_16810,N_16680);
or U16926 (N_16926,N_16593,N_16264);
nor U16927 (N_16927,N_16488,N_16870);
xor U16928 (N_16928,N_16554,N_16378);
nand U16929 (N_16929,N_16404,N_16284);
and U16930 (N_16930,N_16514,N_16381);
nor U16931 (N_16931,N_16515,N_16474);
nand U16932 (N_16932,N_16261,N_16569);
nand U16933 (N_16933,N_16445,N_16805);
nor U16934 (N_16934,N_16555,N_16721);
nor U16935 (N_16935,N_16824,N_16344);
or U16936 (N_16936,N_16630,N_16460);
or U16937 (N_16937,N_16709,N_16492);
and U16938 (N_16938,N_16457,N_16252);
and U16939 (N_16939,N_16706,N_16794);
and U16940 (N_16940,N_16545,N_16871);
nand U16941 (N_16941,N_16549,N_16856);
and U16942 (N_16942,N_16331,N_16635);
or U16943 (N_16943,N_16803,N_16556);
nand U16944 (N_16944,N_16351,N_16440);
xor U16945 (N_16945,N_16461,N_16448);
or U16946 (N_16946,N_16482,N_16831);
xor U16947 (N_16947,N_16639,N_16772);
xnor U16948 (N_16948,N_16411,N_16747);
and U16949 (N_16949,N_16499,N_16739);
nand U16950 (N_16950,N_16731,N_16860);
xor U16951 (N_16951,N_16872,N_16266);
and U16952 (N_16952,N_16578,N_16386);
nor U16953 (N_16953,N_16776,N_16336);
or U16954 (N_16954,N_16740,N_16666);
xor U16955 (N_16955,N_16478,N_16652);
xnor U16956 (N_16956,N_16357,N_16531);
and U16957 (N_16957,N_16727,N_16339);
nand U16958 (N_16958,N_16426,N_16840);
and U16959 (N_16959,N_16614,N_16624);
xor U16960 (N_16960,N_16703,N_16390);
or U16961 (N_16961,N_16821,N_16797);
nand U16962 (N_16962,N_16501,N_16251);
nor U16963 (N_16963,N_16255,N_16450);
or U16964 (N_16964,N_16723,N_16682);
and U16965 (N_16965,N_16687,N_16738);
nand U16966 (N_16966,N_16358,N_16695);
and U16967 (N_16967,N_16330,N_16628);
nor U16968 (N_16968,N_16784,N_16349);
xnor U16969 (N_16969,N_16564,N_16305);
nand U16970 (N_16970,N_16423,N_16328);
or U16971 (N_16971,N_16527,N_16744);
or U16972 (N_16972,N_16730,N_16487);
xor U16973 (N_16973,N_16434,N_16674);
or U16974 (N_16974,N_16800,N_16584);
nor U16975 (N_16975,N_16313,N_16780);
or U16976 (N_16976,N_16362,N_16466);
nor U16977 (N_16977,N_16866,N_16310);
nor U16978 (N_16978,N_16346,N_16459);
nand U16979 (N_16979,N_16807,N_16646);
xor U16980 (N_16980,N_16502,N_16394);
and U16981 (N_16981,N_16427,N_16708);
nor U16982 (N_16982,N_16409,N_16290);
nor U16983 (N_16983,N_16678,N_16382);
and U16984 (N_16984,N_16338,N_16672);
xnor U16985 (N_16985,N_16612,N_16464);
nor U16986 (N_16986,N_16283,N_16658);
and U16987 (N_16987,N_16413,N_16701);
and U16988 (N_16988,N_16317,N_16428);
or U16989 (N_16989,N_16376,N_16335);
nor U16990 (N_16990,N_16833,N_16609);
nor U16991 (N_16991,N_16551,N_16513);
and U16992 (N_16992,N_16799,N_16361);
xnor U16993 (N_16993,N_16688,N_16408);
xnor U16994 (N_16994,N_16256,N_16653);
nand U16995 (N_16995,N_16713,N_16476);
or U16996 (N_16996,N_16650,N_16846);
xnor U16997 (N_16997,N_16401,N_16663);
nand U16998 (N_16998,N_16304,N_16698);
or U16999 (N_16999,N_16528,N_16685);
xor U17000 (N_17000,N_16733,N_16267);
or U17001 (N_17001,N_16268,N_16425);
and U17002 (N_17002,N_16299,N_16371);
xor U17003 (N_17003,N_16302,N_16590);
nand U17004 (N_17004,N_16864,N_16493);
or U17005 (N_17005,N_16485,N_16446);
and U17006 (N_17006,N_16683,N_16562);
nand U17007 (N_17007,N_16717,N_16817);
xnor U17008 (N_17008,N_16391,N_16316);
nand U17009 (N_17009,N_16771,N_16785);
nand U17010 (N_17010,N_16533,N_16379);
and U17011 (N_17011,N_16599,N_16742);
and U17012 (N_17012,N_16757,N_16645);
xor U17013 (N_17013,N_16762,N_16640);
and U17014 (N_17014,N_16815,N_16566);
xnor U17015 (N_17015,N_16469,N_16377);
or U17016 (N_17016,N_16432,N_16874);
and U17017 (N_17017,N_16465,N_16670);
nand U17018 (N_17018,N_16788,N_16659);
nor U17019 (N_17019,N_16286,N_16292);
or U17020 (N_17020,N_16873,N_16664);
xor U17021 (N_17021,N_16836,N_16539);
nor U17022 (N_17022,N_16791,N_16694);
xor U17023 (N_17023,N_16570,N_16326);
nand U17024 (N_17024,N_16581,N_16705);
and U17025 (N_17025,N_16340,N_16301);
and U17026 (N_17026,N_16312,N_16720);
nor U17027 (N_17027,N_16818,N_16272);
nor U17028 (N_17028,N_16295,N_16521);
and U17029 (N_17029,N_16565,N_16603);
nor U17030 (N_17030,N_16366,N_16853);
xor U17031 (N_17031,N_16477,N_16796);
nor U17032 (N_17032,N_16406,N_16443);
and U17033 (N_17033,N_16452,N_16368);
xnor U17034 (N_17034,N_16337,N_16479);
and U17035 (N_17035,N_16436,N_16319);
nand U17036 (N_17036,N_16315,N_16275);
nand U17037 (N_17037,N_16588,N_16572);
xor U17038 (N_17038,N_16816,N_16484);
or U17039 (N_17039,N_16591,N_16827);
or U17040 (N_17040,N_16508,N_16547);
nand U17041 (N_17041,N_16447,N_16861);
nand U17042 (N_17042,N_16250,N_16396);
nor U17043 (N_17043,N_16577,N_16431);
nor U17044 (N_17044,N_16296,N_16288);
nand U17045 (N_17045,N_16322,N_16520);
and U17046 (N_17046,N_16610,N_16616);
xor U17047 (N_17047,N_16407,N_16468);
nand U17048 (N_17048,N_16595,N_16412);
or U17049 (N_17049,N_16617,N_16696);
and U17050 (N_17050,N_16768,N_16475);
nor U17051 (N_17051,N_16398,N_16458);
nand U17052 (N_17052,N_16712,N_16661);
xor U17053 (N_17053,N_16667,N_16838);
and U17054 (N_17054,N_16324,N_16829);
xnor U17055 (N_17055,N_16636,N_16370);
nand U17056 (N_17056,N_16669,N_16352);
xor U17057 (N_17057,N_16522,N_16632);
nand U17058 (N_17058,N_16654,N_16395);
or U17059 (N_17059,N_16571,N_16751);
nor U17060 (N_17060,N_16618,N_16297);
nand U17061 (N_17061,N_16318,N_16380);
nor U17062 (N_17062,N_16424,N_16773);
xor U17063 (N_17063,N_16804,N_16648);
nor U17064 (N_17064,N_16576,N_16660);
nor U17065 (N_17065,N_16834,N_16274);
and U17066 (N_17066,N_16765,N_16559);
and U17067 (N_17067,N_16530,N_16309);
or U17068 (N_17068,N_16763,N_16759);
and U17069 (N_17069,N_16835,N_16749);
and U17070 (N_17070,N_16294,N_16830);
nor U17071 (N_17071,N_16473,N_16585);
and U17072 (N_17072,N_16480,N_16845);
nand U17073 (N_17073,N_16393,N_16643);
and U17074 (N_17074,N_16259,N_16825);
nand U17075 (N_17075,N_16470,N_16675);
and U17076 (N_17076,N_16511,N_16433);
or U17077 (N_17077,N_16857,N_16702);
and U17078 (N_17078,N_16764,N_16504);
nand U17079 (N_17079,N_16620,N_16529);
xor U17080 (N_17080,N_16707,N_16525);
or U17081 (N_17081,N_16622,N_16711);
or U17082 (N_17082,N_16621,N_16364);
and U17083 (N_17083,N_16553,N_16582);
nand U17084 (N_17084,N_16679,N_16718);
nand U17085 (N_17085,N_16526,N_16472);
xnor U17086 (N_17086,N_16278,N_16597);
xor U17087 (N_17087,N_16397,N_16282);
and U17088 (N_17088,N_16323,N_16498);
nor U17089 (N_17089,N_16542,N_16269);
or U17090 (N_17090,N_16641,N_16777);
or U17091 (N_17091,N_16644,N_16289);
nor U17092 (N_17092,N_16629,N_16583);
nand U17093 (N_17093,N_16850,N_16419);
xor U17094 (N_17094,N_16392,N_16855);
xnor U17095 (N_17095,N_16347,N_16573);
nor U17096 (N_17096,N_16442,N_16732);
nand U17097 (N_17097,N_16681,N_16761);
and U17098 (N_17098,N_16518,N_16503);
xnor U17099 (N_17099,N_16550,N_16314);
xnor U17100 (N_17100,N_16359,N_16760);
or U17101 (N_17101,N_16500,N_16841);
xor U17102 (N_17102,N_16321,N_16716);
nor U17103 (N_17103,N_16592,N_16449);
nor U17104 (N_17104,N_16775,N_16367);
nand U17105 (N_17105,N_16580,N_16808);
nand U17106 (N_17106,N_16689,N_16291);
nor U17107 (N_17107,N_16563,N_16724);
or U17108 (N_17108,N_16384,N_16287);
nor U17109 (N_17109,N_16844,N_16589);
xor U17110 (N_17110,N_16416,N_16506);
nand U17111 (N_17111,N_16541,N_16662);
xnor U17112 (N_17112,N_16676,N_16741);
or U17113 (N_17113,N_16567,N_16402);
nor U17114 (N_17114,N_16462,N_16806);
nand U17115 (N_17115,N_16750,N_16642);
or U17116 (N_17116,N_16557,N_16544);
or U17117 (N_17117,N_16505,N_16728);
nor U17118 (N_17118,N_16481,N_16311);
xor U17119 (N_17119,N_16859,N_16365);
nand U17120 (N_17120,N_16516,N_16722);
nand U17121 (N_17121,N_16575,N_16471);
xor U17122 (N_17122,N_16363,N_16619);
nand U17123 (N_17123,N_16320,N_16726);
nor U17124 (N_17124,N_16334,N_16536);
nand U17125 (N_17125,N_16253,N_16719);
nand U17126 (N_17126,N_16754,N_16429);
xor U17127 (N_17127,N_16862,N_16778);
nand U17128 (N_17128,N_16496,N_16327);
and U17129 (N_17129,N_16579,N_16673);
xor U17130 (N_17130,N_16686,N_16280);
nand U17131 (N_17131,N_16254,N_16863);
and U17132 (N_17132,N_16270,N_16626);
xor U17133 (N_17133,N_16360,N_16734);
xnor U17134 (N_17134,N_16852,N_16537);
nand U17135 (N_17135,N_16439,N_16453);
and U17136 (N_17136,N_16560,N_16665);
nor U17137 (N_17137,N_16820,N_16837);
xor U17138 (N_17138,N_16355,N_16756);
nor U17139 (N_17139,N_16684,N_16293);
and U17140 (N_17140,N_16444,N_16627);
nor U17141 (N_17141,N_16715,N_16587);
and U17142 (N_17142,N_16273,N_16373);
or U17143 (N_17143,N_16774,N_16258);
nand U17144 (N_17144,N_16746,N_16405);
nor U17145 (N_17145,N_16332,N_16441);
nand U17146 (N_17146,N_16600,N_16745);
nand U17147 (N_17147,N_16769,N_16517);
and U17148 (N_17148,N_16755,N_16437);
xor U17149 (N_17149,N_16842,N_16832);
or U17150 (N_17150,N_16594,N_16607);
or U17151 (N_17151,N_16341,N_16387);
or U17152 (N_17152,N_16490,N_16497);
nor U17153 (N_17153,N_16415,N_16634);
and U17154 (N_17154,N_16422,N_16369);
xnor U17155 (N_17155,N_16507,N_16798);
or U17156 (N_17156,N_16298,N_16421);
or U17157 (N_17157,N_16454,N_16633);
nand U17158 (N_17158,N_16463,N_16651);
nand U17159 (N_17159,N_16604,N_16671);
xnor U17160 (N_17160,N_16789,N_16700);
or U17161 (N_17161,N_16601,N_16333);
or U17162 (N_17162,N_16781,N_16811);
and U17163 (N_17163,N_16329,N_16656);
xnor U17164 (N_17164,N_16828,N_16790);
and U17165 (N_17165,N_16736,N_16510);
or U17166 (N_17166,N_16574,N_16782);
or U17167 (N_17167,N_16389,N_16343);
or U17168 (N_17168,N_16638,N_16704);
nand U17169 (N_17169,N_16606,N_16285);
and U17170 (N_17170,N_16558,N_16735);
nor U17171 (N_17171,N_16649,N_16438);
and U17172 (N_17172,N_16767,N_16350);
and U17173 (N_17173,N_16388,N_16271);
xor U17174 (N_17174,N_16743,N_16839);
nor U17175 (N_17175,N_16865,N_16611);
xnor U17176 (N_17176,N_16598,N_16613);
nand U17177 (N_17177,N_16851,N_16809);
or U17178 (N_17178,N_16279,N_16519);
xor U17179 (N_17179,N_16435,N_16300);
and U17180 (N_17180,N_16813,N_16814);
nor U17181 (N_17181,N_16787,N_16770);
nand U17182 (N_17182,N_16455,N_16495);
nand U17183 (N_17183,N_16456,N_16697);
and U17184 (N_17184,N_16494,N_16281);
xor U17185 (N_17185,N_16383,N_16693);
nand U17186 (N_17186,N_16543,N_16637);
nand U17187 (N_17187,N_16710,N_16258);
xnor U17188 (N_17188,N_16465,N_16290);
xor U17189 (N_17189,N_16369,N_16293);
xnor U17190 (N_17190,N_16368,N_16578);
or U17191 (N_17191,N_16400,N_16489);
nor U17192 (N_17192,N_16858,N_16840);
nor U17193 (N_17193,N_16854,N_16871);
nand U17194 (N_17194,N_16252,N_16443);
nand U17195 (N_17195,N_16578,N_16620);
or U17196 (N_17196,N_16826,N_16675);
xor U17197 (N_17197,N_16254,N_16499);
nand U17198 (N_17198,N_16797,N_16397);
nand U17199 (N_17199,N_16396,N_16492);
nor U17200 (N_17200,N_16369,N_16619);
and U17201 (N_17201,N_16798,N_16575);
and U17202 (N_17202,N_16251,N_16488);
nor U17203 (N_17203,N_16808,N_16253);
nand U17204 (N_17204,N_16466,N_16271);
xnor U17205 (N_17205,N_16456,N_16282);
and U17206 (N_17206,N_16793,N_16476);
xnor U17207 (N_17207,N_16586,N_16677);
xnor U17208 (N_17208,N_16515,N_16397);
nand U17209 (N_17209,N_16443,N_16329);
and U17210 (N_17210,N_16432,N_16493);
xnor U17211 (N_17211,N_16439,N_16747);
or U17212 (N_17212,N_16824,N_16372);
nand U17213 (N_17213,N_16271,N_16325);
xnor U17214 (N_17214,N_16408,N_16359);
nand U17215 (N_17215,N_16849,N_16723);
or U17216 (N_17216,N_16826,N_16751);
and U17217 (N_17217,N_16544,N_16284);
and U17218 (N_17218,N_16808,N_16824);
nor U17219 (N_17219,N_16756,N_16411);
or U17220 (N_17220,N_16361,N_16812);
nor U17221 (N_17221,N_16325,N_16756);
or U17222 (N_17222,N_16792,N_16688);
xnor U17223 (N_17223,N_16386,N_16852);
nand U17224 (N_17224,N_16644,N_16814);
nor U17225 (N_17225,N_16512,N_16448);
nand U17226 (N_17226,N_16852,N_16383);
or U17227 (N_17227,N_16264,N_16603);
nor U17228 (N_17228,N_16749,N_16367);
nand U17229 (N_17229,N_16738,N_16382);
or U17230 (N_17230,N_16459,N_16464);
and U17231 (N_17231,N_16376,N_16603);
nand U17232 (N_17232,N_16730,N_16374);
nor U17233 (N_17233,N_16840,N_16621);
xnor U17234 (N_17234,N_16820,N_16432);
and U17235 (N_17235,N_16758,N_16280);
nand U17236 (N_17236,N_16380,N_16751);
nand U17237 (N_17237,N_16734,N_16679);
xor U17238 (N_17238,N_16864,N_16817);
nor U17239 (N_17239,N_16549,N_16431);
xor U17240 (N_17240,N_16411,N_16839);
xnor U17241 (N_17241,N_16627,N_16396);
and U17242 (N_17242,N_16316,N_16348);
xnor U17243 (N_17243,N_16513,N_16265);
nor U17244 (N_17244,N_16736,N_16581);
nor U17245 (N_17245,N_16404,N_16476);
or U17246 (N_17246,N_16276,N_16756);
and U17247 (N_17247,N_16812,N_16346);
or U17248 (N_17248,N_16602,N_16469);
nor U17249 (N_17249,N_16451,N_16399);
nor U17250 (N_17250,N_16476,N_16639);
and U17251 (N_17251,N_16356,N_16815);
xor U17252 (N_17252,N_16419,N_16413);
xnor U17253 (N_17253,N_16316,N_16466);
and U17254 (N_17254,N_16531,N_16631);
or U17255 (N_17255,N_16401,N_16768);
or U17256 (N_17256,N_16631,N_16786);
xnor U17257 (N_17257,N_16862,N_16759);
nand U17258 (N_17258,N_16763,N_16459);
xor U17259 (N_17259,N_16784,N_16680);
xnor U17260 (N_17260,N_16535,N_16296);
xor U17261 (N_17261,N_16863,N_16477);
nor U17262 (N_17262,N_16532,N_16819);
xor U17263 (N_17263,N_16444,N_16598);
xnor U17264 (N_17264,N_16722,N_16709);
or U17265 (N_17265,N_16604,N_16257);
nor U17266 (N_17266,N_16582,N_16276);
xor U17267 (N_17267,N_16340,N_16861);
nor U17268 (N_17268,N_16303,N_16690);
xnor U17269 (N_17269,N_16421,N_16252);
or U17270 (N_17270,N_16722,N_16466);
or U17271 (N_17271,N_16777,N_16415);
nor U17272 (N_17272,N_16306,N_16790);
and U17273 (N_17273,N_16272,N_16788);
nor U17274 (N_17274,N_16683,N_16812);
nand U17275 (N_17275,N_16554,N_16767);
nand U17276 (N_17276,N_16870,N_16352);
nand U17277 (N_17277,N_16571,N_16854);
and U17278 (N_17278,N_16400,N_16852);
nor U17279 (N_17279,N_16447,N_16518);
nor U17280 (N_17280,N_16839,N_16687);
and U17281 (N_17281,N_16593,N_16869);
xnor U17282 (N_17282,N_16291,N_16807);
nand U17283 (N_17283,N_16336,N_16375);
and U17284 (N_17284,N_16651,N_16300);
or U17285 (N_17285,N_16523,N_16540);
nor U17286 (N_17286,N_16582,N_16768);
nand U17287 (N_17287,N_16633,N_16327);
or U17288 (N_17288,N_16482,N_16266);
or U17289 (N_17289,N_16524,N_16353);
nor U17290 (N_17290,N_16377,N_16775);
or U17291 (N_17291,N_16397,N_16297);
nor U17292 (N_17292,N_16407,N_16443);
xnor U17293 (N_17293,N_16748,N_16566);
nor U17294 (N_17294,N_16448,N_16870);
and U17295 (N_17295,N_16449,N_16272);
xnor U17296 (N_17296,N_16252,N_16579);
or U17297 (N_17297,N_16819,N_16507);
or U17298 (N_17298,N_16759,N_16827);
nand U17299 (N_17299,N_16513,N_16469);
and U17300 (N_17300,N_16280,N_16386);
and U17301 (N_17301,N_16744,N_16660);
nor U17302 (N_17302,N_16718,N_16450);
xor U17303 (N_17303,N_16635,N_16793);
or U17304 (N_17304,N_16332,N_16600);
xnor U17305 (N_17305,N_16366,N_16453);
nand U17306 (N_17306,N_16835,N_16753);
xor U17307 (N_17307,N_16503,N_16871);
xor U17308 (N_17308,N_16696,N_16416);
xnor U17309 (N_17309,N_16615,N_16562);
or U17310 (N_17310,N_16788,N_16674);
or U17311 (N_17311,N_16863,N_16769);
xnor U17312 (N_17312,N_16345,N_16267);
nor U17313 (N_17313,N_16560,N_16355);
or U17314 (N_17314,N_16516,N_16530);
xnor U17315 (N_17315,N_16817,N_16389);
nand U17316 (N_17316,N_16496,N_16370);
xor U17317 (N_17317,N_16654,N_16446);
and U17318 (N_17318,N_16740,N_16272);
nor U17319 (N_17319,N_16373,N_16845);
or U17320 (N_17320,N_16479,N_16461);
and U17321 (N_17321,N_16834,N_16482);
nor U17322 (N_17322,N_16593,N_16458);
and U17323 (N_17323,N_16847,N_16743);
and U17324 (N_17324,N_16432,N_16532);
or U17325 (N_17325,N_16367,N_16656);
xnor U17326 (N_17326,N_16827,N_16424);
xor U17327 (N_17327,N_16288,N_16469);
nand U17328 (N_17328,N_16461,N_16671);
nor U17329 (N_17329,N_16356,N_16613);
or U17330 (N_17330,N_16366,N_16838);
xnor U17331 (N_17331,N_16357,N_16867);
and U17332 (N_17332,N_16756,N_16573);
and U17333 (N_17333,N_16859,N_16531);
nor U17334 (N_17334,N_16845,N_16417);
nand U17335 (N_17335,N_16654,N_16295);
and U17336 (N_17336,N_16600,N_16589);
nor U17337 (N_17337,N_16436,N_16549);
and U17338 (N_17338,N_16353,N_16438);
xnor U17339 (N_17339,N_16605,N_16367);
nand U17340 (N_17340,N_16445,N_16576);
or U17341 (N_17341,N_16355,N_16310);
nor U17342 (N_17342,N_16681,N_16851);
nor U17343 (N_17343,N_16290,N_16304);
nand U17344 (N_17344,N_16469,N_16666);
and U17345 (N_17345,N_16815,N_16512);
and U17346 (N_17346,N_16472,N_16275);
or U17347 (N_17347,N_16567,N_16519);
xor U17348 (N_17348,N_16477,N_16449);
and U17349 (N_17349,N_16462,N_16671);
or U17350 (N_17350,N_16608,N_16771);
and U17351 (N_17351,N_16791,N_16553);
and U17352 (N_17352,N_16328,N_16494);
nand U17353 (N_17353,N_16451,N_16266);
nand U17354 (N_17354,N_16775,N_16360);
xnor U17355 (N_17355,N_16572,N_16524);
xnor U17356 (N_17356,N_16610,N_16823);
or U17357 (N_17357,N_16585,N_16316);
or U17358 (N_17358,N_16722,N_16296);
and U17359 (N_17359,N_16582,N_16842);
or U17360 (N_17360,N_16325,N_16479);
nand U17361 (N_17361,N_16701,N_16845);
nand U17362 (N_17362,N_16711,N_16365);
and U17363 (N_17363,N_16308,N_16707);
and U17364 (N_17364,N_16515,N_16532);
nor U17365 (N_17365,N_16738,N_16639);
xor U17366 (N_17366,N_16438,N_16304);
and U17367 (N_17367,N_16408,N_16704);
or U17368 (N_17368,N_16526,N_16389);
nor U17369 (N_17369,N_16506,N_16526);
and U17370 (N_17370,N_16484,N_16720);
xor U17371 (N_17371,N_16643,N_16358);
or U17372 (N_17372,N_16688,N_16379);
nor U17373 (N_17373,N_16340,N_16638);
nand U17374 (N_17374,N_16370,N_16373);
nand U17375 (N_17375,N_16510,N_16361);
and U17376 (N_17376,N_16504,N_16360);
nand U17377 (N_17377,N_16572,N_16426);
xnor U17378 (N_17378,N_16409,N_16312);
or U17379 (N_17379,N_16273,N_16784);
or U17380 (N_17380,N_16835,N_16830);
and U17381 (N_17381,N_16380,N_16685);
or U17382 (N_17382,N_16863,N_16444);
nor U17383 (N_17383,N_16804,N_16666);
nand U17384 (N_17384,N_16342,N_16572);
and U17385 (N_17385,N_16651,N_16401);
nand U17386 (N_17386,N_16852,N_16436);
nor U17387 (N_17387,N_16419,N_16484);
nand U17388 (N_17388,N_16309,N_16793);
xor U17389 (N_17389,N_16597,N_16488);
nand U17390 (N_17390,N_16659,N_16611);
and U17391 (N_17391,N_16702,N_16286);
nand U17392 (N_17392,N_16529,N_16807);
xor U17393 (N_17393,N_16705,N_16334);
xor U17394 (N_17394,N_16716,N_16296);
nand U17395 (N_17395,N_16352,N_16696);
nand U17396 (N_17396,N_16374,N_16315);
nand U17397 (N_17397,N_16756,N_16843);
or U17398 (N_17398,N_16626,N_16845);
nand U17399 (N_17399,N_16423,N_16565);
and U17400 (N_17400,N_16866,N_16544);
and U17401 (N_17401,N_16736,N_16679);
nor U17402 (N_17402,N_16493,N_16507);
nand U17403 (N_17403,N_16678,N_16749);
and U17404 (N_17404,N_16574,N_16595);
xnor U17405 (N_17405,N_16366,N_16338);
nand U17406 (N_17406,N_16577,N_16481);
and U17407 (N_17407,N_16574,N_16317);
nand U17408 (N_17408,N_16282,N_16784);
nand U17409 (N_17409,N_16324,N_16828);
xor U17410 (N_17410,N_16459,N_16685);
or U17411 (N_17411,N_16602,N_16667);
nand U17412 (N_17412,N_16869,N_16305);
nand U17413 (N_17413,N_16298,N_16314);
xor U17414 (N_17414,N_16612,N_16295);
or U17415 (N_17415,N_16412,N_16383);
xnor U17416 (N_17416,N_16857,N_16730);
and U17417 (N_17417,N_16697,N_16450);
nor U17418 (N_17418,N_16391,N_16266);
and U17419 (N_17419,N_16557,N_16587);
nand U17420 (N_17420,N_16486,N_16447);
and U17421 (N_17421,N_16580,N_16849);
xor U17422 (N_17422,N_16421,N_16484);
or U17423 (N_17423,N_16399,N_16398);
nor U17424 (N_17424,N_16381,N_16636);
nand U17425 (N_17425,N_16583,N_16487);
nand U17426 (N_17426,N_16533,N_16410);
and U17427 (N_17427,N_16503,N_16687);
xor U17428 (N_17428,N_16852,N_16440);
nand U17429 (N_17429,N_16871,N_16713);
nor U17430 (N_17430,N_16851,N_16754);
or U17431 (N_17431,N_16467,N_16485);
or U17432 (N_17432,N_16620,N_16833);
nor U17433 (N_17433,N_16741,N_16611);
or U17434 (N_17434,N_16670,N_16716);
nor U17435 (N_17435,N_16559,N_16531);
and U17436 (N_17436,N_16803,N_16577);
nor U17437 (N_17437,N_16619,N_16691);
xor U17438 (N_17438,N_16368,N_16534);
nand U17439 (N_17439,N_16252,N_16544);
nand U17440 (N_17440,N_16828,N_16593);
or U17441 (N_17441,N_16506,N_16349);
xor U17442 (N_17442,N_16827,N_16833);
xnor U17443 (N_17443,N_16645,N_16631);
nor U17444 (N_17444,N_16388,N_16862);
nand U17445 (N_17445,N_16783,N_16578);
nor U17446 (N_17446,N_16772,N_16793);
nor U17447 (N_17447,N_16816,N_16459);
nor U17448 (N_17448,N_16825,N_16679);
xor U17449 (N_17449,N_16501,N_16739);
nand U17450 (N_17450,N_16408,N_16344);
or U17451 (N_17451,N_16722,N_16514);
nor U17452 (N_17452,N_16403,N_16821);
nand U17453 (N_17453,N_16344,N_16264);
or U17454 (N_17454,N_16767,N_16769);
nand U17455 (N_17455,N_16601,N_16761);
or U17456 (N_17456,N_16582,N_16429);
xnor U17457 (N_17457,N_16312,N_16519);
xor U17458 (N_17458,N_16651,N_16423);
or U17459 (N_17459,N_16405,N_16784);
or U17460 (N_17460,N_16595,N_16729);
or U17461 (N_17461,N_16401,N_16646);
nor U17462 (N_17462,N_16550,N_16288);
nand U17463 (N_17463,N_16754,N_16766);
nand U17464 (N_17464,N_16558,N_16274);
or U17465 (N_17465,N_16757,N_16651);
nor U17466 (N_17466,N_16701,N_16645);
nand U17467 (N_17467,N_16732,N_16859);
xnor U17468 (N_17468,N_16513,N_16385);
or U17469 (N_17469,N_16541,N_16626);
nand U17470 (N_17470,N_16324,N_16821);
nor U17471 (N_17471,N_16821,N_16251);
or U17472 (N_17472,N_16442,N_16676);
and U17473 (N_17473,N_16809,N_16436);
and U17474 (N_17474,N_16437,N_16280);
nor U17475 (N_17475,N_16768,N_16511);
xor U17476 (N_17476,N_16307,N_16330);
and U17477 (N_17477,N_16512,N_16863);
nand U17478 (N_17478,N_16802,N_16710);
xnor U17479 (N_17479,N_16553,N_16709);
nand U17480 (N_17480,N_16397,N_16833);
nor U17481 (N_17481,N_16822,N_16558);
or U17482 (N_17482,N_16798,N_16567);
nor U17483 (N_17483,N_16673,N_16352);
nand U17484 (N_17484,N_16411,N_16612);
nand U17485 (N_17485,N_16511,N_16421);
nand U17486 (N_17486,N_16597,N_16753);
or U17487 (N_17487,N_16796,N_16467);
nor U17488 (N_17488,N_16261,N_16590);
xnor U17489 (N_17489,N_16356,N_16523);
or U17490 (N_17490,N_16827,N_16713);
nand U17491 (N_17491,N_16466,N_16824);
or U17492 (N_17492,N_16787,N_16392);
nand U17493 (N_17493,N_16868,N_16518);
nand U17494 (N_17494,N_16835,N_16861);
xor U17495 (N_17495,N_16435,N_16521);
xnor U17496 (N_17496,N_16319,N_16775);
nand U17497 (N_17497,N_16576,N_16285);
xor U17498 (N_17498,N_16632,N_16653);
or U17499 (N_17499,N_16719,N_16461);
nor U17500 (N_17500,N_17101,N_17185);
and U17501 (N_17501,N_17052,N_17199);
nand U17502 (N_17502,N_16913,N_17079);
xor U17503 (N_17503,N_17462,N_17464);
and U17504 (N_17504,N_17339,N_17457);
xor U17505 (N_17505,N_17120,N_17121);
and U17506 (N_17506,N_17084,N_17206);
and U17507 (N_17507,N_17355,N_17393);
nand U17508 (N_17508,N_17481,N_17201);
nand U17509 (N_17509,N_17466,N_17423);
nor U17510 (N_17510,N_17492,N_16953);
and U17511 (N_17511,N_17286,N_16993);
and U17512 (N_17512,N_17277,N_16977);
nand U17513 (N_17513,N_16925,N_17032);
xnor U17514 (N_17514,N_17496,N_17318);
nor U17515 (N_17515,N_17219,N_16957);
and U17516 (N_17516,N_17227,N_16916);
and U17517 (N_17517,N_17241,N_17159);
and U17518 (N_17518,N_16894,N_17328);
xor U17519 (N_17519,N_17148,N_17461);
xor U17520 (N_17520,N_17158,N_17088);
and U17521 (N_17521,N_16958,N_16891);
or U17522 (N_17522,N_17107,N_17347);
or U17523 (N_17523,N_17261,N_17278);
nor U17524 (N_17524,N_17141,N_17443);
or U17525 (N_17525,N_16912,N_17291);
or U17526 (N_17526,N_17209,N_17060);
xnor U17527 (N_17527,N_17155,N_16908);
nand U17528 (N_17528,N_17388,N_16939);
or U17529 (N_17529,N_17190,N_16878);
and U17530 (N_17530,N_17086,N_17062);
nand U17531 (N_17531,N_17303,N_17389);
nand U17532 (N_17532,N_17354,N_17138);
nand U17533 (N_17533,N_17090,N_17267);
nand U17534 (N_17534,N_17013,N_17256);
nor U17535 (N_17535,N_17498,N_17372);
and U17536 (N_17536,N_17245,N_17030);
nor U17537 (N_17537,N_17401,N_17251);
and U17538 (N_17538,N_17011,N_17211);
and U17539 (N_17539,N_17285,N_16984);
and U17540 (N_17540,N_17330,N_17017);
and U17541 (N_17541,N_17234,N_16933);
nand U17542 (N_17542,N_16889,N_17273);
xnor U17543 (N_17543,N_17037,N_17447);
xor U17544 (N_17544,N_17175,N_17203);
xor U17545 (N_17545,N_17288,N_17078);
and U17546 (N_17546,N_16879,N_17123);
nor U17547 (N_17547,N_17276,N_17257);
nand U17548 (N_17548,N_17025,N_17191);
nand U17549 (N_17549,N_17322,N_17197);
nor U17550 (N_17550,N_16905,N_17095);
nand U17551 (N_17551,N_17394,N_16959);
and U17552 (N_17552,N_17207,N_17230);
nor U17553 (N_17553,N_17183,N_17452);
and U17554 (N_17554,N_17173,N_17387);
nor U17555 (N_17555,N_17246,N_17231);
and U17556 (N_17556,N_16962,N_16979);
or U17557 (N_17557,N_17048,N_16981);
nand U17558 (N_17558,N_16971,N_17218);
and U17559 (N_17559,N_17437,N_16972);
nand U17560 (N_17560,N_17365,N_17022);
nand U17561 (N_17561,N_17270,N_17043);
nand U17562 (N_17562,N_17317,N_17242);
nand U17563 (N_17563,N_17491,N_17152);
nand U17564 (N_17564,N_17340,N_17314);
nand U17565 (N_17565,N_17055,N_16915);
and U17566 (N_17566,N_17200,N_16928);
nand U17567 (N_17567,N_17254,N_17195);
or U17568 (N_17568,N_17140,N_17331);
xnor U17569 (N_17569,N_16999,N_17028);
nand U17570 (N_17570,N_17224,N_17091);
nor U17571 (N_17571,N_17327,N_17005);
nor U17572 (N_17572,N_17379,N_17012);
or U17573 (N_17573,N_17098,N_17410);
nor U17574 (N_17574,N_16927,N_17475);
and U17575 (N_17575,N_16918,N_17332);
nor U17576 (N_17576,N_17470,N_17264);
and U17577 (N_17577,N_17223,N_17336);
or U17578 (N_17578,N_17016,N_17417);
nor U17579 (N_17579,N_16934,N_16944);
xnor U17580 (N_17580,N_17193,N_16964);
or U17581 (N_17581,N_16976,N_17066);
or U17582 (N_17582,N_17194,N_16998);
nor U17583 (N_17583,N_17186,N_16883);
nor U17584 (N_17584,N_16911,N_17063);
and U17585 (N_17585,N_17479,N_16881);
or U17586 (N_17586,N_17050,N_17490);
nor U17587 (N_17587,N_17391,N_17212);
nand U17588 (N_17588,N_17471,N_17253);
or U17589 (N_17589,N_17036,N_17056);
nor U17590 (N_17590,N_17117,N_17071);
or U17591 (N_17591,N_17239,N_17020);
xor U17592 (N_17592,N_17029,N_17129);
and U17593 (N_17593,N_17236,N_17077);
and U17594 (N_17594,N_16922,N_17039);
and U17595 (N_17595,N_17405,N_17301);
nand U17596 (N_17596,N_17374,N_16965);
or U17597 (N_17597,N_17493,N_16986);
xnor U17598 (N_17598,N_17400,N_17100);
or U17599 (N_17599,N_17164,N_17358);
and U17600 (N_17600,N_16968,N_17179);
nand U17601 (N_17601,N_17220,N_17364);
and U17602 (N_17602,N_17381,N_17166);
nor U17603 (N_17603,N_17312,N_17484);
xor U17604 (N_17604,N_17404,N_17344);
nor U17605 (N_17605,N_17165,N_17263);
xnor U17606 (N_17606,N_16983,N_17049);
xnor U17607 (N_17607,N_17359,N_17161);
or U17608 (N_17608,N_17248,N_17403);
nand U17609 (N_17609,N_17109,N_17040);
and U17610 (N_17610,N_17237,N_17238);
and U17611 (N_17611,N_17311,N_17167);
and U17612 (N_17612,N_16956,N_17349);
or U17613 (N_17613,N_17127,N_16980);
nand U17614 (N_17614,N_17455,N_17162);
xnor U17615 (N_17615,N_17178,N_17142);
or U17616 (N_17616,N_17444,N_17059);
xnor U17617 (N_17617,N_17368,N_17177);
or U17618 (N_17618,N_16929,N_17292);
nand U17619 (N_17619,N_17143,N_16975);
xor U17620 (N_17620,N_17080,N_17135);
and U17621 (N_17621,N_17069,N_17181);
nand U17622 (N_17622,N_17448,N_17010);
and U17623 (N_17623,N_17441,N_17092);
xor U17624 (N_17624,N_17415,N_17021);
xor U17625 (N_17625,N_17478,N_17275);
or U17626 (N_17626,N_17395,N_17294);
nor U17627 (N_17627,N_17293,N_17385);
and U17628 (N_17628,N_17150,N_17382);
nand U17629 (N_17629,N_16909,N_16880);
xor U17630 (N_17630,N_17076,N_17124);
or U17631 (N_17631,N_16895,N_16949);
nor U17632 (N_17632,N_17134,N_17169);
nand U17633 (N_17633,N_17045,N_17260);
or U17634 (N_17634,N_17002,N_17074);
nor U17635 (N_17635,N_17065,N_17271);
or U17636 (N_17636,N_17073,N_17133);
and U17637 (N_17637,N_16945,N_17419);
or U17638 (N_17638,N_17182,N_16943);
nand U17639 (N_17639,N_17465,N_17420);
nor U17640 (N_17640,N_17422,N_17439);
xnor U17641 (N_17641,N_17371,N_17172);
or U17642 (N_17642,N_17108,N_17309);
xor U17643 (N_17643,N_17433,N_16936);
or U17644 (N_17644,N_17132,N_17126);
nand U17645 (N_17645,N_17287,N_17247);
and U17646 (N_17646,N_17310,N_16921);
xnor U17647 (N_17647,N_16969,N_17226);
nand U17648 (N_17648,N_17451,N_17054);
xor U17649 (N_17649,N_17110,N_17151);
and U17650 (N_17650,N_17214,N_17154);
xor U17651 (N_17651,N_16893,N_17337);
xnor U17652 (N_17652,N_17229,N_16950);
and U17653 (N_17653,N_17348,N_17325);
nand U17654 (N_17654,N_17118,N_17341);
or U17655 (N_17655,N_17192,N_17034);
or U17656 (N_17656,N_17035,N_17146);
or U17657 (N_17657,N_17367,N_16876);
xor U17658 (N_17658,N_17488,N_17407);
nand U17659 (N_17659,N_17042,N_17213);
and U17660 (N_17660,N_17087,N_17027);
nor U17661 (N_17661,N_17189,N_17357);
nor U17662 (N_17662,N_17431,N_16884);
or U17663 (N_17663,N_17047,N_17397);
xnor U17664 (N_17664,N_17305,N_16952);
xnor U17665 (N_17665,N_17473,N_17390);
nor U17666 (N_17666,N_17346,N_17250);
nor U17667 (N_17667,N_16995,N_17075);
or U17668 (N_17668,N_16937,N_17283);
xor U17669 (N_17669,N_17083,N_17157);
and U17670 (N_17670,N_17009,N_17103);
or U17671 (N_17671,N_16886,N_17085);
or U17672 (N_17672,N_17068,N_17072);
nor U17673 (N_17673,N_16892,N_16898);
or U17674 (N_17674,N_16966,N_17232);
or U17675 (N_17675,N_17061,N_16951);
and U17676 (N_17676,N_17064,N_17144);
xor U17677 (N_17677,N_17255,N_16938);
and U17678 (N_17678,N_16982,N_16994);
nor U17679 (N_17679,N_17244,N_17221);
or U17680 (N_17680,N_17398,N_17352);
nor U17681 (N_17681,N_17031,N_17435);
nor U17682 (N_17682,N_17014,N_17113);
nor U17683 (N_17683,N_17252,N_17188);
and U17684 (N_17684,N_17116,N_16985);
nand U17685 (N_17685,N_16978,N_17137);
nand U17686 (N_17686,N_16877,N_17122);
nand U17687 (N_17687,N_17233,N_17119);
nand U17688 (N_17688,N_17225,N_17460);
xor U17689 (N_17689,N_16946,N_17187);
and U17690 (N_17690,N_16903,N_16899);
xor U17691 (N_17691,N_17081,N_17326);
xor U17692 (N_17692,N_16923,N_17483);
and U17693 (N_17693,N_17295,N_17476);
and U17694 (N_17694,N_17089,N_17139);
xor U17695 (N_17695,N_17033,N_16890);
and U17696 (N_17696,N_17321,N_17006);
or U17697 (N_17697,N_17363,N_17297);
nor U17698 (N_17698,N_17243,N_16990);
nor U17699 (N_17699,N_17386,N_17442);
nor U17700 (N_17700,N_17411,N_17015);
nand U17701 (N_17701,N_17424,N_17338);
and U17702 (N_17702,N_16973,N_17174);
and U17703 (N_17703,N_17215,N_17376);
xnor U17704 (N_17704,N_17111,N_17004);
and U17705 (N_17705,N_17362,N_17485);
nand U17706 (N_17706,N_17313,N_17414);
nand U17707 (N_17707,N_17449,N_17105);
and U17708 (N_17708,N_17259,N_17114);
nand U17709 (N_17709,N_17196,N_16974);
and U17710 (N_17710,N_17216,N_17494);
and U17711 (N_17711,N_17380,N_16896);
nand U17712 (N_17712,N_17289,N_17003);
and U17713 (N_17713,N_17370,N_17041);
nor U17714 (N_17714,N_17279,N_16888);
and U17715 (N_17715,N_17269,N_16941);
or U17716 (N_17716,N_16924,N_17302);
xnor U17717 (N_17717,N_17290,N_17320);
nor U17718 (N_17718,N_17416,N_17168);
or U17719 (N_17719,N_17274,N_16882);
nor U17720 (N_17720,N_17459,N_17497);
nor U17721 (N_17721,N_17057,N_17115);
or U17722 (N_17722,N_17472,N_17499);
xor U17723 (N_17723,N_17335,N_17366);
nor U17724 (N_17724,N_17425,N_17184);
xnor U17725 (N_17725,N_16907,N_17298);
and U17726 (N_17726,N_16935,N_17130);
nand U17727 (N_17727,N_17044,N_17384);
nor U17728 (N_17728,N_16954,N_17268);
xnor U17729 (N_17729,N_17350,N_16930);
nor U17730 (N_17730,N_17217,N_17281);
nand U17731 (N_17731,N_17046,N_17205);
or U17732 (N_17732,N_17486,N_17378);
xor U17733 (N_17733,N_17453,N_17282);
or U17734 (N_17734,N_17323,N_17051);
nand U17735 (N_17735,N_16970,N_17440);
or U17736 (N_17736,N_17399,N_17334);
or U17737 (N_17737,N_16906,N_17429);
and U17738 (N_17738,N_17058,N_17128);
nor U17739 (N_17739,N_16897,N_17300);
nor U17740 (N_17740,N_17094,N_16961);
and U17741 (N_17741,N_16987,N_17007);
or U17742 (N_17742,N_17136,N_17019);
nand U17743 (N_17743,N_17023,N_17000);
nand U17744 (N_17744,N_16926,N_16920);
nand U17745 (N_17745,N_17067,N_17463);
nand U17746 (N_17746,N_17304,N_17333);
and U17747 (N_17747,N_17436,N_17106);
or U17748 (N_17748,N_17489,N_17383);
xor U17749 (N_17749,N_17147,N_17373);
nand U17750 (N_17750,N_17445,N_17038);
xnor U17751 (N_17751,N_16901,N_17171);
or U17752 (N_17752,N_17222,N_17480);
nand U17753 (N_17753,N_16989,N_17099);
or U17754 (N_17754,N_17208,N_17163);
nor U17755 (N_17755,N_17495,N_17375);
xnor U17756 (N_17756,N_17369,N_17026);
nor U17757 (N_17757,N_17249,N_17170);
nor U17758 (N_17758,N_17125,N_17024);
xnor U17759 (N_17759,N_17299,N_16887);
xnor U17760 (N_17760,N_17351,N_16917);
and U17761 (N_17761,N_17342,N_16919);
nor U17762 (N_17762,N_17458,N_17198);
nand U17763 (N_17763,N_17432,N_17306);
nor U17764 (N_17764,N_17353,N_17284);
and U17765 (N_17765,N_17396,N_16988);
or U17766 (N_17766,N_17426,N_17412);
nor U17767 (N_17767,N_16947,N_16967);
and U17768 (N_17768,N_17093,N_17240);
nor U17769 (N_17769,N_17377,N_17104);
or U17770 (N_17770,N_17324,N_17082);
nor U17771 (N_17771,N_16948,N_17053);
xor U17772 (N_17772,N_16902,N_17409);
and U17773 (N_17773,N_16996,N_17319);
nor U17774 (N_17774,N_16904,N_16900);
and U17775 (N_17775,N_16960,N_17430);
or U17776 (N_17776,N_17474,N_17112);
or U17777 (N_17777,N_17156,N_17070);
or U17778 (N_17778,N_16963,N_17131);
nor U17779 (N_17779,N_17018,N_17329);
nor U17780 (N_17780,N_16931,N_17202);
xnor U17781 (N_17781,N_17482,N_16991);
nor U17782 (N_17782,N_17446,N_16992);
or U17783 (N_17783,N_17356,N_17413);
nand U17784 (N_17784,N_17468,N_17272);
xor U17785 (N_17785,N_17427,N_17180);
nand U17786 (N_17786,N_16942,N_17160);
or U17787 (N_17787,N_17296,N_17467);
xor U17788 (N_17788,N_17450,N_17153);
or U17789 (N_17789,N_17361,N_17262);
xnor U17790 (N_17790,N_17307,N_17316);
nand U17791 (N_17791,N_17418,N_17392);
nand U17792 (N_17792,N_17345,N_17280);
xnor U17793 (N_17793,N_16940,N_16997);
nand U17794 (N_17794,N_17210,N_17408);
and U17795 (N_17795,N_17477,N_17315);
nand U17796 (N_17796,N_16910,N_17456);
and U17797 (N_17797,N_17228,N_17428);
nand U17798 (N_17798,N_17421,N_17487);
xnor U17799 (N_17799,N_17406,N_17097);
and U17800 (N_17800,N_17308,N_17149);
xor U17801 (N_17801,N_17204,N_17258);
nor U17802 (N_17802,N_16955,N_17096);
or U17803 (N_17803,N_17008,N_17343);
nor U17804 (N_17804,N_17102,N_17360);
and U17805 (N_17805,N_17265,N_16914);
or U17806 (N_17806,N_17001,N_17402);
and U17807 (N_17807,N_17434,N_17176);
xnor U17808 (N_17808,N_17145,N_17454);
nor U17809 (N_17809,N_17266,N_16932);
nand U17810 (N_17810,N_17235,N_17438);
xor U17811 (N_17811,N_16885,N_17469);
xnor U17812 (N_17812,N_16875,N_17377);
xnor U17813 (N_17813,N_17459,N_17038);
or U17814 (N_17814,N_17453,N_17249);
or U17815 (N_17815,N_17148,N_17033);
nor U17816 (N_17816,N_17492,N_17374);
or U17817 (N_17817,N_16915,N_17012);
xnor U17818 (N_17818,N_17324,N_17101);
nor U17819 (N_17819,N_16959,N_16975);
xor U17820 (N_17820,N_17099,N_17339);
nor U17821 (N_17821,N_17050,N_16991);
nor U17822 (N_17822,N_16914,N_17001);
nand U17823 (N_17823,N_16915,N_16951);
and U17824 (N_17824,N_17080,N_16897);
nand U17825 (N_17825,N_17129,N_17495);
nor U17826 (N_17826,N_17146,N_17132);
and U17827 (N_17827,N_17421,N_17295);
nand U17828 (N_17828,N_17082,N_17129);
xor U17829 (N_17829,N_17059,N_17381);
nor U17830 (N_17830,N_17387,N_17028);
nor U17831 (N_17831,N_17196,N_17045);
or U17832 (N_17832,N_17021,N_16965);
xnor U17833 (N_17833,N_17340,N_16959);
xnor U17834 (N_17834,N_17177,N_17495);
xnor U17835 (N_17835,N_17187,N_17358);
or U17836 (N_17836,N_17311,N_17140);
nor U17837 (N_17837,N_17231,N_17479);
nand U17838 (N_17838,N_17335,N_17442);
xor U17839 (N_17839,N_17280,N_16886);
nand U17840 (N_17840,N_17489,N_16905);
nand U17841 (N_17841,N_17467,N_16993);
or U17842 (N_17842,N_17078,N_17463);
and U17843 (N_17843,N_17326,N_17245);
xor U17844 (N_17844,N_17130,N_17220);
nand U17845 (N_17845,N_17499,N_16908);
and U17846 (N_17846,N_17205,N_17092);
and U17847 (N_17847,N_17289,N_17485);
nor U17848 (N_17848,N_17193,N_17210);
xnor U17849 (N_17849,N_17004,N_16883);
nor U17850 (N_17850,N_16961,N_17197);
nor U17851 (N_17851,N_17015,N_16905);
nor U17852 (N_17852,N_17320,N_17387);
or U17853 (N_17853,N_17372,N_17391);
or U17854 (N_17854,N_17183,N_17342);
xor U17855 (N_17855,N_17056,N_17224);
nor U17856 (N_17856,N_17464,N_16881);
nand U17857 (N_17857,N_17285,N_17404);
nand U17858 (N_17858,N_17227,N_17007);
and U17859 (N_17859,N_16912,N_16958);
nor U17860 (N_17860,N_17160,N_17410);
and U17861 (N_17861,N_17050,N_17491);
or U17862 (N_17862,N_17285,N_17042);
nand U17863 (N_17863,N_16946,N_16955);
xor U17864 (N_17864,N_17227,N_17280);
nor U17865 (N_17865,N_17385,N_16993);
or U17866 (N_17866,N_17007,N_17361);
nand U17867 (N_17867,N_17173,N_17181);
xor U17868 (N_17868,N_17249,N_17017);
xor U17869 (N_17869,N_16971,N_16975);
or U17870 (N_17870,N_17237,N_16981);
nand U17871 (N_17871,N_17337,N_17114);
or U17872 (N_17872,N_17372,N_16966);
xor U17873 (N_17873,N_17059,N_17393);
xnor U17874 (N_17874,N_17126,N_17466);
nand U17875 (N_17875,N_17062,N_17297);
nand U17876 (N_17876,N_16877,N_16901);
and U17877 (N_17877,N_16877,N_17014);
nand U17878 (N_17878,N_17457,N_17087);
and U17879 (N_17879,N_16915,N_17011);
or U17880 (N_17880,N_17281,N_17402);
nor U17881 (N_17881,N_16896,N_17326);
nand U17882 (N_17882,N_17342,N_17092);
and U17883 (N_17883,N_17264,N_17483);
or U17884 (N_17884,N_17116,N_17413);
and U17885 (N_17885,N_17024,N_17450);
nor U17886 (N_17886,N_17157,N_16947);
nor U17887 (N_17887,N_17234,N_17013);
and U17888 (N_17888,N_16946,N_17379);
and U17889 (N_17889,N_17153,N_17295);
xnor U17890 (N_17890,N_17070,N_16894);
nand U17891 (N_17891,N_16928,N_17126);
nor U17892 (N_17892,N_17394,N_16948);
nand U17893 (N_17893,N_17122,N_17395);
nor U17894 (N_17894,N_17488,N_16925);
nand U17895 (N_17895,N_17462,N_17150);
and U17896 (N_17896,N_17329,N_17395);
nand U17897 (N_17897,N_17392,N_17313);
or U17898 (N_17898,N_17240,N_17316);
xor U17899 (N_17899,N_17036,N_17011);
nand U17900 (N_17900,N_17292,N_16980);
nor U17901 (N_17901,N_17221,N_17358);
and U17902 (N_17902,N_17122,N_17437);
xnor U17903 (N_17903,N_17151,N_16947);
nand U17904 (N_17904,N_17280,N_16975);
or U17905 (N_17905,N_17233,N_17403);
nor U17906 (N_17906,N_17011,N_17352);
nor U17907 (N_17907,N_17041,N_17427);
and U17908 (N_17908,N_16950,N_17437);
and U17909 (N_17909,N_17356,N_17056);
nand U17910 (N_17910,N_17224,N_17214);
nor U17911 (N_17911,N_17439,N_17254);
nand U17912 (N_17912,N_17306,N_17019);
nor U17913 (N_17913,N_17160,N_17233);
nand U17914 (N_17914,N_16990,N_17357);
xor U17915 (N_17915,N_17355,N_17299);
and U17916 (N_17916,N_17086,N_17447);
and U17917 (N_17917,N_17034,N_16978);
xnor U17918 (N_17918,N_17340,N_17410);
xor U17919 (N_17919,N_17213,N_17115);
or U17920 (N_17920,N_17214,N_17345);
nand U17921 (N_17921,N_17245,N_17243);
xnor U17922 (N_17922,N_16924,N_17303);
and U17923 (N_17923,N_17465,N_17159);
or U17924 (N_17924,N_17296,N_17165);
or U17925 (N_17925,N_17317,N_17336);
xor U17926 (N_17926,N_16917,N_17297);
nor U17927 (N_17927,N_17193,N_17090);
nand U17928 (N_17928,N_17097,N_16953);
and U17929 (N_17929,N_17205,N_17254);
nand U17930 (N_17930,N_16932,N_17417);
nand U17931 (N_17931,N_17086,N_17434);
or U17932 (N_17932,N_17359,N_17265);
and U17933 (N_17933,N_16904,N_17023);
nand U17934 (N_17934,N_17058,N_17034);
xor U17935 (N_17935,N_16944,N_17276);
nand U17936 (N_17936,N_17152,N_17416);
or U17937 (N_17937,N_17293,N_17299);
or U17938 (N_17938,N_17498,N_17361);
xnor U17939 (N_17939,N_17054,N_17293);
xnor U17940 (N_17940,N_17109,N_17354);
nand U17941 (N_17941,N_17325,N_16883);
nand U17942 (N_17942,N_17086,N_17416);
and U17943 (N_17943,N_16939,N_17147);
or U17944 (N_17944,N_17251,N_17204);
nor U17945 (N_17945,N_17158,N_17125);
nand U17946 (N_17946,N_16994,N_17445);
or U17947 (N_17947,N_17390,N_16970);
or U17948 (N_17948,N_16991,N_17072);
nor U17949 (N_17949,N_16965,N_17451);
and U17950 (N_17950,N_17016,N_17248);
nand U17951 (N_17951,N_17065,N_17198);
or U17952 (N_17952,N_17488,N_17467);
nor U17953 (N_17953,N_17055,N_16881);
xor U17954 (N_17954,N_17297,N_17452);
nand U17955 (N_17955,N_17438,N_16888);
xor U17956 (N_17956,N_17012,N_17312);
or U17957 (N_17957,N_17412,N_16940);
nand U17958 (N_17958,N_17007,N_17338);
nor U17959 (N_17959,N_17164,N_17381);
or U17960 (N_17960,N_16992,N_16974);
xnor U17961 (N_17961,N_17159,N_17213);
and U17962 (N_17962,N_16909,N_17338);
xnor U17963 (N_17963,N_17319,N_17311);
xor U17964 (N_17964,N_16929,N_16943);
nor U17965 (N_17965,N_17006,N_17131);
and U17966 (N_17966,N_17039,N_17143);
nand U17967 (N_17967,N_17472,N_17314);
and U17968 (N_17968,N_16936,N_17270);
or U17969 (N_17969,N_17038,N_17119);
nor U17970 (N_17970,N_16877,N_17236);
xnor U17971 (N_17971,N_17320,N_17311);
xnor U17972 (N_17972,N_17226,N_17331);
nand U17973 (N_17973,N_17275,N_17201);
nor U17974 (N_17974,N_17431,N_17319);
and U17975 (N_17975,N_17231,N_17454);
nor U17976 (N_17976,N_17412,N_17203);
nand U17977 (N_17977,N_16985,N_17094);
or U17978 (N_17978,N_17003,N_17190);
nand U17979 (N_17979,N_17244,N_17251);
nor U17980 (N_17980,N_17373,N_17182);
nor U17981 (N_17981,N_17352,N_16904);
and U17982 (N_17982,N_17170,N_16898);
nor U17983 (N_17983,N_17106,N_17365);
and U17984 (N_17984,N_17218,N_17458);
and U17985 (N_17985,N_17395,N_16967);
nand U17986 (N_17986,N_17100,N_17039);
and U17987 (N_17987,N_17450,N_16967);
xnor U17988 (N_17988,N_16923,N_16890);
nand U17989 (N_17989,N_17277,N_17218);
and U17990 (N_17990,N_17477,N_17220);
and U17991 (N_17991,N_17170,N_17464);
or U17992 (N_17992,N_17041,N_17193);
xor U17993 (N_17993,N_17184,N_16916);
and U17994 (N_17994,N_17204,N_17375);
xor U17995 (N_17995,N_16976,N_17006);
and U17996 (N_17996,N_17124,N_17148);
or U17997 (N_17997,N_17474,N_17496);
or U17998 (N_17998,N_17312,N_17112);
nand U17999 (N_17999,N_17214,N_17385);
xnor U18000 (N_18000,N_17363,N_17416);
nand U18001 (N_18001,N_17447,N_17172);
or U18002 (N_18002,N_17364,N_17452);
or U18003 (N_18003,N_17005,N_17389);
or U18004 (N_18004,N_17449,N_17312);
or U18005 (N_18005,N_17091,N_17319);
or U18006 (N_18006,N_17048,N_17160);
or U18007 (N_18007,N_17278,N_17221);
and U18008 (N_18008,N_16930,N_16974);
or U18009 (N_18009,N_17478,N_17486);
nor U18010 (N_18010,N_17363,N_17065);
xnor U18011 (N_18011,N_17056,N_17497);
xnor U18012 (N_18012,N_17323,N_17450);
and U18013 (N_18013,N_17230,N_16908);
or U18014 (N_18014,N_16938,N_17121);
xor U18015 (N_18015,N_17039,N_17137);
nand U18016 (N_18016,N_17405,N_17112);
or U18017 (N_18017,N_17082,N_17496);
and U18018 (N_18018,N_17292,N_17376);
and U18019 (N_18019,N_17202,N_17269);
xnor U18020 (N_18020,N_17499,N_17329);
and U18021 (N_18021,N_17391,N_17012);
nand U18022 (N_18022,N_17298,N_16928);
nand U18023 (N_18023,N_17461,N_17394);
xnor U18024 (N_18024,N_17371,N_16999);
and U18025 (N_18025,N_16912,N_17074);
or U18026 (N_18026,N_16903,N_16985);
xor U18027 (N_18027,N_17271,N_17233);
nand U18028 (N_18028,N_17270,N_17295);
nand U18029 (N_18029,N_16972,N_17157);
nor U18030 (N_18030,N_17305,N_16936);
nor U18031 (N_18031,N_17173,N_17076);
nor U18032 (N_18032,N_16942,N_17342);
and U18033 (N_18033,N_17467,N_17403);
nand U18034 (N_18034,N_17322,N_16944);
or U18035 (N_18035,N_16954,N_16920);
nand U18036 (N_18036,N_17424,N_17113);
xnor U18037 (N_18037,N_17106,N_17024);
or U18038 (N_18038,N_17151,N_16975);
nand U18039 (N_18039,N_17356,N_17189);
or U18040 (N_18040,N_16983,N_17477);
xnor U18041 (N_18041,N_17004,N_16897);
or U18042 (N_18042,N_16910,N_17271);
nand U18043 (N_18043,N_16895,N_17328);
or U18044 (N_18044,N_17141,N_17310);
or U18045 (N_18045,N_17442,N_17139);
nor U18046 (N_18046,N_17364,N_16876);
nor U18047 (N_18047,N_16962,N_16886);
xnor U18048 (N_18048,N_17420,N_17470);
nand U18049 (N_18049,N_17214,N_16917);
nand U18050 (N_18050,N_17324,N_17052);
nand U18051 (N_18051,N_17366,N_17044);
nor U18052 (N_18052,N_17258,N_16947);
nand U18053 (N_18053,N_17204,N_17327);
nor U18054 (N_18054,N_17154,N_17271);
and U18055 (N_18055,N_16897,N_17321);
or U18056 (N_18056,N_17021,N_17178);
nor U18057 (N_18057,N_17220,N_17437);
nand U18058 (N_18058,N_17476,N_17160);
and U18059 (N_18059,N_17088,N_17047);
nor U18060 (N_18060,N_17059,N_17169);
nor U18061 (N_18061,N_17470,N_17150);
xnor U18062 (N_18062,N_17022,N_17469);
and U18063 (N_18063,N_17376,N_16897);
and U18064 (N_18064,N_16983,N_17121);
nor U18065 (N_18065,N_17085,N_17466);
or U18066 (N_18066,N_17377,N_16966);
nand U18067 (N_18067,N_16996,N_17082);
or U18068 (N_18068,N_16944,N_17486);
xnor U18069 (N_18069,N_17061,N_17028);
xnor U18070 (N_18070,N_17161,N_17183);
nand U18071 (N_18071,N_17252,N_17288);
xor U18072 (N_18072,N_17080,N_17383);
nand U18073 (N_18073,N_17168,N_17174);
and U18074 (N_18074,N_17317,N_17049);
nand U18075 (N_18075,N_17359,N_17444);
or U18076 (N_18076,N_16996,N_17379);
and U18077 (N_18077,N_17072,N_17099);
nor U18078 (N_18078,N_17140,N_17277);
nor U18079 (N_18079,N_17278,N_17204);
and U18080 (N_18080,N_16968,N_17408);
nor U18081 (N_18081,N_17328,N_17470);
nor U18082 (N_18082,N_17171,N_16994);
nand U18083 (N_18083,N_17200,N_17029);
nor U18084 (N_18084,N_17291,N_17212);
and U18085 (N_18085,N_17048,N_17391);
xnor U18086 (N_18086,N_17030,N_16996);
or U18087 (N_18087,N_17245,N_16979);
and U18088 (N_18088,N_16895,N_17353);
nor U18089 (N_18089,N_17321,N_17033);
nand U18090 (N_18090,N_17439,N_17216);
xor U18091 (N_18091,N_17451,N_17212);
or U18092 (N_18092,N_17158,N_17409);
xor U18093 (N_18093,N_17248,N_17179);
nor U18094 (N_18094,N_17463,N_17036);
xor U18095 (N_18095,N_17235,N_17143);
nand U18096 (N_18096,N_17453,N_17343);
nand U18097 (N_18097,N_17072,N_17107);
nand U18098 (N_18098,N_16987,N_17303);
and U18099 (N_18099,N_17416,N_17146);
nor U18100 (N_18100,N_17277,N_17243);
xnor U18101 (N_18101,N_17205,N_17481);
nor U18102 (N_18102,N_16891,N_17335);
xor U18103 (N_18103,N_17413,N_16938);
xnor U18104 (N_18104,N_17093,N_17237);
nor U18105 (N_18105,N_17402,N_16890);
xnor U18106 (N_18106,N_17481,N_16958);
and U18107 (N_18107,N_16980,N_16947);
and U18108 (N_18108,N_17326,N_17392);
or U18109 (N_18109,N_17292,N_16927);
nand U18110 (N_18110,N_17424,N_17120);
nand U18111 (N_18111,N_16897,N_16987);
and U18112 (N_18112,N_17157,N_17254);
nand U18113 (N_18113,N_17107,N_17181);
nand U18114 (N_18114,N_17204,N_17388);
nand U18115 (N_18115,N_16995,N_16925);
nor U18116 (N_18116,N_17033,N_16970);
xnor U18117 (N_18117,N_16977,N_17444);
nand U18118 (N_18118,N_17437,N_16919);
or U18119 (N_18119,N_17135,N_17309);
or U18120 (N_18120,N_17223,N_16966);
nand U18121 (N_18121,N_17184,N_17423);
nor U18122 (N_18122,N_17269,N_17432);
nor U18123 (N_18123,N_16939,N_17127);
xnor U18124 (N_18124,N_17295,N_17328);
and U18125 (N_18125,N_18089,N_17956);
or U18126 (N_18126,N_17950,N_17713);
or U18127 (N_18127,N_17906,N_17552);
nor U18128 (N_18128,N_17776,N_18120);
and U18129 (N_18129,N_17784,N_17993);
nand U18130 (N_18130,N_17888,N_17883);
and U18131 (N_18131,N_17611,N_17971);
and U18132 (N_18132,N_18098,N_17852);
nand U18133 (N_18133,N_17685,N_18039);
or U18134 (N_18134,N_17551,N_18015);
nor U18135 (N_18135,N_17988,N_18105);
nand U18136 (N_18136,N_17810,N_17651);
or U18137 (N_18137,N_17840,N_17858);
or U18138 (N_18138,N_17924,N_17601);
and U18139 (N_18139,N_17597,N_17679);
or U18140 (N_18140,N_17815,N_17925);
and U18141 (N_18141,N_17905,N_17580);
nor U18142 (N_18142,N_17828,N_17579);
and U18143 (N_18143,N_17664,N_17959);
nand U18144 (N_18144,N_18114,N_17766);
xor U18145 (N_18145,N_18021,N_17943);
and U18146 (N_18146,N_17737,N_17812);
xor U18147 (N_18147,N_17500,N_17650);
xor U18148 (N_18148,N_17518,N_18005);
nor U18149 (N_18149,N_18095,N_17897);
nor U18150 (N_18150,N_17787,N_17548);
or U18151 (N_18151,N_17671,N_18123);
xor U18152 (N_18152,N_17504,N_18102);
nand U18153 (N_18153,N_17600,N_17907);
nor U18154 (N_18154,N_17822,N_17602);
nand U18155 (N_18155,N_17527,N_17770);
nand U18156 (N_18156,N_17657,N_17534);
nor U18157 (N_18157,N_18010,N_17649);
and U18158 (N_18158,N_17636,N_17797);
xnor U18159 (N_18159,N_17790,N_17989);
xor U18160 (N_18160,N_17873,N_17684);
xor U18161 (N_18161,N_17767,N_17529);
xnor U18162 (N_18162,N_17506,N_17798);
nand U18163 (N_18163,N_17744,N_18042);
nand U18164 (N_18164,N_17922,N_18020);
nor U18165 (N_18165,N_17522,N_17878);
or U18166 (N_18166,N_18079,N_17753);
and U18167 (N_18167,N_17505,N_17708);
or U18168 (N_18168,N_17808,N_17793);
or U18169 (N_18169,N_17992,N_17917);
nor U18170 (N_18170,N_17741,N_17544);
xnor U18171 (N_18171,N_17855,N_18029);
xor U18172 (N_18172,N_17947,N_18101);
nand U18173 (N_18173,N_17613,N_17738);
and U18174 (N_18174,N_17598,N_17550);
nor U18175 (N_18175,N_17641,N_18071);
nand U18176 (N_18176,N_17759,N_17707);
and U18177 (N_18177,N_18043,N_17977);
nor U18178 (N_18178,N_17789,N_17817);
xor U18179 (N_18179,N_17524,N_18117);
and U18180 (N_18180,N_17760,N_17903);
and U18181 (N_18181,N_17909,N_17990);
or U18182 (N_18182,N_17612,N_17694);
xor U18183 (N_18183,N_17614,N_17898);
or U18184 (N_18184,N_18003,N_17867);
xor U18185 (N_18185,N_17692,N_17618);
nor U18186 (N_18186,N_17582,N_17591);
nand U18187 (N_18187,N_17982,N_18053);
nor U18188 (N_18188,N_18004,N_17740);
nand U18189 (N_18189,N_17985,N_17837);
xnor U18190 (N_18190,N_17845,N_17691);
or U18191 (N_18191,N_17821,N_18007);
and U18192 (N_18192,N_17973,N_17607);
nand U18193 (N_18193,N_18121,N_17934);
or U18194 (N_18194,N_18001,N_17722);
xor U18195 (N_18195,N_17592,N_17997);
and U18196 (N_18196,N_17951,N_18055);
and U18197 (N_18197,N_17663,N_17652);
nand U18198 (N_18198,N_17718,N_17512);
xor U18199 (N_18199,N_17751,N_18023);
and U18200 (N_18200,N_18027,N_17964);
nor U18201 (N_18201,N_17944,N_17528);
nand U18202 (N_18202,N_17764,N_17953);
and U18203 (N_18203,N_17577,N_17929);
xnor U18204 (N_18204,N_17847,N_18031);
nor U18205 (N_18205,N_17732,N_17520);
xor U18206 (N_18206,N_18110,N_18017);
or U18207 (N_18207,N_17996,N_17511);
and U18208 (N_18208,N_17761,N_17616);
nand U18209 (N_18209,N_17714,N_17891);
nor U18210 (N_18210,N_17555,N_18062);
xor U18211 (N_18211,N_18111,N_17653);
nand U18212 (N_18212,N_18035,N_17674);
and U18213 (N_18213,N_17879,N_17886);
or U18214 (N_18214,N_18049,N_17742);
xor U18215 (N_18215,N_17892,N_17687);
xor U18216 (N_18216,N_17806,N_17557);
nand U18217 (N_18217,N_17573,N_17863);
xnor U18218 (N_18218,N_17615,N_17622);
nor U18219 (N_18219,N_18124,N_17626);
or U18220 (N_18220,N_18002,N_17771);
and U18221 (N_18221,N_17517,N_17726);
nand U18222 (N_18222,N_18030,N_18032);
nand U18223 (N_18223,N_17583,N_18006);
nand U18224 (N_18224,N_17609,N_17778);
nand U18225 (N_18225,N_18060,N_18013);
nand U18226 (N_18226,N_17834,N_18107);
xnor U18227 (N_18227,N_18091,N_17836);
or U18228 (N_18228,N_17927,N_17594);
and U18229 (N_18229,N_17590,N_17918);
nor U18230 (N_18230,N_17632,N_17937);
and U18231 (N_18231,N_17794,N_18066);
nand U18232 (N_18232,N_17763,N_17525);
nor U18233 (N_18233,N_17667,N_18059);
nor U18234 (N_18234,N_17814,N_17786);
nor U18235 (N_18235,N_17772,N_17725);
nand U18236 (N_18236,N_17755,N_17606);
or U18237 (N_18237,N_17887,N_17781);
nor U18238 (N_18238,N_17588,N_17890);
nand U18239 (N_18239,N_17757,N_18088);
and U18240 (N_18240,N_17541,N_17853);
nor U18241 (N_18241,N_18051,N_17746);
nor U18242 (N_18242,N_17670,N_17800);
nand U18243 (N_18243,N_17859,N_17716);
nor U18244 (N_18244,N_17889,N_17818);
xnor U18245 (N_18245,N_17710,N_18008);
or U18246 (N_18246,N_17928,N_17975);
nor U18247 (N_18247,N_17948,N_17914);
and U18248 (N_18248,N_17962,N_17659);
nor U18249 (N_18249,N_17904,N_17532);
xnor U18250 (N_18250,N_17709,N_17967);
nand U18251 (N_18251,N_18054,N_17578);
or U18252 (N_18252,N_18026,N_17645);
and U18253 (N_18253,N_17874,N_18108);
and U18254 (N_18254,N_17570,N_18009);
or U18255 (N_18255,N_18058,N_17976);
nand U18256 (N_18256,N_17830,N_17549);
or U18257 (N_18257,N_18064,N_18093);
xnor U18258 (N_18258,N_17644,N_17969);
nor U18259 (N_18259,N_17823,N_17819);
and U18260 (N_18260,N_18085,N_17980);
xnor U18261 (N_18261,N_17727,N_18068);
and U18262 (N_18262,N_17567,N_17768);
nor U18263 (N_18263,N_17523,N_17593);
and U18264 (N_18264,N_17756,N_18073);
nor U18265 (N_18265,N_17515,N_17884);
and U18266 (N_18266,N_17688,N_17734);
nand U18267 (N_18267,N_17783,N_17595);
nand U18268 (N_18268,N_17563,N_17900);
or U18269 (N_18269,N_17862,N_17844);
nor U18270 (N_18270,N_18113,N_17882);
nand U18271 (N_18271,N_17605,N_17695);
and U18272 (N_18272,N_17829,N_17516);
and U18273 (N_18273,N_17963,N_17940);
or U18274 (N_18274,N_18080,N_17938);
nand U18275 (N_18275,N_17868,N_17748);
nand U18276 (N_18276,N_17676,N_17678);
or U18277 (N_18277,N_17665,N_17805);
nor U18278 (N_18278,N_17639,N_17728);
xnor U18279 (N_18279,N_17585,N_17655);
and U18280 (N_18280,N_17696,N_17777);
nor U18281 (N_18281,N_18099,N_18046);
and U18282 (N_18282,N_17720,N_17824);
nor U18283 (N_18283,N_17724,N_17958);
nand U18284 (N_18284,N_17832,N_17954);
nor U18285 (N_18285,N_17546,N_17893);
nor U18286 (N_18286,N_17865,N_17625);
and U18287 (N_18287,N_17683,N_17677);
and U18288 (N_18288,N_17635,N_18103);
nand U18289 (N_18289,N_17535,N_17536);
nand U18290 (N_18290,N_17885,N_17656);
or U18291 (N_18291,N_17876,N_17881);
or U18292 (N_18292,N_17995,N_17672);
nand U18293 (N_18293,N_17843,N_18104);
nand U18294 (N_18294,N_18045,N_18096);
xor U18295 (N_18295,N_17902,N_17848);
and U18296 (N_18296,N_18022,N_18116);
nand U18297 (N_18297,N_17796,N_17589);
nand U18298 (N_18298,N_17745,N_17991);
nor U18299 (N_18299,N_17507,N_17825);
nand U18300 (N_18300,N_17508,N_17599);
nand U18301 (N_18301,N_18052,N_17773);
and U18302 (N_18302,N_17941,N_17935);
xor U18303 (N_18303,N_17701,N_18014);
or U18304 (N_18304,N_17712,N_17983);
or U18305 (N_18305,N_17831,N_17556);
nand U18306 (N_18306,N_17634,N_17895);
xor U18307 (N_18307,N_17752,N_17526);
and U18308 (N_18308,N_18000,N_17946);
and U18309 (N_18309,N_17542,N_17920);
xor U18310 (N_18310,N_17801,N_17921);
nor U18311 (N_18311,N_18112,N_17566);
xnor U18312 (N_18312,N_17539,N_17561);
or U18313 (N_18313,N_17916,N_17621);
nand U18314 (N_18314,N_17804,N_17503);
xor U18315 (N_18315,N_17637,N_17608);
nor U18316 (N_18316,N_17700,N_17610);
or U18317 (N_18317,N_17877,N_17735);
xnor U18318 (N_18318,N_17864,N_17519);
nand U18319 (N_18319,N_18050,N_17998);
nor U18320 (N_18320,N_17627,N_17559);
nor U18321 (N_18321,N_18028,N_17623);
and U18322 (N_18322,N_17970,N_17681);
xor U18323 (N_18323,N_18033,N_18092);
xor U18324 (N_18324,N_17620,N_17624);
and U18325 (N_18325,N_17564,N_18038);
and U18326 (N_18326,N_17514,N_18081);
nand U18327 (N_18327,N_17533,N_17849);
or U18328 (N_18328,N_18044,N_17658);
and U18329 (N_18329,N_17870,N_18072);
nor U18330 (N_18330,N_17638,N_18087);
and U18331 (N_18331,N_17788,N_17510);
or U18332 (N_18332,N_17699,N_17972);
nor U18333 (N_18333,N_17999,N_17587);
and U18334 (N_18334,N_18047,N_17913);
nand U18335 (N_18335,N_17565,N_17568);
nand U18336 (N_18336,N_18075,N_17880);
or U18337 (N_18337,N_17690,N_17723);
or U18338 (N_18338,N_17986,N_17939);
or U18339 (N_18339,N_17711,N_17662);
or U18340 (N_18340,N_18100,N_17680);
or U18341 (N_18341,N_17633,N_17571);
and U18342 (N_18342,N_17617,N_17811);
and U18343 (N_18343,N_17799,N_17509);
or U18344 (N_18344,N_17926,N_17730);
and U18345 (N_18345,N_17697,N_17747);
or U18346 (N_18346,N_17803,N_18036);
xor U18347 (N_18347,N_17931,N_17932);
or U18348 (N_18348,N_17553,N_17743);
nor U18349 (N_18349,N_17540,N_17547);
and U18350 (N_18350,N_17543,N_17693);
nand U18351 (N_18351,N_17974,N_17596);
and U18352 (N_18352,N_18037,N_17576);
or U18353 (N_18353,N_17762,N_17705);
xor U18354 (N_18354,N_17899,N_18019);
xnor U18355 (N_18355,N_17846,N_17686);
nor U18356 (N_18356,N_17558,N_17733);
xnor U18357 (N_18357,N_17660,N_17850);
or U18358 (N_18358,N_17936,N_17765);
or U18359 (N_18359,N_17802,N_17966);
xor U18360 (N_18360,N_17758,N_17682);
or U18361 (N_18361,N_17739,N_18082);
xor U18362 (N_18362,N_17961,N_17908);
and U18363 (N_18363,N_18024,N_18057);
nand U18364 (N_18364,N_18118,N_17955);
xor U18365 (N_18365,N_18070,N_18122);
and U18366 (N_18366,N_17875,N_17668);
and U18367 (N_18367,N_17957,N_17640);
and U18368 (N_18368,N_17630,N_17872);
or U18369 (N_18369,N_17643,N_18106);
xor U18370 (N_18370,N_17642,N_18109);
nand U18371 (N_18371,N_17704,N_18012);
xor U18372 (N_18372,N_17648,N_18065);
xnor U18373 (N_18373,N_17866,N_17978);
nand U18374 (N_18374,N_17675,N_18119);
nor U18375 (N_18375,N_17912,N_17820);
or U18376 (N_18376,N_17979,N_17513);
or U18377 (N_18377,N_17545,N_18011);
and U18378 (N_18378,N_18067,N_17839);
xnor U18379 (N_18379,N_18090,N_17689);
and U18380 (N_18380,N_17581,N_17715);
and U18381 (N_18381,N_17749,N_18040);
and U18382 (N_18382,N_18069,N_17827);
or U18383 (N_18383,N_18078,N_18034);
nand U18384 (N_18384,N_17554,N_17833);
nor U18385 (N_18385,N_17856,N_17968);
and U18386 (N_18386,N_17574,N_17901);
nor U18387 (N_18387,N_17666,N_17619);
nand U18388 (N_18388,N_17861,N_17719);
and U18389 (N_18389,N_17569,N_18084);
nand U18390 (N_18390,N_17942,N_17792);
nand U18391 (N_18391,N_18074,N_17807);
xor U18392 (N_18392,N_17629,N_17702);
and U18393 (N_18393,N_17562,N_17706);
nand U18394 (N_18394,N_17838,N_17949);
nand U18395 (N_18395,N_17560,N_17530);
or U18396 (N_18396,N_17631,N_17857);
xnor U18397 (N_18397,N_17721,N_18076);
xor U18398 (N_18398,N_17894,N_17911);
nand U18399 (N_18399,N_17919,N_17994);
nor U18400 (N_18400,N_17782,N_17775);
nand U18401 (N_18401,N_17779,N_18061);
nor U18402 (N_18402,N_17731,N_17628);
nor U18403 (N_18403,N_17930,N_17603);
xor U18404 (N_18404,N_17869,N_17816);
nand U18405 (N_18405,N_18077,N_17646);
nor U18406 (N_18406,N_18094,N_17960);
nand U18407 (N_18407,N_17896,N_17502);
or U18408 (N_18408,N_17785,N_18086);
or U18409 (N_18409,N_17791,N_17521);
and U18410 (N_18410,N_18048,N_17729);
and U18411 (N_18411,N_18063,N_17860);
nand U18412 (N_18412,N_17537,N_18018);
or U18413 (N_18413,N_17736,N_17584);
or U18414 (N_18414,N_17809,N_18016);
xnor U18415 (N_18415,N_17769,N_17754);
nor U18416 (N_18416,N_18115,N_17842);
nand U18417 (N_18417,N_17915,N_18083);
nand U18418 (N_18418,N_17774,N_17572);
and U18419 (N_18419,N_17780,N_17945);
nor U18420 (N_18420,N_18041,N_17717);
and U18421 (N_18421,N_17871,N_17661);
nand U18422 (N_18422,N_17835,N_17854);
xor U18423 (N_18423,N_17586,N_17952);
nand U18424 (N_18424,N_17669,N_17841);
or U18425 (N_18425,N_17703,N_17933);
nor U18426 (N_18426,N_17987,N_17981);
or U18427 (N_18427,N_17851,N_17910);
and U18428 (N_18428,N_17647,N_17826);
xnor U18429 (N_18429,N_17531,N_18056);
and U18430 (N_18430,N_17750,N_18097);
or U18431 (N_18431,N_17795,N_17813);
nand U18432 (N_18432,N_18025,N_17501);
nand U18433 (N_18433,N_17673,N_17984);
and U18434 (N_18434,N_17538,N_17575);
nor U18435 (N_18435,N_17965,N_17654);
and U18436 (N_18436,N_17698,N_17923);
nor U18437 (N_18437,N_17604,N_17844);
nor U18438 (N_18438,N_17640,N_17584);
xor U18439 (N_18439,N_17673,N_17848);
nand U18440 (N_18440,N_17501,N_17507);
nand U18441 (N_18441,N_17976,N_17964);
or U18442 (N_18442,N_17925,N_17856);
or U18443 (N_18443,N_18092,N_18115);
nand U18444 (N_18444,N_17879,N_17807);
nand U18445 (N_18445,N_17504,N_17709);
nand U18446 (N_18446,N_17632,N_17817);
xor U18447 (N_18447,N_17688,N_18023);
xnor U18448 (N_18448,N_17580,N_17668);
nand U18449 (N_18449,N_17790,N_17873);
and U18450 (N_18450,N_17511,N_17748);
or U18451 (N_18451,N_18055,N_17641);
nand U18452 (N_18452,N_17999,N_17691);
nor U18453 (N_18453,N_17771,N_17821);
nor U18454 (N_18454,N_17701,N_17621);
nand U18455 (N_18455,N_17729,N_17787);
and U18456 (N_18456,N_17765,N_17887);
xor U18457 (N_18457,N_17765,N_17667);
xor U18458 (N_18458,N_17569,N_17541);
nor U18459 (N_18459,N_17808,N_17751);
nand U18460 (N_18460,N_17987,N_17632);
or U18461 (N_18461,N_17733,N_18072);
nand U18462 (N_18462,N_17797,N_17716);
nor U18463 (N_18463,N_17563,N_18104);
and U18464 (N_18464,N_17880,N_17994);
or U18465 (N_18465,N_18021,N_17745);
or U18466 (N_18466,N_17851,N_17899);
nor U18467 (N_18467,N_18060,N_18053);
nor U18468 (N_18468,N_18031,N_18014);
nand U18469 (N_18469,N_17892,N_18058);
and U18470 (N_18470,N_17927,N_17545);
nor U18471 (N_18471,N_17533,N_18099);
xnor U18472 (N_18472,N_17547,N_17890);
and U18473 (N_18473,N_17696,N_17919);
nand U18474 (N_18474,N_18006,N_17538);
xor U18475 (N_18475,N_17517,N_17584);
and U18476 (N_18476,N_17602,N_17925);
or U18477 (N_18477,N_17920,N_17968);
xnor U18478 (N_18478,N_18082,N_17747);
or U18479 (N_18479,N_17773,N_18063);
or U18480 (N_18480,N_17815,N_17783);
and U18481 (N_18481,N_18009,N_17502);
nand U18482 (N_18482,N_17535,N_17645);
or U18483 (N_18483,N_17623,N_18023);
or U18484 (N_18484,N_17764,N_17597);
and U18485 (N_18485,N_18092,N_17606);
nor U18486 (N_18486,N_17757,N_18073);
nand U18487 (N_18487,N_17501,N_17946);
or U18488 (N_18488,N_17677,N_17964);
or U18489 (N_18489,N_18022,N_17905);
or U18490 (N_18490,N_17686,N_17886);
or U18491 (N_18491,N_17737,N_17746);
xor U18492 (N_18492,N_17599,N_17675);
or U18493 (N_18493,N_17807,N_17731);
and U18494 (N_18494,N_17768,N_18083);
xnor U18495 (N_18495,N_17642,N_17559);
xor U18496 (N_18496,N_18074,N_17518);
nor U18497 (N_18497,N_17919,N_17704);
or U18498 (N_18498,N_17821,N_18043);
or U18499 (N_18499,N_17588,N_17649);
nor U18500 (N_18500,N_17585,N_17617);
nand U18501 (N_18501,N_18028,N_17821);
nor U18502 (N_18502,N_17537,N_17645);
nand U18503 (N_18503,N_17788,N_18087);
xor U18504 (N_18504,N_17988,N_17760);
nor U18505 (N_18505,N_17564,N_17533);
xnor U18506 (N_18506,N_17600,N_17795);
and U18507 (N_18507,N_17987,N_18079);
nand U18508 (N_18508,N_17876,N_18026);
nand U18509 (N_18509,N_17573,N_17968);
nand U18510 (N_18510,N_17789,N_17894);
and U18511 (N_18511,N_17540,N_17910);
and U18512 (N_18512,N_18045,N_17888);
and U18513 (N_18513,N_17721,N_18121);
and U18514 (N_18514,N_17731,N_17653);
and U18515 (N_18515,N_17998,N_17976);
nand U18516 (N_18516,N_17511,N_17881);
or U18517 (N_18517,N_17636,N_17562);
or U18518 (N_18518,N_17801,N_17689);
and U18519 (N_18519,N_17797,N_18001);
and U18520 (N_18520,N_18083,N_18123);
nor U18521 (N_18521,N_18001,N_17768);
nand U18522 (N_18522,N_17549,N_17727);
and U18523 (N_18523,N_18104,N_17604);
or U18524 (N_18524,N_17710,N_17580);
nor U18525 (N_18525,N_18046,N_17532);
or U18526 (N_18526,N_18085,N_17872);
nor U18527 (N_18527,N_17807,N_17752);
xor U18528 (N_18528,N_17916,N_17818);
and U18529 (N_18529,N_17734,N_17923);
nor U18530 (N_18530,N_17565,N_17508);
or U18531 (N_18531,N_18038,N_18067);
nand U18532 (N_18532,N_17851,N_17962);
nand U18533 (N_18533,N_17728,N_18059);
nand U18534 (N_18534,N_17820,N_17587);
or U18535 (N_18535,N_17993,N_17749);
nor U18536 (N_18536,N_17525,N_18074);
nand U18537 (N_18537,N_17734,N_17547);
or U18538 (N_18538,N_18044,N_17763);
xor U18539 (N_18539,N_17943,N_17989);
nor U18540 (N_18540,N_17551,N_17547);
nand U18541 (N_18541,N_17638,N_17964);
nand U18542 (N_18542,N_17586,N_18118);
xnor U18543 (N_18543,N_17624,N_18077);
or U18544 (N_18544,N_17610,N_17628);
nand U18545 (N_18545,N_17559,N_17847);
or U18546 (N_18546,N_17778,N_18096);
nor U18547 (N_18547,N_17962,N_17663);
or U18548 (N_18548,N_18023,N_17821);
or U18549 (N_18549,N_18120,N_18032);
nand U18550 (N_18550,N_17513,N_17686);
and U18551 (N_18551,N_17760,N_17643);
and U18552 (N_18552,N_17608,N_18017);
nor U18553 (N_18553,N_17896,N_17618);
xor U18554 (N_18554,N_18021,N_18029);
nor U18555 (N_18555,N_17641,N_17896);
nor U18556 (N_18556,N_18013,N_18046);
nor U18557 (N_18557,N_17822,N_17577);
nand U18558 (N_18558,N_17848,N_17890);
or U18559 (N_18559,N_17973,N_17773);
xor U18560 (N_18560,N_17530,N_17650);
and U18561 (N_18561,N_17814,N_17778);
or U18562 (N_18562,N_17922,N_17823);
xnor U18563 (N_18563,N_18006,N_17751);
and U18564 (N_18564,N_17653,N_18109);
nand U18565 (N_18565,N_18039,N_17523);
and U18566 (N_18566,N_18107,N_17861);
xnor U18567 (N_18567,N_17893,N_17891);
or U18568 (N_18568,N_18124,N_17562);
nor U18569 (N_18569,N_17537,N_17843);
or U18570 (N_18570,N_18003,N_17996);
or U18571 (N_18571,N_17511,N_17841);
xor U18572 (N_18572,N_17723,N_17925);
nor U18573 (N_18573,N_18022,N_17780);
nor U18574 (N_18574,N_18026,N_17533);
nand U18575 (N_18575,N_17519,N_17725);
xor U18576 (N_18576,N_17673,N_17910);
and U18577 (N_18577,N_17675,N_17988);
or U18578 (N_18578,N_17893,N_18022);
xnor U18579 (N_18579,N_17567,N_17837);
nor U18580 (N_18580,N_17716,N_17688);
nand U18581 (N_18581,N_18075,N_17805);
xnor U18582 (N_18582,N_17570,N_18074);
xor U18583 (N_18583,N_17819,N_17883);
nor U18584 (N_18584,N_17714,N_17828);
or U18585 (N_18585,N_17723,N_17764);
nor U18586 (N_18586,N_18022,N_17730);
nand U18587 (N_18587,N_17797,N_17922);
xor U18588 (N_18588,N_17731,N_17880);
xor U18589 (N_18589,N_17840,N_18035);
nor U18590 (N_18590,N_17978,N_18040);
nor U18591 (N_18591,N_17542,N_17862);
xnor U18592 (N_18592,N_17587,N_17540);
and U18593 (N_18593,N_17533,N_17882);
and U18594 (N_18594,N_17871,N_18067);
nand U18595 (N_18595,N_17851,N_17985);
xnor U18596 (N_18596,N_18065,N_17561);
or U18597 (N_18597,N_17606,N_17916);
nor U18598 (N_18598,N_18082,N_17980);
nor U18599 (N_18599,N_17896,N_17809);
and U18600 (N_18600,N_17882,N_17923);
nand U18601 (N_18601,N_17845,N_18019);
or U18602 (N_18602,N_17503,N_17929);
or U18603 (N_18603,N_17931,N_18032);
or U18604 (N_18604,N_17714,N_18046);
and U18605 (N_18605,N_18090,N_18061);
or U18606 (N_18606,N_17608,N_17991);
and U18607 (N_18607,N_17937,N_18078);
nand U18608 (N_18608,N_18085,N_17982);
or U18609 (N_18609,N_18036,N_18030);
xnor U18610 (N_18610,N_17514,N_17891);
nand U18611 (N_18611,N_17553,N_17920);
or U18612 (N_18612,N_17744,N_17855);
nand U18613 (N_18613,N_17588,N_17762);
nor U18614 (N_18614,N_17604,N_18091);
nand U18615 (N_18615,N_17826,N_17671);
nand U18616 (N_18616,N_17910,N_17517);
nor U18617 (N_18617,N_18048,N_17930);
nor U18618 (N_18618,N_17533,N_17877);
or U18619 (N_18619,N_17747,N_17864);
nor U18620 (N_18620,N_18071,N_18085);
and U18621 (N_18621,N_17586,N_18104);
xor U18622 (N_18622,N_18029,N_17652);
and U18623 (N_18623,N_17730,N_17618);
nand U18624 (N_18624,N_17984,N_17603);
nand U18625 (N_18625,N_17501,N_17614);
nand U18626 (N_18626,N_17644,N_17925);
nand U18627 (N_18627,N_17581,N_17985);
nor U18628 (N_18628,N_17679,N_17757);
and U18629 (N_18629,N_17591,N_17995);
and U18630 (N_18630,N_17871,N_17663);
nor U18631 (N_18631,N_17593,N_17874);
nand U18632 (N_18632,N_17660,N_17769);
nand U18633 (N_18633,N_18091,N_17830);
xor U18634 (N_18634,N_17509,N_18063);
nor U18635 (N_18635,N_18092,N_18112);
or U18636 (N_18636,N_17641,N_18089);
nand U18637 (N_18637,N_17529,N_18113);
nor U18638 (N_18638,N_17688,N_17998);
nand U18639 (N_18639,N_18117,N_18037);
xor U18640 (N_18640,N_17915,N_18001);
or U18641 (N_18641,N_17859,N_17684);
nor U18642 (N_18642,N_18100,N_17522);
nor U18643 (N_18643,N_17636,N_17710);
or U18644 (N_18644,N_17851,N_18048);
or U18645 (N_18645,N_17632,N_17749);
and U18646 (N_18646,N_17568,N_17542);
nor U18647 (N_18647,N_17723,N_17627);
nor U18648 (N_18648,N_17547,N_17818);
and U18649 (N_18649,N_17839,N_18056);
and U18650 (N_18650,N_18053,N_17657);
and U18651 (N_18651,N_17566,N_17791);
nor U18652 (N_18652,N_17947,N_17523);
nand U18653 (N_18653,N_17848,N_17988);
and U18654 (N_18654,N_17842,N_17815);
or U18655 (N_18655,N_17680,N_17772);
xnor U18656 (N_18656,N_18068,N_18070);
nand U18657 (N_18657,N_17633,N_17695);
xor U18658 (N_18658,N_18011,N_17875);
nand U18659 (N_18659,N_17910,N_17511);
nand U18660 (N_18660,N_18084,N_18091);
nor U18661 (N_18661,N_17680,N_17641);
and U18662 (N_18662,N_17748,N_17603);
and U18663 (N_18663,N_17713,N_17848);
nand U18664 (N_18664,N_18098,N_18009);
or U18665 (N_18665,N_17821,N_17672);
nor U18666 (N_18666,N_17819,N_17660);
or U18667 (N_18667,N_17750,N_17697);
or U18668 (N_18668,N_17519,N_17796);
nand U18669 (N_18669,N_18117,N_18085);
and U18670 (N_18670,N_17931,N_17594);
nor U18671 (N_18671,N_18053,N_17745);
nor U18672 (N_18672,N_17722,N_17816);
and U18673 (N_18673,N_17974,N_17875);
nor U18674 (N_18674,N_17698,N_17983);
xor U18675 (N_18675,N_18038,N_17955);
xnor U18676 (N_18676,N_17889,N_17991);
and U18677 (N_18677,N_17681,N_17930);
nand U18678 (N_18678,N_18095,N_17719);
nand U18679 (N_18679,N_17558,N_17729);
xor U18680 (N_18680,N_17591,N_17993);
nand U18681 (N_18681,N_17669,N_17695);
or U18682 (N_18682,N_17807,N_17798);
nand U18683 (N_18683,N_17849,N_18063);
or U18684 (N_18684,N_18117,N_17920);
nor U18685 (N_18685,N_18076,N_17761);
nand U18686 (N_18686,N_18071,N_17797);
or U18687 (N_18687,N_17744,N_17952);
and U18688 (N_18688,N_17772,N_18075);
or U18689 (N_18689,N_18084,N_18008);
nor U18690 (N_18690,N_17596,N_17606);
nand U18691 (N_18691,N_17861,N_18100);
xor U18692 (N_18692,N_18011,N_17812);
xnor U18693 (N_18693,N_17517,N_17625);
and U18694 (N_18694,N_17868,N_17558);
xor U18695 (N_18695,N_18026,N_17557);
nand U18696 (N_18696,N_17545,N_17729);
and U18697 (N_18697,N_18068,N_18016);
or U18698 (N_18698,N_17936,N_17701);
and U18699 (N_18699,N_17716,N_17535);
or U18700 (N_18700,N_17645,N_17520);
nand U18701 (N_18701,N_17573,N_17881);
nand U18702 (N_18702,N_17765,N_17656);
or U18703 (N_18703,N_17604,N_17537);
xnor U18704 (N_18704,N_17542,N_18000);
and U18705 (N_18705,N_17566,N_17841);
or U18706 (N_18706,N_17641,N_17903);
xnor U18707 (N_18707,N_17662,N_17823);
xor U18708 (N_18708,N_17846,N_17842);
nand U18709 (N_18709,N_17619,N_17873);
xor U18710 (N_18710,N_18092,N_17886);
or U18711 (N_18711,N_17812,N_17932);
nand U18712 (N_18712,N_18057,N_17907);
nor U18713 (N_18713,N_17945,N_17841);
nand U18714 (N_18714,N_18074,N_17587);
nor U18715 (N_18715,N_17851,N_17675);
xor U18716 (N_18716,N_17636,N_17748);
and U18717 (N_18717,N_17632,N_18036);
nand U18718 (N_18718,N_17877,N_18031);
xnor U18719 (N_18719,N_18096,N_17577);
and U18720 (N_18720,N_17959,N_17572);
and U18721 (N_18721,N_18040,N_17887);
and U18722 (N_18722,N_17783,N_17891);
nor U18723 (N_18723,N_17627,N_17996);
and U18724 (N_18724,N_17812,N_18100);
nand U18725 (N_18725,N_18121,N_17859);
nand U18726 (N_18726,N_17904,N_17853);
nor U18727 (N_18727,N_18068,N_17546);
nor U18728 (N_18728,N_17568,N_18050);
or U18729 (N_18729,N_17598,N_17526);
xor U18730 (N_18730,N_17769,N_18023);
or U18731 (N_18731,N_17940,N_17987);
xnor U18732 (N_18732,N_17828,N_17573);
or U18733 (N_18733,N_17658,N_17627);
and U18734 (N_18734,N_18082,N_17986);
or U18735 (N_18735,N_18050,N_17508);
and U18736 (N_18736,N_17697,N_18053);
xnor U18737 (N_18737,N_17686,N_17877);
nor U18738 (N_18738,N_17868,N_17816);
nor U18739 (N_18739,N_17731,N_17550);
nor U18740 (N_18740,N_17964,N_17948);
and U18741 (N_18741,N_17521,N_18027);
xnor U18742 (N_18742,N_17575,N_18002);
nor U18743 (N_18743,N_17877,N_17714);
or U18744 (N_18744,N_17582,N_17620);
and U18745 (N_18745,N_17943,N_17627);
and U18746 (N_18746,N_17564,N_18055);
and U18747 (N_18747,N_18003,N_17880);
xor U18748 (N_18748,N_17596,N_17589);
and U18749 (N_18749,N_18050,N_17852);
nand U18750 (N_18750,N_18694,N_18465);
or U18751 (N_18751,N_18512,N_18641);
and U18752 (N_18752,N_18405,N_18546);
nor U18753 (N_18753,N_18608,N_18436);
nand U18754 (N_18754,N_18262,N_18470);
nand U18755 (N_18755,N_18565,N_18586);
xor U18756 (N_18756,N_18476,N_18592);
or U18757 (N_18757,N_18369,N_18496);
xnor U18758 (N_18758,N_18399,N_18441);
nand U18759 (N_18759,N_18708,N_18202);
and U18760 (N_18760,N_18269,N_18386);
xnor U18761 (N_18761,N_18668,N_18696);
nor U18762 (N_18762,N_18205,N_18324);
nand U18763 (N_18763,N_18398,N_18401);
and U18764 (N_18764,N_18515,N_18477);
nor U18765 (N_18765,N_18161,N_18204);
and U18766 (N_18766,N_18139,N_18278);
nand U18767 (N_18767,N_18435,N_18687);
and U18768 (N_18768,N_18638,N_18260);
and U18769 (N_18769,N_18553,N_18360);
nand U18770 (N_18770,N_18737,N_18368);
and U18771 (N_18771,N_18646,N_18390);
xor U18772 (N_18772,N_18140,N_18653);
or U18773 (N_18773,N_18388,N_18573);
nand U18774 (N_18774,N_18662,N_18245);
nand U18775 (N_18775,N_18525,N_18303);
nor U18776 (N_18776,N_18527,N_18718);
xor U18777 (N_18777,N_18517,N_18666);
nand U18778 (N_18778,N_18232,N_18634);
and U18779 (N_18779,N_18376,N_18611);
xnor U18780 (N_18780,N_18313,N_18615);
and U18781 (N_18781,N_18463,N_18178);
nand U18782 (N_18782,N_18621,N_18670);
and U18783 (N_18783,N_18287,N_18373);
nand U18784 (N_18784,N_18133,N_18511);
nor U18785 (N_18785,N_18551,N_18251);
xnor U18786 (N_18786,N_18567,N_18366);
nand U18787 (N_18787,N_18200,N_18295);
nor U18788 (N_18788,N_18524,N_18654);
xor U18789 (N_18789,N_18167,N_18280);
nor U18790 (N_18790,N_18539,N_18258);
or U18791 (N_18791,N_18695,N_18259);
and U18792 (N_18792,N_18354,N_18307);
and U18793 (N_18793,N_18682,N_18249);
nand U18794 (N_18794,N_18176,N_18520);
or U18795 (N_18795,N_18271,N_18219);
and U18796 (N_18796,N_18595,N_18177);
nand U18797 (N_18797,N_18603,N_18721);
nand U18798 (N_18798,N_18510,N_18692);
or U18799 (N_18799,N_18424,N_18207);
nor U18800 (N_18800,N_18327,N_18183);
nand U18801 (N_18801,N_18344,N_18558);
nor U18802 (N_18802,N_18227,N_18648);
and U18803 (N_18803,N_18663,N_18628);
nand U18804 (N_18804,N_18364,N_18206);
or U18805 (N_18805,N_18691,N_18469);
xor U18806 (N_18806,N_18690,N_18328);
and U18807 (N_18807,N_18652,N_18700);
or U18808 (N_18808,N_18371,N_18671);
and U18809 (N_18809,N_18361,N_18238);
and U18810 (N_18810,N_18452,N_18711);
and U18811 (N_18811,N_18316,N_18148);
nor U18812 (N_18812,N_18735,N_18460);
nand U18813 (N_18813,N_18334,N_18554);
xnor U18814 (N_18814,N_18739,N_18385);
or U18815 (N_18815,N_18427,N_18677);
xnor U18816 (N_18816,N_18490,N_18623);
xor U18817 (N_18817,N_18560,N_18555);
nand U18818 (N_18818,N_18577,N_18459);
xor U18819 (N_18819,N_18346,N_18365);
xnor U18820 (N_18820,N_18732,N_18387);
or U18821 (N_18821,N_18297,N_18283);
nand U18822 (N_18822,N_18449,N_18636);
nor U18823 (N_18823,N_18162,N_18188);
nor U18824 (N_18824,N_18584,N_18717);
nor U18825 (N_18825,N_18409,N_18741);
nor U18826 (N_18826,N_18518,N_18175);
nor U18827 (N_18827,N_18285,N_18521);
nand U18828 (N_18828,N_18263,N_18506);
nand U18829 (N_18829,N_18571,N_18343);
xor U18830 (N_18830,N_18348,N_18442);
nor U18831 (N_18831,N_18288,N_18645);
or U18832 (N_18832,N_18186,N_18617);
or U18833 (N_18833,N_18362,N_18400);
nor U18834 (N_18834,N_18557,N_18268);
and U18835 (N_18835,N_18302,N_18314);
nor U18836 (N_18836,N_18282,N_18128);
nand U18837 (N_18837,N_18256,N_18208);
nor U18838 (N_18838,N_18604,N_18247);
nand U18839 (N_18839,N_18193,N_18154);
and U18840 (N_18840,N_18438,N_18516);
xnor U18841 (N_18841,N_18315,N_18531);
xnor U18842 (N_18842,N_18533,N_18145);
nand U18843 (N_18843,N_18632,N_18325);
and U18844 (N_18844,N_18530,N_18704);
xor U18845 (N_18845,N_18359,N_18679);
nand U18846 (N_18846,N_18716,N_18504);
nor U18847 (N_18847,N_18684,N_18333);
nand U18848 (N_18848,N_18607,N_18151);
nand U18849 (N_18849,N_18683,N_18473);
nor U18850 (N_18850,N_18456,N_18412);
or U18851 (N_18851,N_18480,N_18619);
xor U18852 (N_18852,N_18216,N_18620);
nor U18853 (N_18853,N_18432,N_18300);
xnor U18854 (N_18854,N_18326,N_18444);
nand U18855 (N_18855,N_18657,N_18417);
nand U18856 (N_18856,N_18706,N_18498);
xnor U18857 (N_18857,N_18129,N_18199);
nor U18858 (N_18858,N_18411,N_18130);
nor U18859 (N_18859,N_18351,N_18413);
or U18860 (N_18860,N_18160,N_18612);
or U18861 (N_18861,N_18445,N_18426);
nor U18862 (N_18862,N_18185,N_18507);
or U18863 (N_18863,N_18404,N_18164);
nand U18864 (N_18864,N_18353,N_18450);
nor U18865 (N_18865,N_18481,N_18570);
or U18866 (N_18866,N_18730,N_18242);
or U18867 (N_18867,N_18748,N_18680);
xnor U18868 (N_18868,N_18709,N_18749);
xnor U18869 (N_18869,N_18126,N_18593);
xnor U18870 (N_18870,N_18211,N_18181);
nor U18871 (N_18871,N_18701,N_18228);
nand U18872 (N_18872,N_18578,N_18736);
and U18873 (N_18873,N_18502,N_18276);
nor U18874 (N_18874,N_18493,N_18575);
nor U18875 (N_18875,N_18743,N_18250);
and U18876 (N_18876,N_18392,N_18471);
and U18877 (N_18877,N_18298,N_18236);
xor U18878 (N_18878,N_18522,N_18255);
nand U18879 (N_18879,N_18155,N_18394);
and U18880 (N_18880,N_18728,N_18630);
or U18881 (N_18881,N_18273,N_18487);
or U18882 (N_18882,N_18726,N_18430);
or U18883 (N_18883,N_18453,N_18734);
or U18884 (N_18884,N_18448,N_18168);
xnor U18885 (N_18885,N_18655,N_18309);
or U18886 (N_18886,N_18174,N_18220);
xor U18887 (N_18887,N_18261,N_18545);
nor U18888 (N_18888,N_18135,N_18616);
nand U18889 (N_18889,N_18637,N_18720);
nand U18890 (N_18890,N_18580,N_18585);
nor U18891 (N_18891,N_18624,N_18402);
or U18892 (N_18892,N_18447,N_18396);
and U18893 (N_18893,N_18279,N_18566);
xor U18894 (N_18894,N_18340,N_18606);
xnor U18895 (N_18895,N_18727,N_18489);
or U18896 (N_18896,N_18363,N_18254);
nand U18897 (N_18897,N_18383,N_18681);
and U18898 (N_18898,N_18213,N_18547);
xnor U18899 (N_18899,N_18159,N_18134);
nor U18900 (N_18900,N_18229,N_18674);
nor U18901 (N_18901,N_18375,N_18639);
or U18902 (N_18902,N_18622,N_18458);
and U18903 (N_18903,N_18724,N_18618);
nand U18904 (N_18904,N_18503,N_18591);
nor U18905 (N_18905,N_18688,N_18661);
nand U18906 (N_18906,N_18322,N_18237);
nor U18907 (N_18907,N_18635,N_18329);
and U18908 (N_18908,N_18132,N_18141);
and U18909 (N_18909,N_18197,N_18416);
and U18910 (N_18910,N_18492,N_18572);
and U18911 (N_18911,N_18166,N_18330);
nor U18912 (N_18912,N_18576,N_18425);
or U18913 (N_18913,N_18455,N_18240);
or U18914 (N_18914,N_18715,N_18568);
nor U18915 (N_18915,N_18305,N_18380);
xor U18916 (N_18916,N_18731,N_18395);
xor U18917 (N_18917,N_18464,N_18293);
nand U18918 (N_18918,N_18644,N_18339);
and U18919 (N_18919,N_18308,N_18640);
nor U18920 (N_18920,N_18446,N_18180);
and U18921 (N_18921,N_18310,N_18574);
nor U18922 (N_18922,N_18556,N_18163);
or U18923 (N_18923,N_18597,N_18138);
or U18924 (N_18924,N_18609,N_18610);
xnor U18925 (N_18925,N_18534,N_18614);
nor U18926 (N_18926,N_18342,N_18519);
nor U18927 (N_18927,N_18579,N_18590);
xnor U18928 (N_18928,N_18284,N_18550);
or U18929 (N_18929,N_18149,N_18352);
nand U18930 (N_18930,N_18370,N_18233);
xor U18931 (N_18931,N_18198,N_18311);
nor U18932 (N_18932,N_18719,N_18678);
or U18933 (N_18933,N_18257,N_18513);
xnor U18934 (N_18934,N_18291,N_18439);
nand U18935 (N_18935,N_18431,N_18171);
nand U18936 (N_18936,N_18685,N_18127);
nand U18937 (N_18937,N_18461,N_18350);
xnor U18938 (N_18938,N_18482,N_18332);
or U18939 (N_18939,N_18218,N_18408);
xor U18940 (N_18940,N_18582,N_18722);
or U18941 (N_18941,N_18642,N_18173);
nand U18942 (N_18942,N_18523,N_18665);
or U18943 (N_18943,N_18182,N_18746);
and U18944 (N_18944,N_18146,N_18144);
nand U18945 (N_18945,N_18323,N_18686);
xnor U18946 (N_18946,N_18170,N_18600);
xnor U18947 (N_18947,N_18158,N_18419);
nor U18948 (N_18948,N_18429,N_18601);
and U18949 (N_18949,N_18223,N_18406);
or U18950 (N_18950,N_18699,N_18649);
nand U18951 (N_18951,N_18347,N_18629);
and U18952 (N_18952,N_18485,N_18358);
nand U18953 (N_18953,N_18381,N_18296);
or U18954 (N_18954,N_18698,N_18289);
and U18955 (N_18955,N_18658,N_18673);
xor U18956 (N_18956,N_18239,N_18418);
nand U18957 (N_18957,N_18131,N_18264);
xnor U18958 (N_18958,N_18421,N_18397);
or U18959 (N_18959,N_18253,N_18594);
or U18960 (N_18960,N_18312,N_18336);
nor U18961 (N_18961,N_18475,N_18462);
and U18962 (N_18962,N_18707,N_18451);
nor U18963 (N_18963,N_18187,N_18742);
nand U18964 (N_18964,N_18226,N_18184);
and U18965 (N_18965,N_18466,N_18136);
nand U18966 (N_18966,N_18349,N_18659);
and U18967 (N_18967,N_18367,N_18745);
xor U18968 (N_18968,N_18542,N_18357);
nand U18969 (N_18969,N_18201,N_18667);
nand U18970 (N_18970,N_18337,N_18189);
nand U18971 (N_18971,N_18246,N_18423);
nand U18972 (N_18972,N_18474,N_18468);
or U18973 (N_18973,N_18338,N_18602);
or U18974 (N_18974,N_18647,N_18633);
or U18975 (N_18975,N_18403,N_18304);
and U18976 (N_18976,N_18631,N_18740);
nand U18977 (N_18977,N_18689,N_18266);
and U18978 (N_18978,N_18221,N_18703);
nor U18979 (N_18979,N_18378,N_18235);
nand U18980 (N_18980,N_18286,N_18301);
nand U18981 (N_18981,N_18203,N_18529);
or U18982 (N_18982,N_18713,N_18248);
nand U18983 (N_18983,N_18548,N_18588);
xnor U18984 (N_18984,N_18705,N_18596);
or U18985 (N_18985,N_18627,N_18526);
xor U18986 (N_18986,N_18650,N_18230);
or U18987 (N_18987,N_18672,N_18693);
nor U18988 (N_18988,N_18244,N_18299);
or U18989 (N_18989,N_18669,N_18562);
xor U18990 (N_18990,N_18275,N_18434);
and U18991 (N_18991,N_18643,N_18472);
xnor U18992 (N_18992,N_18483,N_18345);
xnor U18993 (N_18993,N_18660,N_18433);
or U18994 (N_18994,N_18467,N_18150);
or U18995 (N_18995,N_18497,N_18415);
or U18996 (N_18996,N_18729,N_18147);
nand U18997 (N_18997,N_18191,N_18505);
and U18998 (N_18998,N_18538,N_18137);
and U18999 (N_18999,N_18142,N_18454);
or U19000 (N_19000,N_18552,N_18428);
xnor U19001 (N_19001,N_18536,N_18222);
xnor U19002 (N_19002,N_18389,N_18664);
nor U19003 (N_19003,N_18491,N_18535);
xnor U19004 (N_19004,N_18613,N_18290);
or U19005 (N_19005,N_18723,N_18212);
or U19006 (N_19006,N_18318,N_18563);
nor U19007 (N_19007,N_18599,N_18320);
and U19008 (N_19008,N_18231,N_18281);
xnor U19009 (N_19009,N_18581,N_18192);
and U19010 (N_19010,N_18440,N_18501);
xnor U19011 (N_19011,N_18319,N_18437);
or U19012 (N_19012,N_18210,N_18478);
or U19013 (N_19013,N_18420,N_18587);
or U19014 (N_19014,N_18374,N_18407);
or U19015 (N_19015,N_18241,N_18274);
nor U19016 (N_19016,N_18532,N_18157);
xnor U19017 (N_19017,N_18294,N_18514);
or U19018 (N_19018,N_18410,N_18528);
and U19019 (N_19019,N_18651,N_18321);
or U19020 (N_19020,N_18165,N_18153);
and U19021 (N_19021,N_18341,N_18355);
and U19022 (N_19022,N_18559,N_18252);
and U19023 (N_19023,N_18143,N_18195);
nand U19024 (N_19024,N_18457,N_18156);
nand U19025 (N_19025,N_18744,N_18725);
or U19026 (N_19026,N_18443,N_18152);
and U19027 (N_19027,N_18179,N_18382);
or U19028 (N_19028,N_18626,N_18292);
nor U19029 (N_19029,N_18209,N_18196);
nand U19030 (N_19030,N_18277,N_18317);
xnor U19031 (N_19031,N_18270,N_18561);
nand U19032 (N_19032,N_18422,N_18549);
nor U19033 (N_19033,N_18267,N_18564);
xnor U19034 (N_19034,N_18676,N_18625);
xnor U19035 (N_19035,N_18656,N_18172);
nand U19036 (N_19036,N_18537,N_18125);
nor U19037 (N_19037,N_18214,N_18499);
or U19038 (N_19038,N_18272,N_18306);
nand U19039 (N_19039,N_18509,N_18605);
nand U19040 (N_19040,N_18190,N_18379);
or U19041 (N_19041,N_18331,N_18217);
nor U19042 (N_19042,N_18494,N_18377);
xnor U19043 (N_19043,N_18488,N_18712);
or U19044 (N_19044,N_18169,N_18508);
or U19045 (N_19045,N_18710,N_18747);
nand U19046 (N_19046,N_18335,N_18356);
and U19047 (N_19047,N_18589,N_18215);
and U19048 (N_19048,N_18479,N_18372);
xor U19049 (N_19049,N_18384,N_18540);
xor U19050 (N_19050,N_18500,N_18265);
xnor U19051 (N_19051,N_18714,N_18486);
nand U19052 (N_19052,N_18738,N_18414);
xnor U19053 (N_19053,N_18391,N_18194);
xnor U19054 (N_19054,N_18675,N_18224);
and U19055 (N_19055,N_18234,N_18225);
or U19056 (N_19056,N_18598,N_18544);
and U19057 (N_19057,N_18393,N_18569);
nand U19058 (N_19058,N_18543,N_18243);
or U19059 (N_19059,N_18541,N_18697);
or U19060 (N_19060,N_18484,N_18583);
nand U19061 (N_19061,N_18702,N_18495);
nand U19062 (N_19062,N_18733,N_18170);
or U19063 (N_19063,N_18176,N_18531);
and U19064 (N_19064,N_18462,N_18211);
nor U19065 (N_19065,N_18438,N_18360);
nand U19066 (N_19066,N_18612,N_18204);
and U19067 (N_19067,N_18479,N_18711);
xor U19068 (N_19068,N_18549,N_18337);
or U19069 (N_19069,N_18395,N_18492);
xor U19070 (N_19070,N_18419,N_18587);
xor U19071 (N_19071,N_18227,N_18632);
and U19072 (N_19072,N_18298,N_18254);
or U19073 (N_19073,N_18498,N_18664);
or U19074 (N_19074,N_18353,N_18413);
or U19075 (N_19075,N_18251,N_18295);
xor U19076 (N_19076,N_18557,N_18700);
nand U19077 (N_19077,N_18738,N_18364);
or U19078 (N_19078,N_18717,N_18384);
or U19079 (N_19079,N_18381,N_18362);
or U19080 (N_19080,N_18345,N_18276);
or U19081 (N_19081,N_18661,N_18580);
and U19082 (N_19082,N_18370,N_18502);
nand U19083 (N_19083,N_18596,N_18493);
or U19084 (N_19084,N_18146,N_18236);
or U19085 (N_19085,N_18581,N_18343);
and U19086 (N_19086,N_18432,N_18509);
and U19087 (N_19087,N_18396,N_18342);
xnor U19088 (N_19088,N_18491,N_18413);
and U19089 (N_19089,N_18291,N_18485);
xor U19090 (N_19090,N_18135,N_18195);
nor U19091 (N_19091,N_18553,N_18229);
xnor U19092 (N_19092,N_18574,N_18620);
and U19093 (N_19093,N_18642,N_18644);
and U19094 (N_19094,N_18567,N_18612);
nand U19095 (N_19095,N_18516,N_18238);
nand U19096 (N_19096,N_18323,N_18180);
nor U19097 (N_19097,N_18728,N_18411);
or U19098 (N_19098,N_18299,N_18372);
and U19099 (N_19099,N_18332,N_18629);
or U19100 (N_19100,N_18504,N_18367);
or U19101 (N_19101,N_18407,N_18717);
or U19102 (N_19102,N_18411,N_18568);
nor U19103 (N_19103,N_18189,N_18199);
nand U19104 (N_19104,N_18490,N_18615);
nand U19105 (N_19105,N_18448,N_18345);
and U19106 (N_19106,N_18551,N_18443);
or U19107 (N_19107,N_18631,N_18247);
or U19108 (N_19108,N_18400,N_18299);
nor U19109 (N_19109,N_18385,N_18313);
xor U19110 (N_19110,N_18476,N_18588);
nand U19111 (N_19111,N_18229,N_18545);
xor U19112 (N_19112,N_18284,N_18490);
xor U19113 (N_19113,N_18439,N_18562);
or U19114 (N_19114,N_18525,N_18286);
nand U19115 (N_19115,N_18163,N_18624);
nand U19116 (N_19116,N_18226,N_18141);
nand U19117 (N_19117,N_18517,N_18278);
xor U19118 (N_19118,N_18219,N_18612);
nand U19119 (N_19119,N_18161,N_18229);
and U19120 (N_19120,N_18697,N_18295);
xor U19121 (N_19121,N_18325,N_18353);
nor U19122 (N_19122,N_18699,N_18430);
and U19123 (N_19123,N_18159,N_18201);
or U19124 (N_19124,N_18425,N_18299);
nor U19125 (N_19125,N_18697,N_18392);
nand U19126 (N_19126,N_18476,N_18571);
nand U19127 (N_19127,N_18521,N_18168);
and U19128 (N_19128,N_18603,N_18643);
or U19129 (N_19129,N_18711,N_18181);
nor U19130 (N_19130,N_18577,N_18447);
or U19131 (N_19131,N_18711,N_18577);
nor U19132 (N_19132,N_18469,N_18137);
and U19133 (N_19133,N_18427,N_18137);
and U19134 (N_19134,N_18545,N_18493);
nand U19135 (N_19135,N_18222,N_18619);
and U19136 (N_19136,N_18666,N_18560);
nand U19137 (N_19137,N_18414,N_18196);
or U19138 (N_19138,N_18545,N_18689);
xor U19139 (N_19139,N_18246,N_18589);
or U19140 (N_19140,N_18686,N_18288);
nand U19141 (N_19141,N_18411,N_18298);
nand U19142 (N_19142,N_18410,N_18713);
and U19143 (N_19143,N_18379,N_18466);
and U19144 (N_19144,N_18722,N_18681);
and U19145 (N_19145,N_18418,N_18616);
or U19146 (N_19146,N_18371,N_18435);
and U19147 (N_19147,N_18699,N_18308);
nor U19148 (N_19148,N_18519,N_18302);
or U19149 (N_19149,N_18229,N_18495);
xor U19150 (N_19150,N_18283,N_18411);
and U19151 (N_19151,N_18592,N_18481);
xnor U19152 (N_19152,N_18724,N_18303);
xor U19153 (N_19153,N_18323,N_18452);
nand U19154 (N_19154,N_18480,N_18220);
or U19155 (N_19155,N_18680,N_18449);
nand U19156 (N_19156,N_18193,N_18519);
xor U19157 (N_19157,N_18426,N_18334);
xor U19158 (N_19158,N_18583,N_18607);
nor U19159 (N_19159,N_18128,N_18535);
or U19160 (N_19160,N_18673,N_18160);
xnor U19161 (N_19161,N_18218,N_18257);
and U19162 (N_19162,N_18311,N_18335);
or U19163 (N_19163,N_18727,N_18646);
nand U19164 (N_19164,N_18207,N_18294);
and U19165 (N_19165,N_18201,N_18242);
and U19166 (N_19166,N_18600,N_18398);
or U19167 (N_19167,N_18531,N_18749);
nand U19168 (N_19168,N_18192,N_18254);
nor U19169 (N_19169,N_18488,N_18329);
and U19170 (N_19170,N_18376,N_18706);
nor U19171 (N_19171,N_18684,N_18581);
nand U19172 (N_19172,N_18688,N_18332);
nor U19173 (N_19173,N_18743,N_18136);
or U19174 (N_19174,N_18166,N_18599);
or U19175 (N_19175,N_18511,N_18580);
and U19176 (N_19176,N_18243,N_18367);
or U19177 (N_19177,N_18546,N_18541);
or U19178 (N_19178,N_18550,N_18285);
nand U19179 (N_19179,N_18353,N_18415);
nand U19180 (N_19180,N_18315,N_18345);
xor U19181 (N_19181,N_18267,N_18713);
or U19182 (N_19182,N_18161,N_18624);
and U19183 (N_19183,N_18636,N_18719);
nor U19184 (N_19184,N_18312,N_18627);
and U19185 (N_19185,N_18274,N_18552);
nand U19186 (N_19186,N_18380,N_18263);
and U19187 (N_19187,N_18746,N_18176);
nor U19188 (N_19188,N_18152,N_18191);
xor U19189 (N_19189,N_18673,N_18473);
and U19190 (N_19190,N_18343,N_18219);
nand U19191 (N_19191,N_18258,N_18435);
and U19192 (N_19192,N_18210,N_18384);
or U19193 (N_19193,N_18417,N_18531);
or U19194 (N_19194,N_18447,N_18579);
or U19195 (N_19195,N_18676,N_18549);
or U19196 (N_19196,N_18268,N_18433);
and U19197 (N_19197,N_18675,N_18368);
nand U19198 (N_19198,N_18639,N_18339);
nand U19199 (N_19199,N_18619,N_18728);
xor U19200 (N_19200,N_18314,N_18506);
xor U19201 (N_19201,N_18135,N_18597);
or U19202 (N_19202,N_18270,N_18505);
or U19203 (N_19203,N_18385,N_18170);
nor U19204 (N_19204,N_18399,N_18250);
nor U19205 (N_19205,N_18673,N_18398);
nand U19206 (N_19206,N_18166,N_18346);
and U19207 (N_19207,N_18251,N_18261);
nor U19208 (N_19208,N_18284,N_18189);
nand U19209 (N_19209,N_18304,N_18490);
xor U19210 (N_19210,N_18564,N_18269);
or U19211 (N_19211,N_18211,N_18690);
nor U19212 (N_19212,N_18490,N_18397);
and U19213 (N_19213,N_18278,N_18141);
nor U19214 (N_19214,N_18738,N_18498);
or U19215 (N_19215,N_18434,N_18479);
nand U19216 (N_19216,N_18673,N_18589);
xnor U19217 (N_19217,N_18286,N_18429);
and U19218 (N_19218,N_18441,N_18290);
and U19219 (N_19219,N_18270,N_18320);
nand U19220 (N_19220,N_18516,N_18571);
xor U19221 (N_19221,N_18678,N_18401);
nand U19222 (N_19222,N_18616,N_18137);
and U19223 (N_19223,N_18280,N_18473);
xor U19224 (N_19224,N_18314,N_18234);
and U19225 (N_19225,N_18507,N_18207);
and U19226 (N_19226,N_18430,N_18152);
nor U19227 (N_19227,N_18562,N_18730);
and U19228 (N_19228,N_18383,N_18453);
or U19229 (N_19229,N_18406,N_18650);
xor U19230 (N_19230,N_18240,N_18629);
xnor U19231 (N_19231,N_18448,N_18335);
and U19232 (N_19232,N_18247,N_18283);
xor U19233 (N_19233,N_18394,N_18596);
or U19234 (N_19234,N_18265,N_18647);
or U19235 (N_19235,N_18362,N_18517);
nand U19236 (N_19236,N_18518,N_18645);
or U19237 (N_19237,N_18512,N_18645);
xor U19238 (N_19238,N_18305,N_18550);
nor U19239 (N_19239,N_18557,N_18422);
or U19240 (N_19240,N_18692,N_18535);
and U19241 (N_19241,N_18459,N_18283);
or U19242 (N_19242,N_18320,N_18664);
xor U19243 (N_19243,N_18302,N_18307);
or U19244 (N_19244,N_18285,N_18302);
and U19245 (N_19245,N_18427,N_18654);
nand U19246 (N_19246,N_18148,N_18163);
or U19247 (N_19247,N_18612,N_18189);
nand U19248 (N_19248,N_18133,N_18739);
nand U19249 (N_19249,N_18400,N_18690);
nand U19250 (N_19250,N_18396,N_18712);
xor U19251 (N_19251,N_18439,N_18235);
xnor U19252 (N_19252,N_18749,N_18193);
or U19253 (N_19253,N_18482,N_18424);
and U19254 (N_19254,N_18215,N_18273);
and U19255 (N_19255,N_18319,N_18245);
xor U19256 (N_19256,N_18403,N_18320);
or U19257 (N_19257,N_18608,N_18741);
nand U19258 (N_19258,N_18634,N_18260);
or U19259 (N_19259,N_18324,N_18749);
xnor U19260 (N_19260,N_18422,N_18463);
and U19261 (N_19261,N_18482,N_18262);
nor U19262 (N_19262,N_18488,N_18553);
and U19263 (N_19263,N_18252,N_18283);
nand U19264 (N_19264,N_18284,N_18637);
nand U19265 (N_19265,N_18706,N_18238);
and U19266 (N_19266,N_18521,N_18598);
xor U19267 (N_19267,N_18295,N_18695);
nor U19268 (N_19268,N_18180,N_18356);
xnor U19269 (N_19269,N_18689,N_18331);
nand U19270 (N_19270,N_18142,N_18718);
and U19271 (N_19271,N_18703,N_18631);
nand U19272 (N_19272,N_18275,N_18736);
and U19273 (N_19273,N_18186,N_18449);
or U19274 (N_19274,N_18227,N_18445);
nand U19275 (N_19275,N_18527,N_18514);
and U19276 (N_19276,N_18223,N_18383);
nand U19277 (N_19277,N_18569,N_18150);
xnor U19278 (N_19278,N_18323,N_18176);
and U19279 (N_19279,N_18416,N_18610);
nor U19280 (N_19280,N_18243,N_18617);
or U19281 (N_19281,N_18587,N_18466);
and U19282 (N_19282,N_18520,N_18512);
or U19283 (N_19283,N_18165,N_18698);
nand U19284 (N_19284,N_18550,N_18712);
xor U19285 (N_19285,N_18318,N_18699);
nor U19286 (N_19286,N_18620,N_18193);
or U19287 (N_19287,N_18440,N_18251);
nand U19288 (N_19288,N_18214,N_18159);
or U19289 (N_19289,N_18514,N_18300);
or U19290 (N_19290,N_18741,N_18271);
and U19291 (N_19291,N_18170,N_18743);
nand U19292 (N_19292,N_18295,N_18621);
or U19293 (N_19293,N_18276,N_18520);
or U19294 (N_19294,N_18583,N_18501);
xnor U19295 (N_19295,N_18199,N_18266);
xor U19296 (N_19296,N_18584,N_18466);
nand U19297 (N_19297,N_18542,N_18275);
or U19298 (N_19298,N_18659,N_18672);
or U19299 (N_19299,N_18670,N_18460);
or U19300 (N_19300,N_18409,N_18306);
or U19301 (N_19301,N_18743,N_18255);
nand U19302 (N_19302,N_18472,N_18203);
or U19303 (N_19303,N_18347,N_18169);
and U19304 (N_19304,N_18407,N_18661);
and U19305 (N_19305,N_18564,N_18567);
nor U19306 (N_19306,N_18441,N_18208);
or U19307 (N_19307,N_18329,N_18184);
xnor U19308 (N_19308,N_18622,N_18717);
or U19309 (N_19309,N_18202,N_18500);
and U19310 (N_19310,N_18433,N_18157);
or U19311 (N_19311,N_18167,N_18475);
or U19312 (N_19312,N_18651,N_18370);
nor U19313 (N_19313,N_18284,N_18494);
xor U19314 (N_19314,N_18274,N_18219);
or U19315 (N_19315,N_18281,N_18254);
xor U19316 (N_19316,N_18527,N_18595);
or U19317 (N_19317,N_18203,N_18184);
nor U19318 (N_19318,N_18441,N_18196);
xor U19319 (N_19319,N_18725,N_18156);
xnor U19320 (N_19320,N_18433,N_18422);
or U19321 (N_19321,N_18616,N_18400);
nand U19322 (N_19322,N_18633,N_18729);
or U19323 (N_19323,N_18532,N_18405);
nand U19324 (N_19324,N_18476,N_18454);
xor U19325 (N_19325,N_18368,N_18217);
nand U19326 (N_19326,N_18249,N_18394);
xor U19327 (N_19327,N_18195,N_18399);
nor U19328 (N_19328,N_18328,N_18567);
nand U19329 (N_19329,N_18509,N_18234);
xnor U19330 (N_19330,N_18276,N_18140);
xnor U19331 (N_19331,N_18692,N_18502);
and U19332 (N_19332,N_18732,N_18298);
nand U19333 (N_19333,N_18169,N_18723);
nor U19334 (N_19334,N_18476,N_18722);
or U19335 (N_19335,N_18169,N_18354);
or U19336 (N_19336,N_18151,N_18161);
xnor U19337 (N_19337,N_18196,N_18396);
nor U19338 (N_19338,N_18615,N_18605);
nand U19339 (N_19339,N_18165,N_18579);
nor U19340 (N_19340,N_18678,N_18339);
nor U19341 (N_19341,N_18418,N_18541);
and U19342 (N_19342,N_18622,N_18401);
nor U19343 (N_19343,N_18631,N_18143);
nor U19344 (N_19344,N_18345,N_18412);
xnor U19345 (N_19345,N_18577,N_18530);
nor U19346 (N_19346,N_18194,N_18153);
xnor U19347 (N_19347,N_18165,N_18675);
and U19348 (N_19348,N_18420,N_18173);
nor U19349 (N_19349,N_18607,N_18490);
or U19350 (N_19350,N_18625,N_18566);
xor U19351 (N_19351,N_18264,N_18446);
xor U19352 (N_19352,N_18309,N_18534);
and U19353 (N_19353,N_18357,N_18654);
xnor U19354 (N_19354,N_18488,N_18572);
and U19355 (N_19355,N_18727,N_18586);
xor U19356 (N_19356,N_18214,N_18210);
xor U19357 (N_19357,N_18686,N_18640);
xor U19358 (N_19358,N_18286,N_18450);
and U19359 (N_19359,N_18171,N_18337);
nor U19360 (N_19360,N_18576,N_18347);
or U19361 (N_19361,N_18129,N_18637);
nand U19362 (N_19362,N_18454,N_18362);
and U19363 (N_19363,N_18718,N_18399);
nand U19364 (N_19364,N_18361,N_18491);
nand U19365 (N_19365,N_18333,N_18673);
or U19366 (N_19366,N_18575,N_18159);
nand U19367 (N_19367,N_18430,N_18443);
or U19368 (N_19368,N_18279,N_18373);
and U19369 (N_19369,N_18512,N_18221);
and U19370 (N_19370,N_18531,N_18539);
nand U19371 (N_19371,N_18227,N_18161);
and U19372 (N_19372,N_18405,N_18669);
and U19373 (N_19373,N_18723,N_18234);
xnor U19374 (N_19374,N_18505,N_18236);
nand U19375 (N_19375,N_18976,N_19038);
xnor U19376 (N_19376,N_19280,N_19103);
nand U19377 (N_19377,N_18830,N_19279);
nor U19378 (N_19378,N_18891,N_18769);
xnor U19379 (N_19379,N_19067,N_19239);
and U19380 (N_19380,N_18906,N_19299);
xnor U19381 (N_19381,N_19025,N_18867);
or U19382 (N_19382,N_19137,N_19310);
or U19383 (N_19383,N_19153,N_19043);
and U19384 (N_19384,N_19223,N_19284);
nand U19385 (N_19385,N_18839,N_18890);
nand U19386 (N_19386,N_19057,N_19085);
xnor U19387 (N_19387,N_19018,N_19350);
and U19388 (N_19388,N_18824,N_19076);
xor U19389 (N_19389,N_19050,N_18899);
xnor U19390 (N_19390,N_18852,N_18962);
xnor U19391 (N_19391,N_18878,N_19119);
nor U19392 (N_19392,N_19300,N_18975);
or U19393 (N_19393,N_19361,N_18799);
xnor U19394 (N_19394,N_19194,N_19078);
or U19395 (N_19395,N_19183,N_19068);
or U19396 (N_19396,N_19154,N_18866);
and U19397 (N_19397,N_18970,N_18996);
nor U19398 (N_19398,N_19215,N_19210);
or U19399 (N_19399,N_19247,N_18893);
and U19400 (N_19400,N_19147,N_18993);
nand U19401 (N_19401,N_19218,N_18951);
and U19402 (N_19402,N_18889,N_19165);
and U19403 (N_19403,N_19164,N_19285);
nor U19404 (N_19404,N_19358,N_19344);
nand U19405 (N_19405,N_19090,N_19357);
or U19406 (N_19406,N_19211,N_19092);
or U19407 (N_19407,N_18948,N_19229);
and U19408 (N_19408,N_18800,N_19347);
and U19409 (N_19409,N_19008,N_19161);
and U19410 (N_19410,N_19248,N_19323);
xor U19411 (N_19411,N_18916,N_19116);
nor U19412 (N_19412,N_19151,N_18759);
or U19413 (N_19413,N_19332,N_19065);
nor U19414 (N_19414,N_19301,N_18917);
xor U19415 (N_19415,N_18922,N_19261);
or U19416 (N_19416,N_18757,N_19062);
nand U19417 (N_19417,N_18949,N_19288);
or U19418 (N_19418,N_19349,N_19077);
nor U19419 (N_19419,N_19101,N_18971);
nand U19420 (N_19420,N_19338,N_18877);
nor U19421 (N_19421,N_18921,N_19345);
nand U19422 (N_19422,N_18946,N_19040);
nor U19423 (N_19423,N_18904,N_18765);
xor U19424 (N_19424,N_18811,N_19172);
and U19425 (N_19425,N_19331,N_18766);
nor U19426 (N_19426,N_18752,N_18809);
and U19427 (N_19427,N_19179,N_18911);
and U19428 (N_19428,N_18961,N_19024);
xor U19429 (N_19429,N_19100,N_19204);
and U19430 (N_19430,N_18858,N_19305);
xor U19431 (N_19431,N_19139,N_19199);
nor U19432 (N_19432,N_19023,N_19182);
xor U19433 (N_19433,N_19083,N_19028);
xnor U19434 (N_19434,N_18837,N_18872);
and U19435 (N_19435,N_19333,N_19328);
xnor U19436 (N_19436,N_18793,N_18771);
nand U19437 (N_19437,N_18941,N_19200);
nor U19438 (N_19438,N_19070,N_19264);
nor U19439 (N_19439,N_18826,N_18779);
xnor U19440 (N_19440,N_19041,N_18843);
nand U19441 (N_19441,N_18859,N_19011);
nor U19442 (N_19442,N_19074,N_19155);
or U19443 (N_19443,N_19181,N_19242);
or U19444 (N_19444,N_18784,N_18959);
or U19445 (N_19445,N_19112,N_19001);
nand U19446 (N_19446,N_18855,N_18810);
and U19447 (N_19447,N_19069,N_18817);
xnor U19448 (N_19448,N_19118,N_18767);
nor U19449 (N_19449,N_19304,N_19167);
nor U19450 (N_19450,N_19340,N_19162);
nor U19451 (N_19451,N_18907,N_19108);
nand U19452 (N_19452,N_18992,N_18838);
nand U19453 (N_19453,N_18945,N_19031);
nand U19454 (N_19454,N_18968,N_19311);
and U19455 (N_19455,N_19273,N_18832);
nand U19456 (N_19456,N_18823,N_18818);
nor U19457 (N_19457,N_19291,N_19262);
and U19458 (N_19458,N_18815,N_19005);
and U19459 (N_19459,N_19292,N_18820);
nand U19460 (N_19460,N_19370,N_19134);
and U19461 (N_19461,N_19277,N_19205);
xnor U19462 (N_19462,N_19135,N_19207);
or U19463 (N_19463,N_19079,N_18896);
xnor U19464 (N_19464,N_19243,N_18750);
nand U19465 (N_19465,N_19208,N_18788);
xnor U19466 (N_19466,N_18913,N_19368);
and U19467 (N_19467,N_19145,N_18955);
xor U19468 (N_19468,N_18834,N_19187);
nand U19469 (N_19469,N_19244,N_19056);
xor U19470 (N_19470,N_19237,N_18930);
nor U19471 (N_19471,N_18887,N_18812);
nand U19472 (N_19472,N_19163,N_18933);
xor U19473 (N_19473,N_18997,N_19255);
nor U19474 (N_19474,N_18984,N_18846);
nor U19475 (N_19475,N_18861,N_19158);
nor U19476 (N_19476,N_18895,N_19221);
xor U19477 (N_19477,N_19317,N_18844);
and U19478 (N_19478,N_19166,N_19289);
nor U19479 (N_19479,N_19193,N_19206);
nand U19480 (N_19480,N_19130,N_19259);
xnor U19481 (N_19481,N_19294,N_19348);
xor U19482 (N_19482,N_19306,N_19086);
nor U19483 (N_19483,N_18883,N_18853);
nand U19484 (N_19484,N_19203,N_19327);
nor U19485 (N_19485,N_18956,N_18927);
nand U19486 (N_19486,N_19125,N_19274);
nand U19487 (N_19487,N_18847,N_18792);
and U19488 (N_19488,N_18821,N_19335);
nand U19489 (N_19489,N_18778,N_19060);
and U19490 (N_19490,N_18775,N_18776);
nor U19491 (N_19491,N_18768,N_19019);
and U19492 (N_19492,N_18786,N_19231);
xor U19493 (N_19493,N_18967,N_18937);
nand U19494 (N_19494,N_19293,N_19282);
nand U19495 (N_19495,N_18915,N_19087);
xnor U19496 (N_19496,N_18787,N_18963);
or U19497 (N_19497,N_19270,N_19250);
and U19498 (N_19498,N_19230,N_18989);
and U19499 (N_19499,N_19141,N_18923);
xor U19500 (N_19500,N_19322,N_18785);
nor U19501 (N_19501,N_19089,N_19283);
xnor U19502 (N_19502,N_19022,N_19110);
nand U19503 (N_19503,N_18762,N_19275);
and U19504 (N_19504,N_18790,N_18851);
or U19505 (N_19505,N_18990,N_18802);
nand U19506 (N_19506,N_18944,N_19029);
nand U19507 (N_19507,N_19126,N_18758);
nor U19508 (N_19508,N_19149,N_19140);
and U19509 (N_19509,N_19003,N_19296);
xnor U19510 (N_19510,N_19160,N_18873);
nor U19511 (N_19511,N_19354,N_19257);
nor U19512 (N_19512,N_19342,N_18777);
nor U19513 (N_19513,N_19346,N_18957);
xor U19514 (N_19514,N_18881,N_19298);
nor U19515 (N_19515,N_19343,N_19114);
and U19516 (N_19516,N_19326,N_18804);
nand U19517 (N_19517,N_18979,N_18860);
nor U19518 (N_19518,N_18870,N_18986);
or U19519 (N_19519,N_18991,N_19044);
and U19520 (N_19520,N_18874,N_19096);
nor U19521 (N_19521,N_19364,N_19012);
or U19522 (N_19522,N_18836,N_18931);
and U19523 (N_19523,N_19321,N_18876);
nand U19524 (N_19524,N_19088,N_18958);
nand U19525 (N_19525,N_19104,N_19272);
and U19526 (N_19526,N_19026,N_18763);
and U19527 (N_19527,N_18950,N_18869);
nor U19528 (N_19528,N_19302,N_19233);
xor U19529 (N_19529,N_18995,N_18914);
nor U19530 (N_19530,N_18938,N_19325);
or U19531 (N_19531,N_19117,N_19109);
and U19532 (N_19532,N_19314,N_18791);
nor U19533 (N_19533,N_19152,N_19316);
nor U19534 (N_19534,N_19032,N_19016);
nor U19535 (N_19535,N_19303,N_19020);
or U19536 (N_19536,N_18978,N_19168);
xnor U19537 (N_19537,N_19170,N_19127);
nor U19538 (N_19538,N_19055,N_18863);
or U19539 (N_19539,N_18875,N_19099);
nand U19540 (N_19540,N_19120,N_18789);
and U19541 (N_19541,N_18756,N_19312);
xor U19542 (N_19542,N_18828,N_18935);
and U19543 (N_19543,N_18934,N_18928);
nand U19544 (N_19544,N_18833,N_18973);
nor U19545 (N_19545,N_18761,N_19045);
nor U19546 (N_19546,N_18902,N_18982);
or U19547 (N_19547,N_19202,N_19241);
xnor U19548 (N_19548,N_19105,N_19013);
and U19549 (N_19549,N_19171,N_19146);
and U19550 (N_19550,N_19186,N_19269);
and U19551 (N_19551,N_19226,N_19320);
or U19552 (N_19552,N_19128,N_18829);
or U19553 (N_19553,N_19124,N_19004);
xnor U19554 (N_19554,N_19198,N_19192);
and U19555 (N_19555,N_19021,N_18926);
and U19556 (N_19556,N_18856,N_18754);
or U19557 (N_19557,N_19220,N_18783);
xor U19558 (N_19558,N_19196,N_19049);
nor U19559 (N_19559,N_19010,N_18831);
or U19560 (N_19560,N_18857,N_18888);
xor U19561 (N_19561,N_18764,N_18901);
xnor U19562 (N_19562,N_18920,N_19066);
or U19563 (N_19563,N_18980,N_18868);
or U19564 (N_19564,N_19365,N_19271);
nand U19565 (N_19565,N_19330,N_19093);
and U19566 (N_19566,N_18942,N_19318);
or U19567 (N_19567,N_19295,N_19156);
or U19568 (N_19568,N_19334,N_19249);
nor U19569 (N_19569,N_19138,N_18835);
nor U19570 (N_19570,N_18772,N_19268);
xor U19571 (N_19571,N_18912,N_18849);
and U19572 (N_19572,N_18987,N_19058);
nand U19573 (N_19573,N_19366,N_18947);
or U19574 (N_19574,N_19121,N_19142);
nand U19575 (N_19575,N_18994,N_19191);
and U19576 (N_19576,N_19097,N_18903);
nor U19577 (N_19577,N_19341,N_19176);
xnor U19578 (N_19578,N_19209,N_19260);
or U19579 (N_19579,N_19132,N_18964);
xor U19580 (N_19580,N_19102,N_19039);
and U19581 (N_19581,N_18862,N_19190);
and U19582 (N_19582,N_19113,N_18825);
nor U19583 (N_19583,N_19228,N_18977);
and U19584 (N_19584,N_19048,N_19094);
or U19585 (N_19585,N_18885,N_18753);
xor U19586 (N_19586,N_19222,N_18880);
nand U19587 (N_19587,N_19173,N_18774);
xnor U19588 (N_19588,N_18755,N_19053);
xnor U19589 (N_19589,N_19315,N_19189);
xor U19590 (N_19590,N_18966,N_18919);
xnor U19591 (N_19591,N_18988,N_18770);
nand U19592 (N_19592,N_18816,N_19148);
xnor U19593 (N_19593,N_19174,N_18794);
and U19594 (N_19594,N_19051,N_19355);
nor U19595 (N_19595,N_18819,N_18939);
xor U19596 (N_19596,N_18796,N_19232);
and U19597 (N_19597,N_18905,N_19219);
xor U19598 (N_19598,N_19336,N_19033);
and U19599 (N_19599,N_19224,N_19324);
xor U19600 (N_19600,N_19238,N_18751);
nor U19601 (N_19601,N_19253,N_19015);
or U19602 (N_19602,N_19072,N_19374);
and U19603 (N_19603,N_19007,N_19256);
nor U19604 (N_19604,N_18918,N_19000);
and U19605 (N_19605,N_18865,N_18960);
xnor U19606 (N_19606,N_19278,N_19236);
xor U19607 (N_19607,N_18854,N_19184);
nor U19608 (N_19608,N_19235,N_19061);
and U19609 (N_19609,N_18892,N_18882);
nor U19610 (N_19610,N_18925,N_18943);
and U19611 (N_19611,N_19265,N_19240);
nand U19612 (N_19612,N_19360,N_19267);
or U19613 (N_19613,N_19046,N_19014);
xor U19614 (N_19614,N_18886,N_18952);
xnor U19615 (N_19615,N_19245,N_19201);
nand U19616 (N_19616,N_18822,N_18999);
and U19617 (N_19617,N_19054,N_19185);
nor U19618 (N_19618,N_18841,N_18936);
xor U19619 (N_19619,N_18798,N_19002);
nor U19620 (N_19620,N_19106,N_18780);
xnor U19621 (N_19621,N_19175,N_19212);
xnor U19622 (N_19622,N_19254,N_19107);
xnor U19623 (N_19623,N_19286,N_19136);
xor U19624 (N_19624,N_19082,N_19178);
nand U19625 (N_19625,N_19351,N_18840);
xor U19626 (N_19626,N_19372,N_19246);
nand U19627 (N_19627,N_19006,N_18940);
and U19628 (N_19628,N_18908,N_19263);
nand U19629 (N_19629,N_18897,N_19071);
nand U19630 (N_19630,N_19367,N_19214);
and U19631 (N_19631,N_18781,N_19266);
and U19632 (N_19632,N_19225,N_19159);
or U19633 (N_19633,N_18807,N_19091);
and U19634 (N_19634,N_18814,N_18909);
nand U19635 (N_19635,N_19115,N_19339);
xnor U19636 (N_19636,N_18827,N_18898);
nand U19637 (N_19637,N_19098,N_19371);
or U19638 (N_19638,N_19290,N_19063);
nor U19639 (N_19639,N_19297,N_18801);
or U19640 (N_19640,N_18954,N_19059);
and U19641 (N_19641,N_19133,N_18965);
nor U19642 (N_19642,N_19177,N_19227);
or U19643 (N_19643,N_19150,N_19037);
xor U19644 (N_19644,N_19197,N_19251);
or U19645 (N_19645,N_19144,N_19123);
or U19646 (N_19646,N_19035,N_19009);
nor U19647 (N_19647,N_19359,N_19213);
nand U19648 (N_19648,N_19075,N_18797);
nor U19649 (N_19649,N_18924,N_19180);
nor U19650 (N_19650,N_19373,N_19129);
nor U19651 (N_19651,N_19188,N_18894);
xor U19652 (N_19652,N_19362,N_18782);
or U19653 (N_19653,N_19095,N_19042);
or U19654 (N_19654,N_18864,N_18953);
nor U19655 (N_19655,N_18972,N_19308);
nand U19656 (N_19656,N_19369,N_19027);
nand U19657 (N_19657,N_18932,N_19131);
xor U19658 (N_19658,N_19080,N_19047);
nor U19659 (N_19659,N_19169,N_19353);
nand U19660 (N_19660,N_19307,N_18773);
and U19661 (N_19661,N_18884,N_19034);
nand U19662 (N_19662,N_18929,N_18848);
nor U19663 (N_19663,N_18974,N_18910);
and U19664 (N_19664,N_19052,N_18803);
or U19665 (N_19665,N_18795,N_18805);
nand U19666 (N_19666,N_19319,N_19036);
and U19667 (N_19667,N_18998,N_19143);
nand U19668 (N_19668,N_19122,N_18983);
xor U19669 (N_19669,N_19111,N_18842);
or U19670 (N_19670,N_18981,N_19356);
or U19671 (N_19671,N_19017,N_19313);
nand U19672 (N_19672,N_19234,N_19073);
xnor U19673 (N_19673,N_19309,N_19363);
or U19674 (N_19674,N_19030,N_19081);
nand U19675 (N_19675,N_19276,N_18871);
nand U19676 (N_19676,N_19352,N_19217);
and U19677 (N_19677,N_18845,N_19157);
and U19678 (N_19678,N_19281,N_19258);
and U19679 (N_19679,N_18850,N_18813);
nor U19680 (N_19680,N_19329,N_18879);
xnor U19681 (N_19681,N_19216,N_19287);
nand U19682 (N_19682,N_18969,N_18760);
nor U19683 (N_19683,N_19084,N_19064);
nor U19684 (N_19684,N_18806,N_19252);
and U19685 (N_19685,N_19195,N_19337);
nand U19686 (N_19686,N_18900,N_18985);
xnor U19687 (N_19687,N_18808,N_19005);
or U19688 (N_19688,N_19082,N_19105);
xnor U19689 (N_19689,N_19091,N_19287);
nor U19690 (N_19690,N_18769,N_18816);
nor U19691 (N_19691,N_19286,N_19124);
and U19692 (N_19692,N_18796,N_19203);
or U19693 (N_19693,N_18830,N_18979);
and U19694 (N_19694,N_19267,N_18922);
or U19695 (N_19695,N_19010,N_19302);
and U19696 (N_19696,N_18908,N_19193);
nor U19697 (N_19697,N_18873,N_18987);
xor U19698 (N_19698,N_19068,N_19250);
xnor U19699 (N_19699,N_19042,N_18872);
nor U19700 (N_19700,N_18795,N_19274);
and U19701 (N_19701,N_19294,N_19072);
nor U19702 (N_19702,N_19270,N_18918);
and U19703 (N_19703,N_19286,N_18789);
nor U19704 (N_19704,N_18918,N_18979);
nand U19705 (N_19705,N_19140,N_19092);
xor U19706 (N_19706,N_18842,N_18936);
nor U19707 (N_19707,N_18857,N_18880);
nand U19708 (N_19708,N_18830,N_18784);
nor U19709 (N_19709,N_19307,N_18809);
nand U19710 (N_19710,N_18884,N_19142);
nand U19711 (N_19711,N_18859,N_19323);
nor U19712 (N_19712,N_19176,N_19253);
or U19713 (N_19713,N_19225,N_19145);
xor U19714 (N_19714,N_19145,N_18757);
xor U19715 (N_19715,N_19153,N_19304);
or U19716 (N_19716,N_19184,N_19144);
nand U19717 (N_19717,N_19032,N_19373);
xor U19718 (N_19718,N_19322,N_19110);
or U19719 (N_19719,N_18994,N_19118);
xnor U19720 (N_19720,N_19264,N_19239);
nor U19721 (N_19721,N_19356,N_19100);
or U19722 (N_19722,N_18940,N_18773);
nand U19723 (N_19723,N_19191,N_19232);
nor U19724 (N_19724,N_19165,N_19319);
or U19725 (N_19725,N_18844,N_18944);
xnor U19726 (N_19726,N_19202,N_19173);
nor U19727 (N_19727,N_18885,N_19040);
and U19728 (N_19728,N_19072,N_19057);
xnor U19729 (N_19729,N_19164,N_18772);
nand U19730 (N_19730,N_18893,N_19124);
xor U19731 (N_19731,N_19336,N_18939);
nor U19732 (N_19732,N_19086,N_18886);
or U19733 (N_19733,N_19000,N_18936);
xnor U19734 (N_19734,N_18864,N_19307);
or U19735 (N_19735,N_18835,N_18890);
nor U19736 (N_19736,N_19010,N_19229);
or U19737 (N_19737,N_19199,N_18892);
nor U19738 (N_19738,N_19034,N_19093);
nor U19739 (N_19739,N_19167,N_18925);
xor U19740 (N_19740,N_19345,N_19339);
nor U19741 (N_19741,N_19330,N_19172);
nand U19742 (N_19742,N_19001,N_18806);
nand U19743 (N_19743,N_18831,N_19107);
nor U19744 (N_19744,N_18752,N_19055);
and U19745 (N_19745,N_18810,N_18786);
nand U19746 (N_19746,N_18852,N_18821);
nor U19747 (N_19747,N_18933,N_18982);
nand U19748 (N_19748,N_19198,N_18760);
xnor U19749 (N_19749,N_19019,N_18865);
xor U19750 (N_19750,N_19317,N_18771);
and U19751 (N_19751,N_19112,N_19103);
and U19752 (N_19752,N_18967,N_19358);
or U19753 (N_19753,N_18838,N_18833);
xnor U19754 (N_19754,N_18859,N_18896);
and U19755 (N_19755,N_19163,N_19317);
and U19756 (N_19756,N_19145,N_19155);
or U19757 (N_19757,N_18906,N_18979);
nand U19758 (N_19758,N_18898,N_19217);
xor U19759 (N_19759,N_18877,N_19007);
or U19760 (N_19760,N_19371,N_19066);
xor U19761 (N_19761,N_19313,N_18845);
or U19762 (N_19762,N_19172,N_19178);
and U19763 (N_19763,N_18783,N_19030);
or U19764 (N_19764,N_18828,N_18770);
or U19765 (N_19765,N_19219,N_19140);
nand U19766 (N_19766,N_18773,N_18949);
nor U19767 (N_19767,N_19337,N_19270);
nor U19768 (N_19768,N_18807,N_19177);
nand U19769 (N_19769,N_19004,N_19064);
or U19770 (N_19770,N_19200,N_19219);
or U19771 (N_19771,N_18998,N_18814);
nand U19772 (N_19772,N_19005,N_19313);
xnor U19773 (N_19773,N_19343,N_19096);
or U19774 (N_19774,N_18764,N_18854);
and U19775 (N_19775,N_18767,N_18789);
nand U19776 (N_19776,N_19192,N_18947);
xnor U19777 (N_19777,N_18830,N_19085);
or U19778 (N_19778,N_19256,N_19371);
xor U19779 (N_19779,N_19281,N_19010);
nand U19780 (N_19780,N_19358,N_19310);
nor U19781 (N_19781,N_18847,N_18955);
nor U19782 (N_19782,N_18880,N_19169);
or U19783 (N_19783,N_19361,N_18855);
nor U19784 (N_19784,N_19327,N_18957);
or U19785 (N_19785,N_19013,N_19275);
or U19786 (N_19786,N_19163,N_19060);
nor U19787 (N_19787,N_18785,N_19269);
nand U19788 (N_19788,N_18950,N_18892);
and U19789 (N_19789,N_19032,N_19218);
nor U19790 (N_19790,N_18813,N_18972);
or U19791 (N_19791,N_19344,N_19268);
and U19792 (N_19792,N_18835,N_19090);
or U19793 (N_19793,N_18876,N_18966);
nor U19794 (N_19794,N_19150,N_18882);
nor U19795 (N_19795,N_18759,N_18979);
xnor U19796 (N_19796,N_19165,N_19295);
or U19797 (N_19797,N_19213,N_18973);
nor U19798 (N_19798,N_18854,N_19163);
nand U19799 (N_19799,N_19301,N_19082);
nand U19800 (N_19800,N_19172,N_19040);
nor U19801 (N_19801,N_19208,N_19094);
nor U19802 (N_19802,N_18927,N_19067);
xnor U19803 (N_19803,N_19142,N_19288);
nor U19804 (N_19804,N_19006,N_19005);
or U19805 (N_19805,N_18883,N_19321);
or U19806 (N_19806,N_19079,N_18838);
or U19807 (N_19807,N_19158,N_19050);
and U19808 (N_19808,N_18814,N_18804);
xor U19809 (N_19809,N_19350,N_19122);
xnor U19810 (N_19810,N_19271,N_18837);
xor U19811 (N_19811,N_19230,N_19288);
xnor U19812 (N_19812,N_19024,N_19257);
nand U19813 (N_19813,N_19359,N_18940);
nand U19814 (N_19814,N_19325,N_19311);
xor U19815 (N_19815,N_18998,N_19303);
or U19816 (N_19816,N_18765,N_18970);
nand U19817 (N_19817,N_18929,N_19359);
xnor U19818 (N_19818,N_19081,N_18812);
and U19819 (N_19819,N_18995,N_18881);
xor U19820 (N_19820,N_18771,N_18939);
nor U19821 (N_19821,N_19034,N_19323);
and U19822 (N_19822,N_18754,N_19286);
or U19823 (N_19823,N_19134,N_19168);
or U19824 (N_19824,N_18784,N_19187);
and U19825 (N_19825,N_19311,N_18824);
xor U19826 (N_19826,N_18951,N_18772);
nand U19827 (N_19827,N_18891,N_19244);
or U19828 (N_19828,N_19129,N_19257);
xor U19829 (N_19829,N_19171,N_19204);
nor U19830 (N_19830,N_19148,N_18987);
nor U19831 (N_19831,N_18818,N_19362);
nand U19832 (N_19832,N_19283,N_19193);
xor U19833 (N_19833,N_19206,N_18889);
nand U19834 (N_19834,N_19189,N_18794);
xnor U19835 (N_19835,N_19115,N_19324);
or U19836 (N_19836,N_19092,N_18854);
and U19837 (N_19837,N_19120,N_18933);
and U19838 (N_19838,N_18853,N_19368);
and U19839 (N_19839,N_19013,N_19272);
xor U19840 (N_19840,N_19006,N_18784);
and U19841 (N_19841,N_18779,N_19173);
nand U19842 (N_19842,N_18957,N_19335);
xor U19843 (N_19843,N_19244,N_18789);
xor U19844 (N_19844,N_18846,N_19058);
nand U19845 (N_19845,N_19299,N_18832);
nand U19846 (N_19846,N_19351,N_18855);
nand U19847 (N_19847,N_19174,N_19344);
xor U19848 (N_19848,N_19323,N_18935);
or U19849 (N_19849,N_18789,N_19147);
and U19850 (N_19850,N_19155,N_19168);
nand U19851 (N_19851,N_18890,N_19104);
or U19852 (N_19852,N_19077,N_19092);
xor U19853 (N_19853,N_19301,N_18759);
and U19854 (N_19854,N_19373,N_19226);
nand U19855 (N_19855,N_19052,N_19345);
xnor U19856 (N_19856,N_19125,N_19234);
nor U19857 (N_19857,N_19082,N_19192);
and U19858 (N_19858,N_19292,N_19037);
nand U19859 (N_19859,N_18958,N_19368);
or U19860 (N_19860,N_19024,N_19013);
and U19861 (N_19861,N_18912,N_19240);
and U19862 (N_19862,N_18773,N_19080);
and U19863 (N_19863,N_18846,N_19310);
nand U19864 (N_19864,N_19318,N_18806);
and U19865 (N_19865,N_19175,N_18849);
xnor U19866 (N_19866,N_18936,N_19093);
and U19867 (N_19867,N_19365,N_19177);
nor U19868 (N_19868,N_19238,N_18903);
nand U19869 (N_19869,N_18994,N_19031);
nand U19870 (N_19870,N_19340,N_18789);
or U19871 (N_19871,N_18751,N_19076);
nand U19872 (N_19872,N_19150,N_19205);
nand U19873 (N_19873,N_18815,N_18954);
xnor U19874 (N_19874,N_18867,N_19175);
xnor U19875 (N_19875,N_18827,N_19167);
or U19876 (N_19876,N_19077,N_19299);
nand U19877 (N_19877,N_18922,N_19006);
nand U19878 (N_19878,N_18937,N_19309);
nor U19879 (N_19879,N_19211,N_18827);
nor U19880 (N_19880,N_18918,N_19145);
nor U19881 (N_19881,N_19233,N_19215);
xor U19882 (N_19882,N_19153,N_19182);
or U19883 (N_19883,N_19066,N_19191);
nand U19884 (N_19884,N_19123,N_19273);
nand U19885 (N_19885,N_19027,N_19020);
nor U19886 (N_19886,N_19281,N_19200);
nor U19887 (N_19887,N_19344,N_18996);
xnor U19888 (N_19888,N_19007,N_18948);
or U19889 (N_19889,N_19093,N_18886);
and U19890 (N_19890,N_19231,N_18795);
nor U19891 (N_19891,N_19172,N_19004);
and U19892 (N_19892,N_19095,N_19274);
nand U19893 (N_19893,N_19053,N_19347);
nor U19894 (N_19894,N_18772,N_19069);
nand U19895 (N_19895,N_19068,N_19207);
and U19896 (N_19896,N_18783,N_18968);
xnor U19897 (N_19897,N_18798,N_19273);
nand U19898 (N_19898,N_18763,N_19296);
nand U19899 (N_19899,N_18847,N_18901);
and U19900 (N_19900,N_18951,N_18903);
nand U19901 (N_19901,N_19084,N_19019);
nand U19902 (N_19902,N_18777,N_19274);
nor U19903 (N_19903,N_19153,N_19097);
or U19904 (N_19904,N_19059,N_19137);
or U19905 (N_19905,N_18930,N_19256);
xnor U19906 (N_19906,N_19357,N_19335);
nor U19907 (N_19907,N_19283,N_19041);
nor U19908 (N_19908,N_19253,N_18952);
and U19909 (N_19909,N_19250,N_18792);
and U19910 (N_19910,N_19132,N_19066);
xor U19911 (N_19911,N_18984,N_18752);
or U19912 (N_19912,N_19179,N_19214);
xnor U19913 (N_19913,N_19225,N_19363);
nor U19914 (N_19914,N_18880,N_19277);
nand U19915 (N_19915,N_19183,N_19370);
or U19916 (N_19916,N_19309,N_18986);
nor U19917 (N_19917,N_18774,N_19280);
and U19918 (N_19918,N_19198,N_19102);
nor U19919 (N_19919,N_19262,N_19189);
nor U19920 (N_19920,N_19097,N_19166);
nand U19921 (N_19921,N_18880,N_18961);
and U19922 (N_19922,N_19013,N_19327);
xnor U19923 (N_19923,N_18855,N_19347);
nand U19924 (N_19924,N_18911,N_19265);
nand U19925 (N_19925,N_19282,N_19062);
and U19926 (N_19926,N_18948,N_19342);
xor U19927 (N_19927,N_19139,N_18887);
or U19928 (N_19928,N_18966,N_18854);
nand U19929 (N_19929,N_18805,N_18994);
nand U19930 (N_19930,N_19275,N_18785);
nor U19931 (N_19931,N_19230,N_19016);
and U19932 (N_19932,N_18896,N_19033);
xor U19933 (N_19933,N_18985,N_19228);
nor U19934 (N_19934,N_18966,N_18929);
and U19935 (N_19935,N_18865,N_18764);
or U19936 (N_19936,N_19368,N_19072);
nand U19937 (N_19937,N_19070,N_19018);
nor U19938 (N_19938,N_19357,N_18923);
and U19939 (N_19939,N_18953,N_19112);
or U19940 (N_19940,N_19156,N_18800);
xnor U19941 (N_19941,N_18839,N_18873);
and U19942 (N_19942,N_18801,N_19110);
or U19943 (N_19943,N_19017,N_18854);
and U19944 (N_19944,N_18929,N_19373);
nor U19945 (N_19945,N_18812,N_19166);
and U19946 (N_19946,N_19238,N_19078);
nand U19947 (N_19947,N_18825,N_18920);
or U19948 (N_19948,N_18790,N_18874);
and U19949 (N_19949,N_18870,N_18866);
xor U19950 (N_19950,N_19365,N_18833);
xor U19951 (N_19951,N_19025,N_19330);
nor U19952 (N_19952,N_19227,N_19305);
xnor U19953 (N_19953,N_19331,N_18881);
or U19954 (N_19954,N_19236,N_19006);
xnor U19955 (N_19955,N_19117,N_19315);
nor U19956 (N_19956,N_18946,N_19250);
xnor U19957 (N_19957,N_19304,N_18959);
xor U19958 (N_19958,N_19281,N_18979);
or U19959 (N_19959,N_18756,N_18837);
or U19960 (N_19960,N_19303,N_19004);
nor U19961 (N_19961,N_18971,N_18899);
xnor U19962 (N_19962,N_18763,N_19332);
or U19963 (N_19963,N_18891,N_18915);
and U19964 (N_19964,N_19165,N_19292);
xor U19965 (N_19965,N_18877,N_18950);
xor U19966 (N_19966,N_18942,N_19107);
nand U19967 (N_19967,N_18982,N_18919);
nand U19968 (N_19968,N_19348,N_18991);
xnor U19969 (N_19969,N_18768,N_19111);
or U19970 (N_19970,N_18985,N_18793);
nor U19971 (N_19971,N_19221,N_19138);
nor U19972 (N_19972,N_19368,N_19052);
and U19973 (N_19973,N_18759,N_19064);
xnor U19974 (N_19974,N_19368,N_18874);
xnor U19975 (N_19975,N_19367,N_19329);
xor U19976 (N_19976,N_18820,N_18784);
nand U19977 (N_19977,N_18911,N_19201);
nor U19978 (N_19978,N_18883,N_18924);
xor U19979 (N_19979,N_18952,N_19349);
xnor U19980 (N_19980,N_19183,N_19107);
or U19981 (N_19981,N_19206,N_19089);
nand U19982 (N_19982,N_19374,N_18779);
nor U19983 (N_19983,N_19265,N_19069);
nor U19984 (N_19984,N_19133,N_18947);
or U19985 (N_19985,N_19185,N_18992);
or U19986 (N_19986,N_19241,N_18885);
and U19987 (N_19987,N_19226,N_19138);
xor U19988 (N_19988,N_19078,N_19073);
nor U19989 (N_19989,N_19224,N_19250);
nand U19990 (N_19990,N_18977,N_19351);
or U19991 (N_19991,N_19003,N_19105);
xnor U19992 (N_19992,N_19371,N_19042);
and U19993 (N_19993,N_18755,N_18945);
nand U19994 (N_19994,N_19069,N_19236);
nor U19995 (N_19995,N_18866,N_19094);
nor U19996 (N_19996,N_19224,N_18940);
nand U19997 (N_19997,N_18800,N_19264);
xnor U19998 (N_19998,N_18936,N_18928);
nand U19999 (N_19999,N_19282,N_19274);
or U20000 (N_20000,N_19844,N_19820);
nand U20001 (N_20001,N_19647,N_19639);
or U20002 (N_20002,N_19990,N_19825);
and U20003 (N_20003,N_19695,N_19493);
nand U20004 (N_20004,N_19551,N_19710);
and U20005 (N_20005,N_19883,N_19386);
and U20006 (N_20006,N_19747,N_19524);
and U20007 (N_20007,N_19583,N_19866);
xnor U20008 (N_20008,N_19927,N_19575);
nor U20009 (N_20009,N_19724,N_19542);
nand U20010 (N_20010,N_19599,N_19926);
nand U20011 (N_20011,N_19988,N_19787);
nor U20012 (N_20012,N_19512,N_19955);
nor U20013 (N_20013,N_19431,N_19778);
xor U20014 (N_20014,N_19970,N_19548);
nor U20015 (N_20015,N_19401,N_19856);
and U20016 (N_20016,N_19488,N_19385);
xnor U20017 (N_20017,N_19454,N_19879);
xnor U20018 (N_20018,N_19411,N_19703);
nand U20019 (N_20019,N_19752,N_19499);
nand U20020 (N_20020,N_19800,N_19887);
nand U20021 (N_20021,N_19419,N_19545);
xnor U20022 (N_20022,N_19643,N_19992);
nor U20023 (N_20023,N_19514,N_19464);
or U20024 (N_20024,N_19562,N_19607);
and U20025 (N_20025,N_19918,N_19427);
nor U20026 (N_20026,N_19793,N_19726);
nand U20027 (N_20027,N_19693,N_19819);
nor U20028 (N_20028,N_19953,N_19447);
xnor U20029 (N_20029,N_19899,N_19977);
nand U20030 (N_20030,N_19855,N_19680);
nand U20031 (N_20031,N_19826,N_19640);
xor U20032 (N_20032,N_19500,N_19396);
xor U20033 (N_20033,N_19596,N_19413);
or U20034 (N_20034,N_19768,N_19730);
nand U20035 (N_20035,N_19457,N_19487);
or U20036 (N_20036,N_19719,N_19389);
or U20037 (N_20037,N_19400,N_19506);
xor U20038 (N_20038,N_19571,N_19723);
xor U20039 (N_20039,N_19763,N_19445);
xor U20040 (N_20040,N_19424,N_19520);
and U20041 (N_20041,N_19980,N_19534);
or U20042 (N_20042,N_19472,N_19452);
xnor U20043 (N_20043,N_19983,N_19789);
nor U20044 (N_20044,N_19982,N_19409);
xnor U20045 (N_20045,N_19868,N_19631);
xor U20046 (N_20046,N_19378,N_19909);
xnor U20047 (N_20047,N_19377,N_19957);
nand U20048 (N_20048,N_19662,N_19854);
nor U20049 (N_20049,N_19381,N_19456);
nand U20050 (N_20050,N_19432,N_19753);
and U20051 (N_20051,N_19830,N_19679);
nand U20052 (N_20052,N_19558,N_19960);
nor U20053 (N_20053,N_19886,N_19717);
xnor U20054 (N_20054,N_19942,N_19857);
nor U20055 (N_20055,N_19503,N_19928);
and U20056 (N_20056,N_19792,N_19589);
nand U20057 (N_20057,N_19627,N_19523);
and U20058 (N_20058,N_19473,N_19847);
or U20059 (N_20059,N_19751,N_19897);
and U20060 (N_20060,N_19564,N_19686);
xor U20061 (N_20061,N_19766,N_19754);
xor U20062 (N_20062,N_19528,N_19803);
nor U20063 (N_20063,N_19496,N_19463);
xnor U20064 (N_20064,N_19905,N_19991);
and U20065 (N_20065,N_19430,N_19568);
or U20066 (N_20066,N_19544,N_19872);
xnor U20067 (N_20067,N_19739,N_19654);
xnor U20068 (N_20068,N_19943,N_19848);
nor U20069 (N_20069,N_19834,N_19837);
xnor U20070 (N_20070,N_19592,N_19870);
nor U20071 (N_20071,N_19467,N_19637);
nor U20072 (N_20072,N_19458,N_19880);
and U20073 (N_20073,N_19881,N_19549);
nor U20074 (N_20074,N_19774,N_19698);
nor U20075 (N_20075,N_19835,N_19963);
nand U20076 (N_20076,N_19407,N_19900);
nand U20077 (N_20077,N_19522,N_19961);
nand U20078 (N_20078,N_19418,N_19944);
nand U20079 (N_20079,N_19938,N_19644);
xnor U20080 (N_20080,N_19972,N_19921);
xnor U20081 (N_20081,N_19814,N_19746);
or U20082 (N_20082,N_19605,N_19843);
xnor U20083 (N_20083,N_19392,N_19838);
xor U20084 (N_20084,N_19799,N_19441);
xnor U20085 (N_20085,N_19553,N_19380);
xor U20086 (N_20086,N_19450,N_19901);
nand U20087 (N_20087,N_19517,N_19593);
or U20088 (N_20088,N_19600,N_19451);
nor U20089 (N_20089,N_19875,N_19440);
nor U20090 (N_20090,N_19770,N_19586);
nand U20091 (N_20091,N_19635,N_19802);
nand U20092 (N_20092,N_19994,N_19869);
or U20093 (N_20093,N_19507,N_19925);
or U20094 (N_20094,N_19779,N_19864);
nor U20095 (N_20095,N_19560,N_19630);
or U20096 (N_20096,N_19391,N_19606);
nand U20097 (N_20097,N_19767,N_19794);
xor U20098 (N_20098,N_19669,N_19860);
nand U20099 (N_20099,N_19394,N_19891);
nand U20100 (N_20100,N_19948,N_19771);
nor U20101 (N_20101,N_19438,N_19602);
nor U20102 (N_20102,N_19581,N_19998);
or U20103 (N_20103,N_19813,N_19632);
and U20104 (N_20104,N_19516,N_19713);
nor U20105 (N_20105,N_19384,N_19665);
nand U20106 (N_20106,N_19975,N_19812);
or U20107 (N_20107,N_19859,N_19995);
nand U20108 (N_20108,N_19483,N_19999);
nand U20109 (N_20109,N_19976,N_19591);
nor U20110 (N_20110,N_19375,N_19660);
xor U20111 (N_20111,N_19379,N_19540);
xor U20112 (N_20112,N_19444,N_19688);
xor U20113 (N_20113,N_19687,N_19700);
and U20114 (N_20114,N_19478,N_19397);
or U20115 (N_20115,N_19922,N_19408);
nand U20116 (N_20116,N_19421,N_19645);
or U20117 (N_20117,N_19762,N_19930);
or U20118 (N_20118,N_19704,N_19505);
or U20119 (N_20119,N_19395,N_19436);
nand U20120 (N_20120,N_19890,N_19462);
xnor U20121 (N_20121,N_19615,N_19967);
or U20122 (N_20122,N_19797,N_19584);
or U20123 (N_20123,N_19657,N_19941);
nand U20124 (N_20124,N_19557,N_19477);
or U20125 (N_20125,N_19958,N_19946);
xnor U20126 (N_20126,N_19543,N_19978);
nand U20127 (N_20127,N_19788,N_19468);
nor U20128 (N_20128,N_19775,N_19617);
nor U20129 (N_20129,N_19908,N_19486);
nand U20130 (N_20130,N_19613,N_19780);
or U20131 (N_20131,N_19561,N_19707);
nand U20132 (N_20132,N_19822,N_19737);
nor U20133 (N_20133,N_19484,N_19842);
nor U20134 (N_20134,N_19845,N_19810);
xor U20135 (N_20135,N_19933,N_19877);
or U20136 (N_20136,N_19674,N_19715);
and U20137 (N_20137,N_19410,N_19388);
nor U20138 (N_20138,N_19935,N_19986);
nand U20139 (N_20139,N_19659,N_19449);
and U20140 (N_20140,N_19728,N_19885);
or U20141 (N_20141,N_19656,N_19910);
nor U20142 (N_20142,N_19422,N_19936);
nand U20143 (N_20143,N_19965,N_19572);
or U20144 (N_20144,N_19609,N_19677);
or U20145 (N_20145,N_19858,N_19460);
xor U20146 (N_20146,N_19750,N_19588);
and U20147 (N_20147,N_19603,N_19634);
nor U20148 (N_20148,N_19650,N_19711);
nand U20149 (N_20149,N_19547,N_19433);
or U20150 (N_20150,N_19849,N_19578);
xnor U20151 (N_20151,N_19809,N_19479);
or U20152 (N_20152,N_19954,N_19823);
nor U20153 (N_20153,N_19696,N_19896);
and U20154 (N_20154,N_19989,N_19985);
xnor U20155 (N_20155,N_19741,N_19511);
nand U20156 (N_20156,N_19783,N_19790);
and U20157 (N_20157,N_19757,N_19390);
xor U20158 (N_20158,N_19490,N_19836);
nor U20159 (N_20159,N_19818,N_19435);
nor U20160 (N_20160,N_19601,N_19673);
nor U20161 (N_20161,N_19996,N_19405);
or U20162 (N_20162,N_19567,N_19807);
or U20163 (N_20163,N_19608,N_19668);
nor U20164 (N_20164,N_19889,N_19971);
nor U20165 (N_20165,N_19555,N_19867);
and U20166 (N_20166,N_19618,N_19882);
nand U20167 (N_20167,N_19876,N_19956);
nor U20168 (N_20168,N_19716,N_19945);
xor U20169 (N_20169,N_19725,N_19756);
or U20170 (N_20170,N_19667,N_19485);
nand U20171 (N_20171,N_19937,N_19539);
and U20172 (N_20172,N_19808,N_19939);
nand U20173 (N_20173,N_19626,N_19940);
xnor U20174 (N_20174,N_19689,N_19559);
nand U20175 (N_20175,N_19697,N_19777);
and U20176 (N_20176,N_19556,N_19832);
or U20177 (N_20177,N_19769,N_19437);
nand U20178 (N_20178,N_19376,N_19573);
and U20179 (N_20179,N_19442,N_19641);
nand U20180 (N_20180,N_19898,N_19504);
nor U20181 (N_20181,N_19453,N_19736);
xnor U20182 (N_20182,N_19519,N_19611);
nor U20183 (N_20183,N_19681,N_19892);
xnor U20184 (N_20184,N_19469,N_19675);
or U20185 (N_20185,N_19932,N_19466);
nor U20186 (N_20186,N_19950,N_19840);
nand U20187 (N_20187,N_19651,N_19692);
or U20188 (N_20188,N_19587,N_19633);
nand U20189 (N_20189,N_19476,N_19624);
xnor U20190 (N_20190,N_19598,N_19904);
nor U20191 (N_20191,N_19597,N_19805);
xnor U20192 (N_20192,N_19722,N_19744);
nor U20193 (N_20193,N_19806,N_19629);
and U20194 (N_20194,N_19964,N_19538);
or U20195 (N_20195,N_19612,N_19829);
nor U20196 (N_20196,N_19745,N_19984);
nand U20197 (N_20197,N_19798,N_19917);
xnor U20198 (N_20198,N_19906,N_19495);
and U20199 (N_20199,N_19663,N_19729);
nor U20200 (N_20200,N_19748,N_19404);
nand U20201 (N_20201,N_19535,N_19853);
nand U20202 (N_20202,N_19833,N_19434);
xor U20203 (N_20203,N_19417,N_19852);
xnor U20204 (N_20204,N_19920,N_19947);
nor U20205 (N_20205,N_19480,N_19590);
nand U20206 (N_20206,N_19796,N_19530);
xor U20207 (N_20207,N_19694,N_19570);
and U20208 (N_20208,N_19907,N_19742);
and U20209 (N_20209,N_19727,N_19552);
and U20210 (N_20210,N_19509,N_19678);
nor U20211 (N_20211,N_19721,N_19732);
xor U20212 (N_20212,N_19655,N_19865);
or U20213 (N_20213,N_19894,N_19585);
and U20214 (N_20214,N_19448,N_19474);
nand U20215 (N_20215,N_19735,N_19546);
nor U20216 (N_20216,N_19594,N_19811);
nand U20217 (N_20217,N_19387,N_19903);
xor U20218 (N_20218,N_19893,N_19861);
or U20219 (N_20219,N_19577,N_19670);
or U20220 (N_20220,N_19653,N_19664);
nor U20221 (N_20221,N_19383,N_19816);
and U20222 (N_20222,N_19979,N_19574);
xnor U20223 (N_20223,N_19428,N_19621);
xor U20224 (N_20224,N_19974,N_19489);
xor U20225 (N_20225,N_19515,N_19821);
and U20226 (N_20226,N_19781,N_19661);
or U20227 (N_20227,N_19582,N_19525);
and U20228 (N_20228,N_19720,N_19702);
xor U20229 (N_20229,N_19772,N_19537);
or U20230 (N_20230,N_19649,N_19828);
or U20231 (N_20231,N_19862,N_19863);
nor U20232 (N_20232,N_19443,N_19705);
nor U20233 (N_20233,N_19446,N_19393);
or U20234 (N_20234,N_19931,N_19526);
nand U20235 (N_20235,N_19824,N_19563);
nor U20236 (N_20236,N_19439,N_19682);
xor U20237 (N_20237,N_19878,N_19536);
xor U20238 (N_20238,N_19981,N_19492);
nor U20239 (N_20239,N_19403,N_19733);
or U20240 (N_20240,N_19973,N_19416);
or U20241 (N_20241,N_19912,N_19646);
or U20242 (N_20242,N_19471,N_19773);
nand U20243 (N_20243,N_19642,N_19420);
and U20244 (N_20244,N_19614,N_19951);
xor U20245 (N_20245,N_19871,N_19671);
nor U20246 (N_20246,N_19414,N_19786);
nand U20247 (N_20247,N_19801,N_19482);
nor U20248 (N_20248,N_19541,N_19412);
nor U20249 (N_20249,N_19902,N_19652);
or U20250 (N_20250,N_19791,N_19884);
nand U20251 (N_20251,N_19565,N_19576);
nand U20252 (N_20252,N_19580,N_19740);
nor U20253 (N_20253,N_19616,N_19683);
nand U20254 (N_20254,N_19815,N_19648);
or U20255 (N_20255,N_19604,N_19949);
and U20256 (N_20256,N_19784,N_19758);
or U20257 (N_20257,N_19888,N_19491);
nand U20258 (N_20258,N_19966,N_19731);
and U20259 (N_20259,N_19481,N_19636);
xnor U20260 (N_20260,N_19494,N_19708);
nand U20261 (N_20261,N_19610,N_19382);
and U20262 (N_20262,N_19851,N_19399);
nand U20263 (N_20263,N_19817,N_19701);
and U20264 (N_20264,N_19415,N_19513);
xnor U20265 (N_20265,N_19685,N_19827);
nor U20266 (N_20266,N_19398,N_19924);
xnor U20267 (N_20267,N_19738,N_19423);
xnor U20268 (N_20268,N_19923,N_19426);
and U20269 (N_20269,N_19993,N_19841);
and U20270 (N_20270,N_19531,N_19501);
xor U20271 (N_20271,N_19529,N_19914);
nand U20272 (N_20272,N_19690,N_19795);
or U20273 (N_20273,N_19839,N_19402);
and U20274 (N_20274,N_19622,N_19913);
or U20275 (N_20275,N_19497,N_19658);
and U20276 (N_20276,N_19508,N_19962);
nor U20277 (N_20277,N_19846,N_19804);
or U20278 (N_20278,N_19997,N_19566);
or U20279 (N_20279,N_19969,N_19510);
nor U20280 (N_20280,N_19595,N_19734);
nand U20281 (N_20281,N_19952,N_19625);
and U20282 (N_20282,N_19850,N_19579);
or U20283 (N_20283,N_19470,N_19718);
nand U20284 (N_20284,N_19706,N_19498);
xor U20285 (N_20285,N_19455,N_19628);
xnor U20286 (N_20286,N_19915,N_19776);
xnor U20287 (N_20287,N_19968,N_19874);
xnor U20288 (N_20288,N_19521,N_19672);
or U20289 (N_20289,N_19765,N_19919);
nand U20290 (N_20290,N_19465,N_19533);
and U20291 (N_20291,N_19475,N_19623);
nand U20292 (N_20292,N_19502,N_19684);
or U20293 (N_20293,N_19873,N_19461);
nor U20294 (N_20294,N_19911,N_19785);
xor U20295 (N_20295,N_19638,N_19550);
nor U20296 (N_20296,N_19699,N_19764);
nor U20297 (N_20297,N_19712,N_19691);
nor U20298 (N_20298,N_19709,N_19676);
or U20299 (N_20299,N_19743,N_19934);
and U20300 (N_20300,N_19761,N_19569);
nor U20301 (N_20301,N_19987,N_19759);
nand U20302 (N_20302,N_19532,N_19619);
nand U20303 (N_20303,N_19760,N_19749);
or U20304 (N_20304,N_19666,N_19959);
nand U20305 (N_20305,N_19429,N_19831);
nand U20306 (N_20306,N_19916,N_19518);
nor U20307 (N_20307,N_19895,N_19929);
nand U20308 (N_20308,N_19714,N_19459);
or U20309 (N_20309,N_19406,N_19527);
or U20310 (N_20310,N_19755,N_19620);
and U20311 (N_20311,N_19554,N_19782);
or U20312 (N_20312,N_19425,N_19636);
or U20313 (N_20313,N_19706,N_19977);
xor U20314 (N_20314,N_19950,N_19390);
and U20315 (N_20315,N_19407,N_19887);
nor U20316 (N_20316,N_19837,N_19498);
nand U20317 (N_20317,N_19399,N_19765);
and U20318 (N_20318,N_19868,N_19376);
xnor U20319 (N_20319,N_19660,N_19725);
nor U20320 (N_20320,N_19750,N_19910);
and U20321 (N_20321,N_19642,N_19662);
nor U20322 (N_20322,N_19503,N_19579);
nand U20323 (N_20323,N_19752,N_19725);
and U20324 (N_20324,N_19411,N_19665);
or U20325 (N_20325,N_19509,N_19428);
or U20326 (N_20326,N_19442,N_19843);
xor U20327 (N_20327,N_19575,N_19588);
nor U20328 (N_20328,N_19409,N_19389);
nor U20329 (N_20329,N_19775,N_19934);
xor U20330 (N_20330,N_19831,N_19514);
or U20331 (N_20331,N_19568,N_19404);
nor U20332 (N_20332,N_19628,N_19778);
and U20333 (N_20333,N_19604,N_19844);
or U20334 (N_20334,N_19995,N_19551);
nor U20335 (N_20335,N_19573,N_19815);
and U20336 (N_20336,N_19686,N_19445);
nand U20337 (N_20337,N_19385,N_19576);
and U20338 (N_20338,N_19677,N_19516);
or U20339 (N_20339,N_19643,N_19490);
and U20340 (N_20340,N_19850,N_19448);
nor U20341 (N_20341,N_19629,N_19983);
nor U20342 (N_20342,N_19915,N_19639);
nor U20343 (N_20343,N_19412,N_19675);
xnor U20344 (N_20344,N_19545,N_19913);
nand U20345 (N_20345,N_19932,N_19519);
and U20346 (N_20346,N_19444,N_19459);
xnor U20347 (N_20347,N_19870,N_19532);
xor U20348 (N_20348,N_19600,N_19485);
nand U20349 (N_20349,N_19476,N_19927);
nand U20350 (N_20350,N_19651,N_19390);
xnor U20351 (N_20351,N_19745,N_19626);
or U20352 (N_20352,N_19819,N_19846);
and U20353 (N_20353,N_19664,N_19796);
or U20354 (N_20354,N_19660,N_19526);
and U20355 (N_20355,N_19802,N_19985);
nor U20356 (N_20356,N_19455,N_19521);
nand U20357 (N_20357,N_19629,N_19685);
xor U20358 (N_20358,N_19814,N_19951);
xnor U20359 (N_20359,N_19956,N_19672);
or U20360 (N_20360,N_19866,N_19689);
or U20361 (N_20361,N_19508,N_19736);
or U20362 (N_20362,N_19879,N_19984);
or U20363 (N_20363,N_19809,N_19922);
nand U20364 (N_20364,N_19765,N_19909);
nor U20365 (N_20365,N_19821,N_19906);
nand U20366 (N_20366,N_19995,N_19837);
xor U20367 (N_20367,N_19604,N_19674);
and U20368 (N_20368,N_19427,N_19947);
xor U20369 (N_20369,N_19998,N_19611);
nand U20370 (N_20370,N_19958,N_19533);
and U20371 (N_20371,N_19571,N_19846);
and U20372 (N_20372,N_19817,N_19517);
nor U20373 (N_20373,N_19517,N_19932);
nor U20374 (N_20374,N_19983,N_19952);
xnor U20375 (N_20375,N_19428,N_19978);
nand U20376 (N_20376,N_19892,N_19878);
nor U20377 (N_20377,N_19477,N_19710);
nand U20378 (N_20378,N_19388,N_19942);
or U20379 (N_20379,N_19974,N_19855);
and U20380 (N_20380,N_19945,N_19923);
nand U20381 (N_20381,N_19992,N_19856);
or U20382 (N_20382,N_19886,N_19601);
nor U20383 (N_20383,N_19761,N_19676);
or U20384 (N_20384,N_19830,N_19552);
nor U20385 (N_20385,N_19483,N_19723);
nand U20386 (N_20386,N_19532,N_19460);
and U20387 (N_20387,N_19409,N_19468);
nand U20388 (N_20388,N_19933,N_19859);
and U20389 (N_20389,N_19650,N_19752);
nand U20390 (N_20390,N_19743,N_19449);
or U20391 (N_20391,N_19491,N_19872);
xor U20392 (N_20392,N_19403,N_19538);
nand U20393 (N_20393,N_19961,N_19999);
nand U20394 (N_20394,N_19960,N_19962);
or U20395 (N_20395,N_19805,N_19550);
and U20396 (N_20396,N_19422,N_19718);
xor U20397 (N_20397,N_19917,N_19665);
and U20398 (N_20398,N_19938,N_19955);
nand U20399 (N_20399,N_19787,N_19927);
nor U20400 (N_20400,N_19939,N_19906);
nor U20401 (N_20401,N_19505,N_19518);
or U20402 (N_20402,N_19553,N_19843);
or U20403 (N_20403,N_19710,N_19683);
xor U20404 (N_20404,N_19611,N_19595);
or U20405 (N_20405,N_19480,N_19861);
xnor U20406 (N_20406,N_19899,N_19639);
nand U20407 (N_20407,N_19549,N_19846);
nor U20408 (N_20408,N_19896,N_19760);
or U20409 (N_20409,N_19473,N_19753);
xnor U20410 (N_20410,N_19714,N_19998);
and U20411 (N_20411,N_19463,N_19510);
or U20412 (N_20412,N_19470,N_19949);
xnor U20413 (N_20413,N_19972,N_19956);
and U20414 (N_20414,N_19697,N_19496);
nor U20415 (N_20415,N_19952,N_19724);
nand U20416 (N_20416,N_19700,N_19814);
nand U20417 (N_20417,N_19799,N_19941);
nand U20418 (N_20418,N_19450,N_19437);
nor U20419 (N_20419,N_19743,N_19724);
nor U20420 (N_20420,N_19727,N_19488);
xor U20421 (N_20421,N_19605,N_19690);
or U20422 (N_20422,N_19442,N_19887);
nand U20423 (N_20423,N_19597,N_19673);
and U20424 (N_20424,N_19586,N_19558);
nor U20425 (N_20425,N_19520,N_19411);
xnor U20426 (N_20426,N_19588,N_19724);
and U20427 (N_20427,N_19946,N_19957);
nand U20428 (N_20428,N_19487,N_19654);
xor U20429 (N_20429,N_19775,N_19869);
nand U20430 (N_20430,N_19460,N_19482);
nor U20431 (N_20431,N_19623,N_19649);
and U20432 (N_20432,N_19840,N_19784);
nand U20433 (N_20433,N_19707,N_19514);
xnor U20434 (N_20434,N_19706,N_19960);
and U20435 (N_20435,N_19761,N_19923);
xor U20436 (N_20436,N_19646,N_19627);
nor U20437 (N_20437,N_19744,N_19642);
nand U20438 (N_20438,N_19707,N_19742);
or U20439 (N_20439,N_19806,N_19650);
and U20440 (N_20440,N_19700,N_19598);
xnor U20441 (N_20441,N_19613,N_19652);
nand U20442 (N_20442,N_19908,N_19472);
or U20443 (N_20443,N_19441,N_19805);
and U20444 (N_20444,N_19961,N_19459);
or U20445 (N_20445,N_19456,N_19808);
and U20446 (N_20446,N_19798,N_19550);
and U20447 (N_20447,N_19819,N_19750);
nand U20448 (N_20448,N_19703,N_19641);
xnor U20449 (N_20449,N_19526,N_19909);
and U20450 (N_20450,N_19449,N_19486);
nand U20451 (N_20451,N_19654,N_19955);
or U20452 (N_20452,N_19510,N_19582);
nor U20453 (N_20453,N_19883,N_19639);
and U20454 (N_20454,N_19524,N_19640);
nor U20455 (N_20455,N_19776,N_19619);
and U20456 (N_20456,N_19794,N_19753);
nor U20457 (N_20457,N_19803,N_19795);
nand U20458 (N_20458,N_19525,N_19762);
nor U20459 (N_20459,N_19861,N_19676);
or U20460 (N_20460,N_19682,N_19619);
nand U20461 (N_20461,N_19578,N_19633);
xnor U20462 (N_20462,N_19412,N_19923);
nand U20463 (N_20463,N_19801,N_19839);
or U20464 (N_20464,N_19452,N_19710);
xor U20465 (N_20465,N_19856,N_19886);
xnor U20466 (N_20466,N_19680,N_19379);
or U20467 (N_20467,N_19537,N_19450);
nand U20468 (N_20468,N_19686,N_19377);
or U20469 (N_20469,N_19432,N_19454);
or U20470 (N_20470,N_19547,N_19531);
or U20471 (N_20471,N_19663,N_19938);
nand U20472 (N_20472,N_19721,N_19531);
or U20473 (N_20473,N_19466,N_19602);
xor U20474 (N_20474,N_19466,N_19908);
nand U20475 (N_20475,N_19803,N_19398);
and U20476 (N_20476,N_19446,N_19668);
or U20477 (N_20477,N_19414,N_19924);
nor U20478 (N_20478,N_19987,N_19857);
and U20479 (N_20479,N_19930,N_19392);
xnor U20480 (N_20480,N_19954,N_19617);
and U20481 (N_20481,N_19866,N_19499);
or U20482 (N_20482,N_19553,N_19437);
xor U20483 (N_20483,N_19709,N_19697);
and U20484 (N_20484,N_19630,N_19900);
nor U20485 (N_20485,N_19820,N_19931);
and U20486 (N_20486,N_19699,N_19645);
or U20487 (N_20487,N_19425,N_19504);
or U20488 (N_20488,N_19901,N_19950);
and U20489 (N_20489,N_19758,N_19819);
nand U20490 (N_20490,N_19959,N_19900);
and U20491 (N_20491,N_19481,N_19845);
nor U20492 (N_20492,N_19529,N_19763);
xnor U20493 (N_20493,N_19543,N_19607);
and U20494 (N_20494,N_19776,N_19640);
nand U20495 (N_20495,N_19807,N_19918);
or U20496 (N_20496,N_19810,N_19887);
nor U20497 (N_20497,N_19390,N_19481);
nor U20498 (N_20498,N_19854,N_19659);
nand U20499 (N_20499,N_19798,N_19983);
or U20500 (N_20500,N_19538,N_19757);
xnor U20501 (N_20501,N_19511,N_19958);
or U20502 (N_20502,N_19837,N_19635);
nor U20503 (N_20503,N_19615,N_19754);
nand U20504 (N_20504,N_19856,N_19642);
nor U20505 (N_20505,N_19720,N_19901);
xnor U20506 (N_20506,N_19873,N_19619);
or U20507 (N_20507,N_19375,N_19383);
nor U20508 (N_20508,N_19644,N_19779);
nand U20509 (N_20509,N_19536,N_19868);
and U20510 (N_20510,N_19921,N_19674);
or U20511 (N_20511,N_19719,N_19539);
or U20512 (N_20512,N_19636,N_19573);
nor U20513 (N_20513,N_19652,N_19453);
xnor U20514 (N_20514,N_19864,N_19916);
nand U20515 (N_20515,N_19498,N_19766);
and U20516 (N_20516,N_19426,N_19988);
and U20517 (N_20517,N_19844,N_19822);
or U20518 (N_20518,N_19563,N_19567);
nand U20519 (N_20519,N_19848,N_19415);
or U20520 (N_20520,N_19773,N_19535);
nand U20521 (N_20521,N_19426,N_19680);
xor U20522 (N_20522,N_19435,N_19606);
or U20523 (N_20523,N_19613,N_19411);
nand U20524 (N_20524,N_19827,N_19556);
nor U20525 (N_20525,N_19467,N_19411);
xor U20526 (N_20526,N_19795,N_19447);
nand U20527 (N_20527,N_19999,N_19438);
or U20528 (N_20528,N_19627,N_19848);
and U20529 (N_20529,N_19670,N_19689);
and U20530 (N_20530,N_19913,N_19659);
nor U20531 (N_20531,N_19844,N_19528);
xnor U20532 (N_20532,N_19599,N_19391);
or U20533 (N_20533,N_19435,N_19579);
and U20534 (N_20534,N_19459,N_19530);
nor U20535 (N_20535,N_19539,N_19403);
or U20536 (N_20536,N_19865,N_19408);
or U20537 (N_20537,N_19772,N_19732);
xnor U20538 (N_20538,N_19712,N_19876);
nor U20539 (N_20539,N_19669,N_19906);
xor U20540 (N_20540,N_19680,N_19730);
xnor U20541 (N_20541,N_19826,N_19440);
nor U20542 (N_20542,N_19981,N_19954);
xor U20543 (N_20543,N_19566,N_19708);
and U20544 (N_20544,N_19992,N_19436);
and U20545 (N_20545,N_19617,N_19848);
nand U20546 (N_20546,N_19385,N_19520);
nor U20547 (N_20547,N_19576,N_19407);
or U20548 (N_20548,N_19569,N_19425);
nand U20549 (N_20549,N_19493,N_19494);
and U20550 (N_20550,N_19964,N_19434);
or U20551 (N_20551,N_19820,N_19681);
nand U20552 (N_20552,N_19424,N_19702);
or U20553 (N_20553,N_19881,N_19964);
nand U20554 (N_20554,N_19916,N_19857);
or U20555 (N_20555,N_19592,N_19884);
xnor U20556 (N_20556,N_19705,N_19745);
or U20557 (N_20557,N_19760,N_19388);
nand U20558 (N_20558,N_19768,N_19637);
and U20559 (N_20559,N_19786,N_19743);
nor U20560 (N_20560,N_19390,N_19895);
nand U20561 (N_20561,N_19647,N_19494);
or U20562 (N_20562,N_19659,N_19439);
or U20563 (N_20563,N_19804,N_19808);
or U20564 (N_20564,N_19545,N_19750);
xnor U20565 (N_20565,N_19478,N_19535);
nand U20566 (N_20566,N_19462,N_19595);
or U20567 (N_20567,N_19392,N_19974);
nand U20568 (N_20568,N_19484,N_19542);
nand U20569 (N_20569,N_19671,N_19967);
or U20570 (N_20570,N_19721,N_19618);
and U20571 (N_20571,N_19635,N_19983);
and U20572 (N_20572,N_19546,N_19899);
or U20573 (N_20573,N_19785,N_19923);
nor U20574 (N_20574,N_19771,N_19881);
and U20575 (N_20575,N_19810,N_19415);
and U20576 (N_20576,N_19563,N_19957);
nor U20577 (N_20577,N_19949,N_19532);
or U20578 (N_20578,N_19402,N_19947);
nor U20579 (N_20579,N_19447,N_19507);
and U20580 (N_20580,N_19957,N_19999);
or U20581 (N_20581,N_19946,N_19467);
and U20582 (N_20582,N_19958,N_19805);
nand U20583 (N_20583,N_19415,N_19376);
nor U20584 (N_20584,N_19940,N_19864);
xor U20585 (N_20585,N_19756,N_19902);
xor U20586 (N_20586,N_19644,N_19398);
nand U20587 (N_20587,N_19581,N_19886);
or U20588 (N_20588,N_19623,N_19446);
nor U20589 (N_20589,N_19651,N_19558);
xnor U20590 (N_20590,N_19886,N_19720);
nand U20591 (N_20591,N_19557,N_19750);
nand U20592 (N_20592,N_19641,N_19644);
or U20593 (N_20593,N_19965,N_19517);
nor U20594 (N_20594,N_19462,N_19870);
nor U20595 (N_20595,N_19994,N_19420);
or U20596 (N_20596,N_19796,N_19784);
nor U20597 (N_20597,N_19524,N_19673);
and U20598 (N_20598,N_19674,N_19780);
or U20599 (N_20599,N_19677,N_19916);
and U20600 (N_20600,N_19965,N_19875);
nand U20601 (N_20601,N_19567,N_19754);
and U20602 (N_20602,N_19758,N_19878);
and U20603 (N_20603,N_19390,N_19722);
nand U20604 (N_20604,N_19635,N_19575);
nand U20605 (N_20605,N_19975,N_19999);
xnor U20606 (N_20606,N_19527,N_19740);
and U20607 (N_20607,N_19999,N_19718);
xor U20608 (N_20608,N_19897,N_19394);
nor U20609 (N_20609,N_19524,N_19634);
and U20610 (N_20610,N_19736,N_19403);
nor U20611 (N_20611,N_19933,N_19449);
or U20612 (N_20612,N_19764,N_19897);
and U20613 (N_20613,N_19621,N_19873);
or U20614 (N_20614,N_19801,N_19968);
nor U20615 (N_20615,N_19759,N_19504);
and U20616 (N_20616,N_19539,N_19714);
and U20617 (N_20617,N_19453,N_19546);
nand U20618 (N_20618,N_19630,N_19555);
and U20619 (N_20619,N_19804,N_19956);
nand U20620 (N_20620,N_19917,N_19614);
nor U20621 (N_20621,N_19472,N_19734);
nor U20622 (N_20622,N_19754,N_19826);
nand U20623 (N_20623,N_19550,N_19445);
nand U20624 (N_20624,N_19669,N_19830);
xor U20625 (N_20625,N_20000,N_20500);
nand U20626 (N_20626,N_20168,N_20102);
nor U20627 (N_20627,N_20189,N_20257);
nand U20628 (N_20628,N_20336,N_20536);
or U20629 (N_20629,N_20303,N_20018);
nor U20630 (N_20630,N_20067,N_20527);
xor U20631 (N_20631,N_20528,N_20581);
xor U20632 (N_20632,N_20237,N_20170);
nand U20633 (N_20633,N_20120,N_20017);
xnor U20634 (N_20634,N_20546,N_20137);
and U20635 (N_20635,N_20006,N_20413);
and U20636 (N_20636,N_20525,N_20555);
nor U20637 (N_20637,N_20521,N_20343);
xor U20638 (N_20638,N_20394,N_20033);
nand U20639 (N_20639,N_20201,N_20330);
nor U20640 (N_20640,N_20534,N_20472);
nor U20641 (N_20641,N_20198,N_20136);
nand U20642 (N_20642,N_20200,N_20299);
nor U20643 (N_20643,N_20434,N_20600);
or U20644 (N_20644,N_20428,N_20476);
nor U20645 (N_20645,N_20441,N_20350);
or U20646 (N_20646,N_20422,N_20453);
xor U20647 (N_20647,N_20072,N_20554);
nor U20648 (N_20648,N_20518,N_20001);
nand U20649 (N_20649,N_20552,N_20030);
and U20650 (N_20650,N_20231,N_20583);
xor U20651 (N_20651,N_20221,N_20541);
xnor U20652 (N_20652,N_20055,N_20436);
and U20653 (N_20653,N_20310,N_20161);
nand U20654 (N_20654,N_20376,N_20175);
nand U20655 (N_20655,N_20213,N_20107);
xor U20656 (N_20656,N_20289,N_20308);
and U20657 (N_20657,N_20331,N_20283);
xor U20658 (N_20658,N_20108,N_20080);
or U20659 (N_20659,N_20409,N_20235);
or U20660 (N_20660,N_20066,N_20022);
nor U20661 (N_20661,N_20362,N_20182);
or U20662 (N_20662,N_20034,N_20370);
xnor U20663 (N_20663,N_20256,N_20602);
or U20664 (N_20664,N_20291,N_20451);
xor U20665 (N_20665,N_20227,N_20010);
nand U20666 (N_20666,N_20269,N_20332);
xnor U20667 (N_20667,N_20079,N_20512);
nor U20668 (N_20668,N_20277,N_20319);
nand U20669 (N_20669,N_20402,N_20239);
or U20670 (N_20670,N_20421,N_20224);
or U20671 (N_20671,N_20333,N_20391);
or U20672 (N_20672,N_20622,N_20106);
nor U20673 (N_20673,N_20075,N_20188);
nor U20674 (N_20674,N_20342,N_20234);
nor U20675 (N_20675,N_20570,N_20608);
nand U20676 (N_20676,N_20290,N_20426);
nand U20677 (N_20677,N_20216,N_20389);
nor U20678 (N_20678,N_20569,N_20432);
nor U20679 (N_20679,N_20065,N_20048);
nor U20680 (N_20680,N_20183,N_20077);
xnor U20681 (N_20681,N_20267,N_20186);
xnor U20682 (N_20682,N_20516,N_20438);
nor U20683 (N_20683,N_20060,N_20191);
or U20684 (N_20684,N_20381,N_20105);
or U20685 (N_20685,N_20217,N_20026);
nand U20686 (N_20686,N_20014,N_20420);
xor U20687 (N_20687,N_20069,N_20222);
nand U20688 (N_20688,N_20568,N_20341);
and U20689 (N_20689,N_20440,N_20247);
and U20690 (N_20690,N_20494,N_20450);
nor U20691 (N_20691,N_20011,N_20495);
nand U20692 (N_20692,N_20276,N_20579);
or U20693 (N_20693,N_20351,N_20225);
and U20694 (N_20694,N_20144,N_20061);
nor U20695 (N_20695,N_20240,N_20544);
xnor U20696 (N_20696,N_20535,N_20326);
xnor U20697 (N_20697,N_20181,N_20088);
or U20698 (N_20698,N_20236,N_20455);
or U20699 (N_20699,N_20160,N_20559);
nand U20700 (N_20700,N_20529,N_20028);
xor U20701 (N_20701,N_20177,N_20359);
nand U20702 (N_20702,N_20003,N_20334);
xor U20703 (N_20703,N_20412,N_20244);
and U20704 (N_20704,N_20415,N_20074);
xor U20705 (N_20705,N_20178,N_20086);
and U20706 (N_20706,N_20251,N_20539);
and U20707 (N_20707,N_20242,N_20171);
and U20708 (N_20708,N_20273,N_20449);
xnor U20709 (N_20709,N_20238,N_20265);
or U20710 (N_20710,N_20384,N_20286);
or U20711 (N_20711,N_20329,N_20561);
nor U20712 (N_20712,N_20123,N_20353);
or U20713 (N_20713,N_20112,N_20511);
or U20714 (N_20714,N_20126,N_20617);
nor U20715 (N_20715,N_20169,N_20173);
nor U20716 (N_20716,N_20513,N_20278);
nand U20717 (N_20717,N_20514,N_20547);
nand U20718 (N_20718,N_20063,N_20280);
xor U20719 (N_20719,N_20557,N_20281);
or U20720 (N_20720,N_20416,N_20604);
and U20721 (N_20721,N_20232,N_20057);
xnor U20722 (N_20722,N_20612,N_20530);
nor U20723 (N_20723,N_20425,N_20548);
and U20724 (N_20724,N_20346,N_20328);
and U20725 (N_20725,N_20383,N_20486);
nor U20726 (N_20726,N_20520,N_20035);
nor U20727 (N_20727,N_20611,N_20214);
and U20728 (N_20728,N_20430,N_20262);
nand U20729 (N_20729,N_20101,N_20574);
nor U20730 (N_20730,N_20228,N_20388);
and U20731 (N_20731,N_20380,N_20143);
or U20732 (N_20732,N_20162,N_20233);
or U20733 (N_20733,N_20406,N_20407);
nor U20734 (N_20734,N_20468,N_20203);
nand U20735 (N_20735,N_20208,N_20373);
and U20736 (N_20736,N_20571,N_20135);
xor U20737 (N_20737,N_20124,N_20129);
xnor U20738 (N_20738,N_20163,N_20410);
xor U20739 (N_20739,N_20385,N_20176);
xnor U20740 (N_20740,N_20305,N_20504);
nand U20741 (N_20741,N_20192,N_20607);
xor U20742 (N_20742,N_20323,N_20053);
and U20743 (N_20743,N_20306,N_20372);
or U20744 (N_20744,N_20081,N_20493);
or U20745 (N_20745,N_20496,N_20253);
and U20746 (N_20746,N_20365,N_20459);
xor U20747 (N_20747,N_20575,N_20586);
nand U20748 (N_20748,N_20464,N_20447);
nor U20749 (N_20749,N_20565,N_20545);
nor U20750 (N_20750,N_20068,N_20109);
nor U20751 (N_20751,N_20230,N_20386);
nand U20752 (N_20752,N_20400,N_20324);
or U20753 (N_20753,N_20471,N_20510);
nand U20754 (N_20754,N_20431,N_20322);
nand U20755 (N_20755,N_20437,N_20229);
or U20756 (N_20756,N_20049,N_20258);
xnor U20757 (N_20757,N_20263,N_20615);
and U20758 (N_20758,N_20138,N_20078);
or U20759 (N_20759,N_20128,N_20429);
or U20760 (N_20760,N_20364,N_20111);
or U20761 (N_20761,N_20016,N_20499);
nor U20762 (N_20762,N_20497,N_20556);
xor U20763 (N_20763,N_20122,N_20311);
nand U20764 (N_20764,N_20134,N_20392);
xor U20765 (N_20765,N_20272,N_20573);
and U20766 (N_20766,N_20195,N_20113);
nand U20767 (N_20767,N_20375,N_20279);
nand U20768 (N_20768,N_20369,N_20368);
nand U20769 (N_20769,N_20588,N_20467);
and U20770 (N_20770,N_20302,N_20300);
nor U20771 (N_20771,N_20096,N_20358);
nor U20772 (N_20772,N_20264,N_20180);
and U20773 (N_20773,N_20360,N_20226);
nor U20774 (N_20774,N_20349,N_20241);
or U20775 (N_20775,N_20427,N_20452);
xnor U20776 (N_20776,N_20344,N_20008);
xor U20777 (N_20777,N_20515,N_20193);
nand U20778 (N_20778,N_20537,N_20533);
xor U20779 (N_20779,N_20318,N_20505);
or U20780 (N_20780,N_20398,N_20356);
nor U20781 (N_20781,N_20097,N_20205);
or U20782 (N_20782,N_20338,N_20531);
or U20783 (N_20783,N_20393,N_20184);
nand U20784 (N_20784,N_20288,N_20352);
or U20785 (N_20785,N_20019,N_20595);
and U20786 (N_20786,N_20032,N_20021);
xnor U20787 (N_20787,N_20139,N_20484);
or U20788 (N_20788,N_20395,N_20592);
nor U20789 (N_20789,N_20149,N_20024);
or U20790 (N_20790,N_20621,N_20605);
or U20791 (N_20791,N_20444,N_20414);
xor U20792 (N_20792,N_20462,N_20485);
xnor U20793 (N_20793,N_20355,N_20606);
or U20794 (N_20794,N_20619,N_20419);
nor U20795 (N_20795,N_20020,N_20089);
xnor U20796 (N_20796,N_20131,N_20293);
or U20797 (N_20797,N_20587,N_20446);
xnor U20798 (N_20798,N_20582,N_20598);
nand U20799 (N_20799,N_20327,N_20073);
nor U20800 (N_20800,N_20085,N_20609);
and U20801 (N_20801,N_20140,N_20524);
and U20802 (N_20802,N_20295,N_20039);
nand U20803 (N_20803,N_20479,N_20147);
nand U20804 (N_20804,N_20558,N_20165);
nand U20805 (N_20805,N_20296,N_20519);
xor U20806 (N_20806,N_20268,N_20478);
nand U20807 (N_20807,N_20614,N_20270);
xor U20808 (N_20808,N_20560,N_20076);
and U20809 (N_20809,N_20481,N_20155);
and U20810 (N_20810,N_20005,N_20127);
and U20811 (N_20811,N_20248,N_20297);
nand U20812 (N_20812,N_20091,N_20087);
and U20813 (N_20813,N_20474,N_20058);
and U20814 (N_20814,N_20204,N_20553);
and U20815 (N_20815,N_20418,N_20218);
nor U20816 (N_20816,N_20354,N_20567);
or U20817 (N_20817,N_20133,N_20501);
nor U20818 (N_20818,N_20146,N_20040);
or U20819 (N_20819,N_20509,N_20317);
xor U20820 (N_20820,N_20532,N_20357);
nand U20821 (N_20821,N_20463,N_20597);
xor U20822 (N_20822,N_20260,N_20118);
xor U20823 (N_20823,N_20220,N_20282);
or U20824 (N_20824,N_20599,N_20526);
and U20825 (N_20825,N_20461,N_20490);
xor U20826 (N_20826,N_20207,N_20275);
or U20827 (N_20827,N_20564,N_20578);
nand U20828 (N_20828,N_20209,N_20114);
or U20829 (N_20829,N_20397,N_20340);
or U20830 (N_20830,N_20002,N_20448);
and U20831 (N_20831,N_20488,N_20004);
nand U20832 (N_20832,N_20050,N_20196);
nand U20833 (N_20833,N_20036,N_20543);
or U20834 (N_20834,N_20550,N_20245);
nor U20835 (N_20835,N_20590,N_20266);
xor U20836 (N_20836,N_20156,N_20377);
nor U20837 (N_20837,N_20435,N_20417);
nor U20838 (N_20838,N_20202,N_20287);
and U20839 (N_20839,N_20292,N_20012);
nor U20840 (N_20840,N_20007,N_20577);
and U20841 (N_20841,N_20572,N_20603);
nand U20842 (N_20842,N_20285,N_20041);
or U20843 (N_20843,N_20199,N_20460);
and U20844 (N_20844,N_20094,N_20580);
nand U20845 (N_20845,N_20145,N_20366);
nor U20846 (N_20846,N_20104,N_20158);
and U20847 (N_20847,N_20132,N_20348);
nor U20848 (N_20848,N_20454,N_20445);
and U20849 (N_20849,N_20387,N_20092);
nor U20850 (N_20850,N_20411,N_20623);
or U20851 (N_20851,N_20491,N_20480);
nor U20852 (N_20852,N_20401,N_20037);
and U20853 (N_20853,N_20506,N_20616);
and U20854 (N_20854,N_20507,N_20125);
and U20855 (N_20855,N_20103,N_20059);
xnor U20856 (N_20856,N_20027,N_20093);
nor U20857 (N_20857,N_20082,N_20215);
nand U20858 (N_20858,N_20254,N_20307);
or U20859 (N_20859,N_20013,N_20054);
and U20860 (N_20860,N_20423,N_20009);
and U20861 (N_20861,N_20274,N_20584);
xor U20862 (N_20862,N_20403,N_20259);
xor U20863 (N_20863,N_20363,N_20371);
or U20864 (N_20864,N_20456,N_20433);
xnor U20865 (N_20865,N_20115,N_20071);
nor U20866 (N_20866,N_20031,N_20457);
nor U20867 (N_20867,N_20255,N_20110);
nor U20868 (N_20868,N_20052,N_20470);
nor U20869 (N_20869,N_20045,N_20206);
nand U20870 (N_20870,N_20172,N_20190);
nand U20871 (N_20871,N_20439,N_20374);
xnor U20872 (N_20872,N_20601,N_20469);
nand U20873 (N_20873,N_20185,N_20084);
and U20874 (N_20874,N_20150,N_20339);
and U20875 (N_20875,N_20298,N_20566);
xor U20876 (N_20876,N_20424,N_20522);
nor U20877 (N_20877,N_20047,N_20025);
nor U20878 (N_20878,N_20154,N_20367);
and U20879 (N_20879,N_20624,N_20100);
and U20880 (N_20880,N_20443,N_20179);
nor U20881 (N_20881,N_20502,N_20489);
and U20882 (N_20882,N_20166,N_20117);
xnor U20883 (N_20883,N_20261,N_20396);
nand U20884 (N_20884,N_20315,N_20314);
and U20885 (N_20885,N_20508,N_20064);
nand U20886 (N_20886,N_20187,N_20090);
nand U20887 (N_20887,N_20159,N_20157);
nor U20888 (N_20888,N_20466,N_20458);
or U20889 (N_20889,N_20405,N_20465);
nand U20890 (N_20890,N_20141,N_20116);
or U20891 (N_20891,N_20316,N_20473);
nand U20892 (N_20892,N_20294,N_20325);
nand U20893 (N_20893,N_20210,N_20042);
or U20894 (N_20894,N_20249,N_20345);
or U20895 (N_20895,N_20098,N_20596);
xnor U20896 (N_20896,N_20503,N_20099);
nor U20897 (N_20897,N_20593,N_20378);
and U20898 (N_20898,N_20442,N_20591);
nand U20899 (N_20899,N_20618,N_20194);
xor U20900 (N_20900,N_20038,N_20492);
nor U20901 (N_20901,N_20337,N_20549);
nor U20902 (N_20902,N_20540,N_20211);
or U20903 (N_20903,N_20152,N_20121);
nand U20904 (N_20904,N_20223,N_20361);
and U20905 (N_20905,N_20610,N_20301);
and U20906 (N_20906,N_20482,N_20271);
nor U20907 (N_20907,N_20219,N_20284);
nand U20908 (N_20908,N_20197,N_20167);
nand U20909 (N_20909,N_20051,N_20562);
nor U20910 (N_20910,N_20044,N_20309);
nor U20911 (N_20911,N_20589,N_20404);
nand U20912 (N_20912,N_20119,N_20174);
nor U20913 (N_20913,N_20250,N_20585);
xnor U20914 (N_20914,N_20576,N_20320);
xnor U20915 (N_20915,N_20408,N_20538);
and U20916 (N_20916,N_20312,N_20475);
xnor U20917 (N_20917,N_20083,N_20095);
nand U20918 (N_20918,N_20563,N_20243);
xnor U20919 (N_20919,N_20542,N_20379);
or U20920 (N_20920,N_20062,N_20551);
nand U20921 (N_20921,N_20523,N_20382);
nor U20922 (N_20922,N_20023,N_20252);
nand U20923 (N_20923,N_20620,N_20321);
and U20924 (N_20924,N_20517,N_20594);
and U20925 (N_20925,N_20153,N_20151);
nand U20926 (N_20926,N_20043,N_20483);
or U20927 (N_20927,N_20015,N_20046);
nor U20928 (N_20928,N_20142,N_20029);
xor U20929 (N_20929,N_20613,N_20212);
or U20930 (N_20930,N_20148,N_20477);
xor U20931 (N_20931,N_20347,N_20399);
or U20932 (N_20932,N_20056,N_20130);
nor U20933 (N_20933,N_20304,N_20498);
or U20934 (N_20934,N_20390,N_20070);
xor U20935 (N_20935,N_20313,N_20487);
or U20936 (N_20936,N_20164,N_20246);
or U20937 (N_20937,N_20335,N_20529);
nor U20938 (N_20938,N_20576,N_20598);
or U20939 (N_20939,N_20527,N_20314);
nand U20940 (N_20940,N_20201,N_20268);
xor U20941 (N_20941,N_20060,N_20293);
xnor U20942 (N_20942,N_20600,N_20594);
nor U20943 (N_20943,N_20290,N_20021);
xnor U20944 (N_20944,N_20008,N_20610);
nor U20945 (N_20945,N_20272,N_20345);
nor U20946 (N_20946,N_20206,N_20615);
xor U20947 (N_20947,N_20621,N_20373);
nor U20948 (N_20948,N_20592,N_20564);
or U20949 (N_20949,N_20533,N_20014);
and U20950 (N_20950,N_20513,N_20531);
xnor U20951 (N_20951,N_20137,N_20317);
nand U20952 (N_20952,N_20094,N_20583);
xor U20953 (N_20953,N_20059,N_20559);
xor U20954 (N_20954,N_20379,N_20377);
and U20955 (N_20955,N_20283,N_20500);
and U20956 (N_20956,N_20271,N_20067);
xnor U20957 (N_20957,N_20307,N_20020);
nand U20958 (N_20958,N_20160,N_20615);
or U20959 (N_20959,N_20541,N_20144);
and U20960 (N_20960,N_20347,N_20374);
or U20961 (N_20961,N_20321,N_20183);
or U20962 (N_20962,N_20308,N_20281);
and U20963 (N_20963,N_20300,N_20176);
xnor U20964 (N_20964,N_20608,N_20206);
nor U20965 (N_20965,N_20346,N_20517);
nand U20966 (N_20966,N_20425,N_20407);
and U20967 (N_20967,N_20566,N_20457);
nor U20968 (N_20968,N_20340,N_20514);
xor U20969 (N_20969,N_20190,N_20523);
or U20970 (N_20970,N_20293,N_20537);
and U20971 (N_20971,N_20061,N_20037);
or U20972 (N_20972,N_20591,N_20044);
nand U20973 (N_20973,N_20412,N_20346);
or U20974 (N_20974,N_20035,N_20528);
xor U20975 (N_20975,N_20218,N_20536);
or U20976 (N_20976,N_20425,N_20043);
nand U20977 (N_20977,N_20211,N_20292);
and U20978 (N_20978,N_20160,N_20281);
and U20979 (N_20979,N_20065,N_20017);
or U20980 (N_20980,N_20198,N_20525);
and U20981 (N_20981,N_20327,N_20294);
xor U20982 (N_20982,N_20113,N_20118);
and U20983 (N_20983,N_20419,N_20338);
nand U20984 (N_20984,N_20584,N_20179);
nand U20985 (N_20985,N_20570,N_20409);
and U20986 (N_20986,N_20282,N_20512);
and U20987 (N_20987,N_20176,N_20008);
nor U20988 (N_20988,N_20022,N_20498);
nand U20989 (N_20989,N_20387,N_20045);
and U20990 (N_20990,N_20487,N_20542);
nor U20991 (N_20991,N_20466,N_20433);
and U20992 (N_20992,N_20097,N_20355);
nand U20993 (N_20993,N_20233,N_20239);
and U20994 (N_20994,N_20125,N_20023);
nor U20995 (N_20995,N_20114,N_20397);
or U20996 (N_20996,N_20451,N_20188);
nor U20997 (N_20997,N_20379,N_20421);
or U20998 (N_20998,N_20458,N_20064);
nor U20999 (N_20999,N_20076,N_20464);
or U21000 (N_21000,N_20130,N_20140);
or U21001 (N_21001,N_20621,N_20117);
or U21002 (N_21002,N_20095,N_20287);
xor U21003 (N_21003,N_20114,N_20300);
and U21004 (N_21004,N_20399,N_20218);
and U21005 (N_21005,N_20480,N_20009);
xor U21006 (N_21006,N_20496,N_20200);
and U21007 (N_21007,N_20251,N_20552);
and U21008 (N_21008,N_20542,N_20608);
nor U21009 (N_21009,N_20573,N_20621);
and U21010 (N_21010,N_20091,N_20601);
and U21011 (N_21011,N_20335,N_20356);
nor U21012 (N_21012,N_20534,N_20554);
nor U21013 (N_21013,N_20156,N_20208);
and U21014 (N_21014,N_20257,N_20064);
and U21015 (N_21015,N_20398,N_20329);
nand U21016 (N_21016,N_20390,N_20457);
xnor U21017 (N_21017,N_20225,N_20050);
and U21018 (N_21018,N_20575,N_20410);
and U21019 (N_21019,N_20602,N_20305);
or U21020 (N_21020,N_20614,N_20377);
and U21021 (N_21021,N_20173,N_20309);
xor U21022 (N_21022,N_20026,N_20036);
nand U21023 (N_21023,N_20100,N_20587);
xnor U21024 (N_21024,N_20386,N_20024);
nand U21025 (N_21025,N_20374,N_20280);
nand U21026 (N_21026,N_20321,N_20524);
nand U21027 (N_21027,N_20182,N_20621);
nor U21028 (N_21028,N_20316,N_20179);
xor U21029 (N_21029,N_20555,N_20300);
nor U21030 (N_21030,N_20209,N_20159);
and U21031 (N_21031,N_20125,N_20472);
nand U21032 (N_21032,N_20415,N_20255);
xor U21033 (N_21033,N_20337,N_20171);
xnor U21034 (N_21034,N_20570,N_20372);
or U21035 (N_21035,N_20325,N_20389);
xnor U21036 (N_21036,N_20011,N_20017);
nor U21037 (N_21037,N_20553,N_20325);
nand U21038 (N_21038,N_20322,N_20116);
or U21039 (N_21039,N_20541,N_20087);
nand U21040 (N_21040,N_20371,N_20616);
and U21041 (N_21041,N_20183,N_20349);
nor U21042 (N_21042,N_20594,N_20204);
xnor U21043 (N_21043,N_20515,N_20350);
nor U21044 (N_21044,N_20470,N_20409);
or U21045 (N_21045,N_20138,N_20077);
nand U21046 (N_21046,N_20608,N_20133);
nor U21047 (N_21047,N_20065,N_20294);
or U21048 (N_21048,N_20593,N_20133);
or U21049 (N_21049,N_20290,N_20495);
nand U21050 (N_21050,N_20393,N_20111);
xnor U21051 (N_21051,N_20314,N_20424);
xor U21052 (N_21052,N_20202,N_20201);
nor U21053 (N_21053,N_20288,N_20240);
or U21054 (N_21054,N_20050,N_20156);
nor U21055 (N_21055,N_20035,N_20602);
and U21056 (N_21056,N_20263,N_20209);
nand U21057 (N_21057,N_20224,N_20274);
xor U21058 (N_21058,N_20413,N_20369);
nor U21059 (N_21059,N_20402,N_20112);
nor U21060 (N_21060,N_20010,N_20405);
or U21061 (N_21061,N_20452,N_20407);
xor U21062 (N_21062,N_20381,N_20034);
xor U21063 (N_21063,N_20082,N_20597);
xor U21064 (N_21064,N_20254,N_20023);
nand U21065 (N_21065,N_20552,N_20224);
and U21066 (N_21066,N_20227,N_20173);
nor U21067 (N_21067,N_20269,N_20479);
or U21068 (N_21068,N_20073,N_20600);
nor U21069 (N_21069,N_20292,N_20271);
nand U21070 (N_21070,N_20579,N_20437);
or U21071 (N_21071,N_20143,N_20480);
nand U21072 (N_21072,N_20264,N_20223);
and U21073 (N_21073,N_20514,N_20604);
nor U21074 (N_21074,N_20351,N_20396);
or U21075 (N_21075,N_20050,N_20319);
or U21076 (N_21076,N_20417,N_20264);
or U21077 (N_21077,N_20416,N_20142);
nor U21078 (N_21078,N_20330,N_20508);
or U21079 (N_21079,N_20248,N_20130);
nand U21080 (N_21080,N_20302,N_20064);
or U21081 (N_21081,N_20213,N_20300);
nand U21082 (N_21082,N_20244,N_20489);
nand U21083 (N_21083,N_20023,N_20396);
xnor U21084 (N_21084,N_20223,N_20390);
nand U21085 (N_21085,N_20288,N_20619);
nor U21086 (N_21086,N_20607,N_20392);
nor U21087 (N_21087,N_20113,N_20608);
nand U21088 (N_21088,N_20203,N_20130);
or U21089 (N_21089,N_20203,N_20610);
nand U21090 (N_21090,N_20599,N_20252);
nand U21091 (N_21091,N_20253,N_20601);
nor U21092 (N_21092,N_20152,N_20179);
xnor U21093 (N_21093,N_20601,N_20450);
and U21094 (N_21094,N_20496,N_20373);
nand U21095 (N_21095,N_20479,N_20443);
nor U21096 (N_21096,N_20613,N_20196);
nor U21097 (N_21097,N_20302,N_20054);
xor U21098 (N_21098,N_20261,N_20129);
and U21099 (N_21099,N_20245,N_20580);
xnor U21100 (N_21100,N_20222,N_20001);
nand U21101 (N_21101,N_20441,N_20162);
nand U21102 (N_21102,N_20019,N_20284);
xor U21103 (N_21103,N_20318,N_20050);
or U21104 (N_21104,N_20315,N_20375);
nand U21105 (N_21105,N_20299,N_20079);
xnor U21106 (N_21106,N_20465,N_20230);
xor U21107 (N_21107,N_20425,N_20212);
xnor U21108 (N_21108,N_20539,N_20240);
and U21109 (N_21109,N_20054,N_20273);
and U21110 (N_21110,N_20202,N_20084);
and U21111 (N_21111,N_20242,N_20164);
xor U21112 (N_21112,N_20422,N_20212);
nor U21113 (N_21113,N_20573,N_20495);
nor U21114 (N_21114,N_20075,N_20113);
nand U21115 (N_21115,N_20422,N_20457);
or U21116 (N_21116,N_20336,N_20326);
and U21117 (N_21117,N_20001,N_20588);
xnor U21118 (N_21118,N_20084,N_20514);
nand U21119 (N_21119,N_20600,N_20102);
xor U21120 (N_21120,N_20319,N_20447);
and U21121 (N_21121,N_20351,N_20590);
xnor U21122 (N_21122,N_20137,N_20243);
or U21123 (N_21123,N_20063,N_20616);
and U21124 (N_21124,N_20409,N_20374);
or U21125 (N_21125,N_20124,N_20121);
and U21126 (N_21126,N_20177,N_20011);
or U21127 (N_21127,N_20060,N_20585);
nand U21128 (N_21128,N_20062,N_20425);
nand U21129 (N_21129,N_20292,N_20126);
xnor U21130 (N_21130,N_20475,N_20431);
xnor U21131 (N_21131,N_20107,N_20220);
or U21132 (N_21132,N_20531,N_20205);
nor U21133 (N_21133,N_20248,N_20566);
nand U21134 (N_21134,N_20360,N_20267);
nor U21135 (N_21135,N_20521,N_20099);
xor U21136 (N_21136,N_20489,N_20466);
nand U21137 (N_21137,N_20152,N_20062);
nor U21138 (N_21138,N_20223,N_20136);
and U21139 (N_21139,N_20094,N_20439);
and U21140 (N_21140,N_20381,N_20624);
or U21141 (N_21141,N_20621,N_20617);
and U21142 (N_21142,N_20307,N_20541);
or U21143 (N_21143,N_20081,N_20056);
and U21144 (N_21144,N_20208,N_20517);
and U21145 (N_21145,N_20116,N_20456);
nand U21146 (N_21146,N_20538,N_20618);
and U21147 (N_21147,N_20184,N_20347);
nand U21148 (N_21148,N_20148,N_20000);
or U21149 (N_21149,N_20273,N_20089);
xor U21150 (N_21150,N_20128,N_20263);
and U21151 (N_21151,N_20234,N_20093);
and U21152 (N_21152,N_20210,N_20343);
xor U21153 (N_21153,N_20124,N_20005);
and U21154 (N_21154,N_20164,N_20269);
and U21155 (N_21155,N_20183,N_20211);
or U21156 (N_21156,N_20187,N_20278);
nor U21157 (N_21157,N_20460,N_20576);
xor U21158 (N_21158,N_20310,N_20000);
nand U21159 (N_21159,N_20307,N_20067);
nor U21160 (N_21160,N_20502,N_20015);
xnor U21161 (N_21161,N_20367,N_20430);
nand U21162 (N_21162,N_20514,N_20090);
and U21163 (N_21163,N_20014,N_20146);
and U21164 (N_21164,N_20551,N_20080);
xor U21165 (N_21165,N_20029,N_20320);
nor U21166 (N_21166,N_20598,N_20480);
xor U21167 (N_21167,N_20072,N_20282);
or U21168 (N_21168,N_20419,N_20011);
nand U21169 (N_21169,N_20175,N_20130);
nand U21170 (N_21170,N_20317,N_20432);
nor U21171 (N_21171,N_20149,N_20202);
nor U21172 (N_21172,N_20528,N_20395);
or U21173 (N_21173,N_20406,N_20527);
or U21174 (N_21174,N_20025,N_20087);
xnor U21175 (N_21175,N_20317,N_20154);
nor U21176 (N_21176,N_20363,N_20455);
xnor U21177 (N_21177,N_20054,N_20404);
nand U21178 (N_21178,N_20385,N_20575);
and U21179 (N_21179,N_20144,N_20549);
or U21180 (N_21180,N_20347,N_20072);
or U21181 (N_21181,N_20077,N_20328);
nand U21182 (N_21182,N_20192,N_20623);
nor U21183 (N_21183,N_20189,N_20319);
nand U21184 (N_21184,N_20024,N_20462);
nor U21185 (N_21185,N_20234,N_20132);
nor U21186 (N_21186,N_20506,N_20021);
and U21187 (N_21187,N_20231,N_20476);
xor U21188 (N_21188,N_20144,N_20269);
and U21189 (N_21189,N_20248,N_20021);
or U21190 (N_21190,N_20259,N_20178);
xnor U21191 (N_21191,N_20227,N_20333);
xor U21192 (N_21192,N_20024,N_20425);
xor U21193 (N_21193,N_20098,N_20233);
xnor U21194 (N_21194,N_20319,N_20110);
or U21195 (N_21195,N_20013,N_20500);
and U21196 (N_21196,N_20158,N_20014);
or U21197 (N_21197,N_20562,N_20127);
and U21198 (N_21198,N_20001,N_20525);
and U21199 (N_21199,N_20513,N_20593);
or U21200 (N_21200,N_20288,N_20229);
and U21201 (N_21201,N_20026,N_20464);
nand U21202 (N_21202,N_20560,N_20280);
nor U21203 (N_21203,N_20193,N_20041);
or U21204 (N_21204,N_20439,N_20337);
nor U21205 (N_21205,N_20601,N_20073);
or U21206 (N_21206,N_20331,N_20063);
and U21207 (N_21207,N_20309,N_20513);
and U21208 (N_21208,N_20057,N_20461);
and U21209 (N_21209,N_20512,N_20264);
or U21210 (N_21210,N_20318,N_20172);
nand U21211 (N_21211,N_20372,N_20129);
xnor U21212 (N_21212,N_20574,N_20104);
xnor U21213 (N_21213,N_20199,N_20192);
xor U21214 (N_21214,N_20482,N_20586);
nand U21215 (N_21215,N_20463,N_20244);
or U21216 (N_21216,N_20339,N_20237);
nand U21217 (N_21217,N_20306,N_20425);
nand U21218 (N_21218,N_20270,N_20121);
and U21219 (N_21219,N_20370,N_20020);
xnor U21220 (N_21220,N_20483,N_20617);
nand U21221 (N_21221,N_20446,N_20023);
nor U21222 (N_21222,N_20337,N_20514);
nor U21223 (N_21223,N_20548,N_20502);
xor U21224 (N_21224,N_20282,N_20436);
nand U21225 (N_21225,N_20266,N_20389);
and U21226 (N_21226,N_20045,N_20098);
or U21227 (N_21227,N_20485,N_20454);
and U21228 (N_21228,N_20422,N_20246);
nand U21229 (N_21229,N_20162,N_20485);
xnor U21230 (N_21230,N_20366,N_20601);
and U21231 (N_21231,N_20066,N_20036);
nor U21232 (N_21232,N_20365,N_20529);
xnor U21233 (N_21233,N_20266,N_20258);
and U21234 (N_21234,N_20184,N_20411);
or U21235 (N_21235,N_20118,N_20571);
xnor U21236 (N_21236,N_20193,N_20335);
and U21237 (N_21237,N_20342,N_20132);
or U21238 (N_21238,N_20507,N_20049);
xor U21239 (N_21239,N_20346,N_20504);
and U21240 (N_21240,N_20288,N_20616);
xnor U21241 (N_21241,N_20109,N_20417);
and U21242 (N_21242,N_20119,N_20507);
or U21243 (N_21243,N_20300,N_20212);
nor U21244 (N_21244,N_20257,N_20332);
or U21245 (N_21245,N_20395,N_20024);
xnor U21246 (N_21246,N_20345,N_20405);
and U21247 (N_21247,N_20218,N_20034);
nor U21248 (N_21248,N_20303,N_20199);
nor U21249 (N_21249,N_20112,N_20303);
nor U21250 (N_21250,N_20833,N_21059);
or U21251 (N_21251,N_21205,N_20687);
or U21252 (N_21252,N_20739,N_21200);
and U21253 (N_21253,N_20671,N_21120);
or U21254 (N_21254,N_21169,N_20946);
xor U21255 (N_21255,N_20903,N_20679);
nand U21256 (N_21256,N_20939,N_21082);
and U21257 (N_21257,N_20738,N_20862);
nand U21258 (N_21258,N_20930,N_21209);
nor U21259 (N_21259,N_21030,N_21119);
or U21260 (N_21260,N_21098,N_20987);
and U21261 (N_21261,N_21087,N_20649);
nand U21262 (N_21262,N_20711,N_21151);
xnor U21263 (N_21263,N_20696,N_21029);
xnor U21264 (N_21264,N_20960,N_21016);
nor U21265 (N_21265,N_20742,N_20702);
nor U21266 (N_21266,N_20958,N_20855);
xnor U21267 (N_21267,N_20873,N_21074);
and U21268 (N_21268,N_20654,N_20749);
nor U21269 (N_21269,N_20854,N_20916);
nand U21270 (N_21270,N_20648,N_21076);
or U21271 (N_21271,N_20819,N_21010);
nand U21272 (N_21272,N_21034,N_21245);
and U21273 (N_21273,N_20662,N_20999);
and U21274 (N_21274,N_21242,N_20945);
nand U21275 (N_21275,N_20674,N_20911);
or U21276 (N_21276,N_20970,N_20975);
and U21277 (N_21277,N_20974,N_20844);
nor U21278 (N_21278,N_20751,N_21086);
nand U21279 (N_21279,N_20697,N_21116);
nand U21280 (N_21280,N_21056,N_21071);
nor U21281 (N_21281,N_21094,N_20796);
nand U21282 (N_21282,N_21130,N_21182);
or U21283 (N_21283,N_20898,N_20949);
nand U21284 (N_21284,N_20994,N_20691);
nand U21285 (N_21285,N_20758,N_20972);
and U21286 (N_21286,N_20744,N_20721);
nor U21287 (N_21287,N_20954,N_20772);
or U21288 (N_21288,N_20966,N_21051);
xor U21289 (N_21289,N_21229,N_21234);
and U21290 (N_21290,N_21241,N_20646);
and U21291 (N_21291,N_20664,N_20809);
nor U21292 (N_21292,N_20735,N_21045);
xnor U21293 (N_21293,N_20821,N_20889);
nand U21294 (N_21294,N_21238,N_20813);
nor U21295 (N_21295,N_20703,N_20732);
xor U21296 (N_21296,N_20912,N_21044);
and U21297 (N_21297,N_20978,N_21002);
or U21298 (N_21298,N_20938,N_20667);
or U21299 (N_21299,N_21084,N_21054);
or U21300 (N_21300,N_21025,N_21220);
nand U21301 (N_21301,N_21068,N_20681);
xor U21302 (N_21302,N_21052,N_21136);
or U21303 (N_21303,N_21118,N_20715);
nor U21304 (N_21304,N_20773,N_20668);
nand U21305 (N_21305,N_20766,N_21000);
or U21306 (N_21306,N_20767,N_20980);
and U21307 (N_21307,N_20686,N_21104);
and U21308 (N_21308,N_20811,N_20810);
and U21309 (N_21309,N_20861,N_21058);
nor U21310 (N_21310,N_21228,N_21127);
xor U21311 (N_21311,N_21176,N_20657);
nor U21312 (N_21312,N_20940,N_20942);
and U21313 (N_21313,N_20841,N_21036);
or U21314 (N_21314,N_20706,N_20734);
xor U21315 (N_21315,N_20753,N_20656);
or U21316 (N_21316,N_20757,N_21175);
nor U21317 (N_21317,N_21223,N_20745);
or U21318 (N_21318,N_20948,N_20924);
nand U21319 (N_21319,N_21244,N_21005);
nor U21320 (N_21320,N_20723,N_20842);
or U21321 (N_21321,N_20909,N_21188);
or U21322 (N_21322,N_21167,N_20799);
or U21323 (N_21323,N_20719,N_21201);
xnor U21324 (N_21324,N_20802,N_21124);
or U21325 (N_21325,N_20776,N_20857);
nand U21326 (N_21326,N_20786,N_21077);
nand U21327 (N_21327,N_21100,N_21021);
xnor U21328 (N_21328,N_21221,N_20806);
or U21329 (N_21329,N_20902,N_20878);
xnor U21330 (N_21330,N_21199,N_20793);
or U21331 (N_21331,N_20965,N_20957);
xnor U21332 (N_21332,N_20659,N_21011);
and U21333 (N_21333,N_20777,N_20641);
xor U21334 (N_21334,N_20655,N_20666);
xnor U21335 (N_21335,N_21121,N_21164);
xor U21336 (N_21336,N_20736,N_21180);
nor U21337 (N_21337,N_21227,N_20929);
xor U21338 (N_21338,N_20881,N_21183);
and U21339 (N_21339,N_20825,N_21125);
xor U21340 (N_21340,N_21111,N_20997);
nand U21341 (N_21341,N_20684,N_20725);
and U21342 (N_21342,N_20823,N_21143);
or U21343 (N_21343,N_20710,N_21191);
and U21344 (N_21344,N_21133,N_20636);
nor U21345 (N_21345,N_21023,N_21018);
nor U21346 (N_21346,N_20762,N_21114);
nor U21347 (N_21347,N_20625,N_21152);
xor U21348 (N_21348,N_21017,N_20820);
nand U21349 (N_21349,N_21075,N_20993);
and U21350 (N_21350,N_20784,N_21091);
or U21351 (N_21351,N_21181,N_21173);
or U21352 (N_21352,N_20683,N_20678);
and U21353 (N_21353,N_21050,N_20778);
and U21354 (N_21354,N_21078,N_20952);
nor U21355 (N_21355,N_21240,N_21177);
nand U21356 (N_21356,N_21232,N_20906);
xnor U21357 (N_21357,N_20673,N_20728);
xnor U21358 (N_21358,N_20992,N_21083);
xnor U21359 (N_21359,N_20832,N_21207);
xnor U21360 (N_21360,N_20866,N_20890);
xor U21361 (N_21361,N_20722,N_21093);
nand U21362 (N_21362,N_21105,N_20801);
nor U21363 (N_21363,N_21186,N_20724);
or U21364 (N_21364,N_20869,N_20926);
or U21365 (N_21365,N_20921,N_20707);
or U21366 (N_21366,N_20677,N_20635);
nand U21367 (N_21367,N_20849,N_20733);
or U21368 (N_21368,N_21080,N_21189);
and U21369 (N_21369,N_21069,N_20834);
xor U21370 (N_21370,N_21128,N_20934);
xor U21371 (N_21371,N_21063,N_20913);
and U21372 (N_21372,N_21032,N_21003);
and U21373 (N_21373,N_20918,N_21145);
xor U21374 (N_21374,N_21148,N_20631);
nand U21375 (N_21375,N_21190,N_21024);
or U21376 (N_21376,N_21212,N_20851);
nand U21377 (N_21377,N_20872,N_21088);
and U21378 (N_21378,N_21066,N_20914);
and U21379 (N_21379,N_21060,N_20863);
or U21380 (N_21380,N_21217,N_20689);
and U21381 (N_21381,N_20840,N_21043);
xor U21382 (N_21382,N_21197,N_21213);
or U21383 (N_21383,N_21172,N_21141);
xnor U21384 (N_21384,N_21149,N_21135);
and U21385 (N_21385,N_20893,N_20676);
nor U21386 (N_21386,N_21062,N_20729);
and U21387 (N_21387,N_20865,N_20953);
nand U21388 (N_21388,N_20627,N_20877);
xnor U21389 (N_21389,N_21057,N_20637);
xor U21390 (N_21390,N_20685,N_20800);
xnor U21391 (N_21391,N_20737,N_21165);
nor U21392 (N_21392,N_21004,N_20829);
xor U21393 (N_21393,N_21219,N_21211);
xnor U21394 (N_21394,N_20850,N_20752);
or U21395 (N_21395,N_20956,N_20748);
or U21396 (N_21396,N_21147,N_21142);
xor U21397 (N_21397,N_20640,N_21047);
and U21398 (N_21398,N_20812,N_20884);
and U21399 (N_21399,N_20629,N_21067);
or U21400 (N_21400,N_21184,N_20870);
and U21401 (N_21401,N_21112,N_20962);
xor U21402 (N_21402,N_21028,N_20920);
nor U21403 (N_21403,N_20955,N_20838);
and U21404 (N_21404,N_20808,N_20860);
nand U21405 (N_21405,N_20897,N_21019);
or U21406 (N_21406,N_20986,N_21239);
xor U21407 (N_21407,N_20991,N_21014);
or U21408 (N_21408,N_20647,N_20937);
or U21409 (N_21409,N_20643,N_20756);
or U21410 (N_21410,N_20791,N_20781);
nand U21411 (N_21411,N_20818,N_20936);
nand U21412 (N_21412,N_21150,N_21122);
nor U21413 (N_21413,N_20682,N_20699);
or U21414 (N_21414,N_20690,N_21138);
or U21415 (N_21415,N_21026,N_21132);
nor U21416 (N_21416,N_20983,N_21170);
xnor U21417 (N_21417,N_20754,N_20848);
and U21418 (N_21418,N_20891,N_20988);
and U21419 (N_21419,N_20634,N_21162);
nor U21420 (N_21420,N_20705,N_21095);
xor U21421 (N_21421,N_21048,N_20971);
xnor U21422 (N_21422,N_21117,N_21085);
nand U21423 (N_21423,N_20713,N_20933);
xnor U21424 (N_21424,N_20894,N_20651);
xnor U21425 (N_21425,N_20831,N_20700);
or U21426 (N_21426,N_21102,N_20899);
nor U21427 (N_21427,N_20922,N_21161);
nor U21428 (N_21428,N_21160,N_20822);
xor U21429 (N_21429,N_20680,N_20915);
or U21430 (N_21430,N_21031,N_21099);
and U21431 (N_21431,N_20882,N_20868);
and U21432 (N_21432,N_21230,N_20704);
nor U21433 (N_21433,N_20886,N_21070);
or U21434 (N_21434,N_20910,N_20900);
or U21435 (N_21435,N_20653,N_20874);
nor U21436 (N_21436,N_21187,N_20720);
xnor U21437 (N_21437,N_20935,N_21163);
and U21438 (N_21438,N_21178,N_21129);
or U21439 (N_21439,N_21049,N_21109);
xnor U21440 (N_21440,N_21065,N_21215);
nor U21441 (N_21441,N_21210,N_20905);
and U21442 (N_21442,N_21154,N_20963);
nor U21443 (N_21443,N_20787,N_20765);
and U21444 (N_21444,N_20714,N_20969);
nor U21445 (N_21445,N_20780,N_20759);
xor U21446 (N_21446,N_20947,N_20904);
or U21447 (N_21447,N_20814,N_20964);
nand U21448 (N_21448,N_21249,N_21137);
xor U21449 (N_21449,N_20709,N_20803);
nand U21450 (N_21450,N_21020,N_20642);
xor U21451 (N_21451,N_21103,N_20750);
and U21452 (N_21452,N_20896,N_20928);
or U21453 (N_21453,N_20712,N_21146);
xor U21454 (N_21454,N_21222,N_21134);
and U21455 (N_21455,N_20650,N_20645);
nand U21456 (N_21456,N_21153,N_20984);
or U21457 (N_21457,N_20917,N_20695);
or U21458 (N_21458,N_20764,N_20967);
nor U21459 (N_21459,N_21022,N_21140);
and U21460 (N_21460,N_21101,N_21041);
nand U21461 (N_21461,N_21131,N_20856);
nor U21462 (N_21462,N_21224,N_20785);
and U21463 (N_21463,N_20768,N_21090);
xnor U21464 (N_21464,N_20731,N_21168);
and U21465 (N_21465,N_20977,N_20741);
and U21466 (N_21466,N_21092,N_20830);
or U21467 (N_21467,N_20726,N_20788);
nor U21468 (N_21468,N_21246,N_20846);
nand U21469 (N_21469,N_21206,N_21193);
or U21470 (N_21470,N_20716,N_20839);
nand U21471 (N_21471,N_21144,N_20774);
nand U21472 (N_21472,N_21123,N_20845);
and U21473 (N_21473,N_20740,N_20760);
xnor U21474 (N_21474,N_20730,N_20998);
and U21475 (N_21475,N_21007,N_21073);
or U21476 (N_21476,N_21243,N_20816);
and U21477 (N_21477,N_20805,N_20927);
nand U21478 (N_21478,N_21115,N_20989);
nand U21479 (N_21479,N_21156,N_20626);
nor U21480 (N_21480,N_21248,N_21008);
nor U21481 (N_21481,N_21089,N_20919);
nor U21482 (N_21482,N_20782,N_21126);
or U21483 (N_21483,N_20853,N_20644);
nor U21484 (N_21484,N_21108,N_20888);
nor U21485 (N_21485,N_20794,N_20828);
xnor U21486 (N_21486,N_21055,N_21195);
xor U21487 (N_21487,N_21040,N_20652);
nand U21488 (N_21488,N_21097,N_20835);
or U21489 (N_21489,N_20923,N_20661);
nand U21490 (N_21490,N_20982,N_20961);
xor U21491 (N_21491,N_20901,N_20824);
nor U21492 (N_21492,N_21113,N_20995);
nand U21493 (N_21493,N_21196,N_21012);
and U21494 (N_21494,N_20694,N_20792);
nand U21495 (N_21495,N_20864,N_21009);
and U21496 (N_21496,N_20826,N_20769);
or U21497 (N_21497,N_21096,N_20718);
nand U21498 (N_21498,N_21174,N_20672);
or U21499 (N_21499,N_21001,N_20979);
and U21500 (N_21500,N_21192,N_21237);
xor U21501 (N_21501,N_20632,N_20795);
nand U21502 (N_21502,N_21158,N_20827);
nand U21503 (N_21503,N_21081,N_20951);
or U21504 (N_21504,N_21233,N_21015);
nand U21505 (N_21505,N_20943,N_20698);
or U21506 (N_21506,N_21208,N_21203);
and U21507 (N_21507,N_20633,N_21235);
nor U21508 (N_21508,N_20996,N_20675);
xnor U21509 (N_21509,N_21046,N_21006);
xnor U21510 (N_21510,N_20883,N_21110);
nand U21511 (N_21511,N_20670,N_21039);
or U21512 (N_21512,N_21185,N_21236);
and U21513 (N_21513,N_20638,N_21079);
and U21514 (N_21514,N_20743,N_21226);
xnor U21515 (N_21515,N_20660,N_20859);
or U21516 (N_21516,N_20968,N_21064);
nor U21517 (N_21517,N_20847,N_20908);
xnor U21518 (N_21518,N_21053,N_20771);
nand U21519 (N_21519,N_21166,N_20892);
or U21520 (N_21520,N_20867,N_21061);
nor U21521 (N_21521,N_20708,N_20973);
or U21522 (N_21522,N_20925,N_20779);
nor U21523 (N_21523,N_20693,N_20858);
nor U21524 (N_21524,N_20658,N_20941);
or U21525 (N_21525,N_21231,N_20746);
and U21526 (N_21526,N_20887,N_20797);
nand U21527 (N_21527,N_20663,N_21033);
nor U21528 (N_21528,N_20976,N_20836);
nor U21529 (N_21529,N_21037,N_20837);
nand U21530 (N_21530,N_21179,N_21216);
nand U21531 (N_21531,N_21204,N_20692);
and U21532 (N_21532,N_20815,N_21214);
and U21533 (N_21533,N_21247,N_20665);
xnor U21534 (N_21534,N_20985,N_21139);
and U21535 (N_21535,N_20944,N_21171);
xor U21536 (N_21536,N_20798,N_21107);
nand U21537 (N_21537,N_20817,N_20789);
nand U21538 (N_21538,N_20807,N_20885);
and U21539 (N_21539,N_20895,N_21159);
nand U21540 (N_21540,N_21155,N_21035);
nand U21541 (N_21541,N_21198,N_20727);
nand U21542 (N_21542,N_20630,N_20775);
and U21543 (N_21543,N_20790,N_21194);
or U21544 (N_21544,N_21225,N_20763);
nor U21545 (N_21545,N_20717,N_20990);
nand U21546 (N_21546,N_20959,N_21157);
and U21547 (N_21547,N_20852,N_20871);
and U21548 (N_21548,N_20639,N_20783);
and U21549 (N_21549,N_20747,N_21106);
nand U21550 (N_21550,N_20761,N_21202);
nor U21551 (N_21551,N_21042,N_21072);
nand U21552 (N_21552,N_20755,N_20843);
or U21553 (N_21553,N_21038,N_20688);
or U21554 (N_21554,N_21218,N_20879);
xor U21555 (N_21555,N_20981,N_20880);
and U21556 (N_21556,N_20876,N_20701);
nor U21557 (N_21557,N_20907,N_20804);
nand U21558 (N_21558,N_21013,N_20932);
and U21559 (N_21559,N_20669,N_20931);
nand U21560 (N_21560,N_20770,N_20875);
xnor U21561 (N_21561,N_20950,N_20628);
xor U21562 (N_21562,N_21027,N_20674);
nor U21563 (N_21563,N_20748,N_20787);
nor U21564 (N_21564,N_20952,N_20959);
xor U21565 (N_21565,N_21037,N_20746);
nand U21566 (N_21566,N_20810,N_21011);
xor U21567 (N_21567,N_21130,N_21138);
nand U21568 (N_21568,N_20730,N_20770);
nand U21569 (N_21569,N_21059,N_20756);
or U21570 (N_21570,N_20878,N_20814);
or U21571 (N_21571,N_21052,N_21143);
xor U21572 (N_21572,N_21083,N_21202);
xnor U21573 (N_21573,N_21017,N_20751);
nand U21574 (N_21574,N_20860,N_20648);
nor U21575 (N_21575,N_20958,N_20646);
xor U21576 (N_21576,N_20848,N_20719);
or U21577 (N_21577,N_21031,N_20981);
xor U21578 (N_21578,N_21101,N_20888);
or U21579 (N_21579,N_20839,N_20878);
xnor U21580 (N_21580,N_20777,N_21193);
nand U21581 (N_21581,N_21151,N_20921);
and U21582 (N_21582,N_20956,N_21117);
xnor U21583 (N_21583,N_20905,N_20770);
xor U21584 (N_21584,N_20833,N_21103);
xor U21585 (N_21585,N_21088,N_21046);
nor U21586 (N_21586,N_20692,N_21043);
xnor U21587 (N_21587,N_20976,N_20864);
nor U21588 (N_21588,N_20772,N_20908);
nor U21589 (N_21589,N_20699,N_20910);
and U21590 (N_21590,N_21233,N_20677);
xor U21591 (N_21591,N_20765,N_20884);
and U21592 (N_21592,N_20695,N_21175);
and U21593 (N_21593,N_20761,N_20919);
nor U21594 (N_21594,N_21066,N_21045);
nor U21595 (N_21595,N_21020,N_20767);
nand U21596 (N_21596,N_20627,N_21213);
xnor U21597 (N_21597,N_21189,N_21114);
nand U21598 (N_21598,N_20802,N_21026);
xnor U21599 (N_21599,N_20778,N_20673);
or U21600 (N_21600,N_20781,N_20631);
nand U21601 (N_21601,N_20885,N_20675);
xnor U21602 (N_21602,N_20785,N_21015);
nand U21603 (N_21603,N_20954,N_20634);
nor U21604 (N_21604,N_20688,N_21244);
and U21605 (N_21605,N_21064,N_20744);
xor U21606 (N_21606,N_20693,N_20981);
nor U21607 (N_21607,N_20926,N_21084);
and U21608 (N_21608,N_20646,N_20746);
or U21609 (N_21609,N_20904,N_21095);
nand U21610 (N_21610,N_20665,N_20707);
or U21611 (N_21611,N_20845,N_21065);
xor U21612 (N_21612,N_21205,N_21111);
and U21613 (N_21613,N_21146,N_21129);
or U21614 (N_21614,N_20726,N_21243);
xor U21615 (N_21615,N_20925,N_21080);
nor U21616 (N_21616,N_20723,N_20916);
and U21617 (N_21617,N_21012,N_21214);
or U21618 (N_21618,N_20655,N_21035);
and U21619 (N_21619,N_20881,N_21201);
nor U21620 (N_21620,N_21131,N_20790);
and U21621 (N_21621,N_20892,N_21087);
nor U21622 (N_21622,N_21145,N_20694);
nor U21623 (N_21623,N_21049,N_20631);
nor U21624 (N_21624,N_21033,N_20667);
or U21625 (N_21625,N_20902,N_21235);
xor U21626 (N_21626,N_20994,N_20856);
nor U21627 (N_21627,N_20751,N_20649);
nor U21628 (N_21628,N_20872,N_20820);
xnor U21629 (N_21629,N_21170,N_21151);
nand U21630 (N_21630,N_20853,N_20931);
nor U21631 (N_21631,N_20729,N_20898);
xor U21632 (N_21632,N_21027,N_21096);
or U21633 (N_21633,N_21075,N_21055);
nor U21634 (N_21634,N_20690,N_20672);
or U21635 (N_21635,N_21122,N_21071);
or U21636 (N_21636,N_20979,N_21221);
nand U21637 (N_21637,N_21014,N_21009);
nand U21638 (N_21638,N_20901,N_20832);
xnor U21639 (N_21639,N_21118,N_20753);
or U21640 (N_21640,N_20855,N_21158);
xor U21641 (N_21641,N_20938,N_21227);
or U21642 (N_21642,N_20727,N_20732);
nor U21643 (N_21643,N_21113,N_20703);
nor U21644 (N_21644,N_20737,N_20794);
or U21645 (N_21645,N_20842,N_21124);
nand U21646 (N_21646,N_21002,N_21237);
nor U21647 (N_21647,N_20737,N_20830);
nor U21648 (N_21648,N_20852,N_20987);
nand U21649 (N_21649,N_20631,N_20910);
and U21650 (N_21650,N_21094,N_21127);
and U21651 (N_21651,N_20948,N_20976);
or U21652 (N_21652,N_20717,N_20732);
nand U21653 (N_21653,N_20692,N_21014);
and U21654 (N_21654,N_20878,N_21111);
nor U21655 (N_21655,N_20781,N_21186);
nor U21656 (N_21656,N_21175,N_20975);
nand U21657 (N_21657,N_21144,N_21168);
and U21658 (N_21658,N_20685,N_20797);
xor U21659 (N_21659,N_20878,N_21024);
nand U21660 (N_21660,N_20706,N_20927);
nor U21661 (N_21661,N_21164,N_20838);
nand U21662 (N_21662,N_21021,N_20654);
nand U21663 (N_21663,N_21168,N_20941);
nand U21664 (N_21664,N_21052,N_20814);
nand U21665 (N_21665,N_21086,N_20833);
and U21666 (N_21666,N_20776,N_20634);
or U21667 (N_21667,N_20693,N_21148);
nand U21668 (N_21668,N_21184,N_21194);
nor U21669 (N_21669,N_20658,N_20882);
and U21670 (N_21670,N_20754,N_20692);
or U21671 (N_21671,N_20743,N_20651);
nor U21672 (N_21672,N_20906,N_20949);
or U21673 (N_21673,N_21229,N_20980);
xnor U21674 (N_21674,N_20979,N_20753);
xnor U21675 (N_21675,N_21160,N_21150);
nand U21676 (N_21676,N_20833,N_20913);
nor U21677 (N_21677,N_20680,N_21061);
xor U21678 (N_21678,N_21109,N_21067);
nand U21679 (N_21679,N_20901,N_20740);
nand U21680 (N_21680,N_20740,N_20724);
xnor U21681 (N_21681,N_20897,N_21077);
nor U21682 (N_21682,N_20879,N_21051);
xor U21683 (N_21683,N_20946,N_20714);
nand U21684 (N_21684,N_21062,N_20682);
or U21685 (N_21685,N_20860,N_20692);
xor U21686 (N_21686,N_21193,N_21145);
xnor U21687 (N_21687,N_20882,N_20890);
or U21688 (N_21688,N_20807,N_21060);
or U21689 (N_21689,N_20768,N_20944);
xor U21690 (N_21690,N_20855,N_20870);
xnor U21691 (N_21691,N_21127,N_21076);
nor U21692 (N_21692,N_21072,N_21041);
or U21693 (N_21693,N_21205,N_20964);
or U21694 (N_21694,N_21241,N_21084);
or U21695 (N_21695,N_20965,N_21188);
nor U21696 (N_21696,N_21002,N_21080);
xnor U21697 (N_21697,N_20739,N_20908);
nor U21698 (N_21698,N_20651,N_20644);
nor U21699 (N_21699,N_20752,N_20832);
nor U21700 (N_21700,N_20855,N_20935);
and U21701 (N_21701,N_20695,N_21096);
nand U21702 (N_21702,N_20716,N_20919);
xor U21703 (N_21703,N_20678,N_20771);
nor U21704 (N_21704,N_20831,N_20974);
nand U21705 (N_21705,N_21049,N_20766);
xnor U21706 (N_21706,N_20671,N_20628);
nand U21707 (N_21707,N_21063,N_21228);
and U21708 (N_21708,N_21140,N_20697);
xnor U21709 (N_21709,N_21055,N_21028);
nor U21710 (N_21710,N_21038,N_20861);
nor U21711 (N_21711,N_21107,N_20705);
nor U21712 (N_21712,N_20818,N_21065);
xnor U21713 (N_21713,N_20978,N_20711);
nand U21714 (N_21714,N_21092,N_20904);
and U21715 (N_21715,N_21073,N_20645);
nor U21716 (N_21716,N_20818,N_20846);
and U21717 (N_21717,N_20744,N_20816);
nor U21718 (N_21718,N_21035,N_21080);
xnor U21719 (N_21719,N_21178,N_20970);
xnor U21720 (N_21720,N_20965,N_21039);
xor U21721 (N_21721,N_21056,N_21167);
nor U21722 (N_21722,N_21022,N_20911);
nand U21723 (N_21723,N_20742,N_20721);
xor U21724 (N_21724,N_21036,N_21076);
nand U21725 (N_21725,N_21241,N_20700);
or U21726 (N_21726,N_20812,N_20858);
and U21727 (N_21727,N_20774,N_20675);
nor U21728 (N_21728,N_21066,N_21065);
and U21729 (N_21729,N_21220,N_21106);
or U21730 (N_21730,N_21234,N_20773);
and U21731 (N_21731,N_21007,N_20883);
nand U21732 (N_21732,N_21113,N_20912);
xor U21733 (N_21733,N_21196,N_20799);
xor U21734 (N_21734,N_20871,N_20727);
xnor U21735 (N_21735,N_21247,N_20667);
nor U21736 (N_21736,N_21132,N_20997);
nor U21737 (N_21737,N_21218,N_20742);
nor U21738 (N_21738,N_20989,N_21052);
xnor U21739 (N_21739,N_20914,N_20646);
nand U21740 (N_21740,N_20725,N_20859);
or U21741 (N_21741,N_21146,N_20964);
nor U21742 (N_21742,N_20677,N_20742);
xnor U21743 (N_21743,N_21075,N_20744);
or U21744 (N_21744,N_21005,N_21022);
nand U21745 (N_21745,N_21042,N_20898);
nand U21746 (N_21746,N_20852,N_21029);
and U21747 (N_21747,N_20822,N_20779);
xnor U21748 (N_21748,N_21019,N_21238);
and U21749 (N_21749,N_20890,N_21004);
nor U21750 (N_21750,N_20865,N_21216);
nor U21751 (N_21751,N_20926,N_21082);
and U21752 (N_21752,N_20941,N_21116);
or U21753 (N_21753,N_20777,N_20764);
or U21754 (N_21754,N_21175,N_21129);
and U21755 (N_21755,N_20978,N_20886);
nand U21756 (N_21756,N_20782,N_21069);
xor U21757 (N_21757,N_20772,N_20834);
xor U21758 (N_21758,N_21000,N_21215);
and U21759 (N_21759,N_20627,N_20962);
and U21760 (N_21760,N_20699,N_21127);
or U21761 (N_21761,N_21108,N_21043);
nand U21762 (N_21762,N_21238,N_20789);
nand U21763 (N_21763,N_21009,N_20966);
or U21764 (N_21764,N_20747,N_20863);
xor U21765 (N_21765,N_21118,N_20835);
xor U21766 (N_21766,N_20641,N_20838);
or U21767 (N_21767,N_20717,N_21151);
nand U21768 (N_21768,N_20999,N_20864);
or U21769 (N_21769,N_20887,N_20834);
nor U21770 (N_21770,N_20819,N_21169);
or U21771 (N_21771,N_20709,N_20963);
nor U21772 (N_21772,N_21109,N_21192);
nor U21773 (N_21773,N_20855,N_20671);
or U21774 (N_21774,N_20752,N_21085);
xor U21775 (N_21775,N_20783,N_20893);
or U21776 (N_21776,N_20773,N_21155);
xor U21777 (N_21777,N_20929,N_20708);
nand U21778 (N_21778,N_20746,N_20627);
xor U21779 (N_21779,N_20923,N_21124);
nand U21780 (N_21780,N_20739,N_20840);
xnor U21781 (N_21781,N_20973,N_20831);
xnor U21782 (N_21782,N_21074,N_21170);
nand U21783 (N_21783,N_20652,N_21051);
or U21784 (N_21784,N_21113,N_21095);
and U21785 (N_21785,N_20772,N_21139);
nand U21786 (N_21786,N_21087,N_20648);
and U21787 (N_21787,N_20933,N_20787);
xor U21788 (N_21788,N_20702,N_20986);
or U21789 (N_21789,N_20838,N_20805);
nand U21790 (N_21790,N_20852,N_20654);
nand U21791 (N_21791,N_20750,N_20972);
xor U21792 (N_21792,N_20755,N_20816);
xor U21793 (N_21793,N_20810,N_21171);
nand U21794 (N_21794,N_20842,N_20670);
or U21795 (N_21795,N_20761,N_20650);
xnor U21796 (N_21796,N_21232,N_20714);
xnor U21797 (N_21797,N_21080,N_20732);
nand U21798 (N_21798,N_20766,N_20926);
or U21799 (N_21799,N_21240,N_20697);
or U21800 (N_21800,N_21126,N_21128);
xor U21801 (N_21801,N_20960,N_20783);
xnor U21802 (N_21802,N_21192,N_20717);
xnor U21803 (N_21803,N_20760,N_20765);
xor U21804 (N_21804,N_21115,N_20943);
or U21805 (N_21805,N_20649,N_21072);
nor U21806 (N_21806,N_21056,N_20935);
xnor U21807 (N_21807,N_20760,N_20925);
and U21808 (N_21808,N_20651,N_20714);
nor U21809 (N_21809,N_20829,N_21079);
xnor U21810 (N_21810,N_20940,N_20900);
and U21811 (N_21811,N_20711,N_20739);
or U21812 (N_21812,N_20764,N_20927);
and U21813 (N_21813,N_20836,N_21087);
and U21814 (N_21814,N_21128,N_21249);
and U21815 (N_21815,N_20929,N_21130);
nand U21816 (N_21816,N_20773,N_20880);
or U21817 (N_21817,N_20626,N_20927);
nor U21818 (N_21818,N_20752,N_20962);
or U21819 (N_21819,N_20981,N_20660);
xnor U21820 (N_21820,N_20828,N_21185);
or U21821 (N_21821,N_20945,N_20858);
and U21822 (N_21822,N_21152,N_21122);
nor U21823 (N_21823,N_20918,N_20763);
nand U21824 (N_21824,N_21085,N_20896);
nor U21825 (N_21825,N_20678,N_21173);
xnor U21826 (N_21826,N_21107,N_20788);
nor U21827 (N_21827,N_20890,N_20690);
or U21828 (N_21828,N_20692,N_20832);
or U21829 (N_21829,N_21054,N_20780);
and U21830 (N_21830,N_20898,N_20920);
or U21831 (N_21831,N_20949,N_20705);
and U21832 (N_21832,N_20689,N_20964);
nor U21833 (N_21833,N_21119,N_20715);
or U21834 (N_21834,N_20960,N_21230);
xor U21835 (N_21835,N_21112,N_20830);
xnor U21836 (N_21836,N_21048,N_21065);
and U21837 (N_21837,N_20814,N_20668);
or U21838 (N_21838,N_21023,N_20863);
nand U21839 (N_21839,N_20902,N_20787);
nor U21840 (N_21840,N_20660,N_21015);
and U21841 (N_21841,N_21176,N_20924);
nand U21842 (N_21842,N_20834,N_21017);
xor U21843 (N_21843,N_21118,N_21249);
nand U21844 (N_21844,N_21062,N_21161);
nand U21845 (N_21845,N_20811,N_21017);
nand U21846 (N_21846,N_21077,N_20702);
nor U21847 (N_21847,N_20640,N_20826);
nand U21848 (N_21848,N_20886,N_20625);
or U21849 (N_21849,N_20786,N_20639);
nand U21850 (N_21850,N_21091,N_21243);
xor U21851 (N_21851,N_20914,N_21112);
and U21852 (N_21852,N_20775,N_20637);
and U21853 (N_21853,N_20668,N_20917);
or U21854 (N_21854,N_20688,N_21163);
and U21855 (N_21855,N_21026,N_21189);
nand U21856 (N_21856,N_21024,N_20686);
nand U21857 (N_21857,N_20692,N_20823);
nand U21858 (N_21858,N_20736,N_21248);
nand U21859 (N_21859,N_20649,N_20829);
nand U21860 (N_21860,N_20884,N_20776);
nand U21861 (N_21861,N_20663,N_21174);
nand U21862 (N_21862,N_20921,N_21143);
or U21863 (N_21863,N_20670,N_21224);
and U21864 (N_21864,N_20947,N_21168);
nor U21865 (N_21865,N_20639,N_20697);
or U21866 (N_21866,N_21137,N_21031);
nor U21867 (N_21867,N_20935,N_20911);
or U21868 (N_21868,N_21129,N_20749);
nand U21869 (N_21869,N_20688,N_21007);
and U21870 (N_21870,N_20632,N_21136);
or U21871 (N_21871,N_20654,N_20740);
or U21872 (N_21872,N_21206,N_20809);
nand U21873 (N_21873,N_21024,N_21060);
nor U21874 (N_21874,N_21120,N_20861);
or U21875 (N_21875,N_21668,N_21529);
xnor U21876 (N_21876,N_21686,N_21331);
nor U21877 (N_21877,N_21637,N_21583);
and U21878 (N_21878,N_21791,N_21417);
nand U21879 (N_21879,N_21850,N_21253);
nor U21880 (N_21880,N_21636,N_21369);
xnor U21881 (N_21881,N_21391,N_21265);
or U21882 (N_21882,N_21344,N_21804);
and U21883 (N_21883,N_21345,N_21749);
or U21884 (N_21884,N_21267,N_21298);
nor U21885 (N_21885,N_21680,N_21666);
and U21886 (N_21886,N_21523,N_21468);
nand U21887 (N_21887,N_21827,N_21752);
or U21888 (N_21888,N_21574,N_21536);
nor U21889 (N_21889,N_21742,N_21792);
xnor U21890 (N_21890,N_21593,N_21826);
or U21891 (N_21891,N_21712,N_21720);
nand U21892 (N_21892,N_21403,N_21342);
nand U21893 (N_21893,N_21348,N_21415);
nor U21894 (N_21894,N_21589,N_21546);
nor U21895 (N_21895,N_21856,N_21643);
and U21896 (N_21896,N_21553,N_21429);
and U21897 (N_21897,N_21765,N_21829);
or U21898 (N_21898,N_21616,N_21721);
nand U21899 (N_21899,N_21484,N_21469);
nor U21900 (N_21900,N_21295,N_21596);
and U21901 (N_21901,N_21754,N_21423);
and U21902 (N_21902,N_21603,N_21520);
nand U21903 (N_21903,N_21266,N_21702);
or U21904 (N_21904,N_21602,N_21800);
and U21905 (N_21905,N_21674,N_21845);
nor U21906 (N_21906,N_21388,N_21554);
and U21907 (N_21907,N_21573,N_21504);
or U21908 (N_21908,N_21870,N_21635);
nand U21909 (N_21909,N_21544,N_21435);
nor U21910 (N_21910,N_21537,N_21491);
and U21911 (N_21911,N_21700,N_21328);
nor U21912 (N_21912,N_21625,N_21412);
nand U21913 (N_21913,N_21698,N_21381);
xnor U21914 (N_21914,N_21492,N_21681);
xnor U21915 (N_21915,N_21785,N_21379);
nor U21916 (N_21916,N_21356,N_21640);
or U21917 (N_21917,N_21578,N_21839);
nand U21918 (N_21918,N_21313,N_21287);
or U21919 (N_21919,N_21495,N_21542);
nand U21920 (N_21920,N_21746,N_21658);
nand U21921 (N_21921,N_21263,N_21694);
or U21922 (N_21922,N_21866,N_21816);
and U21923 (N_21923,N_21372,N_21591);
nand U21924 (N_21924,N_21463,N_21617);
and U21925 (N_21925,N_21599,N_21517);
nor U21926 (N_21926,N_21564,N_21652);
or U21927 (N_21927,N_21766,N_21418);
nor U21928 (N_21928,N_21286,N_21366);
or U21929 (N_21929,N_21789,N_21446);
nand U21930 (N_21930,N_21319,N_21270);
and U21931 (N_21931,N_21424,N_21704);
xnor U21932 (N_21932,N_21790,N_21659);
xnor U21933 (N_21933,N_21844,N_21292);
nand U21934 (N_21934,N_21683,N_21330);
or U21935 (N_21935,N_21701,N_21459);
nor U21936 (N_21936,N_21695,N_21571);
xnor U21937 (N_21937,N_21586,N_21824);
xnor U21938 (N_21938,N_21868,N_21370);
nand U21939 (N_21939,N_21610,N_21736);
nor U21940 (N_21940,N_21281,N_21312);
nor U21941 (N_21941,N_21663,N_21503);
nor U21942 (N_21942,N_21540,N_21541);
xor U21943 (N_21943,N_21394,N_21709);
or U21944 (N_21944,N_21706,N_21732);
or U21945 (N_21945,N_21615,N_21814);
and U21946 (N_21946,N_21279,N_21645);
nor U21947 (N_21947,N_21285,N_21632);
and U21948 (N_21948,N_21724,N_21289);
nand U21949 (N_21949,N_21641,N_21430);
or U21950 (N_21950,N_21773,N_21399);
nand U21951 (N_21951,N_21561,N_21427);
xnor U21952 (N_21952,N_21303,N_21329);
nor U21953 (N_21953,N_21408,N_21558);
or U21954 (N_21954,N_21605,N_21679);
and U21955 (N_21955,N_21453,N_21487);
and U21956 (N_21956,N_21299,N_21664);
or U21957 (N_21957,N_21860,N_21449);
nor U21958 (N_21958,N_21481,N_21690);
nor U21959 (N_21959,N_21339,N_21414);
nand U21960 (N_21960,N_21264,N_21568);
xnor U21961 (N_21961,N_21456,N_21570);
xnor U21962 (N_21962,N_21304,N_21556);
nor U21963 (N_21963,N_21361,N_21387);
nor U21964 (N_21964,N_21390,N_21822);
nand U21965 (N_21965,N_21563,N_21751);
or U21966 (N_21966,N_21691,N_21318);
xnor U21967 (N_21967,N_21707,N_21806);
nand U21968 (N_21968,N_21606,N_21256);
nor U21969 (N_21969,N_21572,N_21472);
nand U21970 (N_21970,N_21715,N_21257);
and U21971 (N_21971,N_21815,N_21421);
and U21972 (N_21972,N_21848,N_21431);
nor U21973 (N_21973,N_21741,N_21618);
nor U21974 (N_21974,N_21714,N_21364);
nand U21975 (N_21975,N_21823,N_21750);
xor U21976 (N_21976,N_21708,N_21581);
or U21977 (N_21977,N_21857,N_21522);
and U21978 (N_21978,N_21629,N_21598);
and U21979 (N_21979,N_21585,N_21667);
or U21980 (N_21980,N_21505,N_21350);
nand U21981 (N_21981,N_21808,N_21478);
xnor U21982 (N_21982,N_21722,N_21547);
or U21983 (N_21983,N_21461,N_21307);
nand U21984 (N_21984,N_21382,N_21803);
or U21985 (N_21985,N_21252,N_21510);
or U21986 (N_21986,N_21833,N_21644);
and U21987 (N_21987,N_21254,N_21349);
or U21988 (N_21988,N_21550,N_21675);
nor U21989 (N_21989,N_21689,N_21498);
nor U21990 (N_21990,N_21305,N_21863);
or U21991 (N_21991,N_21768,N_21282);
or U21992 (N_21992,N_21314,N_21828);
or U21993 (N_21993,N_21405,N_21273);
xor U21994 (N_21994,N_21802,N_21549);
and U21995 (N_21995,N_21384,N_21569);
or U21996 (N_21996,N_21419,N_21502);
nor U21997 (N_21997,N_21486,N_21797);
or U21998 (N_21998,N_21255,N_21728);
nor U21999 (N_21999,N_21796,N_21716);
nand U22000 (N_22000,N_21682,N_21335);
and U22001 (N_22001,N_21718,N_21843);
xnor U22002 (N_22002,N_21801,N_21788);
nand U22003 (N_22003,N_21539,N_21406);
nand U22004 (N_22004,N_21422,N_21493);
or U22005 (N_22005,N_21723,N_21525);
xor U22006 (N_22006,N_21853,N_21466);
nor U22007 (N_22007,N_21783,N_21250);
nor U22008 (N_22008,N_21385,N_21473);
and U22009 (N_22009,N_21464,N_21509);
nand U22010 (N_22010,N_21836,N_21867);
or U22011 (N_22011,N_21496,N_21395);
nand U22012 (N_22012,N_21308,N_21793);
nor U22013 (N_22013,N_21410,N_21315);
and U22014 (N_22014,N_21297,N_21460);
nand U22015 (N_22015,N_21326,N_21368);
and U22016 (N_22016,N_21398,N_21347);
or U22017 (N_22017,N_21874,N_21518);
or U22018 (N_22018,N_21759,N_21321);
nand U22019 (N_22019,N_21499,N_21677);
nand U22020 (N_22020,N_21743,N_21411);
or U22021 (N_22021,N_21609,N_21393);
and U22022 (N_22022,N_21514,N_21837);
nor U22023 (N_22023,N_21590,N_21819);
xor U22024 (N_22024,N_21450,N_21438);
nand U22025 (N_22025,N_21726,N_21780);
nor U22026 (N_22026,N_21727,N_21811);
nor U22027 (N_22027,N_21620,N_21374);
or U22028 (N_22028,N_21653,N_21705);
nor U22029 (N_22029,N_21807,N_21784);
and U22030 (N_22030,N_21872,N_21357);
nor U22031 (N_22031,N_21283,N_21662);
and U22032 (N_22032,N_21745,N_21275);
xor U22033 (N_22033,N_21696,N_21612);
nand U22034 (N_22034,N_21434,N_21389);
nor U22035 (N_22035,N_21258,N_21650);
nor U22036 (N_22036,N_21734,N_21291);
nand U22037 (N_22037,N_21762,N_21300);
and U22038 (N_22038,N_21482,N_21656);
or U22039 (N_22039,N_21738,N_21655);
nor U22040 (N_22040,N_21642,N_21634);
and U22041 (N_22041,N_21565,N_21407);
xnor U22042 (N_22042,N_21601,N_21302);
or U22043 (N_22043,N_21757,N_21392);
nand U22044 (N_22044,N_21756,N_21306);
xor U22045 (N_22045,N_21772,N_21343);
and U22046 (N_22046,N_21622,N_21584);
xnor U22047 (N_22047,N_21862,N_21794);
nand U22048 (N_22048,N_21530,N_21771);
and U22049 (N_22049,N_21293,N_21864);
nand U22050 (N_22050,N_21769,N_21760);
nand U22051 (N_22051,N_21351,N_21594);
and U22052 (N_22052,N_21671,N_21755);
and U22053 (N_22053,N_21735,N_21559);
or U22054 (N_22054,N_21770,N_21334);
nor U22055 (N_22055,N_21621,N_21508);
and U22056 (N_22056,N_21810,N_21521);
nor U22057 (N_22057,N_21851,N_21692);
and U22058 (N_22058,N_21327,N_21432);
xor U22059 (N_22059,N_21404,N_21336);
and U22060 (N_22060,N_21433,N_21355);
or U22061 (N_22061,N_21873,N_21767);
nor U22062 (N_22062,N_21847,N_21488);
or U22063 (N_22063,N_21623,N_21480);
nand U22064 (N_22064,N_21676,N_21619);
nor U22065 (N_22065,N_21274,N_21363);
or U22066 (N_22066,N_21462,N_21665);
or U22067 (N_22067,N_21557,N_21323);
or U22068 (N_22068,N_21448,N_21776);
nor U22069 (N_22069,N_21513,N_21841);
nand U22070 (N_22070,N_21575,N_21608);
nor U22071 (N_22071,N_21562,N_21805);
or U22072 (N_22072,N_21582,N_21470);
nand U22073 (N_22073,N_21346,N_21485);
or U22074 (N_22074,N_21373,N_21775);
or U22075 (N_22075,N_21251,N_21567);
or U22076 (N_22076,N_21296,N_21744);
xor U22077 (N_22077,N_21380,N_21719);
xnor U22078 (N_22078,N_21442,N_21693);
xnor U22079 (N_22079,N_21638,N_21260);
and U22080 (N_22080,N_21465,N_21731);
or U22081 (N_22081,N_21436,N_21383);
and U22082 (N_22082,N_21428,N_21628);
and U22083 (N_22083,N_21661,N_21786);
nand U22084 (N_22084,N_21507,N_21301);
xnor U22085 (N_22085,N_21376,N_21820);
xor U22086 (N_22086,N_21511,N_21580);
nor U22087 (N_22087,N_21842,N_21284);
or U22088 (N_22088,N_21604,N_21579);
xnor U22089 (N_22089,N_21340,N_21577);
and U22090 (N_22090,N_21400,N_21798);
nand U22091 (N_22091,N_21479,N_21276);
or U22092 (N_22092,N_21871,N_21758);
nand U22093 (N_22093,N_21576,N_21277);
or U22094 (N_22094,N_21402,N_21633);
nor U22095 (N_22095,N_21262,N_21725);
or U22096 (N_22096,N_21533,N_21458);
xor U22097 (N_22097,N_21795,N_21821);
xnor U22098 (N_22098,N_21648,N_21474);
and U22099 (N_22099,N_21316,N_21774);
and U22100 (N_22100,N_21812,N_21288);
and U22101 (N_22101,N_21528,N_21455);
or U22102 (N_22102,N_21861,N_21830);
or U22103 (N_22103,N_21747,N_21386);
nand U22104 (N_22104,N_21475,N_21371);
or U22105 (N_22105,N_21451,N_21437);
xor U22106 (N_22106,N_21516,N_21678);
nand U22107 (N_22107,N_21699,N_21268);
nand U22108 (N_22108,N_21501,N_21778);
and U22109 (N_22109,N_21259,N_21278);
xnor U22110 (N_22110,N_21269,N_21443);
and U22111 (N_22111,N_21684,N_21338);
xor U22112 (N_22112,N_21809,N_21838);
nor U22113 (N_22113,N_21365,N_21855);
and U22114 (N_22114,N_21748,N_21739);
xor U22115 (N_22115,N_21654,N_21627);
nor U22116 (N_22116,N_21818,N_21595);
nor U22117 (N_22117,N_21717,N_21761);
nand U22118 (N_22118,N_21697,N_21534);
xnor U22119 (N_22119,N_21703,N_21729);
and U22120 (N_22120,N_21500,N_21813);
xor U22121 (N_22121,N_21832,N_21865);
and U22122 (N_22122,N_21280,N_21753);
nand U22123 (N_22123,N_21733,N_21614);
nor U22124 (N_22124,N_21560,N_21597);
and U22125 (N_22125,N_21613,N_21825);
nor U22126 (N_22126,N_21730,N_21272);
nand U22127 (N_22127,N_21854,N_21490);
or U22128 (N_22128,N_21489,N_21763);
nand U22129 (N_22129,N_21713,N_21631);
nand U22130 (N_22130,N_21324,N_21483);
nor U22131 (N_22131,N_21846,N_21362);
xor U22132 (N_22132,N_21647,N_21333);
xor U22133 (N_22133,N_21588,N_21454);
xnor U22134 (N_22134,N_21271,N_21452);
xnor U22135 (N_22135,N_21543,N_21869);
nand U22136 (N_22136,N_21587,N_21425);
or U22137 (N_22137,N_21685,N_21261);
and U22138 (N_22138,N_21600,N_21515);
or U22139 (N_22139,N_21859,N_21317);
nand U22140 (N_22140,N_21710,N_21607);
xor U22141 (N_22141,N_21378,N_21782);
nand U22142 (N_22142,N_21440,N_21592);
nand U22143 (N_22143,N_21441,N_21524);
nor U22144 (N_22144,N_21512,N_21341);
xor U22145 (N_22145,N_21737,N_21416);
xor U22146 (N_22146,N_21396,N_21467);
nor U22147 (N_22147,N_21626,N_21624);
and U22148 (N_22148,N_21294,N_21360);
nand U22149 (N_22149,N_21444,N_21552);
and U22150 (N_22150,N_21840,N_21477);
nor U22151 (N_22151,N_21651,N_21781);
xor U22152 (N_22152,N_21377,N_21457);
nor U22153 (N_22153,N_21311,N_21354);
and U22154 (N_22154,N_21413,N_21310);
and U22155 (N_22155,N_21367,N_21657);
nor U22156 (N_22156,N_21777,N_21669);
xnor U22157 (N_22157,N_21538,N_21353);
nand U22158 (N_22158,N_21611,N_21787);
or U22159 (N_22159,N_21325,N_21630);
and U22160 (N_22160,N_21834,N_21526);
nand U22161 (N_22161,N_21849,N_21639);
and U22162 (N_22162,N_21476,N_21858);
nand U22163 (N_22163,N_21426,N_21337);
nor U22164 (N_22164,N_21497,N_21551);
nor U22165 (N_22165,N_21670,N_21320);
and U22166 (N_22166,N_21447,N_21660);
and U22167 (N_22167,N_21835,N_21401);
or U22168 (N_22168,N_21409,N_21740);
or U22169 (N_22169,N_21352,N_21687);
or U22170 (N_22170,N_21445,N_21852);
nand U22171 (N_22171,N_21817,N_21358);
and U22172 (N_22172,N_21673,N_21322);
or U22173 (N_22173,N_21359,N_21779);
nor U22174 (N_22174,N_21375,N_21646);
or U22175 (N_22175,N_21420,N_21535);
xor U22176 (N_22176,N_21555,N_21548);
or U22177 (N_22177,N_21672,N_21290);
nand U22178 (N_22178,N_21545,N_21711);
nor U22179 (N_22179,N_21309,N_21527);
xnor U22180 (N_22180,N_21506,N_21649);
nor U22181 (N_22181,N_21332,N_21532);
xnor U22182 (N_22182,N_21688,N_21397);
xnor U22183 (N_22183,N_21831,N_21764);
or U22184 (N_22184,N_21471,N_21531);
or U22185 (N_22185,N_21494,N_21799);
or U22186 (N_22186,N_21519,N_21439);
xor U22187 (N_22187,N_21566,N_21591);
and U22188 (N_22188,N_21744,N_21726);
xnor U22189 (N_22189,N_21397,N_21386);
xnor U22190 (N_22190,N_21854,N_21317);
xor U22191 (N_22191,N_21734,N_21613);
nor U22192 (N_22192,N_21443,N_21606);
xor U22193 (N_22193,N_21428,N_21790);
nor U22194 (N_22194,N_21381,N_21845);
or U22195 (N_22195,N_21474,N_21693);
nand U22196 (N_22196,N_21297,N_21389);
and U22197 (N_22197,N_21388,N_21640);
or U22198 (N_22198,N_21576,N_21512);
and U22199 (N_22199,N_21390,N_21465);
nor U22200 (N_22200,N_21635,N_21713);
xnor U22201 (N_22201,N_21760,N_21744);
nand U22202 (N_22202,N_21414,N_21518);
xnor U22203 (N_22203,N_21743,N_21293);
or U22204 (N_22204,N_21313,N_21840);
or U22205 (N_22205,N_21818,N_21871);
or U22206 (N_22206,N_21354,N_21651);
nor U22207 (N_22207,N_21465,N_21344);
nor U22208 (N_22208,N_21833,N_21516);
nor U22209 (N_22209,N_21274,N_21829);
xnor U22210 (N_22210,N_21651,N_21871);
xor U22211 (N_22211,N_21759,N_21527);
xnor U22212 (N_22212,N_21597,N_21766);
xnor U22213 (N_22213,N_21643,N_21268);
and U22214 (N_22214,N_21325,N_21316);
xor U22215 (N_22215,N_21752,N_21736);
nand U22216 (N_22216,N_21394,N_21413);
xor U22217 (N_22217,N_21451,N_21827);
xnor U22218 (N_22218,N_21772,N_21696);
or U22219 (N_22219,N_21355,N_21790);
nand U22220 (N_22220,N_21356,N_21613);
or U22221 (N_22221,N_21516,N_21738);
nand U22222 (N_22222,N_21821,N_21780);
or U22223 (N_22223,N_21357,N_21454);
nor U22224 (N_22224,N_21393,N_21441);
xnor U22225 (N_22225,N_21582,N_21308);
nor U22226 (N_22226,N_21359,N_21489);
or U22227 (N_22227,N_21345,N_21684);
or U22228 (N_22228,N_21813,N_21414);
and U22229 (N_22229,N_21313,N_21389);
or U22230 (N_22230,N_21312,N_21348);
xnor U22231 (N_22231,N_21491,N_21760);
and U22232 (N_22232,N_21416,N_21446);
or U22233 (N_22233,N_21360,N_21434);
and U22234 (N_22234,N_21328,N_21783);
and U22235 (N_22235,N_21579,N_21315);
and U22236 (N_22236,N_21548,N_21825);
xnor U22237 (N_22237,N_21420,N_21385);
xnor U22238 (N_22238,N_21520,N_21684);
or U22239 (N_22239,N_21775,N_21597);
xor U22240 (N_22240,N_21710,N_21849);
nor U22241 (N_22241,N_21271,N_21451);
or U22242 (N_22242,N_21525,N_21589);
xnor U22243 (N_22243,N_21310,N_21403);
or U22244 (N_22244,N_21852,N_21257);
xnor U22245 (N_22245,N_21641,N_21844);
and U22246 (N_22246,N_21725,N_21469);
nor U22247 (N_22247,N_21631,N_21422);
or U22248 (N_22248,N_21661,N_21266);
nor U22249 (N_22249,N_21562,N_21750);
and U22250 (N_22250,N_21340,N_21256);
nor U22251 (N_22251,N_21659,N_21699);
nand U22252 (N_22252,N_21713,N_21821);
nor U22253 (N_22253,N_21560,N_21825);
and U22254 (N_22254,N_21656,N_21477);
and U22255 (N_22255,N_21774,N_21814);
nor U22256 (N_22256,N_21378,N_21265);
nor U22257 (N_22257,N_21263,N_21421);
and U22258 (N_22258,N_21294,N_21725);
xnor U22259 (N_22259,N_21596,N_21765);
nand U22260 (N_22260,N_21693,N_21259);
and U22261 (N_22261,N_21756,N_21588);
and U22262 (N_22262,N_21499,N_21710);
nand U22263 (N_22263,N_21263,N_21484);
nor U22264 (N_22264,N_21336,N_21615);
and U22265 (N_22265,N_21785,N_21536);
nand U22266 (N_22266,N_21874,N_21351);
or U22267 (N_22267,N_21763,N_21599);
nor U22268 (N_22268,N_21441,N_21553);
xnor U22269 (N_22269,N_21252,N_21722);
xnor U22270 (N_22270,N_21756,N_21707);
nand U22271 (N_22271,N_21561,N_21870);
nand U22272 (N_22272,N_21732,N_21445);
or U22273 (N_22273,N_21319,N_21774);
or U22274 (N_22274,N_21392,N_21793);
or U22275 (N_22275,N_21678,N_21357);
nor U22276 (N_22276,N_21441,N_21492);
nor U22277 (N_22277,N_21669,N_21590);
nand U22278 (N_22278,N_21355,N_21867);
nand U22279 (N_22279,N_21694,N_21630);
nor U22280 (N_22280,N_21332,N_21344);
nand U22281 (N_22281,N_21840,N_21432);
and U22282 (N_22282,N_21665,N_21783);
nand U22283 (N_22283,N_21730,N_21348);
nand U22284 (N_22284,N_21711,N_21610);
or U22285 (N_22285,N_21462,N_21269);
nand U22286 (N_22286,N_21440,N_21588);
xnor U22287 (N_22287,N_21376,N_21789);
or U22288 (N_22288,N_21574,N_21819);
or U22289 (N_22289,N_21533,N_21739);
xor U22290 (N_22290,N_21362,N_21844);
xnor U22291 (N_22291,N_21586,N_21636);
nor U22292 (N_22292,N_21378,N_21831);
nand U22293 (N_22293,N_21539,N_21586);
and U22294 (N_22294,N_21717,N_21416);
nand U22295 (N_22295,N_21271,N_21408);
nand U22296 (N_22296,N_21574,N_21519);
and U22297 (N_22297,N_21840,N_21763);
nand U22298 (N_22298,N_21572,N_21769);
and U22299 (N_22299,N_21372,N_21367);
and U22300 (N_22300,N_21522,N_21814);
and U22301 (N_22301,N_21609,N_21866);
nor U22302 (N_22302,N_21267,N_21273);
and U22303 (N_22303,N_21370,N_21319);
or U22304 (N_22304,N_21728,N_21777);
nand U22305 (N_22305,N_21739,N_21528);
or U22306 (N_22306,N_21702,N_21631);
and U22307 (N_22307,N_21665,N_21376);
xnor U22308 (N_22308,N_21294,N_21461);
or U22309 (N_22309,N_21818,N_21752);
xor U22310 (N_22310,N_21458,N_21869);
xor U22311 (N_22311,N_21817,N_21607);
and U22312 (N_22312,N_21701,N_21491);
or U22313 (N_22313,N_21846,N_21722);
nor U22314 (N_22314,N_21518,N_21593);
and U22315 (N_22315,N_21389,N_21292);
and U22316 (N_22316,N_21386,N_21656);
nand U22317 (N_22317,N_21302,N_21496);
nand U22318 (N_22318,N_21626,N_21349);
and U22319 (N_22319,N_21528,N_21333);
xor U22320 (N_22320,N_21345,N_21304);
nand U22321 (N_22321,N_21589,N_21660);
xor U22322 (N_22322,N_21644,N_21635);
and U22323 (N_22323,N_21765,N_21390);
nor U22324 (N_22324,N_21520,N_21330);
and U22325 (N_22325,N_21268,N_21770);
nand U22326 (N_22326,N_21491,N_21502);
or U22327 (N_22327,N_21738,N_21716);
nor U22328 (N_22328,N_21645,N_21713);
and U22329 (N_22329,N_21648,N_21870);
nor U22330 (N_22330,N_21721,N_21729);
nor U22331 (N_22331,N_21482,N_21443);
or U22332 (N_22332,N_21375,N_21518);
or U22333 (N_22333,N_21455,N_21313);
nor U22334 (N_22334,N_21359,N_21728);
nor U22335 (N_22335,N_21347,N_21579);
xnor U22336 (N_22336,N_21811,N_21653);
or U22337 (N_22337,N_21556,N_21766);
nor U22338 (N_22338,N_21467,N_21405);
and U22339 (N_22339,N_21274,N_21645);
or U22340 (N_22340,N_21337,N_21860);
nand U22341 (N_22341,N_21279,N_21488);
nand U22342 (N_22342,N_21435,N_21443);
or U22343 (N_22343,N_21478,N_21711);
xnor U22344 (N_22344,N_21458,N_21863);
nand U22345 (N_22345,N_21869,N_21537);
nor U22346 (N_22346,N_21353,N_21640);
and U22347 (N_22347,N_21261,N_21706);
nand U22348 (N_22348,N_21672,N_21260);
nor U22349 (N_22349,N_21650,N_21657);
xnor U22350 (N_22350,N_21525,N_21675);
xor U22351 (N_22351,N_21821,N_21783);
nor U22352 (N_22352,N_21687,N_21415);
and U22353 (N_22353,N_21668,N_21611);
nand U22354 (N_22354,N_21358,N_21515);
nand U22355 (N_22355,N_21575,N_21676);
xor U22356 (N_22356,N_21664,N_21274);
or U22357 (N_22357,N_21411,N_21574);
and U22358 (N_22358,N_21433,N_21408);
nor U22359 (N_22359,N_21383,N_21294);
and U22360 (N_22360,N_21353,N_21662);
and U22361 (N_22361,N_21262,N_21614);
or U22362 (N_22362,N_21796,N_21389);
xnor U22363 (N_22363,N_21730,N_21488);
and U22364 (N_22364,N_21677,N_21831);
or U22365 (N_22365,N_21352,N_21590);
nand U22366 (N_22366,N_21592,N_21575);
and U22367 (N_22367,N_21564,N_21259);
or U22368 (N_22368,N_21383,N_21508);
xor U22369 (N_22369,N_21578,N_21636);
and U22370 (N_22370,N_21293,N_21438);
or U22371 (N_22371,N_21813,N_21432);
and U22372 (N_22372,N_21767,N_21496);
nor U22373 (N_22373,N_21481,N_21610);
xor U22374 (N_22374,N_21843,N_21800);
or U22375 (N_22375,N_21554,N_21852);
and U22376 (N_22376,N_21527,N_21257);
or U22377 (N_22377,N_21736,N_21729);
and U22378 (N_22378,N_21844,N_21771);
or U22379 (N_22379,N_21669,N_21679);
or U22380 (N_22380,N_21578,N_21523);
or U22381 (N_22381,N_21535,N_21703);
xor U22382 (N_22382,N_21795,N_21675);
nor U22383 (N_22383,N_21287,N_21605);
nand U22384 (N_22384,N_21425,N_21797);
nor U22385 (N_22385,N_21398,N_21823);
or U22386 (N_22386,N_21789,N_21819);
and U22387 (N_22387,N_21619,N_21530);
nand U22388 (N_22388,N_21303,N_21297);
or U22389 (N_22389,N_21370,N_21442);
and U22390 (N_22390,N_21719,N_21438);
or U22391 (N_22391,N_21574,N_21853);
nand U22392 (N_22392,N_21324,N_21540);
xnor U22393 (N_22393,N_21843,N_21831);
nand U22394 (N_22394,N_21459,N_21607);
nand U22395 (N_22395,N_21355,N_21292);
or U22396 (N_22396,N_21531,N_21810);
and U22397 (N_22397,N_21365,N_21302);
or U22398 (N_22398,N_21404,N_21253);
or U22399 (N_22399,N_21301,N_21693);
nand U22400 (N_22400,N_21528,N_21719);
nand U22401 (N_22401,N_21490,N_21355);
xor U22402 (N_22402,N_21476,N_21430);
xor U22403 (N_22403,N_21754,N_21861);
nand U22404 (N_22404,N_21500,N_21606);
nand U22405 (N_22405,N_21390,N_21268);
or U22406 (N_22406,N_21563,N_21344);
nand U22407 (N_22407,N_21811,N_21796);
or U22408 (N_22408,N_21692,N_21647);
nor U22409 (N_22409,N_21470,N_21557);
nand U22410 (N_22410,N_21576,N_21356);
or U22411 (N_22411,N_21478,N_21656);
nand U22412 (N_22412,N_21690,N_21303);
and U22413 (N_22413,N_21826,N_21434);
nor U22414 (N_22414,N_21360,N_21785);
nor U22415 (N_22415,N_21590,N_21743);
xor U22416 (N_22416,N_21433,N_21352);
and U22417 (N_22417,N_21869,N_21290);
nand U22418 (N_22418,N_21676,N_21568);
nand U22419 (N_22419,N_21297,N_21545);
nor U22420 (N_22420,N_21427,N_21322);
nand U22421 (N_22421,N_21352,N_21348);
xor U22422 (N_22422,N_21819,N_21449);
nor U22423 (N_22423,N_21472,N_21451);
and U22424 (N_22424,N_21616,N_21753);
xor U22425 (N_22425,N_21586,N_21615);
and U22426 (N_22426,N_21460,N_21717);
nand U22427 (N_22427,N_21710,N_21623);
nand U22428 (N_22428,N_21262,N_21803);
nand U22429 (N_22429,N_21349,N_21289);
or U22430 (N_22430,N_21710,N_21616);
or U22431 (N_22431,N_21705,N_21671);
and U22432 (N_22432,N_21375,N_21259);
or U22433 (N_22433,N_21793,N_21746);
nand U22434 (N_22434,N_21670,N_21291);
and U22435 (N_22435,N_21643,N_21779);
xnor U22436 (N_22436,N_21456,N_21697);
and U22437 (N_22437,N_21487,N_21659);
and U22438 (N_22438,N_21721,N_21661);
or U22439 (N_22439,N_21781,N_21597);
or U22440 (N_22440,N_21861,N_21700);
xor U22441 (N_22441,N_21417,N_21392);
nor U22442 (N_22442,N_21682,N_21294);
xor U22443 (N_22443,N_21572,N_21492);
and U22444 (N_22444,N_21560,N_21755);
and U22445 (N_22445,N_21437,N_21498);
or U22446 (N_22446,N_21436,N_21793);
nand U22447 (N_22447,N_21689,N_21521);
and U22448 (N_22448,N_21300,N_21459);
and U22449 (N_22449,N_21641,N_21476);
nor U22450 (N_22450,N_21735,N_21254);
or U22451 (N_22451,N_21632,N_21446);
and U22452 (N_22452,N_21296,N_21607);
xor U22453 (N_22453,N_21524,N_21273);
or U22454 (N_22454,N_21674,N_21742);
nand U22455 (N_22455,N_21348,N_21816);
nand U22456 (N_22456,N_21740,N_21689);
and U22457 (N_22457,N_21619,N_21298);
nand U22458 (N_22458,N_21852,N_21790);
and U22459 (N_22459,N_21709,N_21516);
and U22460 (N_22460,N_21437,N_21276);
nand U22461 (N_22461,N_21254,N_21874);
nor U22462 (N_22462,N_21253,N_21415);
xnor U22463 (N_22463,N_21668,N_21630);
nor U22464 (N_22464,N_21824,N_21858);
nand U22465 (N_22465,N_21804,N_21350);
xnor U22466 (N_22466,N_21820,N_21313);
and U22467 (N_22467,N_21617,N_21523);
or U22468 (N_22468,N_21335,N_21722);
xnor U22469 (N_22469,N_21360,N_21637);
nor U22470 (N_22470,N_21557,N_21830);
xnor U22471 (N_22471,N_21265,N_21702);
and U22472 (N_22472,N_21606,N_21531);
xor U22473 (N_22473,N_21441,N_21829);
nand U22474 (N_22474,N_21270,N_21380);
or U22475 (N_22475,N_21693,N_21494);
or U22476 (N_22476,N_21564,N_21766);
nor U22477 (N_22477,N_21312,N_21662);
and U22478 (N_22478,N_21580,N_21745);
nor U22479 (N_22479,N_21618,N_21541);
nor U22480 (N_22480,N_21659,N_21641);
nand U22481 (N_22481,N_21407,N_21681);
and U22482 (N_22482,N_21822,N_21483);
and U22483 (N_22483,N_21516,N_21817);
nor U22484 (N_22484,N_21747,N_21512);
nor U22485 (N_22485,N_21814,N_21724);
nor U22486 (N_22486,N_21411,N_21845);
and U22487 (N_22487,N_21383,N_21663);
nand U22488 (N_22488,N_21541,N_21842);
or U22489 (N_22489,N_21555,N_21446);
xnor U22490 (N_22490,N_21756,N_21535);
xor U22491 (N_22491,N_21531,N_21266);
nand U22492 (N_22492,N_21520,N_21373);
nor U22493 (N_22493,N_21520,N_21689);
and U22494 (N_22494,N_21554,N_21720);
nor U22495 (N_22495,N_21714,N_21541);
nor U22496 (N_22496,N_21578,N_21588);
nand U22497 (N_22497,N_21690,N_21779);
or U22498 (N_22498,N_21256,N_21464);
xor U22499 (N_22499,N_21505,N_21468);
nor U22500 (N_22500,N_22482,N_22027);
nor U22501 (N_22501,N_22394,N_22297);
nor U22502 (N_22502,N_22356,N_22035);
and U22503 (N_22503,N_22073,N_21916);
and U22504 (N_22504,N_22148,N_22327);
or U22505 (N_22505,N_22338,N_22071);
nand U22506 (N_22506,N_21929,N_22026);
nor U22507 (N_22507,N_22168,N_22305);
xnor U22508 (N_22508,N_22334,N_22090);
nand U22509 (N_22509,N_22199,N_22295);
or U22510 (N_22510,N_22084,N_22300);
and U22511 (N_22511,N_21901,N_22006);
or U22512 (N_22512,N_22422,N_22389);
and U22513 (N_22513,N_21955,N_22047);
nand U22514 (N_22514,N_22485,N_22321);
xnor U22515 (N_22515,N_22149,N_22140);
or U22516 (N_22516,N_22183,N_22014);
nor U22517 (N_22517,N_22000,N_22491);
xor U22518 (N_22518,N_22442,N_22102);
nor U22519 (N_22519,N_21974,N_22311);
xnor U22520 (N_22520,N_21898,N_22196);
nor U22521 (N_22521,N_22056,N_22087);
xnor U22522 (N_22522,N_22478,N_21952);
nand U22523 (N_22523,N_21875,N_21956);
nor U22524 (N_22524,N_22432,N_22162);
nand U22525 (N_22525,N_22113,N_22314);
nand U22526 (N_22526,N_21909,N_21993);
nor U22527 (N_22527,N_21996,N_22043);
nand U22528 (N_22528,N_22246,N_22384);
nand U22529 (N_22529,N_22150,N_22299);
xor U22530 (N_22530,N_22424,N_22318);
or U22531 (N_22531,N_22271,N_22267);
or U22532 (N_22532,N_21938,N_22120);
or U22533 (N_22533,N_21928,N_22023);
nand U22534 (N_22534,N_22391,N_22274);
or U22535 (N_22535,N_21919,N_22032);
xor U22536 (N_22536,N_22307,N_22059);
or U22537 (N_22537,N_22171,N_22348);
or U22538 (N_22538,N_22228,N_22283);
or U22539 (N_22539,N_22407,N_22291);
nor U22540 (N_22540,N_22446,N_22017);
nor U22541 (N_22541,N_22202,N_22405);
and U22542 (N_22542,N_22116,N_22031);
and U22543 (N_22543,N_22088,N_21908);
nand U22544 (N_22544,N_22178,N_22414);
nand U22545 (N_22545,N_22040,N_22055);
and U22546 (N_22546,N_22365,N_22357);
and U22547 (N_22547,N_22490,N_22133);
xor U22548 (N_22548,N_22494,N_22119);
nor U22549 (N_22549,N_22203,N_22306);
xnor U22550 (N_22550,N_22046,N_22107);
and U22551 (N_22551,N_22492,N_22235);
or U22552 (N_22552,N_22099,N_22118);
nor U22553 (N_22553,N_22256,N_22335);
or U22554 (N_22554,N_22159,N_22262);
or U22555 (N_22555,N_22117,N_22220);
or U22556 (N_22556,N_22433,N_22114);
nand U22557 (N_22557,N_22170,N_22497);
nor U22558 (N_22558,N_22244,N_22319);
xnor U22559 (N_22559,N_21918,N_21933);
nor U22560 (N_22560,N_22060,N_22331);
and U22561 (N_22561,N_22209,N_21985);
or U22562 (N_22562,N_22280,N_22393);
and U22563 (N_22563,N_22142,N_21926);
or U22564 (N_22564,N_22222,N_22434);
or U22565 (N_22565,N_22363,N_22320);
or U22566 (N_22566,N_22112,N_22163);
nand U22567 (N_22567,N_22350,N_22138);
or U22568 (N_22568,N_21992,N_21950);
nand U22569 (N_22569,N_22083,N_22210);
nor U22570 (N_22570,N_22459,N_22428);
nor U22571 (N_22571,N_22065,N_22408);
and U22572 (N_22572,N_22077,N_22259);
nor U22573 (N_22573,N_21946,N_21945);
and U22574 (N_22574,N_22011,N_21991);
nor U22575 (N_22575,N_22039,N_22156);
and U22576 (N_22576,N_22215,N_22447);
nand U22577 (N_22577,N_22330,N_22078);
nor U22578 (N_22578,N_22021,N_22252);
nor U22579 (N_22579,N_22160,N_22097);
and U22580 (N_22580,N_22127,N_22284);
nand U22581 (N_22581,N_22075,N_22377);
and U22582 (N_22582,N_22450,N_21960);
or U22583 (N_22583,N_22421,N_22460);
nor U22584 (N_22584,N_22385,N_21983);
or U22585 (N_22585,N_22469,N_22126);
or U22586 (N_22586,N_21981,N_22315);
nor U22587 (N_22587,N_22234,N_22361);
xor U22588 (N_22588,N_22376,N_21972);
or U22589 (N_22589,N_21911,N_22044);
and U22590 (N_22590,N_22332,N_22192);
and U22591 (N_22591,N_21995,N_22019);
xnor U22592 (N_22592,N_22495,N_22205);
nand U22593 (N_22593,N_22470,N_22211);
or U22594 (N_22594,N_22227,N_22223);
nor U22595 (N_22595,N_22301,N_22191);
and U22596 (N_22596,N_22456,N_22404);
or U22597 (N_22597,N_22237,N_21903);
nor U22598 (N_22598,N_22395,N_22008);
nor U22599 (N_22599,N_21998,N_22416);
or U22600 (N_22600,N_22474,N_22415);
nand U22601 (N_22601,N_22129,N_22337);
xnor U22602 (N_22602,N_21971,N_21947);
or U22603 (N_22603,N_21883,N_22176);
and U22604 (N_22604,N_22290,N_22037);
nor U22605 (N_22605,N_22190,N_22009);
nor U22606 (N_22606,N_22342,N_21891);
or U22607 (N_22607,N_21962,N_21917);
nor U22608 (N_22608,N_21895,N_22188);
xor U22609 (N_22609,N_22136,N_22058);
and U22610 (N_22610,N_22134,N_22184);
or U22611 (N_22611,N_22169,N_21969);
and U22612 (N_22612,N_22147,N_22464);
and U22613 (N_22613,N_22488,N_22275);
nor U22614 (N_22614,N_22076,N_22177);
xnor U22615 (N_22615,N_22304,N_22152);
nor U22616 (N_22616,N_22195,N_22351);
nand U22617 (N_22617,N_22364,N_22238);
xor U22618 (N_22618,N_22022,N_22413);
xor U22619 (N_22619,N_22208,N_21968);
nand U22620 (N_22620,N_22198,N_22093);
nand U22621 (N_22621,N_22095,N_21984);
or U22622 (N_22622,N_22336,N_22236);
nor U22623 (N_22623,N_22325,N_22279);
and U22624 (N_22624,N_22108,N_22067);
and U22625 (N_22625,N_22427,N_21966);
nand U22626 (N_22626,N_22001,N_22483);
nor U22627 (N_22627,N_22172,N_22398);
nand U22628 (N_22628,N_22457,N_22346);
nor U22629 (N_22629,N_22294,N_22182);
nand U22630 (N_22630,N_22388,N_22368);
xnor U22631 (N_22631,N_22232,N_22317);
xor U22632 (N_22632,N_22371,N_22029);
nand U22633 (N_22633,N_22204,N_22358);
xnor U22634 (N_22634,N_22092,N_22224);
and U22635 (N_22635,N_22481,N_22323);
nand U22636 (N_22636,N_21897,N_22231);
xnor U22637 (N_22637,N_22461,N_22080);
and U22638 (N_22638,N_22050,N_22179);
and U22639 (N_22639,N_22465,N_21900);
or U22640 (N_22640,N_22310,N_21951);
or U22641 (N_22641,N_22165,N_22139);
and U22642 (N_22642,N_22241,N_22091);
xnor U22643 (N_22643,N_22402,N_22226);
xnor U22644 (N_22644,N_22146,N_22423);
xnor U22645 (N_22645,N_22396,N_22069);
nor U22646 (N_22646,N_22042,N_22033);
nand U22647 (N_22647,N_22486,N_22344);
xnor U22648 (N_22648,N_21920,N_22125);
nand U22649 (N_22649,N_22089,N_22004);
xnor U22650 (N_22650,N_22201,N_22189);
and U22651 (N_22651,N_22467,N_22400);
xor U22652 (N_22652,N_22372,N_21925);
xor U22653 (N_22653,N_22286,N_22441);
or U22654 (N_22654,N_22499,N_22034);
xnor U22655 (N_22655,N_22063,N_22454);
nor U22656 (N_22656,N_22479,N_22229);
or U22657 (N_22657,N_21913,N_22403);
and U22658 (N_22658,N_22141,N_22166);
and U22659 (N_22659,N_21880,N_22362);
nand U22660 (N_22660,N_21878,N_22249);
or U22661 (N_22661,N_21905,N_22436);
nor U22662 (N_22662,N_22130,N_22386);
xor U22663 (N_22663,N_22322,N_22086);
and U22664 (N_22664,N_22397,N_22105);
nor U22665 (N_22665,N_22016,N_22287);
xnor U22666 (N_22666,N_22013,N_21943);
nand U22667 (N_22667,N_22349,N_21927);
xnor U22668 (N_22668,N_22473,N_22135);
and U22669 (N_22669,N_22145,N_21914);
nor U22670 (N_22670,N_21934,N_22155);
and U22671 (N_22671,N_22266,N_22217);
nor U22672 (N_22672,N_21931,N_22419);
and U22673 (N_22673,N_22045,N_21949);
nand U22674 (N_22674,N_22174,N_22018);
and U22675 (N_22675,N_22082,N_22072);
and U22676 (N_22676,N_21941,N_22298);
nand U22677 (N_22677,N_22057,N_22281);
xnor U22678 (N_22678,N_22472,N_22066);
nand U22679 (N_22679,N_22339,N_22242);
nor U22680 (N_22680,N_22366,N_21893);
and U22681 (N_22681,N_21935,N_22187);
nor U22682 (N_22682,N_22124,N_22079);
xor U22683 (N_22683,N_21963,N_22316);
or U22684 (N_22684,N_22333,N_22024);
and U22685 (N_22685,N_21953,N_22420);
or U22686 (N_22686,N_22173,N_22341);
and U22687 (N_22687,N_22100,N_21930);
or U22688 (N_22688,N_21989,N_21973);
nor U22689 (N_22689,N_22484,N_22186);
and U22690 (N_22690,N_22128,N_22425);
or U22691 (N_22691,N_21889,N_22326);
and U22692 (N_22692,N_21904,N_22276);
nand U22693 (N_22693,N_22193,N_22430);
and U22694 (N_22694,N_22435,N_22122);
nand U22695 (N_22695,N_22378,N_22282);
or U22696 (N_22696,N_21890,N_21978);
or U22697 (N_22697,N_22104,N_21997);
nor U22698 (N_22698,N_22381,N_21954);
and U22699 (N_22699,N_21948,N_22392);
nand U22700 (N_22700,N_22268,N_21937);
or U22701 (N_22701,N_21921,N_22496);
or U22702 (N_22702,N_22121,N_22289);
and U22703 (N_22703,N_22213,N_21885);
xor U22704 (N_22704,N_22005,N_21967);
xnor U22705 (N_22705,N_21976,N_22049);
nand U22706 (N_22706,N_21886,N_22015);
or U22707 (N_22707,N_22458,N_22328);
and U22708 (N_22708,N_22028,N_22302);
or U22709 (N_22709,N_22219,N_21977);
xor U22710 (N_22710,N_22367,N_21994);
xnor U22711 (N_22711,N_22345,N_22218);
or U22712 (N_22712,N_22062,N_22106);
and U22713 (N_22713,N_21987,N_22094);
nor U22714 (N_22714,N_22151,N_22401);
nor U22715 (N_22715,N_21906,N_22216);
nand U22716 (N_22716,N_22101,N_21988);
nor U22717 (N_22717,N_22418,N_22370);
or U22718 (N_22718,N_21961,N_21986);
or U22719 (N_22719,N_22185,N_22257);
xor U22720 (N_22720,N_22054,N_22448);
nor U22721 (N_22721,N_22374,N_22489);
nor U22722 (N_22722,N_22383,N_22477);
or U22723 (N_22723,N_22053,N_22175);
nor U22724 (N_22724,N_22352,N_21894);
nand U22725 (N_22725,N_22233,N_22260);
or U22726 (N_22726,N_22269,N_21942);
nor U22727 (N_22727,N_22272,N_22463);
nand U22728 (N_22728,N_22429,N_22221);
and U22729 (N_22729,N_22411,N_22230);
nor U22730 (N_22730,N_21999,N_22359);
and U22731 (N_22731,N_22003,N_22096);
nor U22732 (N_22732,N_22030,N_21959);
or U22733 (N_22733,N_22288,N_22343);
and U22734 (N_22734,N_22110,N_22197);
and U22735 (N_22735,N_21965,N_22417);
or U22736 (N_22736,N_22245,N_22412);
nand U22737 (N_22737,N_22445,N_21907);
nand U22738 (N_22738,N_22041,N_22303);
nand U22739 (N_22739,N_22250,N_22292);
and U22740 (N_22740,N_22194,N_22387);
and U22741 (N_22741,N_22061,N_22111);
or U22742 (N_22742,N_22243,N_22466);
nand U22743 (N_22743,N_22153,N_22158);
nor U22744 (N_22744,N_22437,N_22103);
or U22745 (N_22745,N_22253,N_22426);
xor U22746 (N_22746,N_22453,N_21879);
nand U22747 (N_22747,N_22439,N_22085);
or U22748 (N_22748,N_21958,N_22382);
nor U22749 (N_22749,N_22240,N_21970);
xor U22750 (N_22750,N_22180,N_22048);
xnor U22751 (N_22751,N_21939,N_22264);
xor U22752 (N_22752,N_22144,N_21902);
xnor U22753 (N_22753,N_22360,N_22308);
xor U22754 (N_22754,N_21915,N_22143);
nand U22755 (N_22755,N_22263,N_22431);
nand U22756 (N_22756,N_22010,N_21912);
nand U22757 (N_22757,N_22476,N_21892);
nand U22758 (N_22758,N_22002,N_21910);
xnor U22759 (N_22759,N_22167,N_22410);
nand U22760 (N_22760,N_22329,N_21990);
xnor U22761 (N_22761,N_22390,N_21944);
and U22762 (N_22762,N_22064,N_22277);
nor U22763 (N_22763,N_21896,N_22131);
xor U22764 (N_22764,N_22293,N_22020);
or U22765 (N_22765,N_22285,N_22247);
or U22766 (N_22766,N_22468,N_21979);
xnor U22767 (N_22767,N_22443,N_22137);
nand U22768 (N_22768,N_22254,N_22296);
nand U22769 (N_22769,N_22455,N_22132);
nand U22770 (N_22770,N_21957,N_22115);
xor U22771 (N_22771,N_21899,N_22379);
xor U22772 (N_22772,N_22212,N_22052);
xor U22773 (N_22773,N_22265,N_22475);
nor U22774 (N_22774,N_22493,N_22340);
xnor U22775 (N_22775,N_21876,N_22206);
and U22776 (N_22776,N_21924,N_21884);
xnor U22777 (N_22777,N_21980,N_22181);
xnor U22778 (N_22778,N_21964,N_22098);
and U22779 (N_22779,N_22462,N_22025);
nor U22780 (N_22780,N_22154,N_22038);
nor U22781 (N_22781,N_22369,N_22157);
nor U22782 (N_22782,N_22012,N_22354);
nor U22783 (N_22783,N_22081,N_22375);
nor U22784 (N_22784,N_22313,N_22444);
nand U22785 (N_22785,N_22498,N_22355);
xor U22786 (N_22786,N_22207,N_22070);
nand U22787 (N_22787,N_21932,N_22273);
and U22788 (N_22788,N_21982,N_22214);
or U22789 (N_22789,N_22406,N_21936);
or U22790 (N_22790,N_22373,N_22440);
nand U22791 (N_22791,N_22164,N_22074);
nand U22792 (N_22792,N_22161,N_22200);
and U22793 (N_22793,N_22051,N_22270);
or U22794 (N_22794,N_22123,N_21877);
and U22795 (N_22795,N_22258,N_22309);
xor U22796 (N_22796,N_22487,N_21923);
xor U22797 (N_22797,N_22347,N_21881);
or U22798 (N_22798,N_21940,N_22068);
nor U22799 (N_22799,N_22225,N_22248);
xor U22800 (N_22800,N_22452,N_21922);
nand U22801 (N_22801,N_22324,N_22255);
or U22802 (N_22802,N_22036,N_22449);
nor U22803 (N_22803,N_21888,N_22278);
and U22804 (N_22804,N_22251,N_22261);
xor U22805 (N_22805,N_22480,N_22312);
nor U22806 (N_22806,N_22451,N_22109);
xnor U22807 (N_22807,N_22239,N_21882);
xnor U22808 (N_22808,N_22471,N_22438);
or U22809 (N_22809,N_22399,N_21975);
nor U22810 (N_22810,N_22353,N_22380);
xnor U22811 (N_22811,N_21887,N_22409);
nand U22812 (N_22812,N_22007,N_22491);
xor U22813 (N_22813,N_22431,N_21957);
xor U22814 (N_22814,N_22109,N_21964);
or U22815 (N_22815,N_21917,N_22319);
and U22816 (N_22816,N_22176,N_22283);
nor U22817 (N_22817,N_21886,N_22316);
nor U22818 (N_22818,N_22399,N_22083);
xor U22819 (N_22819,N_22293,N_22310);
xnor U22820 (N_22820,N_22361,N_22393);
nor U22821 (N_22821,N_21961,N_22303);
and U22822 (N_22822,N_22382,N_21877);
and U22823 (N_22823,N_22408,N_21934);
and U22824 (N_22824,N_22275,N_21935);
nor U22825 (N_22825,N_22432,N_22352);
nand U22826 (N_22826,N_22105,N_22311);
nand U22827 (N_22827,N_22073,N_22294);
nand U22828 (N_22828,N_22030,N_21999);
or U22829 (N_22829,N_22281,N_21958);
xnor U22830 (N_22830,N_22497,N_22251);
or U22831 (N_22831,N_22189,N_21989);
nand U22832 (N_22832,N_21981,N_22213);
xor U22833 (N_22833,N_22215,N_22229);
or U22834 (N_22834,N_21993,N_22208);
nand U22835 (N_22835,N_22473,N_21960);
and U22836 (N_22836,N_22227,N_22068);
or U22837 (N_22837,N_22140,N_21914);
nand U22838 (N_22838,N_22431,N_22478);
xor U22839 (N_22839,N_22000,N_22071);
xnor U22840 (N_22840,N_22165,N_22102);
nand U22841 (N_22841,N_22168,N_21961);
nand U22842 (N_22842,N_22181,N_22302);
xor U22843 (N_22843,N_22216,N_22488);
nand U22844 (N_22844,N_22210,N_22147);
xor U22845 (N_22845,N_22473,N_21958);
nand U22846 (N_22846,N_22377,N_21946);
xor U22847 (N_22847,N_22101,N_22431);
or U22848 (N_22848,N_22006,N_22482);
nand U22849 (N_22849,N_22151,N_22071);
or U22850 (N_22850,N_22415,N_22093);
xnor U22851 (N_22851,N_22106,N_22460);
and U22852 (N_22852,N_22221,N_22208);
or U22853 (N_22853,N_22398,N_22068);
and U22854 (N_22854,N_22028,N_21944);
nor U22855 (N_22855,N_22282,N_22018);
or U22856 (N_22856,N_22141,N_22330);
nor U22857 (N_22857,N_22129,N_21907);
or U22858 (N_22858,N_22155,N_22291);
xnor U22859 (N_22859,N_22315,N_21939);
xor U22860 (N_22860,N_22212,N_22398);
xnor U22861 (N_22861,N_22199,N_22097);
nor U22862 (N_22862,N_21878,N_22163);
and U22863 (N_22863,N_22062,N_22319);
xor U22864 (N_22864,N_22455,N_22292);
xor U22865 (N_22865,N_22200,N_22113);
xor U22866 (N_22866,N_22404,N_22399);
or U22867 (N_22867,N_21960,N_22118);
xor U22868 (N_22868,N_22153,N_21896);
xor U22869 (N_22869,N_22279,N_22041);
or U22870 (N_22870,N_22092,N_22166);
xor U22871 (N_22871,N_21956,N_22354);
and U22872 (N_22872,N_22038,N_21903);
xnor U22873 (N_22873,N_22034,N_22446);
and U22874 (N_22874,N_21919,N_22159);
nand U22875 (N_22875,N_21985,N_21971);
nand U22876 (N_22876,N_21999,N_22225);
nand U22877 (N_22877,N_22351,N_22377);
nand U22878 (N_22878,N_22415,N_22164);
or U22879 (N_22879,N_22138,N_22467);
nand U22880 (N_22880,N_22341,N_22258);
nand U22881 (N_22881,N_22439,N_22463);
nand U22882 (N_22882,N_22182,N_22164);
and U22883 (N_22883,N_22440,N_22004);
and U22884 (N_22884,N_22196,N_22157);
and U22885 (N_22885,N_22303,N_22113);
nand U22886 (N_22886,N_22010,N_22263);
nand U22887 (N_22887,N_22498,N_22090);
nor U22888 (N_22888,N_22430,N_22099);
nor U22889 (N_22889,N_22495,N_22043);
or U22890 (N_22890,N_22242,N_22484);
nand U22891 (N_22891,N_22117,N_22468);
xor U22892 (N_22892,N_22318,N_22441);
nand U22893 (N_22893,N_22061,N_22225);
xnor U22894 (N_22894,N_22465,N_22010);
nand U22895 (N_22895,N_22081,N_22434);
or U22896 (N_22896,N_22197,N_22166);
xnor U22897 (N_22897,N_21892,N_21968);
or U22898 (N_22898,N_22050,N_22116);
nor U22899 (N_22899,N_22140,N_22029);
nand U22900 (N_22900,N_22180,N_22464);
nand U22901 (N_22901,N_22036,N_22106);
xor U22902 (N_22902,N_22186,N_21905);
xnor U22903 (N_22903,N_22091,N_21947);
xor U22904 (N_22904,N_22438,N_22277);
or U22905 (N_22905,N_22072,N_22099);
xnor U22906 (N_22906,N_22149,N_22194);
xnor U22907 (N_22907,N_22311,N_22123);
xnor U22908 (N_22908,N_22228,N_22363);
or U22909 (N_22909,N_22097,N_22472);
xnor U22910 (N_22910,N_21989,N_22147);
nor U22911 (N_22911,N_22397,N_22182);
and U22912 (N_22912,N_22147,N_22474);
or U22913 (N_22913,N_22157,N_22073);
nor U22914 (N_22914,N_22296,N_22291);
and U22915 (N_22915,N_22099,N_22266);
nor U22916 (N_22916,N_22456,N_21882);
xor U22917 (N_22917,N_22208,N_21895);
xor U22918 (N_22918,N_22138,N_22245);
nand U22919 (N_22919,N_22024,N_22281);
nor U22920 (N_22920,N_21984,N_22032);
nand U22921 (N_22921,N_22403,N_22257);
or U22922 (N_22922,N_22124,N_21983);
nand U22923 (N_22923,N_22233,N_22006);
or U22924 (N_22924,N_21966,N_22356);
xor U22925 (N_22925,N_21937,N_22346);
and U22926 (N_22926,N_22132,N_22084);
nand U22927 (N_22927,N_22221,N_22161);
nand U22928 (N_22928,N_22372,N_22441);
nand U22929 (N_22929,N_22205,N_22484);
nand U22930 (N_22930,N_22419,N_22000);
and U22931 (N_22931,N_22224,N_21897);
and U22932 (N_22932,N_22427,N_22087);
xor U22933 (N_22933,N_21900,N_22378);
nor U22934 (N_22934,N_21902,N_22183);
xnor U22935 (N_22935,N_22304,N_22465);
xnor U22936 (N_22936,N_22276,N_22103);
or U22937 (N_22937,N_22139,N_22237);
and U22938 (N_22938,N_21984,N_22288);
xor U22939 (N_22939,N_21943,N_21928);
xnor U22940 (N_22940,N_22393,N_22405);
nor U22941 (N_22941,N_22269,N_22086);
xnor U22942 (N_22942,N_22305,N_22354);
and U22943 (N_22943,N_22075,N_21944);
xnor U22944 (N_22944,N_21989,N_22145);
and U22945 (N_22945,N_22259,N_22215);
xnor U22946 (N_22946,N_21969,N_22279);
xor U22947 (N_22947,N_22219,N_22050);
xnor U22948 (N_22948,N_22228,N_21960);
nor U22949 (N_22949,N_22049,N_21882);
xnor U22950 (N_22950,N_22224,N_22176);
xor U22951 (N_22951,N_22494,N_22283);
nor U22952 (N_22952,N_22394,N_22334);
and U22953 (N_22953,N_22341,N_22265);
nand U22954 (N_22954,N_21958,N_22233);
or U22955 (N_22955,N_22322,N_22071);
nand U22956 (N_22956,N_22135,N_22188);
nand U22957 (N_22957,N_22449,N_21982);
xnor U22958 (N_22958,N_21993,N_22427);
xor U22959 (N_22959,N_21975,N_22338);
nor U22960 (N_22960,N_22257,N_22062);
nor U22961 (N_22961,N_22336,N_22369);
nand U22962 (N_22962,N_21975,N_22366);
and U22963 (N_22963,N_22276,N_21916);
xnor U22964 (N_22964,N_22227,N_22490);
nor U22965 (N_22965,N_22392,N_22371);
nand U22966 (N_22966,N_22349,N_22335);
xor U22967 (N_22967,N_21891,N_21936);
or U22968 (N_22968,N_22122,N_22247);
nor U22969 (N_22969,N_21961,N_21934);
nor U22970 (N_22970,N_22435,N_22091);
and U22971 (N_22971,N_22013,N_22297);
nor U22972 (N_22972,N_21935,N_22264);
or U22973 (N_22973,N_22049,N_22370);
and U22974 (N_22974,N_22118,N_22269);
nor U22975 (N_22975,N_21933,N_22164);
xor U22976 (N_22976,N_22370,N_22153);
and U22977 (N_22977,N_22381,N_22168);
nand U22978 (N_22978,N_22470,N_22274);
nor U22979 (N_22979,N_21890,N_21941);
nand U22980 (N_22980,N_22372,N_22327);
or U22981 (N_22981,N_21936,N_21905);
nor U22982 (N_22982,N_22279,N_22438);
and U22983 (N_22983,N_21911,N_22186);
nand U22984 (N_22984,N_21946,N_22402);
and U22985 (N_22985,N_22271,N_22210);
nor U22986 (N_22986,N_22250,N_21937);
nor U22987 (N_22987,N_22357,N_22250);
or U22988 (N_22988,N_22290,N_22267);
nor U22989 (N_22989,N_22266,N_22290);
nand U22990 (N_22990,N_21958,N_22332);
or U22991 (N_22991,N_22270,N_22410);
nand U22992 (N_22992,N_22024,N_22116);
nand U22993 (N_22993,N_22090,N_22162);
or U22994 (N_22994,N_22135,N_22101);
xnor U22995 (N_22995,N_22288,N_22344);
xnor U22996 (N_22996,N_21932,N_22021);
xor U22997 (N_22997,N_22070,N_22433);
or U22998 (N_22998,N_21927,N_22440);
nand U22999 (N_22999,N_22374,N_22143);
and U23000 (N_23000,N_22013,N_22299);
nand U23001 (N_23001,N_22175,N_22124);
and U23002 (N_23002,N_22168,N_22426);
or U23003 (N_23003,N_22213,N_21976);
xor U23004 (N_23004,N_22461,N_22320);
or U23005 (N_23005,N_22366,N_22191);
xor U23006 (N_23006,N_22478,N_21987);
nand U23007 (N_23007,N_21928,N_21897);
xnor U23008 (N_23008,N_22289,N_22185);
and U23009 (N_23009,N_21905,N_21897);
nand U23010 (N_23010,N_22091,N_22425);
xor U23011 (N_23011,N_22453,N_22326);
nor U23012 (N_23012,N_21894,N_22447);
nand U23013 (N_23013,N_22287,N_22001);
nor U23014 (N_23014,N_22114,N_22039);
and U23015 (N_23015,N_22449,N_22065);
nor U23016 (N_23016,N_22478,N_22278);
xor U23017 (N_23017,N_22180,N_22239);
and U23018 (N_23018,N_22167,N_22076);
or U23019 (N_23019,N_21977,N_22234);
nand U23020 (N_23020,N_22484,N_22326);
xnor U23021 (N_23021,N_21960,N_22065);
nor U23022 (N_23022,N_22489,N_22150);
nand U23023 (N_23023,N_22391,N_21878);
nand U23024 (N_23024,N_22401,N_22347);
or U23025 (N_23025,N_22088,N_21922);
nand U23026 (N_23026,N_22300,N_21903);
xor U23027 (N_23027,N_22274,N_22206);
nor U23028 (N_23028,N_22444,N_22198);
xnor U23029 (N_23029,N_22355,N_22217);
and U23030 (N_23030,N_22084,N_22466);
nand U23031 (N_23031,N_22016,N_21989);
xor U23032 (N_23032,N_22426,N_22370);
and U23033 (N_23033,N_22102,N_22096);
xor U23034 (N_23034,N_22242,N_22480);
xor U23035 (N_23035,N_22076,N_22161);
xnor U23036 (N_23036,N_22381,N_22270);
xnor U23037 (N_23037,N_22079,N_22347);
xor U23038 (N_23038,N_22224,N_22321);
nand U23039 (N_23039,N_22037,N_22122);
nand U23040 (N_23040,N_22226,N_22308);
nor U23041 (N_23041,N_22337,N_22063);
and U23042 (N_23042,N_21915,N_21939);
xor U23043 (N_23043,N_22446,N_22359);
and U23044 (N_23044,N_22349,N_21941);
or U23045 (N_23045,N_21895,N_22325);
xnor U23046 (N_23046,N_22216,N_22095);
xnor U23047 (N_23047,N_22021,N_22311);
nand U23048 (N_23048,N_22021,N_22281);
nor U23049 (N_23049,N_22152,N_22452);
nand U23050 (N_23050,N_22216,N_22121);
nand U23051 (N_23051,N_21881,N_22033);
xor U23052 (N_23052,N_21996,N_22071);
and U23053 (N_23053,N_21950,N_22167);
xor U23054 (N_23054,N_22181,N_22084);
nor U23055 (N_23055,N_22399,N_22337);
nor U23056 (N_23056,N_22090,N_21907);
or U23057 (N_23057,N_22363,N_22173);
xnor U23058 (N_23058,N_21901,N_21934);
nor U23059 (N_23059,N_21941,N_22158);
nor U23060 (N_23060,N_22142,N_22016);
xnor U23061 (N_23061,N_22230,N_22379);
xor U23062 (N_23062,N_22183,N_22255);
xnor U23063 (N_23063,N_22274,N_21887);
nand U23064 (N_23064,N_22356,N_22496);
xnor U23065 (N_23065,N_21936,N_22141);
nand U23066 (N_23066,N_22365,N_22014);
and U23067 (N_23067,N_22299,N_22263);
or U23068 (N_23068,N_22420,N_22276);
nand U23069 (N_23069,N_21994,N_22094);
nand U23070 (N_23070,N_22291,N_22366);
and U23071 (N_23071,N_22495,N_22225);
and U23072 (N_23072,N_22469,N_22170);
or U23073 (N_23073,N_22020,N_22085);
xor U23074 (N_23074,N_22127,N_22199);
and U23075 (N_23075,N_21894,N_22076);
nor U23076 (N_23076,N_22204,N_22266);
and U23077 (N_23077,N_22309,N_21956);
and U23078 (N_23078,N_22240,N_22266);
or U23079 (N_23079,N_22031,N_22396);
xor U23080 (N_23080,N_22045,N_22488);
xnor U23081 (N_23081,N_22339,N_21888);
nor U23082 (N_23082,N_22304,N_22342);
nor U23083 (N_23083,N_22261,N_22201);
or U23084 (N_23084,N_22374,N_22032);
nor U23085 (N_23085,N_22157,N_22375);
xnor U23086 (N_23086,N_22498,N_21916);
nand U23087 (N_23087,N_22205,N_22399);
nand U23088 (N_23088,N_21909,N_22326);
xnor U23089 (N_23089,N_21964,N_22021);
nand U23090 (N_23090,N_21892,N_22132);
or U23091 (N_23091,N_21991,N_22134);
and U23092 (N_23092,N_22401,N_22293);
or U23093 (N_23093,N_22426,N_22248);
and U23094 (N_23094,N_22248,N_22333);
xor U23095 (N_23095,N_22393,N_21979);
xnor U23096 (N_23096,N_22065,N_22004);
nor U23097 (N_23097,N_22305,N_22213);
nand U23098 (N_23098,N_21972,N_22215);
nor U23099 (N_23099,N_22221,N_22206);
xnor U23100 (N_23100,N_22336,N_22465);
or U23101 (N_23101,N_22214,N_21887);
and U23102 (N_23102,N_21930,N_22069);
xnor U23103 (N_23103,N_22495,N_22060);
nand U23104 (N_23104,N_22350,N_22441);
nand U23105 (N_23105,N_22352,N_22393);
nand U23106 (N_23106,N_22048,N_22430);
or U23107 (N_23107,N_22155,N_22499);
and U23108 (N_23108,N_22089,N_22015);
nor U23109 (N_23109,N_22100,N_21892);
nand U23110 (N_23110,N_21933,N_21953);
or U23111 (N_23111,N_22299,N_22199);
nand U23112 (N_23112,N_21997,N_22317);
nand U23113 (N_23113,N_21972,N_22371);
xnor U23114 (N_23114,N_22129,N_22258);
or U23115 (N_23115,N_22058,N_22125);
nand U23116 (N_23116,N_22061,N_22308);
or U23117 (N_23117,N_22472,N_21893);
or U23118 (N_23118,N_22132,N_22299);
xor U23119 (N_23119,N_21960,N_22244);
and U23120 (N_23120,N_22324,N_22437);
or U23121 (N_23121,N_22040,N_22160);
nand U23122 (N_23122,N_21943,N_22435);
nand U23123 (N_23123,N_22081,N_21968);
nor U23124 (N_23124,N_22127,N_22467);
or U23125 (N_23125,N_23031,N_22790);
xor U23126 (N_23126,N_22989,N_22895);
nand U23127 (N_23127,N_22578,N_22738);
nand U23128 (N_23128,N_22540,N_22651);
and U23129 (N_23129,N_22556,N_22656);
nor U23130 (N_23130,N_23028,N_22691);
or U23131 (N_23131,N_22543,N_23067);
or U23132 (N_23132,N_22580,N_22686);
nor U23133 (N_23133,N_22774,N_23024);
or U23134 (N_23134,N_22727,N_22632);
or U23135 (N_23135,N_22865,N_22677);
or U23136 (N_23136,N_22645,N_22652);
nand U23137 (N_23137,N_23098,N_23030);
nand U23138 (N_23138,N_22679,N_22600);
nand U23139 (N_23139,N_22689,N_23042);
and U23140 (N_23140,N_22539,N_22570);
xnor U23141 (N_23141,N_22897,N_23088);
nand U23142 (N_23142,N_22620,N_22856);
xnor U23143 (N_23143,N_22968,N_22757);
nor U23144 (N_23144,N_22951,N_22735);
nor U23145 (N_23145,N_23117,N_22532);
nand U23146 (N_23146,N_22877,N_22695);
and U23147 (N_23147,N_22665,N_22885);
nor U23148 (N_23148,N_22502,N_23040);
or U23149 (N_23149,N_23010,N_22805);
and U23150 (N_23150,N_23096,N_22998);
or U23151 (N_23151,N_23105,N_22924);
nand U23152 (N_23152,N_22752,N_22987);
or U23153 (N_23153,N_23035,N_22908);
nand U23154 (N_23154,N_23112,N_23116);
nand U23155 (N_23155,N_22820,N_23120);
xnor U23156 (N_23156,N_22607,N_22704);
nor U23157 (N_23157,N_22911,N_22575);
or U23158 (N_23158,N_23013,N_22546);
nand U23159 (N_23159,N_22929,N_22749);
xor U23160 (N_23160,N_22558,N_22581);
or U23161 (N_23161,N_22693,N_22669);
nor U23162 (N_23162,N_22974,N_22734);
nand U23163 (N_23163,N_23051,N_22697);
and U23164 (N_23164,N_22729,N_22746);
xnor U23165 (N_23165,N_23084,N_23121);
or U23166 (N_23166,N_22522,N_22896);
nand U23167 (N_23167,N_22643,N_22508);
or U23168 (N_23168,N_22939,N_22780);
or U23169 (N_23169,N_22721,N_23036);
xor U23170 (N_23170,N_22703,N_22694);
or U23171 (N_23171,N_23069,N_23110);
xnor U23172 (N_23172,N_22609,N_22542);
or U23173 (N_23173,N_23063,N_22850);
xnor U23174 (N_23174,N_23052,N_22615);
xnor U23175 (N_23175,N_22849,N_22829);
nor U23176 (N_23176,N_22655,N_22916);
nor U23177 (N_23177,N_22573,N_22934);
nor U23178 (N_23178,N_23057,N_22904);
xor U23179 (N_23179,N_22874,N_22720);
nor U23180 (N_23180,N_22664,N_22952);
nor U23181 (N_23181,N_23075,N_22634);
xnor U23182 (N_23182,N_23044,N_22517);
nor U23183 (N_23183,N_22725,N_23007);
and U23184 (N_23184,N_22733,N_22574);
and U23185 (N_23185,N_22893,N_22776);
and U23186 (N_23186,N_23006,N_22981);
xnor U23187 (N_23187,N_22960,N_23073);
or U23188 (N_23188,N_23047,N_22722);
xor U23189 (N_23189,N_22838,N_22595);
or U23190 (N_23190,N_22777,N_22894);
nor U23191 (N_23191,N_22657,N_22597);
xor U23192 (N_23192,N_22771,N_22547);
and U23193 (N_23193,N_23003,N_22631);
or U23194 (N_23194,N_22617,N_22699);
xor U23195 (N_23195,N_22994,N_23078);
nand U23196 (N_23196,N_23104,N_22843);
or U23197 (N_23197,N_23050,N_22822);
nor U23198 (N_23198,N_22674,N_22766);
nand U23199 (N_23199,N_22726,N_22943);
nand U23200 (N_23200,N_23111,N_22909);
or U23201 (N_23201,N_22804,N_22966);
nand U23202 (N_23202,N_22710,N_22637);
xnor U23203 (N_23203,N_22940,N_22767);
or U23204 (N_23204,N_22922,N_23018);
xnor U23205 (N_23205,N_22844,N_22673);
and U23206 (N_23206,N_22684,N_22898);
or U23207 (N_23207,N_22588,N_22654);
nor U23208 (N_23208,N_22983,N_22836);
nand U23209 (N_23209,N_22602,N_23022);
or U23210 (N_23210,N_23068,N_22971);
or U23211 (N_23211,N_22832,N_22923);
and U23212 (N_23212,N_22944,N_22649);
and U23213 (N_23213,N_22785,N_22511);
or U23214 (N_23214,N_23101,N_22680);
nand U23215 (N_23215,N_22685,N_22533);
and U23216 (N_23216,N_22984,N_23083);
nor U23217 (N_23217,N_23027,N_23056);
and U23218 (N_23218,N_22878,N_22913);
nor U23219 (N_23219,N_22853,N_22708);
or U23220 (N_23220,N_22819,N_22789);
nand U23221 (N_23221,N_22584,N_22612);
or U23222 (N_23222,N_22642,N_22910);
and U23223 (N_23223,N_22667,N_22826);
nand U23224 (N_23224,N_22606,N_22891);
or U23225 (N_23225,N_22628,N_23034);
or U23226 (N_23226,N_22577,N_22509);
and U23227 (N_23227,N_22641,N_23107);
or U23228 (N_23228,N_22763,N_22518);
xnor U23229 (N_23229,N_22847,N_22881);
nand U23230 (N_23230,N_22650,N_22696);
nor U23231 (N_23231,N_22963,N_22964);
or U23232 (N_23232,N_22801,N_22662);
and U23233 (N_23233,N_22997,N_23005);
nand U23234 (N_23234,N_22995,N_22839);
nand U23235 (N_23235,N_22961,N_22589);
or U23236 (N_23236,N_22553,N_22527);
or U23237 (N_23237,N_22567,N_22562);
nor U23238 (N_23238,N_22736,N_22985);
xor U23239 (N_23239,N_22690,N_23061);
or U23240 (N_23240,N_22803,N_22846);
or U23241 (N_23241,N_23020,N_22630);
or U23242 (N_23242,N_22792,N_23065);
or U23243 (N_23243,N_23114,N_22914);
nand U23244 (N_23244,N_22737,N_22698);
nand U23245 (N_23245,N_22870,N_22753);
nor U23246 (N_23246,N_23118,N_22858);
xnor U23247 (N_23247,N_22902,N_22793);
and U23248 (N_23248,N_22831,N_23011);
or U23249 (N_23249,N_22765,N_23087);
and U23250 (N_23250,N_22503,N_22937);
xnor U23251 (N_23251,N_22958,N_22975);
and U23252 (N_23252,N_23025,N_23095);
xor U23253 (N_23253,N_22730,N_22957);
xor U23254 (N_23254,N_22992,N_22841);
and U23255 (N_23255,N_23072,N_23026);
xor U23256 (N_23256,N_22755,N_22592);
nor U23257 (N_23257,N_22756,N_22571);
and U23258 (N_23258,N_22932,N_22927);
nand U23259 (N_23259,N_22507,N_22837);
nand U23260 (N_23260,N_22824,N_22644);
nor U23261 (N_23261,N_22977,N_22811);
xor U23262 (N_23262,N_22770,N_22918);
nand U23263 (N_23263,N_22613,N_23081);
nor U23264 (N_23264,N_22524,N_22921);
nor U23265 (N_23265,N_22683,N_22751);
and U23266 (N_23266,N_22842,N_22519);
or U23267 (N_23267,N_22619,N_22828);
and U23268 (N_23268,N_22544,N_23054);
nand U23269 (N_23269,N_23039,N_22892);
nand U23270 (N_23270,N_22768,N_22969);
xnor U23271 (N_23271,N_22851,N_22808);
xor U23272 (N_23272,N_22692,N_22795);
and U23273 (N_23273,N_22993,N_22744);
or U23274 (N_23274,N_22723,N_23080);
or U23275 (N_23275,N_22535,N_22718);
xor U23276 (N_23276,N_22627,N_22557);
nor U23277 (N_23277,N_22798,N_22707);
nand U23278 (N_23278,N_22879,N_22552);
and U23279 (N_23279,N_23038,N_22802);
or U23280 (N_23280,N_22840,N_22986);
nor U23281 (N_23281,N_22864,N_22903);
xnor U23282 (N_23282,N_22618,N_22525);
nand U23283 (N_23283,N_22947,N_22545);
nand U23284 (N_23284,N_23097,N_22705);
xor U23285 (N_23285,N_22639,N_22742);
nand U23286 (N_23286,N_22919,N_22868);
and U23287 (N_23287,N_22782,N_22605);
and U23288 (N_23288,N_22833,N_22827);
nor U23289 (N_23289,N_22555,N_22636);
nor U23290 (N_23290,N_23091,N_23048);
xor U23291 (N_23291,N_23041,N_22779);
nand U23292 (N_23292,N_22576,N_22528);
and U23293 (N_23293,N_22549,N_22905);
and U23294 (N_23294,N_22954,N_22701);
nand U23295 (N_23295,N_22728,N_22979);
nor U23296 (N_23296,N_22962,N_22594);
xnor U23297 (N_23297,N_22633,N_22712);
nand U23298 (N_23298,N_22970,N_22663);
xnor U23299 (N_23299,N_22658,N_22586);
nand U23300 (N_23300,N_22635,N_22772);
nor U23301 (N_23301,N_23113,N_22817);
xor U23302 (N_23302,N_23000,N_22711);
nand U23303 (N_23303,N_22603,N_22714);
xor U23304 (N_23304,N_22906,N_22815);
xnor U23305 (N_23305,N_22860,N_22596);
and U23306 (N_23306,N_22816,N_22501);
xnor U23307 (N_23307,N_22506,N_22516);
or U23308 (N_23308,N_22758,N_22813);
or U23309 (N_23309,N_22800,N_22794);
xor U23310 (N_23310,N_22526,N_22702);
nor U23311 (N_23311,N_22797,N_22505);
xor U23312 (N_23312,N_23037,N_22861);
nand U23313 (N_23313,N_22973,N_22942);
or U23314 (N_23314,N_22880,N_22599);
or U23315 (N_23315,N_22762,N_22671);
nand U23316 (N_23316,N_22713,N_23077);
xor U23317 (N_23317,N_22668,N_22883);
xnor U23318 (N_23318,N_23066,N_22585);
xor U23319 (N_23319,N_22551,N_23093);
nor U23320 (N_23320,N_23124,N_23090);
and U23321 (N_23321,N_23032,N_22887);
xor U23322 (N_23322,N_22621,N_23046);
and U23323 (N_23323,N_23086,N_22513);
and U23324 (N_23324,N_22791,N_22716);
and U23325 (N_23325,N_22852,N_22807);
or U23326 (N_23326,N_22821,N_22926);
and U23327 (N_23327,N_22748,N_22788);
or U23328 (N_23328,N_22715,N_23059);
or U23329 (N_23329,N_22786,N_22610);
nand U23330 (N_23330,N_22717,N_22564);
or U23331 (N_23331,N_22611,N_22743);
nor U23332 (N_23332,N_22536,N_23021);
or U23333 (N_23333,N_22561,N_22796);
and U23334 (N_23334,N_22626,N_23058);
nand U23335 (N_23335,N_22855,N_22523);
xor U23336 (N_23336,N_22972,N_22629);
xor U23337 (N_23337,N_22530,N_23008);
nand U23338 (N_23338,N_22991,N_22799);
nor U23339 (N_23339,N_22862,N_22700);
xnor U23340 (N_23340,N_22681,N_22566);
nand U23341 (N_23341,N_22559,N_22835);
and U23342 (N_23342,N_22955,N_22745);
and U23343 (N_23343,N_22568,N_22622);
and U23344 (N_23344,N_22598,N_22915);
nor U23345 (N_23345,N_22608,N_22569);
or U23346 (N_23346,N_22616,N_22741);
or U23347 (N_23347,N_22818,N_23100);
xor U23348 (N_23348,N_22625,N_22541);
and U23349 (N_23349,N_22912,N_22809);
xnor U23350 (N_23350,N_22783,N_22806);
and U23351 (N_23351,N_22537,N_23108);
or U23352 (N_23352,N_22988,N_22933);
or U23353 (N_23353,N_22882,N_22931);
nand U23354 (N_23354,N_23122,N_22706);
and U23355 (N_23355,N_22941,N_22948);
and U23356 (N_23356,N_22732,N_23009);
nand U23357 (N_23357,N_22560,N_22648);
or U23358 (N_23358,N_22583,N_23014);
nand U23359 (N_23359,N_23094,N_22830);
nand U23360 (N_23360,N_23123,N_22928);
and U23361 (N_23361,N_22510,N_22687);
or U23362 (N_23362,N_22675,N_23045);
nand U23363 (N_23363,N_22709,N_22810);
xnor U23364 (N_23364,N_22872,N_22747);
or U23365 (N_23365,N_22901,N_22959);
nand U23366 (N_23366,N_22884,N_23015);
xnor U23367 (N_23367,N_23089,N_22890);
or U23368 (N_23368,N_23109,N_22731);
or U23369 (N_23369,N_22646,N_23029);
nor U23370 (N_23370,N_22764,N_23071);
xnor U23371 (N_23371,N_22859,N_22812);
xnor U23372 (N_23372,N_22572,N_22682);
nand U23373 (N_23373,N_23102,N_22531);
and U23374 (N_23374,N_22548,N_22873);
nor U23375 (N_23375,N_22653,N_22759);
nor U23376 (N_23376,N_22688,N_22867);
nor U23377 (N_23377,N_23082,N_22512);
nand U23378 (N_23378,N_22678,N_22949);
nor U23379 (N_23379,N_22866,N_22554);
or U23380 (N_23380,N_22950,N_22604);
xnor U23381 (N_23381,N_22888,N_22515);
and U23382 (N_23382,N_22784,N_22848);
and U23383 (N_23383,N_22967,N_22672);
xnor U23384 (N_23384,N_22857,N_22869);
and U23385 (N_23385,N_22920,N_22769);
nand U23386 (N_23386,N_23119,N_22787);
nand U23387 (N_23387,N_23103,N_22760);
and U23388 (N_23388,N_22871,N_22781);
nor U23389 (N_23389,N_22579,N_22565);
xor U23390 (N_23390,N_23043,N_23099);
nand U23391 (N_23391,N_23049,N_22660);
and U23392 (N_23392,N_22936,N_22863);
or U23393 (N_23393,N_22754,N_23001);
and U23394 (N_23394,N_22623,N_22990);
nand U23395 (N_23395,N_22582,N_23055);
xor U23396 (N_23396,N_22538,N_22534);
xnor U23397 (N_23397,N_22875,N_22825);
nand U23398 (N_23398,N_22999,N_23079);
nor U23399 (N_23399,N_22661,N_23023);
xnor U23400 (N_23400,N_22775,N_23115);
xnor U23401 (N_23401,N_22773,N_22946);
and U23402 (N_23402,N_22823,N_22976);
and U23403 (N_23403,N_23019,N_22945);
xor U23404 (N_23404,N_23017,N_22591);
xnor U23405 (N_23405,N_22719,N_22587);
nand U23406 (N_23406,N_22520,N_22956);
nand U23407 (N_23407,N_22925,N_22638);
or U23408 (N_23408,N_22876,N_23016);
and U23409 (N_23409,N_22978,N_23053);
nand U23410 (N_23410,N_23106,N_22500);
or U23411 (N_23411,N_22899,N_22521);
or U23412 (N_23412,N_22563,N_22659);
xnor U23413 (N_23413,N_22982,N_22900);
and U23414 (N_23414,N_22965,N_23002);
and U23415 (N_23415,N_23012,N_23033);
nor U23416 (N_23416,N_22886,N_22514);
nor U23417 (N_23417,N_22614,N_22550);
xnor U23418 (N_23418,N_22647,N_23085);
and U23419 (N_23419,N_22624,N_22504);
nand U23420 (N_23420,N_22889,N_22834);
or U23421 (N_23421,N_23070,N_22953);
nor U23422 (N_23422,N_22529,N_22724);
nand U23423 (N_23423,N_22670,N_22938);
or U23424 (N_23424,N_22778,N_22845);
or U23425 (N_23425,N_22996,N_22593);
nor U23426 (N_23426,N_22935,N_23092);
xor U23427 (N_23427,N_22676,N_23004);
xnor U23428 (N_23428,N_22907,N_23060);
xor U23429 (N_23429,N_22601,N_23062);
nand U23430 (N_23430,N_22640,N_22917);
and U23431 (N_23431,N_22739,N_23064);
nor U23432 (N_23432,N_22761,N_22980);
nor U23433 (N_23433,N_22930,N_22750);
nand U23434 (N_23434,N_22814,N_23076);
or U23435 (N_23435,N_22590,N_22666);
nor U23436 (N_23436,N_23074,N_22740);
or U23437 (N_23437,N_22854,N_22718);
and U23438 (N_23438,N_22748,N_22892);
xor U23439 (N_23439,N_22854,N_23063);
nand U23440 (N_23440,N_22871,N_22646);
and U23441 (N_23441,N_22533,N_22586);
nor U23442 (N_23442,N_23085,N_22779);
xor U23443 (N_23443,N_22539,N_22536);
or U23444 (N_23444,N_22578,N_22848);
and U23445 (N_23445,N_23070,N_22588);
nand U23446 (N_23446,N_23077,N_22593);
xor U23447 (N_23447,N_22716,N_22651);
nand U23448 (N_23448,N_22503,N_22537);
nor U23449 (N_23449,N_23029,N_22502);
xnor U23450 (N_23450,N_23043,N_22840);
nand U23451 (N_23451,N_22873,N_22685);
nor U23452 (N_23452,N_22876,N_22999);
nand U23453 (N_23453,N_22782,N_22841);
nor U23454 (N_23454,N_22932,N_23050);
nand U23455 (N_23455,N_22666,N_22897);
nor U23456 (N_23456,N_23005,N_22935);
or U23457 (N_23457,N_22667,N_22942);
or U23458 (N_23458,N_22930,N_23055);
nand U23459 (N_23459,N_22904,N_22859);
nor U23460 (N_23460,N_23110,N_22973);
or U23461 (N_23461,N_22765,N_22975);
nand U23462 (N_23462,N_22621,N_22628);
nand U23463 (N_23463,N_22510,N_22537);
nor U23464 (N_23464,N_22974,N_22607);
nor U23465 (N_23465,N_22556,N_23121);
nand U23466 (N_23466,N_22889,N_23111);
or U23467 (N_23467,N_22546,N_22896);
nor U23468 (N_23468,N_22642,N_22584);
nand U23469 (N_23469,N_22950,N_22744);
or U23470 (N_23470,N_22593,N_22573);
nor U23471 (N_23471,N_22616,N_23001);
and U23472 (N_23472,N_23091,N_23004);
nand U23473 (N_23473,N_22628,N_22574);
and U23474 (N_23474,N_23007,N_22748);
xor U23475 (N_23475,N_22518,N_23012);
nand U23476 (N_23476,N_22612,N_22800);
nor U23477 (N_23477,N_22858,N_22833);
nor U23478 (N_23478,N_22808,N_22998);
or U23479 (N_23479,N_22614,N_22886);
and U23480 (N_23480,N_22896,N_22519);
or U23481 (N_23481,N_23053,N_22728);
xor U23482 (N_23482,N_23011,N_23014);
nor U23483 (N_23483,N_23083,N_22754);
and U23484 (N_23484,N_23055,N_23122);
nor U23485 (N_23485,N_22561,N_22786);
xnor U23486 (N_23486,N_22990,N_22515);
and U23487 (N_23487,N_22947,N_22848);
and U23488 (N_23488,N_22606,N_23042);
nand U23489 (N_23489,N_22919,N_22723);
and U23490 (N_23490,N_22962,N_23027);
and U23491 (N_23491,N_22606,N_22936);
or U23492 (N_23492,N_22881,N_22675);
nand U23493 (N_23493,N_22603,N_22517);
nor U23494 (N_23494,N_22884,N_23095);
or U23495 (N_23495,N_22634,N_22515);
nand U23496 (N_23496,N_22955,N_22871);
nand U23497 (N_23497,N_22528,N_22523);
nor U23498 (N_23498,N_22755,N_23112);
nor U23499 (N_23499,N_22701,N_22672);
xnor U23500 (N_23500,N_22785,N_22868);
nor U23501 (N_23501,N_22568,N_22560);
nor U23502 (N_23502,N_22660,N_22554);
nand U23503 (N_23503,N_22951,N_22543);
nor U23504 (N_23504,N_22738,N_22769);
and U23505 (N_23505,N_22787,N_22879);
and U23506 (N_23506,N_23062,N_22535);
nor U23507 (N_23507,N_22691,N_22983);
and U23508 (N_23508,N_22506,N_23006);
and U23509 (N_23509,N_23035,N_22580);
xnor U23510 (N_23510,N_22733,N_22815);
xor U23511 (N_23511,N_22923,N_22932);
or U23512 (N_23512,N_22640,N_23049);
or U23513 (N_23513,N_22824,N_22543);
nor U23514 (N_23514,N_22888,N_23026);
nand U23515 (N_23515,N_22781,N_22628);
nand U23516 (N_23516,N_22953,N_22954);
xor U23517 (N_23517,N_22505,N_22743);
nand U23518 (N_23518,N_22804,N_22926);
nor U23519 (N_23519,N_22528,N_22899);
and U23520 (N_23520,N_22558,N_23107);
nand U23521 (N_23521,N_22624,N_22606);
xnor U23522 (N_23522,N_22902,N_22553);
and U23523 (N_23523,N_22522,N_23023);
or U23524 (N_23524,N_22741,N_22503);
xor U23525 (N_23525,N_22610,N_22948);
nand U23526 (N_23526,N_22697,N_22740);
nand U23527 (N_23527,N_22817,N_22834);
nand U23528 (N_23528,N_22980,N_22599);
nor U23529 (N_23529,N_22904,N_23013);
nand U23530 (N_23530,N_22917,N_22630);
xor U23531 (N_23531,N_23048,N_22591);
and U23532 (N_23532,N_22770,N_22929);
nor U23533 (N_23533,N_22526,N_22947);
nor U23534 (N_23534,N_22943,N_23049);
nor U23535 (N_23535,N_23075,N_22561);
and U23536 (N_23536,N_23082,N_23057);
or U23537 (N_23537,N_23089,N_22853);
and U23538 (N_23538,N_22688,N_22514);
nor U23539 (N_23539,N_22617,N_22718);
and U23540 (N_23540,N_22790,N_23094);
nor U23541 (N_23541,N_22899,N_22943);
and U23542 (N_23542,N_22548,N_22993);
nor U23543 (N_23543,N_22627,N_22962);
or U23544 (N_23544,N_22978,N_22581);
or U23545 (N_23545,N_22807,N_22974);
or U23546 (N_23546,N_23111,N_22733);
and U23547 (N_23547,N_23010,N_22933);
or U23548 (N_23548,N_22774,N_22868);
nand U23549 (N_23549,N_23033,N_22729);
or U23550 (N_23550,N_22694,N_22741);
and U23551 (N_23551,N_22613,N_22789);
or U23552 (N_23552,N_23089,N_22972);
and U23553 (N_23553,N_22752,N_23077);
or U23554 (N_23554,N_23014,N_22812);
nor U23555 (N_23555,N_22525,N_22544);
or U23556 (N_23556,N_23064,N_22750);
nor U23557 (N_23557,N_22746,N_23050);
nor U23558 (N_23558,N_22882,N_23080);
or U23559 (N_23559,N_22615,N_23026);
or U23560 (N_23560,N_22646,N_23015);
nor U23561 (N_23561,N_22993,N_22697);
nor U23562 (N_23562,N_22719,N_22674);
xor U23563 (N_23563,N_22887,N_23042);
xor U23564 (N_23564,N_22816,N_22697);
nand U23565 (N_23565,N_22655,N_22639);
nor U23566 (N_23566,N_22554,N_22988);
or U23567 (N_23567,N_23098,N_22879);
and U23568 (N_23568,N_22771,N_23097);
or U23569 (N_23569,N_22546,N_22775);
xor U23570 (N_23570,N_22668,N_22805);
or U23571 (N_23571,N_22579,N_23017);
or U23572 (N_23572,N_22554,N_22602);
xor U23573 (N_23573,N_22872,N_22893);
and U23574 (N_23574,N_22674,N_22936);
or U23575 (N_23575,N_22815,N_22659);
or U23576 (N_23576,N_22701,N_22775);
xor U23577 (N_23577,N_22959,N_22566);
or U23578 (N_23578,N_22789,N_22973);
nand U23579 (N_23579,N_22833,N_22685);
xor U23580 (N_23580,N_22849,N_23086);
or U23581 (N_23581,N_23116,N_23120);
nor U23582 (N_23582,N_23028,N_22834);
nand U23583 (N_23583,N_22695,N_22927);
and U23584 (N_23584,N_22617,N_22803);
xnor U23585 (N_23585,N_22733,N_22971);
nor U23586 (N_23586,N_22878,N_22556);
xor U23587 (N_23587,N_22684,N_22607);
xnor U23588 (N_23588,N_23112,N_22611);
nand U23589 (N_23589,N_22924,N_22841);
or U23590 (N_23590,N_23041,N_22570);
or U23591 (N_23591,N_22709,N_22889);
nand U23592 (N_23592,N_22711,N_22823);
and U23593 (N_23593,N_22930,N_22982);
or U23594 (N_23594,N_22976,N_22622);
and U23595 (N_23595,N_23115,N_23006);
or U23596 (N_23596,N_22757,N_23097);
or U23597 (N_23597,N_22787,N_22728);
nand U23598 (N_23598,N_22554,N_22976);
nand U23599 (N_23599,N_22598,N_22945);
nor U23600 (N_23600,N_22702,N_22745);
xnor U23601 (N_23601,N_22978,N_22888);
xnor U23602 (N_23602,N_22866,N_23014);
nand U23603 (N_23603,N_22647,N_22652);
nor U23604 (N_23604,N_22708,N_23036);
and U23605 (N_23605,N_22630,N_22713);
nand U23606 (N_23606,N_22825,N_22665);
or U23607 (N_23607,N_22786,N_23061);
nor U23608 (N_23608,N_23023,N_22870);
nand U23609 (N_23609,N_22851,N_22799);
or U23610 (N_23610,N_23020,N_22997);
and U23611 (N_23611,N_22803,N_22618);
nor U23612 (N_23612,N_22735,N_22684);
or U23613 (N_23613,N_22512,N_23038);
nand U23614 (N_23614,N_22777,N_22687);
and U23615 (N_23615,N_23122,N_23034);
xnor U23616 (N_23616,N_22893,N_22952);
and U23617 (N_23617,N_22604,N_22628);
or U23618 (N_23618,N_22527,N_22667);
and U23619 (N_23619,N_22562,N_22692);
nor U23620 (N_23620,N_22945,N_22787);
or U23621 (N_23621,N_22981,N_22685);
nor U23622 (N_23622,N_22819,N_22805);
nor U23623 (N_23623,N_23059,N_22993);
xnor U23624 (N_23624,N_23096,N_23108);
nor U23625 (N_23625,N_22909,N_22683);
xor U23626 (N_23626,N_23114,N_22858);
nor U23627 (N_23627,N_22750,N_22577);
or U23628 (N_23628,N_22614,N_22768);
xnor U23629 (N_23629,N_22586,N_22957);
and U23630 (N_23630,N_22794,N_22696);
and U23631 (N_23631,N_22677,N_22672);
nor U23632 (N_23632,N_22552,N_22516);
xor U23633 (N_23633,N_22791,N_22656);
nor U23634 (N_23634,N_23048,N_23023);
nor U23635 (N_23635,N_22616,N_22829);
or U23636 (N_23636,N_22819,N_23113);
and U23637 (N_23637,N_22522,N_22826);
nand U23638 (N_23638,N_23053,N_22843);
nor U23639 (N_23639,N_22553,N_22668);
nor U23640 (N_23640,N_22838,N_23058);
or U23641 (N_23641,N_23001,N_22570);
xor U23642 (N_23642,N_22760,N_22812);
and U23643 (N_23643,N_22739,N_22864);
xnor U23644 (N_23644,N_23093,N_22918);
xnor U23645 (N_23645,N_22707,N_23008);
and U23646 (N_23646,N_22882,N_22530);
and U23647 (N_23647,N_22543,N_22680);
xnor U23648 (N_23648,N_22624,N_23002);
nand U23649 (N_23649,N_22948,N_22685);
xor U23650 (N_23650,N_23012,N_22940);
xor U23651 (N_23651,N_22665,N_22514);
and U23652 (N_23652,N_23002,N_22823);
and U23653 (N_23653,N_22874,N_22985);
nand U23654 (N_23654,N_23081,N_22545);
and U23655 (N_23655,N_22694,N_23016);
nor U23656 (N_23656,N_22762,N_22810);
xor U23657 (N_23657,N_22710,N_22909);
xor U23658 (N_23658,N_22919,N_22677);
and U23659 (N_23659,N_22516,N_22751);
or U23660 (N_23660,N_22803,N_23004);
and U23661 (N_23661,N_22951,N_23008);
nand U23662 (N_23662,N_23104,N_22692);
nand U23663 (N_23663,N_23075,N_23057);
or U23664 (N_23664,N_23102,N_22961);
and U23665 (N_23665,N_22959,N_23046);
nor U23666 (N_23666,N_22658,N_22743);
and U23667 (N_23667,N_23037,N_22807);
or U23668 (N_23668,N_22874,N_23035);
xnor U23669 (N_23669,N_22883,N_22860);
and U23670 (N_23670,N_23001,N_22973);
nor U23671 (N_23671,N_22556,N_22573);
and U23672 (N_23672,N_23062,N_23047);
nand U23673 (N_23673,N_22766,N_22821);
and U23674 (N_23674,N_23015,N_22907);
or U23675 (N_23675,N_22847,N_23074);
and U23676 (N_23676,N_23055,N_22657);
xnor U23677 (N_23677,N_22863,N_22500);
nand U23678 (N_23678,N_22797,N_22635);
nand U23679 (N_23679,N_23046,N_23096);
xor U23680 (N_23680,N_22739,N_22636);
nor U23681 (N_23681,N_22564,N_22660);
nor U23682 (N_23682,N_22525,N_22715);
xor U23683 (N_23683,N_22536,N_22772);
or U23684 (N_23684,N_22976,N_22643);
and U23685 (N_23685,N_22854,N_23124);
nor U23686 (N_23686,N_22734,N_22793);
and U23687 (N_23687,N_23065,N_22812);
xnor U23688 (N_23688,N_22724,N_23013);
and U23689 (N_23689,N_22885,N_22550);
or U23690 (N_23690,N_23068,N_22602);
or U23691 (N_23691,N_23012,N_23041);
nor U23692 (N_23692,N_23061,N_22660);
or U23693 (N_23693,N_23032,N_23112);
nand U23694 (N_23694,N_22935,N_22845);
xor U23695 (N_23695,N_22768,N_22747);
xnor U23696 (N_23696,N_22617,N_22950);
nand U23697 (N_23697,N_22695,N_22987);
nor U23698 (N_23698,N_23025,N_22551);
nand U23699 (N_23699,N_23049,N_22886);
or U23700 (N_23700,N_22826,N_22825);
xor U23701 (N_23701,N_23053,N_22568);
nor U23702 (N_23702,N_22571,N_23012);
and U23703 (N_23703,N_22707,N_23065);
and U23704 (N_23704,N_22532,N_22689);
nand U23705 (N_23705,N_23022,N_22560);
or U23706 (N_23706,N_22533,N_22805);
and U23707 (N_23707,N_23010,N_22577);
nand U23708 (N_23708,N_22721,N_22829);
nand U23709 (N_23709,N_22506,N_22616);
nor U23710 (N_23710,N_22550,N_22749);
nand U23711 (N_23711,N_22885,N_22580);
nand U23712 (N_23712,N_22817,N_22991);
nor U23713 (N_23713,N_22868,N_22566);
nor U23714 (N_23714,N_22632,N_23115);
xor U23715 (N_23715,N_22820,N_22896);
and U23716 (N_23716,N_22953,N_22944);
nand U23717 (N_23717,N_22797,N_22857);
nand U23718 (N_23718,N_22916,N_22767);
nand U23719 (N_23719,N_22539,N_22779);
and U23720 (N_23720,N_22620,N_22819);
xnor U23721 (N_23721,N_22803,N_23110);
xor U23722 (N_23722,N_22586,N_22988);
nor U23723 (N_23723,N_22709,N_22928);
nand U23724 (N_23724,N_22653,N_23071);
and U23725 (N_23725,N_22615,N_23108);
or U23726 (N_23726,N_22978,N_22983);
or U23727 (N_23727,N_22786,N_23085);
nor U23728 (N_23728,N_22678,N_23108);
or U23729 (N_23729,N_22864,N_23004);
nor U23730 (N_23730,N_22653,N_22805);
xor U23731 (N_23731,N_23121,N_23002);
nor U23732 (N_23732,N_23117,N_22899);
and U23733 (N_23733,N_23103,N_22519);
nor U23734 (N_23734,N_22962,N_22925);
or U23735 (N_23735,N_22794,N_23116);
and U23736 (N_23736,N_22507,N_22754);
nand U23737 (N_23737,N_22757,N_22631);
nor U23738 (N_23738,N_22568,N_23084);
or U23739 (N_23739,N_22746,N_22572);
nand U23740 (N_23740,N_22731,N_23041);
and U23741 (N_23741,N_23026,N_22885);
nor U23742 (N_23742,N_22603,N_22919);
nor U23743 (N_23743,N_22612,N_22995);
nand U23744 (N_23744,N_23028,N_22830);
or U23745 (N_23745,N_23046,N_22534);
and U23746 (N_23746,N_22867,N_22744);
xor U23747 (N_23747,N_23108,N_23053);
nand U23748 (N_23748,N_22870,N_22783);
or U23749 (N_23749,N_22510,N_22564);
nor U23750 (N_23750,N_23228,N_23621);
and U23751 (N_23751,N_23362,N_23534);
nor U23752 (N_23752,N_23277,N_23302);
or U23753 (N_23753,N_23505,N_23490);
xor U23754 (N_23754,N_23227,N_23522);
and U23755 (N_23755,N_23668,N_23198);
nor U23756 (N_23756,N_23253,N_23331);
nor U23757 (N_23757,N_23141,N_23563);
nand U23758 (N_23758,N_23244,N_23521);
nor U23759 (N_23759,N_23514,N_23680);
nor U23760 (N_23760,N_23164,N_23604);
nand U23761 (N_23761,N_23376,N_23530);
nand U23762 (N_23762,N_23600,N_23134);
xor U23763 (N_23763,N_23587,N_23207);
and U23764 (N_23764,N_23373,N_23155);
or U23765 (N_23765,N_23606,N_23154);
and U23766 (N_23766,N_23733,N_23489);
or U23767 (N_23767,N_23144,N_23455);
nor U23768 (N_23768,N_23409,N_23640);
xnor U23769 (N_23769,N_23510,N_23628);
or U23770 (N_23770,N_23473,N_23605);
nand U23771 (N_23771,N_23392,N_23463);
nand U23772 (N_23772,N_23433,N_23389);
or U23773 (N_23773,N_23629,N_23248);
or U23774 (N_23774,N_23745,N_23359);
or U23775 (N_23775,N_23709,N_23503);
and U23776 (N_23776,N_23718,N_23231);
nor U23777 (N_23777,N_23595,N_23625);
nor U23778 (N_23778,N_23260,N_23632);
nor U23779 (N_23779,N_23438,N_23249);
nand U23780 (N_23780,N_23345,N_23289);
nor U23781 (N_23781,N_23715,N_23700);
xnor U23782 (N_23782,N_23375,N_23497);
xor U23783 (N_23783,N_23222,N_23170);
xnor U23784 (N_23784,N_23265,N_23526);
nor U23785 (N_23785,N_23698,N_23471);
and U23786 (N_23786,N_23725,N_23517);
nand U23787 (N_23787,N_23255,N_23370);
and U23788 (N_23788,N_23435,N_23702);
nor U23789 (N_23789,N_23428,N_23531);
nand U23790 (N_23790,N_23315,N_23562);
nor U23791 (N_23791,N_23276,N_23529);
nor U23792 (N_23792,N_23127,N_23136);
or U23793 (N_23793,N_23727,N_23710);
nand U23794 (N_23794,N_23405,N_23568);
and U23795 (N_23795,N_23662,N_23535);
xnor U23796 (N_23796,N_23541,N_23193);
xnor U23797 (N_23797,N_23382,N_23180);
xor U23798 (N_23798,N_23706,N_23419);
or U23799 (N_23799,N_23195,N_23230);
and U23800 (N_23800,N_23267,N_23410);
or U23801 (N_23801,N_23128,N_23468);
xnor U23802 (N_23802,N_23746,N_23460);
nand U23803 (N_23803,N_23487,N_23571);
or U23804 (N_23804,N_23596,N_23318);
or U23805 (N_23805,N_23215,N_23555);
and U23806 (N_23806,N_23486,N_23140);
or U23807 (N_23807,N_23432,N_23186);
nand U23808 (N_23808,N_23300,N_23635);
nor U23809 (N_23809,N_23581,N_23399);
or U23810 (N_23810,N_23643,N_23556);
nor U23811 (N_23811,N_23146,N_23182);
and U23812 (N_23812,N_23566,N_23358);
nand U23813 (N_23813,N_23378,N_23386);
xor U23814 (N_23814,N_23618,N_23393);
and U23815 (N_23815,N_23694,N_23189);
and U23816 (N_23816,N_23678,N_23259);
xnor U23817 (N_23817,N_23360,N_23516);
nand U23818 (N_23818,N_23540,N_23308);
nand U23819 (N_23819,N_23368,N_23351);
or U23820 (N_23820,N_23691,N_23454);
nand U23821 (N_23821,N_23429,N_23477);
xor U23822 (N_23822,N_23594,N_23578);
xnor U23823 (N_23823,N_23731,N_23391);
nor U23824 (N_23824,N_23446,N_23258);
or U23825 (N_23825,N_23603,N_23188);
and U23826 (N_23826,N_23674,N_23537);
nor U23827 (N_23827,N_23655,N_23280);
and U23828 (N_23828,N_23576,N_23584);
nor U23829 (N_23829,N_23609,N_23321);
nor U23830 (N_23830,N_23169,N_23457);
or U23831 (N_23831,N_23427,N_23564);
xnor U23832 (N_23832,N_23695,N_23569);
nor U23833 (N_23833,N_23422,N_23398);
nand U23834 (N_23834,N_23724,N_23484);
nor U23835 (N_23835,N_23664,N_23325);
xnor U23836 (N_23836,N_23323,N_23583);
nand U23837 (N_23837,N_23273,N_23285);
nor U23838 (N_23838,N_23485,N_23340);
xor U23839 (N_23839,N_23671,N_23714);
nor U23840 (N_23840,N_23157,N_23565);
and U23841 (N_23841,N_23234,N_23172);
and U23842 (N_23842,N_23597,N_23243);
and U23843 (N_23843,N_23712,N_23349);
nand U23844 (N_23844,N_23713,N_23421);
nor U23845 (N_23845,N_23616,N_23403);
and U23846 (N_23846,N_23611,N_23573);
or U23847 (N_23847,N_23348,N_23675);
nor U23848 (N_23848,N_23708,N_23462);
xnor U23849 (N_23849,N_23570,N_23699);
nor U23850 (N_23850,N_23687,N_23167);
and U23851 (N_23851,N_23371,N_23685);
nor U23852 (N_23852,N_23523,N_23689);
and U23853 (N_23853,N_23210,N_23365);
nand U23854 (N_23854,N_23447,N_23173);
or U23855 (N_23855,N_23508,N_23139);
nand U23856 (N_23856,N_23147,N_23240);
xnor U23857 (N_23857,N_23175,N_23266);
nand U23858 (N_23858,N_23572,N_23475);
and U23859 (N_23859,N_23590,N_23720);
or U23860 (N_23860,N_23327,N_23636);
nand U23861 (N_23861,N_23661,N_23716);
or U23862 (N_23862,N_23663,N_23498);
xor U23863 (N_23863,N_23177,N_23434);
nor U23864 (N_23864,N_23294,N_23357);
nor U23865 (N_23865,N_23717,N_23693);
or U23866 (N_23866,N_23350,N_23202);
or U23867 (N_23867,N_23297,N_23395);
xor U23868 (N_23868,N_23622,N_23236);
and U23869 (N_23869,N_23748,N_23707);
or U23870 (N_23870,N_23247,N_23326);
xnor U23871 (N_23871,N_23466,N_23665);
and U23872 (N_23872,N_23319,N_23178);
xor U23873 (N_23873,N_23613,N_23203);
and U23874 (N_23874,N_23322,N_23408);
xnor U23875 (N_23875,N_23450,N_23268);
or U23876 (N_23876,N_23374,N_23579);
and U23877 (N_23877,N_23402,N_23347);
xnor U23878 (N_23878,N_23567,N_23291);
and U23879 (N_23879,N_23528,N_23533);
nand U23880 (N_23880,N_23418,N_23299);
nand U23881 (N_23881,N_23292,N_23580);
xnor U23882 (N_23882,N_23238,N_23316);
and U23883 (N_23883,N_23330,N_23163);
nand U23884 (N_23884,N_23204,N_23246);
or U23885 (N_23885,N_23191,N_23549);
and U23886 (N_23886,N_23610,N_23153);
and U23887 (N_23887,N_23271,N_23728);
nand U23888 (N_23888,N_23184,N_23211);
nor U23889 (N_23889,N_23631,N_23217);
nand U23890 (N_23890,N_23262,N_23352);
nand U23891 (N_23891,N_23361,N_23406);
nand U23892 (N_23892,N_23546,N_23667);
or U23893 (N_23893,N_23200,N_23254);
nand U23894 (N_23894,N_23179,N_23619);
xor U23895 (N_23895,N_23142,N_23132);
nand U23896 (N_23896,N_23197,N_23684);
nor U23897 (N_23897,N_23647,N_23317);
xor U23898 (N_23898,N_23151,N_23270);
xor U23899 (N_23899,N_23282,N_23582);
or U23900 (N_23900,N_23506,N_23697);
or U23901 (N_23901,N_23135,N_23721);
or U23902 (N_23902,N_23656,N_23453);
xnor U23903 (N_23903,N_23591,N_23367);
and U23904 (N_23904,N_23500,N_23303);
nor U23905 (N_23905,N_23666,N_23653);
nand U23906 (N_23906,N_23743,N_23617);
nand U23907 (N_23907,N_23288,N_23379);
nor U23908 (N_23908,N_23612,N_23608);
xor U23909 (N_23909,N_23320,N_23607);
or U23910 (N_23910,N_23654,N_23310);
nor U23911 (N_23911,N_23440,N_23328);
or U23912 (N_23912,N_23290,N_23601);
nor U23913 (N_23913,N_23233,N_23148);
nor U23914 (N_23914,N_23423,N_23458);
xor U23915 (N_23915,N_23162,N_23554);
xor U23916 (N_23916,N_23729,N_23441);
or U23917 (N_23917,N_23474,N_23174);
xor U23918 (N_23918,N_23201,N_23354);
or U23919 (N_23919,N_23221,N_23353);
nand U23920 (N_23920,N_23602,N_23652);
or U23921 (N_23921,N_23638,N_23387);
and U23922 (N_23922,N_23150,N_23336);
or U23923 (N_23923,N_23261,N_23559);
and U23924 (N_23924,N_23278,N_23125);
nand U23925 (N_23925,N_23305,N_23333);
and U23926 (N_23926,N_23673,N_23232);
nand U23927 (N_23927,N_23385,N_23677);
and U23928 (N_23928,N_23511,N_23187);
nand U23929 (N_23929,N_23158,N_23730);
and U23930 (N_23930,N_23483,N_23314);
xnor U23931 (N_23931,N_23479,N_23682);
nand U23932 (N_23932,N_23627,N_23459);
or U23933 (N_23933,N_23513,N_23557);
xnor U23934 (N_23934,N_23214,N_23126);
or U23935 (N_23935,N_23704,N_23205);
nand U23936 (N_23936,N_23738,N_23472);
or U23937 (N_23937,N_23329,N_23465);
and U23938 (N_23938,N_23646,N_23507);
nand U23939 (N_23939,N_23156,N_23334);
nand U23940 (N_23940,N_23469,N_23431);
or U23941 (N_23941,N_23493,N_23660);
nand U23942 (N_23942,N_23363,N_23364);
or U23943 (N_23943,N_23192,N_23548);
xnor U23944 (N_23944,N_23341,N_23190);
nand U23945 (N_23945,N_23377,N_23492);
nand U23946 (N_23946,N_23426,N_23245);
and U23947 (N_23947,N_23380,N_23298);
or U23948 (N_23948,N_23586,N_23194);
and U23949 (N_23949,N_23442,N_23252);
nand U23950 (N_23950,N_23553,N_23723);
nand U23951 (N_23951,N_23509,N_23552);
nand U23952 (N_23952,N_23676,N_23400);
or U23953 (N_23953,N_23149,N_23165);
and U23954 (N_23954,N_23335,N_23551);
or U23955 (N_23955,N_23223,N_23213);
or U23956 (N_23956,N_23133,N_23742);
and U23957 (N_23957,N_23496,N_23219);
and U23958 (N_23958,N_23577,N_23525);
nor U23959 (N_23959,N_23589,N_23574);
or U23960 (N_23960,N_23131,N_23160);
or U23961 (N_23961,N_23722,N_23383);
nor U23962 (N_23962,N_23518,N_23279);
and U23963 (N_23963,N_23739,N_23623);
nand U23964 (N_23964,N_23550,N_23626);
nand U23965 (N_23965,N_23332,N_23287);
and U23966 (N_23966,N_23237,N_23649);
or U23967 (N_23967,N_23401,N_23199);
nor U23968 (N_23968,N_23338,N_23679);
and U23969 (N_23969,N_23416,N_23539);
xor U23970 (N_23970,N_23543,N_23672);
or U23971 (N_23971,N_23143,N_23407);
or U23972 (N_23972,N_23394,N_23670);
nand U23973 (N_23973,N_23532,N_23196);
or U23974 (N_23974,N_23747,N_23634);
nand U23975 (N_23975,N_23286,N_23744);
nor U23976 (N_23976,N_23536,N_23235);
nor U23977 (N_23977,N_23415,N_23615);
and U23978 (N_23978,N_23560,N_23637);
nand U23979 (N_23979,N_23397,N_23212);
or U23980 (N_23980,N_23688,N_23501);
or U23981 (N_23981,N_23159,N_23339);
and U23982 (N_23982,N_23686,N_23711);
xor U23983 (N_23983,N_23451,N_23137);
xnor U23984 (N_23984,N_23575,N_23185);
or U23985 (N_23985,N_23424,N_23545);
and U23986 (N_23986,N_23512,N_23592);
nor U23987 (N_23987,N_23251,N_23313);
and U23988 (N_23988,N_23735,N_23726);
nor U23989 (N_23989,N_23547,N_23476);
xor U23990 (N_23990,N_23425,N_23515);
or U23991 (N_23991,N_23456,N_23161);
and U23992 (N_23992,N_23208,N_23482);
nand U23993 (N_23993,N_23741,N_23130);
nand U23994 (N_23994,N_23183,N_23369);
nand U23995 (N_23995,N_23256,N_23705);
nor U23996 (N_23996,N_23176,N_23439);
xnor U23997 (N_23997,N_23464,N_23239);
nor U23998 (N_23998,N_23593,N_23404);
nor U23999 (N_23999,N_23411,N_23620);
xor U24000 (N_24000,N_23225,N_23312);
and U24001 (N_24001,N_23650,N_23413);
nand U24002 (N_24002,N_23412,N_23448);
nand U24003 (N_24003,N_23337,N_23491);
nor U24004 (N_24004,N_23443,N_23430);
xor U24005 (N_24005,N_23372,N_23558);
nand U24006 (N_24006,N_23599,N_23502);
or U24007 (N_24007,N_23274,N_23633);
xor U24008 (N_24008,N_23478,N_23216);
and U24009 (N_24009,N_23293,N_23467);
and U24010 (N_24010,N_23701,N_23346);
or U24011 (N_24011,N_23740,N_23309);
nand U24012 (N_24012,N_23311,N_23324);
nor U24013 (N_24013,N_23356,N_23561);
nand U24014 (N_24014,N_23381,N_23520);
nand U24015 (N_24015,N_23296,N_23295);
or U24016 (N_24016,N_23749,N_23719);
nor U24017 (N_24017,N_23639,N_23734);
or U24018 (N_24018,N_23272,N_23226);
nand U24019 (N_24019,N_23538,N_23692);
xor U24020 (N_24020,N_23269,N_23304);
nand U24021 (N_24021,N_23171,N_23414);
or U24022 (N_24022,N_23281,N_23301);
nand U24023 (N_24023,N_23499,N_23452);
xnor U24024 (N_24024,N_23696,N_23470);
and U24025 (N_24025,N_23651,N_23614);
or U24026 (N_24026,N_23544,N_23461);
xor U24027 (N_24027,N_23284,N_23657);
or U24028 (N_24028,N_23642,N_23396);
and U24029 (N_24029,N_23275,N_23669);
and U24030 (N_24030,N_23645,N_23481);
xor U24031 (N_24031,N_23736,N_23307);
and U24032 (N_24032,N_23263,N_23181);
or U24033 (N_24033,N_23220,N_23737);
or U24034 (N_24034,N_23138,N_23644);
xor U24035 (N_24035,N_23504,N_23366);
xnor U24036 (N_24036,N_23585,N_23519);
xor U24037 (N_24037,N_23658,N_23264);
xnor U24038 (N_24038,N_23641,N_23524);
xnor U24039 (N_24039,N_23343,N_23436);
nor U24040 (N_24040,N_23598,N_23449);
nand U24041 (N_24041,N_23242,N_23206);
nand U24042 (N_24042,N_23229,N_23417);
nor U24043 (N_24043,N_23542,N_23480);
xor U24044 (N_24044,N_23344,N_23257);
or U24045 (N_24045,N_23444,N_23437);
nand U24046 (N_24046,N_23648,N_23494);
xnor U24047 (N_24047,N_23384,N_23703);
nor U24048 (N_24048,N_23683,N_23224);
or U24049 (N_24049,N_23732,N_23390);
xor U24050 (N_24050,N_23355,N_23152);
and U24051 (N_24051,N_23306,N_23145);
or U24052 (N_24052,N_23588,N_23166);
xor U24053 (N_24053,N_23445,N_23250);
nor U24054 (N_24054,N_23129,N_23630);
or U24055 (N_24055,N_23681,N_23218);
nand U24056 (N_24056,N_23624,N_23659);
and U24057 (N_24057,N_23388,N_23168);
nor U24058 (N_24058,N_23527,N_23690);
nor U24059 (N_24059,N_23488,N_23283);
and U24060 (N_24060,N_23241,N_23342);
nor U24061 (N_24061,N_23209,N_23495);
nand U24062 (N_24062,N_23420,N_23530);
nand U24063 (N_24063,N_23332,N_23578);
nand U24064 (N_24064,N_23447,N_23484);
nand U24065 (N_24065,N_23231,N_23732);
xnor U24066 (N_24066,N_23208,N_23675);
nor U24067 (N_24067,N_23142,N_23542);
and U24068 (N_24068,N_23610,N_23552);
or U24069 (N_24069,N_23739,N_23335);
and U24070 (N_24070,N_23547,N_23513);
or U24071 (N_24071,N_23640,N_23708);
nand U24072 (N_24072,N_23622,N_23166);
xnor U24073 (N_24073,N_23156,N_23737);
nand U24074 (N_24074,N_23360,N_23143);
or U24075 (N_24075,N_23735,N_23495);
nor U24076 (N_24076,N_23597,N_23278);
or U24077 (N_24077,N_23673,N_23672);
and U24078 (N_24078,N_23465,N_23251);
nor U24079 (N_24079,N_23260,N_23561);
xnor U24080 (N_24080,N_23478,N_23379);
nand U24081 (N_24081,N_23443,N_23250);
nor U24082 (N_24082,N_23294,N_23458);
nor U24083 (N_24083,N_23238,N_23211);
xnor U24084 (N_24084,N_23601,N_23716);
nor U24085 (N_24085,N_23194,N_23266);
or U24086 (N_24086,N_23468,N_23139);
and U24087 (N_24087,N_23653,N_23483);
nor U24088 (N_24088,N_23344,N_23700);
or U24089 (N_24089,N_23433,N_23130);
xor U24090 (N_24090,N_23746,N_23517);
nor U24091 (N_24091,N_23620,N_23128);
or U24092 (N_24092,N_23324,N_23265);
xor U24093 (N_24093,N_23512,N_23517);
nor U24094 (N_24094,N_23149,N_23129);
nor U24095 (N_24095,N_23418,N_23633);
nor U24096 (N_24096,N_23210,N_23177);
and U24097 (N_24097,N_23399,N_23275);
nand U24098 (N_24098,N_23716,N_23608);
xnor U24099 (N_24099,N_23378,N_23130);
or U24100 (N_24100,N_23614,N_23484);
nor U24101 (N_24101,N_23425,N_23294);
xor U24102 (N_24102,N_23514,N_23294);
xnor U24103 (N_24103,N_23448,N_23718);
nand U24104 (N_24104,N_23171,N_23233);
nor U24105 (N_24105,N_23586,N_23665);
nor U24106 (N_24106,N_23125,N_23385);
nor U24107 (N_24107,N_23171,N_23426);
or U24108 (N_24108,N_23159,N_23266);
xnor U24109 (N_24109,N_23600,N_23523);
nand U24110 (N_24110,N_23710,N_23374);
or U24111 (N_24111,N_23410,N_23268);
or U24112 (N_24112,N_23354,N_23591);
nor U24113 (N_24113,N_23550,N_23732);
or U24114 (N_24114,N_23549,N_23234);
nand U24115 (N_24115,N_23572,N_23162);
and U24116 (N_24116,N_23419,N_23575);
nand U24117 (N_24117,N_23475,N_23576);
xor U24118 (N_24118,N_23286,N_23136);
nor U24119 (N_24119,N_23483,N_23636);
or U24120 (N_24120,N_23247,N_23720);
or U24121 (N_24121,N_23449,N_23250);
and U24122 (N_24122,N_23563,N_23143);
xnor U24123 (N_24123,N_23236,N_23547);
nand U24124 (N_24124,N_23588,N_23420);
xnor U24125 (N_24125,N_23569,N_23647);
nand U24126 (N_24126,N_23201,N_23149);
nor U24127 (N_24127,N_23616,N_23410);
xnor U24128 (N_24128,N_23313,N_23259);
and U24129 (N_24129,N_23463,N_23520);
nor U24130 (N_24130,N_23320,N_23354);
nand U24131 (N_24131,N_23681,N_23473);
xnor U24132 (N_24132,N_23191,N_23241);
xor U24133 (N_24133,N_23298,N_23165);
nor U24134 (N_24134,N_23253,N_23681);
and U24135 (N_24135,N_23462,N_23141);
and U24136 (N_24136,N_23425,N_23461);
and U24137 (N_24137,N_23277,N_23679);
xnor U24138 (N_24138,N_23583,N_23543);
xnor U24139 (N_24139,N_23436,N_23532);
or U24140 (N_24140,N_23715,N_23353);
nor U24141 (N_24141,N_23334,N_23646);
and U24142 (N_24142,N_23217,N_23336);
and U24143 (N_24143,N_23483,N_23723);
xnor U24144 (N_24144,N_23186,N_23694);
nand U24145 (N_24145,N_23432,N_23282);
xor U24146 (N_24146,N_23410,N_23246);
or U24147 (N_24147,N_23224,N_23400);
and U24148 (N_24148,N_23494,N_23128);
xor U24149 (N_24149,N_23276,N_23239);
xnor U24150 (N_24150,N_23566,N_23442);
nor U24151 (N_24151,N_23380,N_23351);
nor U24152 (N_24152,N_23496,N_23630);
nor U24153 (N_24153,N_23261,N_23487);
nand U24154 (N_24154,N_23147,N_23269);
nor U24155 (N_24155,N_23225,N_23214);
nor U24156 (N_24156,N_23157,N_23549);
and U24157 (N_24157,N_23432,N_23269);
xnor U24158 (N_24158,N_23357,N_23567);
or U24159 (N_24159,N_23528,N_23515);
xnor U24160 (N_24160,N_23369,N_23548);
and U24161 (N_24161,N_23526,N_23200);
nand U24162 (N_24162,N_23736,N_23571);
and U24163 (N_24163,N_23661,N_23446);
or U24164 (N_24164,N_23196,N_23478);
nand U24165 (N_24165,N_23331,N_23553);
or U24166 (N_24166,N_23133,N_23549);
or U24167 (N_24167,N_23476,N_23200);
and U24168 (N_24168,N_23620,N_23318);
nor U24169 (N_24169,N_23537,N_23302);
xor U24170 (N_24170,N_23747,N_23602);
nor U24171 (N_24171,N_23366,N_23658);
or U24172 (N_24172,N_23555,N_23623);
xor U24173 (N_24173,N_23151,N_23711);
xor U24174 (N_24174,N_23580,N_23721);
and U24175 (N_24175,N_23447,N_23525);
nor U24176 (N_24176,N_23293,N_23280);
and U24177 (N_24177,N_23428,N_23458);
or U24178 (N_24178,N_23447,N_23308);
and U24179 (N_24179,N_23405,N_23417);
nand U24180 (N_24180,N_23520,N_23704);
and U24181 (N_24181,N_23305,N_23487);
or U24182 (N_24182,N_23684,N_23718);
nor U24183 (N_24183,N_23188,N_23319);
and U24184 (N_24184,N_23671,N_23390);
and U24185 (N_24185,N_23451,N_23246);
nor U24186 (N_24186,N_23414,N_23266);
xor U24187 (N_24187,N_23339,N_23550);
nor U24188 (N_24188,N_23289,N_23153);
or U24189 (N_24189,N_23277,N_23427);
or U24190 (N_24190,N_23291,N_23208);
or U24191 (N_24191,N_23296,N_23701);
and U24192 (N_24192,N_23665,N_23155);
nor U24193 (N_24193,N_23646,N_23294);
and U24194 (N_24194,N_23323,N_23245);
or U24195 (N_24195,N_23246,N_23232);
nand U24196 (N_24196,N_23622,N_23564);
and U24197 (N_24197,N_23695,N_23292);
or U24198 (N_24198,N_23175,N_23531);
or U24199 (N_24199,N_23326,N_23576);
and U24200 (N_24200,N_23143,N_23307);
xnor U24201 (N_24201,N_23686,N_23176);
xnor U24202 (N_24202,N_23162,N_23238);
nand U24203 (N_24203,N_23316,N_23312);
or U24204 (N_24204,N_23515,N_23181);
and U24205 (N_24205,N_23226,N_23554);
nand U24206 (N_24206,N_23171,N_23597);
nor U24207 (N_24207,N_23216,N_23673);
and U24208 (N_24208,N_23392,N_23610);
nor U24209 (N_24209,N_23273,N_23600);
and U24210 (N_24210,N_23439,N_23595);
nor U24211 (N_24211,N_23183,N_23640);
or U24212 (N_24212,N_23688,N_23330);
nor U24213 (N_24213,N_23587,N_23358);
nor U24214 (N_24214,N_23535,N_23267);
nor U24215 (N_24215,N_23374,N_23164);
nor U24216 (N_24216,N_23155,N_23213);
or U24217 (N_24217,N_23638,N_23491);
xnor U24218 (N_24218,N_23363,N_23154);
nand U24219 (N_24219,N_23355,N_23582);
xor U24220 (N_24220,N_23339,N_23520);
nand U24221 (N_24221,N_23665,N_23416);
and U24222 (N_24222,N_23205,N_23383);
nor U24223 (N_24223,N_23421,N_23400);
xor U24224 (N_24224,N_23648,N_23745);
and U24225 (N_24225,N_23329,N_23194);
nand U24226 (N_24226,N_23331,N_23483);
nor U24227 (N_24227,N_23288,N_23578);
or U24228 (N_24228,N_23534,N_23441);
or U24229 (N_24229,N_23624,N_23623);
xor U24230 (N_24230,N_23746,N_23485);
xor U24231 (N_24231,N_23263,N_23171);
xor U24232 (N_24232,N_23390,N_23513);
nand U24233 (N_24233,N_23536,N_23364);
nand U24234 (N_24234,N_23446,N_23380);
and U24235 (N_24235,N_23390,N_23177);
and U24236 (N_24236,N_23656,N_23151);
or U24237 (N_24237,N_23552,N_23618);
and U24238 (N_24238,N_23534,N_23257);
and U24239 (N_24239,N_23289,N_23678);
nand U24240 (N_24240,N_23748,N_23360);
nand U24241 (N_24241,N_23545,N_23492);
or U24242 (N_24242,N_23644,N_23146);
nand U24243 (N_24243,N_23569,N_23540);
and U24244 (N_24244,N_23244,N_23311);
or U24245 (N_24245,N_23345,N_23253);
xnor U24246 (N_24246,N_23748,N_23578);
or U24247 (N_24247,N_23564,N_23441);
xnor U24248 (N_24248,N_23594,N_23358);
xnor U24249 (N_24249,N_23596,N_23201);
and U24250 (N_24250,N_23230,N_23253);
or U24251 (N_24251,N_23128,N_23734);
nand U24252 (N_24252,N_23548,N_23681);
or U24253 (N_24253,N_23724,N_23379);
nor U24254 (N_24254,N_23700,N_23496);
and U24255 (N_24255,N_23200,N_23300);
nor U24256 (N_24256,N_23423,N_23192);
nor U24257 (N_24257,N_23391,N_23144);
nand U24258 (N_24258,N_23332,N_23364);
or U24259 (N_24259,N_23549,N_23714);
and U24260 (N_24260,N_23272,N_23154);
nor U24261 (N_24261,N_23295,N_23192);
xor U24262 (N_24262,N_23516,N_23397);
or U24263 (N_24263,N_23569,N_23570);
xnor U24264 (N_24264,N_23483,N_23421);
nand U24265 (N_24265,N_23472,N_23167);
or U24266 (N_24266,N_23293,N_23213);
and U24267 (N_24267,N_23187,N_23420);
nand U24268 (N_24268,N_23528,N_23529);
xnor U24269 (N_24269,N_23700,N_23363);
nand U24270 (N_24270,N_23155,N_23552);
xnor U24271 (N_24271,N_23480,N_23392);
nand U24272 (N_24272,N_23542,N_23414);
and U24273 (N_24273,N_23338,N_23416);
or U24274 (N_24274,N_23553,N_23383);
xnor U24275 (N_24275,N_23737,N_23214);
nor U24276 (N_24276,N_23669,N_23204);
nand U24277 (N_24277,N_23734,N_23195);
xor U24278 (N_24278,N_23410,N_23590);
and U24279 (N_24279,N_23294,N_23651);
xor U24280 (N_24280,N_23542,N_23289);
xnor U24281 (N_24281,N_23185,N_23193);
nor U24282 (N_24282,N_23612,N_23432);
and U24283 (N_24283,N_23125,N_23206);
and U24284 (N_24284,N_23430,N_23478);
nand U24285 (N_24285,N_23599,N_23373);
and U24286 (N_24286,N_23482,N_23569);
xor U24287 (N_24287,N_23641,N_23237);
nand U24288 (N_24288,N_23672,N_23519);
xor U24289 (N_24289,N_23690,N_23705);
nor U24290 (N_24290,N_23578,N_23227);
or U24291 (N_24291,N_23163,N_23306);
and U24292 (N_24292,N_23526,N_23676);
and U24293 (N_24293,N_23593,N_23656);
or U24294 (N_24294,N_23704,N_23239);
and U24295 (N_24295,N_23375,N_23134);
or U24296 (N_24296,N_23713,N_23219);
nand U24297 (N_24297,N_23175,N_23219);
and U24298 (N_24298,N_23435,N_23737);
nor U24299 (N_24299,N_23422,N_23379);
or U24300 (N_24300,N_23306,N_23714);
or U24301 (N_24301,N_23725,N_23605);
or U24302 (N_24302,N_23578,N_23422);
xor U24303 (N_24303,N_23274,N_23717);
xnor U24304 (N_24304,N_23453,N_23546);
and U24305 (N_24305,N_23715,N_23615);
nor U24306 (N_24306,N_23563,N_23277);
nor U24307 (N_24307,N_23689,N_23567);
xnor U24308 (N_24308,N_23738,N_23348);
and U24309 (N_24309,N_23168,N_23736);
nor U24310 (N_24310,N_23199,N_23438);
xnor U24311 (N_24311,N_23659,N_23662);
or U24312 (N_24312,N_23281,N_23706);
nor U24313 (N_24313,N_23429,N_23716);
nor U24314 (N_24314,N_23452,N_23323);
and U24315 (N_24315,N_23193,N_23282);
nor U24316 (N_24316,N_23249,N_23298);
nand U24317 (N_24317,N_23214,N_23240);
or U24318 (N_24318,N_23608,N_23478);
nor U24319 (N_24319,N_23691,N_23409);
or U24320 (N_24320,N_23183,N_23667);
or U24321 (N_24321,N_23641,N_23282);
nand U24322 (N_24322,N_23489,N_23523);
nor U24323 (N_24323,N_23622,N_23552);
nand U24324 (N_24324,N_23575,N_23650);
xor U24325 (N_24325,N_23216,N_23730);
nand U24326 (N_24326,N_23639,N_23529);
nand U24327 (N_24327,N_23308,N_23555);
or U24328 (N_24328,N_23429,N_23206);
nor U24329 (N_24329,N_23319,N_23387);
and U24330 (N_24330,N_23273,N_23405);
xnor U24331 (N_24331,N_23584,N_23223);
xor U24332 (N_24332,N_23615,N_23213);
or U24333 (N_24333,N_23471,N_23392);
or U24334 (N_24334,N_23578,N_23263);
nand U24335 (N_24335,N_23653,N_23279);
xor U24336 (N_24336,N_23516,N_23442);
nand U24337 (N_24337,N_23244,N_23171);
nor U24338 (N_24338,N_23423,N_23479);
nor U24339 (N_24339,N_23218,N_23429);
nand U24340 (N_24340,N_23606,N_23290);
nand U24341 (N_24341,N_23232,N_23619);
nor U24342 (N_24342,N_23715,N_23271);
xor U24343 (N_24343,N_23582,N_23250);
nor U24344 (N_24344,N_23404,N_23300);
or U24345 (N_24345,N_23649,N_23379);
and U24346 (N_24346,N_23500,N_23425);
and U24347 (N_24347,N_23430,N_23556);
nand U24348 (N_24348,N_23428,N_23154);
nand U24349 (N_24349,N_23333,N_23509);
and U24350 (N_24350,N_23739,N_23389);
and U24351 (N_24351,N_23573,N_23688);
nor U24352 (N_24352,N_23412,N_23541);
nand U24353 (N_24353,N_23284,N_23443);
and U24354 (N_24354,N_23356,N_23424);
xnor U24355 (N_24355,N_23749,N_23397);
or U24356 (N_24356,N_23382,N_23343);
and U24357 (N_24357,N_23364,N_23301);
and U24358 (N_24358,N_23134,N_23573);
nor U24359 (N_24359,N_23435,N_23553);
or U24360 (N_24360,N_23548,N_23419);
or U24361 (N_24361,N_23289,N_23275);
nor U24362 (N_24362,N_23174,N_23733);
and U24363 (N_24363,N_23286,N_23693);
nand U24364 (N_24364,N_23157,N_23412);
xor U24365 (N_24365,N_23362,N_23493);
or U24366 (N_24366,N_23655,N_23127);
nor U24367 (N_24367,N_23477,N_23221);
and U24368 (N_24368,N_23137,N_23280);
nor U24369 (N_24369,N_23222,N_23313);
nor U24370 (N_24370,N_23362,N_23620);
xnor U24371 (N_24371,N_23585,N_23261);
nand U24372 (N_24372,N_23723,N_23281);
nor U24373 (N_24373,N_23239,N_23695);
nand U24374 (N_24374,N_23306,N_23674);
xnor U24375 (N_24375,N_24114,N_24181);
and U24376 (N_24376,N_23983,N_23822);
xor U24377 (N_24377,N_24041,N_24169);
nand U24378 (N_24378,N_24118,N_24321);
xnor U24379 (N_24379,N_24028,N_23935);
nor U24380 (N_24380,N_24127,N_23933);
and U24381 (N_24381,N_24162,N_23898);
and U24382 (N_24382,N_24361,N_24348);
xor U24383 (N_24383,N_23814,N_24196);
and U24384 (N_24384,N_24094,N_23950);
xor U24385 (N_24385,N_24136,N_23896);
xnor U24386 (N_24386,N_24235,N_24208);
or U24387 (N_24387,N_24243,N_24066);
or U24388 (N_24388,N_23886,N_24197);
or U24389 (N_24389,N_24357,N_24022);
xnor U24390 (N_24390,N_23903,N_23978);
nor U24391 (N_24391,N_24339,N_24313);
nor U24392 (N_24392,N_24077,N_24112);
nor U24393 (N_24393,N_24190,N_24288);
xnor U24394 (N_24394,N_24371,N_24219);
nand U24395 (N_24395,N_23956,N_24001);
xnor U24396 (N_24396,N_24218,N_23947);
or U24397 (N_24397,N_23995,N_24257);
nand U24398 (N_24398,N_24278,N_24252);
and U24399 (N_24399,N_23805,N_23877);
and U24400 (N_24400,N_24170,N_24141);
and U24401 (N_24401,N_23803,N_24042);
nor U24402 (N_24402,N_23952,N_23884);
and U24403 (N_24403,N_24120,N_24263);
or U24404 (N_24404,N_23908,N_24211);
and U24405 (N_24405,N_24036,N_24049);
or U24406 (N_24406,N_23821,N_24315);
xnor U24407 (N_24407,N_24018,N_24093);
nand U24408 (N_24408,N_24126,N_24152);
or U24409 (N_24409,N_24102,N_23824);
and U24410 (N_24410,N_23869,N_24054);
nor U24411 (N_24411,N_24097,N_24091);
nor U24412 (N_24412,N_24100,N_24177);
or U24413 (N_24413,N_23763,N_23872);
nor U24414 (N_24414,N_24200,N_24241);
nand U24415 (N_24415,N_23948,N_24184);
and U24416 (N_24416,N_23813,N_23895);
or U24417 (N_24417,N_24106,N_24167);
nor U24418 (N_24418,N_24341,N_23918);
or U24419 (N_24419,N_23907,N_24233);
xor U24420 (N_24420,N_24282,N_24021);
xor U24421 (N_24421,N_24205,N_24363);
nor U24422 (N_24422,N_24270,N_24227);
xnor U24423 (N_24423,N_23919,N_24063);
nor U24424 (N_24424,N_24207,N_23917);
or U24425 (N_24425,N_23836,N_23980);
or U24426 (N_24426,N_24366,N_23960);
and U24427 (N_24427,N_23755,N_24119);
or U24428 (N_24428,N_24080,N_24217);
and U24429 (N_24429,N_23963,N_24151);
or U24430 (N_24430,N_24327,N_24139);
and U24431 (N_24431,N_23796,N_24192);
xnor U24432 (N_24432,N_24116,N_23901);
or U24433 (N_24433,N_24230,N_24331);
nand U24434 (N_24434,N_24237,N_23991);
and U24435 (N_24435,N_23799,N_24103);
and U24436 (N_24436,N_23875,N_23847);
or U24437 (N_24437,N_24277,N_24368);
nand U24438 (N_24438,N_24369,N_24265);
or U24439 (N_24439,N_23756,N_24229);
xor U24440 (N_24440,N_24342,N_23856);
nand U24441 (N_24441,N_24292,N_24158);
or U24442 (N_24442,N_23988,N_24283);
nand U24443 (N_24443,N_23904,N_24068);
nand U24444 (N_24444,N_24291,N_24006);
nand U24445 (N_24445,N_24074,N_24259);
nor U24446 (N_24446,N_24231,N_24053);
xor U24447 (N_24447,N_23926,N_24032);
and U24448 (N_24448,N_23859,N_24297);
nand U24449 (N_24449,N_24084,N_24221);
xor U24450 (N_24450,N_23806,N_23764);
nor U24451 (N_24451,N_24212,N_24060);
or U24452 (N_24452,N_23964,N_24232);
nand U24453 (N_24453,N_23757,N_24191);
and U24454 (N_24454,N_24113,N_24069);
nand U24455 (N_24455,N_23913,N_24023);
and U24456 (N_24456,N_24347,N_24198);
and U24457 (N_24457,N_23879,N_24135);
and U24458 (N_24458,N_24145,N_24256);
and U24459 (N_24459,N_24002,N_23826);
nand U24460 (N_24460,N_23928,N_23934);
nand U24461 (N_24461,N_23795,N_23953);
or U24462 (N_24462,N_24294,N_24076);
nand U24463 (N_24463,N_24370,N_24214);
or U24464 (N_24464,N_23999,N_24209);
nor U24465 (N_24465,N_23974,N_24007);
or U24466 (N_24466,N_24360,N_23835);
or U24467 (N_24467,N_24155,N_24226);
nand U24468 (N_24468,N_23954,N_23838);
or U24469 (N_24469,N_24253,N_24086);
or U24470 (N_24470,N_24104,N_24314);
or U24471 (N_24471,N_24350,N_24052);
or U24472 (N_24472,N_24316,N_24272);
nand U24473 (N_24473,N_24298,N_24183);
nor U24474 (N_24474,N_24260,N_24025);
xor U24475 (N_24475,N_24279,N_24228);
or U24476 (N_24476,N_23979,N_23998);
nand U24477 (N_24477,N_23900,N_24012);
nor U24478 (N_24478,N_23914,N_23930);
nand U24479 (N_24479,N_24179,N_24062);
and U24480 (N_24480,N_23870,N_24180);
nand U24481 (N_24481,N_24204,N_24009);
or U24482 (N_24482,N_23842,N_23815);
nand U24483 (N_24483,N_23792,N_23833);
nor U24484 (N_24484,N_24334,N_23811);
or U24485 (N_24485,N_23817,N_24333);
and U24486 (N_24486,N_23894,N_24317);
nor U24487 (N_24487,N_24193,N_23897);
xnor U24488 (N_24488,N_24329,N_23990);
and U24489 (N_24489,N_24195,N_24171);
nand U24490 (N_24490,N_24199,N_23882);
nand U24491 (N_24491,N_23832,N_23768);
or U24492 (N_24492,N_24345,N_24300);
nor U24493 (N_24493,N_24132,N_23911);
nand U24494 (N_24494,N_24020,N_24040);
or U24495 (N_24495,N_23986,N_23861);
nand U24496 (N_24496,N_24311,N_24138);
xor U24497 (N_24497,N_23767,N_24129);
nor U24498 (N_24498,N_24134,N_24019);
or U24499 (N_24499,N_23965,N_24045);
and U24500 (N_24500,N_23831,N_24144);
xor U24501 (N_24501,N_24206,N_23854);
xor U24502 (N_24502,N_24051,N_23762);
or U24503 (N_24503,N_24261,N_23899);
and U24504 (N_24504,N_24318,N_23793);
xnor U24505 (N_24505,N_23985,N_24026);
and U24506 (N_24506,N_24072,N_24343);
nand U24507 (N_24507,N_23779,N_23946);
and U24508 (N_24508,N_24295,N_24299);
nor U24509 (N_24509,N_24372,N_24148);
and U24510 (N_24510,N_23807,N_24030);
nand U24511 (N_24511,N_23987,N_24223);
and U24512 (N_24512,N_23924,N_24070);
xor U24513 (N_24513,N_24353,N_24065);
nand U24514 (N_24514,N_23945,N_24143);
xor U24515 (N_24515,N_23876,N_23912);
and U24516 (N_24516,N_23932,N_23994);
nor U24517 (N_24517,N_24137,N_23841);
xnor U24518 (N_24518,N_24146,N_24269);
nor U24519 (N_24519,N_23959,N_24271);
nand U24520 (N_24520,N_24203,N_24024);
and U24521 (N_24521,N_24149,N_24367);
and U24522 (N_24522,N_24014,N_24073);
nand U24523 (N_24523,N_24373,N_23750);
or U24524 (N_24524,N_24248,N_23883);
nand U24525 (N_24525,N_23783,N_23961);
and U24526 (N_24526,N_24098,N_23864);
nor U24527 (N_24527,N_24039,N_23789);
nand U24528 (N_24528,N_24322,N_23939);
and U24529 (N_24529,N_24320,N_24255);
or U24530 (N_24530,N_24164,N_23816);
nor U24531 (N_24531,N_23906,N_24185);
xor U24532 (N_24532,N_23851,N_23808);
xor U24533 (N_24533,N_23798,N_23885);
xnor U24534 (N_24534,N_24307,N_23850);
or U24535 (N_24535,N_23958,N_23858);
and U24536 (N_24536,N_23992,N_24029);
or U24537 (N_24537,N_23794,N_24122);
or U24538 (N_24538,N_24374,N_24044);
xnor U24539 (N_24539,N_23938,N_24109);
nor U24540 (N_24540,N_24325,N_23868);
nor U24541 (N_24541,N_24013,N_23774);
xor U24542 (N_24542,N_24038,N_24356);
and U24543 (N_24543,N_24275,N_23787);
and U24544 (N_24544,N_23775,N_24175);
xnor U24545 (N_24545,N_24095,N_24274);
nand U24546 (N_24546,N_24050,N_23893);
xor U24547 (N_24547,N_24215,N_23971);
nor U24548 (N_24548,N_23828,N_24273);
xor U24549 (N_24549,N_23997,N_23830);
and U24550 (N_24550,N_24332,N_23916);
or U24551 (N_24551,N_24128,N_24107);
or U24552 (N_24552,N_23848,N_23878);
nor U24553 (N_24553,N_24092,N_24238);
or U24554 (N_24554,N_23927,N_24188);
and U24555 (N_24555,N_24121,N_23780);
xor U24556 (N_24556,N_23818,N_24064);
xor U24557 (N_24557,N_24174,N_23923);
nand U24558 (N_24558,N_24234,N_24306);
nand U24559 (N_24559,N_24005,N_23951);
nand U24560 (N_24560,N_24096,N_24017);
and U24561 (N_24561,N_24035,N_23782);
or U24562 (N_24562,N_24239,N_24281);
nor U24563 (N_24563,N_24210,N_23769);
xor U24564 (N_24564,N_24078,N_24166);
nand U24565 (N_24565,N_24312,N_24082);
xnor U24566 (N_24566,N_23888,N_23845);
nor U24567 (N_24567,N_24133,N_24186);
or U24568 (N_24568,N_24015,N_23863);
or U24569 (N_24569,N_24266,N_23966);
xnor U24570 (N_24570,N_24157,N_23976);
and U24571 (N_24571,N_24189,N_24236);
xnor U24572 (N_24572,N_23860,N_23855);
xnor U24573 (N_24573,N_23819,N_23772);
nor U24574 (N_24574,N_24124,N_23837);
nor U24575 (N_24575,N_24301,N_23777);
nand U24576 (N_24576,N_24033,N_24027);
or U24577 (N_24577,N_24123,N_24287);
or U24578 (N_24578,N_23871,N_24090);
nor U24579 (N_24579,N_23849,N_23989);
nand U24580 (N_24580,N_23993,N_24289);
nor U24581 (N_24581,N_23944,N_24355);
and U24582 (N_24582,N_24081,N_24351);
xor U24583 (N_24583,N_23902,N_23873);
xor U24584 (N_24584,N_24016,N_23910);
nand U24585 (N_24585,N_23843,N_24099);
and U24586 (N_24586,N_23754,N_24088);
and U24587 (N_24587,N_23791,N_23827);
or U24588 (N_24588,N_24147,N_23776);
nor U24589 (N_24589,N_24303,N_23778);
nor U24590 (N_24590,N_24326,N_24108);
nand U24591 (N_24591,N_23970,N_24328);
nand U24592 (N_24592,N_24250,N_24358);
and U24593 (N_24593,N_24365,N_24349);
nand U24594 (N_24594,N_23874,N_24222);
nor U24595 (N_24595,N_23751,N_23981);
nand U24596 (N_24596,N_24089,N_23786);
xnor U24597 (N_24597,N_24296,N_24059);
and U24598 (N_24598,N_24220,N_23825);
or U24599 (N_24599,N_24061,N_24354);
nor U24600 (N_24600,N_24224,N_23829);
nand U24601 (N_24601,N_23760,N_24110);
xnor U24602 (N_24602,N_24131,N_24225);
or U24603 (N_24603,N_24153,N_24340);
nor U24604 (N_24604,N_23852,N_24216);
xnor U24605 (N_24605,N_24242,N_23909);
or U24606 (N_24606,N_24346,N_23820);
nor U24607 (N_24607,N_24163,N_23801);
or U24608 (N_24608,N_24037,N_23844);
and U24609 (N_24609,N_23785,N_24267);
nor U24610 (N_24610,N_24364,N_23810);
nand U24611 (N_24611,N_24031,N_24067);
and U24612 (N_24612,N_23834,N_23969);
nand U24613 (N_24613,N_24304,N_23770);
nor U24614 (N_24614,N_24285,N_24034);
nor U24615 (N_24615,N_23846,N_23889);
nand U24616 (N_24616,N_24330,N_24240);
or U24617 (N_24617,N_24308,N_24249);
nor U24618 (N_24618,N_24178,N_24105);
or U24619 (N_24619,N_23771,N_24160);
nor U24620 (N_24620,N_23920,N_24008);
nor U24621 (N_24621,N_24173,N_24182);
nand U24622 (N_24622,N_24359,N_24338);
xnor U24623 (N_24623,N_24056,N_24362);
xnor U24624 (N_24624,N_24310,N_24154);
and U24625 (N_24625,N_24245,N_24286);
or U24626 (N_24626,N_23941,N_23865);
and U24627 (N_24627,N_23881,N_24055);
or U24628 (N_24628,N_24202,N_23968);
or U24629 (N_24629,N_24150,N_23784);
or U24630 (N_24630,N_23857,N_24058);
nor U24631 (N_24631,N_24319,N_24057);
nor U24632 (N_24632,N_23758,N_23890);
or U24633 (N_24633,N_24048,N_23892);
or U24634 (N_24634,N_24323,N_23977);
and U24635 (N_24635,N_23800,N_23891);
nor U24636 (N_24636,N_23967,N_23973);
nor U24637 (N_24637,N_23802,N_23972);
nand U24638 (N_24638,N_24262,N_24337);
and U24639 (N_24639,N_24004,N_23936);
nand U24640 (N_24640,N_23996,N_23839);
or U24641 (N_24641,N_23942,N_24258);
and U24642 (N_24642,N_24156,N_23880);
or U24643 (N_24643,N_23790,N_24111);
and U24644 (N_24644,N_24117,N_23921);
xor U24645 (N_24645,N_23797,N_24244);
or U24646 (N_24646,N_23781,N_23940);
xor U24647 (N_24647,N_24142,N_23812);
xnor U24648 (N_24648,N_23943,N_23823);
nor U24649 (N_24649,N_24293,N_24011);
xor U24650 (N_24650,N_24125,N_24290);
nor U24651 (N_24651,N_23925,N_23862);
nor U24652 (N_24652,N_23929,N_24079);
xor U24653 (N_24653,N_24043,N_23761);
and U24654 (N_24654,N_24336,N_24000);
xnor U24655 (N_24655,N_23866,N_24335);
nor U24656 (N_24656,N_23853,N_23962);
nor U24657 (N_24657,N_24115,N_23753);
nand U24658 (N_24658,N_24087,N_24010);
or U24659 (N_24659,N_23887,N_24159);
or U24660 (N_24660,N_24305,N_23867);
nor U24661 (N_24661,N_24176,N_24213);
or U24662 (N_24662,N_23765,N_24101);
xor U24663 (N_24663,N_23931,N_23905);
xor U24664 (N_24664,N_24276,N_24352);
and U24665 (N_24665,N_24083,N_24130);
nor U24666 (N_24666,N_24085,N_23773);
nor U24667 (N_24667,N_24264,N_23752);
nor U24668 (N_24668,N_23840,N_23955);
nand U24669 (N_24669,N_23982,N_23975);
or U24670 (N_24670,N_24324,N_24046);
nor U24671 (N_24671,N_24254,N_24194);
nor U24672 (N_24672,N_23937,N_24047);
xor U24673 (N_24673,N_24201,N_23766);
xnor U24674 (N_24674,N_23915,N_24075);
nor U24675 (N_24675,N_24140,N_24168);
and U24676 (N_24676,N_24165,N_24187);
nor U24677 (N_24677,N_24172,N_24302);
nor U24678 (N_24678,N_24284,N_23759);
nor U24679 (N_24679,N_23804,N_24247);
and U24680 (N_24680,N_23957,N_23984);
or U24681 (N_24681,N_23788,N_24161);
xnor U24682 (N_24682,N_24268,N_24071);
or U24683 (N_24683,N_23922,N_23949);
nor U24684 (N_24684,N_23809,N_24251);
or U24685 (N_24685,N_24344,N_24280);
nor U24686 (N_24686,N_24309,N_24003);
xor U24687 (N_24687,N_24246,N_24320);
nand U24688 (N_24688,N_24354,N_23901);
xnor U24689 (N_24689,N_24245,N_23769);
and U24690 (N_24690,N_24280,N_24048);
and U24691 (N_24691,N_23898,N_23929);
or U24692 (N_24692,N_24206,N_23789);
nor U24693 (N_24693,N_23923,N_24229);
nor U24694 (N_24694,N_23966,N_23977);
nand U24695 (N_24695,N_23992,N_23797);
nor U24696 (N_24696,N_23756,N_23803);
xor U24697 (N_24697,N_24189,N_23829);
nand U24698 (N_24698,N_24042,N_24328);
or U24699 (N_24699,N_24235,N_24341);
nand U24700 (N_24700,N_24066,N_24024);
and U24701 (N_24701,N_23824,N_24251);
xor U24702 (N_24702,N_24367,N_23776);
xnor U24703 (N_24703,N_24001,N_23862);
and U24704 (N_24704,N_24006,N_24146);
and U24705 (N_24705,N_24108,N_24001);
xor U24706 (N_24706,N_24351,N_23942);
or U24707 (N_24707,N_23784,N_24199);
or U24708 (N_24708,N_24327,N_24197);
or U24709 (N_24709,N_23909,N_24116);
nor U24710 (N_24710,N_23807,N_24148);
xnor U24711 (N_24711,N_24190,N_24220);
or U24712 (N_24712,N_24171,N_23864);
nor U24713 (N_24713,N_23791,N_24360);
nor U24714 (N_24714,N_24322,N_24174);
nand U24715 (N_24715,N_24093,N_24042);
and U24716 (N_24716,N_24258,N_23926);
or U24717 (N_24717,N_23856,N_23965);
nor U24718 (N_24718,N_24028,N_23761);
or U24719 (N_24719,N_24315,N_24260);
and U24720 (N_24720,N_23875,N_24220);
nor U24721 (N_24721,N_23899,N_23809);
xnor U24722 (N_24722,N_23771,N_24126);
and U24723 (N_24723,N_24216,N_23846);
xnor U24724 (N_24724,N_24334,N_23793);
or U24725 (N_24725,N_23820,N_24034);
nand U24726 (N_24726,N_24185,N_24298);
xor U24727 (N_24727,N_24070,N_23914);
nand U24728 (N_24728,N_24321,N_24091);
nor U24729 (N_24729,N_24252,N_23843);
nand U24730 (N_24730,N_24278,N_23891);
xor U24731 (N_24731,N_24164,N_24306);
or U24732 (N_24732,N_24121,N_24024);
xnor U24733 (N_24733,N_24088,N_24042);
or U24734 (N_24734,N_24263,N_24176);
nor U24735 (N_24735,N_23957,N_23772);
nand U24736 (N_24736,N_24199,N_24118);
or U24737 (N_24737,N_24350,N_24002);
or U24738 (N_24738,N_23884,N_24068);
xnor U24739 (N_24739,N_24033,N_24149);
and U24740 (N_24740,N_24041,N_24145);
nor U24741 (N_24741,N_23844,N_23775);
and U24742 (N_24742,N_24165,N_23854);
nor U24743 (N_24743,N_23885,N_23950);
nand U24744 (N_24744,N_24024,N_23873);
or U24745 (N_24745,N_24254,N_23768);
nand U24746 (N_24746,N_24328,N_24037);
or U24747 (N_24747,N_24166,N_24311);
and U24748 (N_24748,N_23954,N_23977);
nor U24749 (N_24749,N_24018,N_24142);
nor U24750 (N_24750,N_23818,N_23843);
and U24751 (N_24751,N_24010,N_24272);
nor U24752 (N_24752,N_24057,N_24218);
nand U24753 (N_24753,N_24122,N_23913);
or U24754 (N_24754,N_24101,N_23807);
and U24755 (N_24755,N_24087,N_23943);
and U24756 (N_24756,N_24230,N_23892);
and U24757 (N_24757,N_24289,N_24339);
nand U24758 (N_24758,N_24159,N_23863);
or U24759 (N_24759,N_24294,N_24355);
or U24760 (N_24760,N_23975,N_23802);
xnor U24761 (N_24761,N_24154,N_23862);
nand U24762 (N_24762,N_24363,N_24151);
xnor U24763 (N_24763,N_24210,N_23789);
and U24764 (N_24764,N_24301,N_24104);
xnor U24765 (N_24765,N_24241,N_24089);
nand U24766 (N_24766,N_23858,N_24325);
nor U24767 (N_24767,N_24026,N_24314);
and U24768 (N_24768,N_24164,N_23994);
xnor U24769 (N_24769,N_24303,N_24239);
xor U24770 (N_24770,N_24294,N_24138);
or U24771 (N_24771,N_24283,N_23958);
nor U24772 (N_24772,N_24293,N_24313);
nand U24773 (N_24773,N_24098,N_24338);
xor U24774 (N_24774,N_24346,N_23858);
and U24775 (N_24775,N_23800,N_23775);
nand U24776 (N_24776,N_23860,N_24034);
xor U24777 (N_24777,N_24181,N_24298);
nor U24778 (N_24778,N_24348,N_24350);
nand U24779 (N_24779,N_23892,N_24360);
and U24780 (N_24780,N_23831,N_23756);
or U24781 (N_24781,N_23859,N_23771);
and U24782 (N_24782,N_24116,N_24178);
nor U24783 (N_24783,N_23795,N_24323);
or U24784 (N_24784,N_24164,N_24047);
or U24785 (N_24785,N_23783,N_23826);
nand U24786 (N_24786,N_24150,N_24155);
and U24787 (N_24787,N_23769,N_24137);
and U24788 (N_24788,N_24011,N_24371);
and U24789 (N_24789,N_23959,N_23978);
or U24790 (N_24790,N_23968,N_23901);
or U24791 (N_24791,N_24144,N_24217);
nor U24792 (N_24792,N_23890,N_23919);
or U24793 (N_24793,N_23981,N_24139);
and U24794 (N_24794,N_23843,N_23950);
xnor U24795 (N_24795,N_24206,N_24151);
nand U24796 (N_24796,N_24323,N_24109);
and U24797 (N_24797,N_24270,N_23978);
nor U24798 (N_24798,N_24203,N_24116);
nor U24799 (N_24799,N_24085,N_23852);
or U24800 (N_24800,N_24234,N_24107);
nand U24801 (N_24801,N_24326,N_23864);
nor U24802 (N_24802,N_24195,N_23821);
nor U24803 (N_24803,N_23949,N_24011);
and U24804 (N_24804,N_23785,N_24232);
nor U24805 (N_24805,N_23855,N_23853);
or U24806 (N_24806,N_23811,N_24259);
xor U24807 (N_24807,N_24366,N_23805);
nand U24808 (N_24808,N_24353,N_24066);
xor U24809 (N_24809,N_23843,N_23885);
and U24810 (N_24810,N_24117,N_24202);
or U24811 (N_24811,N_23866,N_24033);
or U24812 (N_24812,N_24321,N_24274);
nand U24813 (N_24813,N_23937,N_23880);
and U24814 (N_24814,N_23909,N_24278);
xor U24815 (N_24815,N_24160,N_23898);
or U24816 (N_24816,N_24133,N_24164);
nand U24817 (N_24817,N_23872,N_23767);
nand U24818 (N_24818,N_23960,N_24320);
xor U24819 (N_24819,N_24228,N_24305);
nor U24820 (N_24820,N_23938,N_24361);
nor U24821 (N_24821,N_24279,N_24352);
xnor U24822 (N_24822,N_24054,N_24209);
or U24823 (N_24823,N_24018,N_24138);
and U24824 (N_24824,N_23848,N_23772);
nor U24825 (N_24825,N_24207,N_23931);
and U24826 (N_24826,N_23986,N_24244);
nor U24827 (N_24827,N_24114,N_24251);
xnor U24828 (N_24828,N_23986,N_23886);
nor U24829 (N_24829,N_23998,N_24116);
or U24830 (N_24830,N_24152,N_24280);
and U24831 (N_24831,N_24284,N_24164);
xor U24832 (N_24832,N_23844,N_23996);
and U24833 (N_24833,N_24052,N_24182);
nor U24834 (N_24834,N_23936,N_23996);
nand U24835 (N_24835,N_23845,N_24203);
nand U24836 (N_24836,N_23939,N_24148);
xnor U24837 (N_24837,N_24236,N_23908);
nand U24838 (N_24838,N_24154,N_24097);
and U24839 (N_24839,N_24300,N_24351);
nand U24840 (N_24840,N_23998,N_24014);
nor U24841 (N_24841,N_24323,N_24025);
nand U24842 (N_24842,N_24123,N_23832);
nand U24843 (N_24843,N_24189,N_24207);
and U24844 (N_24844,N_24233,N_24186);
or U24845 (N_24845,N_24300,N_24316);
nand U24846 (N_24846,N_23998,N_24056);
nand U24847 (N_24847,N_24326,N_23835);
xor U24848 (N_24848,N_24125,N_24087);
nand U24849 (N_24849,N_24225,N_23823);
xnor U24850 (N_24850,N_23889,N_24259);
xnor U24851 (N_24851,N_24090,N_23982);
or U24852 (N_24852,N_24040,N_24300);
and U24853 (N_24853,N_23918,N_24363);
nand U24854 (N_24854,N_24191,N_24373);
or U24855 (N_24855,N_24114,N_24066);
nor U24856 (N_24856,N_24006,N_23835);
or U24857 (N_24857,N_24170,N_23930);
nor U24858 (N_24858,N_24363,N_24055);
or U24859 (N_24859,N_24292,N_24363);
and U24860 (N_24860,N_24030,N_24250);
nor U24861 (N_24861,N_23934,N_24203);
xor U24862 (N_24862,N_24127,N_24336);
and U24863 (N_24863,N_23861,N_23865);
xor U24864 (N_24864,N_24180,N_23823);
nor U24865 (N_24865,N_24204,N_23923);
and U24866 (N_24866,N_24287,N_23832);
and U24867 (N_24867,N_23926,N_24121);
xor U24868 (N_24868,N_23928,N_23753);
xor U24869 (N_24869,N_24194,N_24089);
and U24870 (N_24870,N_24151,N_23784);
or U24871 (N_24871,N_24372,N_23806);
nand U24872 (N_24872,N_24332,N_24046);
nand U24873 (N_24873,N_24102,N_24234);
and U24874 (N_24874,N_24320,N_24100);
nor U24875 (N_24875,N_24346,N_24242);
nor U24876 (N_24876,N_24229,N_23767);
or U24877 (N_24877,N_24363,N_24019);
nor U24878 (N_24878,N_24229,N_24359);
nor U24879 (N_24879,N_23828,N_24351);
nor U24880 (N_24880,N_23780,N_24317);
or U24881 (N_24881,N_23753,N_23888);
or U24882 (N_24882,N_23915,N_23930);
nor U24883 (N_24883,N_24366,N_23923);
and U24884 (N_24884,N_24132,N_24293);
nand U24885 (N_24885,N_23751,N_23945);
nand U24886 (N_24886,N_23764,N_23881);
xnor U24887 (N_24887,N_23985,N_23847);
xor U24888 (N_24888,N_24155,N_23970);
xor U24889 (N_24889,N_24165,N_24048);
nand U24890 (N_24890,N_23806,N_23910);
nand U24891 (N_24891,N_24047,N_24205);
xor U24892 (N_24892,N_24057,N_23759);
nand U24893 (N_24893,N_24023,N_24239);
xor U24894 (N_24894,N_24324,N_24131);
nor U24895 (N_24895,N_24231,N_23916);
or U24896 (N_24896,N_24329,N_24094);
nor U24897 (N_24897,N_23999,N_24290);
xor U24898 (N_24898,N_24099,N_24095);
and U24899 (N_24899,N_23954,N_24373);
nor U24900 (N_24900,N_24132,N_24241);
or U24901 (N_24901,N_23972,N_24189);
or U24902 (N_24902,N_23834,N_23756);
nor U24903 (N_24903,N_24266,N_24374);
xor U24904 (N_24904,N_23753,N_24063);
xor U24905 (N_24905,N_24082,N_23908);
or U24906 (N_24906,N_23781,N_24009);
or U24907 (N_24907,N_23911,N_24140);
nor U24908 (N_24908,N_23901,N_23837);
or U24909 (N_24909,N_24279,N_24169);
nor U24910 (N_24910,N_23824,N_24325);
nor U24911 (N_24911,N_24066,N_23793);
nand U24912 (N_24912,N_24170,N_23781);
and U24913 (N_24913,N_23996,N_23981);
nand U24914 (N_24914,N_23812,N_24297);
xnor U24915 (N_24915,N_24232,N_24030);
xor U24916 (N_24916,N_23888,N_24077);
nor U24917 (N_24917,N_23825,N_23807);
xor U24918 (N_24918,N_23862,N_24150);
xnor U24919 (N_24919,N_24303,N_23770);
nor U24920 (N_24920,N_24272,N_23891);
or U24921 (N_24921,N_24287,N_24003);
nor U24922 (N_24922,N_24072,N_23837);
nor U24923 (N_24923,N_24202,N_24214);
nor U24924 (N_24924,N_24076,N_24083);
xnor U24925 (N_24925,N_24131,N_23971);
nor U24926 (N_24926,N_23904,N_24314);
and U24927 (N_24927,N_24120,N_24169);
nor U24928 (N_24928,N_24113,N_24089);
and U24929 (N_24929,N_24039,N_24292);
nor U24930 (N_24930,N_23772,N_24059);
xor U24931 (N_24931,N_23946,N_23912);
and U24932 (N_24932,N_24182,N_23761);
nor U24933 (N_24933,N_24140,N_23880);
nand U24934 (N_24934,N_24311,N_23950);
nand U24935 (N_24935,N_23805,N_23823);
nor U24936 (N_24936,N_23770,N_24189);
or U24937 (N_24937,N_23804,N_24203);
nand U24938 (N_24938,N_23802,N_23920);
nand U24939 (N_24939,N_24069,N_23961);
nand U24940 (N_24940,N_23861,N_24199);
and U24941 (N_24941,N_24054,N_24057);
or U24942 (N_24942,N_23995,N_23876);
or U24943 (N_24943,N_24356,N_23989);
nand U24944 (N_24944,N_24262,N_24272);
and U24945 (N_24945,N_23963,N_24082);
or U24946 (N_24946,N_24305,N_23977);
or U24947 (N_24947,N_24076,N_24090);
nand U24948 (N_24948,N_24366,N_24056);
xor U24949 (N_24949,N_23868,N_24123);
xnor U24950 (N_24950,N_24115,N_24063);
and U24951 (N_24951,N_24332,N_24073);
xor U24952 (N_24952,N_24230,N_23778);
or U24953 (N_24953,N_24347,N_24254);
xor U24954 (N_24954,N_23933,N_23986);
and U24955 (N_24955,N_24090,N_23772);
nor U24956 (N_24956,N_23923,N_24325);
and U24957 (N_24957,N_24139,N_24291);
or U24958 (N_24958,N_23901,N_23974);
nor U24959 (N_24959,N_23879,N_24015);
nand U24960 (N_24960,N_24155,N_23829);
nor U24961 (N_24961,N_24360,N_24214);
and U24962 (N_24962,N_24242,N_23977);
and U24963 (N_24963,N_24244,N_23971);
xor U24964 (N_24964,N_24126,N_23824);
nor U24965 (N_24965,N_24233,N_23962);
nand U24966 (N_24966,N_24004,N_23963);
or U24967 (N_24967,N_23806,N_24123);
nor U24968 (N_24968,N_24124,N_24201);
nand U24969 (N_24969,N_24231,N_23886);
nor U24970 (N_24970,N_24320,N_24041);
nand U24971 (N_24971,N_24068,N_23795);
and U24972 (N_24972,N_24049,N_23815);
nor U24973 (N_24973,N_23897,N_24081);
or U24974 (N_24974,N_23907,N_23976);
and U24975 (N_24975,N_24022,N_23923);
nand U24976 (N_24976,N_24061,N_23982);
or U24977 (N_24977,N_23775,N_24035);
xnor U24978 (N_24978,N_23998,N_24251);
nand U24979 (N_24979,N_24246,N_23979);
or U24980 (N_24980,N_24015,N_23811);
or U24981 (N_24981,N_24171,N_24123);
nand U24982 (N_24982,N_24070,N_24279);
xor U24983 (N_24983,N_24140,N_23999);
or U24984 (N_24984,N_23780,N_24249);
nor U24985 (N_24985,N_23885,N_23783);
xor U24986 (N_24986,N_23766,N_24026);
nor U24987 (N_24987,N_24322,N_23911);
nand U24988 (N_24988,N_24328,N_24370);
and U24989 (N_24989,N_24261,N_24023);
or U24990 (N_24990,N_23805,N_24314);
nand U24991 (N_24991,N_23755,N_24197);
nand U24992 (N_24992,N_24001,N_23943);
nor U24993 (N_24993,N_23813,N_23916);
nand U24994 (N_24994,N_24158,N_24024);
and U24995 (N_24995,N_23922,N_24197);
xnor U24996 (N_24996,N_24043,N_24337);
or U24997 (N_24997,N_24188,N_24192);
and U24998 (N_24998,N_23863,N_24034);
nand U24999 (N_24999,N_24230,N_24213);
xnor UO_0 (O_0,N_24793,N_24642);
or UO_1 (O_1,N_24712,N_24972);
nor UO_2 (O_2,N_24945,N_24704);
nand UO_3 (O_3,N_24784,N_24548);
nor UO_4 (O_4,N_24834,N_24524);
or UO_5 (O_5,N_24879,N_24990);
nor UO_6 (O_6,N_24933,N_24840);
or UO_7 (O_7,N_24585,N_24765);
nor UO_8 (O_8,N_24976,N_24719);
nor UO_9 (O_9,N_24641,N_24463);
xor UO_10 (O_10,N_24732,N_24671);
nand UO_11 (O_11,N_24583,N_24458);
nand UO_12 (O_12,N_24759,N_24674);
nor UO_13 (O_13,N_24640,N_24918);
nor UO_14 (O_14,N_24632,N_24492);
xnor UO_15 (O_15,N_24917,N_24561);
xor UO_16 (O_16,N_24591,N_24622);
nor UO_17 (O_17,N_24649,N_24549);
nand UO_18 (O_18,N_24695,N_24984);
and UO_19 (O_19,N_24812,N_24810);
nand UO_20 (O_20,N_24938,N_24876);
or UO_21 (O_21,N_24885,N_24489);
xnor UO_22 (O_22,N_24780,N_24958);
and UO_23 (O_23,N_24886,N_24459);
or UO_24 (O_24,N_24543,N_24658);
nand UO_25 (O_25,N_24638,N_24668);
or UO_26 (O_26,N_24673,N_24437);
xor UO_27 (O_27,N_24394,N_24635);
and UO_28 (O_28,N_24397,N_24752);
or UO_29 (O_29,N_24452,N_24686);
xor UO_30 (O_30,N_24837,N_24546);
or UO_31 (O_31,N_24479,N_24851);
or UO_32 (O_32,N_24656,N_24835);
or UO_33 (O_33,N_24628,N_24906);
and UO_34 (O_34,N_24403,N_24779);
nor UO_35 (O_35,N_24598,N_24989);
or UO_36 (O_36,N_24846,N_24946);
nand UO_37 (O_37,N_24692,N_24770);
nor UO_38 (O_38,N_24475,N_24790);
and UO_39 (O_39,N_24845,N_24565);
xor UO_40 (O_40,N_24451,N_24604);
nor UO_41 (O_41,N_24415,N_24574);
nand UO_42 (O_42,N_24731,N_24794);
nor UO_43 (O_43,N_24453,N_24472);
nand UO_44 (O_44,N_24968,N_24637);
xnor UO_45 (O_45,N_24468,N_24380);
and UO_46 (O_46,N_24538,N_24547);
nor UO_47 (O_47,N_24950,N_24690);
nor UO_48 (O_48,N_24934,N_24778);
nor UO_49 (O_49,N_24839,N_24416);
nor UO_50 (O_50,N_24956,N_24439);
xor UO_51 (O_51,N_24923,N_24418);
or UO_52 (O_52,N_24510,N_24662);
nor UO_53 (O_53,N_24469,N_24687);
or UO_54 (O_54,N_24572,N_24723);
nand UO_55 (O_55,N_24422,N_24995);
nor UO_56 (O_56,N_24672,N_24551);
or UO_57 (O_57,N_24733,N_24440);
nand UO_58 (O_58,N_24902,N_24665);
and UO_59 (O_59,N_24775,N_24527);
nand UO_60 (O_60,N_24856,N_24901);
xor UO_61 (O_61,N_24493,N_24587);
and UO_62 (O_62,N_24948,N_24761);
nor UO_63 (O_63,N_24427,N_24998);
nor UO_64 (O_64,N_24657,N_24722);
or UO_65 (O_65,N_24465,N_24831);
xor UO_66 (O_66,N_24434,N_24939);
nand UO_67 (O_67,N_24985,N_24911);
and UO_68 (O_68,N_24407,N_24661);
xor UO_69 (O_69,N_24785,N_24708);
nand UO_70 (O_70,N_24390,N_24398);
nor UO_71 (O_71,N_24825,N_24596);
nor UO_72 (O_72,N_24509,N_24426);
nor UO_73 (O_73,N_24554,N_24436);
nor UO_74 (O_74,N_24983,N_24786);
or UO_75 (O_75,N_24558,N_24400);
or UO_76 (O_76,N_24725,N_24660);
xnor UO_77 (O_77,N_24904,N_24599);
nand UO_78 (O_78,N_24385,N_24776);
nor UO_79 (O_79,N_24826,N_24696);
and UO_80 (O_80,N_24447,N_24644);
or UO_81 (O_81,N_24738,N_24593);
xor UO_82 (O_82,N_24727,N_24772);
and UO_83 (O_83,N_24544,N_24705);
nor UO_84 (O_84,N_24964,N_24613);
or UO_85 (O_85,N_24634,N_24470);
or UO_86 (O_86,N_24997,N_24444);
nor UO_87 (O_87,N_24913,N_24483);
nand UO_88 (O_88,N_24513,N_24858);
xnor UO_89 (O_89,N_24962,N_24566);
and UO_90 (O_90,N_24402,N_24949);
nand UO_91 (O_91,N_24907,N_24454);
nor UO_92 (O_92,N_24645,N_24535);
nand UO_93 (O_93,N_24651,N_24908);
or UO_94 (O_94,N_24860,N_24633);
and UO_95 (O_95,N_24833,N_24497);
and UO_96 (O_96,N_24920,N_24827);
nand UO_97 (O_97,N_24767,N_24707);
or UO_98 (O_98,N_24819,N_24944);
or UO_99 (O_99,N_24464,N_24979);
or UO_100 (O_100,N_24643,N_24986);
xnor UO_101 (O_101,N_24805,N_24391);
xnor UO_102 (O_102,N_24627,N_24910);
nor UO_103 (O_103,N_24814,N_24424);
xor UO_104 (O_104,N_24869,N_24621);
xnor UO_105 (O_105,N_24981,N_24515);
and UO_106 (O_106,N_24430,N_24396);
xor UO_107 (O_107,N_24867,N_24743);
nand UO_108 (O_108,N_24855,N_24376);
and UO_109 (O_109,N_24499,N_24615);
nand UO_110 (O_110,N_24682,N_24735);
nor UO_111 (O_111,N_24431,N_24714);
xnor UO_112 (O_112,N_24853,N_24569);
nor UO_113 (O_113,N_24862,N_24753);
nor UO_114 (O_114,N_24931,N_24954);
and UO_115 (O_115,N_24466,N_24824);
xor UO_116 (O_116,N_24620,N_24881);
nand UO_117 (O_117,N_24386,N_24517);
and UO_118 (O_118,N_24433,N_24650);
or UO_119 (O_119,N_24747,N_24573);
or UO_120 (O_120,N_24874,N_24963);
nor UO_121 (O_121,N_24655,N_24663);
nand UO_122 (O_122,N_24388,N_24844);
and UO_123 (O_123,N_24813,N_24530);
xnor UO_124 (O_124,N_24461,N_24909);
or UO_125 (O_125,N_24863,N_24539);
and UO_126 (O_126,N_24629,N_24670);
or UO_127 (O_127,N_24773,N_24857);
xnor UO_128 (O_128,N_24536,N_24919);
or UO_129 (O_129,N_24659,N_24542);
xnor UO_130 (O_130,N_24519,N_24736);
nand UO_131 (O_131,N_24562,N_24866);
xor UO_132 (O_132,N_24685,N_24699);
nor UO_133 (O_133,N_24847,N_24399);
xnor UO_134 (O_134,N_24854,N_24456);
or UO_135 (O_135,N_24446,N_24442);
nor UO_136 (O_136,N_24612,N_24880);
or UO_137 (O_137,N_24982,N_24496);
or UO_138 (O_138,N_24381,N_24383);
nor UO_139 (O_139,N_24594,N_24889);
and UO_140 (O_140,N_24926,N_24570);
nand UO_141 (O_141,N_24375,N_24413);
xnor UO_142 (O_142,N_24639,N_24597);
nand UO_143 (O_143,N_24841,N_24698);
xnor UO_144 (O_144,N_24905,N_24828);
nor UO_145 (O_145,N_24796,N_24520);
nor UO_146 (O_146,N_24387,N_24420);
or UO_147 (O_147,N_24914,N_24449);
and UO_148 (O_148,N_24611,N_24552);
or UO_149 (O_149,N_24467,N_24838);
nor UO_150 (O_150,N_24384,N_24936);
or UO_151 (O_151,N_24474,N_24807);
and UO_152 (O_152,N_24410,N_24405);
and UO_153 (O_153,N_24382,N_24648);
or UO_154 (O_154,N_24808,N_24471);
or UO_155 (O_155,N_24392,N_24584);
and UO_156 (O_156,N_24891,N_24850);
and UO_157 (O_157,N_24511,N_24969);
and UO_158 (O_158,N_24681,N_24533);
and UO_159 (O_159,N_24757,N_24559);
or UO_160 (O_160,N_24787,N_24664);
nand UO_161 (O_161,N_24927,N_24929);
and UO_162 (O_162,N_24429,N_24614);
or UO_163 (O_163,N_24892,N_24994);
nor UO_164 (O_164,N_24503,N_24978);
xnor UO_165 (O_165,N_24414,N_24528);
or UO_166 (O_166,N_24788,N_24495);
and UO_167 (O_167,N_24993,N_24378);
nand UO_168 (O_168,N_24618,N_24999);
nor UO_169 (O_169,N_24601,N_24996);
and UO_170 (O_170,N_24571,N_24744);
nand UO_171 (O_171,N_24521,N_24746);
or UO_172 (O_172,N_24768,N_24556);
nand UO_173 (O_173,N_24928,N_24646);
xnor UO_174 (O_174,N_24423,N_24771);
nand UO_175 (O_175,N_24729,N_24991);
xnor UO_176 (O_176,N_24488,N_24769);
and UO_177 (O_177,N_24783,N_24829);
or UO_178 (O_178,N_24518,N_24550);
nand UO_179 (O_179,N_24987,N_24797);
nand UO_180 (O_180,N_24677,N_24803);
or UO_181 (O_181,N_24848,N_24425);
nor UO_182 (O_182,N_24580,N_24925);
nand UO_183 (O_183,N_24581,N_24878);
xnor UO_184 (O_184,N_24462,N_24504);
nor UO_185 (O_185,N_24820,N_24966);
or UO_186 (O_186,N_24724,N_24610);
nor UO_187 (O_187,N_24882,N_24448);
and UO_188 (O_188,N_24899,N_24441);
nor UO_189 (O_189,N_24871,N_24417);
and UO_190 (O_190,N_24553,N_24404);
and UO_191 (O_191,N_24395,N_24915);
xnor UO_192 (O_192,N_24478,N_24792);
and UO_193 (O_193,N_24514,N_24700);
or UO_194 (O_194,N_24625,N_24576);
nor UO_195 (O_195,N_24870,N_24711);
nand UO_196 (O_196,N_24653,N_24718);
nand UO_197 (O_197,N_24516,N_24953);
xor UO_198 (O_198,N_24760,N_24975);
or UO_199 (O_199,N_24822,N_24623);
nor UO_200 (O_200,N_24602,N_24716);
or UO_201 (O_201,N_24888,N_24766);
xor UO_202 (O_202,N_24816,N_24408);
and UO_203 (O_203,N_24739,N_24795);
nand UO_204 (O_204,N_24943,N_24647);
xor UO_205 (O_205,N_24842,N_24455);
and UO_206 (O_206,N_24401,N_24774);
xor UO_207 (O_207,N_24849,N_24740);
nor UO_208 (O_208,N_24477,N_24764);
xor UO_209 (O_209,N_24560,N_24941);
nor UO_210 (O_210,N_24630,N_24500);
xor UO_211 (O_211,N_24890,N_24965);
or UO_212 (O_212,N_24756,N_24484);
or UO_213 (O_213,N_24896,N_24491);
and UO_214 (O_214,N_24809,N_24545);
nand UO_215 (O_215,N_24763,N_24877);
and UO_216 (O_216,N_24377,N_24616);
xor UO_217 (O_217,N_24873,N_24749);
or UO_218 (O_218,N_24603,N_24450);
and UO_219 (O_219,N_24804,N_24894);
and UO_220 (O_220,N_24710,N_24865);
xor UO_221 (O_221,N_24534,N_24412);
xor UO_222 (O_222,N_24830,N_24490);
xnor UO_223 (O_223,N_24525,N_24522);
nand UO_224 (O_224,N_24977,N_24460);
and UO_225 (O_225,N_24802,N_24947);
xnor UO_226 (O_226,N_24590,N_24435);
xnor UO_227 (O_227,N_24728,N_24563);
nand UO_228 (O_228,N_24540,N_24980);
and UO_229 (O_229,N_24678,N_24971);
or UO_230 (O_230,N_24811,N_24411);
and UO_231 (O_231,N_24884,N_24959);
or UO_232 (O_232,N_24409,N_24932);
nand UO_233 (O_233,N_24438,N_24501);
and UO_234 (O_234,N_24481,N_24592);
and UO_235 (O_235,N_24758,N_24702);
nor UO_236 (O_236,N_24389,N_24432);
xnor UO_237 (O_237,N_24726,N_24555);
xnor UO_238 (O_238,N_24589,N_24709);
and UO_239 (O_239,N_24961,N_24970);
xor UO_240 (O_240,N_24937,N_24688);
or UO_241 (O_241,N_24379,N_24798);
nand UO_242 (O_242,N_24421,N_24694);
xor UO_243 (O_243,N_24654,N_24823);
and UO_244 (O_244,N_24606,N_24443);
or UO_245 (O_245,N_24512,N_24703);
xor UO_246 (O_246,N_24745,N_24836);
nor UO_247 (O_247,N_24942,N_24737);
or UO_248 (O_248,N_24486,N_24912);
nor UO_249 (O_249,N_24557,N_24693);
nor UO_250 (O_250,N_24532,N_24666);
nor UO_251 (O_251,N_24806,N_24393);
and UO_252 (O_252,N_24895,N_24720);
nand UO_253 (O_253,N_24526,N_24935);
and UO_254 (O_254,N_24679,N_24575);
xnor UO_255 (O_255,N_24617,N_24609);
nand UO_256 (O_256,N_24930,N_24636);
and UO_257 (O_257,N_24782,N_24567);
xnor UO_258 (O_258,N_24588,N_24951);
xnor UO_259 (O_259,N_24974,N_24480);
and UO_260 (O_260,N_24741,N_24476);
or UO_261 (O_261,N_24706,N_24624);
xnor UO_262 (O_262,N_24817,N_24508);
nor UO_263 (O_263,N_24967,N_24777);
and UO_264 (O_264,N_24922,N_24898);
and UO_265 (O_265,N_24529,N_24755);
xnor UO_266 (O_266,N_24537,N_24541);
nand UO_267 (O_267,N_24903,N_24568);
nor UO_268 (O_268,N_24667,N_24843);
nor UO_269 (O_269,N_24924,N_24832);
or UO_270 (O_270,N_24697,N_24502);
nand UO_271 (O_271,N_24940,N_24762);
nand UO_272 (O_272,N_24482,N_24952);
xnor UO_273 (O_273,N_24713,N_24669);
and UO_274 (O_274,N_24631,N_24626);
and UO_275 (O_275,N_24900,N_24715);
nor UO_276 (O_276,N_24680,N_24586);
nor UO_277 (O_277,N_24498,N_24523);
and UO_278 (O_278,N_24485,N_24872);
nand UO_279 (O_279,N_24457,N_24577);
or UO_280 (O_280,N_24683,N_24801);
or UO_281 (O_281,N_24754,N_24689);
nor UO_282 (O_282,N_24608,N_24730);
and UO_283 (O_283,N_24992,N_24887);
xor UO_284 (O_284,N_24564,N_24957);
nand UO_285 (O_285,N_24691,N_24960);
and UO_286 (O_286,N_24619,N_24684);
nand UO_287 (O_287,N_24748,N_24701);
or UO_288 (O_288,N_24505,N_24428);
or UO_289 (O_289,N_24821,N_24955);
xor UO_290 (O_290,N_24406,N_24578);
nor UO_291 (O_291,N_24789,N_24487);
xor UO_292 (O_292,N_24419,N_24818);
nor UO_293 (O_293,N_24791,N_24815);
and UO_294 (O_294,N_24781,N_24897);
nand UO_295 (O_295,N_24652,N_24579);
and UO_296 (O_296,N_24506,N_24799);
xnor UO_297 (O_297,N_24676,N_24531);
or UO_298 (O_298,N_24605,N_24916);
and UO_299 (O_299,N_24721,N_24861);
xor UO_300 (O_300,N_24607,N_24859);
nand UO_301 (O_301,N_24717,N_24473);
nor UO_302 (O_302,N_24494,N_24675);
and UO_303 (O_303,N_24734,N_24582);
xor UO_304 (O_304,N_24921,N_24973);
nand UO_305 (O_305,N_24507,N_24750);
and UO_306 (O_306,N_24864,N_24875);
and UO_307 (O_307,N_24751,N_24988);
and UO_308 (O_308,N_24852,N_24800);
nor UO_309 (O_309,N_24595,N_24742);
or UO_310 (O_310,N_24893,N_24600);
or UO_311 (O_311,N_24445,N_24883);
xor UO_312 (O_312,N_24868,N_24590);
or UO_313 (O_313,N_24639,N_24414);
and UO_314 (O_314,N_24767,N_24713);
or UO_315 (O_315,N_24696,N_24662);
nor UO_316 (O_316,N_24455,N_24547);
nor UO_317 (O_317,N_24908,N_24815);
nand UO_318 (O_318,N_24550,N_24480);
nor UO_319 (O_319,N_24775,N_24391);
xor UO_320 (O_320,N_24652,N_24536);
nand UO_321 (O_321,N_24815,N_24720);
and UO_322 (O_322,N_24448,N_24862);
or UO_323 (O_323,N_24941,N_24995);
nand UO_324 (O_324,N_24984,N_24606);
nor UO_325 (O_325,N_24525,N_24751);
nor UO_326 (O_326,N_24407,N_24464);
and UO_327 (O_327,N_24742,N_24488);
xor UO_328 (O_328,N_24739,N_24642);
nor UO_329 (O_329,N_24642,N_24704);
xor UO_330 (O_330,N_24491,N_24833);
xnor UO_331 (O_331,N_24429,N_24737);
nand UO_332 (O_332,N_24854,N_24883);
xor UO_333 (O_333,N_24758,N_24989);
and UO_334 (O_334,N_24721,N_24712);
or UO_335 (O_335,N_24933,N_24409);
nor UO_336 (O_336,N_24460,N_24768);
xnor UO_337 (O_337,N_24939,N_24890);
xor UO_338 (O_338,N_24932,N_24977);
nor UO_339 (O_339,N_24436,N_24988);
xnor UO_340 (O_340,N_24573,N_24546);
nand UO_341 (O_341,N_24784,N_24604);
or UO_342 (O_342,N_24684,N_24732);
nand UO_343 (O_343,N_24854,N_24977);
nand UO_344 (O_344,N_24476,N_24623);
or UO_345 (O_345,N_24491,N_24530);
or UO_346 (O_346,N_24542,N_24691);
and UO_347 (O_347,N_24630,N_24976);
and UO_348 (O_348,N_24392,N_24833);
and UO_349 (O_349,N_24746,N_24783);
or UO_350 (O_350,N_24889,N_24502);
nor UO_351 (O_351,N_24886,N_24431);
xor UO_352 (O_352,N_24537,N_24747);
xnor UO_353 (O_353,N_24459,N_24487);
or UO_354 (O_354,N_24905,N_24462);
nand UO_355 (O_355,N_24884,N_24991);
and UO_356 (O_356,N_24864,N_24443);
nand UO_357 (O_357,N_24960,N_24817);
xnor UO_358 (O_358,N_24763,N_24432);
and UO_359 (O_359,N_24963,N_24480);
and UO_360 (O_360,N_24982,N_24471);
nor UO_361 (O_361,N_24809,N_24938);
nand UO_362 (O_362,N_24633,N_24705);
nor UO_363 (O_363,N_24461,N_24380);
and UO_364 (O_364,N_24994,N_24986);
or UO_365 (O_365,N_24824,N_24703);
nand UO_366 (O_366,N_24609,N_24508);
and UO_367 (O_367,N_24762,N_24892);
xnor UO_368 (O_368,N_24445,N_24876);
and UO_369 (O_369,N_24998,N_24755);
nand UO_370 (O_370,N_24442,N_24970);
nand UO_371 (O_371,N_24838,N_24503);
or UO_372 (O_372,N_24897,N_24613);
xnor UO_373 (O_373,N_24379,N_24696);
nand UO_374 (O_374,N_24926,N_24397);
xor UO_375 (O_375,N_24693,N_24790);
or UO_376 (O_376,N_24747,N_24791);
nand UO_377 (O_377,N_24763,N_24855);
and UO_378 (O_378,N_24696,N_24516);
and UO_379 (O_379,N_24708,N_24499);
xnor UO_380 (O_380,N_24520,N_24699);
nand UO_381 (O_381,N_24731,N_24658);
nand UO_382 (O_382,N_24458,N_24804);
nor UO_383 (O_383,N_24562,N_24999);
nand UO_384 (O_384,N_24968,N_24625);
and UO_385 (O_385,N_24489,N_24908);
nand UO_386 (O_386,N_24746,N_24446);
nor UO_387 (O_387,N_24467,N_24471);
xnor UO_388 (O_388,N_24411,N_24759);
or UO_389 (O_389,N_24673,N_24708);
and UO_390 (O_390,N_24681,N_24506);
or UO_391 (O_391,N_24401,N_24899);
or UO_392 (O_392,N_24883,N_24581);
nand UO_393 (O_393,N_24793,N_24584);
nor UO_394 (O_394,N_24565,N_24915);
nand UO_395 (O_395,N_24605,N_24423);
nor UO_396 (O_396,N_24635,N_24497);
nor UO_397 (O_397,N_24684,N_24637);
xor UO_398 (O_398,N_24528,N_24730);
xnor UO_399 (O_399,N_24809,N_24381);
nor UO_400 (O_400,N_24664,N_24848);
and UO_401 (O_401,N_24429,N_24559);
nor UO_402 (O_402,N_24694,N_24538);
nand UO_403 (O_403,N_24395,N_24743);
nor UO_404 (O_404,N_24973,N_24428);
nor UO_405 (O_405,N_24823,N_24893);
xnor UO_406 (O_406,N_24746,N_24678);
and UO_407 (O_407,N_24661,N_24394);
or UO_408 (O_408,N_24841,N_24495);
nor UO_409 (O_409,N_24893,N_24571);
nor UO_410 (O_410,N_24556,N_24969);
nor UO_411 (O_411,N_24937,N_24667);
xnor UO_412 (O_412,N_24765,N_24512);
nand UO_413 (O_413,N_24617,N_24720);
nor UO_414 (O_414,N_24484,N_24766);
nor UO_415 (O_415,N_24462,N_24722);
xor UO_416 (O_416,N_24396,N_24466);
nor UO_417 (O_417,N_24943,N_24985);
or UO_418 (O_418,N_24940,N_24463);
nor UO_419 (O_419,N_24465,N_24492);
nand UO_420 (O_420,N_24449,N_24770);
nand UO_421 (O_421,N_24823,N_24470);
xor UO_422 (O_422,N_24819,N_24560);
nor UO_423 (O_423,N_24848,N_24443);
nor UO_424 (O_424,N_24637,N_24612);
nor UO_425 (O_425,N_24471,N_24624);
nor UO_426 (O_426,N_24965,N_24941);
and UO_427 (O_427,N_24656,N_24990);
nor UO_428 (O_428,N_24527,N_24504);
nor UO_429 (O_429,N_24527,N_24689);
or UO_430 (O_430,N_24997,N_24850);
and UO_431 (O_431,N_24636,N_24837);
or UO_432 (O_432,N_24474,N_24790);
and UO_433 (O_433,N_24531,N_24669);
nand UO_434 (O_434,N_24656,N_24536);
xnor UO_435 (O_435,N_24674,N_24467);
xnor UO_436 (O_436,N_24570,N_24932);
nand UO_437 (O_437,N_24526,N_24393);
nor UO_438 (O_438,N_24859,N_24632);
or UO_439 (O_439,N_24906,N_24427);
or UO_440 (O_440,N_24549,N_24384);
nand UO_441 (O_441,N_24705,N_24990);
nor UO_442 (O_442,N_24718,N_24749);
or UO_443 (O_443,N_24796,N_24989);
and UO_444 (O_444,N_24849,N_24954);
or UO_445 (O_445,N_24718,N_24513);
nand UO_446 (O_446,N_24635,N_24676);
or UO_447 (O_447,N_24545,N_24464);
nor UO_448 (O_448,N_24469,N_24577);
xor UO_449 (O_449,N_24448,N_24886);
and UO_450 (O_450,N_24719,N_24860);
nor UO_451 (O_451,N_24565,N_24394);
and UO_452 (O_452,N_24492,N_24411);
and UO_453 (O_453,N_24857,N_24667);
or UO_454 (O_454,N_24406,N_24619);
or UO_455 (O_455,N_24483,N_24993);
nor UO_456 (O_456,N_24779,N_24610);
xor UO_457 (O_457,N_24871,N_24714);
and UO_458 (O_458,N_24978,N_24387);
and UO_459 (O_459,N_24909,N_24375);
nand UO_460 (O_460,N_24743,N_24906);
or UO_461 (O_461,N_24861,N_24617);
or UO_462 (O_462,N_24635,N_24892);
or UO_463 (O_463,N_24497,N_24829);
and UO_464 (O_464,N_24557,N_24774);
nor UO_465 (O_465,N_24849,N_24937);
and UO_466 (O_466,N_24714,N_24659);
nor UO_467 (O_467,N_24526,N_24478);
xnor UO_468 (O_468,N_24403,N_24467);
and UO_469 (O_469,N_24732,N_24579);
nand UO_470 (O_470,N_24519,N_24430);
nand UO_471 (O_471,N_24864,N_24893);
nor UO_472 (O_472,N_24613,N_24521);
xnor UO_473 (O_473,N_24596,N_24656);
and UO_474 (O_474,N_24956,N_24908);
or UO_475 (O_475,N_24636,N_24416);
or UO_476 (O_476,N_24832,N_24558);
nand UO_477 (O_477,N_24793,N_24497);
and UO_478 (O_478,N_24669,N_24390);
or UO_479 (O_479,N_24413,N_24819);
and UO_480 (O_480,N_24597,N_24503);
nor UO_481 (O_481,N_24756,N_24478);
nand UO_482 (O_482,N_24824,N_24952);
nand UO_483 (O_483,N_24400,N_24859);
nor UO_484 (O_484,N_24912,N_24502);
and UO_485 (O_485,N_24402,N_24722);
nand UO_486 (O_486,N_24855,N_24752);
nor UO_487 (O_487,N_24933,N_24760);
nor UO_488 (O_488,N_24594,N_24799);
and UO_489 (O_489,N_24652,N_24699);
xnor UO_490 (O_490,N_24482,N_24665);
or UO_491 (O_491,N_24486,N_24508);
xnor UO_492 (O_492,N_24442,N_24568);
or UO_493 (O_493,N_24951,N_24877);
and UO_494 (O_494,N_24541,N_24543);
or UO_495 (O_495,N_24996,N_24641);
and UO_496 (O_496,N_24457,N_24558);
xnor UO_497 (O_497,N_24576,N_24686);
xor UO_498 (O_498,N_24983,N_24559);
or UO_499 (O_499,N_24999,N_24673);
or UO_500 (O_500,N_24515,N_24837);
or UO_501 (O_501,N_24975,N_24431);
or UO_502 (O_502,N_24675,N_24498);
xnor UO_503 (O_503,N_24748,N_24793);
nor UO_504 (O_504,N_24771,N_24964);
and UO_505 (O_505,N_24719,N_24810);
nor UO_506 (O_506,N_24940,N_24722);
or UO_507 (O_507,N_24526,N_24961);
nor UO_508 (O_508,N_24638,N_24673);
or UO_509 (O_509,N_24763,N_24662);
and UO_510 (O_510,N_24935,N_24709);
xnor UO_511 (O_511,N_24968,N_24442);
and UO_512 (O_512,N_24978,N_24562);
nand UO_513 (O_513,N_24448,N_24529);
xnor UO_514 (O_514,N_24645,N_24723);
nor UO_515 (O_515,N_24747,N_24913);
and UO_516 (O_516,N_24379,N_24689);
and UO_517 (O_517,N_24516,N_24531);
xnor UO_518 (O_518,N_24690,N_24456);
and UO_519 (O_519,N_24706,N_24525);
nor UO_520 (O_520,N_24700,N_24990);
xnor UO_521 (O_521,N_24694,N_24387);
and UO_522 (O_522,N_24849,N_24500);
and UO_523 (O_523,N_24961,N_24559);
xnor UO_524 (O_524,N_24978,N_24438);
xnor UO_525 (O_525,N_24679,N_24776);
or UO_526 (O_526,N_24880,N_24475);
nand UO_527 (O_527,N_24558,N_24992);
xnor UO_528 (O_528,N_24507,N_24449);
or UO_529 (O_529,N_24424,N_24856);
nor UO_530 (O_530,N_24578,N_24789);
and UO_531 (O_531,N_24521,N_24381);
nand UO_532 (O_532,N_24872,N_24873);
nand UO_533 (O_533,N_24416,N_24873);
nand UO_534 (O_534,N_24578,N_24422);
and UO_535 (O_535,N_24953,N_24571);
and UO_536 (O_536,N_24890,N_24568);
nand UO_537 (O_537,N_24675,N_24394);
or UO_538 (O_538,N_24626,N_24478);
nand UO_539 (O_539,N_24871,N_24810);
and UO_540 (O_540,N_24425,N_24558);
xor UO_541 (O_541,N_24413,N_24776);
nor UO_542 (O_542,N_24496,N_24622);
xnor UO_543 (O_543,N_24459,N_24704);
xor UO_544 (O_544,N_24742,N_24795);
nor UO_545 (O_545,N_24551,N_24645);
xnor UO_546 (O_546,N_24542,N_24996);
xor UO_547 (O_547,N_24462,N_24684);
or UO_548 (O_548,N_24472,N_24992);
or UO_549 (O_549,N_24506,N_24755);
and UO_550 (O_550,N_24829,N_24742);
nor UO_551 (O_551,N_24710,N_24689);
nor UO_552 (O_552,N_24399,N_24637);
nor UO_553 (O_553,N_24933,N_24481);
and UO_554 (O_554,N_24764,N_24633);
xor UO_555 (O_555,N_24420,N_24917);
or UO_556 (O_556,N_24730,N_24808);
or UO_557 (O_557,N_24893,N_24974);
nand UO_558 (O_558,N_24688,N_24707);
and UO_559 (O_559,N_24886,N_24570);
nand UO_560 (O_560,N_24580,N_24715);
and UO_561 (O_561,N_24486,N_24706);
and UO_562 (O_562,N_24493,N_24392);
nand UO_563 (O_563,N_24725,N_24503);
nor UO_564 (O_564,N_24727,N_24613);
nor UO_565 (O_565,N_24962,N_24919);
and UO_566 (O_566,N_24626,N_24969);
xnor UO_567 (O_567,N_24917,N_24749);
or UO_568 (O_568,N_24545,N_24741);
or UO_569 (O_569,N_24627,N_24516);
nand UO_570 (O_570,N_24964,N_24710);
nand UO_571 (O_571,N_24636,N_24965);
and UO_572 (O_572,N_24817,N_24570);
xor UO_573 (O_573,N_24433,N_24935);
and UO_574 (O_574,N_24893,N_24859);
xnor UO_575 (O_575,N_24953,N_24468);
or UO_576 (O_576,N_24600,N_24965);
nand UO_577 (O_577,N_24514,N_24896);
or UO_578 (O_578,N_24421,N_24920);
xor UO_579 (O_579,N_24758,N_24849);
nand UO_580 (O_580,N_24920,N_24459);
nand UO_581 (O_581,N_24845,N_24519);
or UO_582 (O_582,N_24885,N_24423);
nor UO_583 (O_583,N_24729,N_24904);
or UO_584 (O_584,N_24659,N_24435);
nand UO_585 (O_585,N_24559,N_24432);
nand UO_586 (O_586,N_24982,N_24530);
and UO_587 (O_587,N_24535,N_24798);
nor UO_588 (O_588,N_24712,N_24636);
nand UO_589 (O_589,N_24522,N_24521);
xnor UO_590 (O_590,N_24762,N_24630);
or UO_591 (O_591,N_24767,N_24985);
nand UO_592 (O_592,N_24512,N_24419);
nand UO_593 (O_593,N_24930,N_24602);
xnor UO_594 (O_594,N_24440,N_24539);
nor UO_595 (O_595,N_24546,N_24876);
or UO_596 (O_596,N_24788,N_24653);
nor UO_597 (O_597,N_24597,N_24563);
or UO_598 (O_598,N_24709,N_24957);
and UO_599 (O_599,N_24755,N_24463);
nand UO_600 (O_600,N_24894,N_24870);
nand UO_601 (O_601,N_24786,N_24672);
nor UO_602 (O_602,N_24451,N_24517);
and UO_603 (O_603,N_24390,N_24818);
and UO_604 (O_604,N_24710,N_24796);
or UO_605 (O_605,N_24578,N_24493);
nor UO_606 (O_606,N_24930,N_24837);
and UO_607 (O_607,N_24512,N_24473);
xnor UO_608 (O_608,N_24758,N_24807);
and UO_609 (O_609,N_24929,N_24526);
xnor UO_610 (O_610,N_24802,N_24524);
nor UO_611 (O_611,N_24748,N_24810);
and UO_612 (O_612,N_24914,N_24974);
xnor UO_613 (O_613,N_24682,N_24788);
xor UO_614 (O_614,N_24962,N_24450);
nor UO_615 (O_615,N_24428,N_24720);
nor UO_616 (O_616,N_24999,N_24941);
and UO_617 (O_617,N_24678,N_24570);
nand UO_618 (O_618,N_24739,N_24947);
xor UO_619 (O_619,N_24977,N_24929);
or UO_620 (O_620,N_24874,N_24711);
xor UO_621 (O_621,N_24594,N_24686);
nor UO_622 (O_622,N_24939,N_24897);
and UO_623 (O_623,N_24969,N_24661);
xnor UO_624 (O_624,N_24382,N_24613);
nand UO_625 (O_625,N_24487,N_24881);
nor UO_626 (O_626,N_24964,N_24509);
xor UO_627 (O_627,N_24478,N_24496);
xor UO_628 (O_628,N_24938,N_24659);
nor UO_629 (O_629,N_24531,N_24845);
nand UO_630 (O_630,N_24595,N_24876);
xnor UO_631 (O_631,N_24946,N_24602);
and UO_632 (O_632,N_24820,N_24896);
nor UO_633 (O_633,N_24889,N_24942);
nand UO_634 (O_634,N_24566,N_24793);
and UO_635 (O_635,N_24387,N_24501);
nand UO_636 (O_636,N_24948,N_24404);
or UO_637 (O_637,N_24864,N_24813);
nand UO_638 (O_638,N_24438,N_24951);
or UO_639 (O_639,N_24396,N_24936);
or UO_640 (O_640,N_24697,N_24933);
and UO_641 (O_641,N_24831,N_24408);
or UO_642 (O_642,N_24513,N_24559);
or UO_643 (O_643,N_24385,N_24681);
nand UO_644 (O_644,N_24407,N_24845);
nand UO_645 (O_645,N_24686,N_24378);
nor UO_646 (O_646,N_24840,N_24520);
or UO_647 (O_647,N_24534,N_24819);
nor UO_648 (O_648,N_24605,N_24917);
and UO_649 (O_649,N_24914,N_24663);
nor UO_650 (O_650,N_24441,N_24544);
xnor UO_651 (O_651,N_24381,N_24522);
or UO_652 (O_652,N_24592,N_24400);
xnor UO_653 (O_653,N_24997,N_24680);
and UO_654 (O_654,N_24907,N_24553);
or UO_655 (O_655,N_24748,N_24770);
nand UO_656 (O_656,N_24454,N_24429);
or UO_657 (O_657,N_24758,N_24975);
nor UO_658 (O_658,N_24704,N_24868);
nand UO_659 (O_659,N_24918,N_24441);
and UO_660 (O_660,N_24916,N_24910);
xor UO_661 (O_661,N_24630,N_24736);
xnor UO_662 (O_662,N_24701,N_24823);
and UO_663 (O_663,N_24446,N_24685);
nor UO_664 (O_664,N_24766,N_24606);
xnor UO_665 (O_665,N_24449,N_24715);
xnor UO_666 (O_666,N_24855,N_24885);
and UO_667 (O_667,N_24742,N_24695);
or UO_668 (O_668,N_24560,N_24643);
and UO_669 (O_669,N_24913,N_24759);
nand UO_670 (O_670,N_24727,N_24523);
or UO_671 (O_671,N_24798,N_24894);
and UO_672 (O_672,N_24691,N_24759);
and UO_673 (O_673,N_24806,N_24708);
or UO_674 (O_674,N_24926,N_24450);
nor UO_675 (O_675,N_24846,N_24764);
or UO_676 (O_676,N_24959,N_24444);
nand UO_677 (O_677,N_24690,N_24911);
nand UO_678 (O_678,N_24709,N_24671);
or UO_679 (O_679,N_24776,N_24927);
and UO_680 (O_680,N_24726,N_24432);
nor UO_681 (O_681,N_24976,N_24457);
and UO_682 (O_682,N_24699,N_24789);
nand UO_683 (O_683,N_24927,N_24991);
or UO_684 (O_684,N_24803,N_24508);
nand UO_685 (O_685,N_24954,N_24981);
and UO_686 (O_686,N_24407,N_24382);
nand UO_687 (O_687,N_24794,N_24419);
nand UO_688 (O_688,N_24473,N_24998);
and UO_689 (O_689,N_24950,N_24590);
nand UO_690 (O_690,N_24663,N_24870);
or UO_691 (O_691,N_24403,N_24460);
or UO_692 (O_692,N_24955,N_24480);
nand UO_693 (O_693,N_24882,N_24985);
or UO_694 (O_694,N_24740,N_24386);
nor UO_695 (O_695,N_24522,N_24677);
and UO_696 (O_696,N_24397,N_24549);
xnor UO_697 (O_697,N_24449,N_24475);
nor UO_698 (O_698,N_24707,N_24775);
xor UO_699 (O_699,N_24846,N_24709);
nor UO_700 (O_700,N_24585,N_24778);
nand UO_701 (O_701,N_24607,N_24535);
or UO_702 (O_702,N_24565,N_24917);
nand UO_703 (O_703,N_24454,N_24874);
xor UO_704 (O_704,N_24862,N_24434);
and UO_705 (O_705,N_24394,N_24759);
xor UO_706 (O_706,N_24798,N_24636);
nor UO_707 (O_707,N_24926,N_24709);
xor UO_708 (O_708,N_24765,N_24624);
xor UO_709 (O_709,N_24810,N_24724);
or UO_710 (O_710,N_24700,N_24862);
xnor UO_711 (O_711,N_24945,N_24396);
xor UO_712 (O_712,N_24472,N_24657);
nand UO_713 (O_713,N_24603,N_24453);
nor UO_714 (O_714,N_24720,N_24400);
nor UO_715 (O_715,N_24971,N_24590);
nand UO_716 (O_716,N_24692,N_24667);
nor UO_717 (O_717,N_24464,N_24588);
or UO_718 (O_718,N_24401,N_24939);
or UO_719 (O_719,N_24642,N_24628);
xnor UO_720 (O_720,N_24698,N_24598);
xor UO_721 (O_721,N_24647,N_24458);
or UO_722 (O_722,N_24920,N_24778);
nand UO_723 (O_723,N_24602,N_24777);
xnor UO_724 (O_724,N_24497,N_24982);
nor UO_725 (O_725,N_24799,N_24619);
xnor UO_726 (O_726,N_24999,N_24755);
or UO_727 (O_727,N_24681,N_24703);
and UO_728 (O_728,N_24972,N_24831);
nand UO_729 (O_729,N_24826,N_24433);
xor UO_730 (O_730,N_24915,N_24782);
nor UO_731 (O_731,N_24883,N_24942);
or UO_732 (O_732,N_24454,N_24848);
nand UO_733 (O_733,N_24544,N_24609);
or UO_734 (O_734,N_24380,N_24592);
xor UO_735 (O_735,N_24461,N_24782);
nand UO_736 (O_736,N_24793,N_24437);
nand UO_737 (O_737,N_24845,N_24641);
xor UO_738 (O_738,N_24620,N_24392);
xor UO_739 (O_739,N_24867,N_24731);
xor UO_740 (O_740,N_24923,N_24385);
nor UO_741 (O_741,N_24797,N_24406);
xnor UO_742 (O_742,N_24784,N_24909);
nand UO_743 (O_743,N_24738,N_24851);
nand UO_744 (O_744,N_24712,N_24402);
nor UO_745 (O_745,N_24908,N_24831);
nor UO_746 (O_746,N_24385,N_24543);
nand UO_747 (O_747,N_24899,N_24914);
and UO_748 (O_748,N_24771,N_24565);
and UO_749 (O_749,N_24754,N_24533);
nand UO_750 (O_750,N_24708,N_24733);
nor UO_751 (O_751,N_24534,N_24963);
nand UO_752 (O_752,N_24766,N_24620);
nor UO_753 (O_753,N_24632,N_24569);
xor UO_754 (O_754,N_24507,N_24967);
or UO_755 (O_755,N_24695,N_24717);
xor UO_756 (O_756,N_24710,N_24390);
nor UO_757 (O_757,N_24816,N_24522);
nand UO_758 (O_758,N_24487,N_24810);
nor UO_759 (O_759,N_24883,N_24745);
nand UO_760 (O_760,N_24463,N_24763);
nor UO_761 (O_761,N_24499,N_24781);
nand UO_762 (O_762,N_24572,N_24979);
nor UO_763 (O_763,N_24583,N_24645);
xnor UO_764 (O_764,N_24584,N_24594);
nand UO_765 (O_765,N_24996,N_24376);
and UO_766 (O_766,N_24799,N_24401);
and UO_767 (O_767,N_24893,N_24900);
xor UO_768 (O_768,N_24601,N_24646);
nor UO_769 (O_769,N_24871,N_24657);
or UO_770 (O_770,N_24442,N_24762);
nand UO_771 (O_771,N_24410,N_24805);
xnor UO_772 (O_772,N_24916,N_24488);
and UO_773 (O_773,N_24823,N_24873);
nand UO_774 (O_774,N_24956,N_24573);
and UO_775 (O_775,N_24739,N_24387);
or UO_776 (O_776,N_24472,N_24950);
nand UO_777 (O_777,N_24451,N_24752);
nor UO_778 (O_778,N_24801,N_24513);
and UO_779 (O_779,N_24747,N_24945);
or UO_780 (O_780,N_24677,N_24862);
or UO_781 (O_781,N_24461,N_24931);
or UO_782 (O_782,N_24621,N_24724);
or UO_783 (O_783,N_24951,N_24733);
or UO_784 (O_784,N_24417,N_24478);
nand UO_785 (O_785,N_24649,N_24886);
nor UO_786 (O_786,N_24861,N_24816);
nor UO_787 (O_787,N_24574,N_24826);
nand UO_788 (O_788,N_24613,N_24994);
or UO_789 (O_789,N_24626,N_24601);
xor UO_790 (O_790,N_24876,N_24706);
and UO_791 (O_791,N_24739,N_24511);
and UO_792 (O_792,N_24940,N_24946);
or UO_793 (O_793,N_24798,N_24820);
nand UO_794 (O_794,N_24613,N_24643);
xnor UO_795 (O_795,N_24521,N_24858);
and UO_796 (O_796,N_24396,N_24906);
and UO_797 (O_797,N_24598,N_24904);
or UO_798 (O_798,N_24521,N_24899);
nand UO_799 (O_799,N_24455,N_24801);
and UO_800 (O_800,N_24419,N_24857);
xor UO_801 (O_801,N_24521,N_24657);
nor UO_802 (O_802,N_24416,N_24459);
nand UO_803 (O_803,N_24480,N_24909);
or UO_804 (O_804,N_24408,N_24506);
xnor UO_805 (O_805,N_24698,N_24892);
xor UO_806 (O_806,N_24516,N_24788);
nor UO_807 (O_807,N_24624,N_24762);
nand UO_808 (O_808,N_24445,N_24960);
xor UO_809 (O_809,N_24823,N_24983);
xnor UO_810 (O_810,N_24785,N_24946);
or UO_811 (O_811,N_24754,N_24960);
and UO_812 (O_812,N_24643,N_24595);
and UO_813 (O_813,N_24474,N_24511);
nand UO_814 (O_814,N_24551,N_24494);
xnor UO_815 (O_815,N_24735,N_24606);
or UO_816 (O_816,N_24978,N_24450);
nor UO_817 (O_817,N_24573,N_24951);
and UO_818 (O_818,N_24595,N_24787);
xor UO_819 (O_819,N_24523,N_24915);
nor UO_820 (O_820,N_24503,N_24681);
xnor UO_821 (O_821,N_24637,N_24994);
nor UO_822 (O_822,N_24646,N_24843);
nand UO_823 (O_823,N_24920,N_24465);
xnor UO_824 (O_824,N_24748,N_24427);
xnor UO_825 (O_825,N_24990,N_24800);
and UO_826 (O_826,N_24376,N_24811);
nor UO_827 (O_827,N_24732,N_24547);
xnor UO_828 (O_828,N_24775,N_24979);
nor UO_829 (O_829,N_24636,N_24792);
and UO_830 (O_830,N_24666,N_24873);
xnor UO_831 (O_831,N_24475,N_24524);
nor UO_832 (O_832,N_24851,N_24818);
nand UO_833 (O_833,N_24763,N_24495);
or UO_834 (O_834,N_24657,N_24709);
and UO_835 (O_835,N_24858,N_24664);
and UO_836 (O_836,N_24929,N_24436);
xor UO_837 (O_837,N_24513,N_24910);
and UO_838 (O_838,N_24627,N_24507);
xnor UO_839 (O_839,N_24773,N_24977);
nor UO_840 (O_840,N_24400,N_24942);
and UO_841 (O_841,N_24521,N_24797);
or UO_842 (O_842,N_24859,N_24997);
xor UO_843 (O_843,N_24563,N_24665);
nand UO_844 (O_844,N_24785,N_24448);
xnor UO_845 (O_845,N_24566,N_24455);
or UO_846 (O_846,N_24431,N_24662);
or UO_847 (O_847,N_24997,N_24880);
nand UO_848 (O_848,N_24786,N_24986);
or UO_849 (O_849,N_24952,N_24757);
or UO_850 (O_850,N_24397,N_24853);
nor UO_851 (O_851,N_24860,N_24451);
and UO_852 (O_852,N_24888,N_24463);
nor UO_853 (O_853,N_24660,N_24952);
or UO_854 (O_854,N_24740,N_24521);
nor UO_855 (O_855,N_24770,N_24870);
and UO_856 (O_856,N_24516,N_24496);
nor UO_857 (O_857,N_24735,N_24972);
xnor UO_858 (O_858,N_24402,N_24541);
nand UO_859 (O_859,N_24728,N_24710);
or UO_860 (O_860,N_24663,N_24487);
nand UO_861 (O_861,N_24485,N_24773);
and UO_862 (O_862,N_24606,N_24436);
and UO_863 (O_863,N_24521,N_24855);
xnor UO_864 (O_864,N_24667,N_24988);
nand UO_865 (O_865,N_24856,N_24829);
nor UO_866 (O_866,N_24577,N_24925);
or UO_867 (O_867,N_24579,N_24917);
nor UO_868 (O_868,N_24905,N_24488);
nand UO_869 (O_869,N_24493,N_24596);
nand UO_870 (O_870,N_24386,N_24591);
nor UO_871 (O_871,N_24984,N_24864);
and UO_872 (O_872,N_24716,N_24452);
nand UO_873 (O_873,N_24592,N_24932);
and UO_874 (O_874,N_24788,N_24542);
nor UO_875 (O_875,N_24510,N_24615);
or UO_876 (O_876,N_24636,N_24740);
nor UO_877 (O_877,N_24672,N_24658);
nand UO_878 (O_878,N_24987,N_24449);
and UO_879 (O_879,N_24554,N_24391);
and UO_880 (O_880,N_24493,N_24979);
or UO_881 (O_881,N_24608,N_24641);
nand UO_882 (O_882,N_24779,N_24525);
and UO_883 (O_883,N_24449,N_24620);
or UO_884 (O_884,N_24639,N_24991);
nand UO_885 (O_885,N_24664,N_24761);
xnor UO_886 (O_886,N_24690,N_24885);
nand UO_887 (O_887,N_24720,N_24497);
and UO_888 (O_888,N_24763,N_24955);
xnor UO_889 (O_889,N_24840,N_24458);
nor UO_890 (O_890,N_24996,N_24506);
or UO_891 (O_891,N_24537,N_24991);
nor UO_892 (O_892,N_24664,N_24960);
and UO_893 (O_893,N_24995,N_24914);
nor UO_894 (O_894,N_24835,N_24940);
xor UO_895 (O_895,N_24785,N_24928);
xnor UO_896 (O_896,N_24629,N_24767);
and UO_897 (O_897,N_24582,N_24426);
or UO_898 (O_898,N_24773,N_24685);
nor UO_899 (O_899,N_24401,N_24756);
nand UO_900 (O_900,N_24393,N_24392);
or UO_901 (O_901,N_24528,N_24644);
nand UO_902 (O_902,N_24674,N_24816);
and UO_903 (O_903,N_24846,N_24756);
or UO_904 (O_904,N_24851,N_24459);
and UO_905 (O_905,N_24604,N_24610);
xor UO_906 (O_906,N_24549,N_24659);
nand UO_907 (O_907,N_24509,N_24579);
and UO_908 (O_908,N_24800,N_24966);
nand UO_909 (O_909,N_24523,N_24591);
nand UO_910 (O_910,N_24384,N_24731);
nor UO_911 (O_911,N_24810,N_24948);
or UO_912 (O_912,N_24448,N_24535);
and UO_913 (O_913,N_24971,N_24784);
xnor UO_914 (O_914,N_24483,N_24400);
nand UO_915 (O_915,N_24824,N_24975);
xnor UO_916 (O_916,N_24674,N_24702);
xor UO_917 (O_917,N_24992,N_24583);
xnor UO_918 (O_918,N_24925,N_24764);
xnor UO_919 (O_919,N_24456,N_24473);
nand UO_920 (O_920,N_24586,N_24807);
or UO_921 (O_921,N_24676,N_24679);
xor UO_922 (O_922,N_24436,N_24447);
nand UO_923 (O_923,N_24630,N_24902);
or UO_924 (O_924,N_24586,N_24818);
nand UO_925 (O_925,N_24796,N_24492);
or UO_926 (O_926,N_24504,N_24468);
nor UO_927 (O_927,N_24693,N_24526);
xor UO_928 (O_928,N_24766,N_24829);
xnor UO_929 (O_929,N_24598,N_24981);
nand UO_930 (O_930,N_24581,N_24871);
and UO_931 (O_931,N_24796,N_24849);
or UO_932 (O_932,N_24544,N_24972);
and UO_933 (O_933,N_24773,N_24967);
nand UO_934 (O_934,N_24683,N_24612);
nor UO_935 (O_935,N_24457,N_24523);
and UO_936 (O_936,N_24473,N_24621);
nor UO_937 (O_937,N_24939,N_24508);
and UO_938 (O_938,N_24684,N_24529);
and UO_939 (O_939,N_24875,N_24422);
nor UO_940 (O_940,N_24377,N_24489);
xnor UO_941 (O_941,N_24806,N_24539);
nand UO_942 (O_942,N_24915,N_24824);
nor UO_943 (O_943,N_24705,N_24720);
and UO_944 (O_944,N_24508,N_24942);
xnor UO_945 (O_945,N_24766,N_24873);
and UO_946 (O_946,N_24927,N_24983);
nand UO_947 (O_947,N_24695,N_24991);
xor UO_948 (O_948,N_24404,N_24610);
or UO_949 (O_949,N_24795,N_24722);
nor UO_950 (O_950,N_24970,N_24547);
and UO_951 (O_951,N_24793,N_24708);
nor UO_952 (O_952,N_24565,N_24746);
and UO_953 (O_953,N_24832,N_24820);
and UO_954 (O_954,N_24957,N_24540);
xor UO_955 (O_955,N_24636,N_24453);
or UO_956 (O_956,N_24438,N_24606);
xor UO_957 (O_957,N_24903,N_24418);
nor UO_958 (O_958,N_24969,N_24809);
nand UO_959 (O_959,N_24964,N_24478);
nand UO_960 (O_960,N_24427,N_24853);
nor UO_961 (O_961,N_24616,N_24518);
and UO_962 (O_962,N_24868,N_24978);
and UO_963 (O_963,N_24570,N_24648);
or UO_964 (O_964,N_24508,N_24738);
xnor UO_965 (O_965,N_24526,N_24465);
and UO_966 (O_966,N_24778,N_24851);
nor UO_967 (O_967,N_24473,N_24458);
and UO_968 (O_968,N_24423,N_24647);
xor UO_969 (O_969,N_24954,N_24447);
xor UO_970 (O_970,N_24561,N_24388);
and UO_971 (O_971,N_24418,N_24527);
or UO_972 (O_972,N_24663,N_24784);
or UO_973 (O_973,N_24707,N_24608);
nor UO_974 (O_974,N_24447,N_24705);
nor UO_975 (O_975,N_24728,N_24813);
nor UO_976 (O_976,N_24384,N_24433);
and UO_977 (O_977,N_24790,N_24838);
nor UO_978 (O_978,N_24641,N_24544);
and UO_979 (O_979,N_24376,N_24992);
or UO_980 (O_980,N_24644,N_24470);
or UO_981 (O_981,N_24535,N_24950);
xor UO_982 (O_982,N_24619,N_24624);
nor UO_983 (O_983,N_24465,N_24607);
nor UO_984 (O_984,N_24538,N_24537);
nor UO_985 (O_985,N_24524,N_24432);
or UO_986 (O_986,N_24718,N_24845);
and UO_987 (O_987,N_24565,N_24932);
nor UO_988 (O_988,N_24466,N_24434);
nand UO_989 (O_989,N_24613,N_24785);
or UO_990 (O_990,N_24891,N_24479);
xnor UO_991 (O_991,N_24955,N_24481);
nand UO_992 (O_992,N_24888,N_24873);
and UO_993 (O_993,N_24660,N_24740);
or UO_994 (O_994,N_24679,N_24608);
nor UO_995 (O_995,N_24514,N_24892);
nor UO_996 (O_996,N_24460,N_24646);
nand UO_997 (O_997,N_24405,N_24757);
xor UO_998 (O_998,N_24561,N_24542);
and UO_999 (O_999,N_24713,N_24967);
xnor UO_1000 (O_1000,N_24673,N_24616);
or UO_1001 (O_1001,N_24891,N_24810);
and UO_1002 (O_1002,N_24827,N_24387);
xor UO_1003 (O_1003,N_24709,N_24386);
nor UO_1004 (O_1004,N_24408,N_24866);
xor UO_1005 (O_1005,N_24642,N_24812);
and UO_1006 (O_1006,N_24854,N_24783);
nor UO_1007 (O_1007,N_24577,N_24952);
and UO_1008 (O_1008,N_24402,N_24826);
xor UO_1009 (O_1009,N_24887,N_24834);
and UO_1010 (O_1010,N_24948,N_24415);
nor UO_1011 (O_1011,N_24697,N_24516);
and UO_1012 (O_1012,N_24982,N_24474);
or UO_1013 (O_1013,N_24498,N_24754);
or UO_1014 (O_1014,N_24828,N_24590);
or UO_1015 (O_1015,N_24802,N_24541);
and UO_1016 (O_1016,N_24867,N_24471);
nand UO_1017 (O_1017,N_24924,N_24420);
and UO_1018 (O_1018,N_24841,N_24902);
or UO_1019 (O_1019,N_24621,N_24958);
and UO_1020 (O_1020,N_24507,N_24384);
nand UO_1021 (O_1021,N_24715,N_24730);
nor UO_1022 (O_1022,N_24594,N_24652);
nand UO_1023 (O_1023,N_24522,N_24494);
and UO_1024 (O_1024,N_24757,N_24961);
or UO_1025 (O_1025,N_24592,N_24895);
nor UO_1026 (O_1026,N_24726,N_24385);
and UO_1027 (O_1027,N_24631,N_24618);
and UO_1028 (O_1028,N_24422,N_24435);
nand UO_1029 (O_1029,N_24576,N_24735);
and UO_1030 (O_1030,N_24703,N_24999);
nor UO_1031 (O_1031,N_24852,N_24511);
and UO_1032 (O_1032,N_24667,N_24900);
nand UO_1033 (O_1033,N_24574,N_24887);
nor UO_1034 (O_1034,N_24556,N_24750);
nand UO_1035 (O_1035,N_24921,N_24661);
or UO_1036 (O_1036,N_24439,N_24483);
and UO_1037 (O_1037,N_24661,N_24770);
or UO_1038 (O_1038,N_24959,N_24780);
or UO_1039 (O_1039,N_24705,N_24883);
nand UO_1040 (O_1040,N_24559,N_24870);
xnor UO_1041 (O_1041,N_24867,N_24894);
or UO_1042 (O_1042,N_24707,N_24542);
nor UO_1043 (O_1043,N_24488,N_24887);
and UO_1044 (O_1044,N_24854,N_24504);
xor UO_1045 (O_1045,N_24916,N_24456);
nand UO_1046 (O_1046,N_24562,N_24903);
nor UO_1047 (O_1047,N_24715,N_24853);
nor UO_1048 (O_1048,N_24532,N_24855);
and UO_1049 (O_1049,N_24879,N_24460);
and UO_1050 (O_1050,N_24911,N_24831);
nand UO_1051 (O_1051,N_24822,N_24809);
nor UO_1052 (O_1052,N_24705,N_24434);
and UO_1053 (O_1053,N_24726,N_24830);
or UO_1054 (O_1054,N_24727,N_24741);
xor UO_1055 (O_1055,N_24891,N_24971);
xor UO_1056 (O_1056,N_24397,N_24993);
nor UO_1057 (O_1057,N_24461,N_24483);
nor UO_1058 (O_1058,N_24943,N_24846);
xor UO_1059 (O_1059,N_24920,N_24979);
xnor UO_1060 (O_1060,N_24869,N_24701);
nor UO_1061 (O_1061,N_24467,N_24536);
nand UO_1062 (O_1062,N_24516,N_24486);
and UO_1063 (O_1063,N_24633,N_24596);
xor UO_1064 (O_1064,N_24798,N_24540);
nand UO_1065 (O_1065,N_24426,N_24611);
and UO_1066 (O_1066,N_24985,N_24595);
or UO_1067 (O_1067,N_24511,N_24454);
xnor UO_1068 (O_1068,N_24826,N_24956);
nand UO_1069 (O_1069,N_24780,N_24611);
xnor UO_1070 (O_1070,N_24577,N_24792);
nor UO_1071 (O_1071,N_24527,N_24949);
nand UO_1072 (O_1072,N_24742,N_24407);
and UO_1073 (O_1073,N_24521,N_24394);
nor UO_1074 (O_1074,N_24623,N_24711);
nor UO_1075 (O_1075,N_24533,N_24744);
nand UO_1076 (O_1076,N_24417,N_24431);
and UO_1077 (O_1077,N_24443,N_24914);
nor UO_1078 (O_1078,N_24757,N_24595);
and UO_1079 (O_1079,N_24736,N_24867);
nor UO_1080 (O_1080,N_24995,N_24510);
nor UO_1081 (O_1081,N_24964,N_24890);
and UO_1082 (O_1082,N_24405,N_24632);
nand UO_1083 (O_1083,N_24747,N_24578);
nor UO_1084 (O_1084,N_24546,N_24933);
xor UO_1085 (O_1085,N_24504,N_24634);
xnor UO_1086 (O_1086,N_24676,N_24590);
or UO_1087 (O_1087,N_24519,N_24380);
and UO_1088 (O_1088,N_24815,N_24541);
or UO_1089 (O_1089,N_24706,N_24461);
or UO_1090 (O_1090,N_24890,N_24725);
nor UO_1091 (O_1091,N_24941,N_24899);
and UO_1092 (O_1092,N_24785,N_24501);
xnor UO_1093 (O_1093,N_24586,N_24771);
nand UO_1094 (O_1094,N_24674,N_24739);
nand UO_1095 (O_1095,N_24978,N_24649);
nor UO_1096 (O_1096,N_24415,N_24514);
nand UO_1097 (O_1097,N_24740,N_24694);
or UO_1098 (O_1098,N_24428,N_24403);
and UO_1099 (O_1099,N_24728,N_24694);
nor UO_1100 (O_1100,N_24675,N_24889);
xor UO_1101 (O_1101,N_24394,N_24652);
nor UO_1102 (O_1102,N_24757,N_24603);
xor UO_1103 (O_1103,N_24966,N_24406);
nand UO_1104 (O_1104,N_24638,N_24565);
xor UO_1105 (O_1105,N_24974,N_24703);
or UO_1106 (O_1106,N_24724,N_24998);
nor UO_1107 (O_1107,N_24736,N_24434);
xor UO_1108 (O_1108,N_24397,N_24705);
or UO_1109 (O_1109,N_24803,N_24802);
and UO_1110 (O_1110,N_24906,N_24687);
xnor UO_1111 (O_1111,N_24669,N_24878);
and UO_1112 (O_1112,N_24706,N_24652);
nand UO_1113 (O_1113,N_24640,N_24425);
nand UO_1114 (O_1114,N_24802,N_24613);
nor UO_1115 (O_1115,N_24408,N_24660);
and UO_1116 (O_1116,N_24967,N_24931);
and UO_1117 (O_1117,N_24553,N_24801);
or UO_1118 (O_1118,N_24863,N_24463);
xnor UO_1119 (O_1119,N_24821,N_24778);
xor UO_1120 (O_1120,N_24664,N_24626);
xnor UO_1121 (O_1121,N_24777,N_24856);
and UO_1122 (O_1122,N_24560,N_24800);
or UO_1123 (O_1123,N_24392,N_24566);
or UO_1124 (O_1124,N_24956,N_24636);
nor UO_1125 (O_1125,N_24768,N_24689);
or UO_1126 (O_1126,N_24494,N_24582);
or UO_1127 (O_1127,N_24713,N_24958);
nor UO_1128 (O_1128,N_24819,N_24739);
nand UO_1129 (O_1129,N_24509,N_24472);
and UO_1130 (O_1130,N_24892,N_24724);
and UO_1131 (O_1131,N_24463,N_24800);
xor UO_1132 (O_1132,N_24554,N_24461);
or UO_1133 (O_1133,N_24486,N_24836);
nand UO_1134 (O_1134,N_24854,N_24727);
or UO_1135 (O_1135,N_24876,N_24919);
nand UO_1136 (O_1136,N_24810,N_24896);
nor UO_1137 (O_1137,N_24657,N_24400);
xor UO_1138 (O_1138,N_24618,N_24854);
nand UO_1139 (O_1139,N_24913,N_24499);
or UO_1140 (O_1140,N_24391,N_24974);
nor UO_1141 (O_1141,N_24701,N_24433);
and UO_1142 (O_1142,N_24751,N_24876);
nand UO_1143 (O_1143,N_24494,N_24401);
nor UO_1144 (O_1144,N_24729,N_24377);
or UO_1145 (O_1145,N_24595,N_24488);
nor UO_1146 (O_1146,N_24587,N_24998);
nor UO_1147 (O_1147,N_24662,N_24551);
nor UO_1148 (O_1148,N_24560,N_24435);
xnor UO_1149 (O_1149,N_24649,N_24652);
nor UO_1150 (O_1150,N_24960,N_24877);
xor UO_1151 (O_1151,N_24670,N_24803);
and UO_1152 (O_1152,N_24629,N_24736);
nor UO_1153 (O_1153,N_24804,N_24407);
nand UO_1154 (O_1154,N_24701,N_24538);
and UO_1155 (O_1155,N_24522,N_24627);
and UO_1156 (O_1156,N_24891,N_24474);
nand UO_1157 (O_1157,N_24625,N_24503);
nand UO_1158 (O_1158,N_24598,N_24422);
nand UO_1159 (O_1159,N_24626,N_24438);
nor UO_1160 (O_1160,N_24631,N_24788);
or UO_1161 (O_1161,N_24966,N_24934);
or UO_1162 (O_1162,N_24711,N_24804);
and UO_1163 (O_1163,N_24738,N_24441);
or UO_1164 (O_1164,N_24824,N_24676);
or UO_1165 (O_1165,N_24772,N_24589);
xnor UO_1166 (O_1166,N_24655,N_24639);
xor UO_1167 (O_1167,N_24522,N_24622);
nand UO_1168 (O_1168,N_24774,N_24993);
nand UO_1169 (O_1169,N_24460,N_24796);
and UO_1170 (O_1170,N_24590,N_24752);
or UO_1171 (O_1171,N_24621,N_24481);
and UO_1172 (O_1172,N_24899,N_24603);
and UO_1173 (O_1173,N_24378,N_24748);
nand UO_1174 (O_1174,N_24406,N_24826);
nand UO_1175 (O_1175,N_24681,N_24465);
and UO_1176 (O_1176,N_24907,N_24922);
nor UO_1177 (O_1177,N_24662,N_24863);
or UO_1178 (O_1178,N_24556,N_24472);
and UO_1179 (O_1179,N_24967,N_24971);
xnor UO_1180 (O_1180,N_24971,N_24822);
nand UO_1181 (O_1181,N_24454,N_24696);
and UO_1182 (O_1182,N_24860,N_24716);
xor UO_1183 (O_1183,N_24647,N_24644);
xnor UO_1184 (O_1184,N_24636,N_24623);
xor UO_1185 (O_1185,N_24523,N_24817);
nand UO_1186 (O_1186,N_24434,N_24591);
nand UO_1187 (O_1187,N_24753,N_24382);
xor UO_1188 (O_1188,N_24586,N_24983);
nor UO_1189 (O_1189,N_24602,N_24804);
xnor UO_1190 (O_1190,N_24486,N_24937);
and UO_1191 (O_1191,N_24807,N_24711);
or UO_1192 (O_1192,N_24426,N_24749);
and UO_1193 (O_1193,N_24607,N_24454);
or UO_1194 (O_1194,N_24886,N_24799);
nand UO_1195 (O_1195,N_24694,N_24490);
or UO_1196 (O_1196,N_24945,N_24609);
or UO_1197 (O_1197,N_24544,N_24963);
nand UO_1198 (O_1198,N_24410,N_24787);
xnor UO_1199 (O_1199,N_24708,N_24606);
nand UO_1200 (O_1200,N_24699,N_24696);
nand UO_1201 (O_1201,N_24629,N_24486);
and UO_1202 (O_1202,N_24501,N_24689);
and UO_1203 (O_1203,N_24900,N_24721);
or UO_1204 (O_1204,N_24432,N_24418);
nor UO_1205 (O_1205,N_24522,N_24868);
or UO_1206 (O_1206,N_24387,N_24392);
and UO_1207 (O_1207,N_24444,N_24858);
and UO_1208 (O_1208,N_24886,N_24837);
nand UO_1209 (O_1209,N_24759,N_24769);
nand UO_1210 (O_1210,N_24951,N_24858);
and UO_1211 (O_1211,N_24731,N_24962);
xor UO_1212 (O_1212,N_24593,N_24430);
or UO_1213 (O_1213,N_24583,N_24703);
and UO_1214 (O_1214,N_24709,N_24856);
nor UO_1215 (O_1215,N_24464,N_24656);
nand UO_1216 (O_1216,N_24830,N_24671);
nand UO_1217 (O_1217,N_24775,N_24748);
nand UO_1218 (O_1218,N_24903,N_24500);
and UO_1219 (O_1219,N_24519,N_24437);
xnor UO_1220 (O_1220,N_24802,N_24855);
and UO_1221 (O_1221,N_24583,N_24434);
nand UO_1222 (O_1222,N_24537,N_24838);
nor UO_1223 (O_1223,N_24845,N_24724);
xor UO_1224 (O_1224,N_24521,N_24722);
or UO_1225 (O_1225,N_24849,N_24663);
nand UO_1226 (O_1226,N_24829,N_24826);
and UO_1227 (O_1227,N_24904,N_24939);
and UO_1228 (O_1228,N_24699,N_24776);
nand UO_1229 (O_1229,N_24568,N_24849);
or UO_1230 (O_1230,N_24389,N_24513);
nand UO_1231 (O_1231,N_24776,N_24513);
nor UO_1232 (O_1232,N_24478,N_24716);
and UO_1233 (O_1233,N_24418,N_24608);
or UO_1234 (O_1234,N_24391,N_24570);
or UO_1235 (O_1235,N_24933,N_24631);
or UO_1236 (O_1236,N_24978,N_24763);
xnor UO_1237 (O_1237,N_24690,N_24405);
xor UO_1238 (O_1238,N_24640,N_24910);
and UO_1239 (O_1239,N_24793,N_24677);
xnor UO_1240 (O_1240,N_24470,N_24910);
nor UO_1241 (O_1241,N_24948,N_24654);
or UO_1242 (O_1242,N_24893,N_24657);
xnor UO_1243 (O_1243,N_24817,N_24566);
xor UO_1244 (O_1244,N_24656,N_24644);
nor UO_1245 (O_1245,N_24607,N_24513);
and UO_1246 (O_1246,N_24457,N_24623);
nor UO_1247 (O_1247,N_24733,N_24417);
nand UO_1248 (O_1248,N_24384,N_24686);
and UO_1249 (O_1249,N_24943,N_24996);
xor UO_1250 (O_1250,N_24955,N_24807);
or UO_1251 (O_1251,N_24457,N_24676);
nor UO_1252 (O_1252,N_24376,N_24423);
nand UO_1253 (O_1253,N_24801,N_24918);
nor UO_1254 (O_1254,N_24527,N_24687);
nand UO_1255 (O_1255,N_24970,N_24546);
nor UO_1256 (O_1256,N_24522,N_24440);
nor UO_1257 (O_1257,N_24490,N_24603);
nor UO_1258 (O_1258,N_24397,N_24596);
nor UO_1259 (O_1259,N_24837,N_24947);
xnor UO_1260 (O_1260,N_24618,N_24794);
nand UO_1261 (O_1261,N_24869,N_24879);
xor UO_1262 (O_1262,N_24513,N_24588);
or UO_1263 (O_1263,N_24908,N_24410);
xnor UO_1264 (O_1264,N_24484,N_24792);
nor UO_1265 (O_1265,N_24988,N_24478);
nor UO_1266 (O_1266,N_24458,N_24580);
or UO_1267 (O_1267,N_24789,N_24444);
xor UO_1268 (O_1268,N_24561,N_24379);
nand UO_1269 (O_1269,N_24784,N_24644);
and UO_1270 (O_1270,N_24882,N_24956);
xor UO_1271 (O_1271,N_24762,N_24873);
nand UO_1272 (O_1272,N_24924,N_24407);
or UO_1273 (O_1273,N_24974,N_24547);
and UO_1274 (O_1274,N_24546,N_24959);
nor UO_1275 (O_1275,N_24905,N_24447);
and UO_1276 (O_1276,N_24701,N_24416);
or UO_1277 (O_1277,N_24673,N_24441);
or UO_1278 (O_1278,N_24840,N_24756);
xnor UO_1279 (O_1279,N_24395,N_24732);
nand UO_1280 (O_1280,N_24450,N_24910);
nor UO_1281 (O_1281,N_24711,N_24529);
xor UO_1282 (O_1282,N_24453,N_24494);
nand UO_1283 (O_1283,N_24587,N_24603);
nor UO_1284 (O_1284,N_24757,N_24896);
and UO_1285 (O_1285,N_24489,N_24775);
xnor UO_1286 (O_1286,N_24633,N_24660);
xnor UO_1287 (O_1287,N_24525,N_24982);
nand UO_1288 (O_1288,N_24780,N_24567);
nor UO_1289 (O_1289,N_24702,N_24648);
nor UO_1290 (O_1290,N_24486,N_24942);
nand UO_1291 (O_1291,N_24706,N_24421);
nor UO_1292 (O_1292,N_24453,N_24971);
xor UO_1293 (O_1293,N_24856,N_24645);
nor UO_1294 (O_1294,N_24447,N_24642);
and UO_1295 (O_1295,N_24922,N_24657);
nor UO_1296 (O_1296,N_24886,N_24382);
nor UO_1297 (O_1297,N_24909,N_24904);
nor UO_1298 (O_1298,N_24656,N_24978);
or UO_1299 (O_1299,N_24541,N_24668);
or UO_1300 (O_1300,N_24675,N_24697);
nand UO_1301 (O_1301,N_24375,N_24760);
and UO_1302 (O_1302,N_24638,N_24661);
and UO_1303 (O_1303,N_24987,N_24943);
xor UO_1304 (O_1304,N_24822,N_24951);
and UO_1305 (O_1305,N_24736,N_24460);
nand UO_1306 (O_1306,N_24825,N_24495);
or UO_1307 (O_1307,N_24969,N_24714);
xnor UO_1308 (O_1308,N_24758,N_24710);
nor UO_1309 (O_1309,N_24743,N_24712);
xnor UO_1310 (O_1310,N_24865,N_24428);
nand UO_1311 (O_1311,N_24766,N_24608);
nand UO_1312 (O_1312,N_24680,N_24725);
or UO_1313 (O_1313,N_24861,N_24983);
or UO_1314 (O_1314,N_24606,N_24913);
xnor UO_1315 (O_1315,N_24886,N_24379);
xnor UO_1316 (O_1316,N_24411,N_24524);
xnor UO_1317 (O_1317,N_24818,N_24670);
nand UO_1318 (O_1318,N_24611,N_24857);
or UO_1319 (O_1319,N_24995,N_24936);
nor UO_1320 (O_1320,N_24573,N_24721);
nor UO_1321 (O_1321,N_24495,N_24886);
xnor UO_1322 (O_1322,N_24721,N_24834);
or UO_1323 (O_1323,N_24852,N_24433);
or UO_1324 (O_1324,N_24826,N_24697);
and UO_1325 (O_1325,N_24842,N_24865);
nor UO_1326 (O_1326,N_24507,N_24665);
xnor UO_1327 (O_1327,N_24552,N_24862);
or UO_1328 (O_1328,N_24993,N_24525);
or UO_1329 (O_1329,N_24595,N_24609);
xnor UO_1330 (O_1330,N_24672,N_24663);
xor UO_1331 (O_1331,N_24780,N_24636);
or UO_1332 (O_1332,N_24926,N_24679);
nor UO_1333 (O_1333,N_24623,N_24406);
and UO_1334 (O_1334,N_24822,N_24442);
and UO_1335 (O_1335,N_24497,N_24430);
xor UO_1336 (O_1336,N_24582,N_24705);
or UO_1337 (O_1337,N_24442,N_24982);
xnor UO_1338 (O_1338,N_24717,N_24934);
and UO_1339 (O_1339,N_24840,N_24738);
xor UO_1340 (O_1340,N_24547,N_24689);
nor UO_1341 (O_1341,N_24568,N_24392);
and UO_1342 (O_1342,N_24826,N_24644);
xnor UO_1343 (O_1343,N_24603,N_24547);
xnor UO_1344 (O_1344,N_24477,N_24728);
xnor UO_1345 (O_1345,N_24822,N_24772);
xnor UO_1346 (O_1346,N_24765,N_24966);
nor UO_1347 (O_1347,N_24909,N_24811);
nand UO_1348 (O_1348,N_24991,N_24498);
and UO_1349 (O_1349,N_24736,N_24976);
nor UO_1350 (O_1350,N_24920,N_24528);
and UO_1351 (O_1351,N_24412,N_24719);
and UO_1352 (O_1352,N_24536,N_24449);
and UO_1353 (O_1353,N_24422,N_24869);
and UO_1354 (O_1354,N_24893,N_24512);
nor UO_1355 (O_1355,N_24818,N_24455);
and UO_1356 (O_1356,N_24378,N_24741);
and UO_1357 (O_1357,N_24995,N_24506);
and UO_1358 (O_1358,N_24451,N_24483);
nand UO_1359 (O_1359,N_24853,N_24800);
and UO_1360 (O_1360,N_24720,N_24527);
or UO_1361 (O_1361,N_24396,N_24990);
and UO_1362 (O_1362,N_24495,N_24688);
or UO_1363 (O_1363,N_24990,N_24821);
nor UO_1364 (O_1364,N_24449,N_24701);
xnor UO_1365 (O_1365,N_24566,N_24693);
xnor UO_1366 (O_1366,N_24396,N_24773);
or UO_1367 (O_1367,N_24594,N_24375);
and UO_1368 (O_1368,N_24708,N_24676);
xor UO_1369 (O_1369,N_24709,N_24653);
or UO_1370 (O_1370,N_24692,N_24624);
and UO_1371 (O_1371,N_24751,N_24668);
or UO_1372 (O_1372,N_24452,N_24739);
nand UO_1373 (O_1373,N_24882,N_24430);
xor UO_1374 (O_1374,N_24702,N_24972);
nor UO_1375 (O_1375,N_24543,N_24455);
and UO_1376 (O_1376,N_24441,N_24893);
nand UO_1377 (O_1377,N_24686,N_24922);
xnor UO_1378 (O_1378,N_24844,N_24803);
and UO_1379 (O_1379,N_24766,N_24551);
and UO_1380 (O_1380,N_24949,N_24902);
xnor UO_1381 (O_1381,N_24516,N_24918);
nor UO_1382 (O_1382,N_24466,N_24914);
nor UO_1383 (O_1383,N_24381,N_24586);
xnor UO_1384 (O_1384,N_24643,N_24774);
nor UO_1385 (O_1385,N_24670,N_24591);
nand UO_1386 (O_1386,N_24428,N_24974);
nand UO_1387 (O_1387,N_24563,N_24466);
nand UO_1388 (O_1388,N_24488,N_24519);
and UO_1389 (O_1389,N_24607,N_24660);
and UO_1390 (O_1390,N_24598,N_24605);
nor UO_1391 (O_1391,N_24861,N_24453);
and UO_1392 (O_1392,N_24464,N_24632);
nor UO_1393 (O_1393,N_24483,N_24620);
and UO_1394 (O_1394,N_24891,N_24699);
xor UO_1395 (O_1395,N_24977,N_24963);
and UO_1396 (O_1396,N_24834,N_24788);
or UO_1397 (O_1397,N_24955,N_24643);
and UO_1398 (O_1398,N_24844,N_24832);
nand UO_1399 (O_1399,N_24641,N_24970);
and UO_1400 (O_1400,N_24472,N_24809);
or UO_1401 (O_1401,N_24716,N_24399);
nor UO_1402 (O_1402,N_24713,N_24606);
or UO_1403 (O_1403,N_24454,N_24734);
or UO_1404 (O_1404,N_24399,N_24754);
or UO_1405 (O_1405,N_24429,N_24717);
nand UO_1406 (O_1406,N_24412,N_24913);
or UO_1407 (O_1407,N_24885,N_24464);
nor UO_1408 (O_1408,N_24572,N_24981);
and UO_1409 (O_1409,N_24399,N_24896);
nor UO_1410 (O_1410,N_24967,N_24457);
nand UO_1411 (O_1411,N_24809,N_24957);
nor UO_1412 (O_1412,N_24665,N_24977);
or UO_1413 (O_1413,N_24512,N_24434);
and UO_1414 (O_1414,N_24883,N_24537);
nor UO_1415 (O_1415,N_24598,N_24774);
or UO_1416 (O_1416,N_24584,N_24419);
nand UO_1417 (O_1417,N_24399,N_24490);
and UO_1418 (O_1418,N_24789,N_24792);
and UO_1419 (O_1419,N_24689,N_24717);
xor UO_1420 (O_1420,N_24996,N_24652);
xnor UO_1421 (O_1421,N_24854,N_24962);
and UO_1422 (O_1422,N_24880,N_24549);
nor UO_1423 (O_1423,N_24888,N_24429);
and UO_1424 (O_1424,N_24807,N_24801);
nand UO_1425 (O_1425,N_24751,N_24871);
nor UO_1426 (O_1426,N_24878,N_24671);
xnor UO_1427 (O_1427,N_24957,N_24614);
xor UO_1428 (O_1428,N_24553,N_24562);
or UO_1429 (O_1429,N_24957,N_24906);
nor UO_1430 (O_1430,N_24553,N_24450);
nor UO_1431 (O_1431,N_24642,N_24887);
nor UO_1432 (O_1432,N_24528,N_24759);
nand UO_1433 (O_1433,N_24684,N_24905);
nor UO_1434 (O_1434,N_24615,N_24727);
xor UO_1435 (O_1435,N_24660,N_24895);
and UO_1436 (O_1436,N_24855,N_24601);
nand UO_1437 (O_1437,N_24776,N_24649);
nand UO_1438 (O_1438,N_24403,N_24387);
or UO_1439 (O_1439,N_24890,N_24855);
nand UO_1440 (O_1440,N_24570,N_24484);
and UO_1441 (O_1441,N_24550,N_24932);
or UO_1442 (O_1442,N_24593,N_24468);
nand UO_1443 (O_1443,N_24728,N_24390);
nand UO_1444 (O_1444,N_24817,N_24735);
nand UO_1445 (O_1445,N_24972,N_24533);
xnor UO_1446 (O_1446,N_24789,N_24548);
and UO_1447 (O_1447,N_24389,N_24694);
xnor UO_1448 (O_1448,N_24840,N_24526);
xnor UO_1449 (O_1449,N_24876,N_24536);
nor UO_1450 (O_1450,N_24664,N_24554);
xnor UO_1451 (O_1451,N_24754,N_24447);
nor UO_1452 (O_1452,N_24473,N_24746);
and UO_1453 (O_1453,N_24837,N_24860);
xor UO_1454 (O_1454,N_24908,N_24747);
and UO_1455 (O_1455,N_24477,N_24814);
nand UO_1456 (O_1456,N_24382,N_24765);
nand UO_1457 (O_1457,N_24384,N_24520);
xor UO_1458 (O_1458,N_24956,N_24837);
nor UO_1459 (O_1459,N_24812,N_24866);
nand UO_1460 (O_1460,N_24515,N_24545);
or UO_1461 (O_1461,N_24679,N_24527);
nor UO_1462 (O_1462,N_24478,N_24683);
xnor UO_1463 (O_1463,N_24644,N_24655);
nor UO_1464 (O_1464,N_24830,N_24392);
nand UO_1465 (O_1465,N_24486,N_24568);
nand UO_1466 (O_1466,N_24614,N_24609);
nand UO_1467 (O_1467,N_24724,N_24387);
or UO_1468 (O_1468,N_24746,N_24596);
and UO_1469 (O_1469,N_24927,N_24551);
nand UO_1470 (O_1470,N_24950,N_24534);
nor UO_1471 (O_1471,N_24456,N_24919);
xnor UO_1472 (O_1472,N_24546,N_24535);
and UO_1473 (O_1473,N_24697,N_24849);
and UO_1474 (O_1474,N_24588,N_24792);
and UO_1475 (O_1475,N_24406,N_24761);
and UO_1476 (O_1476,N_24678,N_24648);
nor UO_1477 (O_1477,N_24377,N_24916);
or UO_1478 (O_1478,N_24468,N_24510);
or UO_1479 (O_1479,N_24875,N_24828);
nor UO_1480 (O_1480,N_24460,N_24478);
nand UO_1481 (O_1481,N_24467,N_24696);
nand UO_1482 (O_1482,N_24657,N_24978);
or UO_1483 (O_1483,N_24713,N_24820);
nor UO_1484 (O_1484,N_24719,N_24730);
nor UO_1485 (O_1485,N_24748,N_24912);
xnor UO_1486 (O_1486,N_24997,N_24663);
nor UO_1487 (O_1487,N_24396,N_24999);
and UO_1488 (O_1488,N_24952,N_24992);
and UO_1489 (O_1489,N_24569,N_24768);
nor UO_1490 (O_1490,N_24488,N_24960);
nor UO_1491 (O_1491,N_24470,N_24650);
and UO_1492 (O_1492,N_24722,N_24894);
nor UO_1493 (O_1493,N_24904,N_24952);
or UO_1494 (O_1494,N_24970,N_24471);
xor UO_1495 (O_1495,N_24448,N_24618);
nor UO_1496 (O_1496,N_24646,N_24570);
or UO_1497 (O_1497,N_24770,N_24761);
nor UO_1498 (O_1498,N_24892,N_24944);
xnor UO_1499 (O_1499,N_24438,N_24763);
and UO_1500 (O_1500,N_24855,N_24892);
nor UO_1501 (O_1501,N_24416,N_24567);
nand UO_1502 (O_1502,N_24452,N_24570);
or UO_1503 (O_1503,N_24863,N_24637);
nand UO_1504 (O_1504,N_24878,N_24377);
nand UO_1505 (O_1505,N_24799,N_24434);
nor UO_1506 (O_1506,N_24985,N_24763);
nor UO_1507 (O_1507,N_24854,N_24784);
nand UO_1508 (O_1508,N_24558,N_24924);
nor UO_1509 (O_1509,N_24816,N_24471);
xor UO_1510 (O_1510,N_24926,N_24874);
xor UO_1511 (O_1511,N_24964,N_24398);
nor UO_1512 (O_1512,N_24714,N_24619);
xnor UO_1513 (O_1513,N_24860,N_24820);
xor UO_1514 (O_1514,N_24394,N_24556);
xnor UO_1515 (O_1515,N_24455,N_24520);
and UO_1516 (O_1516,N_24518,N_24459);
xnor UO_1517 (O_1517,N_24567,N_24579);
or UO_1518 (O_1518,N_24397,N_24464);
or UO_1519 (O_1519,N_24395,N_24702);
or UO_1520 (O_1520,N_24591,N_24898);
and UO_1521 (O_1521,N_24717,N_24564);
and UO_1522 (O_1522,N_24839,N_24737);
xor UO_1523 (O_1523,N_24802,N_24430);
xnor UO_1524 (O_1524,N_24776,N_24846);
nor UO_1525 (O_1525,N_24686,N_24464);
xnor UO_1526 (O_1526,N_24393,N_24710);
nor UO_1527 (O_1527,N_24525,N_24701);
or UO_1528 (O_1528,N_24849,N_24387);
or UO_1529 (O_1529,N_24375,N_24879);
nand UO_1530 (O_1530,N_24886,N_24943);
nor UO_1531 (O_1531,N_24785,N_24871);
nand UO_1532 (O_1532,N_24954,N_24538);
xnor UO_1533 (O_1533,N_24388,N_24468);
nand UO_1534 (O_1534,N_24984,N_24396);
nor UO_1535 (O_1535,N_24952,N_24693);
nor UO_1536 (O_1536,N_24595,N_24613);
and UO_1537 (O_1537,N_24749,N_24826);
nand UO_1538 (O_1538,N_24716,N_24479);
nand UO_1539 (O_1539,N_24493,N_24980);
xnor UO_1540 (O_1540,N_24407,N_24858);
nand UO_1541 (O_1541,N_24767,N_24606);
xnor UO_1542 (O_1542,N_24678,N_24531);
xnor UO_1543 (O_1543,N_24592,N_24835);
nand UO_1544 (O_1544,N_24881,N_24414);
and UO_1545 (O_1545,N_24494,N_24716);
and UO_1546 (O_1546,N_24666,N_24535);
nand UO_1547 (O_1547,N_24875,N_24395);
xnor UO_1548 (O_1548,N_24748,N_24537);
xor UO_1549 (O_1549,N_24641,N_24585);
nand UO_1550 (O_1550,N_24544,N_24408);
and UO_1551 (O_1551,N_24490,N_24802);
and UO_1552 (O_1552,N_24962,N_24753);
or UO_1553 (O_1553,N_24478,N_24826);
and UO_1554 (O_1554,N_24593,N_24417);
nand UO_1555 (O_1555,N_24628,N_24876);
and UO_1556 (O_1556,N_24869,N_24858);
and UO_1557 (O_1557,N_24411,N_24629);
xnor UO_1558 (O_1558,N_24562,N_24609);
and UO_1559 (O_1559,N_24461,N_24791);
xnor UO_1560 (O_1560,N_24739,N_24918);
and UO_1561 (O_1561,N_24862,N_24958);
or UO_1562 (O_1562,N_24991,N_24557);
and UO_1563 (O_1563,N_24827,N_24402);
and UO_1564 (O_1564,N_24973,N_24570);
nor UO_1565 (O_1565,N_24887,N_24687);
and UO_1566 (O_1566,N_24508,N_24572);
or UO_1567 (O_1567,N_24500,N_24916);
nor UO_1568 (O_1568,N_24507,N_24480);
and UO_1569 (O_1569,N_24854,N_24972);
nand UO_1570 (O_1570,N_24979,N_24413);
and UO_1571 (O_1571,N_24736,N_24673);
nand UO_1572 (O_1572,N_24377,N_24698);
and UO_1573 (O_1573,N_24560,N_24977);
nor UO_1574 (O_1574,N_24977,N_24531);
xnor UO_1575 (O_1575,N_24777,N_24972);
nor UO_1576 (O_1576,N_24568,N_24591);
nor UO_1577 (O_1577,N_24668,N_24866);
nand UO_1578 (O_1578,N_24812,N_24516);
xnor UO_1579 (O_1579,N_24950,N_24844);
xor UO_1580 (O_1580,N_24998,N_24574);
xnor UO_1581 (O_1581,N_24744,N_24757);
or UO_1582 (O_1582,N_24649,N_24518);
nand UO_1583 (O_1583,N_24935,N_24510);
xnor UO_1584 (O_1584,N_24846,N_24420);
and UO_1585 (O_1585,N_24541,N_24762);
nand UO_1586 (O_1586,N_24552,N_24842);
and UO_1587 (O_1587,N_24964,N_24856);
nand UO_1588 (O_1588,N_24595,N_24991);
nor UO_1589 (O_1589,N_24992,N_24993);
nor UO_1590 (O_1590,N_24962,N_24504);
or UO_1591 (O_1591,N_24387,N_24460);
xor UO_1592 (O_1592,N_24702,N_24650);
or UO_1593 (O_1593,N_24508,N_24893);
xnor UO_1594 (O_1594,N_24887,N_24645);
and UO_1595 (O_1595,N_24450,N_24844);
nor UO_1596 (O_1596,N_24981,N_24707);
nor UO_1597 (O_1597,N_24651,N_24947);
nand UO_1598 (O_1598,N_24502,N_24945);
nor UO_1599 (O_1599,N_24412,N_24492);
nor UO_1600 (O_1600,N_24693,N_24382);
and UO_1601 (O_1601,N_24990,N_24838);
or UO_1602 (O_1602,N_24416,N_24740);
and UO_1603 (O_1603,N_24820,N_24591);
nand UO_1604 (O_1604,N_24585,N_24858);
xnor UO_1605 (O_1605,N_24687,N_24959);
and UO_1606 (O_1606,N_24397,N_24376);
or UO_1607 (O_1607,N_24936,N_24707);
or UO_1608 (O_1608,N_24386,N_24544);
or UO_1609 (O_1609,N_24599,N_24810);
xnor UO_1610 (O_1610,N_24839,N_24888);
nand UO_1611 (O_1611,N_24726,N_24492);
and UO_1612 (O_1612,N_24881,N_24601);
xnor UO_1613 (O_1613,N_24432,N_24939);
nor UO_1614 (O_1614,N_24569,N_24983);
and UO_1615 (O_1615,N_24388,N_24404);
nand UO_1616 (O_1616,N_24510,N_24996);
or UO_1617 (O_1617,N_24558,N_24706);
or UO_1618 (O_1618,N_24756,N_24764);
or UO_1619 (O_1619,N_24805,N_24960);
nor UO_1620 (O_1620,N_24747,N_24502);
and UO_1621 (O_1621,N_24629,N_24991);
or UO_1622 (O_1622,N_24991,N_24684);
nor UO_1623 (O_1623,N_24513,N_24388);
and UO_1624 (O_1624,N_24510,N_24852);
nor UO_1625 (O_1625,N_24477,N_24473);
and UO_1626 (O_1626,N_24561,N_24397);
or UO_1627 (O_1627,N_24999,N_24565);
or UO_1628 (O_1628,N_24596,N_24985);
xnor UO_1629 (O_1629,N_24852,N_24769);
nand UO_1630 (O_1630,N_24569,N_24598);
nand UO_1631 (O_1631,N_24729,N_24496);
or UO_1632 (O_1632,N_24663,N_24438);
and UO_1633 (O_1633,N_24502,N_24932);
xnor UO_1634 (O_1634,N_24503,N_24405);
xnor UO_1635 (O_1635,N_24400,N_24987);
xnor UO_1636 (O_1636,N_24757,N_24384);
xnor UO_1637 (O_1637,N_24816,N_24724);
nor UO_1638 (O_1638,N_24774,N_24816);
xor UO_1639 (O_1639,N_24849,N_24831);
and UO_1640 (O_1640,N_24895,N_24882);
nand UO_1641 (O_1641,N_24431,N_24905);
nand UO_1642 (O_1642,N_24566,N_24405);
or UO_1643 (O_1643,N_24768,N_24990);
or UO_1644 (O_1644,N_24400,N_24910);
xor UO_1645 (O_1645,N_24399,N_24608);
nand UO_1646 (O_1646,N_24967,N_24874);
nand UO_1647 (O_1647,N_24749,N_24432);
nand UO_1648 (O_1648,N_24473,N_24781);
or UO_1649 (O_1649,N_24583,N_24811);
and UO_1650 (O_1650,N_24834,N_24870);
nor UO_1651 (O_1651,N_24764,N_24600);
xnor UO_1652 (O_1652,N_24997,N_24421);
or UO_1653 (O_1653,N_24900,N_24380);
xor UO_1654 (O_1654,N_24697,N_24743);
xnor UO_1655 (O_1655,N_24476,N_24882);
xor UO_1656 (O_1656,N_24434,N_24543);
xnor UO_1657 (O_1657,N_24663,N_24904);
nor UO_1658 (O_1658,N_24973,N_24940);
nand UO_1659 (O_1659,N_24750,N_24810);
xnor UO_1660 (O_1660,N_24690,N_24997);
and UO_1661 (O_1661,N_24599,N_24674);
nor UO_1662 (O_1662,N_24816,N_24716);
nor UO_1663 (O_1663,N_24425,N_24732);
nor UO_1664 (O_1664,N_24464,N_24929);
nand UO_1665 (O_1665,N_24456,N_24682);
nor UO_1666 (O_1666,N_24863,N_24687);
nor UO_1667 (O_1667,N_24452,N_24380);
or UO_1668 (O_1668,N_24496,N_24705);
nor UO_1669 (O_1669,N_24783,N_24648);
nand UO_1670 (O_1670,N_24807,N_24920);
and UO_1671 (O_1671,N_24865,N_24899);
xnor UO_1672 (O_1672,N_24997,N_24857);
xor UO_1673 (O_1673,N_24999,N_24430);
xnor UO_1674 (O_1674,N_24453,N_24999);
nand UO_1675 (O_1675,N_24636,N_24496);
xnor UO_1676 (O_1676,N_24740,N_24953);
nand UO_1677 (O_1677,N_24883,N_24790);
nand UO_1678 (O_1678,N_24651,N_24975);
nand UO_1679 (O_1679,N_24476,N_24683);
nand UO_1680 (O_1680,N_24979,N_24590);
nand UO_1681 (O_1681,N_24772,N_24831);
or UO_1682 (O_1682,N_24382,N_24732);
and UO_1683 (O_1683,N_24608,N_24557);
xnor UO_1684 (O_1684,N_24419,N_24569);
nor UO_1685 (O_1685,N_24861,N_24638);
nor UO_1686 (O_1686,N_24909,N_24967);
nand UO_1687 (O_1687,N_24558,N_24795);
and UO_1688 (O_1688,N_24529,N_24988);
xor UO_1689 (O_1689,N_24780,N_24535);
nand UO_1690 (O_1690,N_24661,N_24492);
and UO_1691 (O_1691,N_24444,N_24868);
or UO_1692 (O_1692,N_24951,N_24959);
or UO_1693 (O_1693,N_24659,N_24743);
nand UO_1694 (O_1694,N_24755,N_24628);
and UO_1695 (O_1695,N_24955,N_24634);
xnor UO_1696 (O_1696,N_24905,N_24405);
nand UO_1697 (O_1697,N_24837,N_24400);
or UO_1698 (O_1698,N_24984,N_24909);
nand UO_1699 (O_1699,N_24695,N_24952);
nand UO_1700 (O_1700,N_24709,N_24857);
xnor UO_1701 (O_1701,N_24490,N_24535);
or UO_1702 (O_1702,N_24384,N_24567);
nand UO_1703 (O_1703,N_24860,N_24671);
xnor UO_1704 (O_1704,N_24559,N_24918);
and UO_1705 (O_1705,N_24916,N_24465);
nand UO_1706 (O_1706,N_24476,N_24946);
and UO_1707 (O_1707,N_24923,N_24764);
xor UO_1708 (O_1708,N_24641,N_24433);
nor UO_1709 (O_1709,N_24898,N_24856);
and UO_1710 (O_1710,N_24689,N_24654);
nand UO_1711 (O_1711,N_24889,N_24530);
and UO_1712 (O_1712,N_24602,N_24607);
xnor UO_1713 (O_1713,N_24415,N_24739);
and UO_1714 (O_1714,N_24663,N_24891);
and UO_1715 (O_1715,N_24385,N_24722);
nor UO_1716 (O_1716,N_24494,N_24819);
or UO_1717 (O_1717,N_24436,N_24732);
xnor UO_1718 (O_1718,N_24470,N_24484);
or UO_1719 (O_1719,N_24470,N_24513);
nor UO_1720 (O_1720,N_24779,N_24730);
xor UO_1721 (O_1721,N_24674,N_24448);
or UO_1722 (O_1722,N_24828,N_24639);
nor UO_1723 (O_1723,N_24753,N_24539);
nand UO_1724 (O_1724,N_24899,N_24612);
nor UO_1725 (O_1725,N_24521,N_24834);
and UO_1726 (O_1726,N_24718,N_24531);
nand UO_1727 (O_1727,N_24872,N_24612);
nand UO_1728 (O_1728,N_24884,N_24914);
xor UO_1729 (O_1729,N_24417,N_24776);
xor UO_1730 (O_1730,N_24434,N_24770);
nand UO_1731 (O_1731,N_24891,N_24621);
nor UO_1732 (O_1732,N_24979,N_24469);
nor UO_1733 (O_1733,N_24448,N_24690);
nor UO_1734 (O_1734,N_24465,N_24722);
and UO_1735 (O_1735,N_24555,N_24663);
or UO_1736 (O_1736,N_24770,N_24389);
and UO_1737 (O_1737,N_24381,N_24927);
nand UO_1738 (O_1738,N_24681,N_24840);
nand UO_1739 (O_1739,N_24821,N_24637);
nand UO_1740 (O_1740,N_24538,N_24713);
nand UO_1741 (O_1741,N_24565,N_24605);
nand UO_1742 (O_1742,N_24784,N_24863);
xnor UO_1743 (O_1743,N_24776,N_24753);
and UO_1744 (O_1744,N_24901,N_24792);
nor UO_1745 (O_1745,N_24901,N_24956);
nand UO_1746 (O_1746,N_24513,N_24498);
xor UO_1747 (O_1747,N_24687,N_24742);
nor UO_1748 (O_1748,N_24483,N_24814);
and UO_1749 (O_1749,N_24937,N_24446);
nand UO_1750 (O_1750,N_24789,N_24414);
or UO_1751 (O_1751,N_24643,N_24385);
nand UO_1752 (O_1752,N_24456,N_24636);
nor UO_1753 (O_1753,N_24681,N_24640);
nand UO_1754 (O_1754,N_24647,N_24828);
nand UO_1755 (O_1755,N_24788,N_24594);
or UO_1756 (O_1756,N_24966,N_24709);
nor UO_1757 (O_1757,N_24971,N_24906);
xnor UO_1758 (O_1758,N_24647,N_24500);
or UO_1759 (O_1759,N_24691,N_24914);
nand UO_1760 (O_1760,N_24466,N_24438);
nand UO_1761 (O_1761,N_24532,N_24502);
and UO_1762 (O_1762,N_24667,N_24965);
nor UO_1763 (O_1763,N_24788,N_24755);
nand UO_1764 (O_1764,N_24589,N_24720);
nand UO_1765 (O_1765,N_24411,N_24931);
xor UO_1766 (O_1766,N_24824,N_24845);
or UO_1767 (O_1767,N_24918,N_24394);
xnor UO_1768 (O_1768,N_24867,N_24678);
and UO_1769 (O_1769,N_24403,N_24804);
xor UO_1770 (O_1770,N_24674,N_24403);
nor UO_1771 (O_1771,N_24730,N_24416);
or UO_1772 (O_1772,N_24750,N_24926);
xor UO_1773 (O_1773,N_24898,N_24701);
or UO_1774 (O_1774,N_24850,N_24466);
or UO_1775 (O_1775,N_24510,N_24635);
xnor UO_1776 (O_1776,N_24646,N_24607);
and UO_1777 (O_1777,N_24882,N_24677);
xnor UO_1778 (O_1778,N_24916,N_24721);
nor UO_1779 (O_1779,N_24507,N_24917);
nor UO_1780 (O_1780,N_24469,N_24595);
nand UO_1781 (O_1781,N_24897,N_24497);
and UO_1782 (O_1782,N_24788,N_24412);
nand UO_1783 (O_1783,N_24844,N_24755);
xor UO_1784 (O_1784,N_24389,N_24997);
or UO_1785 (O_1785,N_24862,N_24908);
nor UO_1786 (O_1786,N_24605,N_24383);
or UO_1787 (O_1787,N_24755,N_24580);
and UO_1788 (O_1788,N_24871,N_24974);
or UO_1789 (O_1789,N_24475,N_24620);
and UO_1790 (O_1790,N_24745,N_24434);
and UO_1791 (O_1791,N_24968,N_24484);
nand UO_1792 (O_1792,N_24549,N_24759);
or UO_1793 (O_1793,N_24645,N_24402);
and UO_1794 (O_1794,N_24705,N_24536);
nand UO_1795 (O_1795,N_24572,N_24811);
or UO_1796 (O_1796,N_24864,N_24656);
nor UO_1797 (O_1797,N_24615,N_24686);
nor UO_1798 (O_1798,N_24472,N_24952);
nor UO_1799 (O_1799,N_24897,N_24967);
nand UO_1800 (O_1800,N_24463,N_24957);
or UO_1801 (O_1801,N_24390,N_24904);
xnor UO_1802 (O_1802,N_24559,N_24743);
or UO_1803 (O_1803,N_24727,N_24918);
or UO_1804 (O_1804,N_24487,N_24968);
xnor UO_1805 (O_1805,N_24541,N_24734);
nor UO_1806 (O_1806,N_24869,N_24456);
xor UO_1807 (O_1807,N_24742,N_24541);
nor UO_1808 (O_1808,N_24420,N_24825);
xnor UO_1809 (O_1809,N_24830,N_24893);
xnor UO_1810 (O_1810,N_24748,N_24476);
nand UO_1811 (O_1811,N_24491,N_24945);
nand UO_1812 (O_1812,N_24791,N_24435);
and UO_1813 (O_1813,N_24870,N_24973);
xor UO_1814 (O_1814,N_24778,N_24734);
or UO_1815 (O_1815,N_24957,N_24468);
nand UO_1816 (O_1816,N_24525,N_24547);
nand UO_1817 (O_1817,N_24648,N_24499);
or UO_1818 (O_1818,N_24696,N_24841);
nor UO_1819 (O_1819,N_24596,N_24719);
nor UO_1820 (O_1820,N_24591,N_24425);
and UO_1821 (O_1821,N_24870,N_24855);
nand UO_1822 (O_1822,N_24543,N_24792);
xnor UO_1823 (O_1823,N_24852,N_24571);
nand UO_1824 (O_1824,N_24413,N_24903);
and UO_1825 (O_1825,N_24826,N_24477);
nor UO_1826 (O_1826,N_24423,N_24803);
nor UO_1827 (O_1827,N_24414,N_24767);
or UO_1828 (O_1828,N_24683,N_24728);
nand UO_1829 (O_1829,N_24639,N_24669);
nand UO_1830 (O_1830,N_24661,N_24801);
and UO_1831 (O_1831,N_24960,N_24802);
or UO_1832 (O_1832,N_24580,N_24447);
and UO_1833 (O_1833,N_24728,N_24636);
and UO_1834 (O_1834,N_24738,N_24673);
nor UO_1835 (O_1835,N_24995,N_24925);
nand UO_1836 (O_1836,N_24685,N_24778);
nand UO_1837 (O_1837,N_24792,N_24790);
nor UO_1838 (O_1838,N_24458,N_24421);
xnor UO_1839 (O_1839,N_24954,N_24608);
xor UO_1840 (O_1840,N_24982,N_24962);
and UO_1841 (O_1841,N_24570,N_24942);
nor UO_1842 (O_1842,N_24586,N_24378);
nand UO_1843 (O_1843,N_24996,N_24400);
or UO_1844 (O_1844,N_24792,N_24693);
nand UO_1845 (O_1845,N_24471,N_24623);
xnor UO_1846 (O_1846,N_24922,N_24903);
and UO_1847 (O_1847,N_24757,N_24822);
nor UO_1848 (O_1848,N_24978,N_24582);
nor UO_1849 (O_1849,N_24456,N_24841);
xor UO_1850 (O_1850,N_24846,N_24641);
or UO_1851 (O_1851,N_24759,N_24727);
nand UO_1852 (O_1852,N_24458,N_24466);
or UO_1853 (O_1853,N_24479,N_24919);
and UO_1854 (O_1854,N_24998,N_24745);
nor UO_1855 (O_1855,N_24837,N_24621);
and UO_1856 (O_1856,N_24552,N_24816);
nor UO_1857 (O_1857,N_24887,N_24804);
nand UO_1858 (O_1858,N_24627,N_24772);
xnor UO_1859 (O_1859,N_24746,N_24904);
nand UO_1860 (O_1860,N_24536,N_24388);
nor UO_1861 (O_1861,N_24916,N_24954);
nor UO_1862 (O_1862,N_24628,N_24870);
or UO_1863 (O_1863,N_24408,N_24766);
xnor UO_1864 (O_1864,N_24761,N_24599);
nand UO_1865 (O_1865,N_24456,N_24662);
or UO_1866 (O_1866,N_24411,N_24628);
nor UO_1867 (O_1867,N_24907,N_24882);
and UO_1868 (O_1868,N_24492,N_24634);
or UO_1869 (O_1869,N_24991,N_24920);
xor UO_1870 (O_1870,N_24581,N_24970);
or UO_1871 (O_1871,N_24598,N_24870);
nand UO_1872 (O_1872,N_24656,N_24889);
nand UO_1873 (O_1873,N_24973,N_24469);
or UO_1874 (O_1874,N_24994,N_24949);
xnor UO_1875 (O_1875,N_24585,N_24592);
or UO_1876 (O_1876,N_24616,N_24704);
xnor UO_1877 (O_1877,N_24417,N_24652);
or UO_1878 (O_1878,N_24507,N_24963);
nand UO_1879 (O_1879,N_24414,N_24589);
nor UO_1880 (O_1880,N_24705,N_24951);
nand UO_1881 (O_1881,N_24782,N_24818);
xor UO_1882 (O_1882,N_24669,N_24464);
and UO_1883 (O_1883,N_24928,N_24726);
nand UO_1884 (O_1884,N_24952,N_24652);
nor UO_1885 (O_1885,N_24448,N_24521);
xor UO_1886 (O_1886,N_24631,N_24685);
xor UO_1887 (O_1887,N_24556,N_24732);
xor UO_1888 (O_1888,N_24859,N_24928);
nor UO_1889 (O_1889,N_24794,N_24962);
nand UO_1890 (O_1890,N_24628,N_24902);
or UO_1891 (O_1891,N_24416,N_24496);
xnor UO_1892 (O_1892,N_24735,N_24517);
nand UO_1893 (O_1893,N_24782,N_24805);
and UO_1894 (O_1894,N_24943,N_24686);
or UO_1895 (O_1895,N_24497,N_24921);
and UO_1896 (O_1896,N_24663,N_24709);
nor UO_1897 (O_1897,N_24921,N_24788);
nor UO_1898 (O_1898,N_24476,N_24552);
and UO_1899 (O_1899,N_24806,N_24550);
and UO_1900 (O_1900,N_24734,N_24762);
xor UO_1901 (O_1901,N_24465,N_24931);
and UO_1902 (O_1902,N_24920,N_24476);
or UO_1903 (O_1903,N_24606,N_24651);
nor UO_1904 (O_1904,N_24781,N_24820);
nor UO_1905 (O_1905,N_24410,N_24996);
nand UO_1906 (O_1906,N_24999,N_24766);
nor UO_1907 (O_1907,N_24782,N_24597);
nor UO_1908 (O_1908,N_24658,N_24767);
nor UO_1909 (O_1909,N_24868,N_24961);
xnor UO_1910 (O_1910,N_24929,N_24776);
or UO_1911 (O_1911,N_24847,N_24589);
or UO_1912 (O_1912,N_24969,N_24685);
nor UO_1913 (O_1913,N_24893,N_24488);
nor UO_1914 (O_1914,N_24905,N_24976);
or UO_1915 (O_1915,N_24819,N_24507);
nand UO_1916 (O_1916,N_24608,N_24866);
xnor UO_1917 (O_1917,N_24386,N_24550);
nand UO_1918 (O_1918,N_24922,N_24627);
nand UO_1919 (O_1919,N_24507,N_24837);
nor UO_1920 (O_1920,N_24439,N_24414);
or UO_1921 (O_1921,N_24632,N_24762);
nand UO_1922 (O_1922,N_24552,N_24787);
xnor UO_1923 (O_1923,N_24878,N_24442);
nand UO_1924 (O_1924,N_24927,N_24812);
xor UO_1925 (O_1925,N_24848,N_24527);
and UO_1926 (O_1926,N_24448,N_24724);
xor UO_1927 (O_1927,N_24561,N_24675);
nand UO_1928 (O_1928,N_24938,N_24845);
or UO_1929 (O_1929,N_24504,N_24791);
or UO_1930 (O_1930,N_24965,N_24379);
and UO_1931 (O_1931,N_24876,N_24458);
nor UO_1932 (O_1932,N_24660,N_24390);
xnor UO_1933 (O_1933,N_24907,N_24849);
nor UO_1934 (O_1934,N_24531,N_24682);
nand UO_1935 (O_1935,N_24880,N_24590);
nand UO_1936 (O_1936,N_24962,N_24728);
or UO_1937 (O_1937,N_24987,N_24954);
or UO_1938 (O_1938,N_24405,N_24498);
or UO_1939 (O_1939,N_24466,N_24686);
nand UO_1940 (O_1940,N_24570,N_24944);
xor UO_1941 (O_1941,N_24773,N_24815);
or UO_1942 (O_1942,N_24502,N_24808);
or UO_1943 (O_1943,N_24923,N_24864);
and UO_1944 (O_1944,N_24793,N_24653);
nor UO_1945 (O_1945,N_24524,N_24646);
or UO_1946 (O_1946,N_24527,N_24426);
nand UO_1947 (O_1947,N_24515,N_24393);
xor UO_1948 (O_1948,N_24536,N_24684);
nand UO_1949 (O_1949,N_24751,N_24572);
nor UO_1950 (O_1950,N_24562,N_24865);
nand UO_1951 (O_1951,N_24944,N_24834);
and UO_1952 (O_1952,N_24399,N_24923);
or UO_1953 (O_1953,N_24826,N_24958);
nor UO_1954 (O_1954,N_24771,N_24932);
and UO_1955 (O_1955,N_24745,N_24675);
nor UO_1956 (O_1956,N_24421,N_24459);
nor UO_1957 (O_1957,N_24763,N_24854);
xor UO_1958 (O_1958,N_24430,N_24528);
or UO_1959 (O_1959,N_24794,N_24623);
xnor UO_1960 (O_1960,N_24657,N_24909);
xor UO_1961 (O_1961,N_24518,N_24771);
nand UO_1962 (O_1962,N_24939,N_24778);
nor UO_1963 (O_1963,N_24503,N_24784);
nor UO_1964 (O_1964,N_24937,N_24997);
and UO_1965 (O_1965,N_24997,N_24645);
or UO_1966 (O_1966,N_24517,N_24989);
or UO_1967 (O_1967,N_24621,N_24575);
xnor UO_1968 (O_1968,N_24497,N_24863);
or UO_1969 (O_1969,N_24692,N_24942);
and UO_1970 (O_1970,N_24387,N_24872);
nor UO_1971 (O_1971,N_24617,N_24678);
xnor UO_1972 (O_1972,N_24497,N_24386);
nand UO_1973 (O_1973,N_24563,N_24841);
nor UO_1974 (O_1974,N_24784,N_24927);
nand UO_1975 (O_1975,N_24775,N_24897);
nor UO_1976 (O_1976,N_24594,N_24551);
and UO_1977 (O_1977,N_24390,N_24727);
xor UO_1978 (O_1978,N_24571,N_24554);
or UO_1979 (O_1979,N_24484,N_24376);
nor UO_1980 (O_1980,N_24962,N_24886);
or UO_1981 (O_1981,N_24517,N_24778);
or UO_1982 (O_1982,N_24662,N_24573);
and UO_1983 (O_1983,N_24456,N_24774);
nand UO_1984 (O_1984,N_24532,N_24766);
or UO_1985 (O_1985,N_24807,N_24405);
nand UO_1986 (O_1986,N_24395,N_24840);
and UO_1987 (O_1987,N_24636,N_24782);
xor UO_1988 (O_1988,N_24931,N_24709);
nand UO_1989 (O_1989,N_24973,N_24526);
nor UO_1990 (O_1990,N_24676,N_24957);
and UO_1991 (O_1991,N_24445,N_24547);
and UO_1992 (O_1992,N_24556,N_24469);
or UO_1993 (O_1993,N_24595,N_24711);
nor UO_1994 (O_1994,N_24456,N_24380);
nor UO_1995 (O_1995,N_24944,N_24903);
or UO_1996 (O_1996,N_24607,N_24506);
and UO_1997 (O_1997,N_24857,N_24658);
or UO_1998 (O_1998,N_24398,N_24755);
nand UO_1999 (O_1999,N_24512,N_24727);
nor UO_2000 (O_2000,N_24650,N_24560);
or UO_2001 (O_2001,N_24643,N_24832);
nor UO_2002 (O_2002,N_24603,N_24670);
nand UO_2003 (O_2003,N_24736,N_24531);
or UO_2004 (O_2004,N_24681,N_24935);
nor UO_2005 (O_2005,N_24952,N_24588);
nand UO_2006 (O_2006,N_24799,N_24797);
and UO_2007 (O_2007,N_24812,N_24599);
nor UO_2008 (O_2008,N_24622,N_24934);
nand UO_2009 (O_2009,N_24430,N_24867);
or UO_2010 (O_2010,N_24794,N_24677);
nor UO_2011 (O_2011,N_24486,N_24681);
nand UO_2012 (O_2012,N_24645,N_24560);
nor UO_2013 (O_2013,N_24870,N_24636);
xnor UO_2014 (O_2014,N_24735,N_24523);
nor UO_2015 (O_2015,N_24896,N_24856);
xor UO_2016 (O_2016,N_24850,N_24870);
nand UO_2017 (O_2017,N_24915,N_24960);
nor UO_2018 (O_2018,N_24724,N_24453);
nand UO_2019 (O_2019,N_24419,N_24377);
nand UO_2020 (O_2020,N_24728,N_24646);
nand UO_2021 (O_2021,N_24679,N_24610);
or UO_2022 (O_2022,N_24688,N_24440);
nand UO_2023 (O_2023,N_24644,N_24657);
xnor UO_2024 (O_2024,N_24902,N_24797);
xor UO_2025 (O_2025,N_24845,N_24802);
xnor UO_2026 (O_2026,N_24515,N_24944);
xnor UO_2027 (O_2027,N_24907,N_24948);
xnor UO_2028 (O_2028,N_24972,N_24381);
nor UO_2029 (O_2029,N_24530,N_24696);
or UO_2030 (O_2030,N_24697,N_24742);
nor UO_2031 (O_2031,N_24915,N_24790);
nand UO_2032 (O_2032,N_24593,N_24621);
nand UO_2033 (O_2033,N_24488,N_24449);
and UO_2034 (O_2034,N_24534,N_24981);
nand UO_2035 (O_2035,N_24959,N_24636);
and UO_2036 (O_2036,N_24449,N_24923);
nand UO_2037 (O_2037,N_24981,N_24969);
nand UO_2038 (O_2038,N_24981,N_24404);
xnor UO_2039 (O_2039,N_24968,N_24718);
xor UO_2040 (O_2040,N_24595,N_24887);
xnor UO_2041 (O_2041,N_24893,N_24563);
nor UO_2042 (O_2042,N_24668,N_24933);
xnor UO_2043 (O_2043,N_24749,N_24941);
nand UO_2044 (O_2044,N_24860,N_24630);
nor UO_2045 (O_2045,N_24680,N_24862);
xnor UO_2046 (O_2046,N_24654,N_24983);
or UO_2047 (O_2047,N_24805,N_24380);
xor UO_2048 (O_2048,N_24975,N_24434);
or UO_2049 (O_2049,N_24645,N_24672);
or UO_2050 (O_2050,N_24933,N_24450);
or UO_2051 (O_2051,N_24801,N_24378);
or UO_2052 (O_2052,N_24761,N_24609);
nor UO_2053 (O_2053,N_24726,N_24766);
or UO_2054 (O_2054,N_24710,N_24756);
xnor UO_2055 (O_2055,N_24770,N_24913);
xnor UO_2056 (O_2056,N_24965,N_24758);
and UO_2057 (O_2057,N_24805,N_24993);
or UO_2058 (O_2058,N_24411,N_24394);
xnor UO_2059 (O_2059,N_24805,N_24922);
or UO_2060 (O_2060,N_24445,N_24524);
and UO_2061 (O_2061,N_24459,N_24944);
xnor UO_2062 (O_2062,N_24761,N_24377);
nor UO_2063 (O_2063,N_24543,N_24596);
and UO_2064 (O_2064,N_24655,N_24407);
xor UO_2065 (O_2065,N_24886,N_24624);
and UO_2066 (O_2066,N_24655,N_24966);
or UO_2067 (O_2067,N_24496,N_24782);
nand UO_2068 (O_2068,N_24929,N_24997);
nor UO_2069 (O_2069,N_24927,N_24835);
nand UO_2070 (O_2070,N_24868,N_24452);
or UO_2071 (O_2071,N_24951,N_24516);
or UO_2072 (O_2072,N_24513,N_24916);
or UO_2073 (O_2073,N_24950,N_24742);
nor UO_2074 (O_2074,N_24981,N_24911);
and UO_2075 (O_2075,N_24461,N_24971);
xor UO_2076 (O_2076,N_24604,N_24504);
nor UO_2077 (O_2077,N_24406,N_24729);
and UO_2078 (O_2078,N_24381,N_24784);
nor UO_2079 (O_2079,N_24947,N_24630);
or UO_2080 (O_2080,N_24861,N_24574);
or UO_2081 (O_2081,N_24563,N_24870);
xnor UO_2082 (O_2082,N_24892,N_24982);
nor UO_2083 (O_2083,N_24543,N_24456);
or UO_2084 (O_2084,N_24583,N_24781);
xnor UO_2085 (O_2085,N_24560,N_24905);
and UO_2086 (O_2086,N_24935,N_24497);
and UO_2087 (O_2087,N_24412,N_24782);
nand UO_2088 (O_2088,N_24984,N_24510);
xnor UO_2089 (O_2089,N_24898,N_24697);
nand UO_2090 (O_2090,N_24578,N_24441);
or UO_2091 (O_2091,N_24542,N_24412);
nand UO_2092 (O_2092,N_24383,N_24895);
or UO_2093 (O_2093,N_24448,N_24904);
nand UO_2094 (O_2094,N_24575,N_24917);
nor UO_2095 (O_2095,N_24399,N_24447);
and UO_2096 (O_2096,N_24735,N_24578);
nand UO_2097 (O_2097,N_24565,N_24580);
nor UO_2098 (O_2098,N_24516,N_24836);
nand UO_2099 (O_2099,N_24589,N_24517);
xnor UO_2100 (O_2100,N_24955,N_24868);
and UO_2101 (O_2101,N_24893,N_24896);
nand UO_2102 (O_2102,N_24724,N_24679);
or UO_2103 (O_2103,N_24440,N_24456);
or UO_2104 (O_2104,N_24655,N_24735);
nor UO_2105 (O_2105,N_24732,N_24635);
nor UO_2106 (O_2106,N_24387,N_24780);
xor UO_2107 (O_2107,N_24399,N_24814);
xnor UO_2108 (O_2108,N_24999,N_24642);
nand UO_2109 (O_2109,N_24548,N_24407);
nand UO_2110 (O_2110,N_24809,N_24453);
or UO_2111 (O_2111,N_24488,N_24430);
or UO_2112 (O_2112,N_24430,N_24970);
and UO_2113 (O_2113,N_24890,N_24826);
nand UO_2114 (O_2114,N_24414,N_24460);
xor UO_2115 (O_2115,N_24964,N_24936);
nand UO_2116 (O_2116,N_24865,N_24975);
nor UO_2117 (O_2117,N_24758,N_24550);
or UO_2118 (O_2118,N_24886,N_24746);
xnor UO_2119 (O_2119,N_24485,N_24974);
and UO_2120 (O_2120,N_24757,N_24407);
or UO_2121 (O_2121,N_24812,N_24838);
nand UO_2122 (O_2122,N_24772,N_24787);
nor UO_2123 (O_2123,N_24917,N_24846);
or UO_2124 (O_2124,N_24820,N_24845);
nor UO_2125 (O_2125,N_24971,N_24612);
nor UO_2126 (O_2126,N_24932,N_24486);
or UO_2127 (O_2127,N_24538,N_24946);
xor UO_2128 (O_2128,N_24952,N_24690);
or UO_2129 (O_2129,N_24879,N_24474);
xnor UO_2130 (O_2130,N_24646,N_24943);
xnor UO_2131 (O_2131,N_24942,N_24926);
or UO_2132 (O_2132,N_24500,N_24385);
or UO_2133 (O_2133,N_24733,N_24714);
or UO_2134 (O_2134,N_24806,N_24641);
and UO_2135 (O_2135,N_24451,N_24663);
nand UO_2136 (O_2136,N_24879,N_24480);
and UO_2137 (O_2137,N_24779,N_24951);
xor UO_2138 (O_2138,N_24766,N_24518);
nor UO_2139 (O_2139,N_24765,N_24435);
xnor UO_2140 (O_2140,N_24819,N_24491);
and UO_2141 (O_2141,N_24860,N_24386);
xor UO_2142 (O_2142,N_24702,N_24615);
and UO_2143 (O_2143,N_24488,N_24462);
or UO_2144 (O_2144,N_24591,N_24684);
xnor UO_2145 (O_2145,N_24715,N_24558);
xnor UO_2146 (O_2146,N_24376,N_24902);
and UO_2147 (O_2147,N_24830,N_24703);
and UO_2148 (O_2148,N_24985,N_24644);
nor UO_2149 (O_2149,N_24518,N_24497);
nor UO_2150 (O_2150,N_24509,N_24527);
nand UO_2151 (O_2151,N_24786,N_24553);
nand UO_2152 (O_2152,N_24655,N_24926);
nor UO_2153 (O_2153,N_24489,N_24897);
nor UO_2154 (O_2154,N_24401,N_24801);
nor UO_2155 (O_2155,N_24905,N_24449);
and UO_2156 (O_2156,N_24635,N_24956);
xnor UO_2157 (O_2157,N_24935,N_24414);
or UO_2158 (O_2158,N_24440,N_24943);
nor UO_2159 (O_2159,N_24938,N_24945);
or UO_2160 (O_2160,N_24962,N_24948);
nand UO_2161 (O_2161,N_24625,N_24925);
xnor UO_2162 (O_2162,N_24919,N_24761);
nand UO_2163 (O_2163,N_24968,N_24740);
or UO_2164 (O_2164,N_24613,N_24759);
or UO_2165 (O_2165,N_24765,N_24835);
nor UO_2166 (O_2166,N_24461,N_24890);
nor UO_2167 (O_2167,N_24498,N_24559);
nand UO_2168 (O_2168,N_24810,N_24740);
or UO_2169 (O_2169,N_24783,N_24683);
xor UO_2170 (O_2170,N_24837,N_24673);
nor UO_2171 (O_2171,N_24652,N_24529);
or UO_2172 (O_2172,N_24858,N_24863);
nand UO_2173 (O_2173,N_24922,N_24553);
and UO_2174 (O_2174,N_24786,N_24692);
nand UO_2175 (O_2175,N_24876,N_24542);
nand UO_2176 (O_2176,N_24928,N_24488);
or UO_2177 (O_2177,N_24852,N_24690);
or UO_2178 (O_2178,N_24738,N_24542);
and UO_2179 (O_2179,N_24692,N_24836);
xnor UO_2180 (O_2180,N_24830,N_24661);
or UO_2181 (O_2181,N_24524,N_24816);
xnor UO_2182 (O_2182,N_24512,N_24397);
and UO_2183 (O_2183,N_24805,N_24378);
and UO_2184 (O_2184,N_24503,N_24755);
and UO_2185 (O_2185,N_24930,N_24573);
or UO_2186 (O_2186,N_24575,N_24469);
nand UO_2187 (O_2187,N_24819,N_24771);
or UO_2188 (O_2188,N_24579,N_24589);
and UO_2189 (O_2189,N_24378,N_24822);
nor UO_2190 (O_2190,N_24849,N_24635);
nand UO_2191 (O_2191,N_24453,N_24746);
and UO_2192 (O_2192,N_24694,N_24950);
and UO_2193 (O_2193,N_24631,N_24421);
xnor UO_2194 (O_2194,N_24702,N_24392);
and UO_2195 (O_2195,N_24570,N_24384);
xnor UO_2196 (O_2196,N_24784,N_24792);
or UO_2197 (O_2197,N_24811,N_24559);
nor UO_2198 (O_2198,N_24542,N_24851);
nor UO_2199 (O_2199,N_24830,N_24458);
or UO_2200 (O_2200,N_24656,N_24666);
nor UO_2201 (O_2201,N_24742,N_24569);
or UO_2202 (O_2202,N_24411,N_24796);
nor UO_2203 (O_2203,N_24851,N_24527);
and UO_2204 (O_2204,N_24463,N_24412);
nor UO_2205 (O_2205,N_24389,N_24704);
nand UO_2206 (O_2206,N_24862,N_24749);
and UO_2207 (O_2207,N_24419,N_24389);
or UO_2208 (O_2208,N_24987,N_24644);
or UO_2209 (O_2209,N_24792,N_24470);
nand UO_2210 (O_2210,N_24497,N_24934);
and UO_2211 (O_2211,N_24738,N_24456);
nor UO_2212 (O_2212,N_24837,N_24872);
xnor UO_2213 (O_2213,N_24552,N_24460);
nand UO_2214 (O_2214,N_24861,N_24830);
xor UO_2215 (O_2215,N_24928,N_24421);
nand UO_2216 (O_2216,N_24753,N_24551);
xor UO_2217 (O_2217,N_24581,N_24874);
nor UO_2218 (O_2218,N_24796,N_24569);
or UO_2219 (O_2219,N_24599,N_24407);
nand UO_2220 (O_2220,N_24379,N_24431);
or UO_2221 (O_2221,N_24616,N_24657);
xor UO_2222 (O_2222,N_24605,N_24973);
or UO_2223 (O_2223,N_24650,N_24781);
and UO_2224 (O_2224,N_24607,N_24787);
and UO_2225 (O_2225,N_24694,N_24990);
xnor UO_2226 (O_2226,N_24573,N_24886);
or UO_2227 (O_2227,N_24479,N_24922);
nor UO_2228 (O_2228,N_24452,N_24734);
xnor UO_2229 (O_2229,N_24735,N_24653);
and UO_2230 (O_2230,N_24771,N_24669);
nand UO_2231 (O_2231,N_24997,N_24652);
nand UO_2232 (O_2232,N_24658,N_24534);
or UO_2233 (O_2233,N_24724,N_24827);
xor UO_2234 (O_2234,N_24408,N_24557);
xnor UO_2235 (O_2235,N_24960,N_24751);
nand UO_2236 (O_2236,N_24409,N_24563);
xor UO_2237 (O_2237,N_24870,N_24544);
nand UO_2238 (O_2238,N_24637,N_24895);
and UO_2239 (O_2239,N_24400,N_24677);
nor UO_2240 (O_2240,N_24915,N_24999);
and UO_2241 (O_2241,N_24758,N_24884);
nand UO_2242 (O_2242,N_24468,N_24625);
nor UO_2243 (O_2243,N_24945,N_24696);
and UO_2244 (O_2244,N_24461,N_24883);
nor UO_2245 (O_2245,N_24619,N_24389);
or UO_2246 (O_2246,N_24868,N_24502);
nor UO_2247 (O_2247,N_24616,N_24918);
nor UO_2248 (O_2248,N_24996,N_24846);
or UO_2249 (O_2249,N_24661,N_24766);
nor UO_2250 (O_2250,N_24779,N_24669);
or UO_2251 (O_2251,N_24764,N_24571);
xor UO_2252 (O_2252,N_24460,N_24409);
nor UO_2253 (O_2253,N_24437,N_24444);
or UO_2254 (O_2254,N_24627,N_24429);
and UO_2255 (O_2255,N_24415,N_24721);
xnor UO_2256 (O_2256,N_24396,N_24748);
nor UO_2257 (O_2257,N_24721,N_24430);
and UO_2258 (O_2258,N_24917,N_24649);
xor UO_2259 (O_2259,N_24426,N_24645);
xor UO_2260 (O_2260,N_24684,N_24898);
and UO_2261 (O_2261,N_24394,N_24499);
nor UO_2262 (O_2262,N_24504,N_24879);
and UO_2263 (O_2263,N_24607,N_24836);
and UO_2264 (O_2264,N_24987,N_24997);
nand UO_2265 (O_2265,N_24522,N_24896);
or UO_2266 (O_2266,N_24507,N_24850);
xor UO_2267 (O_2267,N_24925,N_24404);
nand UO_2268 (O_2268,N_24785,N_24571);
and UO_2269 (O_2269,N_24515,N_24708);
nor UO_2270 (O_2270,N_24569,N_24963);
or UO_2271 (O_2271,N_24695,N_24830);
and UO_2272 (O_2272,N_24478,N_24724);
nand UO_2273 (O_2273,N_24893,N_24601);
nand UO_2274 (O_2274,N_24874,N_24738);
nand UO_2275 (O_2275,N_24586,N_24436);
nor UO_2276 (O_2276,N_24522,N_24792);
nand UO_2277 (O_2277,N_24916,N_24408);
or UO_2278 (O_2278,N_24648,N_24748);
and UO_2279 (O_2279,N_24841,N_24907);
nand UO_2280 (O_2280,N_24715,N_24985);
nor UO_2281 (O_2281,N_24538,N_24727);
nand UO_2282 (O_2282,N_24525,N_24819);
nor UO_2283 (O_2283,N_24927,N_24968);
nor UO_2284 (O_2284,N_24393,N_24619);
nand UO_2285 (O_2285,N_24947,N_24534);
and UO_2286 (O_2286,N_24699,N_24688);
and UO_2287 (O_2287,N_24451,N_24767);
or UO_2288 (O_2288,N_24495,N_24726);
xnor UO_2289 (O_2289,N_24535,N_24841);
nor UO_2290 (O_2290,N_24753,N_24779);
nand UO_2291 (O_2291,N_24510,N_24416);
and UO_2292 (O_2292,N_24801,N_24724);
xnor UO_2293 (O_2293,N_24684,N_24930);
nor UO_2294 (O_2294,N_24622,N_24860);
nor UO_2295 (O_2295,N_24526,N_24623);
and UO_2296 (O_2296,N_24935,N_24654);
nor UO_2297 (O_2297,N_24551,N_24425);
nand UO_2298 (O_2298,N_24543,N_24768);
or UO_2299 (O_2299,N_24692,N_24993);
and UO_2300 (O_2300,N_24904,N_24963);
nand UO_2301 (O_2301,N_24987,N_24925);
or UO_2302 (O_2302,N_24785,N_24758);
or UO_2303 (O_2303,N_24814,N_24853);
nor UO_2304 (O_2304,N_24482,N_24755);
and UO_2305 (O_2305,N_24375,N_24888);
xnor UO_2306 (O_2306,N_24769,N_24436);
nor UO_2307 (O_2307,N_24605,N_24889);
nand UO_2308 (O_2308,N_24409,N_24508);
nand UO_2309 (O_2309,N_24669,N_24679);
nand UO_2310 (O_2310,N_24515,N_24996);
and UO_2311 (O_2311,N_24984,N_24443);
xnor UO_2312 (O_2312,N_24428,N_24922);
xnor UO_2313 (O_2313,N_24708,N_24881);
xnor UO_2314 (O_2314,N_24945,N_24712);
and UO_2315 (O_2315,N_24917,N_24760);
or UO_2316 (O_2316,N_24444,N_24387);
xor UO_2317 (O_2317,N_24403,N_24588);
xor UO_2318 (O_2318,N_24554,N_24954);
nand UO_2319 (O_2319,N_24849,N_24484);
xor UO_2320 (O_2320,N_24666,N_24770);
nand UO_2321 (O_2321,N_24503,N_24452);
or UO_2322 (O_2322,N_24912,N_24760);
xnor UO_2323 (O_2323,N_24757,N_24868);
nand UO_2324 (O_2324,N_24630,N_24610);
and UO_2325 (O_2325,N_24928,N_24717);
and UO_2326 (O_2326,N_24555,N_24863);
nor UO_2327 (O_2327,N_24566,N_24896);
nor UO_2328 (O_2328,N_24966,N_24644);
and UO_2329 (O_2329,N_24925,N_24453);
nor UO_2330 (O_2330,N_24656,N_24391);
or UO_2331 (O_2331,N_24768,N_24450);
xor UO_2332 (O_2332,N_24576,N_24617);
nor UO_2333 (O_2333,N_24925,N_24412);
nand UO_2334 (O_2334,N_24735,N_24889);
and UO_2335 (O_2335,N_24442,N_24398);
xnor UO_2336 (O_2336,N_24872,N_24417);
xnor UO_2337 (O_2337,N_24558,N_24803);
xor UO_2338 (O_2338,N_24838,N_24665);
or UO_2339 (O_2339,N_24840,N_24668);
nor UO_2340 (O_2340,N_24398,N_24717);
or UO_2341 (O_2341,N_24552,N_24447);
or UO_2342 (O_2342,N_24916,N_24891);
or UO_2343 (O_2343,N_24654,N_24942);
nor UO_2344 (O_2344,N_24653,N_24965);
nand UO_2345 (O_2345,N_24850,N_24460);
or UO_2346 (O_2346,N_24485,N_24689);
and UO_2347 (O_2347,N_24570,N_24914);
nor UO_2348 (O_2348,N_24897,N_24586);
nand UO_2349 (O_2349,N_24996,N_24392);
nand UO_2350 (O_2350,N_24741,N_24789);
nor UO_2351 (O_2351,N_24754,N_24657);
nand UO_2352 (O_2352,N_24792,N_24722);
nor UO_2353 (O_2353,N_24833,N_24945);
nor UO_2354 (O_2354,N_24587,N_24767);
and UO_2355 (O_2355,N_24811,N_24447);
nand UO_2356 (O_2356,N_24767,N_24633);
xor UO_2357 (O_2357,N_24669,N_24416);
xor UO_2358 (O_2358,N_24487,N_24566);
and UO_2359 (O_2359,N_24447,N_24796);
and UO_2360 (O_2360,N_24763,N_24469);
and UO_2361 (O_2361,N_24622,N_24428);
nand UO_2362 (O_2362,N_24475,N_24401);
nor UO_2363 (O_2363,N_24821,N_24667);
and UO_2364 (O_2364,N_24646,N_24440);
nor UO_2365 (O_2365,N_24519,N_24839);
xor UO_2366 (O_2366,N_24440,N_24566);
nand UO_2367 (O_2367,N_24991,N_24641);
nand UO_2368 (O_2368,N_24403,N_24413);
or UO_2369 (O_2369,N_24593,N_24549);
xnor UO_2370 (O_2370,N_24917,N_24586);
and UO_2371 (O_2371,N_24495,N_24876);
xnor UO_2372 (O_2372,N_24860,N_24814);
nor UO_2373 (O_2373,N_24430,N_24570);
nand UO_2374 (O_2374,N_24800,N_24628);
and UO_2375 (O_2375,N_24446,N_24443);
nand UO_2376 (O_2376,N_24440,N_24479);
or UO_2377 (O_2377,N_24512,N_24521);
or UO_2378 (O_2378,N_24690,N_24697);
xnor UO_2379 (O_2379,N_24722,N_24905);
and UO_2380 (O_2380,N_24969,N_24798);
xor UO_2381 (O_2381,N_24731,N_24523);
nand UO_2382 (O_2382,N_24548,N_24533);
nand UO_2383 (O_2383,N_24877,N_24947);
nor UO_2384 (O_2384,N_24679,N_24885);
and UO_2385 (O_2385,N_24394,N_24420);
or UO_2386 (O_2386,N_24847,N_24713);
or UO_2387 (O_2387,N_24420,N_24963);
nand UO_2388 (O_2388,N_24746,N_24954);
xor UO_2389 (O_2389,N_24814,N_24895);
xor UO_2390 (O_2390,N_24655,N_24678);
and UO_2391 (O_2391,N_24950,N_24387);
xor UO_2392 (O_2392,N_24832,N_24392);
nor UO_2393 (O_2393,N_24608,N_24403);
nor UO_2394 (O_2394,N_24904,N_24494);
and UO_2395 (O_2395,N_24858,N_24832);
or UO_2396 (O_2396,N_24521,N_24574);
and UO_2397 (O_2397,N_24677,N_24831);
nand UO_2398 (O_2398,N_24991,N_24694);
or UO_2399 (O_2399,N_24779,N_24658);
nand UO_2400 (O_2400,N_24560,N_24462);
xor UO_2401 (O_2401,N_24900,N_24684);
or UO_2402 (O_2402,N_24506,N_24413);
nand UO_2403 (O_2403,N_24987,N_24658);
and UO_2404 (O_2404,N_24552,N_24612);
nand UO_2405 (O_2405,N_24728,N_24652);
and UO_2406 (O_2406,N_24791,N_24951);
xnor UO_2407 (O_2407,N_24407,N_24849);
xor UO_2408 (O_2408,N_24450,N_24676);
and UO_2409 (O_2409,N_24454,N_24486);
or UO_2410 (O_2410,N_24630,N_24702);
nand UO_2411 (O_2411,N_24690,N_24399);
nor UO_2412 (O_2412,N_24674,N_24395);
nand UO_2413 (O_2413,N_24506,N_24685);
nor UO_2414 (O_2414,N_24896,N_24513);
xnor UO_2415 (O_2415,N_24856,N_24448);
nor UO_2416 (O_2416,N_24965,N_24499);
nor UO_2417 (O_2417,N_24410,N_24638);
or UO_2418 (O_2418,N_24725,N_24877);
xor UO_2419 (O_2419,N_24519,N_24399);
or UO_2420 (O_2420,N_24482,N_24470);
or UO_2421 (O_2421,N_24645,N_24629);
and UO_2422 (O_2422,N_24418,N_24913);
and UO_2423 (O_2423,N_24697,N_24972);
or UO_2424 (O_2424,N_24578,N_24567);
nand UO_2425 (O_2425,N_24866,N_24930);
nand UO_2426 (O_2426,N_24870,N_24768);
nor UO_2427 (O_2427,N_24868,N_24998);
and UO_2428 (O_2428,N_24496,N_24744);
or UO_2429 (O_2429,N_24527,N_24383);
and UO_2430 (O_2430,N_24835,N_24931);
xor UO_2431 (O_2431,N_24919,N_24736);
or UO_2432 (O_2432,N_24502,N_24490);
and UO_2433 (O_2433,N_24560,N_24517);
nand UO_2434 (O_2434,N_24874,N_24745);
nand UO_2435 (O_2435,N_24694,N_24616);
xnor UO_2436 (O_2436,N_24733,N_24861);
xor UO_2437 (O_2437,N_24596,N_24773);
nand UO_2438 (O_2438,N_24978,N_24995);
nor UO_2439 (O_2439,N_24672,N_24851);
nand UO_2440 (O_2440,N_24758,N_24814);
xnor UO_2441 (O_2441,N_24452,N_24471);
nand UO_2442 (O_2442,N_24882,N_24673);
and UO_2443 (O_2443,N_24789,N_24527);
nor UO_2444 (O_2444,N_24521,N_24842);
nand UO_2445 (O_2445,N_24736,N_24564);
xor UO_2446 (O_2446,N_24390,N_24385);
or UO_2447 (O_2447,N_24564,N_24888);
nor UO_2448 (O_2448,N_24642,N_24614);
nand UO_2449 (O_2449,N_24962,N_24821);
xor UO_2450 (O_2450,N_24375,N_24910);
or UO_2451 (O_2451,N_24507,N_24441);
nand UO_2452 (O_2452,N_24723,N_24503);
or UO_2453 (O_2453,N_24714,N_24476);
nand UO_2454 (O_2454,N_24593,N_24539);
xnor UO_2455 (O_2455,N_24510,N_24382);
or UO_2456 (O_2456,N_24551,N_24928);
or UO_2457 (O_2457,N_24995,N_24960);
nand UO_2458 (O_2458,N_24939,N_24746);
nor UO_2459 (O_2459,N_24896,N_24621);
nand UO_2460 (O_2460,N_24706,N_24557);
or UO_2461 (O_2461,N_24539,N_24978);
or UO_2462 (O_2462,N_24535,N_24867);
and UO_2463 (O_2463,N_24775,N_24620);
xnor UO_2464 (O_2464,N_24912,N_24742);
nand UO_2465 (O_2465,N_24490,N_24426);
nor UO_2466 (O_2466,N_24537,N_24529);
nand UO_2467 (O_2467,N_24814,N_24780);
or UO_2468 (O_2468,N_24449,N_24446);
nand UO_2469 (O_2469,N_24668,N_24676);
and UO_2470 (O_2470,N_24612,N_24537);
nor UO_2471 (O_2471,N_24961,N_24727);
or UO_2472 (O_2472,N_24540,N_24463);
and UO_2473 (O_2473,N_24495,N_24638);
nand UO_2474 (O_2474,N_24909,N_24560);
and UO_2475 (O_2475,N_24847,N_24442);
and UO_2476 (O_2476,N_24552,N_24664);
xnor UO_2477 (O_2477,N_24845,N_24677);
xor UO_2478 (O_2478,N_24835,N_24813);
nor UO_2479 (O_2479,N_24530,N_24906);
and UO_2480 (O_2480,N_24641,N_24880);
and UO_2481 (O_2481,N_24488,N_24533);
or UO_2482 (O_2482,N_24901,N_24601);
or UO_2483 (O_2483,N_24917,N_24648);
or UO_2484 (O_2484,N_24900,N_24518);
nand UO_2485 (O_2485,N_24850,N_24961);
nor UO_2486 (O_2486,N_24761,N_24548);
or UO_2487 (O_2487,N_24924,N_24651);
and UO_2488 (O_2488,N_24942,N_24683);
nor UO_2489 (O_2489,N_24475,N_24447);
nor UO_2490 (O_2490,N_24715,N_24417);
nor UO_2491 (O_2491,N_24392,N_24666);
xnor UO_2492 (O_2492,N_24868,N_24656);
or UO_2493 (O_2493,N_24642,N_24856);
and UO_2494 (O_2494,N_24770,N_24653);
nand UO_2495 (O_2495,N_24779,N_24522);
xnor UO_2496 (O_2496,N_24839,N_24968);
nand UO_2497 (O_2497,N_24585,N_24990);
nand UO_2498 (O_2498,N_24770,N_24504);
and UO_2499 (O_2499,N_24665,N_24487);
or UO_2500 (O_2500,N_24964,N_24439);
nand UO_2501 (O_2501,N_24590,N_24829);
and UO_2502 (O_2502,N_24846,N_24880);
and UO_2503 (O_2503,N_24408,N_24960);
or UO_2504 (O_2504,N_24854,N_24764);
and UO_2505 (O_2505,N_24634,N_24730);
and UO_2506 (O_2506,N_24756,N_24588);
nor UO_2507 (O_2507,N_24834,N_24662);
nor UO_2508 (O_2508,N_24641,N_24619);
nand UO_2509 (O_2509,N_24738,N_24680);
or UO_2510 (O_2510,N_24574,N_24912);
and UO_2511 (O_2511,N_24535,N_24836);
nor UO_2512 (O_2512,N_24433,N_24505);
nand UO_2513 (O_2513,N_24598,N_24547);
and UO_2514 (O_2514,N_24376,N_24493);
nand UO_2515 (O_2515,N_24403,N_24945);
nand UO_2516 (O_2516,N_24453,N_24792);
and UO_2517 (O_2517,N_24893,N_24609);
xor UO_2518 (O_2518,N_24522,N_24634);
nand UO_2519 (O_2519,N_24544,N_24561);
nand UO_2520 (O_2520,N_24460,N_24994);
nor UO_2521 (O_2521,N_24786,N_24530);
nand UO_2522 (O_2522,N_24940,N_24640);
nand UO_2523 (O_2523,N_24782,N_24582);
nand UO_2524 (O_2524,N_24516,N_24945);
nor UO_2525 (O_2525,N_24748,N_24697);
nor UO_2526 (O_2526,N_24600,N_24609);
and UO_2527 (O_2527,N_24871,N_24400);
and UO_2528 (O_2528,N_24731,N_24745);
or UO_2529 (O_2529,N_24425,N_24453);
nand UO_2530 (O_2530,N_24668,N_24615);
xnor UO_2531 (O_2531,N_24408,N_24436);
nand UO_2532 (O_2532,N_24764,N_24987);
or UO_2533 (O_2533,N_24399,N_24721);
and UO_2534 (O_2534,N_24962,N_24760);
nand UO_2535 (O_2535,N_24628,N_24587);
nand UO_2536 (O_2536,N_24886,N_24583);
xor UO_2537 (O_2537,N_24837,N_24889);
or UO_2538 (O_2538,N_24386,N_24749);
xor UO_2539 (O_2539,N_24558,N_24694);
xor UO_2540 (O_2540,N_24576,N_24867);
or UO_2541 (O_2541,N_24664,N_24489);
nand UO_2542 (O_2542,N_24775,N_24465);
and UO_2543 (O_2543,N_24559,N_24799);
and UO_2544 (O_2544,N_24862,N_24593);
or UO_2545 (O_2545,N_24821,N_24820);
and UO_2546 (O_2546,N_24742,N_24477);
or UO_2547 (O_2547,N_24499,N_24830);
and UO_2548 (O_2548,N_24561,N_24475);
xor UO_2549 (O_2549,N_24544,N_24862);
and UO_2550 (O_2550,N_24856,N_24742);
or UO_2551 (O_2551,N_24472,N_24925);
and UO_2552 (O_2552,N_24785,N_24894);
nand UO_2553 (O_2553,N_24720,N_24649);
nor UO_2554 (O_2554,N_24466,N_24913);
nor UO_2555 (O_2555,N_24903,N_24380);
nand UO_2556 (O_2556,N_24746,N_24986);
nand UO_2557 (O_2557,N_24987,N_24530);
xnor UO_2558 (O_2558,N_24816,N_24755);
nor UO_2559 (O_2559,N_24674,N_24415);
and UO_2560 (O_2560,N_24699,N_24720);
nor UO_2561 (O_2561,N_24532,N_24552);
xor UO_2562 (O_2562,N_24954,N_24705);
nand UO_2563 (O_2563,N_24502,N_24702);
xor UO_2564 (O_2564,N_24981,N_24614);
xor UO_2565 (O_2565,N_24952,N_24697);
and UO_2566 (O_2566,N_24658,N_24770);
nand UO_2567 (O_2567,N_24473,N_24839);
nand UO_2568 (O_2568,N_24725,N_24568);
nand UO_2569 (O_2569,N_24904,N_24767);
and UO_2570 (O_2570,N_24742,N_24727);
or UO_2571 (O_2571,N_24831,N_24726);
xor UO_2572 (O_2572,N_24927,N_24817);
or UO_2573 (O_2573,N_24631,N_24454);
and UO_2574 (O_2574,N_24514,N_24538);
or UO_2575 (O_2575,N_24891,N_24781);
nor UO_2576 (O_2576,N_24407,N_24961);
nand UO_2577 (O_2577,N_24630,N_24875);
nor UO_2578 (O_2578,N_24551,N_24572);
nand UO_2579 (O_2579,N_24444,N_24798);
xor UO_2580 (O_2580,N_24712,N_24527);
xor UO_2581 (O_2581,N_24653,N_24562);
nor UO_2582 (O_2582,N_24820,N_24395);
nor UO_2583 (O_2583,N_24399,N_24445);
or UO_2584 (O_2584,N_24887,N_24493);
nor UO_2585 (O_2585,N_24865,N_24713);
nor UO_2586 (O_2586,N_24839,N_24463);
or UO_2587 (O_2587,N_24390,N_24576);
nor UO_2588 (O_2588,N_24619,N_24819);
or UO_2589 (O_2589,N_24445,N_24667);
and UO_2590 (O_2590,N_24522,N_24930);
or UO_2591 (O_2591,N_24971,N_24812);
or UO_2592 (O_2592,N_24469,N_24962);
or UO_2593 (O_2593,N_24929,N_24713);
nor UO_2594 (O_2594,N_24393,N_24925);
nand UO_2595 (O_2595,N_24755,N_24634);
or UO_2596 (O_2596,N_24571,N_24830);
nand UO_2597 (O_2597,N_24708,N_24850);
and UO_2598 (O_2598,N_24463,N_24382);
nand UO_2599 (O_2599,N_24775,N_24579);
nand UO_2600 (O_2600,N_24923,N_24517);
xnor UO_2601 (O_2601,N_24709,N_24685);
and UO_2602 (O_2602,N_24845,N_24483);
and UO_2603 (O_2603,N_24651,N_24620);
nor UO_2604 (O_2604,N_24590,N_24526);
nand UO_2605 (O_2605,N_24422,N_24380);
and UO_2606 (O_2606,N_24879,N_24394);
or UO_2607 (O_2607,N_24954,N_24809);
xnor UO_2608 (O_2608,N_24677,N_24423);
xor UO_2609 (O_2609,N_24862,N_24604);
and UO_2610 (O_2610,N_24447,N_24842);
and UO_2611 (O_2611,N_24709,N_24512);
nor UO_2612 (O_2612,N_24836,N_24837);
and UO_2613 (O_2613,N_24815,N_24441);
and UO_2614 (O_2614,N_24777,N_24902);
or UO_2615 (O_2615,N_24891,N_24911);
and UO_2616 (O_2616,N_24927,N_24686);
xor UO_2617 (O_2617,N_24516,N_24656);
and UO_2618 (O_2618,N_24612,N_24930);
nor UO_2619 (O_2619,N_24983,N_24811);
nor UO_2620 (O_2620,N_24901,N_24627);
xor UO_2621 (O_2621,N_24632,N_24785);
nand UO_2622 (O_2622,N_24869,N_24486);
nor UO_2623 (O_2623,N_24629,N_24864);
nor UO_2624 (O_2624,N_24589,N_24419);
and UO_2625 (O_2625,N_24736,N_24683);
xor UO_2626 (O_2626,N_24554,N_24615);
or UO_2627 (O_2627,N_24623,N_24463);
xor UO_2628 (O_2628,N_24565,N_24480);
xor UO_2629 (O_2629,N_24627,N_24997);
xnor UO_2630 (O_2630,N_24411,N_24615);
nor UO_2631 (O_2631,N_24668,N_24563);
and UO_2632 (O_2632,N_24652,N_24978);
nor UO_2633 (O_2633,N_24915,N_24592);
and UO_2634 (O_2634,N_24384,N_24912);
nor UO_2635 (O_2635,N_24434,N_24521);
nor UO_2636 (O_2636,N_24872,N_24601);
xor UO_2637 (O_2637,N_24924,N_24884);
and UO_2638 (O_2638,N_24832,N_24980);
or UO_2639 (O_2639,N_24946,N_24704);
nor UO_2640 (O_2640,N_24438,N_24964);
or UO_2641 (O_2641,N_24979,N_24598);
nand UO_2642 (O_2642,N_24611,N_24493);
nor UO_2643 (O_2643,N_24827,N_24403);
or UO_2644 (O_2644,N_24469,N_24898);
nor UO_2645 (O_2645,N_24435,N_24643);
nor UO_2646 (O_2646,N_24946,N_24589);
or UO_2647 (O_2647,N_24397,N_24547);
or UO_2648 (O_2648,N_24572,N_24682);
xnor UO_2649 (O_2649,N_24483,N_24667);
xnor UO_2650 (O_2650,N_24480,N_24858);
or UO_2651 (O_2651,N_24925,N_24612);
nor UO_2652 (O_2652,N_24445,N_24451);
xor UO_2653 (O_2653,N_24672,N_24567);
nand UO_2654 (O_2654,N_24738,N_24563);
nand UO_2655 (O_2655,N_24724,N_24608);
nor UO_2656 (O_2656,N_24379,N_24722);
nand UO_2657 (O_2657,N_24791,N_24843);
or UO_2658 (O_2658,N_24747,N_24377);
xnor UO_2659 (O_2659,N_24608,N_24490);
nor UO_2660 (O_2660,N_24647,N_24672);
nand UO_2661 (O_2661,N_24743,N_24844);
xor UO_2662 (O_2662,N_24382,N_24777);
xnor UO_2663 (O_2663,N_24922,N_24685);
nand UO_2664 (O_2664,N_24775,N_24402);
nand UO_2665 (O_2665,N_24432,N_24894);
or UO_2666 (O_2666,N_24449,N_24722);
or UO_2667 (O_2667,N_24383,N_24872);
xnor UO_2668 (O_2668,N_24995,N_24788);
nand UO_2669 (O_2669,N_24961,N_24438);
or UO_2670 (O_2670,N_24488,N_24870);
or UO_2671 (O_2671,N_24376,N_24540);
xor UO_2672 (O_2672,N_24502,N_24723);
nand UO_2673 (O_2673,N_24533,N_24832);
and UO_2674 (O_2674,N_24887,N_24873);
xor UO_2675 (O_2675,N_24502,N_24592);
xnor UO_2676 (O_2676,N_24680,N_24755);
or UO_2677 (O_2677,N_24607,N_24915);
or UO_2678 (O_2678,N_24461,N_24770);
xnor UO_2679 (O_2679,N_24939,N_24576);
nor UO_2680 (O_2680,N_24959,N_24838);
nor UO_2681 (O_2681,N_24722,N_24811);
and UO_2682 (O_2682,N_24458,N_24542);
nand UO_2683 (O_2683,N_24741,N_24784);
and UO_2684 (O_2684,N_24461,N_24982);
nor UO_2685 (O_2685,N_24743,N_24820);
xor UO_2686 (O_2686,N_24539,N_24675);
xnor UO_2687 (O_2687,N_24898,N_24782);
and UO_2688 (O_2688,N_24772,N_24947);
or UO_2689 (O_2689,N_24671,N_24843);
and UO_2690 (O_2690,N_24695,N_24410);
and UO_2691 (O_2691,N_24984,N_24985);
xor UO_2692 (O_2692,N_24733,N_24647);
and UO_2693 (O_2693,N_24888,N_24706);
or UO_2694 (O_2694,N_24976,N_24407);
xor UO_2695 (O_2695,N_24497,N_24394);
and UO_2696 (O_2696,N_24682,N_24772);
and UO_2697 (O_2697,N_24531,N_24426);
xor UO_2698 (O_2698,N_24512,N_24950);
nor UO_2699 (O_2699,N_24865,N_24690);
and UO_2700 (O_2700,N_24669,N_24886);
or UO_2701 (O_2701,N_24766,N_24720);
xnor UO_2702 (O_2702,N_24533,N_24628);
nor UO_2703 (O_2703,N_24533,N_24789);
xnor UO_2704 (O_2704,N_24840,N_24858);
or UO_2705 (O_2705,N_24716,N_24965);
nor UO_2706 (O_2706,N_24935,N_24397);
nand UO_2707 (O_2707,N_24947,N_24694);
and UO_2708 (O_2708,N_24783,N_24698);
and UO_2709 (O_2709,N_24895,N_24959);
or UO_2710 (O_2710,N_24550,N_24405);
nand UO_2711 (O_2711,N_24447,N_24881);
xnor UO_2712 (O_2712,N_24419,N_24806);
or UO_2713 (O_2713,N_24655,N_24909);
nand UO_2714 (O_2714,N_24523,N_24793);
nand UO_2715 (O_2715,N_24471,N_24525);
xnor UO_2716 (O_2716,N_24534,N_24581);
and UO_2717 (O_2717,N_24545,N_24971);
and UO_2718 (O_2718,N_24829,N_24697);
xnor UO_2719 (O_2719,N_24668,N_24730);
nand UO_2720 (O_2720,N_24727,N_24761);
xor UO_2721 (O_2721,N_24553,N_24781);
or UO_2722 (O_2722,N_24781,N_24882);
or UO_2723 (O_2723,N_24821,N_24596);
and UO_2724 (O_2724,N_24999,N_24474);
xnor UO_2725 (O_2725,N_24740,N_24697);
nand UO_2726 (O_2726,N_24742,N_24641);
nor UO_2727 (O_2727,N_24555,N_24474);
nor UO_2728 (O_2728,N_24445,N_24861);
xnor UO_2729 (O_2729,N_24777,N_24433);
nor UO_2730 (O_2730,N_24998,N_24535);
and UO_2731 (O_2731,N_24690,N_24534);
and UO_2732 (O_2732,N_24544,N_24962);
xor UO_2733 (O_2733,N_24429,N_24755);
nor UO_2734 (O_2734,N_24703,N_24870);
or UO_2735 (O_2735,N_24720,N_24905);
nor UO_2736 (O_2736,N_24435,N_24473);
xnor UO_2737 (O_2737,N_24944,N_24519);
and UO_2738 (O_2738,N_24486,N_24377);
xnor UO_2739 (O_2739,N_24773,N_24679);
and UO_2740 (O_2740,N_24723,N_24875);
or UO_2741 (O_2741,N_24633,N_24747);
and UO_2742 (O_2742,N_24504,N_24728);
xor UO_2743 (O_2743,N_24879,N_24952);
and UO_2744 (O_2744,N_24415,N_24472);
and UO_2745 (O_2745,N_24495,N_24859);
and UO_2746 (O_2746,N_24705,N_24392);
nand UO_2747 (O_2747,N_24600,N_24516);
nor UO_2748 (O_2748,N_24704,N_24461);
and UO_2749 (O_2749,N_24544,N_24717);
nor UO_2750 (O_2750,N_24651,N_24491);
and UO_2751 (O_2751,N_24620,N_24621);
nand UO_2752 (O_2752,N_24820,N_24664);
nor UO_2753 (O_2753,N_24985,N_24797);
nand UO_2754 (O_2754,N_24996,N_24622);
nand UO_2755 (O_2755,N_24596,N_24715);
nor UO_2756 (O_2756,N_24667,N_24820);
or UO_2757 (O_2757,N_24769,N_24489);
nand UO_2758 (O_2758,N_24798,N_24389);
or UO_2759 (O_2759,N_24767,N_24388);
or UO_2760 (O_2760,N_24901,N_24708);
nand UO_2761 (O_2761,N_24794,N_24984);
or UO_2762 (O_2762,N_24515,N_24750);
xor UO_2763 (O_2763,N_24672,N_24665);
nor UO_2764 (O_2764,N_24574,N_24484);
or UO_2765 (O_2765,N_24679,N_24403);
nand UO_2766 (O_2766,N_24910,N_24504);
xnor UO_2767 (O_2767,N_24572,N_24761);
nor UO_2768 (O_2768,N_24818,N_24931);
xor UO_2769 (O_2769,N_24592,N_24556);
nand UO_2770 (O_2770,N_24380,N_24712);
and UO_2771 (O_2771,N_24912,N_24777);
nor UO_2772 (O_2772,N_24769,N_24421);
nor UO_2773 (O_2773,N_24837,N_24412);
xor UO_2774 (O_2774,N_24964,N_24859);
nor UO_2775 (O_2775,N_24877,N_24576);
nand UO_2776 (O_2776,N_24835,N_24600);
xnor UO_2777 (O_2777,N_24742,N_24461);
and UO_2778 (O_2778,N_24917,N_24746);
and UO_2779 (O_2779,N_24509,N_24815);
nor UO_2780 (O_2780,N_24917,N_24486);
xor UO_2781 (O_2781,N_24879,N_24628);
nor UO_2782 (O_2782,N_24399,N_24596);
or UO_2783 (O_2783,N_24714,N_24721);
nor UO_2784 (O_2784,N_24428,N_24433);
or UO_2785 (O_2785,N_24960,N_24442);
xor UO_2786 (O_2786,N_24818,N_24857);
nand UO_2787 (O_2787,N_24880,N_24973);
xor UO_2788 (O_2788,N_24900,N_24603);
nor UO_2789 (O_2789,N_24830,N_24530);
and UO_2790 (O_2790,N_24573,N_24654);
nor UO_2791 (O_2791,N_24947,N_24733);
or UO_2792 (O_2792,N_24596,N_24451);
and UO_2793 (O_2793,N_24698,N_24971);
xor UO_2794 (O_2794,N_24898,N_24718);
xnor UO_2795 (O_2795,N_24663,N_24558);
nand UO_2796 (O_2796,N_24440,N_24582);
or UO_2797 (O_2797,N_24465,N_24844);
nand UO_2798 (O_2798,N_24387,N_24589);
xor UO_2799 (O_2799,N_24800,N_24910);
nor UO_2800 (O_2800,N_24752,N_24740);
xor UO_2801 (O_2801,N_24667,N_24414);
nor UO_2802 (O_2802,N_24788,N_24660);
nor UO_2803 (O_2803,N_24734,N_24462);
and UO_2804 (O_2804,N_24605,N_24398);
nand UO_2805 (O_2805,N_24973,N_24807);
and UO_2806 (O_2806,N_24567,N_24582);
xnor UO_2807 (O_2807,N_24477,N_24857);
xnor UO_2808 (O_2808,N_24622,N_24488);
xor UO_2809 (O_2809,N_24904,N_24848);
or UO_2810 (O_2810,N_24652,N_24875);
xnor UO_2811 (O_2811,N_24461,N_24955);
nand UO_2812 (O_2812,N_24894,N_24464);
and UO_2813 (O_2813,N_24666,N_24882);
xor UO_2814 (O_2814,N_24932,N_24375);
xnor UO_2815 (O_2815,N_24411,N_24745);
or UO_2816 (O_2816,N_24581,N_24385);
nand UO_2817 (O_2817,N_24949,N_24512);
or UO_2818 (O_2818,N_24974,N_24765);
or UO_2819 (O_2819,N_24939,N_24825);
nand UO_2820 (O_2820,N_24589,N_24722);
nand UO_2821 (O_2821,N_24508,N_24947);
and UO_2822 (O_2822,N_24823,N_24704);
nand UO_2823 (O_2823,N_24751,N_24982);
or UO_2824 (O_2824,N_24976,N_24579);
or UO_2825 (O_2825,N_24624,N_24476);
xnor UO_2826 (O_2826,N_24655,N_24690);
nand UO_2827 (O_2827,N_24758,N_24612);
or UO_2828 (O_2828,N_24842,N_24543);
nand UO_2829 (O_2829,N_24544,N_24710);
xor UO_2830 (O_2830,N_24984,N_24576);
nor UO_2831 (O_2831,N_24716,N_24998);
xnor UO_2832 (O_2832,N_24375,N_24836);
and UO_2833 (O_2833,N_24390,N_24974);
nor UO_2834 (O_2834,N_24512,N_24931);
or UO_2835 (O_2835,N_24748,N_24767);
nor UO_2836 (O_2836,N_24742,N_24778);
xor UO_2837 (O_2837,N_24514,N_24429);
or UO_2838 (O_2838,N_24463,N_24782);
or UO_2839 (O_2839,N_24924,N_24537);
nand UO_2840 (O_2840,N_24983,N_24375);
and UO_2841 (O_2841,N_24732,N_24653);
xnor UO_2842 (O_2842,N_24733,N_24810);
nand UO_2843 (O_2843,N_24587,N_24507);
and UO_2844 (O_2844,N_24744,N_24947);
nor UO_2845 (O_2845,N_24958,N_24598);
xnor UO_2846 (O_2846,N_24670,N_24671);
nor UO_2847 (O_2847,N_24933,N_24654);
nand UO_2848 (O_2848,N_24613,N_24916);
and UO_2849 (O_2849,N_24826,N_24637);
or UO_2850 (O_2850,N_24818,N_24682);
nor UO_2851 (O_2851,N_24377,N_24894);
and UO_2852 (O_2852,N_24826,N_24435);
xor UO_2853 (O_2853,N_24506,N_24697);
or UO_2854 (O_2854,N_24820,N_24934);
and UO_2855 (O_2855,N_24826,N_24413);
nor UO_2856 (O_2856,N_24604,N_24669);
or UO_2857 (O_2857,N_24856,N_24505);
or UO_2858 (O_2858,N_24593,N_24728);
nor UO_2859 (O_2859,N_24708,N_24438);
nor UO_2860 (O_2860,N_24579,N_24642);
or UO_2861 (O_2861,N_24832,N_24835);
and UO_2862 (O_2862,N_24677,N_24974);
and UO_2863 (O_2863,N_24871,N_24957);
xnor UO_2864 (O_2864,N_24581,N_24778);
and UO_2865 (O_2865,N_24813,N_24906);
and UO_2866 (O_2866,N_24387,N_24770);
or UO_2867 (O_2867,N_24909,N_24802);
or UO_2868 (O_2868,N_24950,N_24443);
nor UO_2869 (O_2869,N_24475,N_24552);
and UO_2870 (O_2870,N_24879,N_24671);
and UO_2871 (O_2871,N_24608,N_24794);
xor UO_2872 (O_2872,N_24995,N_24410);
or UO_2873 (O_2873,N_24545,N_24718);
and UO_2874 (O_2874,N_24849,N_24431);
xnor UO_2875 (O_2875,N_24641,N_24885);
or UO_2876 (O_2876,N_24508,N_24871);
xor UO_2877 (O_2877,N_24643,N_24700);
or UO_2878 (O_2878,N_24979,N_24912);
nand UO_2879 (O_2879,N_24877,N_24414);
and UO_2880 (O_2880,N_24655,N_24574);
xor UO_2881 (O_2881,N_24532,N_24946);
nand UO_2882 (O_2882,N_24429,N_24858);
nand UO_2883 (O_2883,N_24834,N_24469);
nand UO_2884 (O_2884,N_24921,N_24758);
nor UO_2885 (O_2885,N_24974,N_24983);
xnor UO_2886 (O_2886,N_24792,N_24766);
and UO_2887 (O_2887,N_24721,N_24482);
xor UO_2888 (O_2888,N_24678,N_24429);
xor UO_2889 (O_2889,N_24509,N_24956);
or UO_2890 (O_2890,N_24667,N_24922);
or UO_2891 (O_2891,N_24505,N_24756);
nand UO_2892 (O_2892,N_24526,N_24882);
xnor UO_2893 (O_2893,N_24858,N_24656);
nor UO_2894 (O_2894,N_24913,N_24796);
nor UO_2895 (O_2895,N_24619,N_24938);
xnor UO_2896 (O_2896,N_24534,N_24940);
nand UO_2897 (O_2897,N_24545,N_24807);
xnor UO_2898 (O_2898,N_24507,N_24926);
nor UO_2899 (O_2899,N_24906,N_24827);
nor UO_2900 (O_2900,N_24852,N_24783);
or UO_2901 (O_2901,N_24828,N_24399);
or UO_2902 (O_2902,N_24760,N_24478);
nor UO_2903 (O_2903,N_24507,N_24473);
or UO_2904 (O_2904,N_24517,N_24751);
nor UO_2905 (O_2905,N_24866,N_24870);
nor UO_2906 (O_2906,N_24425,N_24587);
and UO_2907 (O_2907,N_24882,N_24999);
and UO_2908 (O_2908,N_24396,N_24391);
nor UO_2909 (O_2909,N_24703,N_24625);
xor UO_2910 (O_2910,N_24481,N_24538);
nand UO_2911 (O_2911,N_24764,N_24379);
and UO_2912 (O_2912,N_24887,N_24972);
nand UO_2913 (O_2913,N_24989,N_24426);
nor UO_2914 (O_2914,N_24726,N_24948);
xnor UO_2915 (O_2915,N_24540,N_24459);
or UO_2916 (O_2916,N_24738,N_24438);
and UO_2917 (O_2917,N_24650,N_24440);
nor UO_2918 (O_2918,N_24375,N_24483);
nand UO_2919 (O_2919,N_24928,N_24628);
nor UO_2920 (O_2920,N_24694,N_24630);
and UO_2921 (O_2921,N_24616,N_24901);
nand UO_2922 (O_2922,N_24590,N_24623);
xnor UO_2923 (O_2923,N_24852,N_24474);
nor UO_2924 (O_2924,N_24425,N_24402);
nand UO_2925 (O_2925,N_24655,N_24437);
xnor UO_2926 (O_2926,N_24917,N_24784);
or UO_2927 (O_2927,N_24573,N_24400);
xor UO_2928 (O_2928,N_24578,N_24669);
and UO_2929 (O_2929,N_24454,N_24798);
xor UO_2930 (O_2930,N_24439,N_24988);
or UO_2931 (O_2931,N_24434,N_24395);
nand UO_2932 (O_2932,N_24580,N_24879);
nand UO_2933 (O_2933,N_24413,N_24937);
nand UO_2934 (O_2934,N_24996,N_24792);
nor UO_2935 (O_2935,N_24623,N_24911);
and UO_2936 (O_2936,N_24617,N_24575);
xnor UO_2937 (O_2937,N_24380,N_24886);
nand UO_2938 (O_2938,N_24771,N_24784);
xnor UO_2939 (O_2939,N_24407,N_24731);
and UO_2940 (O_2940,N_24686,N_24408);
nand UO_2941 (O_2941,N_24450,N_24888);
xnor UO_2942 (O_2942,N_24563,N_24648);
nand UO_2943 (O_2943,N_24509,N_24608);
nor UO_2944 (O_2944,N_24839,N_24711);
nand UO_2945 (O_2945,N_24693,N_24499);
nor UO_2946 (O_2946,N_24631,N_24929);
and UO_2947 (O_2947,N_24483,N_24600);
nand UO_2948 (O_2948,N_24941,N_24568);
xor UO_2949 (O_2949,N_24999,N_24804);
nand UO_2950 (O_2950,N_24653,N_24585);
nor UO_2951 (O_2951,N_24387,N_24735);
nand UO_2952 (O_2952,N_24390,N_24513);
xnor UO_2953 (O_2953,N_24983,N_24602);
nor UO_2954 (O_2954,N_24926,N_24962);
nor UO_2955 (O_2955,N_24760,N_24758);
and UO_2956 (O_2956,N_24972,N_24925);
xnor UO_2957 (O_2957,N_24498,N_24417);
or UO_2958 (O_2958,N_24910,N_24384);
nand UO_2959 (O_2959,N_24500,N_24728);
xnor UO_2960 (O_2960,N_24544,N_24953);
or UO_2961 (O_2961,N_24938,N_24904);
xor UO_2962 (O_2962,N_24488,N_24682);
and UO_2963 (O_2963,N_24668,N_24432);
xnor UO_2964 (O_2964,N_24592,N_24403);
nand UO_2965 (O_2965,N_24906,N_24502);
nand UO_2966 (O_2966,N_24548,N_24518);
nand UO_2967 (O_2967,N_24764,N_24375);
or UO_2968 (O_2968,N_24937,N_24575);
and UO_2969 (O_2969,N_24784,N_24580);
nor UO_2970 (O_2970,N_24571,N_24708);
nor UO_2971 (O_2971,N_24592,N_24906);
xnor UO_2972 (O_2972,N_24817,N_24548);
xnor UO_2973 (O_2973,N_24659,N_24979);
xor UO_2974 (O_2974,N_24502,N_24612);
xnor UO_2975 (O_2975,N_24698,N_24614);
or UO_2976 (O_2976,N_24689,N_24775);
nand UO_2977 (O_2977,N_24500,N_24383);
and UO_2978 (O_2978,N_24973,N_24376);
or UO_2979 (O_2979,N_24590,N_24606);
and UO_2980 (O_2980,N_24904,N_24698);
and UO_2981 (O_2981,N_24688,N_24554);
nand UO_2982 (O_2982,N_24431,N_24554);
or UO_2983 (O_2983,N_24868,N_24891);
xnor UO_2984 (O_2984,N_24976,N_24910);
and UO_2985 (O_2985,N_24632,N_24684);
nor UO_2986 (O_2986,N_24622,N_24944);
xor UO_2987 (O_2987,N_24776,N_24405);
nand UO_2988 (O_2988,N_24885,N_24866);
nand UO_2989 (O_2989,N_24630,N_24424);
xor UO_2990 (O_2990,N_24728,N_24797);
and UO_2991 (O_2991,N_24654,N_24621);
nand UO_2992 (O_2992,N_24791,N_24540);
nor UO_2993 (O_2993,N_24891,N_24831);
nor UO_2994 (O_2994,N_24397,N_24632);
and UO_2995 (O_2995,N_24798,N_24558);
or UO_2996 (O_2996,N_24624,N_24750);
and UO_2997 (O_2997,N_24677,N_24653);
and UO_2998 (O_2998,N_24904,N_24520);
or UO_2999 (O_2999,N_24591,N_24496);
endmodule