module basic_2500_25000_3000_10_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nand U0 (N_0,In_869,In_996);
and U1 (N_1,In_1522,In_930);
nor U2 (N_2,In_1310,In_358);
xor U3 (N_3,In_339,In_300);
and U4 (N_4,In_1578,In_695);
xnor U5 (N_5,In_1603,In_879);
and U6 (N_6,In_361,In_1617);
and U7 (N_7,In_373,In_1497);
or U8 (N_8,In_672,In_102);
nor U9 (N_9,In_2346,In_509);
xor U10 (N_10,In_498,In_410);
nand U11 (N_11,In_1303,In_2062);
and U12 (N_12,In_360,In_594);
or U13 (N_13,In_154,In_1656);
nor U14 (N_14,In_1987,In_1835);
nand U15 (N_15,In_602,In_2057);
and U16 (N_16,In_1463,In_2308);
xnor U17 (N_17,In_1168,In_2403);
nor U18 (N_18,In_1169,In_1923);
nor U19 (N_19,In_1081,In_2466);
nor U20 (N_20,In_1045,In_1097);
or U21 (N_21,In_2399,In_124);
or U22 (N_22,In_1745,In_1069);
or U23 (N_23,In_1886,In_1334);
nand U24 (N_24,In_1703,In_1779);
xnor U25 (N_25,In_1063,In_1520);
or U26 (N_26,In_531,In_387);
and U27 (N_27,In_25,In_834);
nor U28 (N_28,In_227,In_1730);
nor U29 (N_29,In_280,In_166);
xnor U30 (N_30,In_2017,In_181);
xor U31 (N_31,In_310,In_61);
nand U32 (N_32,In_1973,In_1751);
nand U33 (N_33,In_1400,In_1856);
xor U34 (N_34,In_1134,In_2342);
nor U35 (N_35,In_887,In_1290);
or U36 (N_36,In_2311,In_2045);
nand U37 (N_37,In_2159,In_27);
and U38 (N_38,In_449,In_1661);
nor U39 (N_39,In_248,In_2186);
nand U40 (N_40,In_1015,In_961);
xor U41 (N_41,In_829,In_2038);
and U42 (N_42,In_1731,In_515);
nor U43 (N_43,In_321,In_1083);
or U44 (N_44,In_109,In_1944);
and U45 (N_45,In_323,In_93);
nor U46 (N_46,In_1061,In_341);
and U47 (N_47,In_344,In_1782);
and U48 (N_48,In_135,In_1472);
or U49 (N_49,In_1786,In_1887);
or U50 (N_50,In_1486,In_2366);
nor U51 (N_51,In_2005,In_1588);
xor U52 (N_52,In_1476,In_616);
nor U53 (N_53,In_612,In_714);
nor U54 (N_54,In_781,In_247);
xnor U55 (N_55,In_2069,In_548);
nand U56 (N_56,In_2206,In_131);
nor U57 (N_57,In_577,In_2445);
or U58 (N_58,In_1021,In_1191);
xnor U59 (N_59,In_1824,In_1874);
xor U60 (N_60,In_1278,In_629);
and U61 (N_61,In_1035,In_653);
nor U62 (N_62,In_10,In_1196);
or U63 (N_63,In_2273,In_290);
or U64 (N_64,In_791,In_1707);
and U65 (N_65,In_1438,In_2245);
and U66 (N_66,In_613,In_841);
or U67 (N_67,In_767,In_1948);
nand U68 (N_68,In_1377,In_2000);
xor U69 (N_69,In_2289,In_2301);
xor U70 (N_70,In_1866,In_719);
xor U71 (N_71,In_306,In_1690);
nand U72 (N_72,In_465,In_2058);
or U73 (N_73,In_1541,In_532);
or U74 (N_74,In_720,In_1820);
nand U75 (N_75,In_660,In_1689);
and U76 (N_76,In_2068,In_1292);
xnor U77 (N_77,In_2156,In_1316);
or U78 (N_78,In_1333,In_412);
and U79 (N_79,In_768,In_876);
nand U80 (N_80,In_1420,In_432);
nand U81 (N_81,In_2034,In_511);
nand U82 (N_82,In_1026,In_1758);
xnor U83 (N_83,In_1324,In_1130);
nor U84 (N_84,In_523,In_426);
xnor U85 (N_85,In_1864,In_2096);
nand U86 (N_86,In_1032,In_1722);
nor U87 (N_87,In_601,In_909);
and U88 (N_88,In_579,In_884);
or U89 (N_89,In_941,In_2182);
and U90 (N_90,In_2386,In_193);
nand U91 (N_91,In_2148,In_152);
nand U92 (N_92,In_1842,In_2398);
nand U93 (N_93,In_2475,In_687);
nor U94 (N_94,In_2,In_1111);
and U95 (N_95,In_1869,In_117);
or U96 (N_96,In_632,In_776);
or U97 (N_97,In_1103,In_1315);
and U98 (N_98,In_2077,In_13);
and U99 (N_99,In_628,In_952);
xnor U100 (N_100,In_1464,In_1589);
nor U101 (N_101,In_1411,In_2056);
or U102 (N_102,In_1900,In_396);
nor U103 (N_103,In_2259,In_526);
or U104 (N_104,In_1117,In_668);
nand U105 (N_105,In_1468,In_67);
xnor U106 (N_106,In_238,In_1633);
nor U107 (N_107,In_2272,In_1955);
and U108 (N_108,In_349,In_984);
nand U109 (N_109,In_1545,In_1488);
nand U110 (N_110,In_5,In_2434);
and U111 (N_111,In_172,In_1637);
or U112 (N_112,In_1296,In_822);
nor U113 (N_113,In_2417,In_1550);
or U114 (N_114,In_419,In_1662);
nand U115 (N_115,In_864,In_529);
xnor U116 (N_116,In_2283,In_987);
or U117 (N_117,In_1154,In_983);
xnor U118 (N_118,In_1294,In_353);
or U119 (N_119,In_902,In_53);
and U120 (N_120,In_1311,In_2185);
nor U121 (N_121,In_492,In_2428);
nor U122 (N_122,In_1428,In_2310);
nand U123 (N_123,In_959,In_922);
and U124 (N_124,In_2369,In_108);
nand U125 (N_125,In_1876,In_1502);
and U126 (N_126,In_1778,In_1006);
or U127 (N_127,In_2339,In_1483);
or U128 (N_128,In_273,In_686);
xnor U129 (N_129,In_2049,In_1408);
and U130 (N_130,In_989,In_2275);
nor U131 (N_131,In_785,In_1052);
nor U132 (N_132,In_76,In_2468);
or U133 (N_133,In_1099,In_1020);
nor U134 (N_134,In_581,In_1905);
or U135 (N_135,In_1078,In_1050);
xnor U136 (N_136,In_596,In_855);
nand U137 (N_137,In_1664,In_2161);
nor U138 (N_138,In_1022,In_1318);
or U139 (N_139,In_1857,In_1110);
and U140 (N_140,In_1638,In_1345);
and U141 (N_141,In_1594,In_372);
nor U142 (N_142,In_267,In_721);
nand U143 (N_143,In_1931,In_1028);
nor U144 (N_144,In_2050,In_1787);
xnor U145 (N_145,In_1821,In_1769);
xor U146 (N_146,In_2480,In_1155);
or U147 (N_147,In_113,In_1434);
nor U148 (N_148,In_404,In_1029);
or U149 (N_149,In_64,In_140);
xnor U150 (N_150,In_2319,In_14);
nand U151 (N_151,In_2157,In_508);
and U152 (N_152,In_26,In_2102);
xnor U153 (N_153,In_1335,In_491);
and U154 (N_154,In_1500,In_593);
and U155 (N_155,In_1806,In_1993);
nor U156 (N_156,In_1659,In_933);
nor U157 (N_157,In_1840,In_843);
nand U158 (N_158,In_467,In_182);
and U159 (N_159,In_132,In_2128);
nor U160 (N_160,In_1912,In_391);
xor U161 (N_161,In_1836,In_2250);
nand U162 (N_162,In_1817,In_1265);
or U163 (N_163,In_47,In_2120);
nand U164 (N_164,In_1425,In_953);
or U165 (N_165,In_106,In_1418);
nor U166 (N_166,In_1366,In_2438);
xor U167 (N_167,In_567,In_728);
and U168 (N_168,In_2484,In_2420);
nand U169 (N_169,In_630,In_545);
nor U170 (N_170,In_2044,In_1627);
xnor U171 (N_171,In_433,In_2370);
nor U172 (N_172,In_1267,In_656);
nor U173 (N_173,In_994,In_2146);
xor U174 (N_174,In_395,In_2177);
and U175 (N_175,In_435,In_201);
or U176 (N_176,In_800,In_3);
nor U177 (N_177,In_572,In_1284);
or U178 (N_178,In_1346,In_2152);
nor U179 (N_179,In_216,In_2201);
nand U180 (N_180,In_2253,In_350);
or U181 (N_181,In_2167,In_1643);
xor U182 (N_182,In_538,In_1381);
or U183 (N_183,In_854,In_2101);
nor U184 (N_184,In_199,In_2293);
or U185 (N_185,In_1775,In_2367);
nor U186 (N_186,In_2383,In_2192);
nor U187 (N_187,In_149,In_1198);
or U188 (N_188,In_425,In_759);
nand U189 (N_189,In_73,In_1270);
or U190 (N_190,In_1357,In_640);
and U191 (N_191,In_1936,In_2224);
nor U192 (N_192,In_928,In_2143);
nor U193 (N_193,In_651,In_303);
and U194 (N_194,In_442,In_1025);
nor U195 (N_195,In_1985,In_705);
and U196 (N_196,In_516,In_1565);
or U197 (N_197,In_1142,In_2204);
or U198 (N_198,In_733,In_1510);
nand U199 (N_199,In_1492,In_2122);
xor U200 (N_200,In_875,In_1162);
xnor U201 (N_201,In_2121,In_48);
nor U202 (N_202,In_1666,In_2215);
nand U203 (N_203,In_145,In_2372);
nand U204 (N_204,In_794,In_220);
nor U205 (N_205,In_1160,In_370);
and U206 (N_206,In_2207,In_696);
xor U207 (N_207,In_1604,In_873);
nor U208 (N_208,In_826,In_211);
and U209 (N_209,In_2309,In_1960);
xor U210 (N_210,In_512,In_1161);
xnor U211 (N_211,In_1060,In_1109);
xnor U212 (N_212,In_1037,In_688);
nor U213 (N_213,In_1048,In_810);
or U214 (N_214,In_877,In_1728);
xor U215 (N_215,In_1555,In_537);
xnor U216 (N_216,In_1808,In_1688);
and U217 (N_217,In_1924,In_1138);
nor U218 (N_218,In_661,In_443);
and U219 (N_219,In_1902,In_1892);
and U220 (N_220,In_926,In_1753);
nand U221 (N_221,In_742,In_2084);
and U222 (N_222,In_2216,In_747);
or U223 (N_223,In_7,In_1450);
xnor U224 (N_224,In_1616,In_481);
and U225 (N_225,In_765,In_2354);
xnor U226 (N_226,In_1564,In_1852);
xor U227 (N_227,In_2375,In_2486);
nand U228 (N_228,In_507,In_1470);
nor U229 (N_229,In_549,In_1071);
nor U230 (N_230,In_1827,In_962);
xor U231 (N_231,In_1772,In_1701);
nor U232 (N_232,In_1274,In_1102);
nor U233 (N_233,In_2035,In_551);
xor U234 (N_234,In_554,In_871);
nand U235 (N_235,In_495,In_1766);
xnor U236 (N_236,In_2287,In_1282);
and U237 (N_237,In_1528,In_459);
nor U238 (N_238,In_223,In_1950);
nand U239 (N_239,In_787,In_725);
nand U240 (N_240,In_753,In_1088);
xnor U241 (N_241,In_1983,In_408);
xor U242 (N_242,In_816,In_1430);
and U243 (N_243,In_1382,In_1040);
nand U244 (N_244,In_0,In_857);
and U245 (N_245,In_423,In_1626);
nand U246 (N_246,In_2088,In_722);
nand U247 (N_247,In_195,In_1585);
nand U248 (N_248,In_2307,In_1937);
nor U249 (N_249,In_775,In_769);
nor U250 (N_250,In_1654,In_1338);
and U251 (N_251,In_148,In_1034);
xnor U252 (N_252,In_853,In_1459);
and U253 (N_253,In_731,In_872);
and U254 (N_254,In_1783,In_649);
or U255 (N_255,In_1790,In_1750);
xnor U256 (N_256,In_1074,In_2411);
xor U257 (N_257,In_215,In_752);
and U258 (N_258,In_729,In_456);
nor U259 (N_259,In_2498,In_1828);
xnor U260 (N_260,In_228,In_944);
and U261 (N_261,In_2297,In_1359);
nand U262 (N_262,In_1653,In_1254);
nand U263 (N_263,In_2104,In_2294);
nand U264 (N_264,In_2132,In_2111);
nor U265 (N_265,In_402,In_1647);
xor U266 (N_266,In_180,In_2391);
or U267 (N_267,In_1066,In_1120);
nor U268 (N_268,In_38,In_1574);
nand U269 (N_269,In_1720,In_1436);
or U270 (N_270,In_50,In_878);
nor U271 (N_271,In_1904,In_700);
xor U272 (N_272,In_1014,In_392);
nor U273 (N_273,In_1737,In_2359);
xor U274 (N_274,In_633,In_2142);
xor U275 (N_275,In_682,In_1628);
nand U276 (N_276,In_2382,In_1132);
nor U277 (N_277,In_207,In_105);
nor U278 (N_278,In_1851,In_1304);
nor U279 (N_279,In_1807,In_107);
nor U280 (N_280,In_689,In_1139);
and U281 (N_281,In_1301,In_2328);
nand U282 (N_282,In_292,In_849);
and U283 (N_283,In_2355,In_1119);
nor U284 (N_284,In_394,In_748);
xnor U285 (N_285,In_803,In_30);
xnor U286 (N_286,In_356,In_1233);
and U287 (N_287,In_1255,In_583);
nand U288 (N_288,In_898,In_244);
or U289 (N_289,In_2336,In_2471);
xor U290 (N_290,In_338,In_539);
nor U291 (N_291,In_643,In_16);
xor U292 (N_292,In_1634,In_1994);
and U293 (N_293,In_204,In_202);
nor U294 (N_294,In_662,In_2011);
xor U295 (N_295,In_1509,In_1477);
nand U296 (N_296,In_2026,In_942);
nand U297 (N_297,In_2223,In_970);
nor U298 (N_298,In_1384,In_1932);
nand U299 (N_299,In_2012,In_1706);
xor U300 (N_300,In_634,In_846);
nand U301 (N_301,In_893,In_2390);
and U302 (N_302,In_190,In_2230);
and U303 (N_303,In_1481,In_19);
nor U304 (N_304,In_1156,In_2335);
nand U305 (N_305,In_226,In_1997);
or U306 (N_306,In_2274,In_276);
nor U307 (N_307,In_165,In_1329);
xor U308 (N_308,In_142,In_990);
or U309 (N_309,In_2353,In_2220);
nor U310 (N_310,In_1496,In_1739);
and U311 (N_311,In_1660,In_1044);
and U312 (N_312,In_403,In_706);
and U313 (N_313,In_351,In_584);
and U314 (N_314,In_1801,In_1249);
nand U315 (N_315,In_1176,In_1457);
xnor U316 (N_316,In_1322,In_1263);
or U317 (N_317,In_1732,In_1018);
or U318 (N_318,In_2254,In_1403);
nor U319 (N_319,In_1406,In_1996);
xor U320 (N_320,In_2109,In_2189);
and U321 (N_321,In_197,In_1979);
and U322 (N_322,In_1184,In_1183);
xor U323 (N_323,In_1893,In_786);
or U324 (N_324,In_694,In_2439);
nand U325 (N_325,In_1646,In_1984);
xor U326 (N_326,In_233,In_897);
nand U327 (N_327,In_1003,In_1552);
or U328 (N_328,In_1221,In_1000);
or U329 (N_329,In_1036,In_1396);
xnor U330 (N_330,In_1543,In_1224);
nor U331 (N_331,In_2315,In_2124);
nor U332 (N_332,In_158,In_1039);
nand U333 (N_333,In_998,In_377);
and U334 (N_334,In_1326,In_1330);
or U335 (N_335,In_938,In_1314);
and U336 (N_336,In_115,In_671);
or U337 (N_337,In_49,In_2350);
or U338 (N_338,In_521,In_122);
or U339 (N_339,In_886,In_141);
nor U340 (N_340,In_737,In_1572);
xor U341 (N_341,In_251,In_525);
nor U342 (N_342,In_1831,In_1587);
nor U343 (N_343,In_2252,In_1651);
and U344 (N_344,In_368,In_2452);
nor U345 (N_345,In_2015,In_1573);
and U346 (N_346,In_792,In_892);
nor U347 (N_347,In_1429,In_451);
xnor U348 (N_348,In_1268,In_2107);
nor U349 (N_349,In_763,In_1070);
nand U350 (N_350,In_272,In_1401);
or U351 (N_351,In_814,In_2208);
nand U352 (N_352,In_2018,In_1173);
nor U353 (N_353,In_609,In_2203);
or U354 (N_354,In_78,In_1388);
or U355 (N_355,In_1352,In_2134);
and U356 (N_356,In_472,In_72);
nor U357 (N_357,In_2174,In_885);
or U358 (N_358,In_607,In_1596);
nor U359 (N_359,In_2173,In_1861);
and U360 (N_360,In_870,In_2340);
or U361 (N_361,In_1291,In_1279);
xor U362 (N_362,In_1741,In_809);
nor U363 (N_363,In_1289,In_1615);
nor U364 (N_364,In_222,In_1792);
nand U365 (N_365,In_191,In_1726);
or U366 (N_366,In_297,In_589);
and U367 (N_367,In_1187,In_421);
nor U368 (N_368,In_482,In_1179);
or U369 (N_369,In_1201,In_1811);
and U370 (N_370,In_995,In_264);
and U371 (N_371,In_1174,In_1131);
nor U372 (N_372,In_179,In_1776);
and U373 (N_373,In_271,In_552);
or U374 (N_374,In_274,In_174);
and U375 (N_375,In_288,In_2071);
nor U376 (N_376,In_417,In_1217);
or U377 (N_377,In_1636,In_1010);
and U378 (N_378,In_1736,In_269);
xnor U379 (N_379,In_1672,In_386);
nor U380 (N_380,In_1079,In_2491);
nand U381 (N_381,In_674,In_1598);
xnor U382 (N_382,In_2488,In_242);
and U383 (N_383,In_1309,In_894);
nand U384 (N_384,In_1523,In_2412);
nand U385 (N_385,In_837,In_2172);
or U386 (N_386,In_17,In_1433);
or U387 (N_387,In_1398,In_278);
nand U388 (N_388,In_390,In_807);
and U389 (N_389,In_1300,In_185);
or U390 (N_390,In_1474,In_831);
nand U391 (N_391,In_452,In_772);
nand U392 (N_392,In_1392,In_1456);
nand U393 (N_393,In_1141,In_1143);
nand U394 (N_394,In_2221,In_836);
nor U395 (N_395,In_947,In_256);
nor U396 (N_396,In_2089,In_1599);
or U397 (N_397,In_1361,In_2037);
nand U398 (N_398,In_2324,In_848);
nand U399 (N_399,In_2269,In_15);
or U400 (N_400,In_200,In_364);
and U401 (N_401,In_503,In_1567);
nand U402 (N_402,In_1729,In_330);
nand U403 (N_403,In_1373,In_1364);
and U404 (N_404,In_441,In_2467);
and U405 (N_405,In_1568,In_980);
or U406 (N_406,In_1675,In_1471);
or U407 (N_407,In_851,In_205);
xor U408 (N_408,In_2461,In_2078);
nand U409 (N_409,In_1992,In_1759);
nand U410 (N_410,In_943,In_1180);
nand U411 (N_411,In_1389,In_1503);
xnor U412 (N_412,In_474,In_192);
or U413 (N_413,In_654,In_988);
nor U414 (N_414,In_868,In_820);
xor U415 (N_415,In_1592,In_744);
nand U416 (N_416,In_240,In_1724);
xnor U417 (N_417,In_1793,In_1687);
nand U418 (N_418,In_289,In_2133);
and U419 (N_419,In_2160,In_2080);
xnor U420 (N_420,In_2075,In_2040);
and U421 (N_421,In_1600,In_2007);
xor U422 (N_422,In_1395,In_1024);
and U423 (N_423,In_119,In_756);
nand U424 (N_424,In_1917,In_2414);
xor U425 (N_425,In_506,In_1883);
and U426 (N_426,In_440,In_1106);
xnor U427 (N_427,In_1645,In_1907);
nor U428 (N_428,In_1487,In_1614);
nor U429 (N_429,In_1941,In_1563);
or U430 (N_430,In_1038,In_1192);
or U431 (N_431,In_576,In_1057);
xor U432 (N_432,In_2257,In_655);
nand U433 (N_433,In_2325,In_85);
or U434 (N_434,In_2415,In_2093);
nor U435 (N_435,In_2406,In_883);
nor U436 (N_436,In_434,In_1721);
nand U437 (N_437,In_1976,In_1605);
nor U438 (N_438,In_1761,In_369);
xnor U439 (N_439,In_1166,In_436);
xor U440 (N_440,In_1974,In_2053);
nand U441 (N_441,In_1723,In_813);
xnor U442 (N_442,In_1190,In_798);
nand U443 (N_443,In_975,In_1575);
nand U444 (N_444,In_2153,In_1073);
xnor U445 (N_445,In_1252,In_2455);
xnor U446 (N_446,In_1505,In_1049);
and U447 (N_447,In_1489,In_2373);
nand U448 (N_448,In_2362,In_1077);
or U449 (N_449,In_1529,In_1952);
nand U450 (N_450,In_1934,In_1409);
nand U451 (N_451,In_1815,In_1966);
or U452 (N_452,In_2384,In_1370);
nor U453 (N_453,In_2169,In_1337);
nand U454 (N_454,In_666,In_1845);
nand U455 (N_455,In_2376,In_2395);
or U456 (N_456,In_281,In_2424);
nor U457 (N_457,In_2258,In_1673);
nand U458 (N_458,In_66,In_2092);
and U459 (N_459,In_736,In_1913);
or U460 (N_460,In_1286,In_856);
or U461 (N_461,In_1989,In_2240);
nor U462 (N_462,In_1964,In_357);
nor U463 (N_463,In_2085,In_1532);
and U464 (N_464,In_951,In_455);
and U465 (N_465,In_665,In_82);
xnor U466 (N_466,In_2267,In_1846);
or U467 (N_467,In_1306,In_912);
xnor U468 (N_468,In_1889,In_1911);
xor U469 (N_469,In_2348,In_1855);
and U470 (N_470,In_1308,In_1242);
nand U471 (N_471,In_555,In_1013);
nand U472 (N_472,In_2227,In_977);
nor U473 (N_473,In_418,In_355);
and U474 (N_474,In_2191,In_218);
or U475 (N_475,In_783,In_1128);
nand U476 (N_476,In_1611,In_1695);
and U477 (N_477,In_2392,In_1449);
nor U478 (N_478,In_401,In_31);
nand U479 (N_479,In_1789,In_2290);
xnor U480 (N_480,In_1865,In_573);
and U481 (N_481,In_279,In_1858);
nand U482 (N_482,In_925,In_1170);
nor U483 (N_483,In_1287,In_949);
nor U484 (N_484,In_1928,In_12);
and U485 (N_485,In_1405,In_914);
or U486 (N_486,In_2377,In_1890);
nand U487 (N_487,In_90,In_493);
or U488 (N_488,In_2113,In_2137);
nor U489 (N_489,In_1546,In_2262);
and U490 (N_490,In_497,In_1098);
xor U491 (N_491,In_1240,In_2260);
or U492 (N_492,In_178,In_1451);
nor U493 (N_493,In_460,In_316);
or U494 (N_494,In_487,In_1946);
or U495 (N_495,In_754,In_1220);
or U496 (N_496,In_1498,In_2371);
xnor U497 (N_497,In_2119,In_778);
xnor U498 (N_498,In_2300,In_1513);
xnor U499 (N_499,In_381,In_830);
and U500 (N_500,In_955,In_684);
nor U501 (N_501,In_1253,In_1348);
nor U502 (N_502,In_2180,In_1453);
or U503 (N_503,In_825,In_692);
nor U504 (N_504,In_934,In_96);
or U505 (N_505,In_2178,In_1704);
xor U506 (N_506,In_2261,In_2014);
xnor U507 (N_507,In_1121,In_863);
and U508 (N_508,In_2465,In_461);
and U509 (N_509,In_2456,In_424);
xnor U510 (N_510,In_563,In_534);
xor U511 (N_511,In_1312,In_1755);
nor U512 (N_512,In_57,In_75);
xnor U513 (N_513,In_1231,In_522);
nand U514 (N_514,In_895,In_478);
or U515 (N_515,In_1631,In_2095);
nand U516 (N_516,In_2442,In_2082);
nand U517 (N_517,In_2090,In_976);
or U518 (N_518,In_1839,In_2433);
xor U519 (N_519,In_1415,In_1264);
or U520 (N_520,In_1484,In_2030);
or U521 (N_521,In_1246,In_77);
or U522 (N_522,In_2114,In_1670);
nand U523 (N_523,In_1908,In_161);
nand U524 (N_524,In_667,In_2422);
or U525 (N_525,In_1927,In_641);
xnor U526 (N_526,In_889,In_1800);
nor U527 (N_527,In_2118,In_1712);
xnor U528 (N_528,In_151,In_1369);
and U529 (N_529,In_348,In_750);
nor U530 (N_530,In_1150,In_1269);
nand U531 (N_531,In_1445,In_1041);
and U532 (N_532,In_544,In_1629);
nor U533 (N_533,In_1482,In_638);
or U534 (N_534,In_237,In_1584);
xor U535 (N_535,In_2276,In_1343);
or U536 (N_536,In_1834,In_2379);
nand U537 (N_537,In_1888,In_1930);
and U538 (N_538,In_1122,In_241);
or U539 (N_539,In_760,In_359);
and U540 (N_540,In_732,In_802);
nand U541 (N_541,In_1347,In_795);
or U542 (N_542,In_1620,In_2234);
nor U543 (N_543,In_1203,In_924);
nor U544 (N_544,In_880,In_1958);
nand U545 (N_545,In_2337,In_1426);
xor U546 (N_546,In_311,In_1208);
or U547 (N_547,In_2016,In_1439);
nand U548 (N_548,In_2318,In_123);
nor U549 (N_549,In_236,In_1404);
or U550 (N_550,In_631,In_1288);
or U551 (N_551,In_1884,In_2304);
or U552 (N_552,In_1794,In_2288);
nor U553 (N_553,In_1458,In_2320);
nor U554 (N_554,In_268,In_2316);
nor U555 (N_555,In_2237,In_301);
or U556 (N_556,In_905,In_917);
nor U557 (N_557,In_378,In_882);
nand U558 (N_558,In_1630,In_1988);
xor U559 (N_559,In_501,In_1681);
and U560 (N_560,In_457,In_2470);
xnor U561 (N_561,In_2451,In_838);
and U562 (N_562,In_1781,In_448);
xnor U563 (N_563,In_39,In_2291);
nor U564 (N_564,In_1495,In_476);
nand U565 (N_565,In_1440,In_1803);
nand U566 (N_566,In_1105,In_1548);
nor U567 (N_567,In_1878,In_1214);
nor U568 (N_568,In_815,In_1277);
and U569 (N_569,In_2212,In_2458);
or U570 (N_570,In_1444,In_1084);
nand U571 (N_571,In_999,In_2219);
nor U572 (N_572,In_285,In_20);
or U573 (N_573,In_1562,In_1914);
and U574 (N_574,In_1788,In_484);
or U575 (N_575,In_1031,In_685);
nand U576 (N_576,In_1257,In_796);
nor U577 (N_577,In_558,In_1746);
and U578 (N_578,In_615,In_2009);
and U579 (N_579,In_134,In_1297);
xnor U580 (N_580,In_1469,In_2426);
or U581 (N_581,In_2404,In_1870);
xnor U582 (N_582,In_2198,In_1918);
xor U583 (N_583,In_1247,In_1579);
xor U584 (N_584,In_2329,In_935);
xor U585 (N_585,In_428,In_717);
xor U586 (N_586,In_2265,In_1027);
and U587 (N_587,In_680,In_1757);
xnor U588 (N_588,In_915,In_806);
nor U589 (N_589,In_991,In_1518);
nor U590 (N_590,In_1982,In_1391);
and U591 (N_591,In_611,In_860);
or U592 (N_592,In_103,In_299);
nand U593 (N_593,In_2231,In_1271);
and U594 (N_594,In_735,In_1260);
or U595 (N_595,In_1877,In_2322);
nor U596 (N_596,In_1602,In_352);
nor U597 (N_597,In_1812,In_439);
or U598 (N_598,In_788,In_2020);
and U599 (N_599,In_133,In_54);
and U600 (N_600,In_295,In_2446);
or U601 (N_601,In_59,In_291);
or U602 (N_602,In_2487,In_125);
nand U603 (N_603,In_1657,In_1671);
nor U604 (N_604,In_407,In_1129);
and U605 (N_605,In_445,In_927);
and U606 (N_606,In_625,In_1205);
xnor U607 (N_607,In_1648,In_691);
xor U608 (N_608,In_1327,In_2247);
nor U609 (N_609,In_950,In_1715);
nor U610 (N_610,In_40,In_104);
nor U611 (N_611,In_600,In_2123);
xor U612 (N_612,In_111,In_1969);
xnor U613 (N_613,In_2479,In_2225);
or U614 (N_614,In_175,In_899);
or U615 (N_615,In_517,In_663);
and U616 (N_616,In_1234,In_1371);
and U617 (N_617,In_2497,In_723);
nand U618 (N_618,In_214,In_1298);
xor U619 (N_619,In_1521,In_245);
and U620 (N_620,In_1698,In_2162);
nand U621 (N_621,In_1228,In_702);
nor U622 (N_622,In_1461,In_405);
nor U623 (N_623,In_130,In_150);
nand U624 (N_624,In_212,In_2388);
and U625 (N_625,In_1962,In_1385);
nor U626 (N_626,In_621,In_2218);
or U627 (N_627,In_159,In_1719);
or U628 (N_628,In_2282,In_2042);
and U629 (N_629,In_1367,In_1076);
and U630 (N_630,In_21,In_1033);
nor U631 (N_631,In_282,In_881);
xor U632 (N_632,In_1171,In_1136);
nor U633 (N_633,In_541,In_1394);
nand U634 (N_634,In_1281,In_1711);
nand U635 (N_635,In_1112,In_1762);
nand U636 (N_636,In_1248,In_56);
or U637 (N_637,In_2469,In_2001);
nor U638 (N_638,In_2457,In_913);
and U639 (N_639,In_1534,In_2485);
or U640 (N_640,In_623,In_1159);
xnor U641 (N_641,In_1780,In_1692);
or U642 (N_642,In_1708,In_755);
nand U643 (N_643,In_1302,In_2495);
and U644 (N_644,In_847,In_1375);
xor U645 (N_645,In_536,In_2063);
or U646 (N_646,In_1624,In_1998);
xnor U647 (N_647,In_1898,In_1251);
xnor U648 (N_648,In_2041,In_206);
and U649 (N_649,In_1770,In_437);
or U650 (N_650,In_1188,In_636);
nor U651 (N_651,In_420,In_530);
and U652 (N_652,In_1530,In_2281);
nand U653 (N_653,In_1847,In_1940);
nor U654 (N_654,In_494,In_726);
xor U655 (N_655,In_1216,In_1691);
nor U656 (N_656,In_1123,In_144);
nand U657 (N_657,In_2277,In_88);
nor U658 (N_658,In_284,In_901);
xor U659 (N_659,In_1319,In_908);
xor U660 (N_660,In_2199,In_2140);
xnor U661 (N_661,In_2387,In_1916);
and U662 (N_662,In_1879,In_2150);
xor U663 (N_663,In_1854,In_693);
or U664 (N_664,In_83,In_198);
nand U665 (N_665,In_2303,In_761);
or U666 (N_666,In_727,In_808);
xnor U667 (N_667,In_642,In_1991);
nor U668 (N_668,In_1305,In_2305);
nand U669 (N_669,In_1199,In_2046);
or U670 (N_670,In_2021,In_1623);
xor U671 (N_671,In_1860,In_382);
nand U672 (N_672,In_2195,In_1957);
nand U673 (N_673,In_2241,In_2421);
nor U674 (N_674,In_1609,In_1213);
xor U675 (N_675,In_136,In_2453);
or U676 (N_676,In_1595,In_920);
nor U677 (N_677,In_698,In_97);
and U678 (N_678,In_1390,In_578);
and U679 (N_679,In_479,In_2222);
xor U680 (N_680,In_1910,In_1089);
xor U681 (N_681,In_932,In_1658);
and U682 (N_682,In_1336,In_213);
or U683 (N_683,In_673,In_1978);
nand U684 (N_684,In_1668,In_1813);
nor U685 (N_685,In_1632,In_707);
nand U686 (N_686,In_160,In_1075);
nor U687 (N_687,In_1683,In_1413);
nand U688 (N_688,In_1140,In_1767);
xor U689 (N_689,In_155,In_1047);
nor U690 (N_690,In_1642,In_1676);
or U691 (N_691,In_1009,In_438);
xnor U692 (N_692,In_287,In_1206);
and U693 (N_693,In_782,In_32);
and U694 (N_694,In_1798,In_724);
nor U695 (N_695,In_1607,In_1921);
nand U696 (N_696,In_637,In_1618);
nor U697 (N_697,In_1432,In_1422);
and U698 (N_698,In_265,In_11);
nor U699 (N_699,In_23,In_547);
xor U700 (N_700,In_2235,In_2345);
nor U701 (N_701,In_690,In_110);
or U702 (N_702,In_2013,In_1397);
nand U703 (N_703,In_966,In_819);
and U704 (N_704,In_1949,In_2449);
and U705 (N_705,In_1591,In_1437);
or U706 (N_706,In_2194,In_1891);
nor U707 (N_707,In_230,In_1072);
and U708 (N_708,In_2149,In_1012);
nand U709 (N_709,In_556,In_1256);
nor U710 (N_710,In_1980,In_780);
nor U711 (N_711,In_1849,In_89);
and U712 (N_712,In_326,In_861);
nor U713 (N_713,In_1118,In_1551);
xor U714 (N_714,In_2279,In_608);
and U715 (N_715,In_2313,In_329);
and U716 (N_716,In_580,In_1922);
and U717 (N_717,In_805,In_804);
or U718 (N_718,In_2130,In_307);
and U719 (N_719,In_1223,In_1531);
nor U720 (N_720,In_712,In_2349);
nand U721 (N_721,In_679,In_1101);
xnor U722 (N_722,In_384,In_1227);
nor U723 (N_723,In_1358,In_2284);
nor U724 (N_724,In_163,In_799);
and U725 (N_725,In_904,In_346);
or U726 (N_726,In_1754,In_367);
nand U727 (N_727,In_2302,In_1621);
nor U728 (N_728,In_327,In_485);
nor U729 (N_729,In_2365,In_1004);
xnor U730 (N_730,In_1011,In_1475);
nand U731 (N_731,In_1442,In_948);
xnor U732 (N_732,In_1734,In_1108);
nor U733 (N_733,In_266,In_960);
nor U734 (N_734,In_147,In_1344);
and U735 (N_735,In_644,In_383);
xor U736 (N_736,In_1895,In_2476);
xor U737 (N_737,In_845,In_1680);
nand U738 (N_738,In_69,In_2147);
and U739 (N_739,In_2083,In_946);
nor U740 (N_740,In_1212,In_1590);
nor U741 (N_741,In_565,In_343);
or U742 (N_742,In_762,In_2246);
xor U743 (N_743,In_463,In_1219);
nand U744 (N_744,In_758,In_1272);
xnor U745 (N_745,In_670,In_337);
or U746 (N_746,In_1321,In_2175);
nand U747 (N_747,In_1756,In_1709);
and U748 (N_748,In_1480,In_1959);
xor U749 (N_749,In_2100,In_1317);
nor U750 (N_750,In_398,In_1519);
and U751 (N_751,In_2179,In_896);
nor U752 (N_752,In_1655,In_1999);
or U753 (N_753,In_1635,In_1717);
or U754 (N_754,In_1593,In_2440);
nor U755 (N_755,In_446,In_2330);
and U756 (N_756,In_553,In_2494);
or U757 (N_757,In_1416,In_2139);
xnor U758 (N_758,In_232,In_1151);
and U759 (N_759,In_1875,In_2165);
or U760 (N_760,In_2437,In_741);
nand U761 (N_761,In_1995,In_890);
xor U762 (N_762,In_1148,In_1115);
or U763 (N_763,In_2205,In_1266);
xnor U764 (N_764,In_1696,In_1819);
or U765 (N_765,In_1938,In_62);
or U766 (N_766,In_2462,In_911);
nand U767 (N_767,In_906,In_2214);
and U768 (N_768,In_1678,In_2483);
or U769 (N_769,In_444,In_2211);
or U770 (N_770,In_2117,In_1862);
and U771 (N_771,In_1055,In_2166);
xor U772 (N_772,In_8,In_711);
xnor U773 (N_773,In_1796,In_1559);
nand U774 (N_774,In_1152,In_2474);
and U775 (N_775,In_1556,In_627);
xnor U776 (N_776,In_305,In_1104);
nand U777 (N_777,In_1501,In_1236);
xor U778 (N_778,In_2429,In_2043);
nand U779 (N_779,In_55,In_399);
or U780 (N_780,In_1981,In_2022);
nor U781 (N_781,In_1059,In_1504);
nor U782 (N_782,In_971,In_2209);
or U783 (N_783,In_1897,In_499);
nor U784 (N_784,In_2202,In_2163);
nand U785 (N_785,In_505,In_588);
nor U786 (N_786,In_2363,In_1951);
nor U787 (N_787,In_294,In_566);
nor U788 (N_788,In_1383,In_1747);
nor U789 (N_789,In_519,In_639);
nand U790 (N_790,In_1417,In_2278);
xnor U791 (N_791,In_1956,In_1163);
or U792 (N_792,In_1525,In_1972);
nand U793 (N_793,In_2447,In_1844);
xor U794 (N_794,In_81,In_749);
or U795 (N_795,In_2423,In_2183);
or U796 (N_796,In_2039,In_1095);
xor U797 (N_797,In_1580,In_683);
and U798 (N_798,In_2292,In_1977);
and U799 (N_799,In_1058,In_319);
nand U800 (N_800,In_2002,In_817);
and U801 (N_801,In_867,In_1393);
and U802 (N_802,In_1524,In_708);
or U803 (N_803,In_2473,In_208);
nand U804 (N_804,In_243,In_2358);
nand U805 (N_805,In_647,In_1885);
nand U806 (N_806,In_1743,In_730);
nor U807 (N_807,In_99,In_2425);
and U808 (N_808,In_98,In_571);
or U809 (N_809,In_225,In_546);
nand U810 (N_810,In_1649,In_2072);
and U811 (N_811,In_1850,In_2158);
nor U812 (N_812,In_1942,In_79);
or U813 (N_813,In_1299,In_1225);
xor U814 (N_814,In_164,In_1560);
xor U815 (N_815,In_1353,In_70);
nand U816 (N_816,In_1053,In_1341);
nand U817 (N_817,In_839,In_2299);
and U818 (N_818,In_2312,In_2338);
and U819 (N_819,In_1181,In_1467);
xnor U820 (N_820,In_1124,In_120);
nor U821 (N_821,In_2444,In_453);
and U822 (N_822,In_176,In_1663);
and U823 (N_823,In_1774,In_1967);
and U824 (N_824,In_2255,In_790);
and U825 (N_825,In_1,In_1410);
and U826 (N_826,In_963,In_1823);
and U827 (N_827,In_751,In_1880);
xor U828 (N_828,In_560,In_622);
and U829 (N_829,In_2419,In_835);
xor U830 (N_830,In_1194,In_2200);
xor U831 (N_831,In_2430,In_833);
and U832 (N_832,In_2187,In_1610);
nand U833 (N_833,In_1705,In_582);
and U834 (N_834,In_557,In_2326);
nor U835 (N_835,In_1016,In_858);
or U836 (N_836,In_513,In_1339);
and U837 (N_837,In_1961,In_1625);
or U838 (N_838,In_1494,In_604);
nand U839 (N_839,In_1280,In_325);
xnor U840 (N_840,In_620,In_1313);
or U841 (N_841,In_1540,In_605);
nor U842 (N_842,In_1046,In_1785);
nor U843 (N_843,In_1064,In_2115);
xor U844 (N_844,In_1873,In_363);
nor U845 (N_845,In_937,In_2496);
xor U846 (N_846,In_929,In_379);
nand U847 (N_847,In_2024,In_1147);
and U848 (N_848,In_993,In_45);
xor U849 (N_849,In_1791,In_597);
nor U850 (N_850,In_112,In_2106);
nand U851 (N_851,In_331,In_2070);
and U852 (N_852,In_2242,In_699);
nor U853 (N_853,In_376,In_1933);
xor U854 (N_854,In_2098,In_183);
and U855 (N_855,In_298,In_1177);
xnor U856 (N_856,In_1340,In_1735);
or U857 (N_857,In_1763,In_253);
and U858 (N_858,In_1536,In_1374);
nand U859 (N_859,In_1975,In_840);
nor U860 (N_860,In_703,In_296);
and U861 (N_861,In_411,In_1107);
nand U862 (N_862,In_261,In_1925);
and U863 (N_863,In_430,In_1909);
or U864 (N_864,In_33,In_1665);
xnor U865 (N_865,In_2493,In_1882);
or U866 (N_866,In_1349,In_1859);
nor U867 (N_867,In_704,In_270);
xor U868 (N_868,In_1554,In_2006);
or U869 (N_869,In_614,In_170);
nand U870 (N_870,In_1512,In_1843);
and U871 (N_871,In_1490,In_945);
or U872 (N_872,In_619,In_1167);
nor U873 (N_873,In_2125,In_1571);
nand U874 (N_874,In_1773,In_309);
nor U875 (N_875,In_1684,In_1583);
and U876 (N_876,In_2145,In_41);
nand U877 (N_877,In_1965,In_1239);
or U878 (N_878,In_1537,In_676);
xnor U879 (N_879,In_1686,In_1215);
xnor U880 (N_880,In_1005,In_2210);
or U881 (N_881,In_801,In_74);
nand U882 (N_882,In_2459,In_1218);
and U883 (N_883,In_2344,In_1853);
nor U884 (N_884,In_1473,In_1896);
nor U885 (N_885,In_2270,In_167);
nor U886 (N_886,In_617,In_1511);
xor U887 (N_887,In_824,In_740);
or U888 (N_888,In_189,In_354);
nor U889 (N_889,In_1829,In_2010);
nand U890 (N_890,In_903,In_1833);
or U891 (N_891,In_1328,In_738);
and U892 (N_892,In_1082,In_2008);
or U893 (N_893,In_2060,In_260);
nand U894 (N_894,In_1986,In_1760);
and U895 (N_895,In_2059,In_648);
nor U896 (N_896,In_1320,In_2317);
nor U897 (N_897,In_1566,In_1507);
xor U898 (N_898,In_489,In_677);
nor U899 (N_899,In_219,In_2331);
xor U900 (N_900,In_2048,In_229);
and U901 (N_901,In_1802,In_2489);
xor U902 (N_902,In_1799,In_789);
nand U903 (N_903,In_2352,In_1085);
xnor U904 (N_904,In_745,In_540);
nor U905 (N_905,In_766,In_811);
nor U906 (N_906,In_978,In_1516);
nand U907 (N_907,In_2170,In_2176);
nand U908 (N_908,In_1929,In_968);
and U909 (N_909,In_2099,In_967);
xnor U910 (N_910,In_1412,In_156);
and U911 (N_911,In_2454,In_1804);
or U912 (N_912,In_598,In_1113);
nand U913 (N_913,In_1158,In_1378);
or U914 (N_914,In_2356,In_2418);
and U915 (N_915,In_2402,In_80);
and U916 (N_916,In_771,In_1460);
nor U917 (N_917,In_1867,In_652);
xor U918 (N_918,In_1332,In_413);
xor U919 (N_919,In_1679,In_645);
xor U920 (N_920,In_1777,In_1365);
nor U921 (N_921,In_777,In_1542);
nand U922 (N_922,In_2236,In_2023);
or U923 (N_923,In_1259,In_1899);
or U924 (N_924,In_6,In_718);
nor U925 (N_925,In_1197,In_2238);
nand U926 (N_926,In_1744,In_2126);
nand U927 (N_927,In_1379,In_2251);
nand U928 (N_928,In_2464,In_259);
and U929 (N_929,In_2393,In_263);
nand U930 (N_930,In_1822,In_2110);
or U931 (N_931,In_770,In_1195);
and U932 (N_932,In_406,In_1479);
or U933 (N_933,In_255,In_2228);
and U934 (N_934,In_2243,In_2019);
or U935 (N_935,In_1448,In_2478);
nor U936 (N_936,In_1019,In_2401);
and U937 (N_937,In_1051,In_454);
nand U938 (N_938,In_956,In_587);
and U939 (N_939,In_2154,In_1126);
nor U940 (N_940,In_664,In_823);
nor U941 (N_941,In_318,In_865);
nand U942 (N_942,In_1508,In_2427);
xnor U943 (N_943,In_187,In_1597);
or U944 (N_944,In_1697,In_592);
xnor U945 (N_945,In_965,In_1752);
and U946 (N_946,In_1211,In_2285);
nand U947 (N_947,In_1462,In_974);
xor U948 (N_948,In_312,In_2264);
nor U949 (N_949,In_678,In_973);
or U950 (N_950,In_1368,In_1086);
or U951 (N_951,In_1443,In_322);
nor U952 (N_952,In_701,In_2378);
and U953 (N_953,In_793,In_972);
xor U954 (N_954,In_1127,In_365);
or U955 (N_955,In_1096,In_342);
nand U956 (N_956,In_866,In_1699);
xor U957 (N_957,In_22,In_535);
nand U958 (N_958,In_469,In_366);
nand U959 (N_959,In_2400,In_2407);
xor U960 (N_960,In_1275,In_1023);
nand U961 (N_961,In_827,In_2054);
nor U962 (N_962,In_1514,In_821);
xor U963 (N_963,In_1091,In_1399);
or U964 (N_964,In_940,In_1466);
nand U965 (N_965,In_328,In_2364);
and U966 (N_966,In_520,In_345);
xnor U967 (N_967,In_1241,In_188);
xnor U968 (N_968,In_2127,In_4);
nor U969 (N_969,In_169,In_2190);
or U970 (N_970,In_340,In_92);
or U971 (N_971,In_2155,In_2248);
nand U972 (N_972,In_477,In_1795);
or U973 (N_973,In_137,In_308);
and U974 (N_974,In_2131,In_2067);
xor U975 (N_975,In_1030,In_2036);
or U976 (N_976,In_1809,In_1295);
nor U977 (N_977,In_1137,In_1674);
and U978 (N_978,In_1435,In_1008);
or U979 (N_979,In_1094,In_1186);
and U980 (N_980,In_1612,In_2472);
or U981 (N_981,In_470,In_335);
nor U982 (N_982,In_1652,In_2066);
and U983 (N_983,In_235,In_1810);
xnor U984 (N_984,In_429,In_332);
or U985 (N_985,In_1165,In_1380);
xnor U986 (N_986,In_1172,In_1446);
nand U987 (N_987,In_504,In_1114);
nand U988 (N_988,In_1553,In_919);
nor U989 (N_989,In_542,In_314);
nand U990 (N_990,In_2394,In_293);
nand U991 (N_991,In_2116,In_1576);
nand U992 (N_992,In_320,In_415);
and U993 (N_993,In_734,In_1100);
or U994 (N_994,In_1407,In_2432);
or U995 (N_995,In_91,In_334);
nor U996 (N_996,In_2443,In_1414);
xor U997 (N_997,In_2296,In_36);
nor U998 (N_998,In_1903,In_1065);
nor U999 (N_999,In_514,In_1331);
nand U1000 (N_1000,In_2396,In_1230);
nor U1001 (N_1001,In_1250,In_1485);
nor U1002 (N_1002,In_1733,In_1387);
or U1003 (N_1003,In_564,In_923);
or U1004 (N_1004,In_1402,In_250);
nand U1005 (N_1005,In_385,In_874);
nor U1006 (N_1006,In_1273,In_715);
or U1007 (N_1007,In_1350,In_209);
or U1008 (N_1008,In_1640,In_2129);
nand U1009 (N_1009,In_1276,In_43);
or U1010 (N_1010,In_203,In_2341);
xor U1011 (N_1011,In_957,In_1954);
nor U1012 (N_1012,In_1149,In_2061);
or U1013 (N_1013,In_431,In_94);
or U1014 (N_1014,In_1185,In_1837);
or U1015 (N_1015,In_1771,In_28);
or U1016 (N_1016,In_1356,In_186);
and U1017 (N_1017,In_336,In_128);
nand U1018 (N_1018,In_568,In_1901);
nor U1019 (N_1019,In_129,In_2405);
and U1020 (N_1020,In_1222,In_986);
or U1021 (N_1021,In_262,In_1558);
or U1022 (N_1022,In_561,In_1764);
and U1023 (N_1023,In_675,In_2413);
nand U1024 (N_1024,In_1202,In_2079);
nor U1025 (N_1025,In_1863,In_2065);
xor U1026 (N_1026,In_669,In_1441);
nor U1027 (N_1027,In_2463,In_2239);
nor U1028 (N_1028,In_812,In_739);
or U1029 (N_1029,In_194,In_650);
or U1030 (N_1030,In_743,In_852);
or U1031 (N_1031,In_380,In_844);
xnor U1032 (N_1032,In_450,In_1641);
nor U1033 (N_1033,In_35,In_2374);
or U1034 (N_1034,In_2051,In_590);
and U1035 (N_1035,In_1007,In_1742);
nand U1036 (N_1036,In_595,In_1238);
or U1037 (N_1037,In_1157,In_86);
or U1038 (N_1038,In_1765,In_985);
and U1039 (N_1039,In_1797,In_2410);
nand U1040 (N_1040,In_606,In_1825);
nor U1041 (N_1041,In_171,In_234);
nand U1042 (N_1042,In_1209,In_657);
nand U1043 (N_1043,In_2333,In_2314);
and U1044 (N_1044,In_1784,In_2441);
nor U1045 (N_1045,In_1805,In_779);
and U1046 (N_1046,In_2361,In_574);
xor U1047 (N_1047,In_1182,In_1832);
or U1048 (N_1048,In_362,In_2492);
xor U1049 (N_1049,In_746,In_2188);
nand U1050 (N_1050,In_510,In_466);
nor U1051 (N_1051,In_1258,In_2029);
nor U1052 (N_1052,In_2031,In_1725);
and U1053 (N_1053,In_954,In_34);
and U1054 (N_1054,In_1325,In_2306);
and U1055 (N_1055,In_1768,In_46);
and U1056 (N_1056,In_1454,In_1561);
xnor U1057 (N_1057,In_2171,In_168);
and U1058 (N_1058,In_1354,In_2087);
xnor U1059 (N_1059,In_939,In_979);
xnor U1060 (N_1060,In_1714,In_1478);
and U1061 (N_1061,In_2323,In_1421);
nor U1062 (N_1062,In_1677,In_2408);
or U1063 (N_1063,In_1718,In_1153);
nand U1064 (N_1064,In_784,In_1748);
nand U1065 (N_1065,In_2450,In_1054);
and U1066 (N_1066,In_1342,In_2108);
or U1067 (N_1067,In_1068,In_2081);
xor U1068 (N_1068,In_570,In_1990);
xor U1069 (N_1069,In_63,In_2064);
xor U1070 (N_1070,In_126,In_2028);
nand U1071 (N_1071,In_315,In_2347);
and U1072 (N_1072,In_1926,In_1816);
nor U1073 (N_1073,In_1920,In_275);
and U1074 (N_1074,In_709,In_374);
nand U1075 (N_1075,In_1818,In_1915);
or U1076 (N_1076,In_1515,In_231);
and U1077 (N_1077,In_1146,In_500);
nand U1078 (N_1078,In_2249,In_2168);
xor U1079 (N_1079,In_1133,In_2321);
nand U1080 (N_1080,In_1947,In_162);
or U1081 (N_1081,In_610,In_1539);
nand U1082 (N_1082,In_862,In_842);
and U1083 (N_1083,In_1738,In_2032);
and U1084 (N_1084,In_1526,In_496);
nand U1085 (N_1085,In_1067,In_464);
nand U1086 (N_1086,In_100,In_116);
or U1087 (N_1087,In_254,In_585);
nand U1088 (N_1088,In_1549,In_1193);
xor U1089 (N_1089,In_1178,In_1943);
xnor U1090 (N_1090,In_2141,In_1606);
or U1091 (N_1091,In_2226,In_1538);
or U1092 (N_1092,In_1970,In_527);
xnor U1093 (N_1093,In_1939,In_2193);
or U1094 (N_1094,In_1307,In_143);
and U1095 (N_1095,In_1639,In_393);
nand U1096 (N_1096,In_1881,In_483);
nand U1097 (N_1097,In_1830,In_177);
xor U1098 (N_1098,In_716,In_2298);
or U1099 (N_1099,In_101,In_1569);
or U1100 (N_1100,In_486,In_524);
nor U1101 (N_1101,In_1713,In_562);
xor U1102 (N_1102,In_2112,In_71);
nor U1103 (N_1103,In_1650,In_1144);
nor U1104 (N_1104,In_246,In_1963);
or U1105 (N_1105,In_1694,In_1868);
or U1106 (N_1106,In_1544,In_2135);
nor U1107 (N_1107,In_2380,In_1740);
and U1108 (N_1108,In_221,In_1581);
and U1109 (N_1109,In_1669,In_528);
xor U1110 (N_1110,In_2073,In_1042);
or U1111 (N_1111,In_2263,In_2385);
nor U1112 (N_1112,In_422,In_1285);
xor U1113 (N_1113,In_1894,In_2244);
nand U1114 (N_1114,In_2448,In_1577);
nor U1115 (N_1115,In_1043,In_958);
and U1116 (N_1116,In_51,In_68);
and U1117 (N_1117,In_2389,In_2105);
and U1118 (N_1118,In_1175,In_1355);
nand U1119 (N_1119,In_2136,In_603);
nand U1120 (N_1120,In_347,In_1090);
xor U1121 (N_1121,In_1535,In_2271);
xor U1122 (N_1122,In_184,In_773);
or U1123 (N_1123,In_375,In_1244);
xor U1124 (N_1124,In_797,In_1235);
nor U1125 (N_1125,In_121,In_981);
nand U1126 (N_1126,In_1919,In_52);
and U1127 (N_1127,In_2233,In_458);
nand U1128 (N_1128,In_1547,In_757);
nand U1129 (N_1129,In_774,In_1557);
and U1130 (N_1130,In_2334,In_543);
xnor U1131 (N_1131,In_1749,In_1351);
nand U1132 (N_1132,In_1693,In_916);
nor U1133 (N_1133,In_646,In_969);
or U1134 (N_1134,In_2435,In_1189);
nand U1135 (N_1135,In_2229,In_157);
nand U1136 (N_1136,In_1491,In_2094);
nor U1137 (N_1137,In_58,In_87);
nor U1138 (N_1138,In_710,In_1871);
xor U1139 (N_1139,In_490,In_389);
or U1140 (N_1140,In_1814,In_828);
nor U1141 (N_1141,In_138,In_2004);
nand U1142 (N_1142,In_2025,In_888);
or U1143 (N_1143,In_2213,In_1533);
xnor U1144 (N_1144,In_1493,In_2368);
and U1145 (N_1145,In_146,In_2003);
and U1146 (N_1146,In_1586,In_1427);
or U1147 (N_1147,In_1360,In_324);
nor U1148 (N_1148,In_891,In_2266);
nor U1149 (N_1149,In_2184,In_1622);
nor U1150 (N_1150,In_2477,In_1710);
xor U1151 (N_1151,In_2256,In_468);
nand U1152 (N_1152,In_2332,In_400);
and U1153 (N_1153,In_1506,In_60);
and U1154 (N_1154,In_2181,In_910);
nand U1155 (N_1155,In_992,In_1226);
xnor U1156 (N_1156,In_2280,In_850);
nor U1157 (N_1157,In_1423,In_1447);
or U1158 (N_1158,In_44,In_1431);
nand U1159 (N_1159,In_2197,In_1125);
and U1160 (N_1160,In_818,In_1465);
nor U1161 (N_1161,In_313,In_409);
xnor U1162 (N_1162,In_210,In_2097);
xnor U1163 (N_1163,In_153,In_388);
and U1164 (N_1164,In_1372,In_1953);
or U1165 (N_1165,In_286,In_559);
nand U1166 (N_1166,In_2086,In_2397);
or U1167 (N_1167,In_1229,In_2103);
xnor U1168 (N_1168,In_2357,In_9);
xnor U1169 (N_1169,In_1283,In_1232);
nand U1170 (N_1170,In_2091,In_1261);
nand U1171 (N_1171,In_1838,In_224);
or U1172 (N_1172,In_42,In_95);
nand U1173 (N_1173,In_2164,In_127);
or U1174 (N_1174,In_2151,In_713);
nor U1175 (N_1175,In_626,In_1608);
xor U1176 (N_1176,In_302,In_1092);
xor U1177 (N_1177,In_473,In_1062);
nand U1178 (N_1178,In_1945,In_624);
or U1179 (N_1179,In_277,In_982);
nand U1180 (N_1180,In_480,In_1002);
xnor U1181 (N_1181,In_1362,In_37);
nor U1182 (N_1182,In_139,In_936);
xnor U1183 (N_1183,In_964,In_2055);
xnor U1184 (N_1184,In_1056,In_1164);
nand U1185 (N_1185,In_2286,In_2431);
or U1186 (N_1186,In_252,In_764);
xnor U1187 (N_1187,In_317,In_2436);
nor U1188 (N_1188,In_1716,In_471);
nor U1189 (N_1189,In_599,In_416);
nor U1190 (N_1190,In_569,In_1017);
xnor U1191 (N_1191,In_1848,In_1700);
nor U1192 (N_1192,In_427,In_2416);
and U1193 (N_1193,In_635,In_1455);
xnor U1194 (N_1194,In_2351,In_1376);
nand U1195 (N_1195,In_1872,In_239);
nand U1196 (N_1196,In_1424,In_304);
or U1197 (N_1197,In_1906,In_2490);
or U1198 (N_1198,In_2268,In_2295);
xnor U1199 (N_1199,In_196,In_18);
or U1200 (N_1200,In_1001,In_1087);
and U1201 (N_1201,In_1527,In_2343);
nor U1202 (N_1202,In_1702,In_533);
xor U1203 (N_1203,In_1582,In_29);
and U1204 (N_1204,In_1204,In_832);
xnor U1205 (N_1205,In_488,In_1971);
and U1206 (N_1206,In_1145,In_258);
nand U1207 (N_1207,In_697,In_2074);
or U1208 (N_1208,In_2047,In_2409);
or U1209 (N_1209,In_1116,In_1323);
xor U1210 (N_1210,In_2144,In_1093);
or U1211 (N_1211,In_2217,In_2196);
xor U1212 (N_1212,In_1613,In_1210);
nand U1213 (N_1213,In_575,In_173);
and U1214 (N_1214,In_907,In_2232);
or U1215 (N_1215,In_1826,In_371);
xnor U1216 (N_1216,In_1452,In_550);
or U1217 (N_1217,In_918,In_333);
or U1218 (N_1218,In_1619,In_257);
xnor U1219 (N_1219,In_1685,In_1363);
or U1220 (N_1220,In_1667,In_1682);
nor U1221 (N_1221,In_591,In_658);
and U1222 (N_1222,In_2027,In_2138);
nor U1223 (N_1223,In_518,In_1499);
and U1224 (N_1224,In_1935,In_921);
nor U1225 (N_1225,In_84,In_2360);
nor U1226 (N_1226,In_1245,In_1200);
nor U1227 (N_1227,In_414,In_2481);
nand U1228 (N_1228,In_397,In_1135);
nor U1229 (N_1229,In_1968,In_114);
nand U1230 (N_1230,In_586,In_1570);
xor U1231 (N_1231,In_618,In_859);
or U1232 (N_1232,In_997,In_462);
and U1233 (N_1233,In_118,In_2076);
and U1234 (N_1234,In_2499,In_931);
or U1235 (N_1235,In_217,In_1601);
xor U1236 (N_1236,In_1419,In_1237);
xnor U1237 (N_1237,In_1080,In_1727);
nor U1238 (N_1238,In_283,In_2052);
nor U1239 (N_1239,In_2033,In_502);
nand U1240 (N_1240,In_1386,In_681);
nor U1241 (N_1241,In_65,In_475);
xnor U1242 (N_1242,In_1207,In_1517);
and U1243 (N_1243,In_2381,In_659);
and U1244 (N_1244,In_24,In_2482);
or U1245 (N_1245,In_900,In_2460);
xnor U1246 (N_1246,In_1644,In_1262);
nor U1247 (N_1247,In_2327,In_1293);
nand U1248 (N_1248,In_249,In_447);
nand U1249 (N_1249,In_1243,In_1841);
or U1250 (N_1250,In_477,In_2239);
nand U1251 (N_1251,In_60,In_2495);
or U1252 (N_1252,In_1929,In_1773);
nand U1253 (N_1253,In_1614,In_1590);
nor U1254 (N_1254,In_21,In_2199);
or U1255 (N_1255,In_335,In_2444);
or U1256 (N_1256,In_170,In_1004);
xnor U1257 (N_1257,In_1381,In_2349);
or U1258 (N_1258,In_700,In_2032);
xnor U1259 (N_1259,In_397,In_840);
xnor U1260 (N_1260,In_2333,In_1922);
nand U1261 (N_1261,In_1061,In_342);
nor U1262 (N_1262,In_2349,In_623);
and U1263 (N_1263,In_1088,In_1896);
or U1264 (N_1264,In_2191,In_1493);
and U1265 (N_1265,In_777,In_2367);
or U1266 (N_1266,In_1037,In_180);
nand U1267 (N_1267,In_1174,In_492);
xnor U1268 (N_1268,In_1660,In_1364);
nand U1269 (N_1269,In_182,In_1674);
or U1270 (N_1270,In_1139,In_214);
and U1271 (N_1271,In_1798,In_1849);
nor U1272 (N_1272,In_1811,In_278);
xor U1273 (N_1273,In_303,In_2079);
nor U1274 (N_1274,In_1897,In_839);
xnor U1275 (N_1275,In_699,In_2225);
or U1276 (N_1276,In_281,In_736);
nand U1277 (N_1277,In_1370,In_1212);
or U1278 (N_1278,In_1401,In_115);
xnor U1279 (N_1279,In_1114,In_881);
and U1280 (N_1280,In_1102,In_1818);
or U1281 (N_1281,In_455,In_429);
xnor U1282 (N_1282,In_1310,In_2368);
nand U1283 (N_1283,In_830,In_471);
nand U1284 (N_1284,In_572,In_356);
xnor U1285 (N_1285,In_505,In_158);
xor U1286 (N_1286,In_106,In_245);
nand U1287 (N_1287,In_873,In_2229);
nand U1288 (N_1288,In_1291,In_1876);
nor U1289 (N_1289,In_329,In_1152);
xnor U1290 (N_1290,In_1051,In_292);
and U1291 (N_1291,In_1703,In_482);
nand U1292 (N_1292,In_136,In_2496);
nor U1293 (N_1293,In_1797,In_1417);
nand U1294 (N_1294,In_112,In_205);
nor U1295 (N_1295,In_1416,In_34);
nor U1296 (N_1296,In_2003,In_1547);
and U1297 (N_1297,In_158,In_1944);
xnor U1298 (N_1298,In_2023,In_647);
nor U1299 (N_1299,In_1509,In_2350);
or U1300 (N_1300,In_1980,In_582);
nor U1301 (N_1301,In_1177,In_1373);
xnor U1302 (N_1302,In_1223,In_437);
nand U1303 (N_1303,In_422,In_2071);
nand U1304 (N_1304,In_1860,In_1044);
nor U1305 (N_1305,In_913,In_523);
xor U1306 (N_1306,In_932,In_440);
and U1307 (N_1307,In_1316,In_2107);
nand U1308 (N_1308,In_1816,In_838);
nor U1309 (N_1309,In_367,In_1814);
or U1310 (N_1310,In_2030,In_1905);
nor U1311 (N_1311,In_993,In_1048);
nand U1312 (N_1312,In_1711,In_1036);
nor U1313 (N_1313,In_202,In_829);
or U1314 (N_1314,In_1239,In_351);
or U1315 (N_1315,In_323,In_1732);
nor U1316 (N_1316,In_2272,In_1807);
nand U1317 (N_1317,In_123,In_2379);
nor U1318 (N_1318,In_2198,In_1252);
xnor U1319 (N_1319,In_959,In_1390);
and U1320 (N_1320,In_2219,In_791);
nor U1321 (N_1321,In_1772,In_2350);
and U1322 (N_1322,In_1370,In_944);
nand U1323 (N_1323,In_1695,In_1425);
or U1324 (N_1324,In_2443,In_2403);
nor U1325 (N_1325,In_2288,In_1043);
or U1326 (N_1326,In_272,In_1923);
and U1327 (N_1327,In_1574,In_2025);
nand U1328 (N_1328,In_704,In_631);
nor U1329 (N_1329,In_56,In_2431);
xnor U1330 (N_1330,In_17,In_1024);
and U1331 (N_1331,In_91,In_85);
nand U1332 (N_1332,In_1076,In_1291);
nor U1333 (N_1333,In_1970,In_382);
xor U1334 (N_1334,In_921,In_36);
xor U1335 (N_1335,In_1416,In_725);
nand U1336 (N_1336,In_564,In_207);
nor U1337 (N_1337,In_428,In_1175);
and U1338 (N_1338,In_1991,In_1427);
and U1339 (N_1339,In_301,In_1628);
nand U1340 (N_1340,In_947,In_726);
and U1341 (N_1341,In_755,In_1752);
or U1342 (N_1342,In_978,In_1560);
nand U1343 (N_1343,In_1323,In_1894);
nor U1344 (N_1344,In_261,In_1863);
xnor U1345 (N_1345,In_1859,In_2286);
xnor U1346 (N_1346,In_1296,In_1179);
and U1347 (N_1347,In_2177,In_995);
xnor U1348 (N_1348,In_280,In_2034);
nand U1349 (N_1349,In_1218,In_1560);
nand U1350 (N_1350,In_502,In_832);
xnor U1351 (N_1351,In_351,In_666);
or U1352 (N_1352,In_12,In_1571);
and U1353 (N_1353,In_2341,In_983);
nand U1354 (N_1354,In_327,In_825);
xnor U1355 (N_1355,In_987,In_1753);
or U1356 (N_1356,In_710,In_1728);
or U1357 (N_1357,In_1566,In_2245);
nand U1358 (N_1358,In_2130,In_2471);
xor U1359 (N_1359,In_309,In_1411);
nor U1360 (N_1360,In_1840,In_715);
or U1361 (N_1361,In_809,In_1940);
or U1362 (N_1362,In_1979,In_1095);
nor U1363 (N_1363,In_516,In_873);
nor U1364 (N_1364,In_1653,In_20);
or U1365 (N_1365,In_603,In_312);
nand U1366 (N_1366,In_2005,In_1794);
and U1367 (N_1367,In_133,In_1118);
or U1368 (N_1368,In_1968,In_18);
and U1369 (N_1369,In_967,In_1807);
xor U1370 (N_1370,In_2277,In_1828);
or U1371 (N_1371,In_1898,In_448);
and U1372 (N_1372,In_2003,In_1820);
nand U1373 (N_1373,In_2053,In_440);
nor U1374 (N_1374,In_627,In_1780);
xnor U1375 (N_1375,In_828,In_1096);
nor U1376 (N_1376,In_1199,In_722);
or U1377 (N_1377,In_1218,In_608);
or U1378 (N_1378,In_2362,In_569);
or U1379 (N_1379,In_1389,In_1854);
xor U1380 (N_1380,In_1380,In_792);
nand U1381 (N_1381,In_2325,In_1854);
xnor U1382 (N_1382,In_809,In_2486);
xnor U1383 (N_1383,In_1958,In_2395);
xnor U1384 (N_1384,In_1321,In_2478);
nor U1385 (N_1385,In_2222,In_2014);
nor U1386 (N_1386,In_833,In_2126);
or U1387 (N_1387,In_2135,In_1005);
and U1388 (N_1388,In_1093,In_2453);
nand U1389 (N_1389,In_232,In_1348);
xnor U1390 (N_1390,In_1816,In_1124);
and U1391 (N_1391,In_193,In_178);
nor U1392 (N_1392,In_1673,In_797);
nand U1393 (N_1393,In_998,In_210);
and U1394 (N_1394,In_42,In_1406);
nor U1395 (N_1395,In_1999,In_1493);
xnor U1396 (N_1396,In_820,In_1843);
and U1397 (N_1397,In_1206,In_1409);
nand U1398 (N_1398,In_2239,In_363);
nand U1399 (N_1399,In_345,In_237);
or U1400 (N_1400,In_2159,In_2086);
or U1401 (N_1401,In_1953,In_1430);
nand U1402 (N_1402,In_327,In_1379);
xnor U1403 (N_1403,In_1263,In_92);
nand U1404 (N_1404,In_1445,In_1477);
nand U1405 (N_1405,In_374,In_318);
and U1406 (N_1406,In_427,In_1561);
nor U1407 (N_1407,In_530,In_1895);
nor U1408 (N_1408,In_479,In_1902);
or U1409 (N_1409,In_2293,In_706);
nand U1410 (N_1410,In_2285,In_2298);
nand U1411 (N_1411,In_1001,In_1290);
xnor U1412 (N_1412,In_373,In_1962);
nand U1413 (N_1413,In_1,In_285);
xor U1414 (N_1414,In_2499,In_1822);
nand U1415 (N_1415,In_464,In_1503);
nand U1416 (N_1416,In_1583,In_423);
nor U1417 (N_1417,In_756,In_1075);
xnor U1418 (N_1418,In_638,In_694);
or U1419 (N_1419,In_165,In_2458);
nor U1420 (N_1420,In_2358,In_397);
and U1421 (N_1421,In_315,In_1468);
and U1422 (N_1422,In_1176,In_633);
or U1423 (N_1423,In_117,In_1057);
nand U1424 (N_1424,In_511,In_327);
nand U1425 (N_1425,In_1875,In_1346);
nand U1426 (N_1426,In_1434,In_776);
and U1427 (N_1427,In_1244,In_1839);
nand U1428 (N_1428,In_77,In_583);
nand U1429 (N_1429,In_1256,In_379);
nor U1430 (N_1430,In_1333,In_775);
or U1431 (N_1431,In_1174,In_2296);
xor U1432 (N_1432,In_1965,In_40);
nor U1433 (N_1433,In_2093,In_537);
nor U1434 (N_1434,In_838,In_963);
and U1435 (N_1435,In_1843,In_419);
or U1436 (N_1436,In_493,In_1351);
and U1437 (N_1437,In_605,In_494);
or U1438 (N_1438,In_2346,In_1190);
nor U1439 (N_1439,In_1779,In_1785);
nor U1440 (N_1440,In_1990,In_708);
and U1441 (N_1441,In_1466,In_217);
nand U1442 (N_1442,In_1184,In_1607);
nand U1443 (N_1443,In_1223,In_842);
and U1444 (N_1444,In_702,In_1467);
or U1445 (N_1445,In_186,In_1195);
nand U1446 (N_1446,In_2011,In_1738);
and U1447 (N_1447,In_1249,In_1948);
xor U1448 (N_1448,In_1894,In_315);
xor U1449 (N_1449,In_2076,In_50);
xnor U1450 (N_1450,In_2324,In_1656);
xor U1451 (N_1451,In_23,In_2088);
nand U1452 (N_1452,In_205,In_1441);
or U1453 (N_1453,In_2451,In_2135);
or U1454 (N_1454,In_492,In_931);
and U1455 (N_1455,In_933,In_276);
and U1456 (N_1456,In_1378,In_806);
nand U1457 (N_1457,In_2151,In_2491);
nand U1458 (N_1458,In_1864,In_1775);
nor U1459 (N_1459,In_66,In_1457);
and U1460 (N_1460,In_103,In_723);
or U1461 (N_1461,In_2248,In_1964);
or U1462 (N_1462,In_128,In_2488);
nand U1463 (N_1463,In_1747,In_409);
xor U1464 (N_1464,In_390,In_2215);
and U1465 (N_1465,In_1189,In_2268);
xnor U1466 (N_1466,In_1248,In_888);
and U1467 (N_1467,In_1797,In_100);
xnor U1468 (N_1468,In_1663,In_1045);
nor U1469 (N_1469,In_644,In_683);
xor U1470 (N_1470,In_2283,In_2401);
or U1471 (N_1471,In_406,In_1823);
or U1472 (N_1472,In_1953,In_809);
nand U1473 (N_1473,In_2351,In_2143);
xnor U1474 (N_1474,In_862,In_1521);
and U1475 (N_1475,In_406,In_1139);
and U1476 (N_1476,In_2280,In_2483);
xor U1477 (N_1477,In_2336,In_603);
nor U1478 (N_1478,In_183,In_25);
nand U1479 (N_1479,In_2050,In_1861);
nand U1480 (N_1480,In_1638,In_1645);
or U1481 (N_1481,In_967,In_554);
or U1482 (N_1482,In_527,In_13);
nand U1483 (N_1483,In_1639,In_5);
and U1484 (N_1484,In_1873,In_2101);
nand U1485 (N_1485,In_1414,In_2341);
and U1486 (N_1486,In_787,In_1235);
or U1487 (N_1487,In_2277,In_1028);
or U1488 (N_1488,In_281,In_581);
nand U1489 (N_1489,In_2093,In_1571);
and U1490 (N_1490,In_1243,In_1213);
and U1491 (N_1491,In_667,In_292);
xor U1492 (N_1492,In_840,In_1266);
or U1493 (N_1493,In_2365,In_1208);
nand U1494 (N_1494,In_471,In_517);
xnor U1495 (N_1495,In_346,In_2290);
or U1496 (N_1496,In_571,In_2264);
nand U1497 (N_1497,In_1996,In_2105);
nor U1498 (N_1498,In_1369,In_1443);
and U1499 (N_1499,In_2230,In_1177);
or U1500 (N_1500,In_1,In_1395);
nor U1501 (N_1501,In_791,In_1224);
and U1502 (N_1502,In_834,In_2300);
or U1503 (N_1503,In_404,In_608);
or U1504 (N_1504,In_1799,In_13);
xor U1505 (N_1505,In_1998,In_84);
nor U1506 (N_1506,In_765,In_714);
xor U1507 (N_1507,In_1370,In_959);
xnor U1508 (N_1508,In_1614,In_561);
or U1509 (N_1509,In_1833,In_575);
xnor U1510 (N_1510,In_1474,In_324);
nand U1511 (N_1511,In_2001,In_2435);
or U1512 (N_1512,In_1177,In_832);
nand U1513 (N_1513,In_1631,In_365);
xnor U1514 (N_1514,In_328,In_1322);
and U1515 (N_1515,In_2017,In_657);
xor U1516 (N_1516,In_1513,In_1068);
or U1517 (N_1517,In_725,In_1006);
or U1518 (N_1518,In_1931,In_2201);
nand U1519 (N_1519,In_1518,In_1760);
xor U1520 (N_1520,In_201,In_2018);
xor U1521 (N_1521,In_1317,In_140);
and U1522 (N_1522,In_1218,In_394);
nand U1523 (N_1523,In_717,In_2246);
and U1524 (N_1524,In_397,In_1491);
and U1525 (N_1525,In_22,In_1277);
and U1526 (N_1526,In_1980,In_1165);
nor U1527 (N_1527,In_120,In_2372);
nor U1528 (N_1528,In_290,In_1459);
or U1529 (N_1529,In_752,In_820);
or U1530 (N_1530,In_98,In_1061);
nand U1531 (N_1531,In_650,In_2030);
and U1532 (N_1532,In_983,In_153);
nand U1533 (N_1533,In_114,In_2241);
xnor U1534 (N_1534,In_2256,In_194);
or U1535 (N_1535,In_54,In_1889);
and U1536 (N_1536,In_1014,In_842);
or U1537 (N_1537,In_1881,In_855);
and U1538 (N_1538,In_151,In_212);
nand U1539 (N_1539,In_2376,In_2333);
or U1540 (N_1540,In_1320,In_303);
and U1541 (N_1541,In_2105,In_169);
and U1542 (N_1542,In_1051,In_2362);
nand U1543 (N_1543,In_35,In_940);
nand U1544 (N_1544,In_512,In_58);
nand U1545 (N_1545,In_897,In_1980);
xnor U1546 (N_1546,In_1791,In_941);
xnor U1547 (N_1547,In_1367,In_255);
nand U1548 (N_1548,In_436,In_829);
nor U1549 (N_1549,In_224,In_68);
xor U1550 (N_1550,In_1054,In_1482);
or U1551 (N_1551,In_984,In_1411);
and U1552 (N_1552,In_49,In_962);
nand U1553 (N_1553,In_1991,In_971);
nor U1554 (N_1554,In_1821,In_2493);
nand U1555 (N_1555,In_1194,In_2225);
or U1556 (N_1556,In_1696,In_2094);
xor U1557 (N_1557,In_1528,In_2244);
nand U1558 (N_1558,In_815,In_200);
and U1559 (N_1559,In_643,In_1713);
xor U1560 (N_1560,In_1470,In_1985);
xor U1561 (N_1561,In_333,In_847);
nand U1562 (N_1562,In_1922,In_449);
nand U1563 (N_1563,In_2037,In_472);
xnor U1564 (N_1564,In_725,In_1667);
xor U1565 (N_1565,In_1190,In_2334);
nand U1566 (N_1566,In_1106,In_2110);
xnor U1567 (N_1567,In_2221,In_2335);
and U1568 (N_1568,In_2492,In_407);
nand U1569 (N_1569,In_756,In_769);
or U1570 (N_1570,In_515,In_1966);
nor U1571 (N_1571,In_1482,In_1621);
xor U1572 (N_1572,In_932,In_792);
nor U1573 (N_1573,In_1019,In_1569);
and U1574 (N_1574,In_271,In_512);
xnor U1575 (N_1575,In_2492,In_2220);
or U1576 (N_1576,In_95,In_651);
and U1577 (N_1577,In_635,In_1392);
xor U1578 (N_1578,In_1157,In_1791);
nor U1579 (N_1579,In_1772,In_664);
nor U1580 (N_1580,In_1315,In_1647);
nand U1581 (N_1581,In_2148,In_508);
or U1582 (N_1582,In_471,In_815);
and U1583 (N_1583,In_1934,In_1231);
nor U1584 (N_1584,In_921,In_1045);
nand U1585 (N_1585,In_1371,In_2029);
or U1586 (N_1586,In_1741,In_1077);
or U1587 (N_1587,In_2396,In_1262);
xnor U1588 (N_1588,In_1746,In_641);
nand U1589 (N_1589,In_1152,In_1220);
and U1590 (N_1590,In_638,In_1987);
xnor U1591 (N_1591,In_1375,In_2296);
xnor U1592 (N_1592,In_1001,In_157);
and U1593 (N_1593,In_654,In_1370);
nor U1594 (N_1594,In_85,In_228);
xor U1595 (N_1595,In_2312,In_572);
and U1596 (N_1596,In_1887,In_1969);
nor U1597 (N_1597,In_2282,In_283);
nor U1598 (N_1598,In_1569,In_992);
or U1599 (N_1599,In_1323,In_2087);
or U1600 (N_1600,In_1662,In_1935);
and U1601 (N_1601,In_5,In_832);
or U1602 (N_1602,In_950,In_2339);
nand U1603 (N_1603,In_1001,In_1488);
xor U1604 (N_1604,In_1782,In_433);
nand U1605 (N_1605,In_1929,In_1552);
nor U1606 (N_1606,In_92,In_1364);
and U1607 (N_1607,In_1416,In_219);
and U1608 (N_1608,In_1495,In_2492);
or U1609 (N_1609,In_1802,In_1239);
nor U1610 (N_1610,In_1691,In_2247);
or U1611 (N_1611,In_1897,In_2387);
xor U1612 (N_1612,In_985,In_370);
nor U1613 (N_1613,In_2100,In_1279);
and U1614 (N_1614,In_472,In_187);
xor U1615 (N_1615,In_1495,In_682);
xor U1616 (N_1616,In_350,In_1957);
nor U1617 (N_1617,In_565,In_1859);
xor U1618 (N_1618,In_1106,In_2073);
nor U1619 (N_1619,In_305,In_1454);
and U1620 (N_1620,In_1126,In_630);
and U1621 (N_1621,In_2327,In_1995);
or U1622 (N_1622,In_1140,In_2464);
nor U1623 (N_1623,In_825,In_1976);
or U1624 (N_1624,In_1591,In_908);
nand U1625 (N_1625,In_1558,In_1350);
xor U1626 (N_1626,In_1738,In_265);
nor U1627 (N_1627,In_685,In_1485);
nand U1628 (N_1628,In_2317,In_1276);
nor U1629 (N_1629,In_471,In_175);
xnor U1630 (N_1630,In_2011,In_1178);
nor U1631 (N_1631,In_1689,In_657);
xor U1632 (N_1632,In_509,In_1206);
nor U1633 (N_1633,In_1403,In_693);
and U1634 (N_1634,In_469,In_1921);
xnor U1635 (N_1635,In_2033,In_2236);
and U1636 (N_1636,In_2298,In_1034);
nor U1637 (N_1637,In_2,In_2431);
and U1638 (N_1638,In_2440,In_29);
xor U1639 (N_1639,In_497,In_1711);
nor U1640 (N_1640,In_631,In_2160);
or U1641 (N_1641,In_2189,In_1338);
nor U1642 (N_1642,In_1458,In_1678);
xor U1643 (N_1643,In_236,In_1084);
xor U1644 (N_1644,In_1832,In_2060);
xnor U1645 (N_1645,In_1453,In_1507);
xnor U1646 (N_1646,In_2487,In_348);
and U1647 (N_1647,In_1176,In_2121);
and U1648 (N_1648,In_1737,In_1268);
and U1649 (N_1649,In_1063,In_1661);
xor U1650 (N_1650,In_355,In_504);
nand U1651 (N_1651,In_1447,In_1819);
or U1652 (N_1652,In_491,In_2092);
and U1653 (N_1653,In_1884,In_774);
or U1654 (N_1654,In_619,In_996);
nor U1655 (N_1655,In_1934,In_379);
nand U1656 (N_1656,In_215,In_791);
nand U1657 (N_1657,In_574,In_1980);
nand U1658 (N_1658,In_236,In_816);
xnor U1659 (N_1659,In_1884,In_1722);
nor U1660 (N_1660,In_2202,In_2118);
and U1661 (N_1661,In_1531,In_751);
nand U1662 (N_1662,In_2102,In_2458);
nor U1663 (N_1663,In_1934,In_2261);
and U1664 (N_1664,In_2365,In_237);
xnor U1665 (N_1665,In_362,In_477);
xnor U1666 (N_1666,In_682,In_1059);
and U1667 (N_1667,In_395,In_1616);
nor U1668 (N_1668,In_940,In_86);
or U1669 (N_1669,In_772,In_2283);
and U1670 (N_1670,In_97,In_2160);
nand U1671 (N_1671,In_2396,In_2089);
xor U1672 (N_1672,In_147,In_767);
xnor U1673 (N_1673,In_1069,In_1527);
xnor U1674 (N_1674,In_2179,In_678);
and U1675 (N_1675,In_683,In_1482);
xnor U1676 (N_1676,In_235,In_2178);
nor U1677 (N_1677,In_1306,In_362);
nand U1678 (N_1678,In_2,In_931);
or U1679 (N_1679,In_925,In_626);
nor U1680 (N_1680,In_1359,In_1496);
nand U1681 (N_1681,In_1903,In_624);
and U1682 (N_1682,In_463,In_784);
or U1683 (N_1683,In_934,In_1786);
and U1684 (N_1684,In_815,In_196);
xnor U1685 (N_1685,In_1826,In_1341);
and U1686 (N_1686,In_1841,In_543);
nor U1687 (N_1687,In_860,In_1239);
nor U1688 (N_1688,In_1241,In_1342);
or U1689 (N_1689,In_1471,In_169);
nor U1690 (N_1690,In_895,In_1786);
xnor U1691 (N_1691,In_211,In_876);
or U1692 (N_1692,In_1940,In_401);
and U1693 (N_1693,In_969,In_200);
and U1694 (N_1694,In_227,In_1256);
nand U1695 (N_1695,In_913,In_183);
nand U1696 (N_1696,In_2387,In_1493);
xor U1697 (N_1697,In_502,In_2438);
or U1698 (N_1698,In_162,In_1757);
nor U1699 (N_1699,In_315,In_35);
nor U1700 (N_1700,In_1818,In_625);
and U1701 (N_1701,In_275,In_1462);
nor U1702 (N_1702,In_1505,In_1790);
nand U1703 (N_1703,In_344,In_1010);
nand U1704 (N_1704,In_651,In_1269);
xnor U1705 (N_1705,In_2334,In_1243);
or U1706 (N_1706,In_1276,In_15);
xnor U1707 (N_1707,In_851,In_1685);
nor U1708 (N_1708,In_2419,In_604);
or U1709 (N_1709,In_2034,In_811);
nor U1710 (N_1710,In_504,In_1767);
xnor U1711 (N_1711,In_1746,In_160);
and U1712 (N_1712,In_1589,In_2387);
and U1713 (N_1713,In_1299,In_1305);
nand U1714 (N_1714,In_835,In_907);
and U1715 (N_1715,In_1712,In_613);
or U1716 (N_1716,In_364,In_406);
nand U1717 (N_1717,In_189,In_2218);
xor U1718 (N_1718,In_2058,In_1887);
and U1719 (N_1719,In_1878,In_1450);
and U1720 (N_1720,In_1233,In_1212);
and U1721 (N_1721,In_1594,In_527);
and U1722 (N_1722,In_503,In_2446);
or U1723 (N_1723,In_2311,In_2249);
xnor U1724 (N_1724,In_894,In_1983);
xnor U1725 (N_1725,In_1290,In_790);
nor U1726 (N_1726,In_1882,In_308);
nor U1727 (N_1727,In_1038,In_1536);
or U1728 (N_1728,In_1888,In_1309);
or U1729 (N_1729,In_1691,In_119);
nand U1730 (N_1730,In_51,In_1492);
or U1731 (N_1731,In_1298,In_1031);
or U1732 (N_1732,In_1019,In_1443);
xor U1733 (N_1733,In_244,In_92);
nand U1734 (N_1734,In_2204,In_2363);
xor U1735 (N_1735,In_1000,In_730);
nor U1736 (N_1736,In_52,In_771);
or U1737 (N_1737,In_2202,In_1256);
and U1738 (N_1738,In_237,In_688);
xor U1739 (N_1739,In_2278,In_458);
nor U1740 (N_1740,In_494,In_191);
and U1741 (N_1741,In_1111,In_2198);
xor U1742 (N_1742,In_1768,In_2035);
nand U1743 (N_1743,In_1466,In_209);
nor U1744 (N_1744,In_1501,In_104);
xor U1745 (N_1745,In_1896,In_570);
xnor U1746 (N_1746,In_1136,In_1430);
nand U1747 (N_1747,In_1944,In_2422);
nor U1748 (N_1748,In_2318,In_1178);
and U1749 (N_1749,In_1671,In_375);
nand U1750 (N_1750,In_766,In_2474);
or U1751 (N_1751,In_1137,In_1036);
xnor U1752 (N_1752,In_54,In_1678);
xor U1753 (N_1753,In_1296,In_101);
xor U1754 (N_1754,In_1058,In_789);
nor U1755 (N_1755,In_1656,In_1056);
nor U1756 (N_1756,In_2279,In_1715);
xor U1757 (N_1757,In_109,In_240);
nor U1758 (N_1758,In_1535,In_356);
nor U1759 (N_1759,In_1158,In_1565);
nor U1760 (N_1760,In_778,In_1966);
nor U1761 (N_1761,In_258,In_1434);
xnor U1762 (N_1762,In_1016,In_546);
xnor U1763 (N_1763,In_2346,In_14);
and U1764 (N_1764,In_883,In_569);
and U1765 (N_1765,In_810,In_1467);
nand U1766 (N_1766,In_1675,In_1374);
or U1767 (N_1767,In_649,In_1951);
nand U1768 (N_1768,In_992,In_2034);
xor U1769 (N_1769,In_658,In_1199);
and U1770 (N_1770,In_1344,In_1246);
xnor U1771 (N_1771,In_414,In_2387);
and U1772 (N_1772,In_1741,In_1272);
nor U1773 (N_1773,In_1943,In_802);
nor U1774 (N_1774,In_1354,In_1684);
or U1775 (N_1775,In_2001,In_1066);
nand U1776 (N_1776,In_469,In_903);
nand U1777 (N_1777,In_1310,In_2089);
or U1778 (N_1778,In_430,In_1725);
nor U1779 (N_1779,In_233,In_1913);
and U1780 (N_1780,In_1139,In_367);
xnor U1781 (N_1781,In_1493,In_1544);
nor U1782 (N_1782,In_788,In_407);
xnor U1783 (N_1783,In_1472,In_2260);
xnor U1784 (N_1784,In_1326,In_146);
xnor U1785 (N_1785,In_1763,In_1210);
xnor U1786 (N_1786,In_1255,In_908);
nand U1787 (N_1787,In_2141,In_937);
nor U1788 (N_1788,In_1086,In_1102);
nor U1789 (N_1789,In_751,In_1577);
nand U1790 (N_1790,In_555,In_2330);
xor U1791 (N_1791,In_447,In_1408);
or U1792 (N_1792,In_1117,In_2302);
nor U1793 (N_1793,In_1270,In_257);
or U1794 (N_1794,In_927,In_1277);
xnor U1795 (N_1795,In_1303,In_1261);
xor U1796 (N_1796,In_1199,In_1911);
nand U1797 (N_1797,In_191,In_933);
nand U1798 (N_1798,In_969,In_132);
xor U1799 (N_1799,In_1942,In_1915);
nor U1800 (N_1800,In_1802,In_2134);
or U1801 (N_1801,In_1394,In_140);
xor U1802 (N_1802,In_1371,In_384);
or U1803 (N_1803,In_644,In_2056);
xnor U1804 (N_1804,In_1350,In_2264);
xor U1805 (N_1805,In_1406,In_2071);
nor U1806 (N_1806,In_1459,In_514);
xnor U1807 (N_1807,In_2191,In_2200);
nor U1808 (N_1808,In_1024,In_1849);
or U1809 (N_1809,In_413,In_1503);
nand U1810 (N_1810,In_484,In_1376);
xor U1811 (N_1811,In_2166,In_1790);
nand U1812 (N_1812,In_1264,In_1142);
and U1813 (N_1813,In_709,In_1731);
and U1814 (N_1814,In_606,In_893);
and U1815 (N_1815,In_2129,In_477);
xor U1816 (N_1816,In_2083,In_42);
or U1817 (N_1817,In_253,In_1663);
and U1818 (N_1818,In_1523,In_1581);
and U1819 (N_1819,In_1839,In_454);
nor U1820 (N_1820,In_830,In_989);
xor U1821 (N_1821,In_1994,In_1459);
nor U1822 (N_1822,In_859,In_59);
xor U1823 (N_1823,In_728,In_379);
xor U1824 (N_1824,In_1008,In_1701);
nand U1825 (N_1825,In_2417,In_181);
nand U1826 (N_1826,In_814,In_930);
nor U1827 (N_1827,In_1740,In_2355);
and U1828 (N_1828,In_2257,In_433);
nand U1829 (N_1829,In_1564,In_1326);
xor U1830 (N_1830,In_693,In_2329);
nor U1831 (N_1831,In_2161,In_1583);
nand U1832 (N_1832,In_362,In_1874);
nor U1833 (N_1833,In_769,In_2349);
or U1834 (N_1834,In_1793,In_1700);
xor U1835 (N_1835,In_886,In_1010);
xnor U1836 (N_1836,In_11,In_493);
and U1837 (N_1837,In_941,In_167);
and U1838 (N_1838,In_1430,In_2138);
or U1839 (N_1839,In_1161,In_1738);
and U1840 (N_1840,In_1943,In_354);
nor U1841 (N_1841,In_687,In_445);
and U1842 (N_1842,In_1133,In_2466);
or U1843 (N_1843,In_573,In_380);
or U1844 (N_1844,In_2320,In_2178);
or U1845 (N_1845,In_153,In_1562);
or U1846 (N_1846,In_97,In_1753);
or U1847 (N_1847,In_2060,In_1360);
xnor U1848 (N_1848,In_1576,In_280);
xnor U1849 (N_1849,In_1414,In_668);
and U1850 (N_1850,In_2169,In_47);
nor U1851 (N_1851,In_1469,In_1532);
or U1852 (N_1852,In_934,In_1642);
nor U1853 (N_1853,In_233,In_1466);
or U1854 (N_1854,In_1367,In_267);
or U1855 (N_1855,In_2422,In_2199);
and U1856 (N_1856,In_202,In_611);
or U1857 (N_1857,In_2107,In_2032);
or U1858 (N_1858,In_1334,In_2288);
or U1859 (N_1859,In_173,In_566);
or U1860 (N_1860,In_1373,In_1542);
xnor U1861 (N_1861,In_791,In_479);
nand U1862 (N_1862,In_128,In_968);
xor U1863 (N_1863,In_971,In_62);
or U1864 (N_1864,In_1422,In_9);
and U1865 (N_1865,In_1681,In_2399);
nand U1866 (N_1866,In_232,In_1066);
xnor U1867 (N_1867,In_901,In_1932);
and U1868 (N_1868,In_2390,In_1839);
nand U1869 (N_1869,In_880,In_260);
and U1870 (N_1870,In_387,In_2216);
nand U1871 (N_1871,In_1634,In_1735);
nor U1872 (N_1872,In_1746,In_1657);
nand U1873 (N_1873,In_1192,In_993);
nor U1874 (N_1874,In_1183,In_1557);
or U1875 (N_1875,In_46,In_2012);
nand U1876 (N_1876,In_1033,In_1378);
nand U1877 (N_1877,In_1645,In_496);
xnor U1878 (N_1878,In_1317,In_2126);
or U1879 (N_1879,In_1485,In_732);
nand U1880 (N_1880,In_2066,In_272);
nor U1881 (N_1881,In_1092,In_2268);
and U1882 (N_1882,In_420,In_841);
xnor U1883 (N_1883,In_1479,In_1009);
or U1884 (N_1884,In_1243,In_1506);
xor U1885 (N_1885,In_1994,In_1738);
xnor U1886 (N_1886,In_1025,In_888);
or U1887 (N_1887,In_283,In_1772);
nand U1888 (N_1888,In_1006,In_1686);
and U1889 (N_1889,In_198,In_231);
and U1890 (N_1890,In_2492,In_962);
nor U1891 (N_1891,In_1393,In_523);
and U1892 (N_1892,In_750,In_1628);
nand U1893 (N_1893,In_1885,In_952);
or U1894 (N_1894,In_2303,In_1698);
nor U1895 (N_1895,In_2216,In_926);
nor U1896 (N_1896,In_2082,In_1684);
xor U1897 (N_1897,In_400,In_2120);
xnor U1898 (N_1898,In_1818,In_675);
nand U1899 (N_1899,In_1675,In_924);
nor U1900 (N_1900,In_715,In_148);
xnor U1901 (N_1901,In_1564,In_1428);
nor U1902 (N_1902,In_1513,In_229);
and U1903 (N_1903,In_1053,In_1840);
or U1904 (N_1904,In_451,In_2353);
and U1905 (N_1905,In_1499,In_652);
or U1906 (N_1906,In_644,In_2255);
xor U1907 (N_1907,In_1368,In_844);
and U1908 (N_1908,In_1330,In_1926);
nand U1909 (N_1909,In_1223,In_698);
nor U1910 (N_1910,In_1986,In_2024);
nand U1911 (N_1911,In_782,In_2396);
and U1912 (N_1912,In_1005,In_405);
and U1913 (N_1913,In_1742,In_2286);
and U1914 (N_1914,In_262,In_128);
nand U1915 (N_1915,In_346,In_410);
nand U1916 (N_1916,In_144,In_1674);
and U1917 (N_1917,In_81,In_1888);
xor U1918 (N_1918,In_761,In_1331);
xnor U1919 (N_1919,In_348,In_486);
and U1920 (N_1920,In_1405,In_1867);
xor U1921 (N_1921,In_131,In_566);
or U1922 (N_1922,In_518,In_737);
and U1923 (N_1923,In_2216,In_192);
nand U1924 (N_1924,In_843,In_410);
xnor U1925 (N_1925,In_2159,In_1711);
xnor U1926 (N_1926,In_1560,In_828);
or U1927 (N_1927,In_6,In_2357);
nand U1928 (N_1928,In_754,In_2016);
nand U1929 (N_1929,In_215,In_1237);
nor U1930 (N_1930,In_724,In_1227);
nand U1931 (N_1931,In_1944,In_1457);
or U1932 (N_1932,In_786,In_2385);
nand U1933 (N_1933,In_287,In_1261);
xor U1934 (N_1934,In_439,In_1058);
or U1935 (N_1935,In_1932,In_2010);
nor U1936 (N_1936,In_1114,In_1819);
nand U1937 (N_1937,In_359,In_54);
xnor U1938 (N_1938,In_1049,In_2076);
or U1939 (N_1939,In_956,In_2381);
or U1940 (N_1940,In_1470,In_1278);
xor U1941 (N_1941,In_1880,In_285);
nand U1942 (N_1942,In_2118,In_1770);
nor U1943 (N_1943,In_1258,In_2218);
and U1944 (N_1944,In_221,In_198);
nor U1945 (N_1945,In_488,In_1875);
and U1946 (N_1946,In_2052,In_1735);
nor U1947 (N_1947,In_1679,In_1484);
xor U1948 (N_1948,In_587,In_2045);
nand U1949 (N_1949,In_368,In_2164);
xor U1950 (N_1950,In_1093,In_1774);
xnor U1951 (N_1951,In_1235,In_960);
or U1952 (N_1952,In_1144,In_2288);
nor U1953 (N_1953,In_1968,In_2136);
nor U1954 (N_1954,In_1291,In_2157);
or U1955 (N_1955,In_2119,In_1605);
xor U1956 (N_1956,In_606,In_2269);
nand U1957 (N_1957,In_799,In_1903);
or U1958 (N_1958,In_1918,In_1612);
xnor U1959 (N_1959,In_1829,In_788);
nand U1960 (N_1960,In_1161,In_745);
xnor U1961 (N_1961,In_2466,In_1779);
nand U1962 (N_1962,In_1135,In_723);
and U1963 (N_1963,In_2066,In_435);
xor U1964 (N_1964,In_784,In_379);
xor U1965 (N_1965,In_1607,In_201);
or U1966 (N_1966,In_1232,In_1204);
nor U1967 (N_1967,In_661,In_364);
nor U1968 (N_1968,In_1931,In_2244);
nor U1969 (N_1969,In_1056,In_638);
nand U1970 (N_1970,In_1917,In_2240);
nor U1971 (N_1971,In_1387,In_774);
or U1972 (N_1972,In_2192,In_1610);
xnor U1973 (N_1973,In_2140,In_639);
xnor U1974 (N_1974,In_355,In_1569);
xnor U1975 (N_1975,In_2258,In_88);
or U1976 (N_1976,In_1414,In_1504);
or U1977 (N_1977,In_393,In_2379);
and U1978 (N_1978,In_338,In_2474);
and U1979 (N_1979,In_2138,In_1774);
and U1980 (N_1980,In_644,In_1091);
nor U1981 (N_1981,In_2391,In_542);
or U1982 (N_1982,In_507,In_67);
and U1983 (N_1983,In_1500,In_705);
xor U1984 (N_1984,In_1285,In_1291);
xor U1985 (N_1985,In_330,In_32);
and U1986 (N_1986,In_609,In_714);
nor U1987 (N_1987,In_143,In_302);
nor U1988 (N_1988,In_1017,In_162);
nand U1989 (N_1989,In_1429,In_1999);
and U1990 (N_1990,In_647,In_293);
and U1991 (N_1991,In_28,In_2209);
nor U1992 (N_1992,In_214,In_2353);
nor U1993 (N_1993,In_2045,In_523);
or U1994 (N_1994,In_1594,In_1056);
or U1995 (N_1995,In_333,In_1463);
nand U1996 (N_1996,In_986,In_424);
or U1997 (N_1997,In_702,In_1166);
xor U1998 (N_1998,In_1404,In_259);
nor U1999 (N_1999,In_1366,In_2049);
xor U2000 (N_2000,In_1165,In_2135);
xnor U2001 (N_2001,In_2432,In_1245);
and U2002 (N_2002,In_95,In_836);
and U2003 (N_2003,In_1658,In_2244);
xor U2004 (N_2004,In_1514,In_2217);
xor U2005 (N_2005,In_1560,In_2420);
xnor U2006 (N_2006,In_2074,In_559);
and U2007 (N_2007,In_1793,In_2143);
or U2008 (N_2008,In_40,In_528);
nand U2009 (N_2009,In_1053,In_245);
and U2010 (N_2010,In_1501,In_2179);
nand U2011 (N_2011,In_1342,In_2368);
and U2012 (N_2012,In_1199,In_2171);
xnor U2013 (N_2013,In_1345,In_609);
and U2014 (N_2014,In_2113,In_2445);
nor U2015 (N_2015,In_1250,In_1670);
or U2016 (N_2016,In_1314,In_865);
nor U2017 (N_2017,In_1680,In_2093);
nor U2018 (N_2018,In_2323,In_1961);
and U2019 (N_2019,In_1919,In_2372);
and U2020 (N_2020,In_591,In_141);
nor U2021 (N_2021,In_1983,In_2351);
nand U2022 (N_2022,In_2190,In_402);
nor U2023 (N_2023,In_925,In_618);
nand U2024 (N_2024,In_2144,In_1773);
xor U2025 (N_2025,In_670,In_357);
xor U2026 (N_2026,In_212,In_1391);
xor U2027 (N_2027,In_345,In_2491);
or U2028 (N_2028,In_1604,In_854);
xor U2029 (N_2029,In_267,In_278);
or U2030 (N_2030,In_2002,In_249);
nor U2031 (N_2031,In_2156,In_43);
and U2032 (N_2032,In_1424,In_1219);
nand U2033 (N_2033,In_1363,In_942);
or U2034 (N_2034,In_18,In_2178);
or U2035 (N_2035,In_2072,In_1688);
or U2036 (N_2036,In_1804,In_1424);
nand U2037 (N_2037,In_2162,In_1031);
xnor U2038 (N_2038,In_145,In_1267);
or U2039 (N_2039,In_579,In_2470);
nor U2040 (N_2040,In_1269,In_385);
or U2041 (N_2041,In_2250,In_1585);
and U2042 (N_2042,In_1183,In_1940);
or U2043 (N_2043,In_2471,In_913);
xor U2044 (N_2044,In_999,In_2107);
nand U2045 (N_2045,In_1826,In_2219);
xor U2046 (N_2046,In_1583,In_2041);
nor U2047 (N_2047,In_372,In_280);
xnor U2048 (N_2048,In_295,In_900);
and U2049 (N_2049,In_1769,In_2000);
nand U2050 (N_2050,In_2368,In_198);
or U2051 (N_2051,In_1627,In_1123);
and U2052 (N_2052,In_2419,In_639);
nor U2053 (N_2053,In_2330,In_1962);
nand U2054 (N_2054,In_2032,In_306);
xnor U2055 (N_2055,In_516,In_2342);
xor U2056 (N_2056,In_2255,In_175);
nor U2057 (N_2057,In_2379,In_1639);
and U2058 (N_2058,In_1209,In_398);
xor U2059 (N_2059,In_494,In_1281);
nand U2060 (N_2060,In_2081,In_1189);
and U2061 (N_2061,In_1785,In_2193);
and U2062 (N_2062,In_2390,In_562);
nand U2063 (N_2063,In_2474,In_2149);
nor U2064 (N_2064,In_273,In_2099);
xor U2065 (N_2065,In_1711,In_1035);
or U2066 (N_2066,In_713,In_1185);
nor U2067 (N_2067,In_16,In_1162);
and U2068 (N_2068,In_95,In_978);
and U2069 (N_2069,In_1031,In_2015);
nand U2070 (N_2070,In_1985,In_1127);
or U2071 (N_2071,In_581,In_1435);
nor U2072 (N_2072,In_2175,In_1862);
nor U2073 (N_2073,In_61,In_1515);
nand U2074 (N_2074,In_1852,In_1935);
nand U2075 (N_2075,In_2452,In_961);
and U2076 (N_2076,In_712,In_933);
or U2077 (N_2077,In_53,In_2100);
and U2078 (N_2078,In_2390,In_173);
and U2079 (N_2079,In_698,In_2431);
nor U2080 (N_2080,In_1660,In_52);
or U2081 (N_2081,In_83,In_1997);
nand U2082 (N_2082,In_1396,In_1418);
nand U2083 (N_2083,In_722,In_1041);
nand U2084 (N_2084,In_1919,In_443);
xnor U2085 (N_2085,In_472,In_1005);
or U2086 (N_2086,In_428,In_1874);
nand U2087 (N_2087,In_679,In_1862);
nor U2088 (N_2088,In_2018,In_290);
xnor U2089 (N_2089,In_2168,In_1284);
and U2090 (N_2090,In_2274,In_1600);
nand U2091 (N_2091,In_1214,In_2257);
nor U2092 (N_2092,In_2468,In_689);
xor U2093 (N_2093,In_116,In_2387);
nor U2094 (N_2094,In_2382,In_601);
nor U2095 (N_2095,In_2104,In_1200);
and U2096 (N_2096,In_1714,In_265);
xor U2097 (N_2097,In_1974,In_1393);
nor U2098 (N_2098,In_678,In_1276);
nor U2099 (N_2099,In_1824,In_221);
nor U2100 (N_2100,In_144,In_2224);
xor U2101 (N_2101,In_892,In_1669);
and U2102 (N_2102,In_1339,In_1157);
nand U2103 (N_2103,In_841,In_1268);
xnor U2104 (N_2104,In_1666,In_1377);
or U2105 (N_2105,In_2033,In_2482);
nand U2106 (N_2106,In_1084,In_740);
nor U2107 (N_2107,In_1580,In_485);
nand U2108 (N_2108,In_177,In_581);
nor U2109 (N_2109,In_1247,In_1203);
xor U2110 (N_2110,In_2227,In_1518);
nand U2111 (N_2111,In_2089,In_1152);
nor U2112 (N_2112,In_819,In_1668);
nor U2113 (N_2113,In_1717,In_39);
nand U2114 (N_2114,In_473,In_2199);
or U2115 (N_2115,In_1339,In_2411);
or U2116 (N_2116,In_1789,In_380);
and U2117 (N_2117,In_1645,In_1332);
nor U2118 (N_2118,In_1281,In_1547);
and U2119 (N_2119,In_2358,In_2449);
nor U2120 (N_2120,In_1184,In_824);
or U2121 (N_2121,In_327,In_2228);
and U2122 (N_2122,In_1327,In_516);
nor U2123 (N_2123,In_2148,In_1081);
or U2124 (N_2124,In_1965,In_530);
nor U2125 (N_2125,In_1307,In_1970);
xor U2126 (N_2126,In_347,In_417);
xnor U2127 (N_2127,In_1026,In_2479);
nor U2128 (N_2128,In_433,In_1914);
nand U2129 (N_2129,In_329,In_528);
xnor U2130 (N_2130,In_470,In_943);
and U2131 (N_2131,In_1974,In_175);
or U2132 (N_2132,In_713,In_1408);
and U2133 (N_2133,In_1846,In_2226);
nand U2134 (N_2134,In_960,In_1024);
and U2135 (N_2135,In_863,In_1020);
xnor U2136 (N_2136,In_612,In_1887);
or U2137 (N_2137,In_894,In_1934);
xor U2138 (N_2138,In_2135,In_1085);
and U2139 (N_2139,In_1779,In_1965);
nor U2140 (N_2140,In_962,In_1031);
nand U2141 (N_2141,In_1843,In_1288);
xnor U2142 (N_2142,In_2058,In_636);
and U2143 (N_2143,In_1319,In_304);
xnor U2144 (N_2144,In_2400,In_2422);
and U2145 (N_2145,In_1441,In_597);
nand U2146 (N_2146,In_1494,In_691);
nor U2147 (N_2147,In_1570,In_511);
nor U2148 (N_2148,In_721,In_572);
nand U2149 (N_2149,In_1112,In_1361);
nand U2150 (N_2150,In_1327,In_2415);
nand U2151 (N_2151,In_1912,In_850);
nand U2152 (N_2152,In_110,In_367);
xnor U2153 (N_2153,In_903,In_1199);
xor U2154 (N_2154,In_12,In_2010);
xor U2155 (N_2155,In_1857,In_242);
and U2156 (N_2156,In_2435,In_1820);
nor U2157 (N_2157,In_217,In_467);
xnor U2158 (N_2158,In_1198,In_775);
xor U2159 (N_2159,In_1929,In_2233);
xor U2160 (N_2160,In_2487,In_157);
nor U2161 (N_2161,In_790,In_2315);
nor U2162 (N_2162,In_2373,In_2303);
or U2163 (N_2163,In_1332,In_1789);
xnor U2164 (N_2164,In_1844,In_261);
xnor U2165 (N_2165,In_420,In_129);
or U2166 (N_2166,In_1876,In_945);
xor U2167 (N_2167,In_1127,In_1690);
nand U2168 (N_2168,In_1170,In_585);
nand U2169 (N_2169,In_2293,In_2223);
and U2170 (N_2170,In_1219,In_1552);
xor U2171 (N_2171,In_1500,In_1518);
nand U2172 (N_2172,In_324,In_1487);
and U2173 (N_2173,In_2401,In_931);
or U2174 (N_2174,In_2184,In_1809);
xnor U2175 (N_2175,In_432,In_2048);
or U2176 (N_2176,In_1153,In_2302);
or U2177 (N_2177,In_1399,In_2114);
nor U2178 (N_2178,In_2235,In_519);
xor U2179 (N_2179,In_1740,In_2312);
or U2180 (N_2180,In_2251,In_513);
xnor U2181 (N_2181,In_1252,In_492);
xor U2182 (N_2182,In_1007,In_225);
or U2183 (N_2183,In_2284,In_1369);
nor U2184 (N_2184,In_1987,In_1105);
and U2185 (N_2185,In_670,In_973);
and U2186 (N_2186,In_1159,In_574);
nand U2187 (N_2187,In_1061,In_1898);
or U2188 (N_2188,In_732,In_1263);
and U2189 (N_2189,In_736,In_1555);
nand U2190 (N_2190,In_2450,In_1201);
nand U2191 (N_2191,In_1337,In_2089);
xor U2192 (N_2192,In_2040,In_945);
and U2193 (N_2193,In_99,In_608);
nor U2194 (N_2194,In_2293,In_1058);
or U2195 (N_2195,In_228,In_1205);
nor U2196 (N_2196,In_1024,In_1215);
nor U2197 (N_2197,In_46,In_2078);
xnor U2198 (N_2198,In_624,In_1196);
and U2199 (N_2199,In_1523,In_2256);
and U2200 (N_2200,In_1456,In_257);
nor U2201 (N_2201,In_670,In_2088);
nand U2202 (N_2202,In_615,In_2368);
and U2203 (N_2203,In_521,In_174);
or U2204 (N_2204,In_868,In_257);
xor U2205 (N_2205,In_2003,In_1050);
and U2206 (N_2206,In_196,In_2498);
nor U2207 (N_2207,In_2051,In_1058);
xnor U2208 (N_2208,In_1132,In_578);
nand U2209 (N_2209,In_94,In_1654);
nand U2210 (N_2210,In_1761,In_1889);
nor U2211 (N_2211,In_318,In_15);
and U2212 (N_2212,In_1984,In_390);
or U2213 (N_2213,In_2313,In_2497);
nand U2214 (N_2214,In_41,In_1816);
xor U2215 (N_2215,In_1443,In_889);
nand U2216 (N_2216,In_664,In_1733);
and U2217 (N_2217,In_2478,In_1915);
nand U2218 (N_2218,In_323,In_2322);
xor U2219 (N_2219,In_820,In_910);
xnor U2220 (N_2220,In_1385,In_1303);
xnor U2221 (N_2221,In_359,In_677);
nor U2222 (N_2222,In_1805,In_1564);
xnor U2223 (N_2223,In_1751,In_637);
and U2224 (N_2224,In_459,In_1609);
xor U2225 (N_2225,In_1602,In_633);
nor U2226 (N_2226,In_1152,In_297);
and U2227 (N_2227,In_2033,In_676);
nand U2228 (N_2228,In_1789,In_2008);
nand U2229 (N_2229,In_286,In_2247);
xnor U2230 (N_2230,In_2254,In_548);
nand U2231 (N_2231,In_629,In_928);
xnor U2232 (N_2232,In_1349,In_2358);
nor U2233 (N_2233,In_1538,In_1085);
or U2234 (N_2234,In_1279,In_738);
and U2235 (N_2235,In_1490,In_1522);
and U2236 (N_2236,In_2083,In_872);
or U2237 (N_2237,In_323,In_1198);
nand U2238 (N_2238,In_2357,In_895);
or U2239 (N_2239,In_1304,In_1624);
nand U2240 (N_2240,In_1613,In_1180);
and U2241 (N_2241,In_1925,In_1100);
and U2242 (N_2242,In_1421,In_2380);
nor U2243 (N_2243,In_1421,In_612);
nand U2244 (N_2244,In_977,In_112);
xor U2245 (N_2245,In_1743,In_627);
or U2246 (N_2246,In_1476,In_262);
or U2247 (N_2247,In_1559,In_2134);
xnor U2248 (N_2248,In_736,In_1088);
nor U2249 (N_2249,In_2192,In_202);
nor U2250 (N_2250,In_2060,In_1958);
xor U2251 (N_2251,In_554,In_1768);
or U2252 (N_2252,In_135,In_2486);
nand U2253 (N_2253,In_2317,In_2336);
nor U2254 (N_2254,In_879,In_384);
nand U2255 (N_2255,In_2291,In_1298);
or U2256 (N_2256,In_160,In_203);
nand U2257 (N_2257,In_764,In_801);
or U2258 (N_2258,In_461,In_1392);
and U2259 (N_2259,In_592,In_394);
and U2260 (N_2260,In_302,In_33);
xor U2261 (N_2261,In_1423,In_79);
or U2262 (N_2262,In_1062,In_2002);
nand U2263 (N_2263,In_1613,In_2369);
xnor U2264 (N_2264,In_1992,In_232);
nand U2265 (N_2265,In_1008,In_2035);
or U2266 (N_2266,In_2169,In_1007);
xnor U2267 (N_2267,In_915,In_2445);
xnor U2268 (N_2268,In_1833,In_2471);
or U2269 (N_2269,In_136,In_2381);
nor U2270 (N_2270,In_584,In_1369);
nor U2271 (N_2271,In_1059,In_190);
nor U2272 (N_2272,In_1784,In_1198);
and U2273 (N_2273,In_1907,In_520);
and U2274 (N_2274,In_24,In_1710);
xor U2275 (N_2275,In_1792,In_1081);
or U2276 (N_2276,In_588,In_1464);
and U2277 (N_2277,In_2371,In_1692);
and U2278 (N_2278,In_433,In_1051);
nor U2279 (N_2279,In_2338,In_1217);
nor U2280 (N_2280,In_39,In_1984);
and U2281 (N_2281,In_1354,In_1637);
nand U2282 (N_2282,In_2243,In_1674);
and U2283 (N_2283,In_141,In_2424);
or U2284 (N_2284,In_1345,In_383);
nand U2285 (N_2285,In_901,In_578);
nand U2286 (N_2286,In_1148,In_1840);
nand U2287 (N_2287,In_463,In_756);
nor U2288 (N_2288,In_2437,In_8);
nand U2289 (N_2289,In_1639,In_1668);
or U2290 (N_2290,In_2267,In_1389);
or U2291 (N_2291,In_1264,In_2039);
xor U2292 (N_2292,In_877,In_340);
nand U2293 (N_2293,In_2305,In_738);
or U2294 (N_2294,In_1997,In_2220);
and U2295 (N_2295,In_558,In_2108);
nand U2296 (N_2296,In_226,In_1596);
nand U2297 (N_2297,In_96,In_900);
and U2298 (N_2298,In_2256,In_1035);
nand U2299 (N_2299,In_226,In_294);
and U2300 (N_2300,In_1886,In_589);
nor U2301 (N_2301,In_1075,In_305);
and U2302 (N_2302,In_2474,In_1713);
nand U2303 (N_2303,In_181,In_467);
xnor U2304 (N_2304,In_566,In_2485);
nor U2305 (N_2305,In_1585,In_2253);
nand U2306 (N_2306,In_659,In_2305);
and U2307 (N_2307,In_365,In_2252);
nor U2308 (N_2308,In_512,In_1663);
nor U2309 (N_2309,In_580,In_1773);
or U2310 (N_2310,In_993,In_1988);
nand U2311 (N_2311,In_199,In_224);
nand U2312 (N_2312,In_596,In_1349);
or U2313 (N_2313,In_1969,In_109);
or U2314 (N_2314,In_164,In_878);
xor U2315 (N_2315,In_1224,In_1408);
xor U2316 (N_2316,In_2147,In_2465);
nor U2317 (N_2317,In_1223,In_2233);
and U2318 (N_2318,In_2059,In_2357);
xor U2319 (N_2319,In_864,In_563);
xnor U2320 (N_2320,In_1860,In_409);
and U2321 (N_2321,In_1934,In_387);
nand U2322 (N_2322,In_908,In_1617);
and U2323 (N_2323,In_1048,In_2158);
xnor U2324 (N_2324,In_642,In_468);
xor U2325 (N_2325,In_2458,In_1888);
nor U2326 (N_2326,In_2197,In_756);
xor U2327 (N_2327,In_1282,In_513);
nand U2328 (N_2328,In_2119,In_2280);
and U2329 (N_2329,In_1473,In_1188);
nand U2330 (N_2330,In_1279,In_966);
nor U2331 (N_2331,In_945,In_1194);
and U2332 (N_2332,In_131,In_1931);
xor U2333 (N_2333,In_2322,In_1924);
and U2334 (N_2334,In_1005,In_74);
or U2335 (N_2335,In_1322,In_182);
or U2336 (N_2336,In_513,In_380);
and U2337 (N_2337,In_349,In_1853);
and U2338 (N_2338,In_2108,In_410);
nor U2339 (N_2339,In_1287,In_1692);
or U2340 (N_2340,In_2171,In_1364);
nand U2341 (N_2341,In_364,In_22);
or U2342 (N_2342,In_1234,In_1242);
or U2343 (N_2343,In_1555,In_1232);
nor U2344 (N_2344,In_298,In_1109);
xnor U2345 (N_2345,In_1538,In_1161);
or U2346 (N_2346,In_424,In_304);
or U2347 (N_2347,In_300,In_535);
or U2348 (N_2348,In_35,In_843);
or U2349 (N_2349,In_2197,In_1728);
nor U2350 (N_2350,In_326,In_1515);
xnor U2351 (N_2351,In_574,In_2417);
nand U2352 (N_2352,In_1201,In_2033);
and U2353 (N_2353,In_2052,In_298);
nand U2354 (N_2354,In_1595,In_1702);
nor U2355 (N_2355,In_1809,In_93);
and U2356 (N_2356,In_284,In_339);
or U2357 (N_2357,In_583,In_1140);
xnor U2358 (N_2358,In_2064,In_693);
nor U2359 (N_2359,In_2229,In_1311);
xnor U2360 (N_2360,In_1024,In_882);
or U2361 (N_2361,In_862,In_1856);
nor U2362 (N_2362,In_1930,In_1340);
xor U2363 (N_2363,In_1538,In_815);
or U2364 (N_2364,In_241,In_2312);
xor U2365 (N_2365,In_565,In_2452);
xor U2366 (N_2366,In_1779,In_1982);
and U2367 (N_2367,In_1191,In_2);
and U2368 (N_2368,In_12,In_353);
nand U2369 (N_2369,In_401,In_650);
and U2370 (N_2370,In_644,In_1159);
nand U2371 (N_2371,In_1351,In_1562);
nor U2372 (N_2372,In_2189,In_1838);
nor U2373 (N_2373,In_1721,In_692);
nor U2374 (N_2374,In_1595,In_2398);
nand U2375 (N_2375,In_1023,In_83);
and U2376 (N_2376,In_404,In_1683);
nand U2377 (N_2377,In_14,In_36);
and U2378 (N_2378,In_2409,In_517);
nand U2379 (N_2379,In_1219,In_110);
or U2380 (N_2380,In_2277,In_183);
or U2381 (N_2381,In_420,In_1941);
and U2382 (N_2382,In_1854,In_101);
nor U2383 (N_2383,In_1301,In_565);
nand U2384 (N_2384,In_1114,In_1361);
nor U2385 (N_2385,In_719,In_1403);
or U2386 (N_2386,In_673,In_1977);
or U2387 (N_2387,In_671,In_1393);
and U2388 (N_2388,In_1430,In_1804);
xor U2389 (N_2389,In_554,In_997);
and U2390 (N_2390,In_541,In_1115);
and U2391 (N_2391,In_500,In_1095);
xnor U2392 (N_2392,In_243,In_192);
or U2393 (N_2393,In_730,In_2189);
and U2394 (N_2394,In_698,In_581);
and U2395 (N_2395,In_2127,In_987);
or U2396 (N_2396,In_1717,In_413);
and U2397 (N_2397,In_2061,In_384);
or U2398 (N_2398,In_1151,In_1082);
nand U2399 (N_2399,In_1009,In_640);
or U2400 (N_2400,In_2168,In_1989);
or U2401 (N_2401,In_1500,In_1172);
nor U2402 (N_2402,In_1015,In_553);
and U2403 (N_2403,In_978,In_610);
or U2404 (N_2404,In_593,In_1753);
or U2405 (N_2405,In_2003,In_1194);
and U2406 (N_2406,In_1484,In_376);
nand U2407 (N_2407,In_970,In_405);
nand U2408 (N_2408,In_447,In_200);
and U2409 (N_2409,In_11,In_1295);
xnor U2410 (N_2410,In_57,In_1289);
nand U2411 (N_2411,In_2438,In_926);
nand U2412 (N_2412,In_2138,In_974);
xor U2413 (N_2413,In_1566,In_323);
or U2414 (N_2414,In_338,In_123);
nand U2415 (N_2415,In_358,In_85);
or U2416 (N_2416,In_1180,In_1190);
nor U2417 (N_2417,In_1717,In_1869);
or U2418 (N_2418,In_1899,In_1752);
nand U2419 (N_2419,In_482,In_632);
xnor U2420 (N_2420,In_189,In_77);
or U2421 (N_2421,In_1152,In_872);
nand U2422 (N_2422,In_1275,In_1443);
and U2423 (N_2423,In_253,In_1507);
nor U2424 (N_2424,In_2368,In_1657);
xnor U2425 (N_2425,In_209,In_313);
or U2426 (N_2426,In_1653,In_873);
xnor U2427 (N_2427,In_1374,In_880);
nor U2428 (N_2428,In_1671,In_2118);
or U2429 (N_2429,In_426,In_2464);
nor U2430 (N_2430,In_428,In_994);
or U2431 (N_2431,In_2029,In_2389);
nand U2432 (N_2432,In_791,In_1323);
and U2433 (N_2433,In_790,In_234);
xnor U2434 (N_2434,In_927,In_1543);
xnor U2435 (N_2435,In_1159,In_2378);
xor U2436 (N_2436,In_303,In_1208);
and U2437 (N_2437,In_611,In_529);
or U2438 (N_2438,In_1710,In_1779);
nor U2439 (N_2439,In_2477,In_488);
and U2440 (N_2440,In_750,In_678);
nor U2441 (N_2441,In_827,In_1780);
xnor U2442 (N_2442,In_1201,In_189);
nor U2443 (N_2443,In_2025,In_906);
nand U2444 (N_2444,In_675,In_1206);
nand U2445 (N_2445,In_2482,In_518);
or U2446 (N_2446,In_2203,In_86);
xnor U2447 (N_2447,In_1439,In_1394);
and U2448 (N_2448,In_2210,In_613);
and U2449 (N_2449,In_1708,In_1007);
nor U2450 (N_2450,In_449,In_2185);
nand U2451 (N_2451,In_1147,In_1351);
xnor U2452 (N_2452,In_1951,In_2181);
xor U2453 (N_2453,In_1397,In_917);
or U2454 (N_2454,In_1731,In_1976);
xor U2455 (N_2455,In_2329,In_1669);
nor U2456 (N_2456,In_2444,In_377);
or U2457 (N_2457,In_1357,In_176);
or U2458 (N_2458,In_1622,In_120);
nor U2459 (N_2459,In_971,In_1809);
or U2460 (N_2460,In_1499,In_1215);
or U2461 (N_2461,In_176,In_2330);
xor U2462 (N_2462,In_597,In_922);
or U2463 (N_2463,In_2447,In_438);
or U2464 (N_2464,In_244,In_1851);
or U2465 (N_2465,In_646,In_1838);
xor U2466 (N_2466,In_1208,In_1574);
xor U2467 (N_2467,In_365,In_424);
nand U2468 (N_2468,In_1305,In_878);
or U2469 (N_2469,In_975,In_2453);
xor U2470 (N_2470,In_1569,In_609);
and U2471 (N_2471,In_95,In_1282);
nand U2472 (N_2472,In_519,In_688);
nor U2473 (N_2473,In_140,In_1927);
nand U2474 (N_2474,In_1428,In_87);
xnor U2475 (N_2475,In_589,In_2284);
nor U2476 (N_2476,In_2443,In_2342);
and U2477 (N_2477,In_1565,In_656);
and U2478 (N_2478,In_1347,In_1593);
and U2479 (N_2479,In_1674,In_2135);
nor U2480 (N_2480,In_1259,In_500);
and U2481 (N_2481,In_550,In_1259);
and U2482 (N_2482,In_26,In_621);
xnor U2483 (N_2483,In_1469,In_1746);
nor U2484 (N_2484,In_257,In_1698);
or U2485 (N_2485,In_947,In_956);
nand U2486 (N_2486,In_978,In_1501);
nand U2487 (N_2487,In_760,In_2070);
xnor U2488 (N_2488,In_1545,In_2026);
xor U2489 (N_2489,In_1477,In_1349);
and U2490 (N_2490,In_2369,In_791);
and U2491 (N_2491,In_538,In_2125);
nand U2492 (N_2492,In_1384,In_1324);
and U2493 (N_2493,In_392,In_991);
nand U2494 (N_2494,In_417,In_1911);
xor U2495 (N_2495,In_1165,In_1503);
xnor U2496 (N_2496,In_2107,In_2042);
and U2497 (N_2497,In_124,In_850);
nand U2498 (N_2498,In_2271,In_2205);
nand U2499 (N_2499,In_1518,In_2209);
nor U2500 (N_2500,N_1722,N_1190);
nor U2501 (N_2501,N_1230,N_1535);
nand U2502 (N_2502,N_1197,N_998);
nand U2503 (N_2503,N_1113,N_2308);
nor U2504 (N_2504,N_2252,N_1804);
nand U2505 (N_2505,N_224,N_464);
or U2506 (N_2506,N_1842,N_715);
nand U2507 (N_2507,N_386,N_199);
xnor U2508 (N_2508,N_830,N_1171);
and U2509 (N_2509,N_679,N_2407);
nor U2510 (N_2510,N_771,N_991);
or U2511 (N_2511,N_688,N_73);
xnor U2512 (N_2512,N_904,N_2019);
xnor U2513 (N_2513,N_1881,N_1703);
xor U2514 (N_2514,N_2422,N_1158);
or U2515 (N_2515,N_241,N_1284);
nand U2516 (N_2516,N_2481,N_406);
or U2517 (N_2517,N_504,N_1093);
or U2518 (N_2518,N_363,N_2180);
xnor U2519 (N_2519,N_460,N_93);
and U2520 (N_2520,N_1925,N_2010);
and U2521 (N_2521,N_1672,N_972);
nor U2522 (N_2522,N_799,N_287);
nor U2523 (N_2523,N_359,N_1721);
and U2524 (N_2524,N_1418,N_1628);
nor U2525 (N_2525,N_2487,N_1243);
nand U2526 (N_2526,N_1958,N_1076);
nand U2527 (N_2527,N_2074,N_1218);
or U2528 (N_2528,N_1392,N_861);
or U2529 (N_2529,N_367,N_635);
xor U2530 (N_2530,N_1050,N_198);
and U2531 (N_2531,N_1936,N_719);
nand U2532 (N_2532,N_742,N_251);
nor U2533 (N_2533,N_1921,N_384);
nand U2534 (N_2534,N_1482,N_1149);
nand U2535 (N_2535,N_2429,N_299);
and U2536 (N_2536,N_1744,N_2021);
xnor U2537 (N_2537,N_146,N_2084);
xnor U2538 (N_2538,N_1588,N_1791);
or U2539 (N_2539,N_54,N_857);
nor U2540 (N_2540,N_1516,N_1521);
nor U2541 (N_2541,N_1009,N_1978);
nand U2542 (N_2542,N_1256,N_321);
and U2543 (N_2543,N_366,N_438);
or U2544 (N_2544,N_2393,N_541);
nand U2545 (N_2545,N_554,N_1123);
nor U2546 (N_2546,N_1550,N_924);
and U2547 (N_2547,N_1705,N_276);
and U2548 (N_2548,N_580,N_2446);
and U2549 (N_2549,N_2050,N_2463);
and U2550 (N_2550,N_1311,N_2207);
nor U2551 (N_2551,N_2317,N_2373);
nand U2552 (N_2552,N_651,N_1956);
nand U2553 (N_2553,N_1655,N_2244);
nor U2554 (N_2554,N_1692,N_1859);
xor U2555 (N_2555,N_2049,N_2182);
nor U2556 (N_2556,N_28,N_1892);
nand U2557 (N_2557,N_1775,N_2167);
or U2558 (N_2558,N_566,N_1984);
or U2559 (N_2559,N_1928,N_2199);
xor U2560 (N_2560,N_600,N_630);
nand U2561 (N_2561,N_2431,N_816);
nor U2562 (N_2562,N_1750,N_2321);
and U2563 (N_2563,N_173,N_472);
and U2564 (N_2564,N_49,N_1203);
and U2565 (N_2565,N_2476,N_2193);
and U2566 (N_2566,N_30,N_394);
and U2567 (N_2567,N_31,N_2192);
or U2568 (N_2568,N_302,N_2117);
nor U2569 (N_2569,N_1668,N_1107);
and U2570 (N_2570,N_1192,N_1678);
nor U2571 (N_2571,N_1572,N_1926);
or U2572 (N_2572,N_1097,N_2283);
nor U2573 (N_2573,N_1834,N_1563);
and U2574 (N_2574,N_2467,N_2189);
nand U2575 (N_2575,N_1031,N_195);
xnor U2576 (N_2576,N_2485,N_255);
xor U2577 (N_2577,N_1150,N_522);
or U2578 (N_2578,N_1346,N_602);
or U2579 (N_2579,N_1480,N_50);
xnor U2580 (N_2580,N_453,N_274);
and U2581 (N_2581,N_2092,N_211);
nor U2582 (N_2582,N_1518,N_398);
xnor U2583 (N_2583,N_2045,N_1752);
xnor U2584 (N_2584,N_1436,N_1843);
nand U2585 (N_2585,N_1904,N_1950);
nor U2586 (N_2586,N_1860,N_974);
or U2587 (N_2587,N_674,N_115);
nand U2588 (N_2588,N_435,N_2079);
and U2589 (N_2589,N_320,N_397);
or U2590 (N_2590,N_434,N_1975);
nand U2591 (N_2591,N_1250,N_41);
xnor U2592 (N_2592,N_956,N_1309);
and U2593 (N_2593,N_1337,N_2368);
or U2594 (N_2594,N_2390,N_947);
and U2595 (N_2595,N_1426,N_1213);
nand U2596 (N_2596,N_687,N_1794);
nor U2597 (N_2597,N_2190,N_2062);
and U2598 (N_2598,N_1157,N_1652);
nand U2599 (N_2599,N_1032,N_98);
or U2600 (N_2600,N_23,N_1607);
nor U2601 (N_2601,N_1347,N_2444);
and U2602 (N_2602,N_576,N_2473);
nor U2603 (N_2603,N_2264,N_758);
nand U2604 (N_2604,N_109,N_1053);
nor U2605 (N_2605,N_2408,N_1144);
nor U2606 (N_2606,N_1078,N_2225);
nor U2607 (N_2607,N_2071,N_1626);
nand U2608 (N_2608,N_1235,N_1786);
and U2609 (N_2609,N_1897,N_1111);
or U2610 (N_2610,N_217,N_1376);
or U2611 (N_2611,N_1627,N_583);
xor U2612 (N_2612,N_1734,N_582);
nand U2613 (N_2613,N_2111,N_370);
xnor U2614 (N_2614,N_569,N_391);
or U2615 (N_2615,N_987,N_650);
xor U2616 (N_2616,N_1452,N_1239);
or U2617 (N_2617,N_806,N_1533);
or U2618 (N_2618,N_551,N_610);
or U2619 (N_2619,N_1109,N_1841);
and U2620 (N_2620,N_2369,N_1382);
xnor U2621 (N_2621,N_596,N_1951);
nand U2622 (N_2622,N_890,N_1911);
nor U2623 (N_2623,N_1504,N_1944);
or U2624 (N_2624,N_706,N_1559);
or U2625 (N_2625,N_2309,N_1151);
xor U2626 (N_2626,N_135,N_38);
nor U2627 (N_2627,N_810,N_63);
nand U2628 (N_2628,N_1275,N_1754);
or U2629 (N_2629,N_2124,N_1642);
or U2630 (N_2630,N_1402,N_1993);
xnor U2631 (N_2631,N_2466,N_1715);
and U2632 (N_2632,N_680,N_1270);
nor U2633 (N_2633,N_228,N_2237);
xor U2634 (N_2634,N_2053,N_2121);
nor U2635 (N_2635,N_247,N_2239);
xor U2636 (N_2636,N_264,N_1933);
xor U2637 (N_2637,N_482,N_1982);
xor U2638 (N_2638,N_1317,N_1593);
nand U2639 (N_2639,N_1524,N_673);
nor U2640 (N_2640,N_1074,N_1315);
xnor U2641 (N_2641,N_933,N_1246);
nand U2642 (N_2642,N_441,N_1938);
xnor U2643 (N_2643,N_1717,N_196);
nor U2644 (N_2644,N_982,N_1994);
xnor U2645 (N_2645,N_1460,N_1294);
and U2646 (N_2646,N_1467,N_1344);
nor U2647 (N_2647,N_2358,N_137);
nor U2648 (N_2648,N_492,N_96);
xor U2649 (N_2649,N_1090,N_727);
and U2650 (N_2650,N_633,N_1731);
nand U2651 (N_2651,N_2277,N_1973);
or U2652 (N_2652,N_2482,N_666);
nand U2653 (N_2653,N_1055,N_332);
nor U2654 (N_2654,N_2093,N_958);
and U2655 (N_2655,N_1289,N_516);
and U2656 (N_2656,N_1654,N_1466);
nand U2657 (N_2657,N_831,N_2007);
nor U2658 (N_2658,N_1539,N_1765);
and U2659 (N_2659,N_1657,N_2307);
nor U2660 (N_2660,N_2426,N_2365);
nor U2661 (N_2661,N_603,N_1531);
nand U2662 (N_2662,N_1199,N_413);
xnor U2663 (N_2663,N_667,N_1831);
nor U2664 (N_2664,N_817,N_14);
and U2665 (N_2665,N_372,N_590);
and U2666 (N_2666,N_166,N_2410);
xnor U2667 (N_2667,N_884,N_1954);
or U2668 (N_2668,N_2331,N_1186);
and U2669 (N_2669,N_2479,N_1512);
or U2670 (N_2670,N_860,N_2069);
or U2671 (N_2671,N_652,N_57);
xnor U2672 (N_2672,N_481,N_918);
xor U2673 (N_2673,N_2102,N_1324);
nand U2674 (N_2674,N_917,N_1306);
and U2675 (N_2675,N_353,N_2371);
nor U2676 (N_2676,N_2300,N_847);
xnor U2677 (N_2677,N_1435,N_1082);
nor U2678 (N_2678,N_1099,N_2278);
and U2679 (N_2679,N_348,N_1699);
and U2680 (N_2680,N_2327,N_685);
and U2681 (N_2681,N_1611,N_2465);
xor U2682 (N_2682,N_2251,N_1704);
nor U2683 (N_2683,N_2144,N_1154);
and U2684 (N_2684,N_1212,N_1671);
and U2685 (N_2685,N_2177,N_2435);
and U2686 (N_2686,N_1995,N_1766);
nor U2687 (N_2687,N_1930,N_735);
nor U2688 (N_2688,N_133,N_794);
or U2689 (N_2689,N_1272,N_835);
nand U2690 (N_2690,N_1903,N_9);
and U2691 (N_2691,N_97,N_1596);
xor U2692 (N_2692,N_1871,N_42);
and U2693 (N_2693,N_517,N_392);
and U2694 (N_2694,N_377,N_1388);
and U2695 (N_2695,N_2209,N_915);
nand U2696 (N_2696,N_486,N_2316);
nand U2697 (N_2697,N_759,N_32);
nand U2698 (N_2698,N_2326,N_1569);
and U2699 (N_2699,N_449,N_2137);
and U2700 (N_2700,N_2459,N_1026);
or U2701 (N_2701,N_2395,N_591);
and U2702 (N_2702,N_2096,N_864);
nand U2703 (N_2703,N_1577,N_1224);
nor U2704 (N_2704,N_1116,N_1266);
and U2705 (N_2705,N_698,N_281);
nand U2706 (N_2706,N_2028,N_190);
and U2707 (N_2707,N_342,N_1019);
nand U2708 (N_2708,N_168,N_1064);
and U2709 (N_2709,N_1906,N_2201);
or U2710 (N_2710,N_1365,N_2115);
and U2711 (N_2711,N_132,N_1856);
and U2712 (N_2712,N_1960,N_2478);
and U2713 (N_2713,N_1378,N_1514);
xnor U2714 (N_2714,N_1812,N_1439);
nor U2715 (N_2715,N_1591,N_92);
nor U2716 (N_2716,N_2200,N_2240);
or U2717 (N_2717,N_709,N_340);
nor U2718 (N_2718,N_1862,N_927);
or U2719 (N_2719,N_978,N_2304);
and U2720 (N_2720,N_2229,N_156);
or U2721 (N_2721,N_1830,N_1404);
and U2722 (N_2722,N_976,N_1542);
nand U2723 (N_2723,N_1736,N_1867);
nand U2724 (N_2724,N_624,N_783);
nor U2725 (N_2725,N_1971,N_2472);
xor U2726 (N_2726,N_1184,N_1983);
nor U2727 (N_2727,N_996,N_1598);
and U2728 (N_2728,N_1422,N_1367);
and U2729 (N_2729,N_1371,N_1264);
and U2730 (N_2730,N_184,N_1789);
nand U2731 (N_2731,N_106,N_1273);
nand U2732 (N_2732,N_665,N_1217);
or U2733 (N_2733,N_2133,N_1268);
or U2734 (N_2734,N_697,N_823);
and U2735 (N_2735,N_1408,N_1229);
or U2736 (N_2736,N_891,N_717);
nor U2737 (N_2737,N_1735,N_162);
nand U2738 (N_2738,N_258,N_2274);
and U2739 (N_2739,N_2039,N_734);
nand U2740 (N_2740,N_1829,N_2445);
nor U2741 (N_2741,N_360,N_445);
nor U2742 (N_2742,N_1413,N_970);
nand U2743 (N_2743,N_171,N_1698);
or U2744 (N_2744,N_722,N_2341);
xnor U2745 (N_2745,N_2403,N_1066);
nor U2746 (N_2746,N_1821,N_2146);
nand U2747 (N_2747,N_344,N_1522);
xor U2748 (N_2748,N_429,N_647);
nand U2749 (N_2749,N_125,N_500);
xnor U2750 (N_2750,N_2234,N_1851);
xor U2751 (N_2751,N_1929,N_1945);
or U2752 (N_2752,N_2103,N_740);
nand U2753 (N_2753,N_2210,N_907);
xor U2754 (N_2754,N_2024,N_975);
nor U2755 (N_2755,N_1648,N_1129);
nand U2756 (N_2756,N_618,N_2017);
and U2757 (N_2757,N_1002,N_1302);
xor U2758 (N_2758,N_2081,N_2352);
and U2759 (N_2759,N_1188,N_2122);
nor U2760 (N_2760,N_1201,N_1262);
or U2761 (N_2761,N_1132,N_440);
nor U2762 (N_2762,N_620,N_1124);
or U2763 (N_2763,N_1981,N_2130);
xor U2764 (N_2764,N_1965,N_1313);
and U2765 (N_2765,N_632,N_2338);
or U2766 (N_2766,N_1156,N_2185);
nor U2767 (N_2767,N_695,N_2033);
or U2768 (N_2768,N_967,N_2227);
and U2769 (N_2769,N_1134,N_1629);
xor U2770 (N_2770,N_757,N_1615);
nor U2771 (N_2771,N_174,N_1549);
or U2772 (N_2772,N_1263,N_1941);
xnor U2773 (N_2773,N_466,N_962);
nor U2774 (N_2774,N_160,N_215);
or U2775 (N_2775,N_311,N_2013);
xor U2776 (N_2776,N_1465,N_1895);
xor U2777 (N_2777,N_37,N_1410);
and U2778 (N_2778,N_1677,N_616);
nor U2779 (N_2779,N_1173,N_916);
xnor U2780 (N_2780,N_658,N_169);
nand U2781 (N_2781,N_693,N_75);
and U2782 (N_2782,N_1205,N_822);
nand U2783 (N_2783,N_382,N_400);
and U2784 (N_2784,N_1327,N_2291);
xnor U2785 (N_2785,N_1281,N_619);
nor U2786 (N_2786,N_1305,N_1145);
nand U2787 (N_2787,N_639,N_1637);
nand U2788 (N_2788,N_739,N_2452);
nand U2789 (N_2789,N_1147,N_520);
xnor U2790 (N_2790,N_219,N_1578);
nand U2791 (N_2791,N_2215,N_2449);
xnor U2792 (N_2792,N_1179,N_1013);
xnor U2793 (N_2793,N_2057,N_1778);
nand U2794 (N_2794,N_462,N_1709);
nand U2795 (N_2795,N_2035,N_724);
nand U2796 (N_2796,N_943,N_1037);
or U2797 (N_2797,N_1809,N_19);
xnor U2798 (N_2798,N_1473,N_1658);
nor U2799 (N_2799,N_1541,N_1152);
xor U2800 (N_2800,N_2401,N_48);
xnor U2801 (N_2801,N_1575,N_1902);
and U2802 (N_2802,N_1363,N_507);
nor U2803 (N_2803,N_1496,N_813);
xnor U2804 (N_2804,N_1373,N_2428);
or U2805 (N_2805,N_2243,N_2443);
nand U2806 (N_2806,N_2391,N_684);
and U2807 (N_2807,N_1101,N_1567);
nand U2808 (N_2808,N_1822,N_2453);
and U2809 (N_2809,N_67,N_1073);
or U2810 (N_2810,N_534,N_1095);
or U2811 (N_2811,N_64,N_1283);
and U2812 (N_2812,N_1661,N_2315);
nor U2813 (N_2813,N_1659,N_505);
nand U2814 (N_2814,N_1247,N_1594);
xnor U2815 (N_2815,N_444,N_256);
and U2816 (N_2816,N_802,N_1085);
xor U2817 (N_2817,N_597,N_1681);
nand U2818 (N_2818,N_833,N_1942);
xnor U2819 (N_2819,N_497,N_2288);
or U2820 (N_2820,N_291,N_1398);
nor U2821 (N_2821,N_1828,N_152);
nor U2822 (N_2822,N_555,N_1308);
xnor U2823 (N_2823,N_932,N_1795);
xor U2824 (N_2824,N_1290,N_1997);
and U2825 (N_2825,N_2415,N_1972);
and U2826 (N_2826,N_2330,N_1837);
nor U2827 (N_2827,N_1343,N_424);
nand U2828 (N_2828,N_1823,N_1599);
nor U2829 (N_2829,N_659,N_1868);
and U2830 (N_2830,N_2249,N_1519);
nand U2831 (N_2831,N_399,N_102);
nor U2832 (N_2832,N_711,N_312);
xnor U2833 (N_2833,N_828,N_804);
or U2834 (N_2834,N_980,N_227);
and U2835 (N_2835,N_1792,N_1348);
nand U2836 (N_2836,N_2179,N_121);
xor U2837 (N_2837,N_1406,N_234);
nand U2838 (N_2838,N_1989,N_1260);
nand U2839 (N_2839,N_712,N_1182);
nand U2840 (N_2840,N_1486,N_105);
nand U2841 (N_2841,N_2191,N_131);
and U2842 (N_2842,N_2499,N_826);
or U2843 (N_2843,N_1310,N_849);
nor U2844 (N_2844,N_1618,N_654);
nor U2845 (N_2845,N_643,N_803);
xor U2846 (N_2846,N_585,N_945);
and U2847 (N_2847,N_147,N_405);
or U2848 (N_2848,N_72,N_553);
or U2849 (N_2849,N_493,N_425);
or U2850 (N_2850,N_252,N_393);
or U2851 (N_2851,N_2483,N_880);
or U2852 (N_2852,N_1852,N_345);
and U2853 (N_2853,N_2236,N_1908);
and U2854 (N_2854,N_1893,N_825);
xnor U2855 (N_2855,N_2165,N_235);
nor U2856 (N_2856,N_494,N_403);
and U2857 (N_2857,N_2231,N_2097);
nor U2858 (N_2858,N_1010,N_936);
or U2859 (N_2859,N_2441,N_754);
xnor U2860 (N_2860,N_2294,N_2153);
or U2861 (N_2861,N_1676,N_1432);
and U2862 (N_2862,N_193,N_1214);
nor U2863 (N_2863,N_751,N_2232);
or U2864 (N_2864,N_237,N_790);
or U2865 (N_2865,N_797,N_1058);
and U2866 (N_2866,N_2344,N_1719);
xnor U2867 (N_2867,N_1146,N_1417);
or U2868 (N_2868,N_990,N_2172);
nor U2869 (N_2869,N_2106,N_692);
nand U2870 (N_2870,N_1356,N_676);
xnor U2871 (N_2871,N_738,N_2470);
xnor U2872 (N_2872,N_454,N_142);
nor U2873 (N_2873,N_2416,N_280);
or U2874 (N_2874,N_528,N_2413);
and U2875 (N_2875,N_81,N_12);
xnor U2876 (N_2876,N_1185,N_1046);
xnor U2877 (N_2877,N_885,N_556);
nor U2878 (N_2878,N_1988,N_1463);
nand U2879 (N_2879,N_2297,N_1219);
nor U2880 (N_2880,N_1877,N_1552);
nor U2881 (N_2881,N_1782,N_2083);
nor U2882 (N_2882,N_1349,N_129);
or U2883 (N_2883,N_1165,N_1853);
xnor U2884 (N_2884,N_2434,N_1189);
nand U2885 (N_2885,N_656,N_2088);
and U2886 (N_2886,N_1314,N_301);
nor U2887 (N_2887,N_713,N_1024);
and U2888 (N_2888,N_856,N_450);
nand U2889 (N_2889,N_1609,N_1445);
xnor U2890 (N_2890,N_1638,N_318);
nand U2891 (N_2891,N_2299,N_1674);
xor U2892 (N_2892,N_766,N_2438);
and U2893 (N_2893,N_310,N_1240);
or U2894 (N_2894,N_2375,N_612);
nand U2895 (N_2895,N_279,N_1040);
and U2896 (N_2896,N_1204,N_1012);
nand U2897 (N_2897,N_2303,N_1481);
nand U2898 (N_2898,N_1211,N_848);
and U2899 (N_2899,N_1104,N_1886);
or U2900 (N_2900,N_1601,N_2089);
or U2901 (N_2901,N_526,N_402);
or U2902 (N_2902,N_447,N_1193);
nor U2903 (N_2903,N_1557,N_273);
xnor U2904 (N_2904,N_2281,N_2197);
nor U2905 (N_2905,N_1056,N_1007);
and U2906 (N_2906,N_1441,N_1469);
nand U2907 (N_2907,N_1774,N_883);
or U2908 (N_2908,N_16,N_509);
nor U2909 (N_2909,N_1168,N_750);
and U2910 (N_2910,N_1336,N_720);
nor U2911 (N_2911,N_346,N_1163);
nor U2912 (N_2912,N_1054,N_1328);
nor U2913 (N_2913,N_1241,N_1511);
xor U2914 (N_2914,N_1641,N_100);
or U2915 (N_2915,N_2094,N_439);
nand U2916 (N_2916,N_2456,N_2109);
or U2917 (N_2917,N_1683,N_786);
or U2918 (N_2918,N_512,N_1548);
nand U2919 (N_2919,N_1375,N_2379);
nand U2920 (N_2920,N_909,N_1350);
or U2921 (N_2921,N_689,N_1632);
nand U2922 (N_2922,N_879,N_1580);
nand U2923 (N_2923,N_1919,N_2168);
xnor U2924 (N_2924,N_2333,N_418);
xnor U2925 (N_2925,N_305,N_2447);
or U2926 (N_2926,N_2376,N_989);
nor U2927 (N_2927,N_163,N_2060);
and U2928 (N_2928,N_894,N_1622);
xor U2929 (N_2929,N_2214,N_1949);
nand U2930 (N_2930,N_1319,N_708);
or U2931 (N_2931,N_113,N_221);
nor U2932 (N_2932,N_1803,N_2034);
and U2933 (N_2933,N_1835,N_1122);
xor U2934 (N_2934,N_561,N_1194);
or U2935 (N_2935,N_1286,N_10);
nor U2936 (N_2936,N_1437,N_1299);
nor U2937 (N_2937,N_396,N_458);
or U2938 (N_2938,N_2388,N_1819);
or U2939 (N_2939,N_545,N_1303);
nor U2940 (N_2940,N_607,N_151);
or U2941 (N_2941,N_809,N_266);
or U2942 (N_2942,N_934,N_1718);
and U2943 (N_2943,N_1503,N_1832);
nor U2944 (N_2944,N_1827,N_1726);
nand U2945 (N_2945,N_1896,N_157);
or U2946 (N_2946,N_7,N_2319);
nor U2947 (N_2947,N_1021,N_859);
nand U2948 (N_2948,N_2009,N_1961);
nand U2949 (N_2949,N_1470,N_415);
and U2950 (N_2950,N_1790,N_1431);
xnor U2951 (N_2951,N_2223,N_2166);
and U2952 (N_2952,N_563,N_858);
and U2953 (N_2953,N_1065,N_1617);
xor U2954 (N_2954,N_1407,N_613);
and U2955 (N_2955,N_546,N_1613);
xor U2956 (N_2956,N_508,N_1636);
nor U2957 (N_2957,N_798,N_671);
and U2958 (N_2958,N_874,N_479);
or U2959 (N_2959,N_476,N_866);
nor U2960 (N_2960,N_2212,N_925);
xor U2961 (N_2961,N_1574,N_21);
nand U2962 (N_2962,N_1833,N_1801);
and U2963 (N_2963,N_22,N_1044);
xnor U2964 (N_2964,N_201,N_2323);
nand U2965 (N_2965,N_1159,N_1811);
and U2966 (N_2966,N_993,N_1566);
nor U2967 (N_2967,N_404,N_260);
xor U2968 (N_2968,N_189,N_1207);
nand U2969 (N_2969,N_69,N_1458);
nand U2970 (N_2970,N_965,N_910);
xnor U2971 (N_2971,N_845,N_1298);
xnor U2972 (N_2972,N_1245,N_2295);
nand U2973 (N_2973,N_335,N_1288);
nand U2974 (N_2974,N_2044,N_1769);
and U2975 (N_2975,N_1321,N_1075);
nor U2976 (N_2976,N_485,N_899);
and U2977 (N_2977,N_1724,N_977);
nand U2978 (N_2978,N_760,N_1568);
and U2979 (N_2979,N_1300,N_71);
nor U2980 (N_2980,N_923,N_1181);
nor U2981 (N_2981,N_82,N_1176);
nor U2982 (N_2982,N_1603,N_183);
nor U2983 (N_2983,N_1720,N_1039);
nor U2984 (N_2984,N_136,N_463);
xnor U2985 (N_2985,N_1669,N_791);
xnor U2986 (N_2986,N_349,N_495);
or U2987 (N_2987,N_1136,N_672);
and U2988 (N_2988,N_981,N_1485);
nor U2989 (N_2989,N_89,N_1633);
and U2990 (N_2990,N_1400,N_746);
or U2991 (N_2991,N_1579,N_457);
and U2992 (N_2992,N_1335,N_2116);
and U2993 (N_2993,N_246,N_1395);
and U2994 (N_2994,N_960,N_1528);
or U2995 (N_2995,N_467,N_1839);
nand U2996 (N_2996,N_1387,N_1425);
or U2997 (N_2997,N_999,N_350);
and U2998 (N_2998,N_593,N_297);
xor U2999 (N_2999,N_1691,N_1106);
nand U3000 (N_3000,N_1934,N_827);
or U3001 (N_3001,N_1377,N_358);
or U3002 (N_3002,N_1962,N_2142);
or U3003 (N_3003,N_2065,N_901);
or U3004 (N_3004,N_1635,N_1475);
xor U3005 (N_3005,N_2157,N_347);
xor U3006 (N_3006,N_627,N_770);
nor U3007 (N_3007,N_1746,N_908);
or U3008 (N_3008,N_498,N_2392);
nand U3009 (N_3009,N_408,N_2173);
or U3010 (N_3010,N_2110,N_2058);
nor U3011 (N_3011,N_390,N_2296);
xnor U3012 (N_3012,N_2363,N_423);
or U3013 (N_3013,N_2397,N_2054);
xor U3014 (N_3014,N_1797,N_1484);
xnor U3015 (N_3015,N_986,N_1035);
and U3016 (N_3016,N_1105,N_839);
xnor U3017 (N_3017,N_2128,N_586);
or U3018 (N_3018,N_780,N_470);
nor U3019 (N_3019,N_1057,N_1079);
or U3020 (N_3020,N_1855,N_657);
and U3021 (N_3021,N_2480,N_490);
or U3022 (N_3022,N_2154,N_2125);
and U3023 (N_3023,N_26,N_304);
nor U3024 (N_3024,N_938,N_1416);
nor U3025 (N_3025,N_1985,N_2382);
nor U3026 (N_3026,N_2343,N_1927);
xnor U3027 (N_3027,N_86,N_1334);
or U3028 (N_3028,N_1816,N_2332);
or U3029 (N_3029,N_1854,N_59);
or U3030 (N_3030,N_2374,N_1330);
or U3031 (N_3031,N_2055,N_868);
nand U3032 (N_3032,N_442,N_805);
xnor U3033 (N_3033,N_6,N_1713);
and U3034 (N_3034,N_767,N_1353);
xor U3035 (N_3035,N_793,N_1543);
xnor U3036 (N_3036,N_1788,N_2404);
nor U3037 (N_3037,N_187,N_1421);
xnor U3038 (N_3038,N_581,N_361);
nand U3039 (N_3039,N_2029,N_298);
nand U3040 (N_3040,N_2170,N_521);
or U3041 (N_3041,N_2078,N_1161);
or U3042 (N_3042,N_776,N_2046);
or U3043 (N_3043,N_953,N_539);
and U3044 (N_3044,N_1225,N_292);
xor U3045 (N_3045,N_542,N_1953);
nand U3046 (N_3046,N_744,N_2005);
xnor U3047 (N_3047,N_1614,N_2155);
or U3048 (N_3048,N_2269,N_2141);
nand U3049 (N_3049,N_180,N_191);
or U3050 (N_3050,N_1228,N_595);
nand U3051 (N_3051,N_2370,N_85);
or U3052 (N_3052,N_368,N_1702);
nor U3053 (N_3053,N_782,N_811);
nor U3054 (N_3054,N_2120,N_2187);
xnor U3055 (N_3055,N_1647,N_774);
nand U3056 (N_3056,N_2112,N_313);
nand U3057 (N_3057,N_589,N_1526);
or U3058 (N_3058,N_1316,N_2131);
or U3059 (N_3059,N_503,N_18);
and U3060 (N_3060,N_78,N_2228);
or U3061 (N_3061,N_240,N_56);
or U3062 (N_3062,N_2276,N_114);
and U3063 (N_3063,N_867,N_1409);
nand U3064 (N_3064,N_118,N_762);
or U3065 (N_3065,N_2086,N_1584);
nor U3066 (N_3066,N_1364,N_378);
nand U3067 (N_3067,N_1495,N_598);
or U3068 (N_3068,N_1068,N_362);
nand U3069 (N_3069,N_242,N_205);
nor U3070 (N_3070,N_309,N_1952);
and U3071 (N_3071,N_2267,N_2256);
xor U3072 (N_3072,N_540,N_1940);
nand U3073 (N_3073,N_814,N_2462);
nor U3074 (N_3074,N_419,N_2381);
nor U3075 (N_3075,N_192,N_2160);
or U3076 (N_3076,N_1741,N_995);
and U3077 (N_3077,N_628,N_1813);
or U3078 (N_3078,N_356,N_642);
or U3079 (N_3079,N_307,N_843);
nor U3080 (N_3080,N_2301,N_1359);
nor U3081 (N_3081,N_1385,N_111);
nand U3082 (N_3082,N_2378,N_412);
nor U3083 (N_3083,N_2147,N_1857);
xor U3084 (N_3084,N_1680,N_2266);
nor U3085 (N_3085,N_968,N_637);
xor U3086 (N_3086,N_897,N_2175);
or U3087 (N_3087,N_1342,N_1894);
nand U3088 (N_3088,N_1725,N_937);
nor U3089 (N_3089,N_1488,N_1527);
nand U3090 (N_3090,N_2275,N_837);
nand U3091 (N_3091,N_1600,N_207);
nand U3092 (N_3092,N_2073,N_1167);
and U3093 (N_3093,N_2002,N_210);
and U3094 (N_3094,N_1478,N_5);
nand U3095 (N_3095,N_515,N_1162);
or U3096 (N_3096,N_11,N_233);
or U3097 (N_3097,N_446,N_1174);
nand U3098 (N_3098,N_1237,N_992);
and U3099 (N_3099,N_79,N_2461);
nor U3100 (N_3100,N_153,N_997);
xnor U3101 (N_3101,N_13,N_2206);
and U3102 (N_3102,N_529,N_58);
xnor U3103 (N_3103,N_426,N_1848);
nor U3104 (N_3104,N_1456,N_119);
xor U3105 (N_3105,N_1667,N_101);
and U3106 (N_3106,N_2328,N_2238);
or U3107 (N_3107,N_471,N_882);
xor U3108 (N_3108,N_1444,N_1459);
xnor U3109 (N_3109,N_2217,N_648);
xor U3110 (N_3110,N_1850,N_2255);
nor U3111 (N_3111,N_1036,N_1779);
nor U3112 (N_3112,N_452,N_2439);
xnor U3113 (N_3113,N_8,N_175);
nor U3114 (N_3114,N_1540,N_784);
nand U3115 (N_3115,N_2164,N_2048);
xor U3116 (N_3116,N_1604,N_1708);
xor U3117 (N_3117,N_1442,N_1625);
xnor U3118 (N_3118,N_1565,N_20);
and U3119 (N_3119,N_1468,N_749);
xnor U3120 (N_3120,N_2196,N_523);
nor U3121 (N_3121,N_2129,N_1255);
and U3122 (N_3122,N_112,N_1238);
nand U3123 (N_3123,N_1297,N_1447);
xnor U3124 (N_3124,N_588,N_1530);
and U3125 (N_3125,N_197,N_716);
or U3126 (N_3126,N_1208,N_1069);
and U3127 (N_3127,N_1963,N_1573);
nor U3128 (N_3128,N_2012,N_1689);
xnor U3129 (N_3129,N_1491,N_2386);
or U3130 (N_3130,N_433,N_682);
nor U3131 (N_3131,N_1826,N_1390);
xor U3132 (N_3132,N_2139,N_2213);
and U3133 (N_3133,N_911,N_765);
nand U3134 (N_3134,N_1501,N_99);
or U3135 (N_3135,N_1818,N_1875);
and U3136 (N_3136,N_572,N_231);
and U3137 (N_3137,N_248,N_1231);
nor U3138 (N_3138,N_1955,N_1307);
xnor U3139 (N_3139,N_2159,N_158);
xor U3140 (N_3140,N_951,N_1651);
or U3141 (N_3141,N_1534,N_186);
or U3142 (N_3142,N_527,N_796);
nor U3143 (N_3143,N_629,N_2140);
or U3144 (N_3144,N_1916,N_2138);
xor U3145 (N_3145,N_355,N_1553);
xnor U3146 (N_3146,N_1340,N_357);
and U3147 (N_3147,N_854,N_1301);
or U3148 (N_3148,N_514,N_465);
nor U3149 (N_3149,N_409,N_1664);
and U3150 (N_3150,N_2184,N_2258);
or U3151 (N_3151,N_778,N_351);
or U3152 (N_3152,N_737,N_188);
nor U3153 (N_3153,N_2286,N_1397);
nor U3154 (N_3154,N_1498,N_1215);
and U3155 (N_3155,N_2220,N_1352);
or U3156 (N_3156,N_1814,N_2027);
or U3157 (N_3157,N_1974,N_605);
nor U3158 (N_3158,N_1049,N_2218);
xor U3159 (N_3159,N_764,N_1061);
xnor U3160 (N_3160,N_24,N_1876);
nand U3161 (N_3161,N_2400,N_1817);
or U3162 (N_3162,N_1991,N_2450);
xor U3163 (N_3163,N_2424,N_1757);
nor U3164 (N_3164,N_1325,N_1840);
or U3165 (N_3165,N_239,N_1236);
or U3166 (N_3166,N_2260,N_2250);
nor U3167 (N_3167,N_104,N_2398);
nor U3168 (N_3168,N_126,N_2489);
nor U3169 (N_3169,N_928,N_1210);
or U3170 (N_3170,N_1610,N_1665);
or U3171 (N_3171,N_718,N_1271);
nand U3172 (N_3172,N_33,N_2366);
nor U3173 (N_3173,N_1198,N_329);
xor U3174 (N_3174,N_203,N_178);
nand U3175 (N_3175,N_1471,N_579);
or U3176 (N_3176,N_25,N_601);
or U3177 (N_3177,N_1379,N_1712);
and U3178 (N_3178,N_2051,N_807);
nor U3179 (N_3179,N_513,N_691);
nand U3180 (N_3180,N_2394,N_1551);
nor U3181 (N_3181,N_2186,N_2272);
and U3182 (N_3182,N_277,N_177);
nand U3183 (N_3183,N_1114,N_1537);
and U3184 (N_3184,N_1621,N_1697);
xnor U3185 (N_3185,N_1362,N_1087);
nand U3186 (N_3186,N_966,N_2246);
or U3187 (N_3187,N_285,N_726);
or U3188 (N_3188,N_83,N_1261);
and U3189 (N_3189,N_636,N_2068);
xnor U3190 (N_3190,N_1368,N_661);
nor U3191 (N_3191,N_2016,N_1924);
xor U3192 (N_3192,N_714,N_939);
and U3193 (N_3193,N_1453,N_1743);
xor U3194 (N_3194,N_1564,N_1429);
and U3195 (N_3195,N_2041,N_2284);
nor U3196 (N_3196,N_2412,N_1092);
or U3197 (N_3197,N_2108,N_1446);
xor U3198 (N_3198,N_1562,N_283);
xor U3199 (N_3199,N_2372,N_204);
xnor U3200 (N_3200,N_138,N_1029);
xor U3201 (N_3201,N_543,N_2474);
nor U3202 (N_3202,N_929,N_2290);
nand U3203 (N_3203,N_518,N_2339);
nor U3204 (N_3204,N_1285,N_1312);
xor U3205 (N_3205,N_1282,N_1003);
or U3206 (N_3206,N_1545,N_1864);
nor U3207 (N_3207,N_2477,N_269);
xnor U3208 (N_3208,N_1538,N_15);
xor U3209 (N_3209,N_322,N_1047);
nand U3210 (N_3210,N_2000,N_1986);
and U3211 (N_3211,N_306,N_1170);
or U3212 (N_3212,N_557,N_2245);
and U3213 (N_3213,N_1755,N_84);
or U3214 (N_3214,N_531,N_27);
nand U3215 (N_3215,N_1084,N_919);
xor U3216 (N_3216,N_1233,N_1126);
xor U3217 (N_3217,N_51,N_655);
or U3218 (N_3218,N_1706,N_284);
xor U3219 (N_3219,N_2101,N_1711);
nor U3220 (N_3220,N_920,N_2451);
nor U3221 (N_3221,N_1202,N_873);
nor U3222 (N_3222,N_232,N_2126);
or U3223 (N_3223,N_2156,N_646);
nor U3224 (N_3224,N_1753,N_2492);
xnor U3225 (N_3225,N_1493,N_779);
nor U3226 (N_3226,N_1131,N_2345);
nor U3227 (N_3227,N_1222,N_1175);
or U3228 (N_3228,N_2364,N_47);
nor U3229 (N_3229,N_756,N_1141);
nor U3230 (N_3230,N_2032,N_461);
and U3231 (N_3231,N_1226,N_1515);
nor U3232 (N_3232,N_123,N_428);
xnor U3233 (N_3233,N_2336,N_1682);
or U3234 (N_3234,N_1383,N_1115);
and U3235 (N_3235,N_1582,N_2334);
nor U3236 (N_3236,N_1968,N_272);
xnor U3237 (N_3237,N_143,N_1060);
nor U3238 (N_3238,N_40,N_343);
or U3239 (N_3239,N_2399,N_2282);
nand U3240 (N_3240,N_2247,N_167);
nor U3241 (N_3241,N_468,N_2104);
and U3242 (N_3242,N_1517,N_2329);
xor U3243 (N_3243,N_2406,N_1694);
nand U3244 (N_3244,N_2488,N_66);
or U3245 (N_3245,N_1849,N_1670);
and U3246 (N_3246,N_2396,N_1434);
nand U3247 (N_3247,N_1380,N_209);
and U3248 (N_3248,N_1164,N_2285);
and U3249 (N_3249,N_55,N_952);
nor U3250 (N_3250,N_753,N_2494);
or U3251 (N_3251,N_2337,N_1663);
xnor U3252 (N_3252,N_2248,N_2095);
xor U3253 (N_3253,N_944,N_1685);
nor U3254 (N_3254,N_1045,N_295);
xor U3255 (N_3255,N_2208,N_2216);
and U3256 (N_3256,N_631,N_1571);
xnor U3257 (N_3257,N_1597,N_2036);
nand U3258 (N_3258,N_1634,N_2423);
or U3259 (N_3259,N_921,N_259);
or U3260 (N_3260,N_1806,N_1232);
nor U3261 (N_3261,N_455,N_573);
nor U3262 (N_3262,N_469,N_1389);
or U3263 (N_3263,N_1544,N_1785);
or U3264 (N_3264,N_1560,N_1980);
and U3265 (N_3265,N_2241,N_110);
nand U3266 (N_3266,N_1883,N_2085);
or U3267 (N_3267,N_294,N_2349);
and U3268 (N_3268,N_1909,N_2158);
or U3269 (N_3269,N_95,N_29);
xnor U3270 (N_3270,N_1401,N_2075);
nand U3271 (N_3271,N_484,N_2497);
or U3272 (N_3272,N_2015,N_140);
and U3273 (N_3273,N_547,N_2312);
xnor U3274 (N_3274,N_1280,N_819);
or U3275 (N_3275,N_1403,N_1957);
nand U3276 (N_3276,N_1443,N_733);
xnor U3277 (N_3277,N_2475,N_1020);
xnor U3278 (N_3278,N_1267,N_2496);
and U3279 (N_3279,N_946,N_43);
nor U3280 (N_3280,N_1172,N_941);
and U3281 (N_3281,N_959,N_1748);
nand U3282 (N_3282,N_379,N_2261);
xor U3283 (N_3283,N_1701,N_65);
nand U3284 (N_3284,N_2263,N_2351);
or U3285 (N_3285,N_2145,N_1138);
and U3286 (N_3286,N_2491,N_983);
xnor U3287 (N_3287,N_1887,N_414);
nand U3288 (N_3288,N_2233,N_478);
or U3289 (N_3289,N_877,N_988);
xor U3290 (N_3290,N_124,N_2134);
nor U3291 (N_3291,N_875,N_1027);
xor U3292 (N_3292,N_1287,N_2359);
and U3293 (N_3293,N_376,N_337);
nor U3294 (N_3294,N_2314,N_1923);
nand U3295 (N_3295,N_2025,N_1177);
nor U3296 (N_3296,N_985,N_369);
or U3297 (N_3297,N_1523,N_510);
xnor U3298 (N_3298,N_336,N_1913);
or U3299 (N_3299,N_263,N_1148);
nand U3300 (N_3300,N_68,N_1624);
or U3301 (N_3301,N_1077,N_2056);
xor U3302 (N_3302,N_243,N_1384);
nand U3303 (N_3303,N_699,N_1687);
xnor U3304 (N_3304,N_1937,N_752);
and U3305 (N_3305,N_1767,N_149);
and U3306 (N_3306,N_900,N_2067);
and U3307 (N_3307,N_1884,N_134);
nor U3308 (N_3308,N_675,N_2495);
nor U3309 (N_3309,N_35,N_1331);
or U3310 (N_3310,N_354,N_1646);
nor U3311 (N_3311,N_2305,N_328);
nand U3312 (N_3312,N_922,N_1023);
nor U3313 (N_3313,N_840,N_1729);
nand U3314 (N_3314,N_4,N_2498);
nand U3315 (N_3315,N_1391,N_1999);
nand U3316 (N_3316,N_293,N_1454);
nor U3317 (N_3317,N_62,N_2457);
xnor U3318 (N_3318,N_575,N_2324);
xor U3319 (N_3319,N_1366,N_387);
nor U3320 (N_3320,N_2148,N_1381);
or U3321 (N_3321,N_536,N_1216);
or U3322 (N_3322,N_1427,N_1497);
or U3323 (N_3323,N_325,N_664);
nor U3324 (N_3324,N_1355,N_1772);
or U3325 (N_3325,N_748,N_2289);
xor U3326 (N_3326,N_544,N_2059);
and U3327 (N_3327,N_17,N_2273);
nand U3328 (N_3328,N_2409,N_1372);
or U3329 (N_3329,N_808,N_788);
xnor U3330 (N_3330,N_747,N_769);
nand U3331 (N_3331,N_926,N_781);
or U3332 (N_3332,N_902,N_2099);
xor U3333 (N_3333,N_60,N_1922);
or U3334 (N_3334,N_571,N_1433);
xnor U3335 (N_3335,N_1561,N_851);
and U3336 (N_3336,N_2335,N_2347);
nor U3337 (N_3337,N_244,N_940);
nor U3338 (N_3338,N_2486,N_45);
nand U3339 (N_3339,N_1351,N_448);
xnor U3340 (N_3340,N_1693,N_930);
or U3341 (N_3341,N_1510,N_853);
nor U3342 (N_3342,N_2417,N_443);
xnor U3343 (N_3343,N_896,N_821);
nor U3344 (N_3344,N_2038,N_364);
or U3345 (N_3345,N_1630,N_2204);
nor U3346 (N_3346,N_422,N_865);
or U3347 (N_3347,N_1872,N_1656);
xnor U3348 (N_3348,N_1135,N_2);
or U3349 (N_3349,N_2136,N_2082);
nand U3350 (N_3350,N_1874,N_1640);
or U3351 (N_3351,N_1461,N_2411);
xnor U3352 (N_3352,N_290,N_824);
and U3353 (N_3353,N_942,N_913);
nor U3354 (N_3354,N_1879,N_1292);
xor U3355 (N_3355,N_592,N_1191);
nor U3356 (N_3356,N_2066,N_1616);
and U3357 (N_3357,N_892,N_289);
nand U3358 (N_3358,N_2471,N_1608);
nor U3359 (N_3359,N_795,N_1004);
or U3360 (N_3360,N_1142,N_2001);
or U3361 (N_3361,N_2222,N_1419);
and U3362 (N_3362,N_2322,N_1590);
nand U3363 (N_3363,N_2203,N_2259);
xnor U3364 (N_3364,N_1341,N_1361);
nor U3365 (N_3365,N_44,N_1592);
or U3366 (N_3366,N_427,N_1808);
nor U3367 (N_3367,N_895,N_649);
xnor U3368 (N_3368,N_1679,N_1244);
nand U3369 (N_3369,N_1979,N_768);
and U3370 (N_3370,N_844,N_1763);
or U3371 (N_3371,N_1730,N_2306);
or U3372 (N_3372,N_772,N_1555);
xnor U3373 (N_3373,N_725,N_46);
nand U3374 (N_3374,N_905,N_1259);
xnor U3375 (N_3375,N_1770,N_288);
nand U3376 (N_3376,N_1898,N_385);
nand U3377 (N_3377,N_2077,N_1589);
xor U3378 (N_3378,N_474,N_755);
nor U3379 (N_3379,N_2030,N_2178);
and U3380 (N_3380,N_1508,N_338);
xor U3381 (N_3381,N_2004,N_732);
or U3382 (N_3382,N_489,N_2464);
or U3383 (N_3383,N_2493,N_331);
or U3384 (N_3384,N_1771,N_1990);
nand U3385 (N_3385,N_2022,N_34);
nor U3386 (N_3386,N_2436,N_2205);
xnor U3387 (N_3387,N_2420,N_139);
and U3388 (N_3388,N_1759,N_130);
nor U3389 (N_3389,N_599,N_1932);
xnor U3390 (N_3390,N_773,N_549);
and U3391 (N_3391,N_1606,N_451);
nand U3392 (N_3392,N_1998,N_1043);
nor U3393 (N_3393,N_838,N_641);
xnor U3394 (N_3394,N_1424,N_2380);
and U3395 (N_3395,N_1000,N_2018);
or U3396 (N_3396,N_1776,N_2320);
nor U3397 (N_3397,N_1546,N_963);
or U3398 (N_3398,N_2202,N_416);
and U3399 (N_3399,N_881,N_660);
nor U3400 (N_3400,N_1118,N_532);
and U3401 (N_3401,N_1970,N_1749);
and U3402 (N_3402,N_1030,N_530);
and U3403 (N_3403,N_1870,N_316);
or U3404 (N_3404,N_2098,N_2114);
and U3405 (N_3405,N_388,N_570);
or U3406 (N_3406,N_410,N_2427);
xor U3407 (N_3407,N_417,N_1304);
and U3408 (N_3408,N_315,N_473);
or U3409 (N_3409,N_1258,N_1083);
or U3410 (N_3410,N_1130,N_1015);
or U3411 (N_3411,N_957,N_730);
or U3412 (N_3412,N_1196,N_2221);
and U3413 (N_3413,N_604,N_52);
and U3414 (N_3414,N_761,N_1326);
nand U3415 (N_3415,N_220,N_1992);
or U3416 (N_3416,N_1278,N_1602);
or U3417 (N_3417,N_568,N_1094);
and U3418 (N_3418,N_1121,N_511);
nor U3419 (N_3419,N_2235,N_1483);
xnor U3420 (N_3420,N_2265,N_2224);
and U3421 (N_3421,N_145,N_801);
or U3422 (N_3422,N_1695,N_1110);
nand U3423 (N_3423,N_842,N_1532);
or U3424 (N_3424,N_729,N_1354);
or U3425 (N_3425,N_1357,N_1052);
nand U3426 (N_3426,N_1996,N_116);
nor U3427 (N_3427,N_1102,N_161);
nor U3428 (N_3428,N_2163,N_949);
and U3429 (N_3429,N_1451,N_1291);
or U3430 (N_3430,N_202,N_225);
nand U3431 (N_3431,N_1824,N_1011);
xor U3432 (N_3432,N_2311,N_1838);
xor U3433 (N_3433,N_1411,N_1917);
xor U3434 (N_3434,N_1062,N_2183);
and U3435 (N_3435,N_1662,N_800);
xor U3436 (N_3436,N_2402,N_2242);
nor U3437 (N_3437,N_1825,N_117);
xnor U3438 (N_3438,N_950,N_475);
or U3439 (N_3439,N_1959,N_2076);
nand U3440 (N_3440,N_254,N_889);
and U3441 (N_3441,N_1345,N_334);
nand U3442 (N_3442,N_669,N_1025);
and U3443 (N_3443,N_127,N_1457);
and U3444 (N_3444,N_1858,N_1899);
and U3445 (N_3445,N_229,N_2405);
or U3446 (N_3446,N_1967,N_2468);
xnor U3447 (N_3447,N_584,N_2135);
xor U3448 (N_3448,N_745,N_261);
nand U3449 (N_3449,N_1946,N_2003);
nand U3450 (N_3450,N_832,N_374);
nor U3451 (N_3451,N_1509,N_1619);
nand U3452 (N_3452,N_1448,N_491);
xor U3453 (N_3453,N_1252,N_670);
or U3454 (N_3454,N_1479,N_562);
nor U3455 (N_3455,N_1987,N_2279);
xnor U3456 (N_3456,N_155,N_159);
xor U3457 (N_3457,N_2268,N_1117);
and U3458 (N_3458,N_1042,N_2127);
nor U3459 (N_3459,N_710,N_2362);
xnor U3460 (N_3460,N_2072,N_2042);
and U3461 (N_3461,N_1947,N_496);
nor U3462 (N_3462,N_1554,N_1133);
xnor U3463 (N_3463,N_2385,N_1091);
or U3464 (N_3464,N_1464,N_2318);
or U3465 (N_3465,N_1318,N_1169);
xnor U3466 (N_3466,N_2293,N_2355);
or U3467 (N_3467,N_2151,N_1254);
or U3468 (N_3468,N_1296,N_931);
nor U3469 (N_3469,N_787,N_212);
or U3470 (N_3470,N_2052,N_267);
xor U3471 (N_3471,N_2230,N_846);
or U3472 (N_3472,N_1462,N_1733);
or U3473 (N_3473,N_519,N_268);
or U3474 (N_3474,N_1861,N_1710);
nor U3475 (N_3475,N_327,N_314);
nor U3476 (N_3476,N_506,N_432);
xnor U3477 (N_3477,N_1873,N_373);
xor U3478 (N_3478,N_1581,N_872);
and U3479 (N_3479,N_1071,N_1847);
and U3480 (N_3480,N_2440,N_1143);
nand U3481 (N_3481,N_2008,N_2357);
xor U3482 (N_3482,N_2353,N_984);
nand U3483 (N_3483,N_1067,N_1505);
xnor U3484 (N_3484,N_994,N_1783);
nand U3485 (N_3485,N_1494,N_1455);
nor U3486 (N_3486,N_2310,N_2442);
nand U3487 (N_3487,N_154,N_1051);
and U3488 (N_3488,N_1490,N_1948);
xnor U3489 (N_3489,N_2361,N_775);
xnor U3490 (N_3490,N_2132,N_2105);
nand U3491 (N_3491,N_2149,N_300);
nor U3492 (N_3492,N_430,N_812);
nor U3493 (N_3493,N_1474,N_1583);
xnor U3494 (N_3494,N_223,N_1166);
nor U3495 (N_3495,N_181,N_1420);
or U3496 (N_3496,N_577,N_2162);
or U3497 (N_3497,N_1796,N_1815);
or U3498 (N_3498,N_1740,N_2354);
nand U3499 (N_3499,N_1103,N_1866);
and U3500 (N_3500,N_2169,N_564);
nand U3501 (N_3501,N_567,N_176);
nand U3502 (N_3502,N_2414,N_1888);
xnor U3503 (N_3503,N_1017,N_1412);
nor U3504 (N_3504,N_2026,N_1070);
nor U3505 (N_3505,N_2325,N_172);
xnor U3506 (N_3506,N_94,N_914);
nand U3507 (N_3507,N_2040,N_2287);
nand U3508 (N_3508,N_1742,N_2257);
or U3509 (N_3509,N_2360,N_1080);
and U3510 (N_3510,N_502,N_179);
xnor U3511 (N_3511,N_640,N_871);
and U3512 (N_3512,N_611,N_108);
and U3513 (N_3513,N_303,N_420);
xnor U3514 (N_3514,N_964,N_948);
xnor U3515 (N_3515,N_265,N_1869);
xor U3516 (N_3516,N_2023,N_2047);
nand U3517 (N_3517,N_480,N_2198);
and U3518 (N_3518,N_1251,N_663);
nand U3519 (N_3519,N_182,N_1605);
or U3520 (N_3520,N_250,N_870);
and U3521 (N_3521,N_863,N_1836);
nand U3522 (N_3522,N_728,N_862);
xor U3523 (N_3523,N_1180,N_1912);
nor U3524 (N_3524,N_1394,N_622);
or U3525 (N_3525,N_1805,N_1525);
nor U3526 (N_3526,N_1773,N_319);
nor U3527 (N_3527,N_1127,N_395);
nand U3528 (N_3528,N_1728,N_1865);
xor U3529 (N_3529,N_888,N_829);
or U3530 (N_3530,N_1249,N_1891);
nor U3531 (N_3531,N_1690,N_1639);
and U3532 (N_3532,N_1333,N_53);
or U3533 (N_3533,N_1449,N_2418);
xor U3534 (N_3534,N_678,N_1799);
nand U3535 (N_3535,N_694,N_898);
nand U3536 (N_3536,N_326,N_763);
nand U3537 (N_3537,N_1028,N_375);
xnor U3538 (N_3538,N_2080,N_1901);
nand U3539 (N_3539,N_855,N_1220);
or U3540 (N_3540,N_2302,N_1977);
xnor U3541 (N_3541,N_2340,N_681);
xor U3542 (N_3542,N_606,N_2342);
xor U3543 (N_3543,N_700,N_1576);
or U3544 (N_3544,N_1863,N_1666);
or U3545 (N_3545,N_1034,N_2433);
nand U3546 (N_3546,N_1119,N_1125);
and U3547 (N_3547,N_820,N_483);
xor U3548 (N_3548,N_1223,N_1585);
or U3549 (N_3549,N_701,N_1358);
xnor U3550 (N_3550,N_1277,N_609);
xnor U3551 (N_3551,N_621,N_954);
xnor U3552 (N_3552,N_741,N_381);
nand U3553 (N_3553,N_286,N_2458);
and U3554 (N_3554,N_3,N_1005);
xnor U3555 (N_3555,N_2298,N_2226);
or U3556 (N_3556,N_1976,N_1137);
or U3557 (N_3557,N_560,N_702);
xor U3558 (N_3558,N_1820,N_906);
xnor U3559 (N_3559,N_436,N_2377);
nor U3560 (N_3560,N_1112,N_1756);
and U3561 (N_3561,N_731,N_2031);
and U3562 (N_3562,N_120,N_1438);
xnor U3563 (N_3563,N_1800,N_1038);
or U3564 (N_3564,N_777,N_785);
and U3565 (N_3565,N_323,N_1643);
xnor U3566 (N_3566,N_1016,N_1048);
nand U3567 (N_3567,N_39,N_76);
and U3568 (N_3568,N_80,N_1506);
xnor U3569 (N_3569,N_615,N_2455);
nor U3570 (N_3570,N_218,N_2432);
nand U3571 (N_3571,N_608,N_1072);
nand U3572 (N_3572,N_1492,N_128);
nand U3573 (N_3573,N_1089,N_1747);
or U3574 (N_3574,N_1178,N_2484);
xnor U3575 (N_3575,N_2262,N_903);
nor U3576 (N_3576,N_371,N_1414);
and U3577 (N_3577,N_1450,N_2425);
nor U3578 (N_3578,N_170,N_2219);
and U3579 (N_3579,N_74,N_736);
or U3580 (N_3580,N_1762,N_912);
nor U3581 (N_3581,N_1269,N_1155);
and U3582 (N_3582,N_1428,N_222);
xnor U3583 (N_3583,N_271,N_1221);
nor U3584 (N_3584,N_638,N_2091);
nor U3585 (N_3585,N_2100,N_1018);
xnor U3586 (N_3586,N_185,N_1935);
nor U3587 (N_3587,N_789,N_499);
xnor U3588 (N_3588,N_365,N_1931);
or U3589 (N_3589,N_1008,N_1499);
nor U3590 (N_3590,N_0,N_1910);
nor U3591 (N_3591,N_2143,N_1472);
and U3592 (N_3592,N_2152,N_1022);
and U3593 (N_3593,N_1882,N_501);
or U3594 (N_3594,N_2292,N_574);
or U3595 (N_3595,N_208,N_1209);
and U3596 (N_3596,N_617,N_1370);
and U3597 (N_3597,N_150,N_626);
nor U3598 (N_3598,N_1764,N_1660);
xnor U3599 (N_3599,N_2090,N_103);
and U3600 (N_3600,N_1033,N_1738);
and U3601 (N_3601,N_141,N_1649);
and U3602 (N_3602,N_324,N_308);
nor U3603 (N_3603,N_61,N_707);
nand U3604 (N_3604,N_1631,N_122);
nor U3605 (N_3605,N_1966,N_815);
nand U3606 (N_3606,N_1612,N_1360);
nor U3607 (N_3607,N_1529,N_2006);
nand U3608 (N_3608,N_1623,N_2419);
nand U3609 (N_3609,N_1696,N_1587);
and U3610 (N_3610,N_2043,N_2356);
and U3611 (N_3611,N_477,N_2194);
or U3612 (N_3612,N_1339,N_704);
and U3613 (N_3613,N_683,N_973);
and U3614 (N_3614,N_2150,N_2421);
and U3615 (N_3615,N_2270,N_317);
nand U3616 (N_3616,N_1374,N_2350);
nand U3617 (N_3617,N_1810,N_1758);
nor U3618 (N_3618,N_792,N_535);
nor U3619 (N_3619,N_36,N_653);
nand U3620 (N_3620,N_194,N_459);
or U3621 (N_3621,N_352,N_1844);
or U3622 (N_3622,N_2348,N_2383);
or U3623 (N_3623,N_1650,N_2011);
nor U3624 (N_3624,N_559,N_1183);
and U3625 (N_3625,N_645,N_87);
and U3626 (N_3626,N_1520,N_282);
or U3627 (N_3627,N_1415,N_2188);
and U3628 (N_3628,N_2070,N_587);
xnor U3629 (N_3629,N_487,N_662);
or U3630 (N_3630,N_1086,N_2176);
nor U3631 (N_3631,N_1586,N_1399);
nand U3632 (N_3632,N_70,N_1393);
or U3633 (N_3633,N_686,N_1500);
nor U3634 (N_3634,N_2313,N_389);
xor U3635 (N_3635,N_893,N_1120);
nand U3636 (N_3636,N_1802,N_206);
nand U3637 (N_3637,N_213,N_2061);
nand U3638 (N_3638,N_1477,N_2490);
and U3639 (N_3639,N_1081,N_77);
and U3640 (N_3640,N_1059,N_1098);
nand U3641 (N_3641,N_2195,N_1100);
and U3642 (N_3642,N_383,N_1536);
and U3643 (N_3643,N_1320,N_1513);
nand U3644 (N_3644,N_1890,N_1338);
xor U3645 (N_3645,N_1900,N_1253);
nand U3646 (N_3646,N_565,N_668);
and U3647 (N_3647,N_1777,N_1195);
nor U3648 (N_3648,N_743,N_1889);
nor U3649 (N_3649,N_1200,N_2113);
xnor U3650 (N_3650,N_330,N_1907);
nor U3651 (N_3651,N_969,N_216);
and U3652 (N_3652,N_262,N_245);
nor U3653 (N_3653,N_257,N_2020);
nand U3654 (N_3654,N_2254,N_1807);
or U3655 (N_3655,N_1279,N_1440);
nand U3656 (N_3656,N_230,N_1969);
nor U3657 (N_3657,N_275,N_703);
and U3658 (N_3658,N_1487,N_1845);
xor U3659 (N_3659,N_1507,N_614);
or U3660 (N_3660,N_1,N_296);
nand U3661 (N_3661,N_1242,N_2181);
nor U3662 (N_3662,N_623,N_594);
nor U3663 (N_3663,N_1644,N_1595);
and U3664 (N_3664,N_270,N_2107);
and U3665 (N_3665,N_1323,N_2469);
and U3666 (N_3666,N_1653,N_2280);
nand U3667 (N_3667,N_1257,N_1686);
and U3668 (N_3668,N_431,N_1716);
nor U3669 (N_3669,N_1673,N_1798);
nand U3670 (N_3670,N_721,N_144);
nand U3671 (N_3671,N_1153,N_2437);
nand U3672 (N_3672,N_1920,N_1234);
nand U3673 (N_3673,N_2171,N_164);
nor U3674 (N_3674,N_1187,N_238);
and U3675 (N_3675,N_696,N_1386);
nor U3676 (N_3676,N_456,N_1041);
nand U3677 (N_3677,N_1723,N_1489);
nand U3678 (N_3678,N_1088,N_2119);
or U3679 (N_3679,N_878,N_1645);
or U3680 (N_3680,N_2174,N_407);
nor U3681 (N_3681,N_1248,N_2448);
xnor U3682 (N_3682,N_1787,N_1139);
xnor U3683 (N_3683,N_1675,N_1684);
and U3684 (N_3684,N_818,N_1430);
xor U3685 (N_3685,N_1405,N_333);
and U3686 (N_3686,N_533,N_1332);
and U3687 (N_3687,N_1014,N_1760);
nand U3688 (N_3688,N_1096,N_107);
nand U3689 (N_3689,N_401,N_634);
nand U3690 (N_3690,N_2389,N_1737);
nor U3691 (N_3691,N_2037,N_1878);
xor U3692 (N_3692,N_165,N_91);
or U3693 (N_3693,N_2430,N_2384);
or U3694 (N_3694,N_2454,N_1423);
nand U3695 (N_3695,N_869,N_2253);
nor U3696 (N_3696,N_1276,N_226);
and U3697 (N_3697,N_1160,N_1707);
nand U3698 (N_3698,N_1128,N_380);
or U3699 (N_3699,N_677,N_886);
xnor U3700 (N_3700,N_1558,N_1688);
xor U3701 (N_3701,N_524,N_1547);
nand U3702 (N_3702,N_690,N_1915);
or U3703 (N_3703,N_1620,N_1227);
and U3704 (N_3704,N_1396,N_1293);
nand U3705 (N_3705,N_88,N_1780);
xor U3706 (N_3706,N_644,N_971);
or U3707 (N_3707,N_961,N_1784);
and U3708 (N_3708,N_1745,N_834);
xor U3709 (N_3709,N_1700,N_1295);
or U3710 (N_3710,N_2367,N_437);
nor U3711 (N_3711,N_1369,N_1761);
and U3712 (N_3712,N_1781,N_2064);
and U3713 (N_3713,N_236,N_548);
xor U3714 (N_3714,N_2014,N_1140);
nand U3715 (N_3715,N_537,N_836);
xnor U3716 (N_3716,N_852,N_1322);
xnor U3717 (N_3717,N_723,N_1108);
and U3718 (N_3718,N_1914,N_1846);
or U3719 (N_3719,N_1556,N_1751);
and U3720 (N_3720,N_2118,N_1880);
nor U3721 (N_3721,N_1768,N_850);
xnor U3722 (N_3722,N_2087,N_979);
nand U3723 (N_3723,N_1714,N_538);
or U3724 (N_3724,N_876,N_1265);
xor U3725 (N_3725,N_1329,N_625);
and U3726 (N_3726,N_1476,N_253);
nor U3727 (N_3727,N_90,N_1739);
and U3728 (N_3728,N_550,N_1006);
nor U3729 (N_3729,N_148,N_552);
nand U3730 (N_3730,N_2460,N_558);
or U3731 (N_3731,N_2387,N_935);
or U3732 (N_3732,N_525,N_1793);
nor U3733 (N_3733,N_1732,N_1570);
and U3734 (N_3734,N_1274,N_214);
or U3735 (N_3735,N_411,N_1206);
nor U3736 (N_3736,N_1063,N_2211);
nand U3737 (N_3737,N_1964,N_421);
nand U3738 (N_3738,N_2063,N_1943);
nor U3739 (N_3739,N_200,N_705);
or U3740 (N_3740,N_955,N_887);
xor U3741 (N_3741,N_1918,N_1939);
nand U3742 (N_3742,N_578,N_278);
nand U3743 (N_3743,N_1885,N_1502);
nand U3744 (N_3744,N_1905,N_249);
or U3745 (N_3745,N_2346,N_1727);
xnor U3746 (N_3746,N_841,N_2123);
and U3747 (N_3747,N_488,N_1001);
nand U3748 (N_3748,N_2271,N_2161);
and U3749 (N_3749,N_339,N_341);
or U3750 (N_3750,N_692,N_2482);
nor U3751 (N_3751,N_712,N_2208);
or U3752 (N_3752,N_1752,N_1750);
nor U3753 (N_3753,N_989,N_312);
xnor U3754 (N_3754,N_490,N_1583);
nor U3755 (N_3755,N_1614,N_2282);
or U3756 (N_3756,N_750,N_1263);
nor U3757 (N_3757,N_2489,N_587);
nand U3758 (N_3758,N_1979,N_1985);
nor U3759 (N_3759,N_1209,N_247);
nand U3760 (N_3760,N_1378,N_1157);
or U3761 (N_3761,N_277,N_2050);
nor U3762 (N_3762,N_262,N_2275);
xnor U3763 (N_3763,N_1152,N_829);
or U3764 (N_3764,N_1063,N_319);
nand U3765 (N_3765,N_2122,N_718);
nor U3766 (N_3766,N_2168,N_760);
or U3767 (N_3767,N_780,N_2376);
and U3768 (N_3768,N_104,N_1560);
nand U3769 (N_3769,N_760,N_1359);
nand U3770 (N_3770,N_2386,N_2377);
nor U3771 (N_3771,N_1186,N_1048);
or U3772 (N_3772,N_2162,N_2211);
xor U3773 (N_3773,N_680,N_2074);
xnor U3774 (N_3774,N_1963,N_1597);
xor U3775 (N_3775,N_2271,N_433);
nor U3776 (N_3776,N_360,N_640);
nor U3777 (N_3777,N_1760,N_2048);
and U3778 (N_3778,N_1359,N_669);
or U3779 (N_3779,N_1524,N_2170);
nand U3780 (N_3780,N_1867,N_1315);
and U3781 (N_3781,N_525,N_1850);
or U3782 (N_3782,N_1612,N_622);
nor U3783 (N_3783,N_2399,N_1302);
xor U3784 (N_3784,N_1407,N_455);
nand U3785 (N_3785,N_963,N_2293);
nand U3786 (N_3786,N_374,N_1338);
nand U3787 (N_3787,N_2289,N_1906);
nand U3788 (N_3788,N_478,N_1583);
and U3789 (N_3789,N_136,N_1376);
nor U3790 (N_3790,N_2273,N_835);
nor U3791 (N_3791,N_115,N_633);
and U3792 (N_3792,N_1809,N_1004);
xnor U3793 (N_3793,N_34,N_1708);
and U3794 (N_3794,N_655,N_2487);
xnor U3795 (N_3795,N_1238,N_133);
nand U3796 (N_3796,N_1746,N_49);
xnor U3797 (N_3797,N_1276,N_2217);
xor U3798 (N_3798,N_2152,N_935);
xnor U3799 (N_3799,N_2241,N_999);
xor U3800 (N_3800,N_548,N_1334);
or U3801 (N_3801,N_450,N_495);
or U3802 (N_3802,N_2012,N_1124);
nand U3803 (N_3803,N_1440,N_2317);
xnor U3804 (N_3804,N_0,N_1821);
nand U3805 (N_3805,N_2100,N_729);
and U3806 (N_3806,N_603,N_975);
and U3807 (N_3807,N_344,N_1348);
nand U3808 (N_3808,N_1507,N_1673);
xnor U3809 (N_3809,N_363,N_138);
xor U3810 (N_3810,N_2096,N_1160);
and U3811 (N_3811,N_711,N_820);
nor U3812 (N_3812,N_1654,N_1533);
and U3813 (N_3813,N_2459,N_583);
nand U3814 (N_3814,N_1020,N_611);
nor U3815 (N_3815,N_917,N_108);
nand U3816 (N_3816,N_1777,N_738);
xnor U3817 (N_3817,N_2306,N_584);
nor U3818 (N_3818,N_943,N_582);
nor U3819 (N_3819,N_1570,N_2491);
or U3820 (N_3820,N_1041,N_1062);
and U3821 (N_3821,N_426,N_164);
or U3822 (N_3822,N_824,N_516);
nor U3823 (N_3823,N_1854,N_2140);
nor U3824 (N_3824,N_1109,N_762);
or U3825 (N_3825,N_1501,N_327);
or U3826 (N_3826,N_1713,N_1748);
nor U3827 (N_3827,N_513,N_1157);
xor U3828 (N_3828,N_1344,N_1879);
xnor U3829 (N_3829,N_762,N_943);
nand U3830 (N_3830,N_2413,N_50);
nor U3831 (N_3831,N_992,N_2478);
and U3832 (N_3832,N_450,N_551);
nor U3833 (N_3833,N_1976,N_1557);
and U3834 (N_3834,N_1529,N_863);
nand U3835 (N_3835,N_1655,N_38);
and U3836 (N_3836,N_215,N_382);
or U3837 (N_3837,N_917,N_208);
nand U3838 (N_3838,N_2333,N_969);
xor U3839 (N_3839,N_964,N_708);
or U3840 (N_3840,N_577,N_2158);
nand U3841 (N_3841,N_2362,N_1485);
xnor U3842 (N_3842,N_1299,N_1202);
nand U3843 (N_3843,N_1175,N_1049);
nor U3844 (N_3844,N_2330,N_2207);
xnor U3845 (N_3845,N_1045,N_1005);
xnor U3846 (N_3846,N_1692,N_175);
or U3847 (N_3847,N_2027,N_1454);
nand U3848 (N_3848,N_1441,N_1124);
xor U3849 (N_3849,N_1187,N_2336);
nor U3850 (N_3850,N_1354,N_1724);
xnor U3851 (N_3851,N_2397,N_1746);
xnor U3852 (N_3852,N_2133,N_490);
xnor U3853 (N_3853,N_48,N_466);
or U3854 (N_3854,N_754,N_1981);
nand U3855 (N_3855,N_2346,N_2345);
and U3856 (N_3856,N_1002,N_497);
or U3857 (N_3857,N_1601,N_796);
nor U3858 (N_3858,N_1114,N_521);
nor U3859 (N_3859,N_1619,N_1136);
nor U3860 (N_3860,N_351,N_115);
nand U3861 (N_3861,N_228,N_1830);
xor U3862 (N_3862,N_1076,N_1701);
nor U3863 (N_3863,N_1494,N_1397);
and U3864 (N_3864,N_1424,N_1723);
and U3865 (N_3865,N_1309,N_1594);
or U3866 (N_3866,N_1539,N_1653);
xor U3867 (N_3867,N_2347,N_1925);
or U3868 (N_3868,N_1225,N_1643);
or U3869 (N_3869,N_300,N_780);
or U3870 (N_3870,N_2406,N_1137);
and U3871 (N_3871,N_2068,N_1077);
or U3872 (N_3872,N_592,N_1129);
xnor U3873 (N_3873,N_230,N_565);
or U3874 (N_3874,N_2309,N_519);
xnor U3875 (N_3875,N_549,N_1695);
and U3876 (N_3876,N_2492,N_194);
or U3877 (N_3877,N_371,N_501);
nand U3878 (N_3878,N_74,N_732);
nor U3879 (N_3879,N_1739,N_912);
and U3880 (N_3880,N_1351,N_139);
xnor U3881 (N_3881,N_235,N_1907);
or U3882 (N_3882,N_2037,N_2095);
or U3883 (N_3883,N_782,N_1427);
and U3884 (N_3884,N_1532,N_477);
nand U3885 (N_3885,N_139,N_21);
nor U3886 (N_3886,N_981,N_2449);
nand U3887 (N_3887,N_966,N_465);
and U3888 (N_3888,N_839,N_2422);
and U3889 (N_3889,N_2293,N_365);
or U3890 (N_3890,N_1631,N_2365);
and U3891 (N_3891,N_51,N_206);
nor U3892 (N_3892,N_1401,N_1276);
nor U3893 (N_3893,N_1769,N_1718);
xnor U3894 (N_3894,N_1105,N_846);
and U3895 (N_3895,N_1532,N_363);
or U3896 (N_3896,N_1983,N_1937);
nand U3897 (N_3897,N_838,N_1842);
xor U3898 (N_3898,N_1002,N_1541);
and U3899 (N_3899,N_1834,N_648);
nand U3900 (N_3900,N_1197,N_669);
nand U3901 (N_3901,N_1408,N_1312);
and U3902 (N_3902,N_4,N_958);
nor U3903 (N_3903,N_406,N_228);
xnor U3904 (N_3904,N_348,N_594);
and U3905 (N_3905,N_262,N_2436);
and U3906 (N_3906,N_497,N_1882);
or U3907 (N_3907,N_1105,N_2107);
nor U3908 (N_3908,N_1339,N_1801);
nor U3909 (N_3909,N_672,N_910);
and U3910 (N_3910,N_1275,N_49);
or U3911 (N_3911,N_1064,N_77);
nand U3912 (N_3912,N_2139,N_362);
nor U3913 (N_3913,N_2389,N_664);
xor U3914 (N_3914,N_2417,N_1822);
xnor U3915 (N_3915,N_2388,N_293);
xor U3916 (N_3916,N_781,N_1052);
and U3917 (N_3917,N_1369,N_1002);
nand U3918 (N_3918,N_529,N_1747);
and U3919 (N_3919,N_553,N_716);
xor U3920 (N_3920,N_1642,N_807);
nor U3921 (N_3921,N_2178,N_1807);
and U3922 (N_3922,N_1669,N_1658);
nand U3923 (N_3923,N_792,N_1827);
nand U3924 (N_3924,N_143,N_1583);
nor U3925 (N_3925,N_1162,N_1593);
and U3926 (N_3926,N_304,N_1192);
xor U3927 (N_3927,N_499,N_232);
and U3928 (N_3928,N_1000,N_2385);
and U3929 (N_3929,N_121,N_2187);
and U3930 (N_3930,N_1931,N_797);
and U3931 (N_3931,N_390,N_2068);
xor U3932 (N_3932,N_38,N_2165);
xor U3933 (N_3933,N_667,N_514);
and U3934 (N_3934,N_702,N_1692);
nand U3935 (N_3935,N_315,N_1688);
or U3936 (N_3936,N_2454,N_987);
nor U3937 (N_3937,N_754,N_1859);
nor U3938 (N_3938,N_2037,N_1168);
nor U3939 (N_3939,N_2361,N_1646);
and U3940 (N_3940,N_2436,N_933);
nor U3941 (N_3941,N_835,N_1055);
nand U3942 (N_3942,N_1170,N_2305);
nand U3943 (N_3943,N_1071,N_1669);
and U3944 (N_3944,N_659,N_938);
xnor U3945 (N_3945,N_1363,N_2131);
and U3946 (N_3946,N_896,N_593);
or U3947 (N_3947,N_1059,N_980);
nor U3948 (N_3948,N_145,N_100);
or U3949 (N_3949,N_460,N_1366);
or U3950 (N_3950,N_2054,N_1742);
and U3951 (N_3951,N_1739,N_25);
nand U3952 (N_3952,N_2483,N_250);
xor U3953 (N_3953,N_2345,N_1017);
nor U3954 (N_3954,N_2105,N_1620);
and U3955 (N_3955,N_786,N_2322);
and U3956 (N_3956,N_1424,N_18);
xor U3957 (N_3957,N_1301,N_880);
xor U3958 (N_3958,N_71,N_443);
nor U3959 (N_3959,N_2454,N_811);
xor U3960 (N_3960,N_384,N_1782);
xor U3961 (N_3961,N_315,N_645);
or U3962 (N_3962,N_2080,N_1196);
nor U3963 (N_3963,N_435,N_1762);
nand U3964 (N_3964,N_642,N_450);
nand U3965 (N_3965,N_1071,N_2053);
or U3966 (N_3966,N_1343,N_888);
nor U3967 (N_3967,N_2420,N_869);
or U3968 (N_3968,N_1748,N_914);
and U3969 (N_3969,N_2338,N_1089);
nand U3970 (N_3970,N_264,N_2127);
xor U3971 (N_3971,N_1609,N_2482);
nand U3972 (N_3972,N_674,N_1810);
xor U3973 (N_3973,N_1793,N_412);
nor U3974 (N_3974,N_1192,N_855);
xnor U3975 (N_3975,N_274,N_174);
or U3976 (N_3976,N_1837,N_1083);
xor U3977 (N_3977,N_913,N_767);
or U3978 (N_3978,N_1824,N_2390);
and U3979 (N_3979,N_2185,N_2358);
or U3980 (N_3980,N_2395,N_666);
or U3981 (N_3981,N_654,N_1930);
nor U3982 (N_3982,N_840,N_1742);
and U3983 (N_3983,N_1562,N_2483);
xnor U3984 (N_3984,N_967,N_1651);
xnor U3985 (N_3985,N_2439,N_1883);
and U3986 (N_3986,N_1933,N_2174);
xor U3987 (N_3987,N_1037,N_391);
nand U3988 (N_3988,N_1971,N_1394);
nor U3989 (N_3989,N_1984,N_2293);
nand U3990 (N_3990,N_1033,N_251);
nand U3991 (N_3991,N_133,N_554);
and U3992 (N_3992,N_1349,N_2063);
or U3993 (N_3993,N_2269,N_1007);
and U3994 (N_3994,N_346,N_1573);
nor U3995 (N_3995,N_1861,N_0);
xor U3996 (N_3996,N_2205,N_89);
or U3997 (N_3997,N_1793,N_127);
nor U3998 (N_3998,N_1047,N_1044);
nand U3999 (N_3999,N_614,N_289);
or U4000 (N_4000,N_695,N_1041);
or U4001 (N_4001,N_1322,N_2054);
xnor U4002 (N_4002,N_829,N_1960);
and U4003 (N_4003,N_385,N_1176);
xor U4004 (N_4004,N_629,N_1585);
xor U4005 (N_4005,N_1926,N_815);
nand U4006 (N_4006,N_228,N_221);
xor U4007 (N_4007,N_1362,N_1049);
xnor U4008 (N_4008,N_1144,N_890);
nand U4009 (N_4009,N_271,N_916);
or U4010 (N_4010,N_1317,N_2256);
or U4011 (N_4011,N_1101,N_1333);
nor U4012 (N_4012,N_1825,N_1621);
xnor U4013 (N_4013,N_2388,N_2236);
nand U4014 (N_4014,N_477,N_1287);
xor U4015 (N_4015,N_947,N_2073);
or U4016 (N_4016,N_918,N_135);
or U4017 (N_4017,N_2146,N_425);
and U4018 (N_4018,N_1418,N_1349);
nor U4019 (N_4019,N_1262,N_2490);
nor U4020 (N_4020,N_2103,N_2386);
nor U4021 (N_4021,N_369,N_2227);
nand U4022 (N_4022,N_796,N_1584);
xor U4023 (N_4023,N_2085,N_2334);
or U4024 (N_4024,N_2234,N_44);
or U4025 (N_4025,N_2040,N_508);
nor U4026 (N_4026,N_1439,N_1360);
and U4027 (N_4027,N_1859,N_27);
or U4028 (N_4028,N_1917,N_994);
nor U4029 (N_4029,N_2312,N_1222);
nand U4030 (N_4030,N_367,N_192);
nand U4031 (N_4031,N_1351,N_1277);
xnor U4032 (N_4032,N_1754,N_1067);
xnor U4033 (N_4033,N_1155,N_2163);
and U4034 (N_4034,N_900,N_1441);
xnor U4035 (N_4035,N_165,N_640);
or U4036 (N_4036,N_779,N_1410);
or U4037 (N_4037,N_556,N_2328);
xnor U4038 (N_4038,N_2436,N_366);
or U4039 (N_4039,N_467,N_2323);
nand U4040 (N_4040,N_1945,N_2077);
nand U4041 (N_4041,N_2118,N_846);
nor U4042 (N_4042,N_41,N_2294);
nor U4043 (N_4043,N_2224,N_1327);
nand U4044 (N_4044,N_1943,N_986);
nand U4045 (N_4045,N_2217,N_2471);
or U4046 (N_4046,N_765,N_2441);
nand U4047 (N_4047,N_2366,N_179);
nor U4048 (N_4048,N_748,N_1100);
nand U4049 (N_4049,N_257,N_2246);
and U4050 (N_4050,N_1153,N_299);
xnor U4051 (N_4051,N_124,N_2315);
and U4052 (N_4052,N_1364,N_958);
nand U4053 (N_4053,N_1868,N_1701);
xnor U4054 (N_4054,N_537,N_534);
and U4055 (N_4055,N_903,N_1826);
or U4056 (N_4056,N_1816,N_2176);
and U4057 (N_4057,N_1036,N_649);
nand U4058 (N_4058,N_2388,N_2386);
nand U4059 (N_4059,N_10,N_1181);
nor U4060 (N_4060,N_1008,N_1016);
nand U4061 (N_4061,N_487,N_1659);
and U4062 (N_4062,N_2241,N_800);
or U4063 (N_4063,N_536,N_1962);
nor U4064 (N_4064,N_1772,N_1844);
nor U4065 (N_4065,N_2121,N_937);
xor U4066 (N_4066,N_1672,N_1497);
and U4067 (N_4067,N_242,N_1053);
nand U4068 (N_4068,N_1592,N_460);
nor U4069 (N_4069,N_1850,N_2431);
xnor U4070 (N_4070,N_1348,N_1201);
nor U4071 (N_4071,N_115,N_983);
xnor U4072 (N_4072,N_910,N_1597);
or U4073 (N_4073,N_48,N_2496);
nor U4074 (N_4074,N_1038,N_2032);
nor U4075 (N_4075,N_2188,N_189);
nand U4076 (N_4076,N_2288,N_807);
and U4077 (N_4077,N_1503,N_19);
nor U4078 (N_4078,N_1718,N_1714);
nor U4079 (N_4079,N_908,N_2333);
nor U4080 (N_4080,N_521,N_28);
and U4081 (N_4081,N_468,N_436);
and U4082 (N_4082,N_459,N_2239);
nor U4083 (N_4083,N_183,N_2002);
xnor U4084 (N_4084,N_1012,N_893);
xor U4085 (N_4085,N_106,N_1369);
nor U4086 (N_4086,N_2052,N_959);
nor U4087 (N_4087,N_970,N_1565);
and U4088 (N_4088,N_2378,N_403);
or U4089 (N_4089,N_2030,N_178);
nand U4090 (N_4090,N_218,N_1417);
or U4091 (N_4091,N_1082,N_1029);
nand U4092 (N_4092,N_477,N_1742);
nor U4093 (N_4093,N_2225,N_1337);
nor U4094 (N_4094,N_315,N_1974);
xnor U4095 (N_4095,N_91,N_2305);
xor U4096 (N_4096,N_1989,N_367);
nor U4097 (N_4097,N_2072,N_1346);
nand U4098 (N_4098,N_672,N_270);
and U4099 (N_4099,N_74,N_174);
nand U4100 (N_4100,N_119,N_575);
or U4101 (N_4101,N_840,N_2203);
nor U4102 (N_4102,N_887,N_1960);
nand U4103 (N_4103,N_2169,N_119);
and U4104 (N_4104,N_1962,N_394);
nand U4105 (N_4105,N_2407,N_1271);
or U4106 (N_4106,N_723,N_791);
xnor U4107 (N_4107,N_714,N_2265);
and U4108 (N_4108,N_852,N_94);
and U4109 (N_4109,N_106,N_1279);
xnor U4110 (N_4110,N_369,N_1443);
or U4111 (N_4111,N_199,N_546);
xor U4112 (N_4112,N_1032,N_212);
nand U4113 (N_4113,N_307,N_1092);
xnor U4114 (N_4114,N_1309,N_2470);
and U4115 (N_4115,N_1729,N_2023);
nor U4116 (N_4116,N_460,N_1734);
xor U4117 (N_4117,N_1085,N_538);
nand U4118 (N_4118,N_160,N_2351);
and U4119 (N_4119,N_601,N_2212);
xnor U4120 (N_4120,N_1526,N_691);
and U4121 (N_4121,N_1327,N_1400);
nor U4122 (N_4122,N_681,N_2127);
and U4123 (N_4123,N_1294,N_229);
nor U4124 (N_4124,N_2451,N_41);
and U4125 (N_4125,N_1849,N_2423);
nand U4126 (N_4126,N_2,N_2146);
nor U4127 (N_4127,N_262,N_1983);
nand U4128 (N_4128,N_1127,N_259);
or U4129 (N_4129,N_116,N_2101);
and U4130 (N_4130,N_2381,N_915);
nor U4131 (N_4131,N_1962,N_2345);
nand U4132 (N_4132,N_486,N_1623);
or U4133 (N_4133,N_456,N_388);
nor U4134 (N_4134,N_1725,N_2025);
xor U4135 (N_4135,N_1362,N_2389);
and U4136 (N_4136,N_2234,N_2289);
nand U4137 (N_4137,N_449,N_647);
xnor U4138 (N_4138,N_729,N_376);
or U4139 (N_4139,N_772,N_1308);
nand U4140 (N_4140,N_696,N_777);
nor U4141 (N_4141,N_749,N_245);
or U4142 (N_4142,N_1057,N_2211);
and U4143 (N_4143,N_1213,N_92);
or U4144 (N_4144,N_765,N_2311);
nor U4145 (N_4145,N_1443,N_1751);
nand U4146 (N_4146,N_433,N_11);
xor U4147 (N_4147,N_1408,N_508);
nand U4148 (N_4148,N_1845,N_40);
and U4149 (N_4149,N_1684,N_1282);
nand U4150 (N_4150,N_1051,N_465);
nand U4151 (N_4151,N_1144,N_455);
xor U4152 (N_4152,N_2113,N_768);
xnor U4153 (N_4153,N_1686,N_490);
xnor U4154 (N_4154,N_1759,N_572);
nand U4155 (N_4155,N_2472,N_2397);
nand U4156 (N_4156,N_2331,N_1549);
nor U4157 (N_4157,N_132,N_413);
nor U4158 (N_4158,N_1741,N_475);
and U4159 (N_4159,N_1682,N_787);
and U4160 (N_4160,N_980,N_182);
nand U4161 (N_4161,N_565,N_1641);
and U4162 (N_4162,N_1857,N_1493);
or U4163 (N_4163,N_694,N_1070);
xnor U4164 (N_4164,N_972,N_2135);
or U4165 (N_4165,N_1497,N_1383);
nand U4166 (N_4166,N_23,N_2429);
and U4167 (N_4167,N_2261,N_1134);
xor U4168 (N_4168,N_374,N_22);
xor U4169 (N_4169,N_461,N_1264);
and U4170 (N_4170,N_1232,N_1517);
and U4171 (N_4171,N_679,N_2380);
nor U4172 (N_4172,N_503,N_1449);
xor U4173 (N_4173,N_416,N_386);
nand U4174 (N_4174,N_1848,N_502);
or U4175 (N_4175,N_1877,N_310);
and U4176 (N_4176,N_929,N_101);
and U4177 (N_4177,N_1394,N_2219);
and U4178 (N_4178,N_1704,N_515);
nor U4179 (N_4179,N_135,N_1248);
nand U4180 (N_4180,N_1065,N_131);
xnor U4181 (N_4181,N_1461,N_124);
nand U4182 (N_4182,N_1710,N_152);
xor U4183 (N_4183,N_2116,N_2295);
nor U4184 (N_4184,N_1631,N_1344);
nand U4185 (N_4185,N_131,N_161);
and U4186 (N_4186,N_675,N_848);
or U4187 (N_4187,N_429,N_2436);
nor U4188 (N_4188,N_1985,N_1639);
or U4189 (N_4189,N_2256,N_1227);
or U4190 (N_4190,N_998,N_1044);
nor U4191 (N_4191,N_259,N_1527);
nand U4192 (N_4192,N_1927,N_1567);
xnor U4193 (N_4193,N_902,N_1072);
nand U4194 (N_4194,N_2150,N_2246);
or U4195 (N_4195,N_1397,N_1037);
xor U4196 (N_4196,N_635,N_1995);
xnor U4197 (N_4197,N_1163,N_2394);
and U4198 (N_4198,N_154,N_320);
xor U4199 (N_4199,N_896,N_1869);
xor U4200 (N_4200,N_399,N_1972);
or U4201 (N_4201,N_1943,N_1489);
and U4202 (N_4202,N_35,N_2032);
nand U4203 (N_4203,N_1183,N_316);
xor U4204 (N_4204,N_1077,N_611);
or U4205 (N_4205,N_974,N_1307);
or U4206 (N_4206,N_1799,N_932);
or U4207 (N_4207,N_1439,N_848);
nand U4208 (N_4208,N_1770,N_1258);
or U4209 (N_4209,N_1987,N_624);
or U4210 (N_4210,N_326,N_2111);
and U4211 (N_4211,N_1172,N_749);
nand U4212 (N_4212,N_1583,N_862);
and U4213 (N_4213,N_2012,N_205);
and U4214 (N_4214,N_487,N_1169);
nand U4215 (N_4215,N_2263,N_1863);
nand U4216 (N_4216,N_619,N_1825);
xor U4217 (N_4217,N_1213,N_54);
and U4218 (N_4218,N_1067,N_2047);
nor U4219 (N_4219,N_825,N_1600);
or U4220 (N_4220,N_1593,N_1873);
nor U4221 (N_4221,N_2415,N_2382);
xnor U4222 (N_4222,N_66,N_1851);
nor U4223 (N_4223,N_2122,N_2495);
or U4224 (N_4224,N_2467,N_1708);
nand U4225 (N_4225,N_1343,N_2006);
nand U4226 (N_4226,N_105,N_1865);
xnor U4227 (N_4227,N_491,N_947);
and U4228 (N_4228,N_345,N_2197);
or U4229 (N_4229,N_221,N_2184);
nand U4230 (N_4230,N_2023,N_457);
and U4231 (N_4231,N_380,N_1792);
and U4232 (N_4232,N_2443,N_1315);
or U4233 (N_4233,N_1063,N_1822);
xnor U4234 (N_4234,N_518,N_2064);
and U4235 (N_4235,N_220,N_634);
and U4236 (N_4236,N_2130,N_1540);
and U4237 (N_4237,N_955,N_900);
nand U4238 (N_4238,N_456,N_895);
xnor U4239 (N_4239,N_1557,N_1521);
xor U4240 (N_4240,N_1328,N_2341);
nor U4241 (N_4241,N_1835,N_803);
and U4242 (N_4242,N_54,N_1732);
nor U4243 (N_4243,N_140,N_708);
nand U4244 (N_4244,N_814,N_2348);
nor U4245 (N_4245,N_1395,N_484);
or U4246 (N_4246,N_700,N_511);
nor U4247 (N_4247,N_1508,N_1674);
or U4248 (N_4248,N_720,N_197);
xnor U4249 (N_4249,N_1419,N_477);
or U4250 (N_4250,N_1951,N_1915);
nand U4251 (N_4251,N_792,N_2335);
or U4252 (N_4252,N_505,N_1562);
or U4253 (N_4253,N_1887,N_1769);
xor U4254 (N_4254,N_1238,N_2298);
or U4255 (N_4255,N_408,N_339);
nor U4256 (N_4256,N_76,N_1991);
nor U4257 (N_4257,N_1319,N_1648);
nand U4258 (N_4258,N_1328,N_525);
nor U4259 (N_4259,N_2494,N_401);
and U4260 (N_4260,N_1602,N_1912);
nor U4261 (N_4261,N_2364,N_883);
or U4262 (N_4262,N_2398,N_1277);
and U4263 (N_4263,N_1163,N_2078);
nor U4264 (N_4264,N_1102,N_1290);
nor U4265 (N_4265,N_201,N_1045);
xor U4266 (N_4266,N_2430,N_2221);
xor U4267 (N_4267,N_1322,N_1464);
or U4268 (N_4268,N_1126,N_673);
xnor U4269 (N_4269,N_654,N_1375);
nand U4270 (N_4270,N_585,N_1922);
or U4271 (N_4271,N_2156,N_2103);
xnor U4272 (N_4272,N_398,N_1272);
nand U4273 (N_4273,N_376,N_594);
nand U4274 (N_4274,N_1253,N_1133);
nor U4275 (N_4275,N_2298,N_301);
nand U4276 (N_4276,N_2492,N_368);
nand U4277 (N_4277,N_969,N_91);
nand U4278 (N_4278,N_164,N_1550);
or U4279 (N_4279,N_2362,N_1923);
or U4280 (N_4280,N_46,N_306);
nand U4281 (N_4281,N_94,N_508);
nand U4282 (N_4282,N_2295,N_1394);
xor U4283 (N_4283,N_309,N_2154);
nor U4284 (N_4284,N_140,N_2317);
nand U4285 (N_4285,N_1196,N_982);
nor U4286 (N_4286,N_423,N_1793);
nor U4287 (N_4287,N_993,N_1564);
nand U4288 (N_4288,N_1026,N_2308);
or U4289 (N_4289,N_1110,N_2238);
nand U4290 (N_4290,N_1941,N_693);
nor U4291 (N_4291,N_1083,N_2284);
and U4292 (N_4292,N_1267,N_234);
or U4293 (N_4293,N_469,N_451);
or U4294 (N_4294,N_890,N_655);
or U4295 (N_4295,N_360,N_1587);
and U4296 (N_4296,N_652,N_2349);
nand U4297 (N_4297,N_1262,N_272);
and U4298 (N_4298,N_565,N_248);
and U4299 (N_4299,N_1056,N_1960);
or U4300 (N_4300,N_1037,N_1273);
nand U4301 (N_4301,N_597,N_2407);
nand U4302 (N_4302,N_1847,N_287);
or U4303 (N_4303,N_1072,N_2468);
xnor U4304 (N_4304,N_1221,N_229);
and U4305 (N_4305,N_1760,N_2388);
nand U4306 (N_4306,N_320,N_737);
and U4307 (N_4307,N_1441,N_2004);
xnor U4308 (N_4308,N_191,N_1515);
nand U4309 (N_4309,N_2227,N_1832);
nand U4310 (N_4310,N_705,N_2425);
nand U4311 (N_4311,N_1781,N_977);
nand U4312 (N_4312,N_1847,N_312);
nor U4313 (N_4313,N_100,N_1500);
xor U4314 (N_4314,N_1378,N_774);
nand U4315 (N_4315,N_1575,N_1170);
xnor U4316 (N_4316,N_2000,N_111);
xnor U4317 (N_4317,N_882,N_2494);
or U4318 (N_4318,N_1958,N_302);
nand U4319 (N_4319,N_1064,N_483);
xor U4320 (N_4320,N_66,N_2041);
nor U4321 (N_4321,N_124,N_1149);
nand U4322 (N_4322,N_2386,N_2124);
xor U4323 (N_4323,N_706,N_520);
or U4324 (N_4324,N_2101,N_1510);
xor U4325 (N_4325,N_1960,N_1472);
and U4326 (N_4326,N_184,N_2407);
nand U4327 (N_4327,N_1865,N_180);
nor U4328 (N_4328,N_2249,N_130);
and U4329 (N_4329,N_1665,N_1735);
nand U4330 (N_4330,N_94,N_2064);
nand U4331 (N_4331,N_1244,N_2232);
nand U4332 (N_4332,N_1949,N_460);
or U4333 (N_4333,N_696,N_1749);
or U4334 (N_4334,N_2494,N_929);
nand U4335 (N_4335,N_1464,N_81);
xor U4336 (N_4336,N_1,N_2252);
or U4337 (N_4337,N_461,N_2180);
nand U4338 (N_4338,N_403,N_597);
or U4339 (N_4339,N_1921,N_1839);
and U4340 (N_4340,N_379,N_647);
or U4341 (N_4341,N_1854,N_2184);
or U4342 (N_4342,N_1039,N_127);
xnor U4343 (N_4343,N_1556,N_1846);
xnor U4344 (N_4344,N_1523,N_1959);
and U4345 (N_4345,N_1089,N_541);
nor U4346 (N_4346,N_1705,N_1850);
or U4347 (N_4347,N_554,N_1027);
nor U4348 (N_4348,N_1370,N_2115);
xor U4349 (N_4349,N_664,N_2338);
and U4350 (N_4350,N_1947,N_64);
and U4351 (N_4351,N_812,N_2446);
nor U4352 (N_4352,N_2044,N_1836);
xor U4353 (N_4353,N_2303,N_1581);
xor U4354 (N_4354,N_1753,N_1939);
or U4355 (N_4355,N_868,N_2130);
nand U4356 (N_4356,N_2419,N_685);
xnor U4357 (N_4357,N_1413,N_1119);
and U4358 (N_4358,N_1191,N_1458);
or U4359 (N_4359,N_257,N_1005);
or U4360 (N_4360,N_778,N_1066);
nor U4361 (N_4361,N_619,N_1723);
or U4362 (N_4362,N_459,N_1869);
xnor U4363 (N_4363,N_1871,N_1387);
nand U4364 (N_4364,N_1748,N_1848);
xor U4365 (N_4365,N_1717,N_1901);
nand U4366 (N_4366,N_1334,N_1360);
nor U4367 (N_4367,N_1392,N_101);
nor U4368 (N_4368,N_270,N_2366);
nand U4369 (N_4369,N_401,N_1486);
xnor U4370 (N_4370,N_892,N_1297);
or U4371 (N_4371,N_351,N_1411);
nand U4372 (N_4372,N_2459,N_2136);
and U4373 (N_4373,N_820,N_744);
or U4374 (N_4374,N_2435,N_1217);
nand U4375 (N_4375,N_1573,N_838);
nand U4376 (N_4376,N_2488,N_1905);
or U4377 (N_4377,N_882,N_146);
and U4378 (N_4378,N_1238,N_691);
xnor U4379 (N_4379,N_1013,N_622);
nand U4380 (N_4380,N_701,N_840);
xor U4381 (N_4381,N_447,N_1989);
nor U4382 (N_4382,N_1754,N_1702);
and U4383 (N_4383,N_522,N_204);
or U4384 (N_4384,N_1211,N_2212);
and U4385 (N_4385,N_699,N_164);
xor U4386 (N_4386,N_2222,N_525);
or U4387 (N_4387,N_378,N_1332);
nand U4388 (N_4388,N_1888,N_2246);
nor U4389 (N_4389,N_642,N_1306);
nor U4390 (N_4390,N_1402,N_1);
nand U4391 (N_4391,N_180,N_208);
nor U4392 (N_4392,N_1138,N_538);
and U4393 (N_4393,N_1683,N_2427);
and U4394 (N_4394,N_2075,N_1286);
xnor U4395 (N_4395,N_1970,N_1928);
or U4396 (N_4396,N_1877,N_1022);
nand U4397 (N_4397,N_465,N_192);
nand U4398 (N_4398,N_1225,N_1290);
and U4399 (N_4399,N_938,N_1063);
nand U4400 (N_4400,N_1942,N_612);
nand U4401 (N_4401,N_1563,N_617);
nor U4402 (N_4402,N_1033,N_1317);
and U4403 (N_4403,N_653,N_1415);
or U4404 (N_4404,N_1226,N_835);
nand U4405 (N_4405,N_2085,N_886);
nor U4406 (N_4406,N_221,N_938);
nand U4407 (N_4407,N_329,N_181);
nor U4408 (N_4408,N_1811,N_1226);
nand U4409 (N_4409,N_1700,N_197);
nand U4410 (N_4410,N_145,N_1658);
nor U4411 (N_4411,N_1407,N_1367);
xnor U4412 (N_4412,N_1307,N_1031);
xor U4413 (N_4413,N_1080,N_739);
and U4414 (N_4414,N_1097,N_30);
and U4415 (N_4415,N_1421,N_2395);
xnor U4416 (N_4416,N_1532,N_1528);
and U4417 (N_4417,N_2344,N_351);
or U4418 (N_4418,N_936,N_79);
nor U4419 (N_4419,N_1728,N_2143);
or U4420 (N_4420,N_1206,N_230);
xor U4421 (N_4421,N_2446,N_1573);
nor U4422 (N_4422,N_205,N_2084);
nand U4423 (N_4423,N_571,N_664);
nand U4424 (N_4424,N_875,N_1818);
xnor U4425 (N_4425,N_167,N_1847);
nand U4426 (N_4426,N_877,N_664);
and U4427 (N_4427,N_825,N_1649);
nand U4428 (N_4428,N_1943,N_2461);
nor U4429 (N_4429,N_71,N_1093);
and U4430 (N_4430,N_85,N_827);
nor U4431 (N_4431,N_1219,N_387);
and U4432 (N_4432,N_1588,N_1375);
xor U4433 (N_4433,N_812,N_1214);
and U4434 (N_4434,N_503,N_2443);
xnor U4435 (N_4435,N_964,N_189);
nor U4436 (N_4436,N_202,N_2241);
nand U4437 (N_4437,N_2048,N_1763);
or U4438 (N_4438,N_624,N_283);
and U4439 (N_4439,N_1628,N_739);
and U4440 (N_4440,N_857,N_2180);
xnor U4441 (N_4441,N_1260,N_467);
nor U4442 (N_4442,N_1059,N_1167);
nor U4443 (N_4443,N_1487,N_1999);
or U4444 (N_4444,N_62,N_619);
xnor U4445 (N_4445,N_2268,N_678);
nor U4446 (N_4446,N_2196,N_2370);
and U4447 (N_4447,N_1004,N_935);
or U4448 (N_4448,N_1026,N_1170);
xor U4449 (N_4449,N_614,N_584);
xnor U4450 (N_4450,N_1159,N_1059);
and U4451 (N_4451,N_1933,N_1939);
nor U4452 (N_4452,N_1937,N_2313);
nand U4453 (N_4453,N_1672,N_1316);
xnor U4454 (N_4454,N_2481,N_1784);
nor U4455 (N_4455,N_816,N_1604);
and U4456 (N_4456,N_119,N_1574);
xnor U4457 (N_4457,N_1589,N_2023);
or U4458 (N_4458,N_998,N_915);
nand U4459 (N_4459,N_366,N_595);
and U4460 (N_4460,N_743,N_1172);
nor U4461 (N_4461,N_2468,N_2325);
nor U4462 (N_4462,N_2143,N_1724);
xor U4463 (N_4463,N_181,N_1986);
nor U4464 (N_4464,N_1414,N_1786);
and U4465 (N_4465,N_993,N_1914);
nand U4466 (N_4466,N_1348,N_92);
xor U4467 (N_4467,N_1955,N_1466);
or U4468 (N_4468,N_1692,N_253);
nand U4469 (N_4469,N_1481,N_405);
or U4470 (N_4470,N_2268,N_493);
nor U4471 (N_4471,N_452,N_291);
nor U4472 (N_4472,N_2173,N_116);
or U4473 (N_4473,N_4,N_1033);
xnor U4474 (N_4474,N_2379,N_392);
and U4475 (N_4475,N_477,N_78);
nor U4476 (N_4476,N_1218,N_61);
xnor U4477 (N_4477,N_2261,N_42);
xnor U4478 (N_4478,N_1746,N_856);
nor U4479 (N_4479,N_710,N_94);
xor U4480 (N_4480,N_633,N_284);
and U4481 (N_4481,N_1353,N_824);
xnor U4482 (N_4482,N_3,N_2453);
nand U4483 (N_4483,N_1255,N_535);
nor U4484 (N_4484,N_1021,N_677);
nor U4485 (N_4485,N_788,N_2165);
nand U4486 (N_4486,N_35,N_1342);
nand U4487 (N_4487,N_1156,N_724);
or U4488 (N_4488,N_679,N_58);
or U4489 (N_4489,N_2292,N_1354);
or U4490 (N_4490,N_230,N_2492);
nand U4491 (N_4491,N_1142,N_1993);
and U4492 (N_4492,N_2486,N_1783);
or U4493 (N_4493,N_1777,N_221);
or U4494 (N_4494,N_1822,N_2286);
nand U4495 (N_4495,N_1574,N_1164);
and U4496 (N_4496,N_1183,N_1260);
nor U4497 (N_4497,N_1416,N_1545);
nand U4498 (N_4498,N_90,N_622);
nor U4499 (N_4499,N_1939,N_1974);
xnor U4500 (N_4500,N_1791,N_1159);
xnor U4501 (N_4501,N_1759,N_1751);
and U4502 (N_4502,N_508,N_237);
xor U4503 (N_4503,N_1760,N_184);
and U4504 (N_4504,N_2128,N_1018);
nand U4505 (N_4505,N_2421,N_1489);
nand U4506 (N_4506,N_1722,N_2122);
xor U4507 (N_4507,N_745,N_183);
xnor U4508 (N_4508,N_438,N_1179);
and U4509 (N_4509,N_2138,N_827);
or U4510 (N_4510,N_533,N_471);
xor U4511 (N_4511,N_446,N_2028);
or U4512 (N_4512,N_2159,N_450);
and U4513 (N_4513,N_14,N_560);
or U4514 (N_4514,N_427,N_756);
and U4515 (N_4515,N_921,N_1941);
nor U4516 (N_4516,N_1731,N_647);
and U4517 (N_4517,N_1319,N_2267);
nand U4518 (N_4518,N_485,N_985);
nand U4519 (N_4519,N_1369,N_877);
nand U4520 (N_4520,N_581,N_504);
nand U4521 (N_4521,N_1269,N_208);
nor U4522 (N_4522,N_444,N_1276);
or U4523 (N_4523,N_410,N_27);
or U4524 (N_4524,N_435,N_1218);
xnor U4525 (N_4525,N_495,N_2377);
nand U4526 (N_4526,N_394,N_353);
or U4527 (N_4527,N_323,N_334);
and U4528 (N_4528,N_1540,N_1156);
or U4529 (N_4529,N_484,N_1480);
nor U4530 (N_4530,N_355,N_1604);
nor U4531 (N_4531,N_1566,N_1164);
nor U4532 (N_4532,N_2187,N_1580);
xnor U4533 (N_4533,N_2020,N_2064);
or U4534 (N_4534,N_2087,N_2088);
or U4535 (N_4535,N_1338,N_754);
nor U4536 (N_4536,N_904,N_1859);
nor U4537 (N_4537,N_1444,N_2037);
xnor U4538 (N_4538,N_533,N_453);
nor U4539 (N_4539,N_1948,N_173);
nand U4540 (N_4540,N_365,N_1959);
and U4541 (N_4541,N_388,N_834);
nor U4542 (N_4542,N_593,N_1529);
xor U4543 (N_4543,N_2028,N_1050);
or U4544 (N_4544,N_625,N_2101);
and U4545 (N_4545,N_686,N_1035);
and U4546 (N_4546,N_1848,N_2008);
xnor U4547 (N_4547,N_1610,N_1118);
xor U4548 (N_4548,N_1549,N_1071);
or U4549 (N_4549,N_2475,N_401);
nand U4550 (N_4550,N_2341,N_68);
and U4551 (N_4551,N_2430,N_1190);
nor U4552 (N_4552,N_270,N_1223);
xnor U4553 (N_4553,N_33,N_928);
and U4554 (N_4554,N_1810,N_2186);
nand U4555 (N_4555,N_384,N_391);
nand U4556 (N_4556,N_2094,N_2265);
nand U4557 (N_4557,N_1726,N_1982);
xnor U4558 (N_4558,N_1301,N_2187);
and U4559 (N_4559,N_2000,N_500);
xnor U4560 (N_4560,N_292,N_1519);
nor U4561 (N_4561,N_702,N_536);
and U4562 (N_4562,N_157,N_1349);
nor U4563 (N_4563,N_2121,N_1746);
and U4564 (N_4564,N_105,N_679);
nor U4565 (N_4565,N_2109,N_1311);
nor U4566 (N_4566,N_1509,N_2317);
or U4567 (N_4567,N_2481,N_686);
nor U4568 (N_4568,N_1743,N_1355);
or U4569 (N_4569,N_1756,N_1853);
nor U4570 (N_4570,N_36,N_1343);
nand U4571 (N_4571,N_1091,N_829);
and U4572 (N_4572,N_155,N_1721);
nor U4573 (N_4573,N_22,N_2132);
and U4574 (N_4574,N_413,N_1779);
nor U4575 (N_4575,N_1376,N_2002);
xnor U4576 (N_4576,N_2159,N_229);
xnor U4577 (N_4577,N_2331,N_1593);
and U4578 (N_4578,N_2221,N_1912);
xor U4579 (N_4579,N_989,N_2051);
and U4580 (N_4580,N_1413,N_1095);
or U4581 (N_4581,N_712,N_1013);
xor U4582 (N_4582,N_464,N_1952);
nand U4583 (N_4583,N_2327,N_2082);
nor U4584 (N_4584,N_545,N_1120);
or U4585 (N_4585,N_1932,N_226);
nand U4586 (N_4586,N_92,N_709);
and U4587 (N_4587,N_899,N_1237);
nor U4588 (N_4588,N_2097,N_781);
or U4589 (N_4589,N_1186,N_2308);
nor U4590 (N_4590,N_1845,N_1027);
xor U4591 (N_4591,N_744,N_1309);
nand U4592 (N_4592,N_1467,N_1870);
nand U4593 (N_4593,N_404,N_1818);
and U4594 (N_4594,N_354,N_1824);
or U4595 (N_4595,N_1509,N_1670);
xnor U4596 (N_4596,N_2250,N_1240);
and U4597 (N_4597,N_2368,N_1062);
xor U4598 (N_4598,N_1002,N_2386);
or U4599 (N_4599,N_907,N_1130);
nand U4600 (N_4600,N_855,N_203);
nand U4601 (N_4601,N_710,N_171);
and U4602 (N_4602,N_1026,N_984);
or U4603 (N_4603,N_424,N_1807);
nor U4604 (N_4604,N_2183,N_1715);
nand U4605 (N_4605,N_663,N_113);
xor U4606 (N_4606,N_2036,N_358);
xor U4607 (N_4607,N_335,N_2027);
nor U4608 (N_4608,N_2308,N_2057);
nand U4609 (N_4609,N_1242,N_1147);
xor U4610 (N_4610,N_507,N_2435);
or U4611 (N_4611,N_2249,N_1520);
nor U4612 (N_4612,N_62,N_597);
or U4613 (N_4613,N_352,N_2131);
nor U4614 (N_4614,N_1088,N_2395);
and U4615 (N_4615,N_1896,N_2360);
or U4616 (N_4616,N_1760,N_1904);
xor U4617 (N_4617,N_800,N_163);
or U4618 (N_4618,N_431,N_42);
or U4619 (N_4619,N_532,N_18);
and U4620 (N_4620,N_307,N_2001);
and U4621 (N_4621,N_2128,N_1025);
nor U4622 (N_4622,N_1898,N_2009);
or U4623 (N_4623,N_1114,N_1495);
xnor U4624 (N_4624,N_917,N_2482);
or U4625 (N_4625,N_2035,N_2258);
nor U4626 (N_4626,N_1225,N_1491);
nor U4627 (N_4627,N_748,N_306);
nand U4628 (N_4628,N_1431,N_1464);
nor U4629 (N_4629,N_2052,N_942);
nand U4630 (N_4630,N_570,N_2478);
nand U4631 (N_4631,N_307,N_566);
and U4632 (N_4632,N_2380,N_1975);
nor U4633 (N_4633,N_814,N_2223);
or U4634 (N_4634,N_1641,N_944);
xor U4635 (N_4635,N_1443,N_2381);
nor U4636 (N_4636,N_1400,N_1037);
nor U4637 (N_4637,N_2371,N_1130);
and U4638 (N_4638,N_689,N_38);
or U4639 (N_4639,N_997,N_1789);
xnor U4640 (N_4640,N_1161,N_1943);
and U4641 (N_4641,N_56,N_13);
nor U4642 (N_4642,N_1382,N_710);
or U4643 (N_4643,N_604,N_234);
and U4644 (N_4644,N_350,N_177);
or U4645 (N_4645,N_2235,N_1791);
nor U4646 (N_4646,N_1903,N_2135);
xor U4647 (N_4647,N_1640,N_2426);
or U4648 (N_4648,N_1689,N_1659);
nor U4649 (N_4649,N_1806,N_477);
or U4650 (N_4650,N_1794,N_677);
xnor U4651 (N_4651,N_1409,N_2495);
xor U4652 (N_4652,N_824,N_694);
nor U4653 (N_4653,N_258,N_2132);
and U4654 (N_4654,N_1500,N_845);
or U4655 (N_4655,N_165,N_1646);
nand U4656 (N_4656,N_1540,N_2135);
and U4657 (N_4657,N_101,N_2282);
xor U4658 (N_4658,N_965,N_961);
and U4659 (N_4659,N_952,N_1972);
nand U4660 (N_4660,N_1474,N_1701);
nor U4661 (N_4661,N_1315,N_269);
or U4662 (N_4662,N_1470,N_737);
nor U4663 (N_4663,N_1912,N_1374);
and U4664 (N_4664,N_528,N_2426);
nor U4665 (N_4665,N_1056,N_2284);
nor U4666 (N_4666,N_2049,N_352);
nand U4667 (N_4667,N_125,N_1925);
and U4668 (N_4668,N_557,N_1261);
xnor U4669 (N_4669,N_1226,N_1751);
and U4670 (N_4670,N_2050,N_1831);
or U4671 (N_4671,N_1867,N_611);
or U4672 (N_4672,N_246,N_724);
and U4673 (N_4673,N_1606,N_908);
and U4674 (N_4674,N_1684,N_1290);
or U4675 (N_4675,N_414,N_155);
or U4676 (N_4676,N_2408,N_1406);
xor U4677 (N_4677,N_1360,N_2340);
xnor U4678 (N_4678,N_1122,N_2383);
or U4679 (N_4679,N_2309,N_1163);
xnor U4680 (N_4680,N_1096,N_886);
or U4681 (N_4681,N_1884,N_676);
and U4682 (N_4682,N_537,N_1972);
xnor U4683 (N_4683,N_1300,N_846);
and U4684 (N_4684,N_593,N_1286);
xor U4685 (N_4685,N_2225,N_1675);
xor U4686 (N_4686,N_1902,N_12);
or U4687 (N_4687,N_1948,N_2058);
nand U4688 (N_4688,N_395,N_2229);
xnor U4689 (N_4689,N_2084,N_1072);
xor U4690 (N_4690,N_59,N_510);
nor U4691 (N_4691,N_524,N_1644);
xor U4692 (N_4692,N_1212,N_712);
and U4693 (N_4693,N_711,N_193);
xnor U4694 (N_4694,N_9,N_2092);
nor U4695 (N_4695,N_978,N_1861);
nor U4696 (N_4696,N_2291,N_1090);
nor U4697 (N_4697,N_1413,N_999);
or U4698 (N_4698,N_690,N_1925);
nand U4699 (N_4699,N_646,N_319);
nand U4700 (N_4700,N_429,N_972);
xnor U4701 (N_4701,N_763,N_2432);
xnor U4702 (N_4702,N_1132,N_631);
nand U4703 (N_4703,N_320,N_1478);
nand U4704 (N_4704,N_564,N_527);
or U4705 (N_4705,N_2021,N_1398);
xnor U4706 (N_4706,N_1932,N_1161);
or U4707 (N_4707,N_2363,N_1286);
or U4708 (N_4708,N_2137,N_674);
xor U4709 (N_4709,N_1385,N_1632);
or U4710 (N_4710,N_1381,N_174);
xnor U4711 (N_4711,N_1275,N_2277);
nor U4712 (N_4712,N_1186,N_730);
or U4713 (N_4713,N_1015,N_1091);
nor U4714 (N_4714,N_655,N_2339);
and U4715 (N_4715,N_605,N_1710);
nand U4716 (N_4716,N_1652,N_634);
xor U4717 (N_4717,N_401,N_1633);
nand U4718 (N_4718,N_849,N_714);
and U4719 (N_4719,N_653,N_468);
and U4720 (N_4720,N_741,N_1009);
xnor U4721 (N_4721,N_2361,N_835);
nor U4722 (N_4722,N_1937,N_1563);
nand U4723 (N_4723,N_1420,N_69);
and U4724 (N_4724,N_1839,N_1190);
nor U4725 (N_4725,N_2099,N_1257);
or U4726 (N_4726,N_1924,N_154);
nand U4727 (N_4727,N_756,N_1589);
xor U4728 (N_4728,N_625,N_2065);
nor U4729 (N_4729,N_2197,N_126);
xnor U4730 (N_4730,N_1289,N_1502);
xor U4731 (N_4731,N_1213,N_1447);
nor U4732 (N_4732,N_1891,N_738);
nand U4733 (N_4733,N_748,N_1080);
nor U4734 (N_4734,N_350,N_1099);
nor U4735 (N_4735,N_259,N_437);
xor U4736 (N_4736,N_1486,N_87);
xor U4737 (N_4737,N_416,N_483);
or U4738 (N_4738,N_1292,N_2429);
nor U4739 (N_4739,N_1474,N_2312);
and U4740 (N_4740,N_296,N_1368);
nor U4741 (N_4741,N_1697,N_372);
or U4742 (N_4742,N_331,N_535);
and U4743 (N_4743,N_1641,N_2386);
nor U4744 (N_4744,N_555,N_1578);
and U4745 (N_4745,N_551,N_9);
xor U4746 (N_4746,N_1249,N_314);
nor U4747 (N_4747,N_1119,N_190);
nor U4748 (N_4748,N_1843,N_202);
nor U4749 (N_4749,N_2416,N_459);
or U4750 (N_4750,N_510,N_2236);
or U4751 (N_4751,N_699,N_886);
and U4752 (N_4752,N_1954,N_1427);
and U4753 (N_4753,N_411,N_2010);
nor U4754 (N_4754,N_1805,N_2058);
xor U4755 (N_4755,N_657,N_1799);
or U4756 (N_4756,N_1670,N_1488);
and U4757 (N_4757,N_897,N_1484);
and U4758 (N_4758,N_1680,N_2120);
nor U4759 (N_4759,N_433,N_931);
nor U4760 (N_4760,N_1716,N_1003);
nand U4761 (N_4761,N_1386,N_105);
and U4762 (N_4762,N_692,N_1563);
nor U4763 (N_4763,N_1008,N_1060);
or U4764 (N_4764,N_263,N_1512);
nand U4765 (N_4765,N_2170,N_697);
nor U4766 (N_4766,N_910,N_160);
or U4767 (N_4767,N_2333,N_1332);
nor U4768 (N_4768,N_632,N_511);
or U4769 (N_4769,N_1582,N_306);
or U4770 (N_4770,N_83,N_2025);
nor U4771 (N_4771,N_556,N_1401);
or U4772 (N_4772,N_2252,N_1669);
xnor U4773 (N_4773,N_1822,N_1647);
nor U4774 (N_4774,N_381,N_80);
nor U4775 (N_4775,N_1076,N_416);
or U4776 (N_4776,N_1828,N_2210);
xor U4777 (N_4777,N_67,N_1938);
and U4778 (N_4778,N_2399,N_2196);
and U4779 (N_4779,N_101,N_538);
nor U4780 (N_4780,N_1017,N_1464);
nor U4781 (N_4781,N_1553,N_772);
nor U4782 (N_4782,N_2375,N_1356);
nor U4783 (N_4783,N_1135,N_218);
and U4784 (N_4784,N_645,N_873);
nor U4785 (N_4785,N_2447,N_174);
nand U4786 (N_4786,N_504,N_1344);
nand U4787 (N_4787,N_1871,N_662);
nor U4788 (N_4788,N_2155,N_948);
and U4789 (N_4789,N_1040,N_2003);
xnor U4790 (N_4790,N_308,N_1905);
and U4791 (N_4791,N_175,N_1802);
and U4792 (N_4792,N_1353,N_246);
nor U4793 (N_4793,N_103,N_1179);
nand U4794 (N_4794,N_1689,N_1046);
nand U4795 (N_4795,N_1823,N_2303);
and U4796 (N_4796,N_1799,N_753);
or U4797 (N_4797,N_1883,N_1774);
and U4798 (N_4798,N_665,N_1237);
nor U4799 (N_4799,N_1419,N_45);
nand U4800 (N_4800,N_2121,N_223);
nor U4801 (N_4801,N_473,N_2125);
xnor U4802 (N_4802,N_0,N_1013);
and U4803 (N_4803,N_1955,N_2207);
nor U4804 (N_4804,N_1727,N_1257);
and U4805 (N_4805,N_238,N_2456);
nand U4806 (N_4806,N_1176,N_2012);
nor U4807 (N_4807,N_977,N_1143);
nor U4808 (N_4808,N_627,N_912);
xor U4809 (N_4809,N_1088,N_2234);
xor U4810 (N_4810,N_2032,N_1522);
and U4811 (N_4811,N_865,N_702);
nor U4812 (N_4812,N_269,N_928);
nand U4813 (N_4813,N_1043,N_1212);
xor U4814 (N_4814,N_2441,N_897);
and U4815 (N_4815,N_12,N_1404);
nor U4816 (N_4816,N_2356,N_63);
xor U4817 (N_4817,N_890,N_596);
or U4818 (N_4818,N_601,N_1443);
xor U4819 (N_4819,N_272,N_2329);
xnor U4820 (N_4820,N_1811,N_1584);
nor U4821 (N_4821,N_2284,N_1740);
xnor U4822 (N_4822,N_584,N_806);
xnor U4823 (N_4823,N_125,N_1388);
and U4824 (N_4824,N_974,N_2381);
xor U4825 (N_4825,N_490,N_538);
nor U4826 (N_4826,N_1676,N_454);
or U4827 (N_4827,N_774,N_2000);
nand U4828 (N_4828,N_1627,N_588);
nand U4829 (N_4829,N_1474,N_1980);
xor U4830 (N_4830,N_2492,N_403);
nand U4831 (N_4831,N_821,N_186);
xor U4832 (N_4832,N_805,N_2001);
nand U4833 (N_4833,N_430,N_362);
and U4834 (N_4834,N_737,N_1990);
and U4835 (N_4835,N_2148,N_1724);
nand U4836 (N_4836,N_2064,N_1749);
xnor U4837 (N_4837,N_683,N_962);
xor U4838 (N_4838,N_1276,N_913);
nand U4839 (N_4839,N_997,N_1238);
xor U4840 (N_4840,N_538,N_1303);
nand U4841 (N_4841,N_2210,N_1463);
or U4842 (N_4842,N_1833,N_1452);
nor U4843 (N_4843,N_2177,N_562);
or U4844 (N_4844,N_1646,N_955);
nor U4845 (N_4845,N_777,N_1149);
and U4846 (N_4846,N_1816,N_2409);
nor U4847 (N_4847,N_664,N_1505);
and U4848 (N_4848,N_1788,N_1636);
nand U4849 (N_4849,N_1273,N_1730);
nor U4850 (N_4850,N_2268,N_2064);
nand U4851 (N_4851,N_120,N_19);
nor U4852 (N_4852,N_1632,N_1637);
xor U4853 (N_4853,N_1378,N_64);
nor U4854 (N_4854,N_2078,N_1923);
xor U4855 (N_4855,N_144,N_2186);
nor U4856 (N_4856,N_1758,N_1961);
nand U4857 (N_4857,N_2257,N_126);
nor U4858 (N_4858,N_2108,N_2083);
and U4859 (N_4859,N_623,N_1496);
or U4860 (N_4860,N_1978,N_2356);
nor U4861 (N_4861,N_1680,N_760);
and U4862 (N_4862,N_2247,N_409);
or U4863 (N_4863,N_316,N_260);
nor U4864 (N_4864,N_415,N_1589);
or U4865 (N_4865,N_1615,N_328);
and U4866 (N_4866,N_765,N_94);
xor U4867 (N_4867,N_2380,N_1075);
nand U4868 (N_4868,N_1690,N_904);
nor U4869 (N_4869,N_970,N_2286);
nand U4870 (N_4870,N_530,N_1481);
or U4871 (N_4871,N_1849,N_1074);
or U4872 (N_4872,N_1012,N_1415);
nor U4873 (N_4873,N_2337,N_2271);
xor U4874 (N_4874,N_1915,N_2483);
nand U4875 (N_4875,N_1449,N_2039);
nand U4876 (N_4876,N_1113,N_1705);
and U4877 (N_4877,N_918,N_1421);
or U4878 (N_4878,N_1169,N_2408);
and U4879 (N_4879,N_1836,N_499);
nor U4880 (N_4880,N_1038,N_223);
or U4881 (N_4881,N_2304,N_231);
nand U4882 (N_4882,N_2363,N_1730);
nand U4883 (N_4883,N_139,N_2288);
or U4884 (N_4884,N_1842,N_1335);
nor U4885 (N_4885,N_2093,N_126);
xor U4886 (N_4886,N_595,N_0);
nor U4887 (N_4887,N_2385,N_1457);
and U4888 (N_4888,N_2252,N_1042);
nand U4889 (N_4889,N_1622,N_2032);
nor U4890 (N_4890,N_1934,N_683);
nand U4891 (N_4891,N_604,N_246);
or U4892 (N_4892,N_1868,N_1098);
xnor U4893 (N_4893,N_299,N_1);
nand U4894 (N_4894,N_596,N_2432);
nand U4895 (N_4895,N_1804,N_1685);
and U4896 (N_4896,N_305,N_1877);
nor U4897 (N_4897,N_775,N_558);
or U4898 (N_4898,N_294,N_1542);
nand U4899 (N_4899,N_1547,N_1643);
and U4900 (N_4900,N_646,N_1586);
or U4901 (N_4901,N_217,N_2265);
and U4902 (N_4902,N_1065,N_599);
or U4903 (N_4903,N_106,N_2320);
or U4904 (N_4904,N_2362,N_777);
and U4905 (N_4905,N_1348,N_1575);
nor U4906 (N_4906,N_2304,N_2134);
xor U4907 (N_4907,N_2218,N_1503);
nor U4908 (N_4908,N_2439,N_236);
nor U4909 (N_4909,N_2244,N_1890);
xor U4910 (N_4910,N_1939,N_2089);
and U4911 (N_4911,N_459,N_612);
xor U4912 (N_4912,N_530,N_514);
xnor U4913 (N_4913,N_2102,N_1501);
nor U4914 (N_4914,N_316,N_1723);
and U4915 (N_4915,N_2130,N_1971);
xnor U4916 (N_4916,N_1423,N_969);
and U4917 (N_4917,N_944,N_1687);
and U4918 (N_4918,N_1105,N_939);
and U4919 (N_4919,N_1842,N_729);
nand U4920 (N_4920,N_1542,N_1071);
and U4921 (N_4921,N_1153,N_59);
nor U4922 (N_4922,N_232,N_916);
xor U4923 (N_4923,N_1216,N_223);
nand U4924 (N_4924,N_999,N_2247);
and U4925 (N_4925,N_1430,N_1354);
nand U4926 (N_4926,N_1673,N_2423);
or U4927 (N_4927,N_164,N_2259);
or U4928 (N_4928,N_1920,N_366);
nor U4929 (N_4929,N_28,N_2127);
nor U4930 (N_4930,N_2390,N_969);
and U4931 (N_4931,N_2300,N_1379);
nand U4932 (N_4932,N_1323,N_1655);
nand U4933 (N_4933,N_1927,N_1806);
nor U4934 (N_4934,N_2315,N_493);
or U4935 (N_4935,N_1886,N_968);
or U4936 (N_4936,N_1352,N_128);
and U4937 (N_4937,N_861,N_1545);
or U4938 (N_4938,N_1304,N_647);
nand U4939 (N_4939,N_2343,N_812);
nand U4940 (N_4940,N_2447,N_1166);
nor U4941 (N_4941,N_1276,N_514);
xor U4942 (N_4942,N_739,N_806);
nand U4943 (N_4943,N_480,N_2480);
and U4944 (N_4944,N_2191,N_1719);
nand U4945 (N_4945,N_9,N_1550);
nor U4946 (N_4946,N_692,N_1047);
nand U4947 (N_4947,N_1519,N_1732);
or U4948 (N_4948,N_2020,N_795);
or U4949 (N_4949,N_2092,N_2166);
nor U4950 (N_4950,N_1381,N_2385);
and U4951 (N_4951,N_1200,N_821);
or U4952 (N_4952,N_363,N_1181);
nand U4953 (N_4953,N_1798,N_1114);
nand U4954 (N_4954,N_2202,N_1337);
or U4955 (N_4955,N_2265,N_1432);
and U4956 (N_4956,N_1495,N_1468);
nor U4957 (N_4957,N_1749,N_2423);
and U4958 (N_4958,N_120,N_1698);
and U4959 (N_4959,N_34,N_471);
or U4960 (N_4960,N_1506,N_1472);
nand U4961 (N_4961,N_2095,N_1061);
xor U4962 (N_4962,N_1681,N_1584);
or U4963 (N_4963,N_2283,N_1592);
and U4964 (N_4964,N_304,N_1081);
nand U4965 (N_4965,N_1030,N_1421);
or U4966 (N_4966,N_252,N_2465);
and U4967 (N_4967,N_961,N_1907);
xor U4968 (N_4968,N_1556,N_1820);
nand U4969 (N_4969,N_947,N_1798);
and U4970 (N_4970,N_2168,N_1786);
or U4971 (N_4971,N_2320,N_136);
or U4972 (N_4972,N_379,N_2267);
nand U4973 (N_4973,N_1685,N_1447);
nor U4974 (N_4974,N_813,N_321);
xnor U4975 (N_4975,N_166,N_560);
nand U4976 (N_4976,N_1903,N_511);
and U4977 (N_4977,N_2363,N_760);
nand U4978 (N_4978,N_2032,N_1651);
and U4979 (N_4979,N_140,N_1804);
nand U4980 (N_4980,N_636,N_116);
nor U4981 (N_4981,N_1788,N_1933);
nand U4982 (N_4982,N_947,N_248);
and U4983 (N_4983,N_1638,N_1305);
nand U4984 (N_4984,N_2328,N_384);
nor U4985 (N_4985,N_854,N_835);
xnor U4986 (N_4986,N_405,N_44);
xor U4987 (N_4987,N_1255,N_163);
or U4988 (N_4988,N_43,N_1001);
nand U4989 (N_4989,N_2337,N_620);
or U4990 (N_4990,N_353,N_1076);
nor U4991 (N_4991,N_61,N_1925);
nor U4992 (N_4992,N_87,N_190);
nand U4993 (N_4993,N_823,N_669);
xor U4994 (N_4994,N_386,N_590);
nor U4995 (N_4995,N_549,N_1273);
and U4996 (N_4996,N_1149,N_1587);
xor U4997 (N_4997,N_1769,N_607);
nand U4998 (N_4998,N_578,N_697);
and U4999 (N_4999,N_1846,N_2190);
and U5000 (N_5000,N_2828,N_4556);
xor U5001 (N_5001,N_3563,N_2525);
and U5002 (N_5002,N_3576,N_4656);
nor U5003 (N_5003,N_3490,N_4717);
xor U5004 (N_5004,N_3163,N_3437);
nor U5005 (N_5005,N_4232,N_4950);
nor U5006 (N_5006,N_3479,N_4244);
or U5007 (N_5007,N_3422,N_4849);
nand U5008 (N_5008,N_3887,N_4105);
or U5009 (N_5009,N_3673,N_2745);
xnor U5010 (N_5010,N_4607,N_4666);
and U5011 (N_5011,N_4502,N_3311);
nand U5012 (N_5012,N_4984,N_4142);
and U5013 (N_5013,N_3614,N_2797);
nor U5014 (N_5014,N_3387,N_4077);
nor U5015 (N_5015,N_3016,N_3849);
xnor U5016 (N_5016,N_4807,N_2990);
xor U5017 (N_5017,N_4458,N_3432);
and U5018 (N_5018,N_4008,N_4185);
or U5019 (N_5019,N_2758,N_3644);
and U5020 (N_5020,N_3678,N_4843);
and U5021 (N_5021,N_3996,N_4390);
nand U5022 (N_5022,N_4327,N_3018);
xor U5023 (N_5023,N_3103,N_4044);
nor U5024 (N_5024,N_4217,N_3752);
nor U5025 (N_5025,N_2904,N_3938);
nand U5026 (N_5026,N_3928,N_4269);
or U5027 (N_5027,N_2910,N_3127);
xnor U5028 (N_5028,N_4226,N_3304);
and U5029 (N_5029,N_4288,N_3917);
or U5030 (N_5030,N_4793,N_4762);
xnor U5031 (N_5031,N_2644,N_3945);
nor U5032 (N_5032,N_4048,N_4419);
nand U5033 (N_5033,N_2515,N_4052);
xnor U5034 (N_5034,N_2920,N_3805);
nand U5035 (N_5035,N_3181,N_3909);
xnor U5036 (N_5036,N_2539,N_2609);
xnor U5037 (N_5037,N_4910,N_4125);
nand U5038 (N_5038,N_2753,N_3014);
nor U5039 (N_5039,N_3662,N_3052);
or U5040 (N_5040,N_3472,N_3816);
or U5041 (N_5041,N_3112,N_3683);
nor U5042 (N_5042,N_3235,N_4735);
nand U5043 (N_5043,N_3225,N_3803);
nand U5044 (N_5044,N_2754,N_2816);
nor U5045 (N_5045,N_3345,N_4034);
xor U5046 (N_5046,N_3626,N_2839);
and U5047 (N_5047,N_3846,N_3725);
nand U5048 (N_5048,N_4119,N_2617);
or U5049 (N_5049,N_4069,N_4084);
nand U5050 (N_5050,N_3790,N_4025);
xor U5051 (N_5051,N_3090,N_2538);
or U5052 (N_5052,N_4505,N_4851);
and U5053 (N_5053,N_3141,N_4115);
nor U5054 (N_5054,N_4176,N_4167);
nand U5055 (N_5055,N_2632,N_3933);
and U5056 (N_5056,N_3366,N_3639);
nand U5057 (N_5057,N_2918,N_3902);
nand U5058 (N_5058,N_2720,N_4597);
and U5059 (N_5059,N_2832,N_3476);
nor U5060 (N_5060,N_4676,N_3426);
or U5061 (N_5061,N_2581,N_2897);
nor U5062 (N_5062,N_2991,N_3972);
and U5063 (N_5063,N_2624,N_3728);
nand U5064 (N_5064,N_4972,N_3810);
nor U5065 (N_5065,N_2824,N_2583);
nor U5066 (N_5066,N_4393,N_3467);
nor U5067 (N_5067,N_3723,N_2967);
and U5068 (N_5068,N_3044,N_2580);
xnor U5069 (N_5069,N_4781,N_4242);
xnor U5070 (N_5070,N_2642,N_4614);
xor U5071 (N_5071,N_4045,N_2606);
xnor U5072 (N_5072,N_2946,N_4492);
xor U5073 (N_5073,N_4079,N_3350);
or U5074 (N_5074,N_2605,N_2659);
nand U5075 (N_5075,N_3677,N_4090);
nand U5076 (N_5076,N_2603,N_4894);
and U5077 (N_5077,N_3844,N_4814);
xor U5078 (N_5078,N_4872,N_4833);
or U5079 (N_5079,N_3986,N_2662);
and U5080 (N_5080,N_3712,N_2995);
xnor U5081 (N_5081,N_3487,N_3824);
nand U5082 (N_5082,N_2727,N_2512);
nor U5083 (N_5083,N_2883,N_3295);
xor U5084 (N_5084,N_2845,N_3078);
and U5085 (N_5085,N_4483,N_3475);
or U5086 (N_5086,N_4938,N_4171);
nand U5087 (N_5087,N_3021,N_4999);
and U5088 (N_5088,N_3518,N_4734);
xnor U5089 (N_5089,N_3305,N_3533);
xor U5090 (N_5090,N_3047,N_4355);
or U5091 (N_5091,N_4058,N_3772);
nand U5092 (N_5092,N_3358,N_3084);
and U5093 (N_5093,N_3959,N_2980);
nor U5094 (N_5094,N_3690,N_3073);
xnor U5095 (N_5095,N_3002,N_2924);
xor U5096 (N_5096,N_2942,N_3099);
nand U5097 (N_5097,N_3540,N_3253);
nand U5098 (N_5098,N_3965,N_3268);
xor U5099 (N_5099,N_3332,N_4690);
and U5100 (N_5100,N_3561,N_3383);
nor U5101 (N_5101,N_3443,N_2909);
and U5102 (N_5102,N_3210,N_2841);
and U5103 (N_5103,N_3411,N_4400);
and U5104 (N_5104,N_3203,N_4943);
or U5105 (N_5105,N_3319,N_3504);
xor U5106 (N_5106,N_3123,N_4435);
nand U5107 (N_5107,N_2589,N_4612);
or U5108 (N_5108,N_3670,N_4399);
xor U5109 (N_5109,N_4006,N_3547);
xor U5110 (N_5110,N_4011,N_4716);
nor U5111 (N_5111,N_2798,N_3624);
xor U5112 (N_5112,N_4673,N_2806);
and U5113 (N_5113,N_4813,N_4160);
or U5114 (N_5114,N_4871,N_2545);
and U5115 (N_5115,N_3605,N_3987);
nand U5116 (N_5116,N_3742,N_2549);
or U5117 (N_5117,N_4291,N_4624);
or U5118 (N_5118,N_3615,N_2755);
and U5119 (N_5119,N_3468,N_4397);
nand U5120 (N_5120,N_2886,N_4737);
xnor U5121 (N_5121,N_2562,N_4574);
nand U5122 (N_5122,N_4481,N_3832);
or U5123 (N_5123,N_3229,N_4819);
xnor U5124 (N_5124,N_4305,N_3284);
xor U5125 (N_5125,N_3734,N_3714);
xnor U5126 (N_5126,N_2976,N_3762);
nand U5127 (N_5127,N_4699,N_3232);
nor U5128 (N_5128,N_4511,N_2922);
or U5129 (N_5129,N_4016,N_2945);
and U5130 (N_5130,N_2533,N_3367);
nor U5131 (N_5131,N_2936,N_3635);
nand U5132 (N_5132,N_3271,N_3687);
nand U5133 (N_5133,N_3226,N_4775);
and U5134 (N_5134,N_3156,N_4776);
nor U5135 (N_5135,N_4739,N_4420);
and U5136 (N_5136,N_4187,N_4777);
nand U5137 (N_5137,N_4946,N_4277);
or U5138 (N_5138,N_4279,N_3630);
nor U5139 (N_5139,N_3224,N_2697);
nor U5140 (N_5140,N_3169,N_4829);
nor U5141 (N_5141,N_4610,N_2628);
xor U5142 (N_5142,N_4310,N_2938);
nand U5143 (N_5143,N_3142,N_2656);
nand U5144 (N_5144,N_2981,N_2953);
and U5145 (N_5145,N_2524,N_4256);
nor U5146 (N_5146,N_2661,N_3019);
xnor U5147 (N_5147,N_4117,N_4152);
nor U5148 (N_5148,N_3006,N_3571);
or U5149 (N_5149,N_4884,N_4248);
xor U5150 (N_5150,N_2688,N_2738);
and U5151 (N_5151,N_4082,N_3372);
and U5152 (N_5152,N_2925,N_3557);
nand U5153 (N_5153,N_4559,N_4101);
and U5154 (N_5154,N_3030,N_3980);
or U5155 (N_5155,N_4875,N_4960);
or U5156 (N_5156,N_2705,N_2588);
and U5157 (N_5157,N_4982,N_3998);
xor U5158 (N_5158,N_3059,N_3981);
nor U5159 (N_5159,N_3149,N_2501);
xor U5160 (N_5160,N_4796,N_4845);
or U5161 (N_5161,N_2627,N_4463);
and U5162 (N_5162,N_4671,N_4694);
or U5163 (N_5163,N_4241,N_3858);
or U5164 (N_5164,N_4402,N_4832);
nand U5165 (N_5165,N_4335,N_3795);
and U5166 (N_5166,N_4484,N_3025);
xnor U5167 (N_5167,N_4792,N_3252);
and U5168 (N_5168,N_3489,N_3275);
nand U5169 (N_5169,N_4906,N_2794);
and U5170 (N_5170,N_3125,N_2633);
nand U5171 (N_5171,N_4204,N_2791);
nand U5172 (N_5172,N_4580,N_2903);
nand U5173 (N_5173,N_4499,N_3401);
or U5174 (N_5174,N_3863,N_3551);
and U5175 (N_5175,N_4951,N_2756);
nand U5176 (N_5176,N_3092,N_3347);
and U5177 (N_5177,N_4401,N_3553);
or U5178 (N_5178,N_3309,N_3348);
nand U5179 (N_5179,N_4467,N_3754);
nor U5180 (N_5180,N_3148,N_3173);
and U5181 (N_5181,N_3427,N_4782);
nor U5182 (N_5182,N_3206,N_2714);
nand U5183 (N_5183,N_3549,N_3128);
nor U5184 (N_5184,N_4616,N_3865);
or U5185 (N_5185,N_2969,N_3056);
and U5186 (N_5186,N_4754,N_4504);
nand U5187 (N_5187,N_3242,N_2666);
nand U5188 (N_5188,N_3536,N_3516);
or U5189 (N_5189,N_4599,N_3133);
and U5190 (N_5190,N_3447,N_3096);
or U5191 (N_5191,N_3595,N_2956);
xnor U5192 (N_5192,N_4664,N_2973);
nor U5193 (N_5193,N_3172,N_4245);
nand U5194 (N_5194,N_4398,N_3336);
or U5195 (N_5195,N_2629,N_4137);
nor U5196 (N_5196,N_2736,N_3953);
and U5197 (N_5197,N_4831,N_3370);
xnor U5198 (N_5198,N_4411,N_3501);
xor U5199 (N_5199,N_3814,N_3743);
nor U5200 (N_5200,N_3669,N_3509);
or U5201 (N_5201,N_4370,N_4095);
xor U5202 (N_5202,N_4562,N_3807);
and U5203 (N_5203,N_3162,N_2689);
or U5204 (N_5204,N_2805,N_4620);
xnor U5205 (N_5205,N_2560,N_2568);
or U5206 (N_5206,N_4609,N_4967);
nor U5207 (N_5207,N_2848,N_3100);
or U5208 (N_5208,N_3377,N_4102);
or U5209 (N_5209,N_2873,N_3759);
nand U5210 (N_5210,N_2680,N_2743);
nor U5211 (N_5211,N_3821,N_3695);
nor U5212 (N_5212,N_4628,N_4622);
nor U5213 (N_5213,N_3218,N_4383);
xnor U5214 (N_5214,N_3730,N_3094);
nor U5215 (N_5215,N_4183,N_3574);
or U5216 (N_5216,N_3622,N_2999);
or U5217 (N_5217,N_3581,N_3646);
or U5218 (N_5218,N_3261,N_3328);
nand U5219 (N_5219,N_2615,N_4635);
xor U5220 (N_5220,N_4979,N_2917);
nand U5221 (N_5221,N_3979,N_2602);
and U5222 (N_5222,N_3700,N_4001);
xnor U5223 (N_5223,N_3789,N_2664);
nor U5224 (N_5224,N_2812,N_4856);
nor U5225 (N_5225,N_4711,N_3943);
and U5226 (N_5226,N_4826,N_2665);
or U5227 (N_5227,N_4027,N_4750);
nor U5228 (N_5228,N_3322,N_3102);
nor U5229 (N_5229,N_2542,N_3698);
or U5230 (N_5230,N_2534,N_3825);
and U5231 (N_5231,N_4104,N_3600);
nand U5232 (N_5232,N_3619,N_3316);
nor U5233 (N_5233,N_2556,N_4643);
xnor U5234 (N_5234,N_4976,N_4852);
or U5235 (N_5235,N_3121,N_4306);
and U5236 (N_5236,N_4605,N_2856);
xor U5237 (N_5237,N_2929,N_3194);
nand U5238 (N_5238,N_4168,N_3641);
or U5239 (N_5239,N_4429,N_3167);
nand U5240 (N_5240,N_4904,N_3711);
nand U5241 (N_5241,N_3636,N_3596);
nand U5242 (N_5242,N_4756,N_4136);
nor U5243 (N_5243,N_4674,N_3282);
nor U5244 (N_5244,N_4692,N_3098);
nor U5245 (N_5245,N_4715,N_3135);
and U5246 (N_5246,N_3732,N_4421);
nor U5247 (N_5247,N_3541,N_3634);
nor U5248 (N_5248,N_4273,N_4560);
nor U5249 (N_5249,N_3245,N_3718);
nand U5250 (N_5250,N_4952,N_4258);
nor U5251 (N_5251,N_3374,N_3891);
nor U5252 (N_5252,N_4338,N_3404);
nand U5253 (N_5253,N_3031,N_4129);
nor U5254 (N_5254,N_2822,N_3150);
nand U5255 (N_5255,N_4047,N_4631);
nor U5256 (N_5256,N_4945,N_4472);
xor U5257 (N_5257,N_2707,N_4858);
and U5258 (N_5258,N_4249,N_2698);
nand U5259 (N_5259,N_4298,N_3330);
nand U5260 (N_5260,N_4391,N_4839);
and U5261 (N_5261,N_2837,N_3942);
nor U5262 (N_5262,N_2671,N_3667);
xnor U5263 (N_5263,N_4287,N_2862);
or U5264 (N_5264,N_4396,N_4278);
xnor U5265 (N_5265,N_3353,N_4169);
xor U5266 (N_5266,N_4377,N_2552);
xnor U5267 (N_5267,N_4521,N_2898);
nor U5268 (N_5268,N_3498,N_4966);
nand U5269 (N_5269,N_3813,N_4961);
xnor U5270 (N_5270,N_4446,N_3423);
nor U5271 (N_5271,N_4758,N_4932);
nor U5272 (N_5272,N_4650,N_4763);
nand U5273 (N_5273,N_4323,N_2882);
nor U5274 (N_5274,N_3567,N_4892);
nand U5275 (N_5275,N_3396,N_4330);
and U5276 (N_5276,N_2987,N_4085);
xnor U5277 (N_5277,N_3837,N_4968);
nand U5278 (N_5278,N_3523,N_4415);
or U5279 (N_5279,N_3244,N_4925);
xor U5280 (N_5280,N_2768,N_4148);
nand U5281 (N_5281,N_2594,N_3817);
nand U5282 (N_5282,N_4205,N_4773);
or U5283 (N_5283,N_2649,N_4641);
or U5284 (N_5284,N_3339,N_2825);
nand U5285 (N_5285,N_4382,N_3623);
and U5286 (N_5286,N_4326,N_2815);
and U5287 (N_5287,N_4811,N_4054);
or U5288 (N_5288,N_2817,N_4667);
or U5289 (N_5289,N_4325,N_2974);
nand U5290 (N_5290,N_3290,N_4088);
nand U5291 (N_5291,N_4726,N_2884);
and U5292 (N_5292,N_3886,N_3856);
or U5293 (N_5293,N_4962,N_3055);
xor U5294 (N_5294,N_3351,N_4710);
nand U5295 (N_5295,N_4658,N_3993);
nor U5296 (N_5296,N_3390,N_3045);
and U5297 (N_5297,N_3659,N_3845);
or U5298 (N_5298,N_3628,N_4886);
nor U5299 (N_5299,N_3081,N_4182);
and U5300 (N_5300,N_4023,N_3964);
nor U5301 (N_5301,N_2803,N_4384);
xor U5302 (N_5302,N_4022,N_2608);
and U5303 (N_5303,N_2701,N_4113);
xnor U5304 (N_5304,N_4779,N_3054);
nor U5305 (N_5305,N_3478,N_3034);
and U5306 (N_5306,N_4501,N_2595);
nand U5307 (N_5307,N_4935,N_3694);
nand U5308 (N_5308,N_3924,N_4426);
or U5309 (N_5309,N_4568,N_3480);
nand U5310 (N_5310,N_2963,N_3531);
or U5311 (N_5311,N_3483,N_3452);
and U5312 (N_5312,N_4495,N_3583);
and U5313 (N_5313,N_4579,N_3913);
nand U5314 (N_5314,N_2826,N_4549);
xnor U5315 (N_5315,N_2639,N_4003);
and U5316 (N_5316,N_3503,N_4324);
xor U5317 (N_5317,N_4451,N_3606);
nand U5318 (N_5318,N_3454,N_3360);
xnor U5319 (N_5319,N_4526,N_4911);
nand U5320 (N_5320,N_3895,N_3604);
nor U5321 (N_5321,N_3970,N_3896);
nand U5322 (N_5322,N_3978,N_3114);
or U5323 (N_5323,N_3313,N_2785);
xor U5324 (N_5324,N_4418,N_4216);
or U5325 (N_5325,N_4440,N_4417);
and U5326 (N_5326,N_4977,N_4311);
nor U5327 (N_5327,N_4144,N_3875);
nor U5328 (N_5328,N_2977,N_3855);
and U5329 (N_5329,N_4770,N_3451);
or U5330 (N_5330,N_3588,N_3804);
nand U5331 (N_5331,N_3269,N_4661);
xnor U5332 (N_5332,N_4862,N_3420);
xor U5333 (N_5333,N_4714,N_3053);
and U5334 (N_5334,N_3082,N_4114);
or U5335 (N_5335,N_3836,N_3838);
xnor U5336 (N_5336,N_3591,N_2939);
nand U5337 (N_5337,N_4410,N_4838);
nand U5338 (N_5338,N_4527,N_2696);
xnor U5339 (N_5339,N_3524,N_3653);
nor U5340 (N_5340,N_4333,N_4140);
xnor U5341 (N_5341,N_3136,N_4198);
nor U5342 (N_5342,N_2699,N_4744);
nor U5343 (N_5343,N_2792,N_4476);
and U5344 (N_5344,N_4747,N_3592);
or U5345 (N_5345,N_3668,N_2637);
nor U5346 (N_5346,N_3930,N_3629);
nand U5347 (N_5347,N_4460,N_3236);
or U5348 (N_5348,N_4316,N_4606);
and U5349 (N_5349,N_3841,N_4141);
nand U5350 (N_5350,N_2682,N_2574);
nand U5351 (N_5351,N_4211,N_4753);
nand U5352 (N_5352,N_3897,N_4123);
and U5353 (N_5353,N_4888,N_4367);
and U5354 (N_5354,N_2687,N_2874);
or U5355 (N_5355,N_4820,N_4809);
or U5356 (N_5356,N_3187,N_4877);
xnor U5357 (N_5357,N_3397,N_2867);
nand U5358 (N_5358,N_2630,N_3257);
nand U5359 (N_5359,N_3948,N_3684);
and U5360 (N_5360,N_2730,N_4060);
xor U5361 (N_5361,N_3147,N_2959);
nand U5362 (N_5362,N_2932,N_3900);
or U5363 (N_5363,N_3392,N_3241);
xnor U5364 (N_5364,N_3657,N_4997);
nor U5365 (N_5365,N_4379,N_4728);
nor U5366 (N_5366,N_3130,N_3934);
nor U5367 (N_5367,N_2590,N_4577);
xor U5368 (N_5368,N_2610,N_4196);
nand U5369 (N_5369,N_2681,N_3376);
xnor U5370 (N_5370,N_4959,N_4145);
or U5371 (N_5371,N_4213,N_4500);
nor U5372 (N_5372,N_3363,N_4608);
and U5373 (N_5373,N_3748,N_4707);
and U5374 (N_5374,N_4172,N_4905);
or U5375 (N_5375,N_3607,N_4083);
nor U5376 (N_5376,N_4318,N_4339);
nor U5377 (N_5377,N_3027,N_2895);
xnor U5378 (N_5378,N_3111,N_4578);
and U5379 (N_5379,N_4810,N_3521);
and U5380 (N_5380,N_3767,N_3165);
xor U5381 (N_5381,N_2514,N_3051);
nor U5382 (N_5382,N_4109,N_3637);
or U5383 (N_5383,N_3949,N_4682);
xnor U5384 (N_5384,N_3876,N_3079);
nor U5385 (N_5385,N_2618,N_4917);
or U5386 (N_5386,N_2535,N_2934);
nor U5387 (N_5387,N_4456,N_4257);
and U5388 (N_5388,N_3024,N_3124);
xor U5389 (N_5389,N_2572,N_2927);
nor U5390 (N_5390,N_3326,N_3508);
or U5391 (N_5391,N_4519,N_3901);
and U5392 (N_5392,N_3435,N_4385);
xor U5393 (N_5393,N_4683,N_2935);
or U5394 (N_5394,N_2717,N_3652);
nor U5395 (N_5395,N_4395,N_3005);
or U5396 (N_5396,N_3113,N_4889);
nor U5397 (N_5397,N_2989,N_3361);
nor U5398 (N_5398,N_3270,N_4271);
nor U5399 (N_5399,N_4828,N_3962);
xnor U5400 (N_5400,N_4882,N_2750);
and U5401 (N_5401,N_2955,N_2773);
nor U5402 (N_5402,N_4538,N_4535);
xor U5403 (N_5403,N_2849,N_4515);
nand U5404 (N_5404,N_4679,N_2529);
and U5405 (N_5405,N_4723,N_2760);
and U5406 (N_5406,N_3442,N_2718);
and U5407 (N_5407,N_3032,N_4774);
nand U5408 (N_5408,N_4471,N_4425);
nor U5409 (N_5409,N_4736,N_2554);
xnor U5410 (N_5410,N_4948,N_4637);
nor U5411 (N_5411,N_4303,N_4342);
xnor U5412 (N_5412,N_4354,N_4569);
xor U5413 (N_5413,N_2952,N_4290);
xnor U5414 (N_5414,N_4441,N_2994);
nand U5415 (N_5415,N_3450,N_3864);
nand U5416 (N_5416,N_4931,N_4755);
xor U5417 (N_5417,N_3449,N_4010);
and U5418 (N_5418,N_4567,N_3794);
or U5419 (N_5419,N_4509,N_2546);
nor U5420 (N_5420,N_3608,N_3212);
and U5421 (N_5421,N_4017,N_3138);
and U5422 (N_5422,N_3932,N_4700);
nor U5423 (N_5423,N_3492,N_4051);
and U5424 (N_5424,N_4223,N_3899);
and U5425 (N_5425,N_3453,N_3413);
and U5426 (N_5426,N_2887,N_4665);
or U5427 (N_5427,N_2695,N_3013);
nor U5428 (N_5428,N_2557,N_3057);
nand U5429 (N_5429,N_2821,N_2737);
nand U5430 (N_5430,N_4955,N_4103);
nand U5431 (N_5431,N_3407,N_4812);
nand U5432 (N_5432,N_4473,N_3170);
and U5433 (N_5433,N_4301,N_3579);
or U5434 (N_5434,N_3424,N_4254);
nor U5435 (N_5435,N_4212,N_3947);
nand U5436 (N_5436,N_4036,N_4029);
or U5437 (N_5437,N_2614,N_3009);
xor U5438 (N_5438,N_2735,N_3317);
nand U5439 (N_5439,N_3799,N_3860);
nand U5440 (N_5440,N_3915,N_3935);
xor U5441 (N_5441,N_3048,N_4281);
nand U5442 (N_5442,N_4076,N_3240);
xnor U5443 (N_5443,N_4970,N_3093);
or U5444 (N_5444,N_4272,N_4804);
nand U5445 (N_5445,N_2643,N_4424);
and U5446 (N_5446,N_3904,N_3775);
or U5447 (N_5447,N_2842,N_3122);
nand U5448 (N_5448,N_3441,N_3246);
nor U5449 (N_5449,N_3815,N_3705);
and U5450 (N_5450,N_4049,N_3087);
xor U5451 (N_5451,N_3765,N_3802);
xor U5452 (N_5452,N_4663,N_3207);
and U5453 (N_5453,N_4146,N_3076);
nor U5454 (N_5454,N_2985,N_3385);
and U5455 (N_5455,N_3859,N_4985);
nand U5456 (N_5456,N_4436,N_4934);
nand U5457 (N_5457,N_4315,N_4590);
nand U5458 (N_5458,N_3343,N_4646);
or U5459 (N_5459,N_4416,N_3249);
nand U5460 (N_5460,N_4879,N_4973);
and U5461 (N_5461,N_4337,N_3538);
and U5462 (N_5462,N_4649,N_3749);
xnor U5463 (N_5463,N_3780,N_2641);
nor U5464 (N_5464,N_3457,N_3602);
or U5465 (N_5465,N_3822,N_3850);
or U5466 (N_5466,N_3688,N_3520);
xor U5467 (N_5467,N_2807,N_4822);
nand U5468 (N_5468,N_4604,N_4963);
or U5469 (N_5469,N_3310,N_4220);
and U5470 (N_5470,N_2547,N_3337);
xnor U5471 (N_5471,N_4947,N_2744);
nand U5472 (N_5472,N_2752,N_3618);
xnor U5473 (N_5473,N_4121,N_3617);
and U5474 (N_5474,N_3408,N_4857);
nand U5475 (N_5475,N_3983,N_3726);
and U5476 (N_5476,N_4514,N_3243);
nand U5477 (N_5477,N_3564,N_4588);
nand U5478 (N_5478,N_4469,N_2520);
nand U5479 (N_5479,N_4722,N_4642);
nand U5480 (N_5480,N_2612,N_3929);
and U5481 (N_5481,N_2777,N_3080);
and U5482 (N_5482,N_4687,N_4228);
or U5483 (N_5483,N_3023,N_4929);
xnor U5484 (N_5484,N_3386,N_3693);
nand U5485 (N_5485,N_4381,N_4994);
nor U5486 (N_5486,N_4799,N_3560);
nand U5487 (N_5487,N_4496,N_4219);
and U5488 (N_5488,N_3126,N_3656);
nor U5489 (N_5489,N_3709,N_2693);
and U5490 (N_5490,N_3968,N_2729);
and U5491 (N_5491,N_4532,N_2933);
nor U5492 (N_5492,N_2719,N_3513);
xor U5493 (N_5493,N_2764,N_3101);
xor U5494 (N_5494,N_4179,N_4644);
or U5495 (N_5495,N_3288,N_4053);
nor U5496 (N_5496,N_2638,N_4173);
nand U5497 (N_5497,N_3399,N_3511);
xnor U5498 (N_5498,N_3593,N_2947);
nand U5499 (N_5499,N_2598,N_3391);
nand U5500 (N_5500,N_4954,N_4127);
nand U5501 (N_5501,N_4971,N_3176);
nand U5502 (N_5502,N_4107,N_4551);
nor U5503 (N_5503,N_2650,N_4874);
nor U5504 (N_5504,N_3756,N_3747);
nand U5505 (N_5505,N_4615,N_3573);
and U5506 (N_5506,N_2746,N_4178);
nand U5507 (N_5507,N_3958,N_2563);
and U5508 (N_5508,N_3505,N_4778);
nand U5509 (N_5509,N_4433,N_3470);
xor U5510 (N_5510,N_4487,N_2732);
nand U5511 (N_5511,N_4294,N_4834);
or U5512 (N_5512,N_2866,N_4485);
nand U5513 (N_5513,N_3888,N_3661);
nand U5514 (N_5514,N_3868,N_4304);
nand U5515 (N_5515,N_4392,N_4203);
nand U5516 (N_5516,N_4540,N_4050);
or U5517 (N_5517,N_3415,N_3037);
or U5518 (N_5518,N_3209,N_4914);
nor U5519 (N_5519,N_3590,N_3258);
nand U5520 (N_5520,N_2799,N_4891);
or U5521 (N_5521,N_2778,N_3828);
nand U5522 (N_5522,N_4409,N_3445);
nor U5523 (N_5523,N_4863,N_3969);
and U5524 (N_5524,N_3004,N_4903);
or U5525 (N_5525,N_2850,N_4825);
xnor U5526 (N_5526,N_2912,N_4126);
nand U5527 (N_5527,N_4513,N_4721);
or U5528 (N_5528,N_4724,N_3455);
nand U5529 (N_5529,N_4771,N_3003);
xor U5530 (N_5530,N_2616,N_4890);
xnor U5531 (N_5531,N_4844,N_3961);
xor U5532 (N_5532,N_4177,N_3405);
nand U5533 (N_5533,N_3830,N_3854);
or U5534 (N_5534,N_4772,N_3281);
nor U5535 (N_5535,N_3826,N_3314);
xnor U5536 (N_5536,N_2790,N_3294);
xnor U5537 (N_5537,N_3355,N_2631);
nor U5538 (N_5538,N_4462,N_2694);
xnor U5539 (N_5539,N_4002,N_4037);
and U5540 (N_5540,N_3717,N_3552);
nand U5541 (N_5541,N_3587,N_3545);
nand U5542 (N_5542,N_4328,N_3211);
nand U5543 (N_5543,N_4366,N_3381);
nor U5544 (N_5544,N_4089,N_4336);
nor U5545 (N_5545,N_2676,N_4803);
nand U5546 (N_5546,N_3190,N_4477);
and U5547 (N_5547,N_4709,N_4474);
nor U5548 (N_5548,N_4633,N_3555);
and U5549 (N_5549,N_2855,N_3597);
and U5550 (N_5550,N_4595,N_3713);
and U5551 (N_5551,N_2857,N_4741);
nand U5552 (N_5552,N_3685,N_2905);
xor U5553 (N_5553,N_4746,N_3327);
xnor U5554 (N_5554,N_2648,N_4885);
nand U5555 (N_5555,N_3650,N_3085);
or U5556 (N_5556,N_2700,N_3689);
nor U5557 (N_5557,N_4209,N_4795);
or U5558 (N_5558,N_4539,N_4743);
nand U5559 (N_5559,N_3421,N_3880);
or U5560 (N_5560,N_3878,N_3342);
nand U5561 (N_5561,N_3352,N_4246);
xor U5562 (N_5562,N_3502,N_2836);
nor U5563 (N_5563,N_4091,N_3853);
and U5564 (N_5564,N_4170,N_2599);
xnor U5565 (N_5565,N_2558,N_3183);
nand U5566 (N_5566,N_2960,N_4252);
xnor U5567 (N_5567,N_3529,N_3192);
nor U5568 (N_5568,N_3633,N_4581);
nand U5569 (N_5569,N_4553,N_3692);
and U5570 (N_5570,N_4861,N_4919);
or U5571 (N_5571,N_3247,N_3308);
nor U5572 (N_5572,N_4701,N_2992);
and U5573 (N_5573,N_3129,N_4237);
nor U5574 (N_5574,N_4131,N_4640);
xor U5575 (N_5575,N_3827,N_2566);
xor U5576 (N_5576,N_4685,N_3640);
nor U5577 (N_5577,N_4043,N_3565);
xnor U5578 (N_5578,N_3776,N_4265);
nor U5579 (N_5579,N_4378,N_4587);
and U5580 (N_5580,N_3798,N_2775);
and U5581 (N_5581,N_3539,N_3686);
and U5582 (N_5582,N_3632,N_3666);
or U5583 (N_5583,N_4757,N_4638);
xnor U5584 (N_5584,N_4403,N_2654);
nor U5585 (N_5585,N_4162,N_3889);
and U5586 (N_5586,N_4752,N_3753);
nor U5587 (N_5587,N_4764,N_2683);
nand U5588 (N_5588,N_4546,N_4712);
xor U5589 (N_5589,N_3763,N_3994);
and U5590 (N_5590,N_3394,N_3627);
nand U5591 (N_5591,N_3940,N_3990);
nor U5592 (N_5592,N_3263,N_3029);
and U5593 (N_5593,N_4835,N_3866);
nor U5594 (N_5594,N_3642,N_4092);
and U5595 (N_5595,N_4541,N_2550);
xor U5596 (N_5596,N_4686,N_4654);
or U5597 (N_5597,N_3459,N_3702);
nor U5598 (N_5598,N_3299,N_4507);
xnor U5599 (N_5599,N_3287,N_4024);
and U5600 (N_5600,N_3189,N_4447);
nand U5601 (N_5601,N_4544,N_4516);
nor U5602 (N_5602,N_2621,N_4789);
and U5603 (N_5603,N_3727,N_2702);
nand U5604 (N_5604,N_3365,N_4864);
nand U5605 (N_5605,N_3967,N_3758);
xnor U5606 (N_5606,N_3164,N_2553);
nand U5607 (N_5607,N_3291,N_3095);
nor U5608 (N_5608,N_3280,N_2875);
and U5609 (N_5609,N_3182,N_3801);
nor U5610 (N_5610,N_4449,N_3621);
nand U5611 (N_5611,N_2658,N_3040);
xor U5612 (N_5612,N_3106,N_3318);
nand U5613 (N_5613,N_4404,N_3298);
nor U5614 (N_5614,N_4450,N_4611);
nor U5615 (N_5615,N_2548,N_3278);
nand U5616 (N_5616,N_2724,N_3616);
xor U5617 (N_5617,N_3526,N_3681);
nand U5618 (N_5618,N_2526,N_2786);
nand U5619 (N_5619,N_2847,N_4927);
nor U5620 (N_5620,N_3231,N_4093);
or U5621 (N_5621,N_4432,N_4585);
xor U5622 (N_5622,N_2762,N_4525);
xor U5623 (N_5623,N_3991,N_2528);
nand U5624 (N_5624,N_2970,N_4528);
and U5625 (N_5625,N_2712,N_2888);
nor U5626 (N_5626,N_2902,N_3586);
nand U5627 (N_5627,N_3575,N_3001);
and U5628 (N_5628,N_2555,N_3843);
or U5629 (N_5629,N_3872,N_4586);
and U5630 (N_5630,N_4916,N_4677);
xnor U5631 (N_5631,N_4593,N_3879);
and U5632 (N_5632,N_2503,N_3160);
or U5633 (N_5633,N_4790,N_4224);
or U5634 (N_5634,N_4986,N_3202);
nor U5635 (N_5635,N_4128,N_4958);
or U5636 (N_5636,N_4243,N_2669);
and U5637 (N_5637,N_3197,N_3323);
xnor U5638 (N_5638,N_3738,N_4555);
nand U5639 (N_5639,N_4880,N_3251);
or U5640 (N_5640,N_4847,N_4815);
nor U5641 (N_5641,N_2722,N_4941);
nand U5642 (N_5642,N_2559,N_4996);
or U5643 (N_5643,N_4718,N_3178);
nand U5644 (N_5644,N_3041,N_3731);
xnor U5645 (N_5645,N_3038,N_4452);
or U5646 (N_5646,N_4731,N_4480);
nor U5647 (N_5647,N_4918,N_2951);
or U5648 (N_5648,N_4523,N_3664);
and U5649 (N_5649,N_3894,N_3871);
nor U5650 (N_5650,N_3851,N_4548);
nand U5651 (N_5651,N_4081,N_2770);
and U5652 (N_5652,N_2761,N_3230);
nor U5653 (N_5653,N_3512,N_3882);
or U5654 (N_5654,N_3699,N_3744);
xnor U5655 (N_5655,N_4376,N_2789);
nand U5656 (N_5656,N_2571,N_2958);
nand U5657 (N_5657,N_3906,N_4075);
and U5658 (N_5658,N_3672,N_2854);
or U5659 (N_5659,N_3679,N_3349);
nor U5660 (N_5660,N_4603,N_3265);
nor U5661 (N_5661,N_3398,N_4348);
and U5662 (N_5662,N_3716,N_3873);
or U5663 (N_5663,N_2870,N_3800);
and U5664 (N_5664,N_3936,N_3312);
nand U5665 (N_5665,N_3572,N_4413);
nand U5666 (N_5666,N_3793,N_4263);
nand U5667 (N_5667,N_4981,N_2865);
nor U5668 (N_5668,N_3168,N_4824);
or U5669 (N_5669,N_4802,N_2863);
xnor U5670 (N_5670,N_2640,N_3375);
and U5671 (N_5671,N_4059,N_2691);
or U5672 (N_5672,N_3153,N_4350);
xnor U5673 (N_5673,N_2541,N_4818);
and U5674 (N_5674,N_2796,N_3649);
nand U5675 (N_5675,N_4647,N_4340);
and U5676 (N_5676,N_3691,N_3022);
or U5677 (N_5677,N_2678,N_4139);
and U5678 (N_5678,N_4454,N_4320);
or U5679 (N_5679,N_2728,N_4936);
xor U5680 (N_5680,N_2578,N_4019);
and U5681 (N_5681,N_3495,N_3783);
xnor U5682 (N_5682,N_4855,N_3198);
xnor U5683 (N_5683,N_4292,N_3771);
xnor U5684 (N_5684,N_4353,N_2930);
xor U5685 (N_5685,N_4895,N_2772);
nand U5686 (N_5686,N_4522,N_2864);
or U5687 (N_5687,N_3020,N_2861);
nor U5688 (N_5688,N_4175,N_3036);
and U5689 (N_5689,N_4227,N_3462);
nand U5690 (N_5690,N_3134,N_3532);
nor U5691 (N_5691,N_4821,N_3982);
xor U5692 (N_5692,N_4445,N_3012);
nor U5693 (N_5693,N_4108,N_2690);
xnor U5694 (N_5694,N_3493,N_3923);
nand U5695 (N_5695,N_3751,N_3184);
nand U5696 (N_5696,N_3497,N_4751);
nand U5697 (N_5697,N_4840,N_4464);
nand U5698 (N_5698,N_3893,N_4576);
nand U5699 (N_5699,N_4349,N_4239);
xnor U5700 (N_5700,N_4021,N_2830);
nand U5701 (N_5701,N_4261,N_4434);
xnor U5702 (N_5702,N_2711,N_3140);
nand U5703 (N_5703,N_4153,N_3809);
xor U5704 (N_5704,N_4422,N_4520);
xnor U5705 (N_5705,N_3465,N_4362);
or U5706 (N_5706,N_3279,N_4867);
or U5707 (N_5707,N_2986,N_3839);
nor U5708 (N_5708,N_3496,N_2591);
nand U5709 (N_5709,N_4769,N_4293);
and U5710 (N_5710,N_2646,N_3819);
or U5711 (N_5711,N_3188,N_4238);
nor U5712 (N_5712,N_2852,N_4184);
xnor U5713 (N_5713,N_3043,N_3007);
and U5714 (N_5714,N_4794,N_3315);
or U5715 (N_5715,N_4455,N_3992);
nand U5716 (N_5716,N_4940,N_4154);
or U5717 (N_5717,N_3359,N_4841);
nand U5718 (N_5718,N_4547,N_4494);
or U5719 (N_5719,N_3289,N_4039);
nor U5720 (N_5720,N_3530,N_4341);
nor U5721 (N_5721,N_4928,N_4708);
or U5722 (N_5722,N_4015,N_4816);
nand U5723 (N_5723,N_4155,N_4465);
xor U5724 (N_5724,N_3733,N_4572);
nand U5725 (N_5725,N_2891,N_2972);
xnor U5726 (N_5726,N_2779,N_2968);
nor U5727 (N_5727,N_3543,N_4459);
nand U5728 (N_5728,N_4639,N_4314);
and U5729 (N_5729,N_2582,N_4688);
and U5730 (N_5730,N_4729,N_4491);
xnor U5731 (N_5731,N_3201,N_2636);
or U5732 (N_5732,N_3482,N_2954);
nand U5733 (N_5733,N_4041,N_4266);
or U5734 (N_5734,N_3239,N_2670);
and U5735 (N_5735,N_2579,N_3546);
and U5736 (N_5736,N_2685,N_2703);
and U5737 (N_5737,N_3985,N_4166);
or U5738 (N_5738,N_4619,N_3369);
xnor U5739 (N_5739,N_3927,N_4247);
nand U5740 (N_5740,N_4046,N_3064);
nor U5741 (N_5741,N_3259,N_3461);
and U5742 (N_5742,N_4475,N_3589);
xnor U5743 (N_5743,N_3217,N_2983);
or U5744 (N_5744,N_2522,N_3919);
or U5745 (N_5745,N_2829,N_4765);
nand U5746 (N_5746,N_2536,N_3861);
nor U5747 (N_5747,N_2843,N_2592);
nand U5748 (N_5748,N_4557,N_4386);
and U5749 (N_5749,N_4926,N_2709);
nor U5750 (N_5750,N_2876,N_4930);
and U5751 (N_5751,N_4668,N_3186);
nor U5752 (N_5752,N_4705,N_2668);
nand U5753 (N_5753,N_3058,N_4302);
or U5754 (N_5754,N_4369,N_3097);
or U5755 (N_5755,N_2962,N_2660);
or U5756 (N_5756,N_3761,N_4827);
xnor U5757 (N_5757,N_2710,N_2811);
and U5758 (N_5758,N_3781,N_2600);
and U5759 (N_5759,N_3870,N_4387);
nand U5760 (N_5760,N_3458,N_2766);
xor U5761 (N_5761,N_3484,N_2667);
xnor U5762 (N_5762,N_4191,N_4748);
and U5763 (N_5763,N_3227,N_2984);
nor U5764 (N_5764,N_3238,N_4038);
nand U5765 (N_5765,N_4788,N_3104);
or U5766 (N_5766,N_4210,N_4307);
nand U5767 (N_5767,N_3537,N_4356);
xor U5768 (N_5768,N_2801,N_4563);
nand U5769 (N_5769,N_3220,N_2810);
and U5770 (N_5770,N_4923,N_2802);
nor U5771 (N_5771,N_4412,N_3515);
nor U5772 (N_5772,N_3017,N_3721);
or U5773 (N_5773,N_2919,N_4000);
nand U5774 (N_5774,N_2907,N_2622);
or U5775 (N_5775,N_4598,N_4870);
nor U5776 (N_5776,N_4924,N_4062);
xnor U5777 (N_5777,N_2788,N_4468);
and U5778 (N_5778,N_2868,N_4031);
and U5779 (N_5779,N_4913,N_3559);
nand U5780 (N_5780,N_2896,N_3110);
nor U5781 (N_5781,N_4749,N_3931);
nand U5782 (N_5782,N_3214,N_3556);
nor U5783 (N_5783,N_2747,N_3439);
nand U5784 (N_5784,N_4321,N_3371);
or U5785 (N_5785,N_3300,N_4235);
or U5786 (N_5786,N_3703,N_4989);
xor U5787 (N_5787,N_4086,N_3329);
nor U5788 (N_5788,N_4545,N_4192);
xor U5789 (N_5789,N_4583,N_4670);
nand U5790 (N_5790,N_2820,N_4357);
or U5791 (N_5791,N_3645,N_4020);
nor U5792 (N_5792,N_4543,N_2506);
nand U5793 (N_5793,N_3831,N_4866);
and U5794 (N_5794,N_3585,N_4457);
nor U5795 (N_5795,N_2531,N_3221);
xnor U5796 (N_5796,N_4231,N_4953);
nand U5797 (N_5797,N_4097,N_4112);
nand U5798 (N_5798,N_2742,N_4837);
nand U5799 (N_5799,N_4817,N_2734);
xor U5800 (N_5800,N_3196,N_3373);
or U5801 (N_5801,N_3655,N_3285);
xnor U5802 (N_5802,N_3382,N_3151);
or U5803 (N_5803,N_4490,N_2626);
xnor U5804 (N_5804,N_2635,N_4066);
and U5805 (N_5805,N_4566,N_2652);
or U5806 (N_5806,N_2611,N_4510);
nor U5807 (N_5807,N_3325,N_3922);
nand U5808 (N_5808,N_4983,N_3764);
or U5809 (N_5809,N_4331,N_3283);
or U5810 (N_5810,N_2677,N_3820);
xor U5811 (N_5811,N_4363,N_3939);
or U5812 (N_5812,N_3808,N_3380);
nor U5813 (N_5813,N_2827,N_2877);
xnor U5814 (N_5814,N_4629,N_4479);
xor U5815 (N_5815,N_3161,N_4506);
nand U5816 (N_5816,N_3584,N_4630);
xnor U5817 (N_5817,N_4589,N_4407);
and U5818 (N_5818,N_3191,N_3558);
nor U5819 (N_5819,N_3433,N_4704);
nor U5820 (N_5820,N_4268,N_2673);
nor U5821 (N_5821,N_4695,N_3812);
nor U5822 (N_5822,N_3941,N_3477);
and U5823 (N_5823,N_3335,N_3926);
xor U5824 (N_5824,N_3774,N_3951);
and U5825 (N_5825,N_4195,N_3430);
nand U5826 (N_5826,N_4240,N_3388);
or U5827 (N_5827,N_4262,N_4899);
or U5828 (N_5828,N_2634,N_4618);
or U5829 (N_5829,N_3674,N_4005);
nand U5830 (N_5830,N_4018,N_2508);
and U5831 (N_5831,N_4786,N_3792);
or U5832 (N_5832,N_4975,N_3334);
nor U5833 (N_5833,N_4651,N_3609);
xor U5834 (N_5834,N_2607,N_4284);
and U5835 (N_5835,N_4698,N_4096);
and U5836 (N_5836,N_4740,N_4846);
or U5837 (N_5837,N_4634,N_2860);
or U5838 (N_5838,N_4594,N_4897);
nand U5839 (N_5839,N_3177,N_3107);
xnor U5840 (N_5840,N_3682,N_4613);
and U5841 (N_5841,N_4201,N_3485);
xor U5842 (N_5842,N_4312,N_2965);
xor U5843 (N_5843,N_4373,N_3925);
and U5844 (N_5844,N_3660,N_2776);
or U5845 (N_5845,N_3975,N_4158);
xor U5846 (N_5846,N_4207,N_3974);
or U5847 (N_5847,N_2858,N_2926);
or U5848 (N_5848,N_2749,N_3704);
and U5849 (N_5849,N_2726,N_4596);
or U5850 (N_5850,N_3663,N_3089);
xor U5851 (N_5851,N_3208,N_3307);
or U5852 (N_5852,N_2885,N_4697);
xnor U5853 (N_5853,N_4498,N_3577);
nand U5854 (N_5854,N_2733,N_2835);
or U5855 (N_5855,N_4759,N_3829);
or U5856 (N_5856,N_4907,N_4253);
nor U5857 (N_5857,N_4601,N_2900);
or U5858 (N_5858,N_4893,N_4733);
nor U5859 (N_5859,N_4197,N_2679);
or U5860 (N_5860,N_4859,N_3708);
nor U5861 (N_5861,N_4783,N_4600);
nand U5862 (N_5862,N_3737,N_3418);
and U5863 (N_5863,N_2878,N_4437);
xnor U5864 (N_5864,N_4466,N_3412);
nor U5865 (N_5865,N_4013,N_3137);
nand U5866 (N_5866,N_3950,N_3301);
or U5867 (N_5867,N_3963,N_3739);
and U5868 (N_5868,N_3954,N_4993);
xor U5869 (N_5869,N_3065,N_4408);
and U5870 (N_5870,N_4842,N_3729);
and U5871 (N_5871,N_3914,N_3088);
or U5872 (N_5872,N_4414,N_3867);
nor U5873 (N_5873,N_2716,N_4898);
nand U5874 (N_5874,N_4389,N_4064);
or U5875 (N_5875,N_4805,N_2996);
or U5876 (N_5876,N_4565,N_3046);
nor U5877 (N_5877,N_3466,N_2982);
nand U5878 (N_5878,N_2979,N_4570);
and U5879 (N_5879,N_4470,N_3857);
or U5880 (N_5880,N_3395,N_4116);
nor U5881 (N_5881,N_4627,N_3223);
nor U5882 (N_5882,N_3364,N_3788);
nor U5883 (N_5883,N_3152,N_2808);
and U5884 (N_5884,N_3431,N_3434);
nand U5885 (N_5885,N_4592,N_4156);
or U5886 (N_5886,N_4965,N_2923);
xor U5887 (N_5887,N_3988,N_3159);
or U5888 (N_5888,N_4534,N_3514);
nand U5889 (N_5889,N_2872,N_3779);
nand U5890 (N_5890,N_3131,N_4602);
or U5891 (N_5891,N_4150,N_4087);
nor U5892 (N_5892,N_3835,N_3818);
nand U5893 (N_5893,N_2957,N_3869);
nand U5894 (N_5894,N_4508,N_4876);
or U5895 (N_5895,N_3204,N_4584);
nand U5896 (N_5896,N_4283,N_4439);
or U5897 (N_5897,N_3568,N_3638);
nand U5898 (N_5898,N_3724,N_2507);
nand U5899 (N_5899,N_3785,N_3784);
nand U5900 (N_5900,N_4151,N_4625);
and U5901 (N_5901,N_3331,N_4453);
nand U5902 (N_5902,N_2731,N_2931);
xnor U5903 (N_5903,N_3676,N_2975);
nand U5904 (N_5904,N_3234,N_2869);
or U5905 (N_5905,N_4987,N_4130);
nor U5906 (N_5906,N_4159,N_4662);
and U5907 (N_5907,N_3074,N_3544);
and U5908 (N_5908,N_2645,N_4099);
xnor U5909 (N_5909,N_2739,N_4234);
and U5910 (N_5910,N_4512,N_4865);
xnor U5911 (N_5911,N_3834,N_4669);
nor U5912 (N_5912,N_3491,N_2943);
nand U5913 (N_5913,N_2800,N_3333);
nand U5914 (N_5914,N_3213,N_2906);
and U5915 (N_5915,N_2518,N_2619);
xnor U5916 (N_5916,N_2809,N_4956);
nor U5917 (N_5917,N_4014,N_3720);
nand U5918 (N_5918,N_3341,N_3995);
nor U5919 (N_5919,N_4488,N_3746);
nand U5920 (N_5920,N_2544,N_3778);
xor U5921 (N_5921,N_3791,N_4067);
or U5922 (N_5922,N_3091,N_4218);
nand U5923 (N_5923,N_3499,N_3379);
nor U5924 (N_5924,N_3340,N_4823);
nor U5925 (N_5925,N_3910,N_3736);
or U5926 (N_5926,N_2575,N_4056);
nor U5927 (N_5927,N_4448,N_4255);
nand U5928 (N_5928,N_4727,N_3302);
nor U5929 (N_5929,N_3069,N_2509);
or U5930 (N_5930,N_4550,N_4028);
and U5931 (N_5931,N_3877,N_4444);
nor U5932 (N_5932,N_3440,N_4042);
xnor U5933 (N_5933,N_4135,N_3448);
or U5934 (N_5934,N_3255,N_3120);
nor U5935 (N_5935,N_4542,N_4297);
xor U5936 (N_5936,N_2823,N_2684);
or U5937 (N_5937,N_3171,N_2530);
nand U5938 (N_5938,N_2880,N_3697);
or U5939 (N_5939,N_2988,N_3425);
and U5940 (N_5940,N_2795,N_4161);
or U5941 (N_5941,N_3000,N_3195);
or U5942 (N_5942,N_4164,N_3145);
or U5943 (N_5943,N_4332,N_4057);
xnor U5944 (N_5944,N_3907,N_4745);
and U5945 (N_5945,N_4896,N_3414);
or U5946 (N_5946,N_4978,N_2625);
or U5947 (N_5947,N_2721,N_2916);
nand U5948 (N_5948,N_3409,N_2782);
nand U5949 (N_5949,N_4937,N_3266);
nand U5950 (N_5950,N_3028,N_2504);
nor U5951 (N_5951,N_2502,N_4360);
nor U5952 (N_5952,N_2675,N_3999);
xor U5953 (N_5953,N_2704,N_3890);
or U5954 (N_5954,N_2767,N_2780);
nand U5955 (N_5955,N_4901,N_2853);
or U5956 (N_5956,N_4980,N_2564);
nor U5957 (N_5957,N_2593,N_3406);
nand U5958 (N_5958,N_4706,N_3921);
or U5959 (N_5959,N_3811,N_2783);
xor U5960 (N_5960,N_3952,N_3750);
nand U5961 (N_5961,N_4990,N_2914);
nor U5962 (N_5962,N_4143,N_4110);
nor U5963 (N_5963,N_3578,N_4351);
xor U5964 (N_5964,N_3157,N_4190);
or U5965 (N_5965,N_4626,N_2998);
nand U5966 (N_5966,N_3651,N_3117);
nor U5967 (N_5967,N_3267,N_3072);
and U5968 (N_5968,N_3216,N_3488);
or U5969 (N_5969,N_3528,N_3671);
nand U5970 (N_5970,N_4225,N_3842);
xnor U5971 (N_5971,N_4881,N_3957);
and U5972 (N_5972,N_3971,N_3410);
nor U5973 (N_5973,N_3428,N_2818);
xor U5974 (N_5974,N_3806,N_4251);
xnor U5975 (N_5975,N_3522,N_3086);
xnor U5976 (N_5976,N_2948,N_4920);
xor U5977 (N_5977,N_4949,N_4442);
nor U5978 (N_5978,N_2831,N_2781);
nand U5979 (N_5979,N_4684,N_4285);
or U5980 (N_5980,N_2672,N_4784);
nor U5981 (N_5981,N_3228,N_4065);
and U5982 (N_5982,N_4558,N_3356);
or U5983 (N_5983,N_3517,N_4322);
and U5984 (N_5984,N_3937,N_2940);
nor U5985 (N_5985,N_3362,N_3446);
and U5986 (N_5986,N_3303,N_3346);
or U5987 (N_5987,N_3068,N_4026);
nor U5988 (N_5988,N_3473,N_2913);
and U5989 (N_5989,N_3033,N_4134);
and U5990 (N_5990,N_3205,N_4394);
xnor U5991 (N_5991,N_4645,N_3321);
xor U5992 (N_5992,N_2725,N_2519);
xnor U5993 (N_5993,N_3139,N_4486);
nor U5994 (N_5994,N_4787,N_4009);
xor U5995 (N_5995,N_3063,N_3008);
or U5996 (N_5996,N_3174,N_4878);
xnor U5997 (N_5997,N_2647,N_4233);
nand U5998 (N_5998,N_3219,N_4974);
nand U5999 (N_5999,N_4365,N_3620);
and U6000 (N_6000,N_3569,N_4657);
or U6001 (N_6001,N_3840,N_2751);
or U6002 (N_6002,N_4478,N_2757);
and U6003 (N_6003,N_2915,N_2715);
or U6004 (N_6004,N_4868,N_4902);
nand U6005 (N_6005,N_4530,N_3654);
and U6006 (N_6006,N_3903,N_3665);
or U6007 (N_6007,N_2949,N_3248);
or U6008 (N_6008,N_2844,N_4068);
or U6009 (N_6009,N_2784,N_4214);
nand U6010 (N_6010,N_3419,N_4681);
or U6011 (N_6011,N_3601,N_3393);
nand U6012 (N_6012,N_3276,N_4995);
and U6013 (N_6013,N_4221,N_3782);
or U6014 (N_6014,N_4236,N_3118);
and U6015 (N_6015,N_4732,N_3984);
xor U6016 (N_6016,N_4275,N_4259);
xor U6017 (N_6017,N_4122,N_4299);
and U6018 (N_6018,N_3525,N_4313);
and U6019 (N_6019,N_4012,N_3757);
or U6020 (N_6020,N_3658,N_3456);
and U6021 (N_6021,N_3956,N_3143);
or U6022 (N_6022,N_4760,N_3471);
xor U6023 (N_6023,N_3550,N_3920);
and U6024 (N_6024,N_2787,N_2601);
or U6025 (N_6025,N_4074,N_3797);
xor U6026 (N_6026,N_4659,N_2961);
nor U6027 (N_6027,N_3011,N_3185);
nor U6028 (N_6028,N_2834,N_4850);
and U6029 (N_6029,N_3680,N_2859);
or U6030 (N_6030,N_2686,N_4270);
and U6031 (N_6031,N_2997,N_4286);
xor U6032 (N_6032,N_4111,N_2708);
nor U6033 (N_6033,N_3696,N_4552);
or U6034 (N_6034,N_4678,N_4564);
nor U6035 (N_6035,N_3146,N_4222);
nor U6036 (N_6036,N_3286,N_3474);
or U6037 (N_6037,N_2771,N_4215);
and U6038 (N_6038,N_4915,N_4489);
nand U6039 (N_6039,N_2584,N_4189);
nand U6040 (N_6040,N_4909,N_3613);
and U6041 (N_6041,N_4004,N_3486);
nor U6042 (N_6042,N_3417,N_2706);
xor U6043 (N_6043,N_3610,N_4423);
nor U6044 (N_6044,N_4371,N_2653);
nor U6045 (N_6045,N_2950,N_4289);
or U6046 (N_6046,N_3510,N_2871);
or U6047 (N_6047,N_4887,N_3823);
and U6048 (N_6048,N_3500,N_2523);
nand U6049 (N_6049,N_4280,N_2577);
and U6050 (N_6050,N_2851,N_2623);
and U6051 (N_6051,N_3892,N_2881);
nor U6052 (N_6052,N_4274,N_2765);
and U6053 (N_6053,N_2793,N_3154);
nand U6054 (N_6054,N_3648,N_4380);
nand U6055 (N_6055,N_4944,N_4680);
xnor U6056 (N_6056,N_2879,N_4998);
xor U6057 (N_6057,N_3594,N_2763);
and U6058 (N_6058,N_4072,N_3580);
nor U6059 (N_6059,N_4055,N_3077);
and U6060 (N_6060,N_4497,N_4720);
nor U6061 (N_6061,N_3116,N_4730);
or U6062 (N_6062,N_3847,N_2819);
and U6063 (N_6063,N_2814,N_4461);
xnor U6064 (N_6064,N_4132,N_3158);
nor U6065 (N_6065,N_4346,N_4991);
xnor U6066 (N_6066,N_3582,N_2723);
or U6067 (N_6067,N_4696,N_2657);
or U6068 (N_6068,N_4186,N_2971);
nor U6069 (N_6069,N_3535,N_4992);
xnor U6070 (N_6070,N_3438,N_3119);
xor U6071 (N_6071,N_4675,N_3918);
and U6072 (N_6072,N_4071,N_2565);
nand U6073 (N_6073,N_4988,N_2655);
nand U6074 (N_6074,N_4742,N_2894);
nor U6075 (N_6075,N_3237,N_2620);
nor U6076 (N_6076,N_2513,N_4617);
xnor U6077 (N_6077,N_4933,N_3643);
nand U6078 (N_6078,N_3060,N_4120);
and U6079 (N_6079,N_4070,N_2908);
xnor U6080 (N_6080,N_3389,N_3848);
nand U6081 (N_6081,N_2774,N_4493);
xor U6082 (N_6082,N_3035,N_4202);
xnor U6083 (N_6083,N_3542,N_3625);
xnor U6084 (N_6084,N_3745,N_2613);
nor U6085 (N_6085,N_2604,N_3222);
nand U6086 (N_6086,N_4347,N_2510);
and U6087 (N_6087,N_2537,N_3144);
or U6088 (N_6088,N_3233,N_4517);
nor U6089 (N_6089,N_4621,N_4061);
or U6090 (N_6090,N_2921,N_3787);
and U6091 (N_6091,N_2748,N_3884);
nor U6092 (N_6092,N_2813,N_3155);
and U6093 (N_6093,N_3908,N_3976);
or U6094 (N_6094,N_4922,N_4427);
nand U6095 (N_6095,N_4032,N_4300);
nand U6096 (N_6096,N_2740,N_4163);
and U6097 (N_6097,N_4713,N_3675);
xnor U6098 (N_6098,N_4344,N_3378);
nor U6099 (N_6099,N_3460,N_4430);
nand U6100 (N_6100,N_4518,N_3254);
xor U6101 (N_6101,N_3946,N_4106);
nor U6102 (N_6102,N_3631,N_4100);
nor U6103 (N_6103,N_4969,N_3306);
and U6104 (N_6104,N_4652,N_3735);
nor U6105 (N_6105,N_2674,N_3570);
or U6106 (N_6106,N_3297,N_4250);
nand U6107 (N_6107,N_2573,N_3766);
nor U6108 (N_6108,N_4188,N_3066);
or U6109 (N_6109,N_2928,N_4094);
nand U6110 (N_6110,N_3050,N_4180);
nand U6111 (N_6111,N_2838,N_2576);
nand U6112 (N_6112,N_2937,N_3338);
xnor U6113 (N_6113,N_3566,N_3755);
or U6114 (N_6114,N_3175,N_3166);
and U6115 (N_6115,N_4780,N_3740);
nor U6116 (N_6116,N_4575,N_2567);
or U6117 (N_6117,N_3777,N_4267);
or U6118 (N_6118,N_4691,N_4702);
nand U6119 (N_6119,N_3026,N_3274);
nor U6120 (N_6120,N_4138,N_4194);
and U6121 (N_6121,N_2569,N_2833);
nand U6122 (N_6122,N_3105,N_2651);
and U6123 (N_6123,N_4801,N_2964);
nand U6124 (N_6124,N_4672,N_3741);
nor U6125 (N_6125,N_4343,N_3885);
xnor U6126 (N_6126,N_4529,N_4368);
and U6127 (N_6127,N_2540,N_4531);
nand U6128 (N_6128,N_4260,N_2521);
nor U6129 (N_6129,N_4352,N_3911);
and U6130 (N_6130,N_3109,N_3272);
or U6131 (N_6131,N_4591,N_3966);
and U6132 (N_6132,N_3067,N_4405);
xnor U6133 (N_6133,N_4157,N_4118);
nand U6134 (N_6134,N_3403,N_3905);
and U6135 (N_6135,N_4939,N_4808);
or U6136 (N_6136,N_3534,N_3611);
nand U6137 (N_6137,N_2759,N_4374);
nor U6138 (N_6138,N_3997,N_4571);
xnor U6139 (N_6139,N_3429,N_4193);
nand U6140 (N_6140,N_3760,N_4725);
nand U6141 (N_6141,N_3115,N_3368);
xnor U6142 (N_6142,N_2527,N_4208);
xnor U6143 (N_6143,N_4860,N_4873);
nand U6144 (N_6144,N_3070,N_3707);
nor U6145 (N_6145,N_2500,N_2505);
xnor U6146 (N_6146,N_4830,N_3796);
and U6147 (N_6147,N_3494,N_4040);
xnor U6148 (N_6148,N_3320,N_3603);
and U6149 (N_6149,N_4174,N_2561);
nor U6150 (N_6150,N_3083,N_4582);
nand U6151 (N_6151,N_4785,N_4766);
nand U6152 (N_6152,N_3527,N_4375);
or U6153 (N_6153,N_3296,N_2586);
or U6154 (N_6154,N_3481,N_3706);
or U6155 (N_6155,N_4098,N_4848);
and U6156 (N_6156,N_4406,N_3554);
xor U6157 (N_6157,N_2517,N_2899);
xor U6158 (N_6158,N_3436,N_3955);
xor U6159 (N_6159,N_3354,N_3200);
nor U6160 (N_6160,N_4359,N_2941);
nor U6161 (N_6161,N_3324,N_4853);
or U6162 (N_6162,N_3519,N_2597);
nor U6163 (N_6163,N_3562,N_3010);
and U6164 (N_6164,N_4768,N_4438);
or U6165 (N_6165,N_3833,N_3179);
and U6166 (N_6166,N_4536,N_3108);
or U6167 (N_6167,N_2911,N_4964);
nand U6168 (N_6168,N_4524,N_3199);
nor U6169 (N_6169,N_4636,N_3898);
nand U6170 (N_6170,N_3977,N_3548);
nor U6171 (N_6171,N_3402,N_3015);
and U6172 (N_6172,N_2587,N_2663);
nand U6173 (N_6173,N_3719,N_4693);
and U6174 (N_6174,N_4791,N_4537);
and U6175 (N_6175,N_2543,N_4806);
nand U6176 (N_6176,N_4428,N_2769);
nor U6177 (N_6177,N_3260,N_3874);
nor U6178 (N_6178,N_4554,N_3881);
or U6179 (N_6179,N_4206,N_3862);
nor U6180 (N_6180,N_2901,N_4648);
nor U6181 (N_6181,N_2840,N_3883);
or U6182 (N_6182,N_4738,N_3989);
or U6183 (N_6183,N_3647,N_3262);
nor U6184 (N_6184,N_4358,N_4623);
and U6185 (N_6185,N_3416,N_3357);
or U6186 (N_6186,N_3469,N_4800);
or U6187 (N_6187,N_2978,N_2570);
nand U6188 (N_6188,N_3944,N_4364);
xor U6189 (N_6189,N_3256,N_4063);
xnor U6190 (N_6190,N_2892,N_3444);
xor U6191 (N_6191,N_3770,N_3599);
xnor U6192 (N_6192,N_4653,N_3075);
xor U6193 (N_6193,N_3507,N_4761);
nand U6194 (N_6194,N_3071,N_4900);
nand U6195 (N_6195,N_4334,N_3773);
nor U6196 (N_6196,N_3612,N_3292);
nor U6197 (N_6197,N_4767,N_3768);
and U6198 (N_6198,N_3215,N_4854);
and U6199 (N_6199,N_4165,N_4443);
xor U6200 (N_6200,N_3722,N_4912);
nand U6201 (N_6201,N_4030,N_4073);
xor U6202 (N_6202,N_4561,N_3293);
and U6203 (N_6203,N_2511,N_4282);
or U6204 (N_6204,N_4719,N_3180);
or U6205 (N_6205,N_3710,N_4035);
xor U6206 (N_6206,N_2993,N_4345);
nand U6207 (N_6207,N_3463,N_2741);
or U6208 (N_6208,N_4317,N_4199);
or U6209 (N_6209,N_3400,N_4264);
and U6210 (N_6210,N_4957,N_3384);
nor U6211 (N_6211,N_2893,N_2846);
or U6212 (N_6212,N_3061,N_4124);
or U6213 (N_6213,N_3132,N_4482);
xnor U6214 (N_6214,N_4308,N_2890);
and U6215 (N_6215,N_4689,N_4533);
and U6216 (N_6216,N_4080,N_4372);
or U6217 (N_6217,N_2966,N_4319);
nor U6218 (N_6218,N_3264,N_4431);
xor U6219 (N_6219,N_3273,N_4329);
and U6220 (N_6220,N_4276,N_3506);
or U6221 (N_6221,N_3193,N_4632);
xor U6222 (N_6222,N_3852,N_4388);
or U6223 (N_6223,N_4942,N_4296);
nor U6224 (N_6224,N_2596,N_2532);
nor U6225 (N_6225,N_3049,N_4836);
nand U6226 (N_6226,N_3769,N_3912);
nand U6227 (N_6227,N_4200,N_4908);
xor U6228 (N_6228,N_3786,N_4797);
nor U6229 (N_6229,N_3973,N_4033);
and U6230 (N_6230,N_2551,N_2516);
nand U6231 (N_6231,N_2585,N_4798);
or U6232 (N_6232,N_4703,N_4869);
and U6233 (N_6233,N_3464,N_4921);
xnor U6234 (N_6234,N_4181,N_3344);
xnor U6235 (N_6235,N_3701,N_4361);
nand U6236 (N_6236,N_3277,N_3715);
nor U6237 (N_6237,N_4147,N_4230);
nor U6238 (N_6238,N_2889,N_2692);
or U6239 (N_6239,N_3039,N_4007);
xor U6240 (N_6240,N_4078,N_4295);
nor U6241 (N_6241,N_4133,N_4149);
and U6242 (N_6242,N_3960,N_3598);
nor U6243 (N_6243,N_4655,N_4503);
xor U6244 (N_6244,N_4309,N_3042);
or U6245 (N_6245,N_4229,N_4883);
nand U6246 (N_6246,N_2804,N_3916);
or U6247 (N_6247,N_3062,N_4573);
or U6248 (N_6248,N_2713,N_3250);
nand U6249 (N_6249,N_2944,N_4660);
nand U6250 (N_6250,N_2996,N_4337);
nand U6251 (N_6251,N_3945,N_4342);
or U6252 (N_6252,N_2716,N_2602);
and U6253 (N_6253,N_2623,N_3179);
and U6254 (N_6254,N_3390,N_2589);
nor U6255 (N_6255,N_2632,N_2839);
nor U6256 (N_6256,N_4608,N_2957);
nand U6257 (N_6257,N_4075,N_3029);
nor U6258 (N_6258,N_3664,N_3794);
and U6259 (N_6259,N_3855,N_2790);
and U6260 (N_6260,N_3199,N_3720);
and U6261 (N_6261,N_4631,N_4420);
nor U6262 (N_6262,N_4820,N_2714);
xor U6263 (N_6263,N_2822,N_3634);
xor U6264 (N_6264,N_3450,N_4202);
or U6265 (N_6265,N_4640,N_3423);
xnor U6266 (N_6266,N_3645,N_4278);
xnor U6267 (N_6267,N_3178,N_4271);
nand U6268 (N_6268,N_2915,N_4391);
or U6269 (N_6269,N_3345,N_4925);
nor U6270 (N_6270,N_4457,N_2561);
nand U6271 (N_6271,N_4605,N_3411);
or U6272 (N_6272,N_3410,N_3327);
nand U6273 (N_6273,N_4841,N_3897);
or U6274 (N_6274,N_3340,N_3251);
nand U6275 (N_6275,N_4527,N_4484);
and U6276 (N_6276,N_3446,N_4671);
and U6277 (N_6277,N_4250,N_3157);
nor U6278 (N_6278,N_2590,N_2754);
nand U6279 (N_6279,N_4104,N_2968);
nand U6280 (N_6280,N_4515,N_4843);
and U6281 (N_6281,N_3851,N_4732);
xor U6282 (N_6282,N_2534,N_4869);
nor U6283 (N_6283,N_3819,N_3905);
nor U6284 (N_6284,N_3423,N_3578);
nand U6285 (N_6285,N_4378,N_3659);
and U6286 (N_6286,N_3548,N_3082);
xnor U6287 (N_6287,N_3724,N_4994);
xor U6288 (N_6288,N_4769,N_2557);
and U6289 (N_6289,N_3818,N_4872);
nand U6290 (N_6290,N_3346,N_2812);
or U6291 (N_6291,N_3051,N_4152);
xnor U6292 (N_6292,N_2599,N_2933);
and U6293 (N_6293,N_3551,N_3325);
xnor U6294 (N_6294,N_3203,N_4985);
and U6295 (N_6295,N_4975,N_4543);
nand U6296 (N_6296,N_3188,N_3716);
or U6297 (N_6297,N_3286,N_3594);
nand U6298 (N_6298,N_2679,N_3099);
xor U6299 (N_6299,N_4131,N_2932);
xnor U6300 (N_6300,N_3002,N_3089);
and U6301 (N_6301,N_4079,N_4977);
or U6302 (N_6302,N_3331,N_4702);
or U6303 (N_6303,N_2979,N_3350);
nor U6304 (N_6304,N_2830,N_4314);
nor U6305 (N_6305,N_2778,N_3951);
and U6306 (N_6306,N_3911,N_3499);
and U6307 (N_6307,N_4164,N_3364);
or U6308 (N_6308,N_4514,N_2974);
or U6309 (N_6309,N_4897,N_4617);
xor U6310 (N_6310,N_4455,N_3068);
nor U6311 (N_6311,N_2552,N_4762);
xnor U6312 (N_6312,N_3078,N_4143);
or U6313 (N_6313,N_4324,N_3652);
xor U6314 (N_6314,N_4193,N_4985);
or U6315 (N_6315,N_4266,N_4546);
or U6316 (N_6316,N_3710,N_4640);
and U6317 (N_6317,N_4534,N_3866);
and U6318 (N_6318,N_4000,N_3456);
and U6319 (N_6319,N_2665,N_2569);
xnor U6320 (N_6320,N_3918,N_4411);
or U6321 (N_6321,N_3208,N_4922);
nor U6322 (N_6322,N_3473,N_3770);
and U6323 (N_6323,N_4267,N_4274);
xnor U6324 (N_6324,N_3900,N_3354);
or U6325 (N_6325,N_4871,N_3000);
and U6326 (N_6326,N_4419,N_3737);
nor U6327 (N_6327,N_4694,N_4909);
and U6328 (N_6328,N_3966,N_3615);
and U6329 (N_6329,N_2698,N_3308);
nor U6330 (N_6330,N_3874,N_3157);
nor U6331 (N_6331,N_4373,N_3186);
xnor U6332 (N_6332,N_2774,N_4840);
and U6333 (N_6333,N_3983,N_3956);
nor U6334 (N_6334,N_3144,N_2607);
nand U6335 (N_6335,N_2938,N_4429);
and U6336 (N_6336,N_3904,N_3990);
nor U6337 (N_6337,N_4890,N_3958);
or U6338 (N_6338,N_4484,N_3225);
and U6339 (N_6339,N_3938,N_4533);
or U6340 (N_6340,N_2790,N_4062);
nand U6341 (N_6341,N_4637,N_2645);
and U6342 (N_6342,N_2663,N_3472);
xor U6343 (N_6343,N_4243,N_3053);
xor U6344 (N_6344,N_4552,N_3740);
and U6345 (N_6345,N_3190,N_4567);
or U6346 (N_6346,N_2580,N_2906);
xnor U6347 (N_6347,N_4578,N_3371);
or U6348 (N_6348,N_4630,N_3206);
and U6349 (N_6349,N_4836,N_3646);
nor U6350 (N_6350,N_4554,N_4850);
xnor U6351 (N_6351,N_4579,N_4455);
nand U6352 (N_6352,N_3232,N_3850);
or U6353 (N_6353,N_4855,N_4754);
or U6354 (N_6354,N_2876,N_3131);
or U6355 (N_6355,N_4707,N_3425);
nand U6356 (N_6356,N_3706,N_3307);
nand U6357 (N_6357,N_3532,N_2741);
nand U6358 (N_6358,N_4370,N_4094);
and U6359 (N_6359,N_3203,N_3373);
xor U6360 (N_6360,N_2765,N_4113);
and U6361 (N_6361,N_4614,N_3880);
xnor U6362 (N_6362,N_4976,N_3845);
xor U6363 (N_6363,N_4109,N_4082);
nand U6364 (N_6364,N_2688,N_3606);
xor U6365 (N_6365,N_4288,N_4881);
or U6366 (N_6366,N_4651,N_4306);
and U6367 (N_6367,N_4219,N_3466);
and U6368 (N_6368,N_4482,N_3466);
xor U6369 (N_6369,N_4722,N_4712);
nor U6370 (N_6370,N_2516,N_4311);
and U6371 (N_6371,N_4060,N_4405);
and U6372 (N_6372,N_2960,N_4534);
or U6373 (N_6373,N_3005,N_3794);
or U6374 (N_6374,N_3255,N_3533);
nor U6375 (N_6375,N_4057,N_4100);
and U6376 (N_6376,N_4307,N_4971);
nand U6377 (N_6377,N_4068,N_3346);
and U6378 (N_6378,N_3177,N_4598);
or U6379 (N_6379,N_4906,N_2844);
or U6380 (N_6380,N_4408,N_2873);
nor U6381 (N_6381,N_2519,N_2547);
or U6382 (N_6382,N_4668,N_3400);
nand U6383 (N_6383,N_4829,N_4783);
xor U6384 (N_6384,N_3974,N_3315);
xnor U6385 (N_6385,N_4570,N_3620);
or U6386 (N_6386,N_3974,N_4054);
nor U6387 (N_6387,N_2923,N_2632);
or U6388 (N_6388,N_4310,N_3304);
and U6389 (N_6389,N_4442,N_4410);
xor U6390 (N_6390,N_4392,N_3090);
or U6391 (N_6391,N_3876,N_3269);
nor U6392 (N_6392,N_2607,N_3619);
nand U6393 (N_6393,N_3132,N_4717);
and U6394 (N_6394,N_4452,N_2758);
and U6395 (N_6395,N_4604,N_3681);
nand U6396 (N_6396,N_3411,N_3739);
or U6397 (N_6397,N_3722,N_3113);
and U6398 (N_6398,N_3677,N_4411);
or U6399 (N_6399,N_4127,N_4270);
nor U6400 (N_6400,N_4264,N_3340);
or U6401 (N_6401,N_3586,N_3588);
and U6402 (N_6402,N_3948,N_2638);
nand U6403 (N_6403,N_3605,N_3234);
nor U6404 (N_6404,N_2978,N_2648);
or U6405 (N_6405,N_3495,N_3710);
and U6406 (N_6406,N_2664,N_3348);
xor U6407 (N_6407,N_3420,N_3086);
nor U6408 (N_6408,N_4248,N_4875);
xnor U6409 (N_6409,N_4123,N_3361);
and U6410 (N_6410,N_4529,N_3882);
or U6411 (N_6411,N_3322,N_2735);
nor U6412 (N_6412,N_3520,N_4092);
xor U6413 (N_6413,N_3598,N_4353);
and U6414 (N_6414,N_2668,N_3290);
nand U6415 (N_6415,N_2893,N_2797);
nand U6416 (N_6416,N_3370,N_4029);
xor U6417 (N_6417,N_3028,N_4610);
or U6418 (N_6418,N_3214,N_4424);
xor U6419 (N_6419,N_3065,N_4131);
xnor U6420 (N_6420,N_4538,N_4807);
and U6421 (N_6421,N_2751,N_3743);
nand U6422 (N_6422,N_2866,N_3695);
xor U6423 (N_6423,N_4067,N_3160);
nor U6424 (N_6424,N_4764,N_4084);
nand U6425 (N_6425,N_3524,N_4099);
or U6426 (N_6426,N_2577,N_3499);
nor U6427 (N_6427,N_4232,N_4674);
xor U6428 (N_6428,N_4410,N_2578);
or U6429 (N_6429,N_3045,N_3995);
or U6430 (N_6430,N_3038,N_3772);
nor U6431 (N_6431,N_4561,N_4127);
or U6432 (N_6432,N_4433,N_4814);
nor U6433 (N_6433,N_4747,N_4901);
or U6434 (N_6434,N_4855,N_2907);
nor U6435 (N_6435,N_4165,N_3387);
and U6436 (N_6436,N_2610,N_4326);
or U6437 (N_6437,N_2621,N_2933);
nand U6438 (N_6438,N_3547,N_3772);
and U6439 (N_6439,N_2542,N_3721);
nor U6440 (N_6440,N_3119,N_3545);
and U6441 (N_6441,N_2663,N_2908);
nand U6442 (N_6442,N_3554,N_3467);
xor U6443 (N_6443,N_2755,N_2801);
nor U6444 (N_6444,N_3098,N_3101);
xnor U6445 (N_6445,N_2969,N_3727);
and U6446 (N_6446,N_4347,N_3844);
xor U6447 (N_6447,N_4098,N_4285);
or U6448 (N_6448,N_3107,N_4435);
or U6449 (N_6449,N_3316,N_2572);
and U6450 (N_6450,N_2635,N_3212);
or U6451 (N_6451,N_4770,N_2624);
xor U6452 (N_6452,N_3380,N_3018);
or U6453 (N_6453,N_3041,N_3467);
and U6454 (N_6454,N_2728,N_3758);
nor U6455 (N_6455,N_4525,N_4785);
and U6456 (N_6456,N_2992,N_4320);
and U6457 (N_6457,N_3277,N_3615);
xnor U6458 (N_6458,N_4155,N_3226);
or U6459 (N_6459,N_3194,N_2590);
nand U6460 (N_6460,N_4777,N_3896);
nor U6461 (N_6461,N_4736,N_3139);
xor U6462 (N_6462,N_4492,N_4398);
xnor U6463 (N_6463,N_3868,N_3813);
nand U6464 (N_6464,N_3844,N_4549);
or U6465 (N_6465,N_4938,N_4225);
or U6466 (N_6466,N_3985,N_4377);
nand U6467 (N_6467,N_4017,N_3896);
xnor U6468 (N_6468,N_3555,N_2886);
nand U6469 (N_6469,N_3906,N_2743);
nor U6470 (N_6470,N_4304,N_4950);
or U6471 (N_6471,N_2814,N_4078);
or U6472 (N_6472,N_3720,N_3801);
and U6473 (N_6473,N_4726,N_2656);
xnor U6474 (N_6474,N_4883,N_4678);
nand U6475 (N_6475,N_4456,N_4989);
nor U6476 (N_6476,N_3724,N_3426);
or U6477 (N_6477,N_4087,N_2939);
and U6478 (N_6478,N_2619,N_3117);
and U6479 (N_6479,N_4993,N_3652);
nand U6480 (N_6480,N_4199,N_4221);
nand U6481 (N_6481,N_3938,N_4103);
or U6482 (N_6482,N_2953,N_4505);
xor U6483 (N_6483,N_2516,N_4817);
and U6484 (N_6484,N_3589,N_3177);
xnor U6485 (N_6485,N_3397,N_4118);
or U6486 (N_6486,N_3853,N_4367);
and U6487 (N_6487,N_4584,N_4723);
or U6488 (N_6488,N_2864,N_2817);
and U6489 (N_6489,N_2645,N_4319);
nand U6490 (N_6490,N_4851,N_2751);
xnor U6491 (N_6491,N_3905,N_2541);
xor U6492 (N_6492,N_3315,N_3665);
and U6493 (N_6493,N_2995,N_4570);
nor U6494 (N_6494,N_4683,N_4374);
nor U6495 (N_6495,N_4871,N_3170);
nor U6496 (N_6496,N_4320,N_4814);
xnor U6497 (N_6497,N_2642,N_2997);
xnor U6498 (N_6498,N_4076,N_4463);
and U6499 (N_6499,N_3111,N_2565);
nand U6500 (N_6500,N_3697,N_3954);
and U6501 (N_6501,N_3000,N_4181);
nor U6502 (N_6502,N_4104,N_2716);
nor U6503 (N_6503,N_4082,N_2764);
xnor U6504 (N_6504,N_3046,N_4508);
and U6505 (N_6505,N_3698,N_2626);
xnor U6506 (N_6506,N_2611,N_3899);
or U6507 (N_6507,N_2840,N_4763);
nand U6508 (N_6508,N_3929,N_2876);
or U6509 (N_6509,N_3925,N_4310);
or U6510 (N_6510,N_3708,N_4800);
nand U6511 (N_6511,N_4815,N_4379);
or U6512 (N_6512,N_4915,N_4466);
nand U6513 (N_6513,N_2893,N_3341);
nand U6514 (N_6514,N_3640,N_2723);
and U6515 (N_6515,N_3434,N_3274);
or U6516 (N_6516,N_4506,N_2980);
nand U6517 (N_6517,N_3660,N_4159);
or U6518 (N_6518,N_2659,N_4553);
nor U6519 (N_6519,N_4257,N_3886);
and U6520 (N_6520,N_4761,N_3573);
and U6521 (N_6521,N_2962,N_2679);
nor U6522 (N_6522,N_3085,N_4836);
and U6523 (N_6523,N_4553,N_3124);
and U6524 (N_6524,N_4444,N_3892);
or U6525 (N_6525,N_3828,N_4631);
or U6526 (N_6526,N_3627,N_3147);
xnor U6527 (N_6527,N_4603,N_4723);
xnor U6528 (N_6528,N_3855,N_4747);
or U6529 (N_6529,N_3648,N_4275);
nand U6530 (N_6530,N_2878,N_4422);
nand U6531 (N_6531,N_2760,N_3744);
and U6532 (N_6532,N_4201,N_4045);
nand U6533 (N_6533,N_4567,N_3370);
xnor U6534 (N_6534,N_4736,N_3177);
and U6535 (N_6535,N_2934,N_3485);
nand U6536 (N_6536,N_3810,N_4119);
and U6537 (N_6537,N_4561,N_3644);
xnor U6538 (N_6538,N_3543,N_3069);
nand U6539 (N_6539,N_4400,N_4164);
nor U6540 (N_6540,N_2823,N_3141);
and U6541 (N_6541,N_3662,N_3403);
nor U6542 (N_6542,N_3521,N_3080);
nand U6543 (N_6543,N_4733,N_3399);
xnor U6544 (N_6544,N_3322,N_4419);
and U6545 (N_6545,N_4615,N_4083);
or U6546 (N_6546,N_3610,N_4254);
nor U6547 (N_6547,N_4550,N_2898);
xnor U6548 (N_6548,N_3230,N_3104);
and U6549 (N_6549,N_4247,N_3012);
and U6550 (N_6550,N_3416,N_2632);
and U6551 (N_6551,N_4247,N_3471);
nand U6552 (N_6552,N_4483,N_2622);
or U6553 (N_6553,N_3078,N_2774);
nand U6554 (N_6554,N_4586,N_4860);
nand U6555 (N_6555,N_4110,N_2862);
nor U6556 (N_6556,N_3758,N_2985);
or U6557 (N_6557,N_3711,N_3497);
or U6558 (N_6558,N_4848,N_3291);
or U6559 (N_6559,N_2558,N_3287);
xnor U6560 (N_6560,N_3654,N_3382);
xnor U6561 (N_6561,N_4349,N_4761);
and U6562 (N_6562,N_4691,N_2964);
xor U6563 (N_6563,N_3757,N_4606);
nor U6564 (N_6564,N_3894,N_4432);
and U6565 (N_6565,N_3402,N_3035);
nand U6566 (N_6566,N_3047,N_4442);
and U6567 (N_6567,N_4537,N_4244);
xor U6568 (N_6568,N_4030,N_4540);
or U6569 (N_6569,N_2657,N_2659);
xnor U6570 (N_6570,N_3428,N_4774);
or U6571 (N_6571,N_4274,N_3156);
and U6572 (N_6572,N_3602,N_3429);
xor U6573 (N_6573,N_4340,N_2512);
nor U6574 (N_6574,N_2650,N_3805);
or U6575 (N_6575,N_4392,N_2544);
or U6576 (N_6576,N_2936,N_3895);
or U6577 (N_6577,N_3548,N_3126);
or U6578 (N_6578,N_2696,N_3169);
nor U6579 (N_6579,N_2982,N_3387);
nor U6580 (N_6580,N_4654,N_4663);
or U6581 (N_6581,N_4166,N_3050);
nor U6582 (N_6582,N_4591,N_3829);
or U6583 (N_6583,N_4802,N_4949);
and U6584 (N_6584,N_3578,N_4677);
xor U6585 (N_6585,N_4379,N_3308);
nor U6586 (N_6586,N_4536,N_3699);
and U6587 (N_6587,N_4895,N_3971);
or U6588 (N_6588,N_4479,N_3299);
or U6589 (N_6589,N_3234,N_3406);
xor U6590 (N_6590,N_4062,N_4367);
xor U6591 (N_6591,N_4872,N_4800);
nand U6592 (N_6592,N_3497,N_2519);
nand U6593 (N_6593,N_3674,N_3673);
and U6594 (N_6594,N_4173,N_4415);
xor U6595 (N_6595,N_4813,N_3971);
nand U6596 (N_6596,N_3062,N_3628);
xnor U6597 (N_6597,N_4937,N_3215);
nand U6598 (N_6598,N_2582,N_3688);
or U6599 (N_6599,N_4434,N_4571);
nor U6600 (N_6600,N_4326,N_3816);
nor U6601 (N_6601,N_3829,N_3909);
xnor U6602 (N_6602,N_2796,N_3924);
and U6603 (N_6603,N_3326,N_4470);
and U6604 (N_6604,N_4106,N_4393);
xor U6605 (N_6605,N_4861,N_3413);
nor U6606 (N_6606,N_3931,N_3616);
and U6607 (N_6607,N_4469,N_3114);
nand U6608 (N_6608,N_2681,N_4994);
nor U6609 (N_6609,N_3822,N_4620);
xnor U6610 (N_6610,N_2645,N_3451);
nor U6611 (N_6611,N_2571,N_3957);
xor U6612 (N_6612,N_4957,N_4044);
xor U6613 (N_6613,N_3840,N_2636);
nor U6614 (N_6614,N_2948,N_3835);
nor U6615 (N_6615,N_2521,N_4894);
nor U6616 (N_6616,N_3555,N_4849);
nor U6617 (N_6617,N_3039,N_4342);
and U6618 (N_6618,N_3696,N_3378);
and U6619 (N_6619,N_3702,N_4108);
nand U6620 (N_6620,N_3936,N_4755);
nand U6621 (N_6621,N_3191,N_4658);
xnor U6622 (N_6622,N_3880,N_2884);
nor U6623 (N_6623,N_3941,N_4639);
and U6624 (N_6624,N_3225,N_4890);
nand U6625 (N_6625,N_3517,N_3316);
xor U6626 (N_6626,N_3676,N_4954);
xor U6627 (N_6627,N_2746,N_4124);
and U6628 (N_6628,N_4645,N_4454);
xor U6629 (N_6629,N_4067,N_3621);
nand U6630 (N_6630,N_4523,N_3987);
xor U6631 (N_6631,N_3532,N_2545);
and U6632 (N_6632,N_2656,N_3778);
nor U6633 (N_6633,N_3360,N_2822);
and U6634 (N_6634,N_4006,N_2822);
nor U6635 (N_6635,N_3449,N_4057);
nand U6636 (N_6636,N_4933,N_4503);
nor U6637 (N_6637,N_4430,N_3587);
nand U6638 (N_6638,N_2740,N_4066);
xor U6639 (N_6639,N_4626,N_4467);
nand U6640 (N_6640,N_2905,N_3653);
nand U6641 (N_6641,N_4154,N_4003);
nor U6642 (N_6642,N_2639,N_4786);
nor U6643 (N_6643,N_3634,N_2606);
nor U6644 (N_6644,N_2944,N_2799);
nand U6645 (N_6645,N_3836,N_4166);
nor U6646 (N_6646,N_3986,N_2775);
nor U6647 (N_6647,N_3042,N_4453);
and U6648 (N_6648,N_4945,N_3341);
nor U6649 (N_6649,N_4196,N_3834);
nor U6650 (N_6650,N_4063,N_4268);
xnor U6651 (N_6651,N_3474,N_4187);
or U6652 (N_6652,N_4011,N_3993);
nor U6653 (N_6653,N_2919,N_4262);
nand U6654 (N_6654,N_4614,N_2581);
xnor U6655 (N_6655,N_3031,N_3374);
or U6656 (N_6656,N_4740,N_3363);
or U6657 (N_6657,N_4266,N_3783);
nand U6658 (N_6658,N_4932,N_2971);
xnor U6659 (N_6659,N_3840,N_2870);
nand U6660 (N_6660,N_3298,N_2640);
or U6661 (N_6661,N_2780,N_2572);
nor U6662 (N_6662,N_3224,N_2752);
or U6663 (N_6663,N_4846,N_4956);
xnor U6664 (N_6664,N_2739,N_2559);
and U6665 (N_6665,N_2717,N_3334);
xnor U6666 (N_6666,N_3223,N_4668);
or U6667 (N_6667,N_3204,N_4622);
nor U6668 (N_6668,N_3979,N_3427);
or U6669 (N_6669,N_3799,N_4975);
nor U6670 (N_6670,N_4484,N_4574);
and U6671 (N_6671,N_4730,N_4158);
or U6672 (N_6672,N_2670,N_2553);
xnor U6673 (N_6673,N_3737,N_4321);
or U6674 (N_6674,N_3681,N_3309);
nand U6675 (N_6675,N_4689,N_4042);
and U6676 (N_6676,N_3867,N_2778);
xor U6677 (N_6677,N_4925,N_3615);
xor U6678 (N_6678,N_4903,N_3895);
nand U6679 (N_6679,N_4504,N_3856);
nand U6680 (N_6680,N_4664,N_4854);
or U6681 (N_6681,N_4211,N_4814);
and U6682 (N_6682,N_2718,N_2824);
and U6683 (N_6683,N_4854,N_4400);
nand U6684 (N_6684,N_4658,N_4500);
or U6685 (N_6685,N_2548,N_4057);
or U6686 (N_6686,N_4859,N_4643);
or U6687 (N_6687,N_4113,N_4601);
xnor U6688 (N_6688,N_4674,N_3359);
nand U6689 (N_6689,N_2880,N_4672);
nand U6690 (N_6690,N_4831,N_4150);
nand U6691 (N_6691,N_2856,N_3566);
or U6692 (N_6692,N_3036,N_3424);
or U6693 (N_6693,N_2751,N_2985);
xor U6694 (N_6694,N_4236,N_2743);
nor U6695 (N_6695,N_4194,N_2681);
nand U6696 (N_6696,N_4184,N_3355);
nand U6697 (N_6697,N_3741,N_4402);
and U6698 (N_6698,N_4084,N_4010);
nand U6699 (N_6699,N_3556,N_4583);
xor U6700 (N_6700,N_3067,N_3713);
and U6701 (N_6701,N_3082,N_4930);
xnor U6702 (N_6702,N_3021,N_2949);
and U6703 (N_6703,N_2872,N_3100);
and U6704 (N_6704,N_4690,N_3472);
nand U6705 (N_6705,N_4446,N_3458);
nor U6706 (N_6706,N_2568,N_4912);
xnor U6707 (N_6707,N_3863,N_3067);
or U6708 (N_6708,N_3453,N_3993);
and U6709 (N_6709,N_2546,N_4730);
or U6710 (N_6710,N_3321,N_2879);
nand U6711 (N_6711,N_4206,N_2938);
and U6712 (N_6712,N_4683,N_2780);
xnor U6713 (N_6713,N_4300,N_3473);
nand U6714 (N_6714,N_3820,N_3701);
or U6715 (N_6715,N_2833,N_4870);
nand U6716 (N_6716,N_4073,N_4597);
nand U6717 (N_6717,N_3520,N_4780);
nand U6718 (N_6718,N_3383,N_4316);
and U6719 (N_6719,N_2580,N_2735);
or U6720 (N_6720,N_3242,N_4356);
xnor U6721 (N_6721,N_3213,N_4340);
nor U6722 (N_6722,N_3171,N_2843);
and U6723 (N_6723,N_3201,N_3110);
or U6724 (N_6724,N_4051,N_2726);
and U6725 (N_6725,N_2722,N_2646);
or U6726 (N_6726,N_3560,N_4335);
nand U6727 (N_6727,N_3900,N_4599);
xor U6728 (N_6728,N_3606,N_2998);
or U6729 (N_6729,N_3862,N_4238);
nor U6730 (N_6730,N_2545,N_4762);
nand U6731 (N_6731,N_3796,N_2712);
xor U6732 (N_6732,N_3523,N_4388);
nor U6733 (N_6733,N_4704,N_4497);
nor U6734 (N_6734,N_4326,N_4957);
xor U6735 (N_6735,N_3802,N_3325);
nand U6736 (N_6736,N_4103,N_4137);
nor U6737 (N_6737,N_3663,N_2888);
or U6738 (N_6738,N_4018,N_3901);
xnor U6739 (N_6739,N_4222,N_4776);
or U6740 (N_6740,N_2994,N_4333);
or U6741 (N_6741,N_4466,N_4851);
and U6742 (N_6742,N_4188,N_4879);
nand U6743 (N_6743,N_3455,N_2550);
xnor U6744 (N_6744,N_3079,N_2897);
or U6745 (N_6745,N_4758,N_2646);
nor U6746 (N_6746,N_2603,N_4577);
or U6747 (N_6747,N_2827,N_4986);
nor U6748 (N_6748,N_2807,N_4999);
or U6749 (N_6749,N_2784,N_3427);
nand U6750 (N_6750,N_3029,N_2821);
and U6751 (N_6751,N_3526,N_3594);
xor U6752 (N_6752,N_4497,N_4686);
and U6753 (N_6753,N_4206,N_4118);
or U6754 (N_6754,N_4747,N_3679);
xnor U6755 (N_6755,N_3827,N_3735);
nor U6756 (N_6756,N_2555,N_3022);
and U6757 (N_6757,N_3682,N_2977);
nor U6758 (N_6758,N_3645,N_4173);
nor U6759 (N_6759,N_4944,N_2647);
nor U6760 (N_6760,N_4416,N_3951);
nor U6761 (N_6761,N_3628,N_3612);
or U6762 (N_6762,N_3970,N_4831);
xor U6763 (N_6763,N_2952,N_3744);
nand U6764 (N_6764,N_3600,N_3248);
or U6765 (N_6765,N_2812,N_3538);
nand U6766 (N_6766,N_4107,N_4162);
nand U6767 (N_6767,N_4224,N_4461);
or U6768 (N_6768,N_4243,N_3830);
xor U6769 (N_6769,N_4439,N_4571);
xor U6770 (N_6770,N_4830,N_4861);
nand U6771 (N_6771,N_2988,N_2704);
or U6772 (N_6772,N_3613,N_3644);
or U6773 (N_6773,N_4786,N_3126);
or U6774 (N_6774,N_3358,N_4280);
and U6775 (N_6775,N_4180,N_3067);
or U6776 (N_6776,N_4316,N_3121);
xnor U6777 (N_6777,N_4005,N_4367);
or U6778 (N_6778,N_4548,N_3989);
nand U6779 (N_6779,N_3366,N_4348);
or U6780 (N_6780,N_3843,N_2885);
nor U6781 (N_6781,N_3982,N_2615);
nand U6782 (N_6782,N_2622,N_4452);
nand U6783 (N_6783,N_3185,N_3790);
nor U6784 (N_6784,N_3109,N_3037);
xor U6785 (N_6785,N_3690,N_4035);
nand U6786 (N_6786,N_2709,N_3518);
xnor U6787 (N_6787,N_4173,N_3079);
or U6788 (N_6788,N_3820,N_2506);
or U6789 (N_6789,N_3364,N_3891);
xnor U6790 (N_6790,N_4168,N_3173);
xnor U6791 (N_6791,N_4901,N_3818);
and U6792 (N_6792,N_3073,N_2656);
xor U6793 (N_6793,N_3894,N_2538);
or U6794 (N_6794,N_4790,N_3691);
xor U6795 (N_6795,N_3700,N_4268);
xnor U6796 (N_6796,N_3841,N_2650);
and U6797 (N_6797,N_4509,N_4150);
nand U6798 (N_6798,N_2801,N_4578);
xnor U6799 (N_6799,N_3643,N_4309);
nand U6800 (N_6800,N_4309,N_4072);
nand U6801 (N_6801,N_3829,N_3337);
and U6802 (N_6802,N_4611,N_3453);
xor U6803 (N_6803,N_3319,N_4707);
or U6804 (N_6804,N_2554,N_4108);
nand U6805 (N_6805,N_3376,N_4486);
xnor U6806 (N_6806,N_2640,N_4449);
xor U6807 (N_6807,N_4396,N_3012);
nand U6808 (N_6808,N_3431,N_4897);
nand U6809 (N_6809,N_4346,N_3229);
and U6810 (N_6810,N_3272,N_2928);
nand U6811 (N_6811,N_4039,N_4953);
xnor U6812 (N_6812,N_3172,N_4162);
or U6813 (N_6813,N_4158,N_4328);
xor U6814 (N_6814,N_4640,N_4751);
nand U6815 (N_6815,N_4738,N_4997);
nand U6816 (N_6816,N_4769,N_4879);
xor U6817 (N_6817,N_3462,N_4827);
xor U6818 (N_6818,N_4047,N_4095);
and U6819 (N_6819,N_3695,N_4651);
nor U6820 (N_6820,N_4295,N_4431);
and U6821 (N_6821,N_4658,N_2979);
nand U6822 (N_6822,N_4525,N_4565);
and U6823 (N_6823,N_3839,N_2960);
or U6824 (N_6824,N_2629,N_3494);
xnor U6825 (N_6825,N_2754,N_2641);
or U6826 (N_6826,N_2961,N_3569);
and U6827 (N_6827,N_3933,N_3000);
nand U6828 (N_6828,N_3222,N_3121);
or U6829 (N_6829,N_3442,N_3459);
nor U6830 (N_6830,N_3806,N_4171);
or U6831 (N_6831,N_4770,N_4527);
or U6832 (N_6832,N_3735,N_3879);
nor U6833 (N_6833,N_3543,N_3316);
and U6834 (N_6834,N_3029,N_2586);
or U6835 (N_6835,N_3896,N_4717);
xor U6836 (N_6836,N_2508,N_3711);
nor U6837 (N_6837,N_3767,N_4380);
nor U6838 (N_6838,N_3540,N_3478);
nand U6839 (N_6839,N_2557,N_4824);
nand U6840 (N_6840,N_4219,N_2859);
or U6841 (N_6841,N_3179,N_3719);
and U6842 (N_6842,N_3664,N_3521);
or U6843 (N_6843,N_2569,N_4834);
nor U6844 (N_6844,N_3966,N_2729);
and U6845 (N_6845,N_3235,N_2594);
xor U6846 (N_6846,N_3009,N_3875);
nand U6847 (N_6847,N_3945,N_4348);
xnor U6848 (N_6848,N_3498,N_3109);
or U6849 (N_6849,N_4311,N_4237);
nand U6850 (N_6850,N_3641,N_3642);
xnor U6851 (N_6851,N_4611,N_3122);
xnor U6852 (N_6852,N_2583,N_3225);
or U6853 (N_6853,N_4026,N_2600);
or U6854 (N_6854,N_4424,N_4384);
nor U6855 (N_6855,N_3347,N_3874);
and U6856 (N_6856,N_2991,N_3634);
nand U6857 (N_6857,N_2703,N_4668);
and U6858 (N_6858,N_2855,N_3721);
xor U6859 (N_6859,N_2835,N_4599);
or U6860 (N_6860,N_4351,N_3119);
nor U6861 (N_6861,N_2541,N_3668);
nor U6862 (N_6862,N_4574,N_2651);
and U6863 (N_6863,N_4706,N_3143);
xnor U6864 (N_6864,N_3706,N_3866);
and U6865 (N_6865,N_3645,N_2916);
xnor U6866 (N_6866,N_3622,N_3359);
nand U6867 (N_6867,N_3494,N_2968);
and U6868 (N_6868,N_4212,N_4158);
and U6869 (N_6869,N_3892,N_3947);
nor U6870 (N_6870,N_2798,N_4025);
xnor U6871 (N_6871,N_3565,N_3407);
nand U6872 (N_6872,N_2741,N_4392);
or U6873 (N_6873,N_3462,N_4527);
nor U6874 (N_6874,N_4211,N_3470);
xnor U6875 (N_6875,N_4234,N_4613);
or U6876 (N_6876,N_2789,N_4480);
nand U6877 (N_6877,N_4246,N_2508);
nor U6878 (N_6878,N_4797,N_4687);
nor U6879 (N_6879,N_4941,N_2693);
or U6880 (N_6880,N_3332,N_3775);
nor U6881 (N_6881,N_3519,N_4067);
or U6882 (N_6882,N_3629,N_3563);
or U6883 (N_6883,N_3571,N_3844);
nand U6884 (N_6884,N_4774,N_3166);
and U6885 (N_6885,N_2875,N_4375);
nand U6886 (N_6886,N_4408,N_3718);
xnor U6887 (N_6887,N_4697,N_4326);
nand U6888 (N_6888,N_3752,N_3488);
xor U6889 (N_6889,N_3742,N_4680);
or U6890 (N_6890,N_3911,N_3841);
and U6891 (N_6891,N_2606,N_4380);
nor U6892 (N_6892,N_4798,N_4310);
nand U6893 (N_6893,N_3013,N_3988);
nand U6894 (N_6894,N_4755,N_4777);
nor U6895 (N_6895,N_4601,N_2894);
and U6896 (N_6896,N_4162,N_3459);
nand U6897 (N_6897,N_3182,N_4410);
nor U6898 (N_6898,N_4868,N_2850);
xnor U6899 (N_6899,N_2944,N_4733);
or U6900 (N_6900,N_4375,N_3516);
xor U6901 (N_6901,N_3804,N_2589);
xnor U6902 (N_6902,N_2887,N_4092);
or U6903 (N_6903,N_4625,N_4367);
nand U6904 (N_6904,N_4727,N_4903);
xor U6905 (N_6905,N_4471,N_2573);
nor U6906 (N_6906,N_3382,N_2918);
and U6907 (N_6907,N_2835,N_4528);
nor U6908 (N_6908,N_4120,N_3447);
nand U6909 (N_6909,N_2712,N_3622);
nor U6910 (N_6910,N_3221,N_3493);
nor U6911 (N_6911,N_3457,N_4068);
or U6912 (N_6912,N_2721,N_3642);
nand U6913 (N_6913,N_3494,N_4359);
and U6914 (N_6914,N_4225,N_4412);
nand U6915 (N_6915,N_3492,N_3473);
nor U6916 (N_6916,N_3938,N_3876);
or U6917 (N_6917,N_2892,N_4538);
or U6918 (N_6918,N_4582,N_2851);
or U6919 (N_6919,N_2553,N_4122);
xor U6920 (N_6920,N_3757,N_3789);
nand U6921 (N_6921,N_2773,N_3057);
nand U6922 (N_6922,N_3726,N_2991);
or U6923 (N_6923,N_2656,N_4321);
and U6924 (N_6924,N_4860,N_3622);
or U6925 (N_6925,N_4738,N_3679);
or U6926 (N_6926,N_3637,N_4454);
nand U6927 (N_6927,N_3788,N_4316);
or U6928 (N_6928,N_2945,N_3221);
nand U6929 (N_6929,N_4009,N_4963);
or U6930 (N_6930,N_2897,N_4565);
nand U6931 (N_6931,N_2623,N_4320);
xor U6932 (N_6932,N_2886,N_3412);
nand U6933 (N_6933,N_4470,N_3872);
and U6934 (N_6934,N_2720,N_4738);
nand U6935 (N_6935,N_2995,N_4868);
xor U6936 (N_6936,N_3610,N_3611);
nand U6937 (N_6937,N_4034,N_3727);
or U6938 (N_6938,N_2605,N_3743);
nor U6939 (N_6939,N_4845,N_2688);
nand U6940 (N_6940,N_3290,N_4218);
xnor U6941 (N_6941,N_4976,N_4288);
nand U6942 (N_6942,N_2697,N_4991);
nand U6943 (N_6943,N_4430,N_4869);
nand U6944 (N_6944,N_2574,N_3761);
xor U6945 (N_6945,N_3870,N_4339);
or U6946 (N_6946,N_2763,N_2545);
nand U6947 (N_6947,N_4127,N_4831);
and U6948 (N_6948,N_4589,N_2845);
nand U6949 (N_6949,N_3508,N_3739);
nand U6950 (N_6950,N_4828,N_4069);
nand U6951 (N_6951,N_3264,N_2658);
or U6952 (N_6952,N_4662,N_3474);
or U6953 (N_6953,N_2662,N_4324);
nor U6954 (N_6954,N_4402,N_3682);
nand U6955 (N_6955,N_4303,N_3644);
xor U6956 (N_6956,N_4883,N_3665);
or U6957 (N_6957,N_2876,N_4032);
nor U6958 (N_6958,N_3828,N_2927);
nor U6959 (N_6959,N_4928,N_4816);
xnor U6960 (N_6960,N_3070,N_3121);
and U6961 (N_6961,N_3050,N_2609);
and U6962 (N_6962,N_3267,N_3839);
nand U6963 (N_6963,N_4185,N_3121);
nor U6964 (N_6964,N_3632,N_2616);
and U6965 (N_6965,N_3819,N_3837);
and U6966 (N_6966,N_4445,N_4376);
nand U6967 (N_6967,N_4589,N_3806);
nand U6968 (N_6968,N_4688,N_3915);
nand U6969 (N_6969,N_2885,N_4418);
and U6970 (N_6970,N_2970,N_4669);
and U6971 (N_6971,N_2729,N_2806);
and U6972 (N_6972,N_4652,N_2964);
nand U6973 (N_6973,N_3568,N_2652);
nor U6974 (N_6974,N_2707,N_2996);
xor U6975 (N_6975,N_2816,N_2985);
and U6976 (N_6976,N_3225,N_3947);
nand U6977 (N_6977,N_2539,N_3017);
and U6978 (N_6978,N_2706,N_3089);
or U6979 (N_6979,N_3643,N_4981);
xor U6980 (N_6980,N_4294,N_4780);
and U6981 (N_6981,N_4101,N_4021);
or U6982 (N_6982,N_2767,N_2909);
nor U6983 (N_6983,N_4598,N_4555);
or U6984 (N_6984,N_3254,N_4154);
and U6985 (N_6985,N_2523,N_4714);
nor U6986 (N_6986,N_3071,N_4144);
nand U6987 (N_6987,N_3302,N_3877);
xor U6988 (N_6988,N_4009,N_4388);
and U6989 (N_6989,N_2586,N_3009);
nor U6990 (N_6990,N_3917,N_3857);
nand U6991 (N_6991,N_4645,N_3728);
or U6992 (N_6992,N_4258,N_3681);
xor U6993 (N_6993,N_4472,N_3193);
nand U6994 (N_6994,N_3626,N_3180);
nor U6995 (N_6995,N_2561,N_4706);
nand U6996 (N_6996,N_3998,N_4706);
or U6997 (N_6997,N_2886,N_4843);
nor U6998 (N_6998,N_3137,N_4440);
nand U6999 (N_6999,N_3868,N_4255);
nor U7000 (N_7000,N_3774,N_3518);
nand U7001 (N_7001,N_2880,N_4933);
or U7002 (N_7002,N_3131,N_4481);
or U7003 (N_7003,N_3389,N_3088);
and U7004 (N_7004,N_4748,N_2777);
nor U7005 (N_7005,N_3524,N_3489);
and U7006 (N_7006,N_4806,N_3510);
nor U7007 (N_7007,N_4747,N_4755);
nor U7008 (N_7008,N_2623,N_3596);
or U7009 (N_7009,N_2835,N_3276);
or U7010 (N_7010,N_3475,N_4936);
or U7011 (N_7011,N_4418,N_3042);
nor U7012 (N_7012,N_4678,N_3120);
or U7013 (N_7013,N_4811,N_3619);
nand U7014 (N_7014,N_4070,N_2925);
or U7015 (N_7015,N_3377,N_4686);
nand U7016 (N_7016,N_3071,N_4319);
nand U7017 (N_7017,N_2997,N_3887);
xnor U7018 (N_7018,N_4895,N_3807);
nand U7019 (N_7019,N_3919,N_3246);
xnor U7020 (N_7020,N_3439,N_4521);
and U7021 (N_7021,N_4992,N_3630);
nor U7022 (N_7022,N_3499,N_4239);
xor U7023 (N_7023,N_3811,N_3371);
and U7024 (N_7024,N_4427,N_4115);
and U7025 (N_7025,N_4959,N_3830);
nor U7026 (N_7026,N_3206,N_3480);
nand U7027 (N_7027,N_3901,N_2566);
or U7028 (N_7028,N_2834,N_3603);
nor U7029 (N_7029,N_3939,N_3835);
or U7030 (N_7030,N_4523,N_2612);
or U7031 (N_7031,N_4230,N_3010);
and U7032 (N_7032,N_4406,N_4793);
xor U7033 (N_7033,N_4488,N_3496);
and U7034 (N_7034,N_3150,N_3288);
xor U7035 (N_7035,N_3549,N_3541);
or U7036 (N_7036,N_3924,N_3459);
and U7037 (N_7037,N_3043,N_3058);
nor U7038 (N_7038,N_4663,N_4028);
and U7039 (N_7039,N_3162,N_4133);
and U7040 (N_7040,N_3723,N_4386);
nand U7041 (N_7041,N_4172,N_2564);
nand U7042 (N_7042,N_2953,N_4370);
nor U7043 (N_7043,N_4688,N_4950);
nand U7044 (N_7044,N_4915,N_3997);
xor U7045 (N_7045,N_3274,N_3525);
or U7046 (N_7046,N_4268,N_3510);
xnor U7047 (N_7047,N_2929,N_4998);
and U7048 (N_7048,N_2935,N_4115);
nor U7049 (N_7049,N_3970,N_3636);
nand U7050 (N_7050,N_4749,N_2660);
xor U7051 (N_7051,N_3601,N_2969);
or U7052 (N_7052,N_4232,N_3001);
and U7053 (N_7053,N_3266,N_2668);
xor U7054 (N_7054,N_4999,N_4797);
nand U7055 (N_7055,N_3156,N_3033);
xor U7056 (N_7056,N_2573,N_4631);
nand U7057 (N_7057,N_2773,N_3031);
nand U7058 (N_7058,N_4717,N_3319);
or U7059 (N_7059,N_2774,N_2865);
and U7060 (N_7060,N_2536,N_3206);
nand U7061 (N_7061,N_2599,N_4174);
or U7062 (N_7062,N_2578,N_4079);
and U7063 (N_7063,N_3142,N_2766);
nand U7064 (N_7064,N_4792,N_4643);
and U7065 (N_7065,N_4294,N_4916);
nand U7066 (N_7066,N_4376,N_3233);
xor U7067 (N_7067,N_4854,N_2672);
xnor U7068 (N_7068,N_3229,N_2919);
xnor U7069 (N_7069,N_3830,N_2968);
xnor U7070 (N_7070,N_3503,N_4407);
xnor U7071 (N_7071,N_2540,N_4874);
nand U7072 (N_7072,N_3133,N_3690);
or U7073 (N_7073,N_4338,N_4008);
nor U7074 (N_7074,N_2912,N_4830);
nand U7075 (N_7075,N_4639,N_2926);
xnor U7076 (N_7076,N_3861,N_3411);
or U7077 (N_7077,N_4947,N_3093);
xor U7078 (N_7078,N_2816,N_2774);
and U7079 (N_7079,N_4913,N_2630);
and U7080 (N_7080,N_3663,N_2974);
nand U7081 (N_7081,N_2882,N_3127);
or U7082 (N_7082,N_3786,N_4558);
nand U7083 (N_7083,N_3280,N_2588);
xnor U7084 (N_7084,N_3473,N_2767);
nand U7085 (N_7085,N_4293,N_3741);
xor U7086 (N_7086,N_2762,N_3005);
nand U7087 (N_7087,N_3554,N_4306);
nor U7088 (N_7088,N_3162,N_2907);
or U7089 (N_7089,N_2666,N_3655);
or U7090 (N_7090,N_4778,N_3580);
nand U7091 (N_7091,N_2929,N_4636);
nand U7092 (N_7092,N_4859,N_4116);
and U7093 (N_7093,N_4605,N_3341);
or U7094 (N_7094,N_2957,N_2937);
nor U7095 (N_7095,N_2997,N_4275);
and U7096 (N_7096,N_4786,N_3078);
and U7097 (N_7097,N_3944,N_3374);
or U7098 (N_7098,N_3593,N_4487);
and U7099 (N_7099,N_3432,N_4849);
xor U7100 (N_7100,N_2937,N_4276);
xor U7101 (N_7101,N_2972,N_4865);
nor U7102 (N_7102,N_2836,N_4809);
or U7103 (N_7103,N_3502,N_4500);
or U7104 (N_7104,N_4862,N_3021);
and U7105 (N_7105,N_2756,N_4083);
nand U7106 (N_7106,N_4011,N_3043);
and U7107 (N_7107,N_3786,N_4796);
and U7108 (N_7108,N_4436,N_3320);
or U7109 (N_7109,N_3733,N_4608);
nand U7110 (N_7110,N_2564,N_3377);
and U7111 (N_7111,N_3419,N_2541);
nand U7112 (N_7112,N_4395,N_4831);
and U7113 (N_7113,N_4119,N_3303);
nor U7114 (N_7114,N_2855,N_3722);
xor U7115 (N_7115,N_3059,N_4737);
nor U7116 (N_7116,N_4169,N_3436);
xor U7117 (N_7117,N_4381,N_3725);
xor U7118 (N_7118,N_4777,N_3993);
nand U7119 (N_7119,N_3429,N_3115);
or U7120 (N_7120,N_3342,N_2801);
nand U7121 (N_7121,N_4297,N_2900);
and U7122 (N_7122,N_3912,N_4691);
and U7123 (N_7123,N_2931,N_3899);
or U7124 (N_7124,N_3235,N_4261);
and U7125 (N_7125,N_3052,N_4290);
nor U7126 (N_7126,N_2806,N_4067);
and U7127 (N_7127,N_3294,N_3983);
and U7128 (N_7128,N_3391,N_4597);
xnor U7129 (N_7129,N_2529,N_4820);
xor U7130 (N_7130,N_4753,N_2560);
xor U7131 (N_7131,N_2951,N_2542);
or U7132 (N_7132,N_3304,N_2688);
nor U7133 (N_7133,N_2889,N_4334);
or U7134 (N_7134,N_3349,N_3397);
nor U7135 (N_7135,N_2738,N_3678);
and U7136 (N_7136,N_2886,N_3207);
and U7137 (N_7137,N_2891,N_2663);
or U7138 (N_7138,N_4894,N_2771);
xor U7139 (N_7139,N_4028,N_4823);
nand U7140 (N_7140,N_3596,N_4389);
nor U7141 (N_7141,N_3349,N_3901);
and U7142 (N_7142,N_4091,N_3242);
xor U7143 (N_7143,N_2506,N_4993);
and U7144 (N_7144,N_2902,N_3428);
nor U7145 (N_7145,N_3286,N_3412);
nor U7146 (N_7146,N_2699,N_4434);
xnor U7147 (N_7147,N_3098,N_4831);
nor U7148 (N_7148,N_2874,N_3405);
nor U7149 (N_7149,N_3289,N_3209);
and U7150 (N_7150,N_3096,N_4183);
and U7151 (N_7151,N_2627,N_4715);
or U7152 (N_7152,N_2737,N_3355);
and U7153 (N_7153,N_3433,N_4812);
xnor U7154 (N_7154,N_3134,N_3362);
and U7155 (N_7155,N_4737,N_3022);
xnor U7156 (N_7156,N_4288,N_4060);
and U7157 (N_7157,N_3128,N_3531);
nor U7158 (N_7158,N_3781,N_2617);
nor U7159 (N_7159,N_4431,N_3860);
nor U7160 (N_7160,N_4066,N_2844);
nor U7161 (N_7161,N_4438,N_4101);
xor U7162 (N_7162,N_2824,N_2743);
and U7163 (N_7163,N_2873,N_4524);
xnor U7164 (N_7164,N_3193,N_4165);
and U7165 (N_7165,N_3418,N_2950);
nand U7166 (N_7166,N_3251,N_4816);
nor U7167 (N_7167,N_3031,N_4024);
and U7168 (N_7168,N_4427,N_3569);
nand U7169 (N_7169,N_4703,N_3246);
xor U7170 (N_7170,N_3901,N_3126);
nor U7171 (N_7171,N_3189,N_4819);
or U7172 (N_7172,N_3441,N_4614);
and U7173 (N_7173,N_4710,N_4400);
xnor U7174 (N_7174,N_2998,N_4912);
and U7175 (N_7175,N_3904,N_4677);
or U7176 (N_7176,N_3943,N_4590);
and U7177 (N_7177,N_2612,N_3179);
nor U7178 (N_7178,N_3878,N_4712);
nand U7179 (N_7179,N_4148,N_4361);
xnor U7180 (N_7180,N_2753,N_4471);
xor U7181 (N_7181,N_4658,N_3736);
nor U7182 (N_7182,N_4102,N_3525);
or U7183 (N_7183,N_4623,N_3002);
nand U7184 (N_7184,N_4705,N_3525);
and U7185 (N_7185,N_2746,N_4539);
nor U7186 (N_7186,N_2840,N_4393);
nor U7187 (N_7187,N_3692,N_4005);
or U7188 (N_7188,N_4325,N_4224);
or U7189 (N_7189,N_4998,N_3752);
and U7190 (N_7190,N_4586,N_2769);
xor U7191 (N_7191,N_3112,N_4242);
nor U7192 (N_7192,N_3161,N_2899);
nand U7193 (N_7193,N_4028,N_3345);
nand U7194 (N_7194,N_2844,N_3886);
and U7195 (N_7195,N_4731,N_3230);
nand U7196 (N_7196,N_3557,N_4809);
or U7197 (N_7197,N_2607,N_4013);
or U7198 (N_7198,N_4568,N_2752);
xnor U7199 (N_7199,N_3123,N_3602);
xnor U7200 (N_7200,N_3532,N_4484);
nor U7201 (N_7201,N_2547,N_4150);
or U7202 (N_7202,N_2810,N_2769);
nand U7203 (N_7203,N_3794,N_2544);
and U7204 (N_7204,N_3529,N_4573);
and U7205 (N_7205,N_3716,N_3803);
and U7206 (N_7206,N_4206,N_4887);
and U7207 (N_7207,N_3874,N_3940);
nor U7208 (N_7208,N_2513,N_2626);
nand U7209 (N_7209,N_4321,N_3785);
nand U7210 (N_7210,N_3319,N_3538);
or U7211 (N_7211,N_4025,N_3069);
xor U7212 (N_7212,N_3170,N_4873);
and U7213 (N_7213,N_4190,N_3428);
or U7214 (N_7214,N_2764,N_2557);
nor U7215 (N_7215,N_4955,N_4037);
or U7216 (N_7216,N_3370,N_4215);
nand U7217 (N_7217,N_4553,N_4181);
nand U7218 (N_7218,N_3447,N_4823);
or U7219 (N_7219,N_4984,N_3911);
nor U7220 (N_7220,N_4447,N_4296);
nor U7221 (N_7221,N_2671,N_3184);
nand U7222 (N_7222,N_4905,N_4522);
nand U7223 (N_7223,N_3317,N_3659);
nand U7224 (N_7224,N_3782,N_4350);
xnor U7225 (N_7225,N_3217,N_4690);
and U7226 (N_7226,N_3067,N_3785);
xor U7227 (N_7227,N_3720,N_2656);
xnor U7228 (N_7228,N_2833,N_2757);
or U7229 (N_7229,N_3423,N_4554);
nor U7230 (N_7230,N_2645,N_4968);
xor U7231 (N_7231,N_4488,N_2934);
or U7232 (N_7232,N_4240,N_3879);
and U7233 (N_7233,N_4892,N_4821);
nor U7234 (N_7234,N_3237,N_3659);
nor U7235 (N_7235,N_2565,N_3548);
or U7236 (N_7236,N_3687,N_3975);
nor U7237 (N_7237,N_4728,N_3882);
or U7238 (N_7238,N_4908,N_3005);
and U7239 (N_7239,N_4405,N_4900);
or U7240 (N_7240,N_3922,N_2550);
xor U7241 (N_7241,N_4358,N_4994);
nand U7242 (N_7242,N_3451,N_4586);
or U7243 (N_7243,N_4232,N_2777);
and U7244 (N_7244,N_4577,N_3265);
nor U7245 (N_7245,N_3754,N_2795);
xor U7246 (N_7246,N_3753,N_3486);
xor U7247 (N_7247,N_2509,N_4852);
or U7248 (N_7248,N_4887,N_3064);
nand U7249 (N_7249,N_4103,N_3671);
or U7250 (N_7250,N_2932,N_4052);
and U7251 (N_7251,N_2667,N_3014);
and U7252 (N_7252,N_2772,N_3010);
or U7253 (N_7253,N_2816,N_3512);
or U7254 (N_7254,N_2657,N_4856);
and U7255 (N_7255,N_2501,N_2506);
and U7256 (N_7256,N_2887,N_2678);
or U7257 (N_7257,N_4274,N_4433);
nand U7258 (N_7258,N_3654,N_4160);
nand U7259 (N_7259,N_2679,N_2934);
nand U7260 (N_7260,N_4704,N_4238);
nor U7261 (N_7261,N_3716,N_4750);
nor U7262 (N_7262,N_2660,N_3525);
nand U7263 (N_7263,N_3984,N_4692);
and U7264 (N_7264,N_4589,N_2511);
xor U7265 (N_7265,N_2989,N_4516);
xnor U7266 (N_7266,N_4067,N_4670);
xor U7267 (N_7267,N_3996,N_4910);
nand U7268 (N_7268,N_3128,N_4402);
nand U7269 (N_7269,N_4843,N_3680);
and U7270 (N_7270,N_2945,N_4013);
and U7271 (N_7271,N_2922,N_3775);
or U7272 (N_7272,N_4183,N_4792);
and U7273 (N_7273,N_4594,N_4852);
nand U7274 (N_7274,N_4725,N_4385);
nor U7275 (N_7275,N_4011,N_4755);
xnor U7276 (N_7276,N_3270,N_4803);
xor U7277 (N_7277,N_4442,N_2717);
nand U7278 (N_7278,N_3103,N_3344);
nand U7279 (N_7279,N_3559,N_2663);
nor U7280 (N_7280,N_4084,N_4162);
xor U7281 (N_7281,N_3138,N_3349);
xor U7282 (N_7282,N_4823,N_4484);
and U7283 (N_7283,N_3286,N_4425);
nand U7284 (N_7284,N_2516,N_2804);
nand U7285 (N_7285,N_4403,N_2768);
and U7286 (N_7286,N_3293,N_3104);
nand U7287 (N_7287,N_4673,N_3563);
and U7288 (N_7288,N_3189,N_4476);
or U7289 (N_7289,N_4797,N_4441);
and U7290 (N_7290,N_2803,N_3450);
or U7291 (N_7291,N_3149,N_3507);
nand U7292 (N_7292,N_4446,N_4512);
nand U7293 (N_7293,N_3578,N_3706);
nand U7294 (N_7294,N_3347,N_3570);
nand U7295 (N_7295,N_2544,N_2783);
xnor U7296 (N_7296,N_3818,N_2972);
and U7297 (N_7297,N_3124,N_2714);
nor U7298 (N_7298,N_3100,N_4793);
nor U7299 (N_7299,N_3376,N_4136);
or U7300 (N_7300,N_2601,N_4568);
and U7301 (N_7301,N_3748,N_3419);
xor U7302 (N_7302,N_3349,N_2790);
and U7303 (N_7303,N_4118,N_4707);
nand U7304 (N_7304,N_4461,N_3430);
nor U7305 (N_7305,N_4865,N_4357);
or U7306 (N_7306,N_3238,N_3104);
xnor U7307 (N_7307,N_3344,N_4968);
and U7308 (N_7308,N_4659,N_4487);
and U7309 (N_7309,N_4600,N_4160);
xnor U7310 (N_7310,N_4278,N_3198);
xor U7311 (N_7311,N_4499,N_2704);
xor U7312 (N_7312,N_4449,N_4393);
xor U7313 (N_7313,N_3138,N_3900);
xor U7314 (N_7314,N_4502,N_4368);
nand U7315 (N_7315,N_4133,N_3493);
nor U7316 (N_7316,N_4836,N_4600);
or U7317 (N_7317,N_3787,N_2721);
or U7318 (N_7318,N_4245,N_4455);
and U7319 (N_7319,N_4044,N_2975);
nand U7320 (N_7320,N_3960,N_3996);
nor U7321 (N_7321,N_3989,N_3720);
xor U7322 (N_7322,N_3514,N_2962);
or U7323 (N_7323,N_4427,N_4426);
nor U7324 (N_7324,N_3406,N_3460);
nand U7325 (N_7325,N_4743,N_4497);
nor U7326 (N_7326,N_4293,N_3727);
nor U7327 (N_7327,N_3282,N_2787);
nor U7328 (N_7328,N_4840,N_4841);
or U7329 (N_7329,N_3929,N_3315);
or U7330 (N_7330,N_3944,N_3340);
or U7331 (N_7331,N_4112,N_3091);
xor U7332 (N_7332,N_2959,N_3353);
xor U7333 (N_7333,N_3873,N_2932);
xnor U7334 (N_7334,N_4994,N_4524);
nor U7335 (N_7335,N_3082,N_2567);
nor U7336 (N_7336,N_4501,N_4002);
or U7337 (N_7337,N_3572,N_2895);
nand U7338 (N_7338,N_3250,N_4468);
or U7339 (N_7339,N_4688,N_4847);
or U7340 (N_7340,N_3156,N_4906);
xor U7341 (N_7341,N_2832,N_3218);
and U7342 (N_7342,N_4594,N_4876);
nand U7343 (N_7343,N_4490,N_2770);
xor U7344 (N_7344,N_2975,N_3994);
xnor U7345 (N_7345,N_3372,N_3926);
xnor U7346 (N_7346,N_3238,N_3048);
and U7347 (N_7347,N_2516,N_4706);
or U7348 (N_7348,N_2809,N_4918);
nand U7349 (N_7349,N_3051,N_2806);
and U7350 (N_7350,N_3789,N_4909);
nor U7351 (N_7351,N_3557,N_3421);
nand U7352 (N_7352,N_4933,N_2776);
and U7353 (N_7353,N_3429,N_4656);
or U7354 (N_7354,N_4609,N_2729);
nor U7355 (N_7355,N_2524,N_3921);
or U7356 (N_7356,N_3504,N_4363);
or U7357 (N_7357,N_4335,N_2730);
xnor U7358 (N_7358,N_4764,N_2767);
nand U7359 (N_7359,N_3988,N_4771);
xor U7360 (N_7360,N_3063,N_2503);
and U7361 (N_7361,N_3502,N_3082);
nor U7362 (N_7362,N_2553,N_4510);
nand U7363 (N_7363,N_2816,N_3570);
nor U7364 (N_7364,N_3267,N_3507);
nand U7365 (N_7365,N_2736,N_2959);
xnor U7366 (N_7366,N_3633,N_4028);
and U7367 (N_7367,N_2539,N_4660);
or U7368 (N_7368,N_3050,N_2928);
or U7369 (N_7369,N_2717,N_2514);
or U7370 (N_7370,N_4796,N_4098);
nor U7371 (N_7371,N_2579,N_4516);
or U7372 (N_7372,N_2953,N_3809);
and U7373 (N_7373,N_3918,N_2753);
or U7374 (N_7374,N_4954,N_4660);
xor U7375 (N_7375,N_2902,N_2758);
nor U7376 (N_7376,N_3741,N_3619);
and U7377 (N_7377,N_4789,N_3239);
or U7378 (N_7378,N_4057,N_3767);
or U7379 (N_7379,N_4649,N_2684);
nor U7380 (N_7380,N_4056,N_3010);
or U7381 (N_7381,N_2677,N_4462);
and U7382 (N_7382,N_3244,N_3262);
and U7383 (N_7383,N_2594,N_2642);
nand U7384 (N_7384,N_3383,N_3028);
xnor U7385 (N_7385,N_3987,N_3769);
and U7386 (N_7386,N_3497,N_3679);
nand U7387 (N_7387,N_3044,N_4871);
nor U7388 (N_7388,N_4917,N_3154);
and U7389 (N_7389,N_4086,N_3809);
xnor U7390 (N_7390,N_2974,N_3695);
nand U7391 (N_7391,N_4001,N_3230);
nor U7392 (N_7392,N_3106,N_3805);
nand U7393 (N_7393,N_4145,N_3364);
or U7394 (N_7394,N_2507,N_4108);
nand U7395 (N_7395,N_4527,N_3601);
xor U7396 (N_7396,N_2620,N_2549);
xor U7397 (N_7397,N_4129,N_4588);
nor U7398 (N_7398,N_4768,N_3871);
xor U7399 (N_7399,N_3666,N_4497);
xor U7400 (N_7400,N_4491,N_4733);
or U7401 (N_7401,N_3200,N_2832);
and U7402 (N_7402,N_4754,N_4904);
and U7403 (N_7403,N_4230,N_3234);
nand U7404 (N_7404,N_4596,N_4804);
and U7405 (N_7405,N_4771,N_2917);
nor U7406 (N_7406,N_4088,N_3580);
nand U7407 (N_7407,N_2750,N_4083);
xnor U7408 (N_7408,N_4751,N_4771);
nand U7409 (N_7409,N_4195,N_3030);
nor U7410 (N_7410,N_4677,N_4608);
xnor U7411 (N_7411,N_2769,N_3670);
nand U7412 (N_7412,N_4198,N_3346);
nand U7413 (N_7413,N_3027,N_4729);
nor U7414 (N_7414,N_3770,N_2890);
nand U7415 (N_7415,N_4968,N_4495);
nor U7416 (N_7416,N_3136,N_4932);
and U7417 (N_7417,N_3849,N_3969);
or U7418 (N_7418,N_4598,N_4518);
or U7419 (N_7419,N_2997,N_3979);
xor U7420 (N_7420,N_4648,N_3815);
or U7421 (N_7421,N_4508,N_3655);
and U7422 (N_7422,N_2870,N_3067);
and U7423 (N_7423,N_3982,N_2954);
nor U7424 (N_7424,N_3450,N_3008);
or U7425 (N_7425,N_2867,N_3081);
and U7426 (N_7426,N_3178,N_4356);
nor U7427 (N_7427,N_3606,N_3894);
nand U7428 (N_7428,N_3039,N_3528);
or U7429 (N_7429,N_4278,N_2536);
or U7430 (N_7430,N_3265,N_3512);
xor U7431 (N_7431,N_3594,N_4031);
nor U7432 (N_7432,N_3799,N_2505);
nand U7433 (N_7433,N_4206,N_3376);
nor U7434 (N_7434,N_3185,N_4403);
nand U7435 (N_7435,N_4406,N_2584);
xor U7436 (N_7436,N_3764,N_4309);
nand U7437 (N_7437,N_3334,N_3282);
and U7438 (N_7438,N_3720,N_3885);
or U7439 (N_7439,N_4178,N_2971);
xor U7440 (N_7440,N_3820,N_3699);
nor U7441 (N_7441,N_3619,N_3758);
nor U7442 (N_7442,N_4939,N_4669);
nor U7443 (N_7443,N_3268,N_2865);
nand U7444 (N_7444,N_4187,N_2982);
nand U7445 (N_7445,N_3959,N_4966);
nor U7446 (N_7446,N_2869,N_2517);
or U7447 (N_7447,N_3080,N_2726);
or U7448 (N_7448,N_2517,N_3692);
nor U7449 (N_7449,N_4765,N_2912);
xor U7450 (N_7450,N_4712,N_4860);
xnor U7451 (N_7451,N_4248,N_3655);
nor U7452 (N_7452,N_2534,N_2899);
nor U7453 (N_7453,N_4039,N_4886);
xnor U7454 (N_7454,N_3702,N_2535);
and U7455 (N_7455,N_4613,N_2740);
or U7456 (N_7456,N_4929,N_4607);
and U7457 (N_7457,N_3424,N_4537);
and U7458 (N_7458,N_4337,N_3534);
nand U7459 (N_7459,N_3061,N_3481);
nor U7460 (N_7460,N_3040,N_3995);
xnor U7461 (N_7461,N_4913,N_4610);
xor U7462 (N_7462,N_4462,N_3166);
nor U7463 (N_7463,N_3771,N_3061);
xor U7464 (N_7464,N_3792,N_3748);
xor U7465 (N_7465,N_3713,N_2777);
and U7466 (N_7466,N_3366,N_3321);
and U7467 (N_7467,N_3195,N_3422);
nand U7468 (N_7468,N_3185,N_3728);
or U7469 (N_7469,N_2837,N_3822);
xor U7470 (N_7470,N_3134,N_4194);
or U7471 (N_7471,N_3951,N_4187);
xor U7472 (N_7472,N_3696,N_2818);
or U7473 (N_7473,N_4136,N_3547);
or U7474 (N_7474,N_3713,N_3434);
or U7475 (N_7475,N_2928,N_3247);
or U7476 (N_7476,N_3950,N_3215);
nor U7477 (N_7477,N_4556,N_3244);
xor U7478 (N_7478,N_4064,N_2914);
or U7479 (N_7479,N_4343,N_4951);
and U7480 (N_7480,N_4847,N_2838);
nor U7481 (N_7481,N_3077,N_3767);
nand U7482 (N_7482,N_3769,N_3954);
xor U7483 (N_7483,N_4163,N_4015);
xnor U7484 (N_7484,N_4986,N_2785);
and U7485 (N_7485,N_4639,N_3532);
nor U7486 (N_7486,N_4804,N_4545);
or U7487 (N_7487,N_3772,N_3024);
and U7488 (N_7488,N_3254,N_3631);
xor U7489 (N_7489,N_2513,N_4987);
nor U7490 (N_7490,N_3180,N_3509);
nand U7491 (N_7491,N_2936,N_3018);
nand U7492 (N_7492,N_3800,N_4465);
or U7493 (N_7493,N_2640,N_3079);
or U7494 (N_7494,N_4281,N_4116);
and U7495 (N_7495,N_4077,N_4015);
and U7496 (N_7496,N_3206,N_2733);
xor U7497 (N_7497,N_4180,N_3386);
or U7498 (N_7498,N_4429,N_4194);
or U7499 (N_7499,N_3932,N_4340);
nand U7500 (N_7500,N_6016,N_7026);
nand U7501 (N_7501,N_5772,N_7292);
or U7502 (N_7502,N_7205,N_6636);
xnor U7503 (N_7503,N_7311,N_7226);
or U7504 (N_7504,N_7279,N_6521);
or U7505 (N_7505,N_5151,N_5918);
nor U7506 (N_7506,N_6781,N_6829);
xnor U7507 (N_7507,N_6845,N_5386);
nor U7508 (N_7508,N_5953,N_6649);
and U7509 (N_7509,N_6396,N_7437);
nor U7510 (N_7510,N_5715,N_6243);
xor U7511 (N_7511,N_6690,N_5216);
and U7512 (N_7512,N_7184,N_6795);
or U7513 (N_7513,N_6998,N_5399);
nor U7514 (N_7514,N_5242,N_6878);
nand U7515 (N_7515,N_7386,N_6473);
nand U7516 (N_7516,N_5334,N_5064);
xor U7517 (N_7517,N_5722,N_7455);
or U7518 (N_7518,N_6325,N_5811);
nand U7519 (N_7519,N_5300,N_6793);
nor U7520 (N_7520,N_5484,N_6430);
xnor U7521 (N_7521,N_5747,N_5585);
nand U7522 (N_7522,N_5054,N_7350);
and U7523 (N_7523,N_6967,N_6848);
xnor U7524 (N_7524,N_5879,N_5223);
and U7525 (N_7525,N_6527,N_5114);
or U7526 (N_7526,N_6093,N_6697);
nand U7527 (N_7527,N_5143,N_6858);
and U7528 (N_7528,N_5600,N_5946);
xnor U7529 (N_7529,N_6515,N_5705);
xor U7530 (N_7530,N_5530,N_5792);
nand U7531 (N_7531,N_5105,N_6782);
nor U7532 (N_7532,N_6134,N_5723);
or U7533 (N_7533,N_6497,N_6284);
nor U7534 (N_7534,N_6030,N_5572);
nor U7535 (N_7535,N_5289,N_5311);
xnor U7536 (N_7536,N_6338,N_7346);
nor U7537 (N_7537,N_7086,N_6202);
nand U7538 (N_7538,N_5767,N_5032);
or U7539 (N_7539,N_7272,N_6850);
nand U7540 (N_7540,N_6227,N_6112);
nor U7541 (N_7541,N_6714,N_6774);
or U7542 (N_7542,N_5661,N_7293);
nor U7543 (N_7543,N_6180,N_6142);
xnor U7544 (N_7544,N_6021,N_6882);
xnor U7545 (N_7545,N_6417,N_6075);
and U7546 (N_7546,N_6276,N_5084);
nand U7547 (N_7547,N_5213,N_5382);
and U7548 (N_7548,N_7207,N_6588);
nand U7549 (N_7549,N_5652,N_5999);
or U7550 (N_7550,N_7446,N_7489);
nand U7551 (N_7551,N_5874,N_7299);
xnor U7552 (N_7552,N_5256,N_6990);
and U7553 (N_7553,N_6218,N_7370);
nor U7554 (N_7554,N_5215,N_7373);
nor U7555 (N_7555,N_6370,N_6116);
nor U7556 (N_7556,N_7122,N_7248);
nor U7557 (N_7557,N_6265,N_6778);
xnor U7558 (N_7558,N_6427,N_6738);
xnor U7559 (N_7559,N_5310,N_6494);
nand U7560 (N_7560,N_6916,N_5196);
nand U7561 (N_7561,N_7430,N_5610);
or U7562 (N_7562,N_7404,N_7075);
xnor U7563 (N_7563,N_5551,N_5915);
nand U7564 (N_7564,N_5886,N_5859);
and U7565 (N_7565,N_6368,N_6268);
nor U7566 (N_7566,N_5616,N_7286);
xor U7567 (N_7567,N_6761,N_7008);
nor U7568 (N_7568,N_5589,N_6522);
nor U7569 (N_7569,N_6905,N_5603);
and U7570 (N_7570,N_5494,N_6443);
and U7571 (N_7571,N_6127,N_6852);
nor U7572 (N_7572,N_6006,N_5955);
nand U7573 (N_7573,N_6864,N_5302);
and U7574 (N_7574,N_5865,N_6216);
or U7575 (N_7575,N_6395,N_6136);
xor U7576 (N_7576,N_5881,N_6766);
nor U7577 (N_7577,N_6971,N_6230);
or U7578 (N_7578,N_7478,N_6183);
nand U7579 (N_7579,N_7260,N_6692);
xnor U7580 (N_7580,N_6656,N_7278);
and U7581 (N_7581,N_5895,N_6593);
nand U7582 (N_7582,N_5158,N_7481);
or U7583 (N_7583,N_6352,N_5303);
nor U7584 (N_7584,N_7179,N_7264);
nor U7585 (N_7585,N_6303,N_7423);
nor U7586 (N_7586,N_6869,N_6996);
xor U7587 (N_7587,N_6658,N_6099);
or U7588 (N_7588,N_5155,N_5570);
nand U7589 (N_7589,N_5081,N_6958);
nor U7590 (N_7590,N_7444,N_7425);
nand U7591 (N_7591,N_5543,N_7103);
xnor U7592 (N_7592,N_5743,N_7325);
or U7593 (N_7593,N_5327,N_5854);
xor U7594 (N_7594,N_6818,N_5470);
or U7595 (N_7595,N_5617,N_6548);
and U7596 (N_7596,N_5248,N_7115);
or U7597 (N_7597,N_5230,N_5748);
and U7598 (N_7598,N_5855,N_5745);
and U7599 (N_7599,N_7062,N_6063);
xnor U7600 (N_7600,N_7309,N_5631);
and U7601 (N_7601,N_5699,N_7335);
and U7602 (N_7602,N_5241,N_7332);
nor U7603 (N_7603,N_6817,N_7051);
nand U7604 (N_7604,N_5940,N_5165);
xnor U7605 (N_7605,N_7084,N_5036);
and U7606 (N_7606,N_6087,N_5059);
xnor U7607 (N_7607,N_5800,N_6000);
xnor U7608 (N_7608,N_5046,N_5683);
xor U7609 (N_7609,N_6643,N_5562);
xnor U7610 (N_7610,N_6010,N_7055);
xor U7611 (N_7611,N_6820,N_5420);
nor U7612 (N_7612,N_7191,N_5313);
nor U7613 (N_7613,N_6675,N_6082);
and U7614 (N_7614,N_6729,N_6269);
xor U7615 (N_7615,N_6982,N_6693);
or U7616 (N_7616,N_6966,N_7022);
nor U7617 (N_7617,N_6399,N_5089);
and U7618 (N_7618,N_5424,N_6271);
nand U7619 (N_7619,N_5137,N_5272);
nor U7620 (N_7620,N_6258,N_5057);
or U7621 (N_7621,N_5167,N_5134);
xnor U7622 (N_7622,N_5473,N_5759);
xnor U7623 (N_7623,N_5243,N_5169);
nand U7624 (N_7624,N_5411,N_6172);
xnor U7625 (N_7625,N_6932,N_5538);
xnor U7626 (N_7626,N_5459,N_6659);
xor U7627 (N_7627,N_7052,N_6550);
xnor U7628 (N_7628,N_5487,N_7208);
and U7629 (N_7629,N_7464,N_5279);
and U7630 (N_7630,N_7372,N_5594);
nand U7631 (N_7631,N_6120,N_5808);
nor U7632 (N_7632,N_7011,N_6144);
xnor U7633 (N_7633,N_5725,N_5132);
nor U7634 (N_7634,N_6193,N_5768);
or U7635 (N_7635,N_6740,N_7067);
xor U7636 (N_7636,N_6737,N_5116);
xnor U7637 (N_7637,N_6613,N_5913);
or U7638 (N_7638,N_7039,N_7210);
xnor U7639 (N_7639,N_7030,N_5344);
and U7640 (N_7640,N_7475,N_7465);
and U7641 (N_7641,N_5878,N_6981);
xor U7642 (N_7642,N_6286,N_5101);
and U7643 (N_7643,N_6107,N_7043);
nor U7644 (N_7644,N_6379,N_6867);
and U7645 (N_7645,N_7237,N_6100);
and U7646 (N_7646,N_7017,N_6005);
nor U7647 (N_7647,N_6745,N_6956);
nand U7648 (N_7648,N_7159,N_6547);
nor U7649 (N_7649,N_6987,N_5995);
nand U7650 (N_7650,N_6054,N_5709);
nand U7651 (N_7651,N_7148,N_5546);
nor U7652 (N_7652,N_5065,N_5210);
or U7653 (N_7653,N_6915,N_5740);
nor U7654 (N_7654,N_5703,N_5188);
and U7655 (N_7655,N_5736,N_6195);
or U7656 (N_7656,N_7046,N_5107);
nand U7657 (N_7657,N_6512,N_6209);
xor U7658 (N_7658,N_6783,N_7190);
or U7659 (N_7659,N_5067,N_6407);
xor U7660 (N_7660,N_6385,N_6194);
xor U7661 (N_7661,N_6211,N_6929);
xor U7662 (N_7662,N_6660,N_6799);
xor U7663 (N_7663,N_6632,N_6534);
nor U7664 (N_7664,N_7170,N_7238);
nand U7665 (N_7665,N_5380,N_7314);
and U7666 (N_7666,N_5754,N_6191);
xnor U7667 (N_7667,N_7076,N_6391);
nand U7668 (N_7668,N_6484,N_5219);
and U7669 (N_7669,N_6712,N_6239);
or U7670 (N_7670,N_7174,N_5030);
nand U7671 (N_7671,N_5283,N_7059);
and U7672 (N_7672,N_5710,N_6415);
nor U7673 (N_7673,N_6498,N_6772);
xor U7674 (N_7674,N_6721,N_5437);
nor U7675 (N_7675,N_7415,N_5891);
or U7676 (N_7676,N_6641,N_7479);
nand U7677 (N_7677,N_6517,N_5672);
and U7678 (N_7678,N_7232,N_5689);
and U7679 (N_7679,N_5117,N_5016);
xnor U7680 (N_7680,N_5047,N_5611);
or U7681 (N_7681,N_7436,N_6700);
nor U7682 (N_7682,N_5477,N_7296);
xor U7683 (N_7683,N_7410,N_6347);
xnor U7684 (N_7684,N_6296,N_6507);
xnor U7685 (N_7685,N_5802,N_6896);
nor U7686 (N_7686,N_6710,N_5471);
nand U7687 (N_7687,N_5247,N_6114);
xnor U7688 (N_7688,N_6167,N_7009);
and U7689 (N_7689,N_6487,N_7355);
xor U7690 (N_7690,N_6836,N_6215);
xnor U7691 (N_7691,N_5025,N_6462);
and U7692 (N_7692,N_6029,N_5154);
or U7693 (N_7693,N_5157,N_5325);
xor U7694 (N_7694,N_7078,N_5385);
nand U7695 (N_7695,N_6015,N_5130);
nand U7696 (N_7696,N_6376,N_5920);
nand U7697 (N_7697,N_6143,N_7164);
and U7698 (N_7698,N_5847,N_6166);
and U7699 (N_7699,N_7048,N_7071);
nand U7700 (N_7700,N_7169,N_5907);
and U7701 (N_7701,N_6023,N_5642);
xor U7702 (N_7702,N_5897,N_6925);
or U7703 (N_7703,N_5189,N_5989);
nand U7704 (N_7704,N_6270,N_5527);
or U7705 (N_7705,N_7428,N_5712);
nand U7706 (N_7706,N_5676,N_6827);
nor U7707 (N_7707,N_6317,N_5875);
or U7708 (N_7708,N_6861,N_5192);
or U7709 (N_7709,N_7198,N_6502);
and U7710 (N_7710,N_5163,N_6383);
nand U7711 (N_7711,N_6868,N_6092);
or U7712 (N_7712,N_6233,N_6404);
nand U7713 (N_7713,N_5852,N_7441);
xnor U7714 (N_7714,N_6957,N_7131);
or U7715 (N_7715,N_5756,N_6685);
nor U7716 (N_7716,N_6559,N_5693);
or U7717 (N_7717,N_6393,N_6965);
nand U7718 (N_7718,N_5402,N_5927);
and U7719 (N_7719,N_5371,N_6314);
and U7720 (N_7720,N_7044,N_7054);
nand U7721 (N_7721,N_6285,N_6595);
xnor U7722 (N_7722,N_5304,N_5894);
or U7723 (N_7723,N_5842,N_6477);
and U7724 (N_7724,N_6111,N_5435);
or U7725 (N_7725,N_7382,N_6475);
nor U7726 (N_7726,N_6549,N_5338);
xor U7727 (N_7727,N_6241,N_5633);
or U7728 (N_7728,N_6267,N_5680);
nor U7729 (N_7729,N_6125,N_7412);
xor U7730 (N_7730,N_5446,N_5977);
and U7731 (N_7731,N_5015,N_6997);
or U7732 (N_7732,N_6942,N_7163);
nor U7733 (N_7733,N_5615,N_7091);
nand U7734 (N_7734,N_5651,N_7168);
nand U7735 (N_7735,N_6717,N_7351);
nand U7736 (N_7736,N_6625,N_5028);
nor U7737 (N_7737,N_5466,N_6968);
and U7738 (N_7738,N_5902,N_6592);
xnor U7739 (N_7739,N_5390,N_7394);
or U7740 (N_7740,N_6913,N_6739);
and U7741 (N_7741,N_5586,N_6574);
and U7742 (N_7742,N_6553,N_6519);
and U7743 (N_7743,N_6500,N_5352);
and U7744 (N_7744,N_6945,N_6678);
and U7745 (N_7745,N_6558,N_5391);
nand U7746 (N_7746,N_7089,N_6071);
and U7747 (N_7747,N_5899,N_5171);
and U7748 (N_7748,N_5412,N_6441);
xnor U7749 (N_7749,N_6482,N_6287);
or U7750 (N_7750,N_5249,N_5587);
and U7751 (N_7751,N_5257,N_5877);
and U7752 (N_7752,N_7391,N_6062);
and U7753 (N_7753,N_6779,N_5893);
and U7754 (N_7754,N_5770,N_5716);
xnor U7755 (N_7755,N_5765,N_7414);
and U7756 (N_7756,N_6851,N_6214);
and U7757 (N_7757,N_5836,N_7105);
or U7758 (N_7758,N_6077,N_5614);
nor U7759 (N_7759,N_5376,N_5039);
or U7760 (N_7760,N_6066,N_6436);
and U7761 (N_7761,N_5975,N_5850);
nand U7762 (N_7762,N_5654,N_7038);
xor U7763 (N_7763,N_7211,N_5641);
and U7764 (N_7764,N_5244,N_6946);
or U7765 (N_7765,N_5845,N_6964);
or U7766 (N_7766,N_6885,N_6505);
xnor U7767 (N_7767,N_7393,N_5483);
xnor U7768 (N_7768,N_5994,N_5100);
nand U7769 (N_7769,N_5834,N_6792);
or U7770 (N_7770,N_5427,N_6131);
and U7771 (N_7771,N_6831,N_6380);
xor U7772 (N_7772,N_5212,N_6872);
or U7773 (N_7773,N_6554,N_5504);
and U7774 (N_7774,N_5450,N_7321);
nor U7775 (N_7775,N_7140,N_6406);
and U7776 (N_7776,N_6833,N_5892);
nand U7777 (N_7777,N_6589,N_7135);
xnor U7778 (N_7778,N_5787,N_6049);
and U7779 (N_7779,N_6065,N_5185);
nor U7780 (N_7780,N_5866,N_5406);
nor U7781 (N_7781,N_5306,N_5305);
or U7782 (N_7782,N_5038,N_5941);
or U7783 (N_7783,N_7406,N_6562);
nor U7784 (N_7784,N_5764,N_6624);
nor U7785 (N_7785,N_6291,N_5111);
nor U7786 (N_7786,N_5438,N_7396);
xor U7787 (N_7787,N_5298,N_5087);
nand U7788 (N_7788,N_6040,N_5726);
nor U7789 (N_7789,N_5801,N_5822);
and U7790 (N_7790,N_6518,N_5627);
and U7791 (N_7791,N_5618,N_5880);
and U7792 (N_7792,N_5246,N_5448);
nand U7793 (N_7793,N_6485,N_5394);
xnor U7794 (N_7794,N_6153,N_5180);
and U7795 (N_7795,N_7186,N_7066);
or U7796 (N_7796,N_6552,N_6642);
xnor U7797 (N_7797,N_7345,N_6826);
and U7798 (N_7798,N_5904,N_7035);
or U7799 (N_7799,N_6033,N_6506);
xor U7800 (N_7800,N_7100,N_5443);
nand U7801 (N_7801,N_6674,N_7294);
nor U7802 (N_7802,N_6392,N_6053);
or U7803 (N_7803,N_5432,N_7124);
or U7804 (N_7804,N_5735,N_7165);
or U7805 (N_7805,N_5049,N_5796);
nor U7806 (N_7806,N_5358,N_5001);
and U7807 (N_7807,N_6622,N_5673);
nand U7808 (N_7808,N_6504,N_6734);
nand U7809 (N_7809,N_7416,N_5308);
nor U7810 (N_7810,N_7120,N_7228);
and U7811 (N_7811,N_6496,N_5602);
nand U7812 (N_7812,N_5541,N_6955);
nand U7813 (N_7813,N_7171,N_6004);
or U7814 (N_7814,N_6930,N_6924);
nand U7815 (N_7815,N_6953,N_7323);
xor U7816 (N_7816,N_6252,N_5199);
nand U7817 (N_7817,N_7023,N_6117);
nor U7818 (N_7818,N_5621,N_6977);
xor U7819 (N_7819,N_6897,N_6264);
and U7820 (N_7820,N_5809,N_6297);
nand U7821 (N_7821,N_6571,N_5009);
nor U7822 (N_7822,N_7007,N_5718);
or U7823 (N_7823,N_5550,N_5156);
xor U7824 (N_7824,N_6476,N_5867);
xnor U7825 (N_7825,N_5079,N_5112);
nand U7826 (N_7826,N_5813,N_7491);
nor U7827 (N_7827,N_5378,N_5685);
nor U7828 (N_7828,N_5564,N_7467);
or U7829 (N_7829,N_6654,N_5119);
nand U7830 (N_7830,N_5947,N_7127);
and U7831 (N_7831,N_5649,N_6031);
and U7832 (N_7832,N_7287,N_5195);
nand U7833 (N_7833,N_7461,N_6587);
xor U7834 (N_7834,N_5912,N_5010);
xnor U7835 (N_7835,N_5348,N_6866);
xnor U7836 (N_7836,N_6979,N_6823);
nor U7837 (N_7837,N_6822,N_5372);
or U7838 (N_7838,N_5949,N_7252);
xor U7839 (N_7839,N_5532,N_7360);
nand U7840 (N_7840,N_6157,N_5981);
or U7841 (N_7841,N_5779,N_5831);
xor U7842 (N_7842,N_6723,N_6152);
and U7843 (N_7843,N_6309,N_6046);
xnor U7844 (N_7844,N_6451,N_7267);
or U7845 (N_7845,N_7126,N_5750);
and U7846 (N_7846,N_5857,N_7063);
or U7847 (N_7847,N_5853,N_6647);
nand U7848 (N_7848,N_6047,N_5403);
nor U7849 (N_7849,N_5301,N_6532);
nand U7850 (N_7850,N_5023,N_5851);
or U7851 (N_7851,N_6640,N_7367);
and U7852 (N_7852,N_7167,N_6203);
xnor U7853 (N_7853,N_7214,N_6057);
nor U7854 (N_7854,N_6280,N_7173);
xor U7855 (N_7855,N_6181,N_5276);
or U7856 (N_7856,N_6089,N_6699);
or U7857 (N_7857,N_5362,N_5198);
and U7858 (N_7858,N_7487,N_6491);
xor U7859 (N_7859,N_5653,N_5200);
xnor U7860 (N_7860,N_6493,N_7216);
xor U7861 (N_7861,N_5284,N_6886);
nand U7862 (N_7862,N_6048,N_5336);
nand U7863 (N_7863,N_6598,N_6350);
nand U7864 (N_7864,N_6008,N_6403);
nand U7865 (N_7865,N_7337,N_6566);
nor U7866 (N_7866,N_5291,N_6735);
nor U7867 (N_7867,N_6807,N_6090);
nand U7868 (N_7868,N_6912,N_5636);
nand U7869 (N_7869,N_6880,N_7096);
and U7870 (N_7870,N_5565,N_5815);
xnor U7871 (N_7871,N_7177,N_6013);
and U7872 (N_7872,N_5667,N_5396);
nor U7873 (N_7873,N_5178,N_5004);
or U7874 (N_7874,N_7324,N_6810);
xor U7875 (N_7875,N_7357,N_6765);
nand U7876 (N_7876,N_5674,N_5969);
nor U7877 (N_7877,N_6097,N_6910);
xor U7878 (N_7878,N_6056,N_6240);
nor U7879 (N_7879,N_7476,N_6121);
and U7880 (N_7880,N_5197,N_5656);
and U7881 (N_7881,N_5806,N_7003);
nor U7882 (N_7882,N_6652,N_5051);
nand U7883 (N_7883,N_6199,N_7098);
nor U7884 (N_7884,N_6386,N_6606);
xor U7885 (N_7885,N_5884,N_6224);
and U7886 (N_7886,N_5882,N_6843);
or U7887 (N_7887,N_6985,N_7195);
and U7888 (N_7888,N_7347,N_6551);
nor U7889 (N_7889,N_7326,N_6110);
and U7890 (N_7890,N_6235,N_6607);
or U7891 (N_7891,N_6422,N_7484);
or U7892 (N_7892,N_7155,N_6938);
nor U7893 (N_7893,N_5960,N_6619);
nand U7894 (N_7894,N_6219,N_5980);
xnor U7895 (N_7895,N_5509,N_5194);
or U7896 (N_7896,N_6537,N_7315);
nor U7897 (N_7897,N_7150,N_6752);
and U7898 (N_7898,N_6342,N_5755);
or U7899 (N_7899,N_6020,N_6648);
or U7900 (N_7900,N_5388,N_6777);
xor U7901 (N_7901,N_5581,N_6095);
and U7902 (N_7902,N_5416,N_7204);
or U7903 (N_7903,N_6797,N_7041);
nor U7904 (N_7904,N_6960,N_5804);
and U7905 (N_7905,N_5374,N_5896);
or U7906 (N_7906,N_5033,N_7320);
nand U7907 (N_7907,N_5395,N_5700);
nand U7908 (N_7908,N_6844,N_5007);
xnor U7909 (N_7909,N_6716,N_6454);
xnor U7910 (N_7910,N_5035,N_6124);
nand U7911 (N_7911,N_7130,N_6159);
or U7912 (N_7912,N_6511,N_6465);
nor U7913 (N_7913,N_5053,N_5552);
or U7914 (N_7914,N_7342,N_5252);
and U7915 (N_7915,N_7364,N_6748);
nor U7916 (N_7916,N_6374,N_5356);
nand U7917 (N_7917,N_5042,N_7276);
and U7918 (N_7918,N_6992,N_6328);
and U7919 (N_7919,N_5871,N_7102);
or U7920 (N_7920,N_5675,N_5445);
nand U7921 (N_7921,N_7015,N_6251);
nand U7922 (N_7922,N_6220,N_5335);
or U7923 (N_7923,N_7443,N_5534);
nand U7924 (N_7924,N_7049,N_5000);
and U7925 (N_7925,N_6446,N_5540);
or U7926 (N_7926,N_6816,N_7136);
xor U7927 (N_7927,N_5906,N_5976);
xnor U7928 (N_7928,N_7318,N_5273);
nand U7929 (N_7929,N_5182,N_5255);
xor U7930 (N_7930,N_6150,N_7322);
nand U7931 (N_7931,N_6129,N_5688);
nand U7932 (N_7932,N_5956,N_7058);
or U7933 (N_7933,N_6510,N_5844);
nor U7934 (N_7934,N_7329,N_5596);
nand U7935 (N_7935,N_7217,N_5500);
nor U7936 (N_7936,N_5934,N_5021);
nor U7937 (N_7937,N_6612,N_7079);
or U7938 (N_7938,N_5330,N_6991);
and U7939 (N_7939,N_5474,N_5456);
or U7940 (N_7940,N_7270,N_5418);
or U7941 (N_7941,N_5545,N_5463);
and U7942 (N_7942,N_6951,N_7439);
nand U7943 (N_7943,N_5331,N_6601);
xor U7944 (N_7944,N_6344,N_7392);
nand U7945 (N_7945,N_5591,N_5074);
or U7946 (N_7946,N_6384,N_5259);
or U7947 (N_7947,N_5662,N_6791);
or U7948 (N_7948,N_7497,N_7451);
nand U7949 (N_7949,N_7339,N_5821);
xnor U7950 (N_7950,N_6324,N_6170);
nor U7951 (N_7951,N_5939,N_7317);
nor U7952 (N_7952,N_6891,N_5864);
and U7953 (N_7953,N_5011,N_7244);
and U7954 (N_7954,N_7014,N_7457);
nand U7955 (N_7955,N_6175,N_5537);
nor U7956 (N_7956,N_6094,N_7285);
xor U7957 (N_7957,N_6911,N_7137);
or U7958 (N_7958,N_7053,N_5141);
nand U7959 (N_7959,N_5398,N_6801);
xnor U7960 (N_7960,N_6664,N_5104);
or U7961 (N_7961,N_7298,N_5783);
nor U7962 (N_7962,N_7001,N_7227);
nand U7963 (N_7963,N_5274,N_7468);
and U7964 (N_7964,N_6316,N_5166);
nor U7965 (N_7965,N_7129,N_6205);
nor U7966 (N_7966,N_6307,N_6546);
or U7967 (N_7967,N_5826,N_5733);
or U7968 (N_7968,N_6130,N_5965);
and U7969 (N_7969,N_7450,N_5098);
and U7970 (N_7970,N_5319,N_6390);
xnor U7971 (N_7971,N_7407,N_6800);
nor U7972 (N_7972,N_5837,N_7398);
or U7973 (N_7973,N_6244,N_5753);
xnor U7974 (N_7974,N_5433,N_6954);
and U7975 (N_7975,N_7250,N_6755);
nor U7976 (N_7976,N_6969,N_7010);
xnor U7977 (N_7977,N_5265,N_7308);
nor U7978 (N_7978,N_7019,N_6151);
nand U7979 (N_7979,N_7376,N_7175);
nor U7980 (N_7980,N_7469,N_7380);
nand U7981 (N_7981,N_6819,N_5397);
xnor U7982 (N_7982,N_5342,N_5440);
and U7983 (N_7983,N_6630,N_5512);
and U7984 (N_7984,N_6530,N_5357);
nor U7985 (N_7985,N_7271,N_5077);
and U7986 (N_7986,N_6043,N_6146);
xnor U7987 (N_7987,N_6017,N_5027);
and U7988 (N_7988,N_6847,N_7256);
nor U7989 (N_7989,N_7132,N_7005);
nor U7990 (N_7990,N_5677,N_5936);
and U7991 (N_7991,N_5945,N_5095);
and U7992 (N_7992,N_6295,N_5522);
xnor U7993 (N_7993,N_5905,N_7133);
and U7994 (N_7994,N_7025,N_7183);
nor U7995 (N_7995,N_5479,N_5365);
nand U7996 (N_7996,N_5052,N_6917);
nor U7997 (N_7997,N_7417,N_5619);
xnor U7998 (N_7998,N_6719,N_5268);
and U7999 (N_7999,N_5092,N_6322);
or U8000 (N_8000,N_5938,N_5341);
xnor U8001 (N_8001,N_5914,N_7146);
and U8002 (N_8002,N_5235,N_6361);
nor U8003 (N_8003,N_5266,N_5961);
xnor U8004 (N_8004,N_5774,N_6545);
nor U8005 (N_8005,N_6616,N_6903);
nor U8006 (N_8006,N_6813,N_5322);
xor U8007 (N_8007,N_6952,N_6382);
or U8008 (N_8008,N_5103,N_5187);
or U8009 (N_8009,N_5597,N_7460);
or U8010 (N_8010,N_6055,N_7379);
xnor U8011 (N_8011,N_7193,N_6771);
nand U8012 (N_8012,N_5580,N_6963);
and U8013 (N_8013,N_7377,N_7004);
nand U8014 (N_8014,N_6689,N_7247);
xor U8015 (N_8015,N_5138,N_5405);
nor U8016 (N_8016,N_6542,N_5655);
xor U8017 (N_8017,N_5353,N_5634);
and U8018 (N_8018,N_6975,N_5436);
xor U8019 (N_8019,N_6661,N_6464);
nand U8020 (N_8020,N_5490,N_6814);
and U8021 (N_8021,N_5840,N_5558);
xnor U8022 (N_8022,N_5560,N_5493);
xnor U8023 (N_8023,N_6154,N_7283);
xor U8024 (N_8024,N_7018,N_6785);
xnor U8025 (N_8025,N_5109,N_7142);
nor U8026 (N_8026,N_6078,N_7427);
and U8027 (N_8027,N_7197,N_5556);
xnor U8028 (N_8028,N_5451,N_6806);
xnor U8029 (N_8029,N_6533,N_7243);
nor U8030 (N_8030,N_5080,N_5535);
nand U8031 (N_8031,N_7161,N_6703);
and U8032 (N_8032,N_5696,N_7378);
or U8033 (N_8033,N_7249,N_7108);
or U8034 (N_8034,N_5296,N_6790);
and U8035 (N_8035,N_7288,N_7157);
xor U8036 (N_8036,N_7234,N_6600);
nor U8037 (N_8037,N_6028,N_6257);
or U8038 (N_8038,N_6927,N_6525);
or U8039 (N_8039,N_5846,N_6081);
or U8040 (N_8040,N_6914,N_6334);
or U8041 (N_8041,N_5607,N_6709);
or U8042 (N_8042,N_6898,N_6989);
nand U8043 (N_8043,N_6926,N_5227);
nor U8044 (N_8044,N_6242,N_7012);
xor U8045 (N_8045,N_7236,N_5697);
xor U8046 (N_8046,N_6459,N_7421);
or U8047 (N_8047,N_7397,N_6186);
nand U8048 (N_8048,N_5773,N_5136);
nor U8049 (N_8049,N_5232,N_5873);
nand U8050 (N_8050,N_6775,N_5024);
nand U8051 (N_8051,N_5521,N_5507);
or U8052 (N_8052,N_5972,N_5088);
and U8053 (N_8053,N_7031,N_6169);
or U8054 (N_8054,N_6604,N_5316);
xnor U8055 (N_8055,N_5229,N_5019);
nor U8056 (N_8056,N_6260,N_6637);
xor U8057 (N_8057,N_6085,N_6884);
nand U8058 (N_8058,N_6478,N_6544);
or U8059 (N_8059,N_7114,N_5663);
and U8060 (N_8060,N_5203,N_6222);
xnor U8061 (N_8061,N_6109,N_7400);
nor U8062 (N_8062,N_7162,N_6277);
and U8063 (N_8063,N_5579,N_6821);
and U8064 (N_8064,N_6160,N_5135);
nand U8065 (N_8065,N_7149,N_6680);
xor U8066 (N_8066,N_6171,N_7006);
and U8067 (N_8067,N_5281,N_7356);
nor U8068 (N_8068,N_7456,N_7110);
or U8069 (N_8069,N_6849,N_6132);
nand U8070 (N_8070,N_7483,N_5208);
and U8071 (N_8071,N_6928,N_6434);
or U8072 (N_8072,N_5048,N_5665);
nor U8073 (N_8073,N_5290,N_7399);
and U8074 (N_8074,N_5225,N_7448);
and U8075 (N_8075,N_5254,N_6207);
nor U8076 (N_8076,N_7362,N_6003);
and U8077 (N_8077,N_6803,N_6340);
or U8078 (N_8078,N_7034,N_6210);
nand U8079 (N_8079,N_5118,N_6306);
xor U8080 (N_8080,N_7212,N_5383);
nand U8081 (N_8081,N_5963,N_5606);
and U8082 (N_8082,N_5812,N_6770);
nor U8083 (N_8083,N_7452,N_7281);
xor U8084 (N_8084,N_5595,N_7463);
nor U8085 (N_8085,N_5567,N_5860);
nor U8086 (N_8086,N_6375,N_5078);
xnor U8087 (N_8087,N_5122,N_6623);
nand U8088 (N_8088,N_6174,N_7125);
or U8089 (N_8089,N_6012,N_5682);
and U8090 (N_8090,N_6934,N_7429);
or U8091 (N_8091,N_6014,N_5339);
and U8092 (N_8092,N_5954,N_6842);
or U8093 (N_8093,N_6450,N_7466);
and U8094 (N_8094,N_6139,N_5161);
nor U8095 (N_8095,N_5455,N_6671);
xor U8096 (N_8096,N_6730,N_5250);
nand U8097 (N_8097,N_7082,N_7353);
xor U8098 (N_8098,N_6348,N_5498);
and U8099 (N_8099,N_5314,N_6586);
or U8100 (N_8100,N_6122,N_5234);
nor U8101 (N_8101,N_7033,N_5986);
and U8102 (N_8102,N_5097,N_5701);
nand U8103 (N_8103,N_6319,N_6261);
nor U8104 (N_8104,N_5911,N_5605);
xnor U8105 (N_8105,N_7061,N_7295);
or U8106 (N_8106,N_6103,N_5499);
nor U8107 (N_8107,N_7368,N_5549);
nor U8108 (N_8108,N_6433,N_5876);
or U8109 (N_8109,N_5093,N_7361);
or U8110 (N_8110,N_6669,N_6610);
nor U8111 (N_8111,N_7057,N_6919);
nor U8112 (N_8112,N_6300,N_5031);
nor U8113 (N_8113,N_6749,N_6560);
or U8114 (N_8114,N_6569,N_6358);
or U8115 (N_8115,N_5669,N_5045);
xnor U8116 (N_8116,N_7266,N_7381);
nor U8117 (N_8117,N_7220,N_5037);
nor U8118 (N_8118,N_5657,N_5422);
or U8119 (N_8119,N_6448,N_7021);
xnor U8120 (N_8120,N_7000,N_5205);
or U8121 (N_8121,N_6133,N_6409);
or U8122 (N_8122,N_5520,N_5501);
and U8123 (N_8123,N_6321,N_5979);
nor U8124 (N_8124,N_7242,N_6304);
nor U8125 (N_8125,N_5544,N_6995);
nand U8126 (N_8126,N_6027,N_7065);
nor U8127 (N_8127,N_5149,N_5069);
nor U8128 (N_8128,N_5909,N_5262);
or U8129 (N_8129,N_6711,N_6278);
or U8130 (N_8130,N_5990,N_5326);
nand U8131 (N_8131,N_6070,N_7192);
nand U8132 (N_8132,N_7490,N_7486);
nand U8133 (N_8133,N_6449,N_6363);
nand U8134 (N_8134,N_6161,N_5513);
nor U8135 (N_8135,N_6986,N_5434);
and U8136 (N_8136,N_5140,N_7420);
nand U8137 (N_8137,N_5209,N_6290);
nor U8138 (N_8138,N_6638,N_6611);
or U8139 (N_8139,N_6067,N_5108);
nand U8140 (N_8140,N_5014,N_5751);
nand U8141 (N_8141,N_6825,N_6688);
or U8142 (N_8142,N_6138,N_5070);
and U8143 (N_8143,N_5307,N_5312);
and U8144 (N_8144,N_7225,N_5278);
or U8145 (N_8145,N_6580,N_5983);
nand U8146 (N_8146,N_5373,N_5978);
nor U8147 (N_8147,N_6538,N_7185);
nor U8148 (N_8148,N_5006,N_5133);
and U8149 (N_8149,N_6389,N_5168);
nor U8150 (N_8150,N_5333,N_5791);
xor U8151 (N_8151,N_5233,N_5423);
or U8152 (N_8152,N_7194,N_6555);
and U8153 (N_8153,N_5147,N_6001);
and U8154 (N_8154,N_6101,N_6754);
or U8155 (N_8155,N_6948,N_5870);
nand U8156 (N_8156,N_5379,N_6556);
nor U8157 (N_8157,N_6044,N_6402);
and U8158 (N_8158,N_5730,N_5449);
xnor U8159 (N_8159,N_5758,N_5387);
and U8160 (N_8160,N_5355,N_6918);
and U8161 (N_8161,N_7087,N_5238);
nor U8162 (N_8162,N_5553,N_5883);
or U8163 (N_8163,N_6950,N_7366);
and U8164 (N_8164,N_6974,N_5719);
nor U8165 (N_8165,N_6411,N_6523);
xor U8166 (N_8166,N_5317,N_5659);
xor U8167 (N_8167,N_7029,N_6509);
nor U8168 (N_8168,N_5583,N_6874);
or U8169 (N_8169,N_5997,N_5777);
nor U8170 (N_8170,N_6708,N_5184);
nor U8171 (N_8171,N_5935,N_5299);
xor U8172 (N_8172,N_6543,N_6855);
xor U8173 (N_8173,N_7447,N_5354);
nand U8174 (N_8174,N_5511,N_7153);
nor U8175 (N_8175,N_6234,N_6335);
xor U8176 (N_8176,N_7401,N_6308);
xnor U8177 (N_8177,N_6731,N_6472);
nor U8178 (N_8178,N_5269,N_6457);
xnor U8179 (N_8179,N_5835,N_5381);
nand U8180 (N_8180,N_5050,N_6492);
and U8181 (N_8181,N_5439,N_6007);
and U8182 (N_8182,N_7369,N_5206);
xor U8183 (N_8183,N_7166,N_7411);
xnor U8184 (N_8184,N_6182,N_7116);
xnor U8185 (N_8185,N_5044,N_6582);
xor U8186 (N_8186,N_6440,N_5153);
nor U8187 (N_8187,N_5760,N_6682);
or U8188 (N_8188,N_5211,N_7387);
nor U8189 (N_8189,N_5343,N_6590);
xor U8190 (N_8190,N_6584,N_5970);
and U8191 (N_8191,N_6875,N_5728);
or U8192 (N_8192,N_5368,N_5624);
xnor U8193 (N_8193,N_5632,N_5810);
xor U8194 (N_8194,N_6428,N_7070);
nor U8195 (N_8195,N_6788,N_5769);
or U8196 (N_8196,N_7172,N_5584);
and U8197 (N_8197,N_5626,N_5516);
or U8198 (N_8198,N_5650,N_6331);
nor U8199 (N_8199,N_5598,N_7301);
nor U8200 (N_8200,N_7221,N_6732);
and U8201 (N_8201,N_6657,N_7310);
nor U8202 (N_8202,N_5838,N_7068);
and U8203 (N_8203,N_7255,N_6113);
and U8204 (N_8204,N_6983,N_5575);
nor U8205 (N_8205,N_5181,N_5741);
or U8206 (N_8206,N_6526,N_6367);
xor U8207 (N_8207,N_5058,N_5932);
or U8208 (N_8208,N_7040,N_6018);
xnor U8209 (N_8209,N_5771,N_7340);
or U8210 (N_8210,N_5441,N_5005);
or U8211 (N_8211,N_5749,N_5820);
and U8212 (N_8212,N_6993,N_5571);
or U8213 (N_8213,N_6663,N_5102);
or U8214 (N_8214,N_5542,N_5622);
or U8215 (N_8215,N_5497,N_5968);
xnor U8216 (N_8216,N_6236,N_5827);
or U8217 (N_8217,N_5679,N_6994);
xor U8218 (N_8218,N_6357,N_6301);
and U8219 (N_8219,N_6865,N_5757);
and U8220 (N_8220,N_5505,N_6333);
and U8221 (N_8221,N_5539,N_7077);
and U8222 (N_8222,N_6147,N_6631);
and U8223 (N_8223,N_7482,N_6603);
nand U8224 (N_8224,N_5734,N_6439);
nand U8225 (N_8225,N_5128,N_5115);
xnor U8226 (N_8226,N_5086,N_5508);
nor U8227 (N_8227,N_5569,N_7085);
and U8228 (N_8228,N_5294,N_5404);
nor U8229 (N_8229,N_7090,N_5987);
and U8230 (N_8230,N_5923,N_5126);
nor U8231 (N_8231,N_6602,N_6315);
nand U8232 (N_8232,N_6573,N_7147);
nand U8233 (N_8233,N_5060,N_6137);
xor U8234 (N_8234,N_6798,N_6597);
nor U8235 (N_8235,N_5055,N_5671);
nand U8236 (N_8236,N_5848,N_6064);
and U8237 (N_8237,N_5264,N_5629);
nand U8238 (N_8238,N_6426,N_7080);
nand U8239 (N_8239,N_6834,N_6293);
or U8240 (N_8240,N_5717,N_6198);
or U8241 (N_8241,N_5106,N_6460);
xnor U8242 (N_8242,N_5431,N_5858);
and U8243 (N_8243,N_7188,N_6811);
or U8244 (N_8244,N_5775,N_7494);
or U8245 (N_8245,N_5476,N_6653);
nor U8246 (N_8246,N_5170,N_7128);
or U8247 (N_8247,N_6453,N_5329);
nand U8248 (N_8248,N_6045,N_5561);
and U8249 (N_8249,N_6780,N_5592);
or U8250 (N_8250,N_6366,N_5599);
xnor U8251 (N_8251,N_5958,N_5407);
and U8252 (N_8252,N_5384,N_6468);
or U8253 (N_8253,N_6341,N_7180);
nor U8254 (N_8254,N_5782,N_7290);
or U8255 (N_8255,N_6086,N_6255);
nand U8256 (N_8256,N_5613,N_5309);
or U8257 (N_8257,N_6197,N_5825);
nand U8258 (N_8258,N_6398,N_6676);
nand U8259 (N_8259,N_5193,N_6581);
xnor U8260 (N_8260,N_6429,N_5690);
xnor U8261 (N_8261,N_6561,N_5514);
nor U8262 (N_8262,N_5351,N_5973);
or U8263 (N_8263,N_5828,N_6320);
and U8264 (N_8264,N_6895,N_5125);
xor U8265 (N_8265,N_5393,N_6050);
and U8266 (N_8266,N_5275,N_7470);
nand U8267 (N_8267,N_5410,N_7303);
nand U8268 (N_8268,N_6628,N_6165);
and U8269 (N_8269,N_6135,N_5781);
and U8270 (N_8270,N_6629,N_6900);
nor U8271 (N_8271,N_6838,N_7442);
and U8272 (N_8272,N_6299,N_5029);
nor U8273 (N_8273,N_5022,N_7106);
nor U8274 (N_8274,N_6349,N_6725);
and U8275 (N_8275,N_6539,N_6026);
xor U8276 (N_8276,N_6360,N_6416);
xor U8277 (N_8277,N_6254,N_6405);
or U8278 (N_8278,N_7316,N_7268);
nand U8279 (N_8279,N_6812,N_5292);
xor U8280 (N_8280,N_6332,N_6796);
nand U8281 (N_8281,N_5401,N_6776);
and U8282 (N_8282,N_7200,N_6456);
and U8283 (N_8283,N_6038,N_6035);
nor U8284 (N_8284,N_5179,N_5462);
or U8285 (N_8285,N_5123,N_6577);
nor U8286 (N_8286,N_5413,N_6196);
and U8287 (N_8287,N_6204,N_6514);
xnor U8288 (N_8288,N_5898,N_7438);
or U8289 (N_8289,N_6906,N_7385);
and U8290 (N_8290,N_5952,N_5625);
nand U8291 (N_8291,N_5465,N_6256);
nand U8292 (N_8292,N_6042,N_6757);
nand U8293 (N_8293,N_7352,N_7224);
or U8294 (N_8294,N_5359,N_6310);
xnor U8295 (N_8295,N_6899,N_5162);
xnor U8296 (N_8296,N_7488,N_6644);
nor U8297 (N_8297,N_5214,N_5593);
or U8298 (N_8298,N_6024,N_5517);
nor U8299 (N_8299,N_6887,N_6435);
or U8300 (N_8300,N_5991,N_6535);
and U8301 (N_8301,N_6673,N_6615);
or U8302 (N_8302,N_5744,N_6715);
xnor U8303 (N_8303,N_6750,N_7097);
xnor U8304 (N_8304,N_5766,N_5495);
xnor U8305 (N_8305,N_6763,N_5776);
nand U8306 (N_8306,N_5347,N_7359);
xor U8307 (N_8307,N_5536,N_6011);
nor U8308 (N_8308,N_6471,N_5096);
or U8309 (N_8309,N_5239,N_5903);
or U8310 (N_8310,N_5183,N_7060);
nand U8311 (N_8311,N_5623,N_6767);
xnor U8312 (N_8312,N_6313,N_7257);
nand U8313 (N_8313,N_5798,N_6208);
or U8314 (N_8314,N_7050,N_7358);
xor U8315 (N_8315,N_7223,N_6520);
and U8316 (N_8316,N_6696,N_6743);
xor U8317 (N_8317,N_6294,N_5062);
xor U8318 (N_8318,N_6904,N_6639);
or U8319 (N_8319,N_7092,N_5349);
and U8320 (N_8320,N_6185,N_6108);
nand U8321 (N_8321,N_5910,N_5489);
xor U8322 (N_8322,N_6479,N_6039);
nor U8323 (N_8323,N_7291,N_5176);
nand U8324 (N_8324,N_5510,N_6618);
or U8325 (N_8325,N_6466,N_6863);
or U8326 (N_8326,N_6149,N_6037);
nor U8327 (N_8327,N_6377,N_6503);
xnor U8328 (N_8328,N_6876,N_7101);
or U8329 (N_8329,N_6741,N_5785);
and U8330 (N_8330,N_7409,N_6356);
and U8331 (N_8331,N_5202,N_6330);
nand U8332 (N_8332,N_5361,N_5464);
and U8333 (N_8333,N_5637,N_5814);
nor U8334 (N_8334,N_5444,N_5066);
and U8335 (N_8335,N_6727,N_6272);
or U8336 (N_8336,N_6158,N_5345);
or U8337 (N_8337,N_6677,N_5467);
and U8338 (N_8338,N_6245,N_6489);
nand U8339 (N_8339,N_5933,N_7134);
nor U8340 (N_8340,N_5400,N_7251);
nor U8341 (N_8341,N_6617,N_5428);
nand U8342 (N_8342,N_5795,N_6177);
xor U8343 (N_8343,N_5492,N_6804);
or U8344 (N_8344,N_6248,N_5453);
nand U8345 (N_8345,N_6226,N_7020);
nor U8346 (N_8346,N_7485,N_5297);
nor U8347 (N_8347,N_5475,N_7330);
or U8348 (N_8348,N_5082,N_6145);
and U8349 (N_8349,N_6759,N_5172);
or U8350 (N_8350,N_6162,N_6854);
xor U8351 (N_8351,N_6418,N_5732);
nor U8352 (N_8352,N_6808,N_6060);
nand U8353 (N_8353,N_6835,N_5930);
nand U8354 (N_8354,N_5590,N_5780);
and U8355 (N_8355,N_5648,N_5687);
and U8356 (N_8356,N_5555,N_5286);
or U8357 (N_8357,N_7282,N_6907);
or U8358 (N_8358,N_6769,N_7045);
and U8359 (N_8359,N_6155,N_5221);
nand U8360 (N_8360,N_5630,N_5830);
and U8361 (N_8361,N_6881,N_6490);
or U8362 (N_8362,N_6323,N_7462);
nand U8363 (N_8363,N_6935,N_5628);
or U8364 (N_8364,N_5488,N_6223);
xnor U8365 (N_8365,N_6355,N_6922);
nor U8366 (N_8366,N_6691,N_5707);
nand U8367 (N_8367,N_6036,N_5708);
nor U8368 (N_8368,N_5002,N_5366);
nand U8369 (N_8369,N_7403,N_7445);
xor U8370 (N_8370,N_6421,N_6292);
or U8371 (N_8371,N_6972,N_5073);
nand U8372 (N_8372,N_6828,N_6096);
nand U8373 (N_8373,N_5515,N_6528);
nor U8374 (N_8374,N_6022,N_5271);
and U8375 (N_8375,N_5974,N_5548);
nor U8376 (N_8376,N_6939,N_6128);
and U8377 (N_8377,N_7156,N_7449);
and U8378 (N_8378,N_5698,N_5794);
nand U8379 (N_8379,N_5967,N_7154);
and U8380 (N_8380,N_5240,N_6200);
xor U8381 (N_8381,N_5786,N_7499);
and U8382 (N_8382,N_5321,N_7331);
or U8383 (N_8383,N_6262,N_6351);
or U8384 (N_8384,N_5658,N_6760);
nand U8385 (N_8385,N_5224,N_5948);
or U8386 (N_8386,N_7144,N_5604);
or U8387 (N_8387,N_6431,N_7307);
and U8388 (N_8388,N_5832,N_5601);
and U8389 (N_8389,N_5929,N_5320);
and U8390 (N_8390,N_6536,N_6856);
nand U8391 (N_8391,N_6650,N_5012);
and U8392 (N_8392,N_5318,N_5888);
nor U8393 (N_8393,N_5890,N_6288);
nor U8394 (N_8394,N_6668,N_6707);
or U8395 (N_8395,N_5573,N_5647);
nor U8396 (N_8396,N_5429,N_6724);
xnor U8397 (N_8397,N_5720,N_6140);
and U8398 (N_8398,N_5643,N_6794);
nand U8399 (N_8399,N_5142,N_5253);
and U8400 (N_8400,N_6118,N_5496);
and U8401 (N_8401,N_6369,N_6187);
xor U8402 (N_8402,N_7280,N_6002);
or U8403 (N_8403,N_6633,N_5419);
or U8404 (N_8404,N_7435,N_5706);
nand U8405 (N_8405,N_5724,N_5201);
nor U8406 (N_8406,N_5263,N_6072);
and U8407 (N_8407,N_6933,N_6184);
nand U8408 (N_8408,N_7458,N_5742);
and U8409 (N_8409,N_7036,N_6713);
and U8410 (N_8410,N_6051,N_5389);
nand U8411 (N_8411,N_6564,N_5578);
xnor U8412 (N_8412,N_5148,N_5788);
and U8413 (N_8413,N_5293,N_6401);
nand U8414 (N_8414,N_7473,N_6705);
nor U8415 (N_8415,N_6787,N_6805);
nand U8416 (N_8416,N_6962,N_5529);
and U8417 (N_8417,N_6921,N_5377);
nand U8418 (N_8418,N_5524,N_7274);
xnor U8419 (N_8419,N_6815,N_6178);
and U8420 (N_8420,N_5478,N_7028);
nor U8421 (N_8421,N_7182,N_6397);
or U8422 (N_8422,N_7109,N_5026);
nor U8423 (N_8423,N_6425,N_5982);
xnor U8424 (N_8424,N_5461,N_7453);
nor U8425 (N_8425,N_6832,N_6944);
nand U8426 (N_8426,N_6846,N_7203);
or U8427 (N_8427,N_5738,N_7081);
or U8428 (N_8428,N_6841,N_6859);
nand U8429 (N_8429,N_5468,N_6988);
xor U8430 (N_8430,N_5346,N_6762);
nand U8431 (N_8431,N_6176,N_5506);
and U8432 (N_8432,N_7123,N_6764);
or U8433 (N_8433,N_6225,N_5729);
or U8434 (N_8434,N_6665,N_6359);
nand U8435 (N_8435,N_5684,N_7258);
or U8436 (N_8436,N_5922,N_7277);
xor U8437 (N_8437,N_7405,N_5121);
xor U8438 (N_8438,N_6452,N_7024);
xor U8439 (N_8439,N_7419,N_7302);
xnor U8440 (N_8440,N_6920,N_7348);
nor U8441 (N_8441,N_6378,N_5925);
nor U8442 (N_8442,N_7418,N_7139);
nor U8443 (N_8443,N_5694,N_5731);
xor U8444 (N_8444,N_5639,N_5280);
xor U8445 (N_8445,N_5094,N_5173);
nor U8446 (N_8446,N_5577,N_5739);
xor U8447 (N_8447,N_6667,N_5417);
nand U8448 (N_8448,N_5328,N_5222);
nand U8449 (N_8449,N_7477,N_6388);
xor U8450 (N_8450,N_6890,N_6483);
or U8451 (N_8451,N_6870,N_6889);
nor U8452 (N_8452,N_6873,N_6557);
nand U8453 (N_8453,N_6608,N_7178);
and U8454 (N_8454,N_5063,N_6733);
nand U8455 (N_8455,N_6579,N_5943);
xor U8456 (N_8456,N_5737,N_6570);
nand U8457 (N_8457,N_7201,N_7113);
nor U8458 (N_8458,N_5713,N_6978);
and U8459 (N_8459,N_7073,N_6445);
xnor U8460 (N_8460,N_6164,N_6474);
nand U8461 (N_8461,N_6901,N_7069);
or U8462 (N_8462,N_6188,N_6751);
or U8463 (N_8463,N_6371,N_5340);
nand U8464 (N_8464,N_5041,N_5962);
nor U8465 (N_8465,N_5146,N_5207);
nand U8466 (N_8466,N_6701,N_5458);
or U8467 (N_8467,N_6508,N_5863);
and U8468 (N_8468,N_5645,N_5139);
or U8469 (N_8469,N_7099,N_5175);
or U8470 (N_8470,N_6470,N_7328);
and U8471 (N_8471,N_6941,N_5704);
and U8472 (N_8472,N_6662,N_6221);
nand U8473 (N_8473,N_7383,N_6892);
xnor U8474 (N_8474,N_5237,N_6148);
or U8475 (N_8475,N_6809,N_6362);
and U8476 (N_8476,N_6698,N_5260);
or U8477 (N_8477,N_7240,N_6432);
nor U8478 (N_8478,N_7181,N_5919);
nor U8479 (N_8479,N_6337,N_7265);
xnor U8480 (N_8480,N_5799,N_6104);
or U8481 (N_8481,N_5083,N_5746);
nand U8482 (N_8482,N_6722,N_6726);
and U8483 (N_8483,N_7215,N_6486);
and U8484 (N_8484,N_7235,N_7424);
nand U8485 (N_8485,N_6862,N_5819);
and U8486 (N_8486,N_5204,N_6626);
nor U8487 (N_8487,N_5408,N_7093);
nor U8488 (N_8488,N_5220,N_6970);
nor U8489 (N_8489,N_5711,N_5992);
nand U8490 (N_8490,N_6666,N_6695);
nor U8491 (N_8491,N_5288,N_6073);
xor U8492 (N_8492,N_5823,N_5251);
and U8493 (N_8493,N_7121,N_6681);
or U8494 (N_8494,N_7304,N_7431);
or U8495 (N_8495,N_5113,N_6032);
and U8496 (N_8496,N_5003,N_5950);
xor U8497 (N_8497,N_6531,N_7319);
or U8498 (N_8498,N_5486,N_7472);
xnor U8499 (N_8499,N_6840,N_6481);
or U8500 (N_8500,N_6179,N_7300);
nand U8501 (N_8501,N_5531,N_7160);
xnor U8502 (N_8502,N_6126,N_6839);
nand U8503 (N_8503,N_7141,N_5442);
nor U8504 (N_8504,N_6651,N_5691);
xor U8505 (N_8505,N_7313,N_5218);
nand U8506 (N_8506,N_6488,N_6084);
xnor U8507 (N_8507,N_6747,N_5099);
nor U8508 (N_8508,N_6442,N_5287);
or U8509 (N_8509,N_6339,N_7119);
nand U8510 (N_8510,N_6412,N_5805);
xnor U8511 (N_8511,N_7344,N_5043);
nor U8512 (N_8512,N_5425,N_6635);
xnor U8513 (N_8513,N_6229,N_7341);
nand U8514 (N_8514,N_5131,N_7107);
nand U8515 (N_8515,N_5392,N_6091);
and U8516 (N_8516,N_6976,N_7395);
nand U8517 (N_8517,N_7176,N_6365);
or U8518 (N_8518,N_5937,N_5124);
nand U8519 (N_8519,N_7094,N_6684);
xor U8520 (N_8520,N_5518,N_7083);
nand U8521 (N_8521,N_5426,N_5817);
xnor U8522 (N_8522,N_6372,N_6250);
and U8523 (N_8523,N_5120,N_6789);
xor U8524 (N_8524,N_5375,N_7143);
or U8525 (N_8525,N_5152,N_5127);
and U8526 (N_8526,N_7088,N_7471);
or U8527 (N_8527,N_6025,N_6408);
xnor U8528 (N_8528,N_6312,N_5363);
xnor U8529 (N_8529,N_7111,N_6061);
nand U8530 (N_8530,N_5861,N_7432);
xor U8531 (N_8531,N_6289,N_6163);
xnor U8532 (N_8532,N_5258,N_6585);
or U8533 (N_8533,N_5901,N_6080);
and U8534 (N_8534,N_6420,N_7246);
nor U8535 (N_8535,N_6575,N_5638);
nand U8536 (N_8536,N_5236,N_7047);
xor U8537 (N_8537,N_5261,N_6387);
nor U8538 (N_8538,N_6583,N_6461);
xor U8539 (N_8539,N_7219,N_5364);
nand U8540 (N_8540,N_5926,N_7338);
xnor U8541 (N_8541,N_7072,N_5964);
and U8542 (N_8542,N_6984,N_5612);
nor U8543 (N_8543,N_5013,N_5491);
xnor U8544 (N_8544,N_6410,N_5277);
nor U8545 (N_8545,N_6524,N_5360);
or U8546 (N_8546,N_7118,N_6565);
nor U8547 (N_8547,N_6516,N_5056);
nor U8548 (N_8548,N_5324,N_6343);
and U8549 (N_8549,N_5818,N_7112);
nand U8550 (N_8550,N_6168,N_5547);
nand U8551 (N_8551,N_5008,N_6894);
nand U8552 (N_8552,N_7259,N_6467);
nand U8553 (N_8553,N_7151,N_7152);
and U8554 (N_8554,N_6326,N_6720);
nor U8555 (N_8555,N_5315,N_5526);
nand U8556 (N_8556,N_5528,N_6327);
xnor U8557 (N_8557,N_6784,N_5159);
or U8558 (N_8558,N_6620,N_6414);
nand U8559 (N_8559,N_6201,N_6444);
or U8560 (N_8560,N_5931,N_5559);
and U8561 (N_8561,N_5957,N_5843);
nor U8562 (N_8562,N_6860,N_5174);
xnor U8563 (N_8563,N_6423,N_5503);
xor U8564 (N_8564,N_7189,N_6877);
nor U8565 (N_8565,N_5695,N_5944);
xnor U8566 (N_8566,N_6883,N_5068);
nor U8567 (N_8567,N_6123,N_5533);
nand U8568 (N_8568,N_6238,N_6702);
or U8569 (N_8569,N_5824,N_5833);
nand U8570 (N_8570,N_6068,N_6706);
and U8571 (N_8571,N_6756,N_5797);
and U8572 (N_8572,N_6058,N_5563);
nor U8573 (N_8573,N_5454,N_5145);
xor U8574 (N_8574,N_5245,N_5686);
and U8575 (N_8575,N_6419,N_5568);
nand U8576 (N_8576,N_5721,N_5485);
and U8577 (N_8577,N_6298,N_5430);
and U8578 (N_8578,N_7275,N_6019);
xnor U8579 (N_8579,N_5447,N_5150);
nand U8580 (N_8580,N_5040,N_5414);
and U8581 (N_8581,N_5996,N_5839);
nand U8582 (N_8582,N_5908,N_7305);
and U8583 (N_8583,N_6305,N_6232);
nor U8584 (N_8584,N_5988,N_6115);
and U8585 (N_8585,N_6102,N_7273);
or U8586 (N_8586,N_5635,N_6364);
nand U8587 (N_8587,N_7261,N_5609);
xnor U8588 (N_8588,N_5337,N_6354);
and U8589 (N_8589,N_7312,N_6672);
and U8590 (N_8590,N_7306,N_6888);
and U8591 (N_8591,N_7297,N_6830);
nand U8592 (N_8592,N_5323,N_5966);
and U8593 (N_8593,N_6704,N_6824);
xor U8594 (N_8594,N_6119,N_7239);
or U8595 (N_8595,N_6893,N_7454);
nand U8596 (N_8596,N_6311,N_6274);
and U8597 (N_8597,N_5034,N_7388);
or U8598 (N_8598,N_6302,N_6645);
nand U8599 (N_8599,N_6083,N_6353);
xnor U8600 (N_8600,N_6999,N_6599);
or U8601 (N_8601,N_6279,N_6237);
nand U8602 (N_8602,N_6283,N_5191);
xor U8603 (N_8603,N_6605,N_6853);
nand U8604 (N_8604,N_6469,N_5640);
nor U8605 (N_8605,N_7013,N_6742);
xnor U8606 (N_8606,N_5917,N_6744);
nor U8607 (N_8607,N_7474,N_5644);
and U8608 (N_8608,N_5714,N_7433);
nand U8609 (N_8609,N_5557,N_5482);
nor U8610 (N_8610,N_5369,N_7389);
or U8611 (N_8611,N_6041,N_7375);
or U8612 (N_8612,N_5091,N_5469);
or U8613 (N_8613,N_6345,N_6253);
xor U8614 (N_8614,N_7138,N_6857);
nor U8615 (N_8615,N_5129,N_6059);
nor U8616 (N_8616,N_6074,N_7032);
or U8617 (N_8617,N_6936,N_6173);
nor U8618 (N_8618,N_6513,N_5702);
xnor U8619 (N_8619,N_7187,N_5681);
or U8620 (N_8620,N_6228,N_7233);
xor U8621 (N_8621,N_7480,N_6156);
or U8622 (N_8622,N_7492,N_6634);
nand U8623 (N_8623,N_6694,N_6273);
or U8624 (N_8624,N_6686,N_7002);
nand U8625 (N_8625,N_5574,N_6034);
or U8626 (N_8626,N_5984,N_5803);
nand U8627 (N_8627,N_5076,N_5457);
or U8628 (N_8628,N_5998,N_6069);
or U8629 (N_8629,N_7104,N_7402);
or U8630 (N_8630,N_6373,N_7384);
or U8631 (N_8631,N_6247,N_7269);
and U8632 (N_8632,N_6940,N_6540);
or U8633 (N_8633,N_5231,N_6231);
and U8634 (N_8634,N_6249,N_7209);
or U8635 (N_8635,N_7440,N_5921);
xnor U8636 (N_8636,N_5862,N_7390);
nand U8637 (N_8637,N_6837,N_6438);
nor U8638 (N_8638,N_6753,N_6961);
and U8639 (N_8639,N_7262,N_5090);
xor U8640 (N_8640,N_6394,N_5763);
or U8641 (N_8641,N_6758,N_6455);
nor U8642 (N_8642,N_5332,N_6576);
or U8643 (N_8643,N_5164,N_6908);
nor U8644 (N_8644,N_5285,N_6594);
xor U8645 (N_8645,N_5620,N_7408);
or U8646 (N_8646,N_6627,N_6192);
nor U8647 (N_8647,N_6947,N_7374);
xor U8648 (N_8648,N_6275,N_5971);
nor U8649 (N_8649,N_7422,N_7349);
and U8650 (N_8650,N_5018,N_5481);
or U8651 (N_8651,N_5409,N_5816);
nand U8652 (N_8652,N_5942,N_7327);
and U8653 (N_8653,N_5849,N_6871);
nand U8654 (N_8654,N_5061,N_7363);
or U8655 (N_8655,N_5789,N_7056);
or U8656 (N_8656,N_5959,N_6572);
nor U8657 (N_8657,N_6768,N_7199);
and U8658 (N_8658,N_6318,N_7333);
nand U8659 (N_8659,N_5762,N_6246);
nor U8660 (N_8660,N_6937,N_7158);
nand U8661 (N_8661,N_6009,N_7074);
xor U8662 (N_8662,N_7218,N_5350);
or U8663 (N_8663,N_7498,N_5576);
nor U8664 (N_8664,N_6400,N_6424);
xor U8665 (N_8665,N_6052,N_6563);
and U8666 (N_8666,N_7354,N_6329);
nor U8667 (N_8667,N_6578,N_6646);
or U8668 (N_8668,N_5144,N_5829);
or U8669 (N_8669,N_5885,N_5415);
xor U8670 (N_8670,N_7042,N_5421);
or U8671 (N_8671,N_5295,N_5190);
xor U8672 (N_8672,N_7016,N_7145);
and U8673 (N_8673,N_5793,N_5924);
nand U8674 (N_8674,N_7230,N_5951);
nand U8675 (N_8675,N_5267,N_6786);
nor U8676 (N_8676,N_6596,N_6959);
nor U8677 (N_8677,N_6529,N_6902);
nand U8678 (N_8678,N_5160,N_6106);
xnor U8679 (N_8679,N_5370,N_6670);
nand U8680 (N_8680,N_5778,N_5270);
nand U8681 (N_8681,N_5085,N_5692);
and U8682 (N_8682,N_6437,N_6568);
and U8683 (N_8683,N_5525,N_7253);
nand U8684 (N_8684,N_7495,N_5668);
nor U8685 (N_8685,N_6879,N_6098);
xor U8686 (N_8686,N_6213,N_5608);
nor U8687 (N_8687,N_5761,N_7434);
and U8688 (N_8688,N_6336,N_7289);
nand U8689 (N_8689,N_5985,N_6501);
xor U8690 (N_8690,N_7213,N_5670);
or U8691 (N_8691,N_6909,N_7037);
nand U8692 (N_8692,N_5666,N_6105);
or U8693 (N_8693,N_6718,N_6683);
xor U8694 (N_8694,N_5460,N_6413);
xnor U8695 (N_8695,N_7413,N_5841);
nor U8696 (N_8696,N_5502,N_7231);
and U8697 (N_8697,N_5072,N_7426);
xnor U8698 (N_8698,N_7496,N_6679);
nor U8699 (N_8699,N_5020,N_5916);
xnor U8700 (N_8700,N_5017,N_6079);
nand U8701 (N_8701,N_5856,N_5784);
xnor U8702 (N_8702,N_6259,N_7371);
nor U8703 (N_8703,N_5588,N_6266);
and U8704 (N_8704,N_7493,N_6949);
nor U8705 (N_8705,N_5889,N_5790);
or U8706 (N_8706,N_5226,N_6728);
nor U8707 (N_8707,N_6687,N_6447);
nand U8708 (N_8708,N_6282,N_7027);
and U8709 (N_8709,N_5872,N_6591);
nor U8710 (N_8710,N_5582,N_7459);
and U8711 (N_8711,N_7336,N_7284);
and U8712 (N_8712,N_5228,N_5452);
xor U8713 (N_8713,N_6923,N_6212);
and U8714 (N_8714,N_5186,N_6480);
nor U8715 (N_8715,N_6263,N_7263);
xor U8716 (N_8716,N_6088,N_7343);
nand U8717 (N_8717,N_6141,N_6281);
and U8718 (N_8718,N_5282,N_7254);
and U8719 (N_8719,N_7196,N_6499);
xor U8720 (N_8720,N_5367,N_5993);
xor U8721 (N_8721,N_5217,N_7334);
and U8722 (N_8722,N_5727,N_5660);
nand U8723 (N_8723,N_5472,N_5519);
nand U8724 (N_8724,N_6773,N_7202);
nand U8725 (N_8725,N_6973,N_5678);
nand U8726 (N_8726,N_6463,N_6346);
or U8727 (N_8727,N_5566,N_7117);
nand U8728 (N_8728,N_5900,N_7241);
nand U8729 (N_8729,N_7229,N_5664);
xnor U8730 (N_8730,N_6458,N_6076);
xnor U8731 (N_8731,N_6736,N_5868);
and U8732 (N_8732,N_7245,N_6206);
xor U8733 (N_8733,N_6217,N_6614);
nand U8734 (N_8734,N_5807,N_6655);
nor U8735 (N_8735,N_6980,N_6189);
nand U8736 (N_8736,N_7222,N_5177);
and U8737 (N_8737,N_7206,N_5887);
xor U8738 (N_8738,N_6802,N_6621);
xor U8739 (N_8739,N_5523,N_6567);
nand U8740 (N_8740,N_5075,N_5928);
xor U8741 (N_8741,N_5110,N_7064);
xnor U8742 (N_8742,N_5752,N_7095);
or U8743 (N_8743,N_6609,N_5554);
nand U8744 (N_8744,N_6943,N_6746);
nand U8745 (N_8745,N_5646,N_5480);
nor U8746 (N_8746,N_7365,N_5869);
xor U8747 (N_8747,N_6381,N_6541);
and U8748 (N_8748,N_6190,N_6495);
xnor U8749 (N_8749,N_5071,N_6931);
xor U8750 (N_8750,N_5379,N_5792);
nor U8751 (N_8751,N_6090,N_5155);
nor U8752 (N_8752,N_5491,N_6961);
nor U8753 (N_8753,N_6906,N_6986);
or U8754 (N_8754,N_7440,N_5566);
xnor U8755 (N_8755,N_5922,N_5683);
nand U8756 (N_8756,N_5650,N_5194);
or U8757 (N_8757,N_5071,N_6212);
nor U8758 (N_8758,N_6919,N_5144);
nor U8759 (N_8759,N_5173,N_6261);
xor U8760 (N_8760,N_6531,N_7469);
nand U8761 (N_8761,N_6441,N_7372);
nand U8762 (N_8762,N_6632,N_6569);
nand U8763 (N_8763,N_7175,N_6493);
xor U8764 (N_8764,N_7136,N_6404);
nor U8765 (N_8765,N_6324,N_7092);
nand U8766 (N_8766,N_6465,N_6162);
or U8767 (N_8767,N_7132,N_5805);
nor U8768 (N_8768,N_7273,N_5959);
nand U8769 (N_8769,N_5127,N_6036);
or U8770 (N_8770,N_5858,N_6505);
xnor U8771 (N_8771,N_7051,N_6294);
nor U8772 (N_8772,N_5643,N_6893);
or U8773 (N_8773,N_6754,N_6940);
nand U8774 (N_8774,N_7374,N_5308);
xor U8775 (N_8775,N_6097,N_6988);
and U8776 (N_8776,N_7060,N_7495);
or U8777 (N_8777,N_6483,N_6138);
nor U8778 (N_8778,N_6061,N_5696);
nor U8779 (N_8779,N_6641,N_6593);
xor U8780 (N_8780,N_6434,N_5373);
nand U8781 (N_8781,N_7417,N_7333);
xor U8782 (N_8782,N_6455,N_5440);
nor U8783 (N_8783,N_5697,N_6963);
nor U8784 (N_8784,N_5921,N_5089);
and U8785 (N_8785,N_7073,N_6703);
xnor U8786 (N_8786,N_5305,N_5569);
and U8787 (N_8787,N_7408,N_6550);
or U8788 (N_8788,N_7056,N_7341);
and U8789 (N_8789,N_6026,N_5314);
xor U8790 (N_8790,N_6034,N_5965);
xnor U8791 (N_8791,N_6979,N_7039);
or U8792 (N_8792,N_5317,N_7364);
and U8793 (N_8793,N_5607,N_6499);
xor U8794 (N_8794,N_6411,N_5013);
xnor U8795 (N_8795,N_7335,N_5401);
nand U8796 (N_8796,N_5436,N_5595);
nor U8797 (N_8797,N_6305,N_6055);
nand U8798 (N_8798,N_6307,N_5177);
and U8799 (N_8799,N_6333,N_5256);
xnor U8800 (N_8800,N_6529,N_5440);
nor U8801 (N_8801,N_5731,N_6631);
nor U8802 (N_8802,N_7028,N_6056);
nor U8803 (N_8803,N_5351,N_6804);
xor U8804 (N_8804,N_6501,N_5385);
nor U8805 (N_8805,N_5503,N_6302);
nand U8806 (N_8806,N_5846,N_7406);
xor U8807 (N_8807,N_5676,N_5254);
or U8808 (N_8808,N_7064,N_6356);
nand U8809 (N_8809,N_5303,N_5291);
nor U8810 (N_8810,N_5655,N_7161);
or U8811 (N_8811,N_6403,N_7085);
nor U8812 (N_8812,N_6138,N_5612);
or U8813 (N_8813,N_6674,N_6364);
or U8814 (N_8814,N_7107,N_5239);
and U8815 (N_8815,N_5731,N_6065);
nor U8816 (N_8816,N_7383,N_5354);
nor U8817 (N_8817,N_5850,N_5050);
nand U8818 (N_8818,N_6503,N_5190);
nand U8819 (N_8819,N_5733,N_6666);
xnor U8820 (N_8820,N_7192,N_6977);
and U8821 (N_8821,N_6372,N_7393);
and U8822 (N_8822,N_7413,N_6926);
nand U8823 (N_8823,N_6851,N_6276);
and U8824 (N_8824,N_7174,N_7152);
or U8825 (N_8825,N_5696,N_5996);
xnor U8826 (N_8826,N_5759,N_7498);
xnor U8827 (N_8827,N_5875,N_6132);
nor U8828 (N_8828,N_5234,N_6530);
and U8829 (N_8829,N_5164,N_5316);
nand U8830 (N_8830,N_5112,N_5057);
or U8831 (N_8831,N_5657,N_5633);
or U8832 (N_8832,N_5844,N_6448);
nand U8833 (N_8833,N_6695,N_5158);
or U8834 (N_8834,N_6664,N_6875);
xor U8835 (N_8835,N_6167,N_5979);
nand U8836 (N_8836,N_5271,N_6986);
or U8837 (N_8837,N_6449,N_7385);
or U8838 (N_8838,N_6688,N_5813);
or U8839 (N_8839,N_5782,N_6043);
xnor U8840 (N_8840,N_6136,N_7294);
and U8841 (N_8841,N_6898,N_6966);
nand U8842 (N_8842,N_6298,N_5974);
nand U8843 (N_8843,N_6283,N_6405);
nand U8844 (N_8844,N_6194,N_7111);
xnor U8845 (N_8845,N_6951,N_6210);
and U8846 (N_8846,N_6287,N_5021);
nand U8847 (N_8847,N_6192,N_5164);
nor U8848 (N_8848,N_6718,N_7335);
or U8849 (N_8849,N_5490,N_5562);
or U8850 (N_8850,N_6129,N_7314);
nor U8851 (N_8851,N_5315,N_6802);
or U8852 (N_8852,N_5249,N_5112);
and U8853 (N_8853,N_6773,N_5146);
nand U8854 (N_8854,N_5369,N_5456);
nand U8855 (N_8855,N_7221,N_5859);
nor U8856 (N_8856,N_6153,N_6006);
xnor U8857 (N_8857,N_6101,N_5309);
nor U8858 (N_8858,N_6927,N_6078);
and U8859 (N_8859,N_5773,N_6660);
xnor U8860 (N_8860,N_7338,N_5184);
nand U8861 (N_8861,N_5735,N_6391);
nand U8862 (N_8862,N_6889,N_6787);
nand U8863 (N_8863,N_5654,N_6511);
or U8864 (N_8864,N_5562,N_6803);
nor U8865 (N_8865,N_6365,N_7179);
or U8866 (N_8866,N_6492,N_5918);
nand U8867 (N_8867,N_6206,N_6641);
xnor U8868 (N_8868,N_5572,N_5920);
and U8869 (N_8869,N_6701,N_6632);
or U8870 (N_8870,N_6315,N_5136);
and U8871 (N_8871,N_6865,N_6077);
or U8872 (N_8872,N_6885,N_6228);
nand U8873 (N_8873,N_5254,N_5514);
nand U8874 (N_8874,N_7382,N_5483);
nor U8875 (N_8875,N_6978,N_6726);
nor U8876 (N_8876,N_5046,N_7293);
or U8877 (N_8877,N_6809,N_7311);
nor U8878 (N_8878,N_6735,N_7056);
and U8879 (N_8879,N_6321,N_7099);
xor U8880 (N_8880,N_5546,N_5670);
or U8881 (N_8881,N_5021,N_6626);
xor U8882 (N_8882,N_6311,N_6191);
or U8883 (N_8883,N_6530,N_5115);
and U8884 (N_8884,N_6490,N_7240);
nor U8885 (N_8885,N_5596,N_5939);
and U8886 (N_8886,N_5267,N_7093);
or U8887 (N_8887,N_5104,N_5215);
xor U8888 (N_8888,N_5962,N_7423);
nor U8889 (N_8889,N_6917,N_6359);
and U8890 (N_8890,N_5243,N_6129);
or U8891 (N_8891,N_6736,N_6948);
and U8892 (N_8892,N_5344,N_5890);
or U8893 (N_8893,N_5126,N_7404);
xnor U8894 (N_8894,N_6762,N_5753);
nand U8895 (N_8895,N_6608,N_5520);
nand U8896 (N_8896,N_6301,N_6843);
nand U8897 (N_8897,N_5814,N_6095);
nor U8898 (N_8898,N_5230,N_5298);
xnor U8899 (N_8899,N_7415,N_6744);
and U8900 (N_8900,N_6090,N_5655);
nand U8901 (N_8901,N_6802,N_7097);
nor U8902 (N_8902,N_6695,N_5430);
and U8903 (N_8903,N_5012,N_7303);
nand U8904 (N_8904,N_5257,N_5849);
or U8905 (N_8905,N_7273,N_6462);
xnor U8906 (N_8906,N_5668,N_5582);
and U8907 (N_8907,N_6083,N_6811);
or U8908 (N_8908,N_5614,N_5916);
or U8909 (N_8909,N_5671,N_6512);
nand U8910 (N_8910,N_5388,N_5242);
nand U8911 (N_8911,N_7377,N_5918);
or U8912 (N_8912,N_5298,N_6368);
nor U8913 (N_8913,N_5859,N_6519);
nand U8914 (N_8914,N_6563,N_6405);
nand U8915 (N_8915,N_6203,N_6587);
and U8916 (N_8916,N_7175,N_7055);
or U8917 (N_8917,N_6818,N_5585);
or U8918 (N_8918,N_7060,N_5233);
and U8919 (N_8919,N_5011,N_5618);
nand U8920 (N_8920,N_6195,N_6028);
or U8921 (N_8921,N_5960,N_6275);
xnor U8922 (N_8922,N_6023,N_5918);
nor U8923 (N_8923,N_6924,N_5589);
xor U8924 (N_8924,N_5235,N_5939);
or U8925 (N_8925,N_5068,N_6530);
nor U8926 (N_8926,N_6958,N_5378);
or U8927 (N_8927,N_6950,N_6489);
nand U8928 (N_8928,N_5764,N_5311);
nor U8929 (N_8929,N_5578,N_6342);
or U8930 (N_8930,N_5425,N_7463);
or U8931 (N_8931,N_6636,N_6866);
or U8932 (N_8932,N_6150,N_5451);
and U8933 (N_8933,N_5713,N_7169);
nor U8934 (N_8934,N_7362,N_6909);
and U8935 (N_8935,N_5917,N_7041);
xor U8936 (N_8936,N_6612,N_6099);
or U8937 (N_8937,N_5338,N_5034);
xnor U8938 (N_8938,N_5450,N_6235);
xnor U8939 (N_8939,N_7351,N_6587);
or U8940 (N_8940,N_7176,N_5160);
and U8941 (N_8941,N_7205,N_7259);
nand U8942 (N_8942,N_5475,N_5563);
nor U8943 (N_8943,N_6046,N_5793);
and U8944 (N_8944,N_6387,N_5807);
xor U8945 (N_8945,N_5811,N_6581);
xor U8946 (N_8946,N_5199,N_7030);
xnor U8947 (N_8947,N_7039,N_6205);
or U8948 (N_8948,N_6015,N_5354);
and U8949 (N_8949,N_5308,N_7263);
nor U8950 (N_8950,N_5634,N_7471);
xor U8951 (N_8951,N_7352,N_6808);
xnor U8952 (N_8952,N_6241,N_5655);
nor U8953 (N_8953,N_6484,N_7250);
nor U8954 (N_8954,N_5000,N_5258);
xor U8955 (N_8955,N_6259,N_5546);
xor U8956 (N_8956,N_6122,N_6296);
nand U8957 (N_8957,N_5573,N_7318);
nand U8958 (N_8958,N_5295,N_5079);
or U8959 (N_8959,N_5942,N_5695);
and U8960 (N_8960,N_7260,N_7481);
nand U8961 (N_8961,N_6898,N_7360);
and U8962 (N_8962,N_6098,N_6378);
xnor U8963 (N_8963,N_5882,N_7497);
xnor U8964 (N_8964,N_5385,N_7463);
or U8965 (N_8965,N_5342,N_6860);
xor U8966 (N_8966,N_5683,N_5004);
or U8967 (N_8967,N_6245,N_6542);
nand U8968 (N_8968,N_5956,N_6996);
xor U8969 (N_8969,N_5354,N_5056);
nor U8970 (N_8970,N_5151,N_5192);
and U8971 (N_8971,N_6602,N_6247);
and U8972 (N_8972,N_5005,N_5003);
and U8973 (N_8973,N_6511,N_5285);
nor U8974 (N_8974,N_7052,N_7269);
nor U8975 (N_8975,N_5675,N_5858);
or U8976 (N_8976,N_6847,N_6214);
or U8977 (N_8977,N_6282,N_6693);
or U8978 (N_8978,N_5239,N_5737);
nand U8979 (N_8979,N_5600,N_5188);
nand U8980 (N_8980,N_7298,N_6134);
and U8981 (N_8981,N_5908,N_6976);
xor U8982 (N_8982,N_5394,N_5018);
nand U8983 (N_8983,N_6197,N_5422);
and U8984 (N_8984,N_5060,N_7134);
or U8985 (N_8985,N_5877,N_7056);
and U8986 (N_8986,N_5009,N_6861);
and U8987 (N_8987,N_6886,N_6935);
nor U8988 (N_8988,N_7002,N_5610);
nor U8989 (N_8989,N_6893,N_5705);
xor U8990 (N_8990,N_6059,N_7371);
or U8991 (N_8991,N_5472,N_6140);
nand U8992 (N_8992,N_5557,N_6572);
and U8993 (N_8993,N_6991,N_5537);
nand U8994 (N_8994,N_7383,N_7285);
or U8995 (N_8995,N_6410,N_5336);
nand U8996 (N_8996,N_6133,N_5128);
nor U8997 (N_8997,N_5879,N_5362);
nor U8998 (N_8998,N_5066,N_6559);
nor U8999 (N_8999,N_6259,N_6153);
nor U9000 (N_9000,N_5099,N_7316);
and U9001 (N_9001,N_5565,N_6713);
xor U9002 (N_9002,N_7132,N_6281);
or U9003 (N_9003,N_6571,N_7083);
and U9004 (N_9004,N_5612,N_6663);
xnor U9005 (N_9005,N_7258,N_5264);
and U9006 (N_9006,N_5120,N_5824);
xnor U9007 (N_9007,N_6907,N_5105);
nand U9008 (N_9008,N_7023,N_6780);
xor U9009 (N_9009,N_7220,N_6434);
nand U9010 (N_9010,N_5661,N_5253);
and U9011 (N_9011,N_5804,N_5747);
or U9012 (N_9012,N_6129,N_6804);
and U9013 (N_9013,N_7062,N_5260);
and U9014 (N_9014,N_5083,N_7157);
xnor U9015 (N_9015,N_6904,N_6762);
nand U9016 (N_9016,N_5866,N_5331);
nand U9017 (N_9017,N_6323,N_6285);
nand U9018 (N_9018,N_6162,N_5655);
xnor U9019 (N_9019,N_5252,N_5546);
xnor U9020 (N_9020,N_5123,N_6352);
xnor U9021 (N_9021,N_7073,N_6731);
xor U9022 (N_9022,N_6062,N_7414);
nor U9023 (N_9023,N_5316,N_5489);
nand U9024 (N_9024,N_6536,N_6929);
nand U9025 (N_9025,N_5362,N_5222);
and U9026 (N_9026,N_5095,N_7110);
or U9027 (N_9027,N_5971,N_6209);
and U9028 (N_9028,N_6728,N_6883);
or U9029 (N_9029,N_7180,N_6807);
xor U9030 (N_9030,N_7346,N_7277);
and U9031 (N_9031,N_5912,N_5510);
or U9032 (N_9032,N_5180,N_7217);
or U9033 (N_9033,N_5872,N_6646);
nand U9034 (N_9034,N_5595,N_6207);
nor U9035 (N_9035,N_5032,N_5478);
xor U9036 (N_9036,N_6559,N_7405);
and U9037 (N_9037,N_7232,N_7129);
nand U9038 (N_9038,N_6741,N_7282);
or U9039 (N_9039,N_5203,N_6696);
xor U9040 (N_9040,N_5277,N_5331);
and U9041 (N_9041,N_6106,N_6282);
xnor U9042 (N_9042,N_6885,N_7397);
nor U9043 (N_9043,N_5902,N_5387);
xnor U9044 (N_9044,N_6093,N_5703);
nor U9045 (N_9045,N_5048,N_5522);
xnor U9046 (N_9046,N_6045,N_6831);
and U9047 (N_9047,N_6280,N_7056);
xnor U9048 (N_9048,N_6580,N_5020);
nor U9049 (N_9049,N_6983,N_5022);
nor U9050 (N_9050,N_6606,N_5123);
nand U9051 (N_9051,N_7364,N_5599);
nor U9052 (N_9052,N_6130,N_7044);
xnor U9053 (N_9053,N_5565,N_5122);
nor U9054 (N_9054,N_6973,N_5247);
xnor U9055 (N_9055,N_5888,N_5089);
xnor U9056 (N_9056,N_5827,N_6490);
or U9057 (N_9057,N_6842,N_7338);
and U9058 (N_9058,N_6982,N_7457);
xnor U9059 (N_9059,N_5776,N_5581);
and U9060 (N_9060,N_6480,N_7477);
nand U9061 (N_9061,N_7043,N_5862);
xor U9062 (N_9062,N_6443,N_6291);
or U9063 (N_9063,N_6855,N_6044);
nand U9064 (N_9064,N_5345,N_5243);
or U9065 (N_9065,N_5560,N_7377);
xnor U9066 (N_9066,N_6738,N_7070);
or U9067 (N_9067,N_7356,N_6688);
nor U9068 (N_9068,N_6189,N_5873);
nor U9069 (N_9069,N_5447,N_6338);
nand U9070 (N_9070,N_5973,N_5021);
and U9071 (N_9071,N_7499,N_5841);
nand U9072 (N_9072,N_6602,N_6955);
or U9073 (N_9073,N_6868,N_7285);
nand U9074 (N_9074,N_6958,N_6725);
xnor U9075 (N_9075,N_5900,N_6664);
and U9076 (N_9076,N_6728,N_6006);
nor U9077 (N_9077,N_7093,N_7054);
nand U9078 (N_9078,N_6745,N_6574);
or U9079 (N_9079,N_6228,N_6193);
nor U9080 (N_9080,N_5785,N_6452);
nand U9081 (N_9081,N_6554,N_7320);
and U9082 (N_9082,N_6611,N_5711);
nor U9083 (N_9083,N_6447,N_6315);
or U9084 (N_9084,N_7348,N_6376);
or U9085 (N_9085,N_5878,N_6882);
and U9086 (N_9086,N_7069,N_6863);
xnor U9087 (N_9087,N_7310,N_6552);
nand U9088 (N_9088,N_6780,N_6897);
xor U9089 (N_9089,N_7421,N_6610);
nor U9090 (N_9090,N_5547,N_6485);
xnor U9091 (N_9091,N_6706,N_5146);
xor U9092 (N_9092,N_6883,N_6398);
nor U9093 (N_9093,N_6908,N_7170);
xnor U9094 (N_9094,N_5607,N_5996);
nand U9095 (N_9095,N_6656,N_5978);
nand U9096 (N_9096,N_5763,N_6828);
and U9097 (N_9097,N_5931,N_6933);
nand U9098 (N_9098,N_7426,N_5817);
or U9099 (N_9099,N_5056,N_6385);
nand U9100 (N_9100,N_6042,N_5984);
and U9101 (N_9101,N_6805,N_5313);
xor U9102 (N_9102,N_6388,N_5620);
nor U9103 (N_9103,N_5114,N_6512);
nor U9104 (N_9104,N_6506,N_5076);
and U9105 (N_9105,N_5339,N_5747);
nand U9106 (N_9106,N_5481,N_7302);
nor U9107 (N_9107,N_7086,N_6737);
nand U9108 (N_9108,N_6830,N_6297);
or U9109 (N_9109,N_5541,N_6507);
or U9110 (N_9110,N_6752,N_6239);
nor U9111 (N_9111,N_6196,N_6923);
xor U9112 (N_9112,N_5741,N_5241);
xnor U9113 (N_9113,N_6403,N_5962);
nor U9114 (N_9114,N_5607,N_6341);
and U9115 (N_9115,N_7196,N_7416);
nand U9116 (N_9116,N_7475,N_7398);
nand U9117 (N_9117,N_5928,N_5666);
or U9118 (N_9118,N_7013,N_6791);
or U9119 (N_9119,N_6957,N_5470);
xnor U9120 (N_9120,N_7402,N_7274);
and U9121 (N_9121,N_6310,N_5896);
nor U9122 (N_9122,N_5203,N_7251);
nand U9123 (N_9123,N_5312,N_7017);
or U9124 (N_9124,N_6005,N_6717);
nand U9125 (N_9125,N_7360,N_7378);
and U9126 (N_9126,N_7353,N_7251);
nor U9127 (N_9127,N_7479,N_6918);
or U9128 (N_9128,N_6341,N_5301);
nor U9129 (N_9129,N_6817,N_7390);
xnor U9130 (N_9130,N_6782,N_7346);
nor U9131 (N_9131,N_5186,N_6229);
nor U9132 (N_9132,N_5376,N_5632);
xor U9133 (N_9133,N_6129,N_5410);
nand U9134 (N_9134,N_5084,N_6766);
and U9135 (N_9135,N_6384,N_7435);
or U9136 (N_9136,N_5260,N_6149);
and U9137 (N_9137,N_5011,N_6870);
xor U9138 (N_9138,N_6631,N_5352);
and U9139 (N_9139,N_5645,N_5227);
nor U9140 (N_9140,N_5417,N_5227);
nor U9141 (N_9141,N_6196,N_5971);
xnor U9142 (N_9142,N_6245,N_5231);
nand U9143 (N_9143,N_6869,N_6013);
nand U9144 (N_9144,N_5061,N_5957);
and U9145 (N_9145,N_5911,N_5644);
and U9146 (N_9146,N_5315,N_7269);
or U9147 (N_9147,N_6632,N_5855);
nand U9148 (N_9148,N_5767,N_5195);
xor U9149 (N_9149,N_7423,N_6300);
nand U9150 (N_9150,N_6343,N_7383);
and U9151 (N_9151,N_6502,N_5542);
nand U9152 (N_9152,N_5229,N_5183);
nand U9153 (N_9153,N_5596,N_6416);
and U9154 (N_9154,N_7463,N_7188);
nand U9155 (N_9155,N_5247,N_5732);
and U9156 (N_9156,N_5492,N_6325);
xor U9157 (N_9157,N_6337,N_5007);
and U9158 (N_9158,N_6523,N_6169);
or U9159 (N_9159,N_7248,N_5910);
and U9160 (N_9160,N_6605,N_7205);
and U9161 (N_9161,N_6951,N_5679);
and U9162 (N_9162,N_5685,N_7413);
and U9163 (N_9163,N_6075,N_6117);
xor U9164 (N_9164,N_5925,N_6728);
nand U9165 (N_9165,N_5560,N_6917);
nor U9166 (N_9166,N_6411,N_5821);
and U9167 (N_9167,N_7021,N_5025);
or U9168 (N_9168,N_5423,N_6407);
nor U9169 (N_9169,N_5410,N_5239);
nor U9170 (N_9170,N_5582,N_5311);
or U9171 (N_9171,N_6016,N_5129);
nor U9172 (N_9172,N_6732,N_5757);
nor U9173 (N_9173,N_6387,N_7259);
or U9174 (N_9174,N_5687,N_6404);
or U9175 (N_9175,N_6480,N_5971);
nor U9176 (N_9176,N_6785,N_5085);
nor U9177 (N_9177,N_6705,N_6341);
nand U9178 (N_9178,N_5627,N_6358);
xor U9179 (N_9179,N_5796,N_6474);
nor U9180 (N_9180,N_5317,N_6541);
nor U9181 (N_9181,N_7347,N_7211);
xnor U9182 (N_9182,N_7108,N_5568);
xor U9183 (N_9183,N_5999,N_5859);
nand U9184 (N_9184,N_5096,N_5477);
xnor U9185 (N_9185,N_5211,N_7044);
and U9186 (N_9186,N_5156,N_7285);
and U9187 (N_9187,N_6432,N_5600);
and U9188 (N_9188,N_5694,N_7083);
xnor U9189 (N_9189,N_6460,N_5793);
xnor U9190 (N_9190,N_6144,N_7045);
xnor U9191 (N_9191,N_5018,N_6884);
xnor U9192 (N_9192,N_6166,N_7086);
xnor U9193 (N_9193,N_6732,N_6136);
nand U9194 (N_9194,N_5758,N_7224);
or U9195 (N_9195,N_7448,N_6826);
or U9196 (N_9196,N_5526,N_5312);
nor U9197 (N_9197,N_6732,N_5803);
or U9198 (N_9198,N_5846,N_6404);
or U9199 (N_9199,N_6755,N_5879);
and U9200 (N_9200,N_6948,N_6312);
and U9201 (N_9201,N_7155,N_5072);
nor U9202 (N_9202,N_5270,N_5094);
xnor U9203 (N_9203,N_6745,N_6436);
nand U9204 (N_9204,N_7055,N_6058);
and U9205 (N_9205,N_6642,N_5054);
nor U9206 (N_9206,N_6164,N_5748);
nor U9207 (N_9207,N_6739,N_6990);
xnor U9208 (N_9208,N_5431,N_6337);
xnor U9209 (N_9209,N_6635,N_7275);
xnor U9210 (N_9210,N_7252,N_7212);
nor U9211 (N_9211,N_5665,N_6409);
and U9212 (N_9212,N_6057,N_5634);
xor U9213 (N_9213,N_6046,N_7401);
and U9214 (N_9214,N_5763,N_7120);
or U9215 (N_9215,N_5831,N_5188);
nor U9216 (N_9216,N_7285,N_5147);
or U9217 (N_9217,N_6788,N_6666);
nand U9218 (N_9218,N_7341,N_5617);
nand U9219 (N_9219,N_5096,N_5677);
nand U9220 (N_9220,N_5512,N_6099);
nand U9221 (N_9221,N_6453,N_7374);
nand U9222 (N_9222,N_6685,N_6923);
nand U9223 (N_9223,N_5295,N_6057);
nor U9224 (N_9224,N_6220,N_6314);
and U9225 (N_9225,N_7319,N_5732);
nand U9226 (N_9226,N_5236,N_6093);
or U9227 (N_9227,N_6620,N_6225);
xor U9228 (N_9228,N_5356,N_5166);
and U9229 (N_9229,N_5337,N_7442);
nor U9230 (N_9230,N_5630,N_6284);
xnor U9231 (N_9231,N_5316,N_7241);
xor U9232 (N_9232,N_5194,N_6683);
nor U9233 (N_9233,N_6099,N_5768);
xor U9234 (N_9234,N_6108,N_6820);
nand U9235 (N_9235,N_6164,N_6699);
nor U9236 (N_9236,N_6377,N_7338);
nand U9237 (N_9237,N_7417,N_6800);
nand U9238 (N_9238,N_6667,N_5037);
xnor U9239 (N_9239,N_6272,N_7424);
xor U9240 (N_9240,N_7033,N_5777);
xor U9241 (N_9241,N_6853,N_6361);
and U9242 (N_9242,N_7446,N_5612);
nor U9243 (N_9243,N_5178,N_6596);
or U9244 (N_9244,N_7065,N_6369);
nor U9245 (N_9245,N_6619,N_5406);
xor U9246 (N_9246,N_5220,N_5730);
and U9247 (N_9247,N_7325,N_5252);
or U9248 (N_9248,N_7343,N_6147);
or U9249 (N_9249,N_7085,N_6817);
xnor U9250 (N_9250,N_6743,N_6738);
xnor U9251 (N_9251,N_5641,N_6354);
nand U9252 (N_9252,N_7151,N_5147);
xor U9253 (N_9253,N_7491,N_6428);
and U9254 (N_9254,N_5297,N_5083);
and U9255 (N_9255,N_6262,N_6253);
xnor U9256 (N_9256,N_6361,N_5497);
or U9257 (N_9257,N_5815,N_7378);
nor U9258 (N_9258,N_5744,N_5112);
xnor U9259 (N_9259,N_7328,N_7094);
and U9260 (N_9260,N_5679,N_6659);
nor U9261 (N_9261,N_6530,N_5247);
or U9262 (N_9262,N_6051,N_7021);
or U9263 (N_9263,N_7483,N_5335);
nor U9264 (N_9264,N_6769,N_5270);
or U9265 (N_9265,N_5898,N_6657);
and U9266 (N_9266,N_5378,N_6026);
xnor U9267 (N_9267,N_6940,N_6637);
xnor U9268 (N_9268,N_5258,N_7125);
xor U9269 (N_9269,N_5676,N_5287);
and U9270 (N_9270,N_5642,N_7490);
or U9271 (N_9271,N_6377,N_5248);
or U9272 (N_9272,N_6540,N_7044);
xor U9273 (N_9273,N_6906,N_5256);
nor U9274 (N_9274,N_5800,N_6345);
nor U9275 (N_9275,N_7102,N_7209);
and U9276 (N_9276,N_7176,N_6416);
and U9277 (N_9277,N_6218,N_6981);
or U9278 (N_9278,N_5413,N_7232);
and U9279 (N_9279,N_6370,N_7109);
or U9280 (N_9280,N_6855,N_5317);
nor U9281 (N_9281,N_5215,N_5535);
nand U9282 (N_9282,N_5512,N_6764);
nor U9283 (N_9283,N_7288,N_5188);
and U9284 (N_9284,N_7415,N_5517);
or U9285 (N_9285,N_5234,N_5295);
nand U9286 (N_9286,N_5777,N_5601);
or U9287 (N_9287,N_5804,N_7046);
nand U9288 (N_9288,N_5016,N_7294);
or U9289 (N_9289,N_6845,N_5560);
or U9290 (N_9290,N_6330,N_7441);
and U9291 (N_9291,N_6936,N_7077);
nor U9292 (N_9292,N_5869,N_6402);
and U9293 (N_9293,N_6822,N_6564);
or U9294 (N_9294,N_5298,N_7477);
xnor U9295 (N_9295,N_5488,N_6656);
xnor U9296 (N_9296,N_5792,N_5207);
nor U9297 (N_9297,N_6253,N_5017);
or U9298 (N_9298,N_7420,N_6914);
xnor U9299 (N_9299,N_5032,N_5944);
nor U9300 (N_9300,N_6653,N_6460);
and U9301 (N_9301,N_7097,N_5097);
nor U9302 (N_9302,N_7039,N_6912);
xnor U9303 (N_9303,N_6222,N_7086);
xnor U9304 (N_9304,N_6901,N_6124);
nor U9305 (N_9305,N_6662,N_6004);
and U9306 (N_9306,N_6442,N_5981);
or U9307 (N_9307,N_6815,N_6619);
or U9308 (N_9308,N_7113,N_5921);
or U9309 (N_9309,N_6681,N_6347);
xor U9310 (N_9310,N_5402,N_6439);
and U9311 (N_9311,N_5828,N_6000);
or U9312 (N_9312,N_7196,N_6345);
or U9313 (N_9313,N_5178,N_6779);
nand U9314 (N_9314,N_5601,N_5110);
or U9315 (N_9315,N_6482,N_5724);
or U9316 (N_9316,N_6075,N_6041);
nor U9317 (N_9317,N_7440,N_7127);
or U9318 (N_9318,N_5403,N_7450);
or U9319 (N_9319,N_6871,N_6925);
nor U9320 (N_9320,N_6290,N_6333);
nand U9321 (N_9321,N_6161,N_5263);
nor U9322 (N_9322,N_5606,N_6641);
nand U9323 (N_9323,N_6966,N_5539);
nor U9324 (N_9324,N_7230,N_7436);
or U9325 (N_9325,N_5355,N_5827);
or U9326 (N_9326,N_7192,N_5590);
nand U9327 (N_9327,N_5586,N_7429);
nor U9328 (N_9328,N_5412,N_7161);
or U9329 (N_9329,N_5248,N_6119);
nor U9330 (N_9330,N_6996,N_6763);
nor U9331 (N_9331,N_6716,N_6326);
xor U9332 (N_9332,N_5139,N_5894);
and U9333 (N_9333,N_6438,N_6611);
xnor U9334 (N_9334,N_6577,N_6844);
nor U9335 (N_9335,N_6616,N_5151);
xnor U9336 (N_9336,N_5375,N_6334);
nand U9337 (N_9337,N_7404,N_5114);
and U9338 (N_9338,N_5830,N_7228);
nand U9339 (N_9339,N_5730,N_5193);
nor U9340 (N_9340,N_5255,N_5149);
nand U9341 (N_9341,N_5155,N_6832);
nor U9342 (N_9342,N_6531,N_7339);
xor U9343 (N_9343,N_5533,N_7320);
xor U9344 (N_9344,N_6633,N_5745);
xor U9345 (N_9345,N_6673,N_6090);
nand U9346 (N_9346,N_6600,N_5578);
nand U9347 (N_9347,N_5848,N_5491);
and U9348 (N_9348,N_7322,N_5215);
and U9349 (N_9349,N_5300,N_7238);
xnor U9350 (N_9350,N_5265,N_5097);
xor U9351 (N_9351,N_7437,N_5905);
nand U9352 (N_9352,N_5266,N_7281);
xnor U9353 (N_9353,N_7075,N_5921);
or U9354 (N_9354,N_6544,N_6968);
xor U9355 (N_9355,N_5107,N_7419);
and U9356 (N_9356,N_7236,N_5388);
nand U9357 (N_9357,N_6979,N_7413);
nand U9358 (N_9358,N_6474,N_6435);
and U9359 (N_9359,N_7097,N_5047);
and U9360 (N_9360,N_5572,N_6421);
and U9361 (N_9361,N_5146,N_5625);
nand U9362 (N_9362,N_6199,N_5043);
xnor U9363 (N_9363,N_5140,N_6974);
nand U9364 (N_9364,N_6675,N_6958);
nor U9365 (N_9365,N_5645,N_5501);
xor U9366 (N_9366,N_5489,N_5084);
xnor U9367 (N_9367,N_6669,N_5318);
or U9368 (N_9368,N_7300,N_6040);
and U9369 (N_9369,N_7075,N_6705);
or U9370 (N_9370,N_5106,N_5711);
or U9371 (N_9371,N_7075,N_6273);
xnor U9372 (N_9372,N_5696,N_5416);
xnor U9373 (N_9373,N_5973,N_6747);
and U9374 (N_9374,N_6649,N_5525);
nand U9375 (N_9375,N_7392,N_6632);
nor U9376 (N_9376,N_6926,N_7253);
and U9377 (N_9377,N_6552,N_5761);
and U9378 (N_9378,N_5766,N_7356);
nand U9379 (N_9379,N_5834,N_6075);
nor U9380 (N_9380,N_6758,N_6385);
nor U9381 (N_9381,N_6800,N_6154);
nor U9382 (N_9382,N_7039,N_6610);
nand U9383 (N_9383,N_7464,N_6603);
nand U9384 (N_9384,N_5474,N_6614);
nand U9385 (N_9385,N_6952,N_6137);
nand U9386 (N_9386,N_7098,N_5088);
and U9387 (N_9387,N_5355,N_6795);
or U9388 (N_9388,N_7317,N_6693);
or U9389 (N_9389,N_5198,N_5345);
nand U9390 (N_9390,N_5030,N_5719);
or U9391 (N_9391,N_6721,N_6414);
xor U9392 (N_9392,N_6263,N_6225);
and U9393 (N_9393,N_7052,N_5159);
xnor U9394 (N_9394,N_5140,N_5577);
nand U9395 (N_9395,N_5086,N_7362);
or U9396 (N_9396,N_6242,N_6237);
xor U9397 (N_9397,N_5161,N_5577);
nand U9398 (N_9398,N_7287,N_5355);
or U9399 (N_9399,N_5840,N_7383);
nor U9400 (N_9400,N_6931,N_6211);
xnor U9401 (N_9401,N_5164,N_5930);
xor U9402 (N_9402,N_5631,N_5291);
xnor U9403 (N_9403,N_5893,N_6722);
and U9404 (N_9404,N_7319,N_5808);
and U9405 (N_9405,N_5518,N_7069);
xnor U9406 (N_9406,N_6686,N_5309);
or U9407 (N_9407,N_6372,N_6571);
nand U9408 (N_9408,N_6004,N_5676);
nand U9409 (N_9409,N_6418,N_6332);
and U9410 (N_9410,N_6843,N_6479);
and U9411 (N_9411,N_7327,N_6290);
nand U9412 (N_9412,N_5202,N_6395);
nand U9413 (N_9413,N_5533,N_6517);
nand U9414 (N_9414,N_5327,N_7471);
and U9415 (N_9415,N_6697,N_6999);
or U9416 (N_9416,N_6645,N_6903);
nand U9417 (N_9417,N_6306,N_6761);
or U9418 (N_9418,N_6922,N_5020);
and U9419 (N_9419,N_6966,N_5232);
or U9420 (N_9420,N_6201,N_5236);
or U9421 (N_9421,N_5890,N_5154);
xor U9422 (N_9422,N_7093,N_5957);
or U9423 (N_9423,N_6083,N_6961);
nand U9424 (N_9424,N_5281,N_6249);
nand U9425 (N_9425,N_6867,N_6790);
and U9426 (N_9426,N_5051,N_6687);
and U9427 (N_9427,N_5976,N_5052);
xnor U9428 (N_9428,N_6143,N_5208);
nor U9429 (N_9429,N_6430,N_5864);
nand U9430 (N_9430,N_5871,N_7265);
nor U9431 (N_9431,N_5864,N_6135);
nor U9432 (N_9432,N_6447,N_7451);
nor U9433 (N_9433,N_7427,N_6999);
xnor U9434 (N_9434,N_6884,N_5505);
or U9435 (N_9435,N_5673,N_5084);
nand U9436 (N_9436,N_7385,N_5121);
xnor U9437 (N_9437,N_5963,N_6028);
or U9438 (N_9438,N_6086,N_5952);
or U9439 (N_9439,N_5212,N_7136);
xor U9440 (N_9440,N_5772,N_5702);
nor U9441 (N_9441,N_7203,N_5243);
or U9442 (N_9442,N_6556,N_5035);
nand U9443 (N_9443,N_6246,N_5168);
xnor U9444 (N_9444,N_7007,N_6855);
nor U9445 (N_9445,N_5083,N_6322);
nor U9446 (N_9446,N_5123,N_7224);
or U9447 (N_9447,N_7398,N_6874);
nor U9448 (N_9448,N_7093,N_5865);
nor U9449 (N_9449,N_7028,N_5124);
or U9450 (N_9450,N_6384,N_5376);
or U9451 (N_9451,N_5308,N_6098);
and U9452 (N_9452,N_5219,N_6606);
nand U9453 (N_9453,N_7150,N_5038);
nand U9454 (N_9454,N_5104,N_6484);
and U9455 (N_9455,N_6605,N_6901);
or U9456 (N_9456,N_5487,N_5735);
xor U9457 (N_9457,N_6726,N_6504);
or U9458 (N_9458,N_6209,N_5451);
nor U9459 (N_9459,N_5566,N_6984);
and U9460 (N_9460,N_7129,N_7239);
and U9461 (N_9461,N_5650,N_5250);
nor U9462 (N_9462,N_6689,N_5088);
xor U9463 (N_9463,N_5778,N_5558);
and U9464 (N_9464,N_7029,N_7314);
nand U9465 (N_9465,N_7011,N_5132);
xnor U9466 (N_9466,N_6061,N_6137);
or U9467 (N_9467,N_5690,N_6901);
or U9468 (N_9468,N_6211,N_5948);
nand U9469 (N_9469,N_5568,N_6861);
nor U9470 (N_9470,N_7081,N_5310);
nor U9471 (N_9471,N_7431,N_7189);
and U9472 (N_9472,N_6949,N_5997);
nand U9473 (N_9473,N_7272,N_6075);
xnor U9474 (N_9474,N_5928,N_6114);
nor U9475 (N_9475,N_7474,N_7112);
nor U9476 (N_9476,N_7421,N_5413);
xnor U9477 (N_9477,N_6262,N_5340);
xor U9478 (N_9478,N_6655,N_7142);
xor U9479 (N_9479,N_6547,N_6434);
nand U9480 (N_9480,N_5394,N_7413);
xor U9481 (N_9481,N_6575,N_6729);
nand U9482 (N_9482,N_5530,N_5017);
or U9483 (N_9483,N_5988,N_5906);
nand U9484 (N_9484,N_6970,N_6011);
or U9485 (N_9485,N_6106,N_5472);
nor U9486 (N_9486,N_5304,N_7258);
and U9487 (N_9487,N_6260,N_7040);
nand U9488 (N_9488,N_7226,N_5273);
or U9489 (N_9489,N_5552,N_5107);
or U9490 (N_9490,N_5964,N_5459);
nor U9491 (N_9491,N_5730,N_7462);
nand U9492 (N_9492,N_5906,N_6733);
and U9493 (N_9493,N_7413,N_7050);
nor U9494 (N_9494,N_5786,N_5390);
nor U9495 (N_9495,N_6859,N_5563);
or U9496 (N_9496,N_6627,N_6542);
nand U9497 (N_9497,N_5692,N_6441);
nand U9498 (N_9498,N_5712,N_6986);
nand U9499 (N_9499,N_6701,N_5069);
xor U9500 (N_9500,N_7475,N_6821);
or U9501 (N_9501,N_6103,N_5581);
nand U9502 (N_9502,N_6545,N_6707);
nor U9503 (N_9503,N_5000,N_5104);
nor U9504 (N_9504,N_7426,N_6653);
nand U9505 (N_9505,N_7279,N_7369);
nand U9506 (N_9506,N_6717,N_5213);
xor U9507 (N_9507,N_7302,N_6963);
nand U9508 (N_9508,N_7232,N_6555);
xor U9509 (N_9509,N_5103,N_5894);
xor U9510 (N_9510,N_7427,N_6895);
xor U9511 (N_9511,N_6941,N_6541);
and U9512 (N_9512,N_7208,N_5390);
nand U9513 (N_9513,N_6747,N_5811);
xor U9514 (N_9514,N_6870,N_5720);
nor U9515 (N_9515,N_5908,N_7428);
and U9516 (N_9516,N_6625,N_5042);
xnor U9517 (N_9517,N_6966,N_5168);
or U9518 (N_9518,N_5661,N_6047);
or U9519 (N_9519,N_5282,N_6404);
nand U9520 (N_9520,N_5398,N_6689);
or U9521 (N_9521,N_6833,N_5348);
or U9522 (N_9522,N_5342,N_7440);
or U9523 (N_9523,N_5882,N_5960);
and U9524 (N_9524,N_6712,N_7389);
nand U9525 (N_9525,N_6620,N_6795);
and U9526 (N_9526,N_7406,N_5969);
xor U9527 (N_9527,N_6620,N_6918);
nor U9528 (N_9528,N_7461,N_6493);
nor U9529 (N_9529,N_5531,N_6357);
nand U9530 (N_9530,N_6853,N_5447);
xnor U9531 (N_9531,N_5597,N_6369);
nor U9532 (N_9532,N_5805,N_7212);
or U9533 (N_9533,N_5180,N_6702);
and U9534 (N_9534,N_7114,N_7487);
xor U9535 (N_9535,N_7368,N_7054);
and U9536 (N_9536,N_6445,N_6861);
xnor U9537 (N_9537,N_7411,N_5662);
xor U9538 (N_9538,N_6773,N_5814);
nand U9539 (N_9539,N_6114,N_5628);
or U9540 (N_9540,N_5281,N_5042);
nor U9541 (N_9541,N_6596,N_5622);
xnor U9542 (N_9542,N_6932,N_6980);
or U9543 (N_9543,N_6721,N_5145);
or U9544 (N_9544,N_7170,N_5441);
xnor U9545 (N_9545,N_6328,N_6622);
xor U9546 (N_9546,N_5999,N_7464);
nor U9547 (N_9547,N_5239,N_5054);
xor U9548 (N_9548,N_5494,N_5208);
and U9549 (N_9549,N_7298,N_5229);
nor U9550 (N_9550,N_6294,N_6181);
and U9551 (N_9551,N_6285,N_7079);
nand U9552 (N_9552,N_5718,N_7209);
nor U9553 (N_9553,N_6891,N_7100);
nor U9554 (N_9554,N_5693,N_5438);
nor U9555 (N_9555,N_6463,N_7088);
and U9556 (N_9556,N_7433,N_5153);
nor U9557 (N_9557,N_5560,N_6004);
xor U9558 (N_9558,N_6488,N_5461);
or U9559 (N_9559,N_7460,N_7016);
and U9560 (N_9560,N_5429,N_5734);
nor U9561 (N_9561,N_5864,N_5603);
xor U9562 (N_9562,N_5848,N_6996);
xor U9563 (N_9563,N_5856,N_7461);
nor U9564 (N_9564,N_5281,N_6772);
or U9565 (N_9565,N_7086,N_7382);
and U9566 (N_9566,N_6371,N_5505);
nor U9567 (N_9567,N_6575,N_6362);
nor U9568 (N_9568,N_6248,N_6529);
and U9569 (N_9569,N_6964,N_6027);
nor U9570 (N_9570,N_7357,N_6483);
or U9571 (N_9571,N_6741,N_6202);
or U9572 (N_9572,N_5426,N_5098);
nor U9573 (N_9573,N_6921,N_5230);
or U9574 (N_9574,N_5853,N_5742);
nor U9575 (N_9575,N_6470,N_5028);
nand U9576 (N_9576,N_7159,N_5233);
and U9577 (N_9577,N_6495,N_7045);
nand U9578 (N_9578,N_6487,N_6873);
and U9579 (N_9579,N_5333,N_5406);
and U9580 (N_9580,N_6309,N_5137);
nor U9581 (N_9581,N_6218,N_6023);
and U9582 (N_9582,N_6249,N_6425);
and U9583 (N_9583,N_5274,N_6206);
xnor U9584 (N_9584,N_6621,N_6816);
xnor U9585 (N_9585,N_6094,N_7263);
nand U9586 (N_9586,N_5545,N_5912);
and U9587 (N_9587,N_7066,N_6718);
xor U9588 (N_9588,N_6207,N_6309);
and U9589 (N_9589,N_6360,N_6810);
xor U9590 (N_9590,N_5817,N_6797);
nand U9591 (N_9591,N_6447,N_5591);
or U9592 (N_9592,N_5133,N_7226);
nand U9593 (N_9593,N_5807,N_5704);
and U9594 (N_9594,N_7107,N_5414);
nand U9595 (N_9595,N_6430,N_5422);
or U9596 (N_9596,N_5511,N_7176);
or U9597 (N_9597,N_7256,N_7227);
and U9598 (N_9598,N_5162,N_5280);
nand U9599 (N_9599,N_7254,N_5700);
xnor U9600 (N_9600,N_5725,N_6310);
nand U9601 (N_9601,N_5511,N_7292);
nand U9602 (N_9602,N_6727,N_7365);
nor U9603 (N_9603,N_5688,N_7328);
nand U9604 (N_9604,N_6275,N_6855);
nand U9605 (N_9605,N_6244,N_5358);
nand U9606 (N_9606,N_7037,N_6649);
and U9607 (N_9607,N_6269,N_7021);
or U9608 (N_9608,N_7493,N_5656);
xor U9609 (N_9609,N_7284,N_5516);
nand U9610 (N_9610,N_7403,N_6052);
xnor U9611 (N_9611,N_6850,N_6176);
or U9612 (N_9612,N_6218,N_5208);
nor U9613 (N_9613,N_6970,N_5827);
nand U9614 (N_9614,N_5185,N_7474);
or U9615 (N_9615,N_7073,N_5570);
nor U9616 (N_9616,N_7290,N_7091);
nor U9617 (N_9617,N_6113,N_5488);
nor U9618 (N_9618,N_6428,N_6252);
or U9619 (N_9619,N_5980,N_6329);
and U9620 (N_9620,N_6079,N_6224);
or U9621 (N_9621,N_6698,N_6276);
nor U9622 (N_9622,N_7022,N_5407);
xnor U9623 (N_9623,N_7132,N_7373);
nand U9624 (N_9624,N_5009,N_5372);
nand U9625 (N_9625,N_5185,N_5133);
and U9626 (N_9626,N_6176,N_6091);
or U9627 (N_9627,N_5495,N_6067);
and U9628 (N_9628,N_6025,N_6454);
nand U9629 (N_9629,N_5970,N_5198);
and U9630 (N_9630,N_6919,N_6293);
xnor U9631 (N_9631,N_5592,N_6983);
or U9632 (N_9632,N_6078,N_7456);
or U9633 (N_9633,N_6747,N_6913);
or U9634 (N_9634,N_7435,N_6555);
xnor U9635 (N_9635,N_6529,N_6043);
nor U9636 (N_9636,N_5805,N_6893);
and U9637 (N_9637,N_5714,N_5496);
nand U9638 (N_9638,N_6943,N_7319);
nand U9639 (N_9639,N_5336,N_5347);
and U9640 (N_9640,N_5779,N_6836);
xor U9641 (N_9641,N_7193,N_5361);
nor U9642 (N_9642,N_6744,N_7000);
and U9643 (N_9643,N_5692,N_5353);
or U9644 (N_9644,N_5593,N_6536);
nand U9645 (N_9645,N_6395,N_6858);
and U9646 (N_9646,N_6369,N_6985);
nand U9647 (N_9647,N_6390,N_5163);
nor U9648 (N_9648,N_7053,N_6097);
nor U9649 (N_9649,N_5432,N_6588);
xnor U9650 (N_9650,N_5213,N_6423);
and U9651 (N_9651,N_5429,N_7111);
nor U9652 (N_9652,N_7383,N_6148);
or U9653 (N_9653,N_6143,N_7496);
or U9654 (N_9654,N_5354,N_5304);
nor U9655 (N_9655,N_6875,N_5980);
nand U9656 (N_9656,N_6359,N_5236);
or U9657 (N_9657,N_5602,N_6861);
or U9658 (N_9658,N_6980,N_5375);
nor U9659 (N_9659,N_6002,N_6377);
and U9660 (N_9660,N_7115,N_5412);
nand U9661 (N_9661,N_6562,N_6279);
xor U9662 (N_9662,N_7106,N_6468);
nand U9663 (N_9663,N_6197,N_6399);
or U9664 (N_9664,N_6715,N_5951);
nand U9665 (N_9665,N_5325,N_7233);
xor U9666 (N_9666,N_5959,N_5412);
xor U9667 (N_9667,N_5723,N_6064);
xnor U9668 (N_9668,N_6881,N_6805);
xor U9669 (N_9669,N_6525,N_5533);
and U9670 (N_9670,N_6760,N_7254);
nor U9671 (N_9671,N_6024,N_6901);
and U9672 (N_9672,N_6755,N_5526);
and U9673 (N_9673,N_5204,N_5539);
nor U9674 (N_9674,N_5855,N_5657);
xor U9675 (N_9675,N_6973,N_5910);
or U9676 (N_9676,N_7205,N_5258);
xnor U9677 (N_9677,N_6275,N_6535);
nor U9678 (N_9678,N_6677,N_7236);
and U9679 (N_9679,N_7427,N_5363);
or U9680 (N_9680,N_5901,N_6548);
nor U9681 (N_9681,N_6696,N_6270);
nor U9682 (N_9682,N_5951,N_7394);
or U9683 (N_9683,N_7388,N_5148);
nor U9684 (N_9684,N_5873,N_6997);
or U9685 (N_9685,N_6533,N_6640);
nor U9686 (N_9686,N_6918,N_5406);
nand U9687 (N_9687,N_6859,N_6394);
xnor U9688 (N_9688,N_6786,N_5787);
or U9689 (N_9689,N_5954,N_6080);
nand U9690 (N_9690,N_7342,N_5051);
nand U9691 (N_9691,N_7151,N_5283);
and U9692 (N_9692,N_5701,N_5168);
or U9693 (N_9693,N_6302,N_6750);
xor U9694 (N_9694,N_6472,N_5728);
nand U9695 (N_9695,N_6384,N_6390);
nand U9696 (N_9696,N_5776,N_6203);
nand U9697 (N_9697,N_5537,N_5366);
xor U9698 (N_9698,N_5545,N_5161);
nor U9699 (N_9699,N_5180,N_5763);
or U9700 (N_9700,N_6128,N_6796);
and U9701 (N_9701,N_5174,N_6987);
xor U9702 (N_9702,N_5223,N_5272);
xnor U9703 (N_9703,N_7122,N_5860);
and U9704 (N_9704,N_6670,N_5476);
nand U9705 (N_9705,N_6972,N_7399);
or U9706 (N_9706,N_5392,N_6408);
nor U9707 (N_9707,N_6022,N_5247);
xor U9708 (N_9708,N_5848,N_6559);
and U9709 (N_9709,N_5827,N_5872);
xor U9710 (N_9710,N_5750,N_7197);
xor U9711 (N_9711,N_6584,N_5403);
nand U9712 (N_9712,N_6402,N_7331);
or U9713 (N_9713,N_5292,N_5553);
nand U9714 (N_9714,N_5967,N_5064);
and U9715 (N_9715,N_6186,N_5752);
and U9716 (N_9716,N_5958,N_6517);
or U9717 (N_9717,N_7230,N_6331);
and U9718 (N_9718,N_7162,N_5262);
nor U9719 (N_9719,N_6487,N_6269);
or U9720 (N_9720,N_7225,N_5619);
nand U9721 (N_9721,N_6804,N_6193);
and U9722 (N_9722,N_6079,N_7185);
nand U9723 (N_9723,N_7258,N_5833);
or U9724 (N_9724,N_5656,N_5588);
nor U9725 (N_9725,N_7393,N_7246);
nand U9726 (N_9726,N_7254,N_6756);
and U9727 (N_9727,N_5369,N_7304);
xnor U9728 (N_9728,N_7272,N_7026);
and U9729 (N_9729,N_7226,N_6452);
nand U9730 (N_9730,N_5982,N_6297);
nor U9731 (N_9731,N_7002,N_5235);
nand U9732 (N_9732,N_5412,N_5427);
nor U9733 (N_9733,N_6261,N_5159);
nand U9734 (N_9734,N_7284,N_6366);
xnor U9735 (N_9735,N_6325,N_5127);
or U9736 (N_9736,N_5159,N_7436);
nor U9737 (N_9737,N_5504,N_6517);
and U9738 (N_9738,N_5831,N_6117);
nand U9739 (N_9739,N_5806,N_7138);
and U9740 (N_9740,N_7421,N_5231);
nand U9741 (N_9741,N_7281,N_6671);
or U9742 (N_9742,N_7223,N_5826);
xnor U9743 (N_9743,N_5294,N_6695);
or U9744 (N_9744,N_5779,N_5563);
or U9745 (N_9745,N_6697,N_6465);
nor U9746 (N_9746,N_6927,N_5601);
and U9747 (N_9747,N_7033,N_6911);
nor U9748 (N_9748,N_5946,N_5487);
xor U9749 (N_9749,N_7448,N_6401);
nand U9750 (N_9750,N_5842,N_6571);
xnor U9751 (N_9751,N_6380,N_7450);
and U9752 (N_9752,N_7173,N_6261);
and U9753 (N_9753,N_7085,N_6026);
nand U9754 (N_9754,N_7280,N_5834);
and U9755 (N_9755,N_6853,N_5927);
xor U9756 (N_9756,N_6452,N_6570);
xnor U9757 (N_9757,N_5832,N_5201);
and U9758 (N_9758,N_5356,N_5391);
xnor U9759 (N_9759,N_5739,N_5453);
or U9760 (N_9760,N_7189,N_6646);
nand U9761 (N_9761,N_5519,N_5275);
or U9762 (N_9762,N_6144,N_6702);
nand U9763 (N_9763,N_6379,N_6393);
and U9764 (N_9764,N_6142,N_7010);
and U9765 (N_9765,N_5577,N_6006);
and U9766 (N_9766,N_5159,N_6171);
or U9767 (N_9767,N_7364,N_7265);
or U9768 (N_9768,N_6920,N_5288);
and U9769 (N_9769,N_5737,N_5960);
and U9770 (N_9770,N_6507,N_5224);
nor U9771 (N_9771,N_5627,N_5491);
xnor U9772 (N_9772,N_6710,N_6533);
nor U9773 (N_9773,N_6856,N_5776);
and U9774 (N_9774,N_5084,N_5903);
and U9775 (N_9775,N_5780,N_6358);
and U9776 (N_9776,N_6997,N_5484);
xor U9777 (N_9777,N_5682,N_7011);
or U9778 (N_9778,N_6346,N_5711);
nand U9779 (N_9779,N_7139,N_6037);
and U9780 (N_9780,N_6034,N_5484);
nor U9781 (N_9781,N_5080,N_5620);
xnor U9782 (N_9782,N_6061,N_5152);
and U9783 (N_9783,N_5379,N_5702);
or U9784 (N_9784,N_5922,N_7188);
xor U9785 (N_9785,N_6915,N_5958);
or U9786 (N_9786,N_7284,N_5875);
xnor U9787 (N_9787,N_7494,N_6150);
nor U9788 (N_9788,N_5669,N_7190);
and U9789 (N_9789,N_5727,N_5255);
or U9790 (N_9790,N_5137,N_6422);
or U9791 (N_9791,N_5376,N_5085);
xor U9792 (N_9792,N_5682,N_5867);
nor U9793 (N_9793,N_5393,N_7020);
nand U9794 (N_9794,N_6007,N_7143);
xor U9795 (N_9795,N_6829,N_6969);
nor U9796 (N_9796,N_5242,N_5885);
nor U9797 (N_9797,N_5795,N_5254);
or U9798 (N_9798,N_6647,N_5461);
nand U9799 (N_9799,N_6254,N_6788);
nand U9800 (N_9800,N_5559,N_5584);
nor U9801 (N_9801,N_5510,N_5605);
xor U9802 (N_9802,N_5933,N_6715);
xnor U9803 (N_9803,N_7227,N_6805);
and U9804 (N_9804,N_5529,N_6728);
nor U9805 (N_9805,N_7236,N_7137);
or U9806 (N_9806,N_7321,N_5560);
and U9807 (N_9807,N_7484,N_5036);
xor U9808 (N_9808,N_5938,N_6835);
or U9809 (N_9809,N_6833,N_5055);
and U9810 (N_9810,N_5493,N_6415);
nand U9811 (N_9811,N_6966,N_6402);
nand U9812 (N_9812,N_6080,N_6334);
or U9813 (N_9813,N_6768,N_5767);
nand U9814 (N_9814,N_5053,N_5707);
xnor U9815 (N_9815,N_7092,N_6905);
and U9816 (N_9816,N_7425,N_7112);
nand U9817 (N_9817,N_5879,N_7300);
and U9818 (N_9818,N_6130,N_6968);
xor U9819 (N_9819,N_6548,N_7279);
or U9820 (N_9820,N_5908,N_6607);
or U9821 (N_9821,N_7294,N_5996);
nor U9822 (N_9822,N_7494,N_5081);
nand U9823 (N_9823,N_7084,N_7025);
nor U9824 (N_9824,N_7101,N_6810);
nor U9825 (N_9825,N_7339,N_7499);
nor U9826 (N_9826,N_7169,N_6112);
xnor U9827 (N_9827,N_7342,N_7415);
nand U9828 (N_9828,N_5005,N_6984);
and U9829 (N_9829,N_5228,N_6465);
nand U9830 (N_9830,N_6242,N_5917);
nor U9831 (N_9831,N_5912,N_6895);
xnor U9832 (N_9832,N_6351,N_7179);
nor U9833 (N_9833,N_5279,N_5858);
nand U9834 (N_9834,N_6583,N_5223);
nand U9835 (N_9835,N_5705,N_5881);
xor U9836 (N_9836,N_6172,N_5923);
or U9837 (N_9837,N_6077,N_6949);
nand U9838 (N_9838,N_6554,N_5267);
nand U9839 (N_9839,N_7117,N_5602);
nor U9840 (N_9840,N_6695,N_5843);
or U9841 (N_9841,N_6558,N_6900);
or U9842 (N_9842,N_6469,N_5221);
nor U9843 (N_9843,N_6461,N_6635);
xnor U9844 (N_9844,N_6289,N_5728);
and U9845 (N_9845,N_5062,N_6144);
or U9846 (N_9846,N_5755,N_5187);
nor U9847 (N_9847,N_6804,N_5146);
or U9848 (N_9848,N_5353,N_5953);
nor U9849 (N_9849,N_6365,N_5799);
xor U9850 (N_9850,N_5883,N_5555);
xnor U9851 (N_9851,N_7030,N_7293);
xnor U9852 (N_9852,N_6604,N_7165);
xor U9853 (N_9853,N_6445,N_7373);
nand U9854 (N_9854,N_6007,N_5017);
nand U9855 (N_9855,N_6882,N_6826);
nand U9856 (N_9856,N_6710,N_5550);
nand U9857 (N_9857,N_7034,N_6305);
and U9858 (N_9858,N_6459,N_5749);
nor U9859 (N_9859,N_6014,N_5565);
and U9860 (N_9860,N_6745,N_5286);
nand U9861 (N_9861,N_6422,N_5924);
or U9862 (N_9862,N_6714,N_6440);
or U9863 (N_9863,N_5358,N_6866);
nor U9864 (N_9864,N_5810,N_6944);
xor U9865 (N_9865,N_5510,N_6539);
xor U9866 (N_9866,N_7341,N_6983);
or U9867 (N_9867,N_6702,N_6673);
or U9868 (N_9868,N_5190,N_6677);
xor U9869 (N_9869,N_6685,N_5306);
nand U9870 (N_9870,N_5485,N_6845);
nand U9871 (N_9871,N_7215,N_7371);
and U9872 (N_9872,N_7398,N_5563);
xor U9873 (N_9873,N_7252,N_5856);
and U9874 (N_9874,N_5996,N_5173);
and U9875 (N_9875,N_6731,N_6056);
or U9876 (N_9876,N_6800,N_5497);
or U9877 (N_9877,N_6058,N_5569);
nor U9878 (N_9878,N_5524,N_7197);
nor U9879 (N_9879,N_6443,N_7110);
or U9880 (N_9880,N_5499,N_7410);
nor U9881 (N_9881,N_6338,N_6077);
xor U9882 (N_9882,N_5243,N_5671);
and U9883 (N_9883,N_7427,N_6946);
nand U9884 (N_9884,N_5870,N_5609);
nor U9885 (N_9885,N_7178,N_6053);
or U9886 (N_9886,N_6658,N_6675);
xnor U9887 (N_9887,N_6865,N_6939);
nand U9888 (N_9888,N_6455,N_5203);
and U9889 (N_9889,N_5642,N_6056);
or U9890 (N_9890,N_6540,N_7304);
nor U9891 (N_9891,N_7088,N_6925);
nor U9892 (N_9892,N_6250,N_6293);
nor U9893 (N_9893,N_5446,N_7236);
or U9894 (N_9894,N_6126,N_6038);
xnor U9895 (N_9895,N_5936,N_7011);
and U9896 (N_9896,N_7300,N_6488);
or U9897 (N_9897,N_6353,N_5773);
nand U9898 (N_9898,N_5381,N_6143);
xnor U9899 (N_9899,N_5496,N_5501);
and U9900 (N_9900,N_6407,N_6670);
nor U9901 (N_9901,N_6490,N_5552);
xnor U9902 (N_9902,N_6660,N_5033);
nor U9903 (N_9903,N_6004,N_6687);
and U9904 (N_9904,N_7250,N_6743);
nor U9905 (N_9905,N_5170,N_5896);
or U9906 (N_9906,N_6645,N_5129);
nor U9907 (N_9907,N_5903,N_6743);
and U9908 (N_9908,N_6017,N_5934);
and U9909 (N_9909,N_6251,N_5625);
and U9910 (N_9910,N_6791,N_6977);
and U9911 (N_9911,N_5506,N_6664);
xnor U9912 (N_9912,N_5167,N_5802);
nand U9913 (N_9913,N_7170,N_7219);
nor U9914 (N_9914,N_7047,N_5831);
nand U9915 (N_9915,N_5583,N_5798);
xnor U9916 (N_9916,N_7351,N_5175);
nor U9917 (N_9917,N_6704,N_5796);
nand U9918 (N_9918,N_5667,N_5856);
and U9919 (N_9919,N_6951,N_5319);
and U9920 (N_9920,N_6975,N_6764);
and U9921 (N_9921,N_7030,N_7409);
or U9922 (N_9922,N_6991,N_6090);
xnor U9923 (N_9923,N_5832,N_7031);
nand U9924 (N_9924,N_5263,N_5929);
nor U9925 (N_9925,N_6186,N_5201);
and U9926 (N_9926,N_7110,N_6223);
xnor U9927 (N_9927,N_5340,N_6515);
nand U9928 (N_9928,N_6321,N_6707);
nor U9929 (N_9929,N_6315,N_5657);
xor U9930 (N_9930,N_6601,N_6089);
and U9931 (N_9931,N_6718,N_5005);
and U9932 (N_9932,N_5169,N_6413);
nand U9933 (N_9933,N_5737,N_6342);
and U9934 (N_9934,N_6750,N_7196);
nor U9935 (N_9935,N_5278,N_5030);
or U9936 (N_9936,N_6135,N_6865);
xor U9937 (N_9937,N_5283,N_7494);
xor U9938 (N_9938,N_5081,N_7109);
or U9939 (N_9939,N_5154,N_7284);
and U9940 (N_9940,N_5877,N_5211);
nor U9941 (N_9941,N_6983,N_6110);
nor U9942 (N_9942,N_6411,N_5382);
and U9943 (N_9943,N_5118,N_5131);
nand U9944 (N_9944,N_5440,N_7175);
or U9945 (N_9945,N_6545,N_6638);
or U9946 (N_9946,N_5490,N_6267);
nand U9947 (N_9947,N_5324,N_7174);
xor U9948 (N_9948,N_6651,N_5401);
xnor U9949 (N_9949,N_6930,N_6656);
nor U9950 (N_9950,N_6736,N_6658);
xnor U9951 (N_9951,N_5847,N_5506);
and U9952 (N_9952,N_7453,N_6608);
xor U9953 (N_9953,N_5957,N_6298);
and U9954 (N_9954,N_7064,N_6616);
nor U9955 (N_9955,N_6420,N_6863);
nor U9956 (N_9956,N_5384,N_7431);
and U9957 (N_9957,N_5884,N_5895);
xnor U9958 (N_9958,N_5873,N_5641);
or U9959 (N_9959,N_5010,N_6977);
nor U9960 (N_9960,N_5652,N_5415);
nand U9961 (N_9961,N_6309,N_5837);
nand U9962 (N_9962,N_6645,N_6341);
xor U9963 (N_9963,N_7343,N_6065);
nor U9964 (N_9964,N_7189,N_6955);
xnor U9965 (N_9965,N_5583,N_6963);
or U9966 (N_9966,N_5440,N_5133);
nor U9967 (N_9967,N_5671,N_6218);
and U9968 (N_9968,N_7337,N_6306);
nand U9969 (N_9969,N_7379,N_6420);
xor U9970 (N_9970,N_6228,N_7328);
xnor U9971 (N_9971,N_6234,N_6487);
nor U9972 (N_9972,N_5285,N_6734);
nand U9973 (N_9973,N_5302,N_6697);
nand U9974 (N_9974,N_5605,N_5819);
and U9975 (N_9975,N_7039,N_7001);
or U9976 (N_9976,N_5399,N_6836);
xor U9977 (N_9977,N_6774,N_5371);
nand U9978 (N_9978,N_5485,N_6349);
nor U9979 (N_9979,N_6519,N_6499);
nand U9980 (N_9980,N_5679,N_5837);
nor U9981 (N_9981,N_7285,N_5052);
xor U9982 (N_9982,N_5768,N_5276);
xnor U9983 (N_9983,N_5689,N_7475);
and U9984 (N_9984,N_6773,N_6250);
nor U9985 (N_9985,N_6389,N_5925);
and U9986 (N_9986,N_6594,N_6926);
or U9987 (N_9987,N_5710,N_5372);
nand U9988 (N_9988,N_5548,N_5810);
nor U9989 (N_9989,N_5984,N_7183);
nor U9990 (N_9990,N_6972,N_6330);
or U9991 (N_9991,N_7054,N_7228);
nand U9992 (N_9992,N_6407,N_6769);
xnor U9993 (N_9993,N_5857,N_7126);
nor U9994 (N_9994,N_5803,N_6914);
xnor U9995 (N_9995,N_7328,N_6100);
nand U9996 (N_9996,N_6221,N_6564);
nand U9997 (N_9997,N_7117,N_6364);
xnor U9998 (N_9998,N_5741,N_7431);
nand U9999 (N_9999,N_5185,N_5202);
nand U10000 (N_10000,N_9514,N_8654);
xor U10001 (N_10001,N_9284,N_8561);
nor U10002 (N_10002,N_8788,N_9449);
nand U10003 (N_10003,N_9918,N_9207);
and U10004 (N_10004,N_8541,N_8142);
nand U10005 (N_10005,N_7771,N_9905);
nor U10006 (N_10006,N_8923,N_7561);
xnor U10007 (N_10007,N_9647,N_7872);
nor U10008 (N_10008,N_9108,N_7877);
nor U10009 (N_10009,N_8609,N_8872);
or U10010 (N_10010,N_7563,N_7927);
and U10011 (N_10011,N_8751,N_9990);
or U10012 (N_10012,N_8421,N_9664);
or U10013 (N_10013,N_8009,N_8667);
nand U10014 (N_10014,N_7728,N_8659);
or U10015 (N_10015,N_8570,N_9555);
and U10016 (N_10016,N_8909,N_7964);
xnor U10017 (N_10017,N_8286,N_8330);
nand U10018 (N_10018,N_9246,N_8798);
nand U10019 (N_10019,N_7693,N_9734);
nor U10020 (N_10020,N_8157,N_7880);
nor U10021 (N_10021,N_7914,N_9817);
or U10022 (N_10022,N_9690,N_8642);
and U10023 (N_10023,N_7580,N_9203);
or U10024 (N_10024,N_7671,N_8753);
nor U10025 (N_10025,N_9457,N_7641);
and U10026 (N_10026,N_9047,N_8450);
nand U10027 (N_10027,N_9065,N_8724);
and U10028 (N_10028,N_8956,N_8482);
or U10029 (N_10029,N_9319,N_7697);
nand U10030 (N_10030,N_8383,N_7604);
nand U10031 (N_10031,N_8817,N_9334);
nand U10032 (N_10032,N_7610,N_9491);
nor U10033 (N_10033,N_7962,N_9811);
xnor U10034 (N_10034,N_9854,N_7768);
xnor U10035 (N_10035,N_7669,N_8981);
nand U10036 (N_10036,N_9240,N_9086);
nand U10037 (N_10037,N_8579,N_9374);
xor U10038 (N_10038,N_8943,N_9581);
nor U10039 (N_10039,N_9949,N_8974);
and U10040 (N_10040,N_9845,N_7609);
or U10041 (N_10041,N_9658,N_9787);
nor U10042 (N_10042,N_8081,N_9216);
nand U10043 (N_10043,N_7786,N_9221);
nor U10044 (N_10044,N_9878,N_7706);
nand U10045 (N_10045,N_7852,N_8436);
xor U10046 (N_10046,N_8804,N_8007);
xor U10047 (N_10047,N_9760,N_8941);
and U10048 (N_10048,N_8344,N_9339);
and U10049 (N_10049,N_8374,N_8841);
and U10050 (N_10050,N_7614,N_8422);
nor U10051 (N_10051,N_8822,N_9999);
and U10052 (N_10052,N_9104,N_9718);
nand U10053 (N_10053,N_8765,N_8268);
and U10054 (N_10054,N_9473,N_9834);
and U10055 (N_10055,N_7874,N_8021);
nand U10056 (N_10056,N_9421,N_9842);
and U10057 (N_10057,N_8229,N_9723);
or U10058 (N_10058,N_9039,N_7683);
xnor U10059 (N_10059,N_8054,N_9631);
nor U10060 (N_10060,N_8707,N_9963);
nor U10061 (N_10061,N_9518,N_9267);
xnor U10062 (N_10062,N_8401,N_9759);
nor U10063 (N_10063,N_8996,N_9057);
nand U10064 (N_10064,N_9560,N_7982);
and U10065 (N_10065,N_8891,N_9448);
xnor U10066 (N_10066,N_9646,N_8321);
and U10067 (N_10067,N_7865,N_9184);
nor U10068 (N_10068,N_9495,N_8039);
xor U10069 (N_10069,N_8773,N_9579);
nand U10070 (N_10070,N_7732,N_7546);
or U10071 (N_10071,N_8698,N_9719);
xor U10072 (N_10072,N_7856,N_9685);
and U10073 (N_10073,N_9347,N_8380);
or U10074 (N_10074,N_8827,N_8256);
xnor U10075 (N_10075,N_9067,N_9577);
and U10076 (N_10076,N_8961,N_7835);
nand U10077 (N_10077,N_7719,N_9767);
nand U10078 (N_10078,N_9937,N_8816);
xnor U10079 (N_10079,N_9014,N_8492);
nand U10080 (N_10080,N_8682,N_9798);
or U10081 (N_10081,N_8728,N_8070);
nand U10082 (N_10082,N_8060,N_9400);
xnor U10083 (N_10083,N_8523,N_8594);
nand U10084 (N_10084,N_8819,N_9135);
nand U10085 (N_10085,N_9125,N_8525);
nor U10086 (N_10086,N_7616,N_9800);
nand U10087 (N_10087,N_9528,N_8219);
or U10088 (N_10088,N_8631,N_8017);
and U10089 (N_10089,N_8145,N_7884);
and U10090 (N_10090,N_9433,N_9585);
nand U10091 (N_10091,N_7944,N_7508);
or U10092 (N_10092,N_7938,N_9792);
nor U10093 (N_10093,N_8494,N_8702);
nand U10094 (N_10094,N_9853,N_8351);
xor U10095 (N_10095,N_9124,N_8512);
nor U10096 (N_10096,N_8314,N_8663);
nor U10097 (N_10097,N_7581,N_8040);
xor U10098 (N_10098,N_8430,N_8411);
and U10099 (N_10099,N_8184,N_7654);
xnor U10100 (N_10100,N_8989,N_8115);
or U10101 (N_10101,N_9253,N_8409);
or U10102 (N_10102,N_7650,N_8098);
nand U10103 (N_10103,N_9139,N_9586);
and U10104 (N_10104,N_9945,N_8095);
and U10105 (N_10105,N_8225,N_8825);
xnor U10106 (N_10106,N_8621,N_7704);
and U10107 (N_10107,N_9699,N_9230);
and U10108 (N_10108,N_9464,N_8024);
nor U10109 (N_10109,N_9417,N_7537);
nand U10110 (N_10110,N_7777,N_9188);
nand U10111 (N_10111,N_8993,N_8417);
or U10112 (N_10112,N_9475,N_7824);
and U10113 (N_10113,N_8213,N_7784);
or U10114 (N_10114,N_9262,N_9698);
or U10115 (N_10115,N_9331,N_8927);
xor U10116 (N_10116,N_8437,N_8121);
nor U10117 (N_10117,N_9046,N_8498);
nand U10118 (N_10118,N_7565,N_8965);
and U10119 (N_10119,N_8771,N_9741);
and U10120 (N_10120,N_7709,N_9915);
or U10121 (N_10121,N_7668,N_8537);
xor U10122 (N_10122,N_9265,N_9415);
or U10123 (N_10123,N_9282,N_8141);
and U10124 (N_10124,N_8487,N_8510);
or U10125 (N_10125,N_7603,N_7601);
and U10126 (N_10126,N_8776,N_8182);
xor U10127 (N_10127,N_8801,N_9471);
and U10128 (N_10128,N_9485,N_8265);
nor U10129 (N_10129,N_9439,N_9494);
and U10130 (N_10130,N_8435,N_8163);
or U10131 (N_10131,N_9481,N_9438);
and U10132 (N_10132,N_9616,N_9502);
nor U10133 (N_10133,N_8556,N_8743);
or U10134 (N_10134,N_7968,N_9396);
and U10135 (N_10135,N_9522,N_8329);
nand U10136 (N_10136,N_9919,N_9006);
or U10137 (N_10137,N_7844,N_7685);
nand U10138 (N_10138,N_8161,N_7550);
and U10139 (N_10139,N_8188,N_7589);
nand U10140 (N_10140,N_7875,N_8360);
nand U10141 (N_10141,N_8467,N_9382);
nor U10142 (N_10142,N_8658,N_9409);
or U10143 (N_10143,N_8979,N_7766);
xnor U10144 (N_10144,N_9486,N_9453);
and U10145 (N_10145,N_9212,N_9368);
or U10146 (N_10146,N_8376,N_9157);
or U10147 (N_10147,N_9287,N_8050);
nor U10148 (N_10148,N_7585,N_9758);
xor U10149 (N_10149,N_7716,N_9511);
nand U10150 (N_10150,N_7901,N_9726);
or U10151 (N_10151,N_8983,N_8287);
nor U10152 (N_10152,N_8307,N_9651);
xor U10153 (N_10153,N_7597,N_7828);
and U10154 (N_10154,N_8878,N_7545);
or U10155 (N_10155,N_7783,N_7710);
nand U10156 (N_10156,N_8544,N_7959);
nor U10157 (N_10157,N_8279,N_8875);
or U10158 (N_10158,N_9826,N_8635);
nand U10159 (N_10159,N_9300,N_9349);
xor U10160 (N_10160,N_7837,N_9615);
nor U10161 (N_10161,N_9932,N_7992);
or U10162 (N_10162,N_9291,N_8230);
xor U10163 (N_10163,N_8859,N_8685);
xor U10164 (N_10164,N_7988,N_8051);
nor U10165 (N_10165,N_8303,N_9200);
nand U10166 (N_10166,N_8873,N_8599);
nand U10167 (N_10167,N_9077,N_9416);
nor U10168 (N_10168,N_8253,N_8883);
nand U10169 (N_10169,N_7691,N_7753);
xor U10170 (N_10170,N_9423,N_7843);
and U10171 (N_10171,N_8269,N_9998);
nor U10172 (N_10172,N_9640,N_8109);
or U10173 (N_10173,N_7969,N_8766);
and U10174 (N_10174,N_7517,N_8908);
nor U10175 (N_10175,N_9372,N_9531);
and U10176 (N_10176,N_9142,N_9425);
xnor U10177 (N_10177,N_9478,N_9732);
nor U10178 (N_10178,N_8010,N_9237);
nor U10179 (N_10179,N_8980,N_8861);
nor U10180 (N_10180,N_9725,N_9796);
nor U10181 (N_10181,N_8049,N_9168);
nor U10182 (N_10182,N_9069,N_9653);
nor U10183 (N_10183,N_9024,N_9628);
xnor U10184 (N_10184,N_8105,N_8839);
or U10185 (N_10185,N_9019,N_9505);
nand U10186 (N_10186,N_8185,N_9973);
nor U10187 (N_10187,N_7736,N_9652);
nand U10188 (N_10188,N_7806,N_9445);
nor U10189 (N_10189,N_9671,N_8002);
and U10190 (N_10190,N_8977,N_8835);
and U10191 (N_10191,N_9170,N_7506);
and U10192 (N_10192,N_8749,N_8308);
or U10193 (N_10193,N_9645,N_8963);
nand U10194 (N_10194,N_9232,N_9928);
xor U10195 (N_10195,N_9789,N_9713);
or U10196 (N_10196,N_8851,N_7810);
nand U10197 (N_10197,N_7755,N_8676);
and U10198 (N_10198,N_9623,N_9575);
nand U10199 (N_10199,N_7793,N_9948);
and U10200 (N_10200,N_8748,N_8154);
or U10201 (N_10201,N_7720,N_8723);
or U10202 (N_10202,N_8805,N_8447);
xor U10203 (N_10203,N_9045,N_9620);
nor U10204 (N_10204,N_9923,N_8104);
nand U10205 (N_10205,N_7808,N_8740);
or U10206 (N_10206,N_7970,N_8388);
and U10207 (N_10207,N_9807,N_8708);
nand U10208 (N_10208,N_9573,N_8140);
and U10209 (N_10209,N_8146,N_8089);
nand U10210 (N_10210,N_8033,N_9783);
nand U10211 (N_10211,N_9041,N_8610);
nor U10212 (N_10212,N_9954,N_7598);
nor U10213 (N_10213,N_8299,N_7788);
or U10214 (N_10214,N_9263,N_8710);
or U10215 (N_10215,N_9407,N_7953);
and U10216 (N_10216,N_8858,N_9410);
xor U10217 (N_10217,N_7756,N_8971);
or U10218 (N_10218,N_8236,N_7807);
xnor U10219 (N_10219,N_8356,N_9824);
xnor U10220 (N_10220,N_9563,N_9822);
and U10221 (N_10221,N_9847,N_7577);
and U10222 (N_10222,N_8426,N_7551);
and U10223 (N_10223,N_9335,N_8480);
nor U10224 (N_10224,N_8699,N_8565);
nand U10225 (N_10225,N_8918,N_9959);
nor U10226 (N_10226,N_9765,N_7511);
or U10227 (N_10227,N_7717,N_9099);
nand U10228 (N_10228,N_8233,N_7935);
xor U10229 (N_10229,N_9898,N_9345);
nor U10230 (N_10230,N_7519,N_8522);
nand U10231 (N_10231,N_8995,N_9538);
and U10232 (N_10232,N_8170,N_9360);
nor U10233 (N_10233,N_9268,N_8591);
nand U10234 (N_10234,N_9774,N_9754);
nand U10235 (N_10235,N_8557,N_9078);
or U10236 (N_10236,N_8155,N_9803);
or U10237 (N_10237,N_7879,N_8453);
and U10238 (N_10238,N_8261,N_9100);
xor U10239 (N_10239,N_7893,N_9264);
nor U10240 (N_10240,N_7592,N_8074);
or U10241 (N_10241,N_7811,N_8317);
and U10242 (N_10242,N_9418,N_9179);
and U10243 (N_10243,N_9249,N_9819);
xor U10244 (N_10244,N_8960,N_8479);
xnor U10245 (N_10245,N_7785,N_9446);
nand U10246 (N_10246,N_8911,N_9189);
nor U10247 (N_10247,N_9540,N_9072);
and U10248 (N_10248,N_9805,N_7859);
xnor U10249 (N_10249,N_9187,N_7599);
nand U10250 (N_10250,N_9700,N_8657);
nor U10251 (N_10251,N_8648,N_9761);
or U10252 (N_10252,N_8386,N_8058);
nand U10253 (N_10253,N_8190,N_9117);
and U10254 (N_10254,N_9317,N_7948);
xnor U10255 (N_10255,N_8359,N_9162);
or U10256 (N_10256,N_8346,N_7946);
and U10257 (N_10257,N_8174,N_9181);
xnor U10258 (N_10258,N_8596,N_8946);
or U10259 (N_10259,N_9378,N_9000);
nor U10260 (N_10260,N_9009,N_9526);
xnor U10261 (N_10261,N_8630,N_9295);
and U10262 (N_10262,N_7532,N_7726);
nor U10263 (N_10263,N_9058,N_7829);
and U10264 (N_10264,N_8331,N_9985);
and U10265 (N_10265,N_8701,N_9280);
xor U10266 (N_10266,N_9670,N_8643);
nand U10267 (N_10267,N_9790,N_8769);
or U10268 (N_10268,N_7882,N_7665);
nand U10269 (N_10269,N_8138,N_8674);
xor U10270 (N_10270,N_8297,N_9244);
or U10271 (N_10271,N_9008,N_7606);
and U10272 (N_10272,N_8905,N_8000);
or U10273 (N_10273,N_8474,N_8071);
and U10274 (N_10274,N_9052,N_9530);
nand U10275 (N_10275,N_8954,N_7708);
and U10276 (N_10276,N_9995,N_7998);
and U10277 (N_10277,N_8845,N_9091);
or U10278 (N_10278,N_9424,N_9716);
and U10279 (N_10279,N_8811,N_8439);
or U10280 (N_10280,N_8128,N_8678);
xor U10281 (N_10281,N_9897,N_8396);
nor U10282 (N_10282,N_9544,N_8921);
xnor U10283 (N_10283,N_7832,N_9140);
and U10284 (N_10284,N_9061,N_8405);
nor U10285 (N_10285,N_9687,N_9654);
xnor U10286 (N_10286,N_9584,N_9984);
or U10287 (N_10287,N_7911,N_9493);
nor U10288 (N_10288,N_9183,N_8836);
xnor U10289 (N_10289,N_9343,N_8466);
nor U10290 (N_10290,N_9250,N_7989);
nor U10291 (N_10291,N_7809,N_8131);
nor U10292 (N_10292,N_8540,N_8477);
nand U10293 (N_10293,N_8410,N_9144);
or U10294 (N_10294,N_8015,N_9498);
xnor U10295 (N_10295,N_7860,N_7981);
xnor U10296 (N_10296,N_7536,N_9946);
or U10297 (N_10297,N_8750,N_8250);
and U10298 (N_10298,N_8777,N_9610);
and U10299 (N_10299,N_9599,N_8536);
xnor U10300 (N_10300,N_7891,N_9027);
and U10301 (N_10301,N_9314,N_9906);
nand U10302 (N_10302,N_8870,N_9341);
and U10303 (N_10303,N_8473,N_9044);
or U10304 (N_10304,N_7887,N_9277);
xor U10305 (N_10305,N_9297,N_9468);
nand U10306 (N_10306,N_8633,N_8720);
and U10307 (N_10307,N_8489,N_8130);
nor U10308 (N_10308,N_9443,N_8907);
and U10309 (N_10309,N_9138,N_8559);
or U10310 (N_10310,N_8944,N_8882);
xnor U10311 (N_10311,N_9380,N_8320);
or U10312 (N_10312,N_8516,N_9888);
or U10313 (N_10313,N_8196,N_8273);
nor U10314 (N_10314,N_7883,N_7727);
nand U10315 (N_10315,N_7666,N_9982);
and U10316 (N_10316,N_7734,N_8829);
xnor U10317 (N_10317,N_8513,N_8520);
or U10318 (N_10318,N_9757,N_8673);
nor U10319 (N_10319,N_9243,N_9567);
nor U10320 (N_10320,N_8719,N_8264);
and U10321 (N_10321,N_9989,N_7707);
and U10322 (N_10322,N_9866,N_8592);
nor U10323 (N_10323,N_8468,N_8550);
nand U10324 (N_10324,N_9739,N_9806);
xor U10325 (N_10325,N_7672,N_9537);
and U10326 (N_10326,N_7885,N_9463);
nand U10327 (N_10327,N_9968,N_9987);
or U10328 (N_10328,N_9876,N_7840);
xor U10329 (N_10329,N_9436,N_7692);
and U10330 (N_10330,N_7584,N_8041);
or U10331 (N_10331,N_9634,N_7869);
nor U10332 (N_10332,N_9483,N_9167);
nor U10333 (N_10333,N_8248,N_7763);
nand U10334 (N_10334,N_8252,N_8456);
and U10335 (N_10335,N_9083,N_9145);
and U10336 (N_10336,N_9333,N_9627);
and U10337 (N_10337,N_8842,N_8246);
and U10338 (N_10338,N_8315,N_8120);
nand U10339 (N_10339,N_8948,N_7853);
or U10340 (N_10340,N_8693,N_8652);
nand U10341 (N_10341,N_7919,N_8132);
or U10342 (N_10342,N_8047,N_9683);
and U10343 (N_10343,N_9500,N_8849);
xor U10344 (N_10344,N_9238,N_7731);
nand U10345 (N_10345,N_9021,N_7512);
or U10346 (N_10346,N_9929,N_9541);
nor U10347 (N_10347,N_9172,N_9241);
nor U10348 (N_10348,N_8847,N_7586);
xor U10349 (N_10349,N_8432,N_7937);
and U10350 (N_10350,N_7956,N_8072);
and U10351 (N_10351,N_9708,N_7881);
nand U10352 (N_10352,N_9311,N_7648);
nor U10353 (N_10353,N_8589,N_9286);
or U10354 (N_10354,N_9804,N_7530);
xor U10355 (N_10355,N_7814,N_8691);
nand U10356 (N_10356,N_8087,N_8533);
nor U10357 (N_10357,N_8932,N_8505);
or U10358 (N_10358,N_7847,N_8784);
nand U10359 (N_10359,N_8363,N_8210);
or U10360 (N_10360,N_8172,N_7676);
nor U10361 (N_10361,N_8222,N_9840);
and U10362 (N_10362,N_7640,N_8152);
or U10363 (N_10363,N_9875,N_8198);
xnor U10364 (N_10364,N_9361,N_9093);
or U10365 (N_10365,N_8355,N_9637);
nor U10366 (N_10366,N_8324,N_9430);
nor U10367 (N_10367,N_9674,N_8731);
nand U10368 (N_10368,N_7928,N_8106);
nor U10369 (N_10369,N_9330,N_8133);
and U10370 (N_10370,N_9829,N_8837);
xor U10371 (N_10371,N_8666,N_8729);
or U10372 (N_10372,N_9626,N_8349);
nor U10373 (N_10373,N_7523,N_9120);
or U10374 (N_10374,N_8451,N_8339);
nand U10375 (N_10375,N_8245,N_9205);
and U10376 (N_10376,N_7588,N_8065);
nand U10377 (N_10377,N_7827,N_8227);
nor U10378 (N_10378,N_8820,N_8280);
nor U10379 (N_10379,N_9729,N_7518);
nor U10380 (N_10380,N_8169,N_9639);
nand U10381 (N_10381,N_7863,N_8367);
nand U10382 (N_10382,N_9961,N_9176);
nor U10383 (N_10383,N_8573,N_7730);
nand U10384 (N_10384,N_7718,N_9768);
and U10385 (N_10385,N_8398,N_9001);
nand U10386 (N_10386,N_8672,N_8695);
nor U10387 (N_10387,N_7943,N_8097);
nand U10388 (N_10388,N_7547,N_8793);
xor U10389 (N_10389,N_9970,N_8916);
xnor U10390 (N_10390,N_7960,N_9354);
or U10391 (N_10391,N_7980,N_8704);
nand U10392 (N_10392,N_9818,N_8919);
nor U10393 (N_10393,N_8413,N_9837);
nor U10394 (N_10394,N_9272,N_9855);
nand U10395 (N_10395,N_9677,N_8073);
nor U10396 (N_10396,N_8312,N_7595);
xor U10397 (N_10397,N_7918,N_9472);
and U10398 (N_10398,N_8900,N_9028);
and U10399 (N_10399,N_9967,N_7765);
nor U10400 (N_10400,N_8787,N_8939);
or U10401 (N_10401,N_8499,N_8902);
nor U10402 (N_10402,N_9026,N_7632);
nand U10403 (N_10403,N_8342,N_8497);
nor U10404 (N_10404,N_7688,N_9398);
xor U10405 (N_10405,N_9163,N_8706);
nand U10406 (N_10406,N_9597,N_8226);
xor U10407 (N_10407,N_9110,N_9160);
nand U10408 (N_10408,N_8276,N_8953);
and U10409 (N_10409,N_9477,N_7607);
nor U10410 (N_10410,N_9568,N_7906);
or U10411 (N_10411,N_8929,N_8554);
and U10412 (N_10412,N_9572,N_9825);
or U10413 (N_10413,N_8962,N_8665);
nor U10414 (N_10414,N_8463,N_8333);
and U10415 (N_10415,N_9031,N_9766);
xnor U10416 (N_10416,N_7673,N_7945);
xor U10417 (N_10417,N_7997,N_8488);
nor U10418 (N_10418,N_7680,N_8562);
nand U10419 (N_10419,N_7789,N_9814);
or U10420 (N_10420,N_7541,N_8752);
nand U10421 (N_10421,N_8271,N_9321);
and U10422 (N_10422,N_9042,N_9583);
and U10423 (N_10423,N_7826,N_8627);
nand U10424 (N_10424,N_9838,N_7534);
or U10425 (N_10425,N_9235,N_9592);
xnor U10426 (N_10426,N_7645,N_9356);
xor U10427 (N_10427,N_9960,N_9289);
and U10428 (N_10428,N_8458,N_9508);
nand U10429 (N_10429,N_7623,N_8868);
or U10430 (N_10430,N_9743,N_8716);
xor U10431 (N_10431,N_9208,N_8700);
nand U10432 (N_10432,N_9185,N_8780);
nor U10433 (N_10433,N_8259,N_9523);
or U10434 (N_10434,N_9704,N_9509);
xor U10435 (N_10435,N_7790,N_9900);
or U10436 (N_10436,N_7721,N_8853);
xor U10437 (N_10437,N_9499,N_8524);
and U10438 (N_10438,N_8402,N_9852);
and U10439 (N_10439,N_9794,N_8906);
and U10440 (N_10440,N_9293,N_7849);
nor U10441 (N_10441,N_7531,N_9223);
or U10442 (N_10442,N_8998,N_8904);
xnor U10443 (N_10443,N_8668,N_8585);
nor U10444 (N_10444,N_8580,N_7993);
nor U10445 (N_10445,N_9059,N_8325);
nor U10446 (N_10446,N_9780,N_7917);
or U10447 (N_10447,N_9388,N_8124);
nand U10448 (N_10448,N_8661,N_7915);
nand U10449 (N_10449,N_9992,N_9089);
or U10450 (N_10450,N_8733,N_9426);
nand U10451 (N_10451,N_9731,N_8866);
and U10452 (N_10452,N_9455,N_8760);
xnor U10453 (N_10453,N_8019,N_7723);
and U10454 (N_10454,N_9942,N_8774);
and U10455 (N_10455,N_7569,N_7501);
or U10456 (N_10456,N_9164,N_8880);
xnor U10457 (N_10457,N_8455,N_9247);
and U10458 (N_10458,N_9827,N_7564);
or U10459 (N_10459,N_8770,N_9112);
nor U10460 (N_10460,N_8738,N_7643);
and U10461 (N_10461,N_9074,N_7583);
or U10462 (N_10462,N_7633,N_7566);
or U10463 (N_10463,N_9283,N_9763);
nor U10464 (N_10464,N_8048,N_8045);
nand U10465 (N_10465,N_8521,N_8119);
xor U10466 (N_10466,N_7841,N_8370);
nand U10467 (N_10467,N_9673,N_8266);
xor U10468 (N_10468,N_8772,N_8571);
xnor U10469 (N_10469,N_8205,N_7582);
nor U10470 (N_10470,N_8149,N_9403);
nand U10471 (N_10471,N_8263,N_9373);
or U10472 (N_10472,N_9375,N_8283);
xnor U10473 (N_10473,N_7752,N_9705);
xnor U10474 (N_10474,N_8506,N_9465);
nand U10475 (N_10475,N_9744,N_9706);
and U10476 (N_10476,N_9482,N_9776);
and U10477 (N_10477,N_7618,N_8741);
xor U10478 (N_10478,N_8290,N_8897);
xor U10479 (N_10479,N_8644,N_8326);
nor U10480 (N_10480,N_9933,N_7504);
nor U10481 (N_10481,N_8181,N_8144);
and U10482 (N_10482,N_7694,N_8208);
nand U10483 (N_10483,N_8076,N_8403);
nor U10484 (N_10484,N_8327,N_8620);
nor U10485 (N_10485,N_8425,N_9503);
xnor U10486 (N_10486,N_9355,N_8898);
or U10487 (N_10487,N_8850,N_8920);
and U10488 (N_10488,N_9381,N_9565);
and U10489 (N_10489,N_8029,N_8877);
nor U10490 (N_10490,N_8353,N_9606);
or U10491 (N_10491,N_8150,N_8624);
or U10492 (N_10492,N_7987,N_9150);
nand U10493 (N_10493,N_7562,N_8235);
and U10494 (N_10494,N_9618,N_9219);
or U10495 (N_10495,N_8539,N_9326);
and U10496 (N_10496,N_8424,N_9778);
xor U10497 (N_10497,N_8176,N_8301);
or U10498 (N_10498,N_8372,N_8608);
nand U10499 (N_10499,N_8257,N_9772);
nor U10500 (N_10500,N_7936,N_7903);
nor U10501 (N_10501,N_7698,N_8147);
xor U10502 (N_10502,N_8053,N_8197);
and U10503 (N_10503,N_8914,N_8517);
nand U10504 (N_10504,N_9159,N_7747);
xnor U10505 (N_10505,N_8282,N_7854);
or U10506 (N_10506,N_8158,N_8064);
nor U10507 (N_10507,N_9411,N_8697);
xor U10508 (N_10508,N_8800,N_7516);
xnor U10509 (N_10509,N_8690,N_8484);
nor U10510 (N_10510,N_8319,N_7897);
and U10511 (N_10511,N_8876,N_9994);
nand U10512 (N_10512,N_8637,N_9841);
nor U10513 (N_10513,N_8978,N_9557);
xnor U10514 (N_10514,N_8959,N_8495);
and U10515 (N_10515,N_8448,N_7667);
and U10516 (N_10516,N_9676,N_7794);
and U10517 (N_10517,N_8808,N_9504);
or U10518 (N_10518,N_8854,N_9534);
nor U10519 (N_10519,N_8457,N_8588);
xor U10520 (N_10520,N_7743,N_8195);
or U10521 (N_10521,N_8481,N_8838);
nor U10522 (N_10522,N_9632,N_8813);
nor U10523 (N_10523,N_8828,N_9966);
and U10524 (N_10524,N_9712,N_8885);
and U10525 (N_10525,N_8881,N_9785);
nand U10526 (N_10526,N_8221,N_8083);
xor U10527 (N_10527,N_8538,N_8936);
or U10528 (N_10528,N_7833,N_8997);
xor U10529 (N_10529,N_7851,N_9979);
nor U10530 (N_10530,N_7801,N_8179);
or U10531 (N_10531,N_9427,N_8471);
nand U10532 (N_10532,N_9691,N_9533);
or U10533 (N_10533,N_8044,N_8419);
nand U10534 (N_10534,N_8304,N_8910);
or U10535 (N_10535,N_9820,N_9958);
nand U10536 (N_10536,N_7750,N_8567);
nand U10537 (N_10537,N_8270,N_9149);
or U10538 (N_10538,N_7681,N_8546);
xor U10539 (N_10539,N_7744,N_9609);
or U10540 (N_10540,N_8404,N_9608);
nor U10541 (N_10541,N_8587,N_9113);
nor U10542 (N_10542,N_9204,N_9656);
nand U10543 (N_10543,N_8306,N_8692);
xnor U10544 (N_10544,N_7861,N_7778);
nand U10545 (N_10545,N_7912,N_8518);
or U10546 (N_10546,N_9920,N_8951);
or U10547 (N_10547,N_7800,N_8091);
xor U10548 (N_10548,N_8846,N_9390);
nor U10549 (N_10549,N_9257,N_9064);
nor U10550 (N_10550,N_9598,N_9285);
xor U10551 (N_10551,N_9893,N_7686);
or U10552 (N_10552,N_7741,N_9600);
nor U10553 (N_10553,N_9020,N_8490);
or U10554 (N_10554,N_9218,N_9489);
or U10555 (N_10555,N_9461,N_8990);
nand U10556 (N_10556,N_7904,N_8328);
nand U10557 (N_10557,N_8651,N_8572);
or U10558 (N_10558,N_8218,N_9351);
and U10559 (N_10559,N_9879,N_8203);
nand U10560 (N_10560,N_8159,N_9332);
nor U10561 (N_10561,N_8732,N_7626);
or U10562 (N_10562,N_8985,N_8392);
and U10563 (N_10563,N_8823,N_7889);
or U10564 (N_10564,N_8177,N_9460);
nand U10565 (N_10565,N_8046,N_8260);
and U10566 (N_10566,N_8440,N_9730);
nand U10567 (N_10567,N_9296,N_9941);
xnor U10568 (N_10568,N_8094,N_9962);
nor U10569 (N_10569,N_7803,N_9454);
xor U10570 (N_10570,N_9738,N_8412);
nand U10571 (N_10571,N_9166,N_9348);
nand U10572 (N_10572,N_8759,N_9603);
or U10573 (N_10573,N_8400,N_8348);
nor U10574 (N_10574,N_9350,N_8187);
or U10575 (N_10575,N_7644,N_7762);
nor U10576 (N_10576,N_8734,N_9322);
nand U10577 (N_10577,N_9607,N_9023);
or U10578 (N_10578,N_9365,N_8206);
nand U10579 (N_10579,N_7831,N_8930);
nand U10580 (N_10580,N_8117,N_7952);
nor U10581 (N_10581,N_8100,N_9714);
nand U10582 (N_10582,N_8462,N_9229);
nand U10583 (N_10583,N_8581,N_7759);
and U10584 (N_10584,N_8892,N_9611);
xor U10585 (N_10585,N_9073,N_8586);
xor U10586 (N_10586,N_8442,N_7751);
and U10587 (N_10587,N_7733,N_8114);
nor U10588 (N_10588,N_9551,N_7554);
xnor U10589 (N_10589,N_8016,N_8703);
xor U10590 (N_10590,N_9178,N_7876);
or U10591 (N_10591,N_9097,N_9234);
or U10592 (N_10592,N_8933,N_9862);
and U10593 (N_10593,N_7514,N_9194);
and U10594 (N_10594,N_7898,N_7999);
and U10595 (N_10595,N_9613,N_7926);
xor U10596 (N_10596,N_8335,N_9672);
nand U10597 (N_10597,N_9101,N_9809);
xor U10598 (N_10598,N_8289,N_8744);
and U10599 (N_10599,N_8519,N_9419);
or U10600 (N_10600,N_7871,N_8530);
nor U10601 (N_10601,N_8136,N_7624);
and U10602 (N_10602,N_8042,N_9895);
nor U10603 (N_10603,N_8852,N_9861);
nor U10604 (N_10604,N_9660,N_8103);
nand U10605 (N_10605,N_7907,N_8783);
xor U10606 (N_10606,N_7653,N_8220);
xor U10607 (N_10607,N_8611,N_9635);
or U10608 (N_10608,N_7700,N_9851);
nand U10609 (N_10609,N_8574,N_7950);
xor U10610 (N_10610,N_8173,N_8284);
xor U10611 (N_10611,N_8949,N_9931);
or U10612 (N_10612,N_9578,N_7925);
nor U10613 (N_10613,N_9927,N_7674);
nand U10614 (N_10614,N_9107,N_9779);
nand U10615 (N_10615,N_9002,N_8646);
or U10616 (N_10616,N_9740,N_8476);
nand U10617 (N_10617,N_9476,N_7812);
or U10618 (N_10618,N_9536,N_8275);
or U10619 (N_10619,N_9310,N_7923);
nand U10620 (N_10620,N_9914,N_8696);
or U10621 (N_10621,N_9562,N_9030);
nor U10622 (N_10622,N_7894,N_9193);
nand U10623 (N_10623,N_9742,N_7590);
xor U10624 (N_10624,N_9561,N_9856);
or U10625 (N_10625,N_8237,N_7933);
nand U10626 (N_10626,N_8156,N_7619);
and U10627 (N_10627,N_7966,N_8415);
nand U10628 (N_10628,N_9082,N_9680);
or U10629 (N_10629,N_8790,N_7748);
and U10630 (N_10630,N_7715,N_8228);
nor U10631 (N_10631,N_8600,N_8578);
and U10632 (N_10632,N_9727,N_8108);
nand U10633 (N_10633,N_7973,N_9554);
xnor U10634 (N_10634,N_8407,N_9007);
nand U10635 (N_10635,N_9126,N_8925);
xnor U10636 (N_10636,N_9733,N_8612);
nor U10637 (N_10637,N_7631,N_9574);
nor U10638 (N_10638,N_9214,N_8414);
nor U10639 (N_10639,N_7983,N_9899);
and U10640 (N_10640,N_7796,N_9891);
and U10641 (N_10641,N_9753,N_7571);
xor U10642 (N_10642,N_8894,N_8232);
and U10643 (N_10643,N_9532,N_9394);
or U10644 (N_10644,N_9196,N_9309);
nand U10645 (N_10645,N_7782,N_9466);
xor U10646 (N_10646,N_8022,N_8318);
nand U10647 (N_10647,N_9955,N_7573);
nor U10648 (N_10648,N_9791,N_7527);
and U10649 (N_10649,N_7627,N_9924);
nor U10650 (N_10650,N_9957,N_9273);
nor U10651 (N_10651,N_8242,N_7820);
nor U10652 (N_10652,N_8247,N_7649);
and U10653 (N_10653,N_8027,N_8028);
nor U10654 (N_10654,N_9642,N_9153);
nand U10655 (N_10655,N_8291,N_8025);
nor U10656 (N_10656,N_9589,N_9487);
or U10657 (N_10657,N_8507,N_8958);
xnor U10658 (N_10658,N_7947,N_8986);
xnor U10659 (N_10659,N_7600,N_7602);
and U10660 (N_10660,N_7539,N_8768);
or U10661 (N_10661,N_9233,N_9337);
or U10662 (N_10662,N_8865,N_8680);
nor U10663 (N_10663,N_8382,N_9549);
nand U10664 (N_10664,N_9944,N_7574);
nand U10665 (N_10665,N_8736,N_8689);
and U10666 (N_10666,N_9633,N_7888);
xor U10667 (N_10667,N_9594,N_9702);
xor U10668 (N_10668,N_9952,N_8343);
nor U10669 (N_10669,N_8341,N_8955);
and U10670 (N_10670,N_8543,N_9062);
nor U10671 (N_10671,N_8515,N_9395);
nor U10672 (N_10672,N_8262,N_7705);
xnor U10673 (N_10673,N_9593,N_7722);
and U10674 (N_10674,N_8496,N_7818);
nor U10675 (N_10675,N_8340,N_8655);
nand U10676 (N_10676,N_8107,N_9749);
xnor U10677 (N_10677,N_9102,N_9865);
nand U10678 (N_10678,N_7746,N_9227);
or U10679 (N_10679,N_8782,N_9217);
and U10680 (N_10680,N_8675,N_9131);
nor U10681 (N_10681,N_8084,N_8189);
nor U10682 (N_10682,N_9515,N_9010);
nor U10683 (N_10683,N_9545,N_9605);
or U10684 (N_10684,N_9972,N_7855);
xnor U10685 (N_10685,N_9867,N_9793);
nand U10686 (N_10686,N_9576,N_8475);
nand U10687 (N_10687,N_8385,N_8534);
nand U10688 (N_10688,N_7757,N_9242);
nand U10689 (N_10689,N_8779,N_8395);
nand U10690 (N_10690,N_7908,N_9174);
xor U10691 (N_10691,N_8192,N_7910);
xor U10692 (N_10692,N_8013,N_9199);
xnor U10693 (N_10693,N_8775,N_8889);
and U10694 (N_10694,N_9892,N_8924);
and U10695 (N_10695,N_8713,N_8653);
xor U10696 (N_10696,N_8298,N_9889);
nor U10697 (N_10697,N_9890,N_9636);
nand U10698 (N_10698,N_8080,N_7714);
nand U10699 (N_10699,N_8619,N_8670);
xor U10700 (N_10700,N_9055,N_9198);
and U10701 (N_10701,N_7500,N_9012);
nand U10702 (N_10702,N_9068,N_8984);
or U10703 (N_10703,N_8406,N_9156);
and U10704 (N_10704,N_7620,N_8310);
nand U10705 (N_10705,N_8761,N_9281);
and U10706 (N_10706,N_7899,N_7994);
xor U10707 (N_10707,N_9520,N_8613);
nor U10708 (N_10708,N_8821,N_8714);
and U10709 (N_10709,N_9516,N_9649);
xor U10710 (N_10710,N_8043,N_9550);
nand U10711 (N_10711,N_9118,N_8802);
xnor U10712 (N_10712,N_9081,N_8444);
and U10713 (N_10713,N_8305,N_8183);
nor U10714 (N_10714,N_7729,N_9590);
or U10715 (N_10715,N_8240,N_8137);
and U10716 (N_10716,N_8088,N_7760);
or U10717 (N_10717,N_7524,N_9921);
or U10718 (N_10718,N_9070,N_9412);
or U10719 (N_10719,N_9588,N_9323);
and U10720 (N_10720,N_9231,N_7678);
and U10721 (N_10721,N_7677,N_7965);
and U10722 (N_10722,N_7684,N_9513);
xnor U10723 (N_10723,N_9088,N_9950);
and U10724 (N_10724,N_9276,N_8758);
or U10725 (N_10725,N_8295,N_9947);
and U10726 (N_10726,N_9885,N_8012);
nor U10727 (N_10727,N_9325,N_8604);
nor U10728 (N_10728,N_8616,N_8576);
nand U10729 (N_10729,N_9748,N_8867);
nand U10730 (N_10730,N_8168,N_9695);
or U10731 (N_10731,N_8617,N_9675);
and U10732 (N_10732,N_9566,N_8746);
nand U10733 (N_10733,N_8035,N_8052);
and U10734 (N_10734,N_9288,N_9721);
and U10735 (N_10735,N_7522,N_8641);
nand U10736 (N_10736,N_8636,N_8994);
and U10737 (N_10737,N_8662,N_8486);
nand U10738 (N_10738,N_9109,N_8542);
or U10739 (N_10739,N_9366,N_8681);
nand U10740 (N_10740,N_9259,N_9621);
or U10741 (N_10741,N_8068,N_9329);
nor U10742 (N_10742,N_7605,N_9147);
and U10743 (N_10743,N_8638,N_9444);
nor U10744 (N_10744,N_8465,N_8472);
nor U10745 (N_10745,N_9991,N_7836);
nand U10746 (N_10746,N_8127,N_8940);
nor U10747 (N_10747,N_9130,N_8201);
or U10748 (N_10748,N_8863,N_8903);
and U10749 (N_10749,N_9029,N_9775);
and U10750 (N_10750,N_7628,N_8938);
xnor U10751 (N_10751,N_9978,N_8739);
or U10752 (N_10752,N_8764,N_8122);
and U10753 (N_10753,N_8056,N_8216);
xor U10754 (N_10754,N_9839,N_7990);
nand U10755 (N_10755,N_8274,N_8148);
nor U10756 (N_10756,N_9441,N_9983);
xor U10757 (N_10757,N_8224,N_8869);
or U10758 (N_10758,N_8552,N_8803);
nor U10759 (N_10759,N_9266,N_7622);
xor U10760 (N_10760,N_8508,N_9539);
xnor U10761 (N_10761,N_9747,N_8762);
or U10762 (N_10762,N_9546,N_9456);
and U10763 (N_10763,N_7922,N_8293);
xor U10764 (N_10764,N_8460,N_7799);
or U10765 (N_10765,N_7661,N_7659);
nor U10766 (N_10766,N_8566,N_8548);
xor U10767 (N_10767,N_7957,N_7774);
nand U10768 (N_10768,N_7892,N_8632);
and U10769 (N_10769,N_8647,N_8129);
nor U10770 (N_10770,N_8514,N_9746);
and U10771 (N_10771,N_8957,N_9836);
nor U10772 (N_10772,N_9559,N_7975);
xor U10773 (N_10773,N_8886,N_7779);
nor U10774 (N_10774,N_8055,N_8926);
and U10775 (N_10775,N_9619,N_7670);
or U10776 (N_10776,N_8755,N_8603);
nand U10777 (N_10777,N_9462,N_9431);
and U10778 (N_10778,N_7868,N_8656);
and U10779 (N_10779,N_9975,N_9857);
and U10780 (N_10780,N_7538,N_9769);
nand U10781 (N_10781,N_9079,N_9490);
nand U10782 (N_10782,N_7510,N_7986);
xnor U10783 (N_10783,N_8211,N_8649);
nand U10784 (N_10784,N_8267,N_7971);
nor U10785 (N_10785,N_9940,N_9090);
xnor U10786 (N_10786,N_9392,N_9141);
nand U10787 (N_10787,N_8175,N_8972);
nand U10788 (N_10788,N_9414,N_8207);
or U10789 (N_10789,N_8915,N_9389);
nor U10790 (N_10790,N_7578,N_9452);
and U10791 (N_10791,N_9450,N_8323);
and U10792 (N_10792,N_9304,N_8857);
nor U10793 (N_10793,N_9013,N_8628);
nand U10794 (N_10794,N_7929,N_9479);
xnor U10795 (N_10795,N_9442,N_9737);
nor U10796 (N_10796,N_9269,N_7594);
nor U10797 (N_10797,N_9016,N_8812);
nor U10798 (N_10798,N_9032,N_9971);
xor U10799 (N_10799,N_9813,N_7815);
nor U10800 (N_10800,N_9771,N_8063);
and U10801 (N_10801,N_9173,N_8679);
nand U10802 (N_10802,N_8569,N_8711);
xor U10803 (N_10803,N_8167,N_8526);
xor U10804 (N_10804,N_8730,N_8584);
nor U10805 (N_10805,N_7544,N_7557);
nand U10806 (N_10806,N_9930,N_9066);
nor U10807 (N_10807,N_8737,N_8202);
nor U10808 (N_10808,N_9239,N_9770);
or U10809 (N_10809,N_8365,N_7775);
xnor U10810 (N_10810,N_9564,N_8964);
nor U10811 (N_10811,N_8031,N_8785);
nand U10812 (N_10812,N_8917,N_8214);
xnor U10813 (N_10813,N_8164,N_7711);
nand U10814 (N_10814,N_8966,N_8618);
or U10815 (N_10815,N_9521,N_9622);
or U10816 (N_10816,N_9161,N_9529);
nand U10817 (N_10817,N_9784,N_7902);
and U10818 (N_10818,N_8030,N_9363);
nand U10819 (N_10819,N_8255,N_9306);
or U10820 (N_10820,N_8387,N_8856);
or U10821 (N_10821,N_8895,N_9724);
nand U10822 (N_10822,N_8969,N_7977);
xnor U10823 (N_10823,N_9186,N_9710);
or U10824 (N_10824,N_8441,N_9969);
and U10825 (N_10825,N_8818,N_8057);
or U10826 (N_10826,N_8888,N_8640);
xor U10827 (N_10827,N_8855,N_7699);
nor U10828 (N_10828,N_8429,N_8922);
xor U10829 (N_10829,N_9226,N_9981);
nor U10830 (N_10830,N_7921,N_9894);
nand U10831 (N_10831,N_9340,N_9106);
nand U10832 (N_10832,N_9111,N_8251);
nand U10833 (N_10833,N_8294,N_8527);
or U10834 (N_10834,N_9034,N_8671);
nand U10835 (N_10835,N_9352,N_9256);
nor U10836 (N_10836,N_8879,N_9225);
nand U10837 (N_10837,N_7740,N_9903);
or U10838 (N_10838,N_8937,N_8241);
nand U10839 (N_10839,N_7560,N_9542);
nor U10840 (N_10840,N_9665,N_7963);
nand U10841 (N_10841,N_9122,N_8135);
and U10842 (N_10842,N_9496,N_7749);
nor U10843 (N_10843,N_9228,N_9507);
xnor U10844 (N_10844,N_8239,N_7636);
nand U10845 (N_10845,N_8893,N_8234);
xor U10846 (N_10846,N_8694,N_8862);
and U10847 (N_10847,N_9916,N_9274);
xor U10848 (N_10848,N_8973,N_9644);
nor U10849 (N_10849,N_8928,N_9376);
nor U10850 (N_10850,N_9402,N_8834);
and U10851 (N_10851,N_9997,N_8090);
nand U10852 (N_10852,N_9255,N_8423);
nand U10853 (N_10853,N_7895,N_7976);
or U10854 (N_10854,N_8334,N_9367);
xor U10855 (N_10855,N_7526,N_8564);
and U10856 (N_10856,N_7725,N_7873);
or U10857 (N_10857,N_8126,N_9114);
nand U10858 (N_10858,N_8092,N_8311);
and U10859 (N_10859,N_9781,N_9751);
nand U10860 (N_10860,N_9934,N_8535);
xnor U10861 (N_10861,N_8366,N_9849);
nand U10862 (N_10862,N_9525,N_9684);
or U10863 (N_10863,N_8717,N_8931);
nand U10864 (N_10864,N_8593,N_9667);
nor U10865 (N_10865,N_9327,N_7764);
xor U10866 (N_10866,N_8354,N_9488);
and U10867 (N_10867,N_7795,N_9773);
or U10868 (N_10868,N_9917,N_8322);
or U10869 (N_10869,N_8864,N_8493);
and U10870 (N_10870,N_9422,N_9964);
nor U10871 (N_10871,N_7575,N_9661);
nor U10872 (N_10872,N_8551,N_8110);
or U10873 (N_10873,N_9527,N_9755);
nand U10874 (N_10874,N_9986,N_7770);
and U10875 (N_10875,N_8278,N_7690);
or U10876 (N_10876,N_9202,N_8884);
nand U10877 (N_10877,N_7629,N_7896);
nand U10878 (N_10878,N_7533,N_8531);
nand U10879 (N_10879,N_8745,N_9220);
nor U10880 (N_10880,N_9270,N_7612);
nand U10881 (N_10881,N_9158,N_8664);
xnor U10882 (N_10882,N_9292,N_8165);
or U10883 (N_10883,N_9802,N_8452);
xor U10884 (N_10884,N_8547,N_8011);
xnor U10885 (N_10885,N_9902,N_7886);
xnor U10886 (N_10886,N_8583,N_8113);
and U10887 (N_10887,N_9926,N_9832);
and U10888 (N_10888,N_9434,N_9711);
xor U10889 (N_10889,N_9084,N_8379);
nand U10890 (N_10890,N_9799,N_9191);
or U10891 (N_10891,N_9816,N_9261);
nor U10892 (N_10892,N_9722,N_9795);
nand U10893 (N_10893,N_8988,N_7570);
or U10894 (N_10894,N_9098,N_8134);
xor U10895 (N_10895,N_7664,N_9629);
and U10896 (N_10896,N_9399,N_7675);
xor U10897 (N_10897,N_8470,N_9116);
nor U10898 (N_10898,N_9548,N_9553);
and U10899 (N_10899,N_8614,N_8602);
and U10900 (N_10900,N_8786,N_7838);
xor U10901 (N_10901,N_7839,N_9386);
and U10902 (N_10902,N_9451,N_9307);
xor U10903 (N_10903,N_9279,N_9543);
nor U10904 (N_10904,N_8338,N_8747);
nor U10905 (N_10905,N_8347,N_8626);
xor U10906 (N_10906,N_8428,N_8558);
and U10907 (N_10907,N_7797,N_7679);
or U10908 (N_10908,N_8077,N_9797);
xor U10909 (N_10909,N_7958,N_8607);
xnor U10910 (N_10910,N_8590,N_8023);
and U10911 (N_10911,N_9886,N_8860);
xnor U10912 (N_10912,N_9121,N_8778);
or U10913 (N_10913,N_7568,N_9484);
nand U10914 (N_10914,N_8622,N_9951);
nor U10915 (N_10915,N_9896,N_8162);
nand U10916 (N_10916,N_8112,N_8810);
nand U10917 (N_10917,N_8003,N_7932);
nand U10918 (N_10918,N_9641,N_9717);
nand U10919 (N_10919,N_9254,N_8116);
nand U10920 (N_10920,N_8004,N_9956);
xnor U10921 (N_10921,N_7703,N_8416);
nand U10922 (N_10922,N_8781,N_8258);
and U10923 (N_10923,N_7529,N_9469);
nand U10924 (N_10924,N_8688,N_7528);
and U10925 (N_10925,N_7916,N_8912);
or U10926 (N_10926,N_8215,N_9353);
and U10927 (N_10927,N_8767,N_7652);
nor U10928 (N_10928,N_8735,N_8143);
nor U10929 (N_10929,N_8935,N_8660);
nand U10930 (N_10930,N_9085,N_7593);
or U10931 (N_10931,N_8391,N_9346);
nand U10932 (N_10932,N_8418,N_9988);
and U10933 (N_10933,N_9133,N_7630);
nor U10934 (N_10934,N_8193,N_8725);
xnor U10935 (N_10935,N_9025,N_9777);
xor U10936 (N_10936,N_9420,N_9524);
and U10937 (N_10937,N_8545,N_9095);
xnor U10938 (N_10938,N_8018,N_9638);
nor U10939 (N_10939,N_7509,N_8244);
or U10940 (N_10940,N_8789,N_7941);
xor U10941 (N_10941,N_9312,N_8634);
or U10942 (N_10942,N_8709,N_9320);
or U10943 (N_10943,N_9440,N_9871);
nand U10944 (N_10944,N_9215,N_7773);
nor U10945 (N_10945,N_9004,N_9943);
and U10946 (N_10946,N_7954,N_8832);
xnor U10947 (N_10947,N_9686,N_8844);
or U10948 (N_10948,N_9308,N_8438);
nand U10949 (N_10949,N_8118,N_8445);
or U10950 (N_10950,N_9883,N_9689);
nand U10951 (N_10951,N_7712,N_9087);
or U10952 (N_10952,N_7996,N_7617);
and U10953 (N_10953,N_8814,N_9192);
xor U10954 (N_10954,N_7742,N_9129);
and U10955 (N_10955,N_7761,N_8449);
nand U10956 (N_10956,N_9209,N_7656);
nor U10957 (N_10957,N_8454,N_7651);
nor U10958 (N_10958,N_7507,N_9874);
xor U10959 (N_10959,N_9175,N_9709);
nand U10960 (N_10960,N_8006,N_8577);
or U10961 (N_10961,N_9571,N_7955);
or U10962 (N_10962,N_8036,N_7931);
nor U10963 (N_10963,N_9909,N_9169);
xor U10964 (N_10964,N_9152,N_8511);
nand U10965 (N_10965,N_9782,N_9197);
nand U10966 (N_10966,N_9036,N_9762);
nand U10967 (N_10967,N_8757,N_9397);
and U10968 (N_10968,N_8199,N_7657);
or U10969 (N_10969,N_9911,N_8687);
or U10970 (N_10970,N_7542,N_8500);
nand U10971 (N_10971,N_9359,N_9552);
nor U10972 (N_10972,N_9063,N_8171);
or U10973 (N_10973,N_7978,N_8826);
and U10974 (N_10974,N_7548,N_8067);
nand U10975 (N_10975,N_8032,N_7842);
or U10976 (N_10976,N_8238,N_8796);
or U10977 (N_10977,N_7587,N_7776);
and U10978 (N_10978,N_9715,N_8361);
xnor U10979 (N_10979,N_9222,N_9510);
nor U10980 (N_10980,N_7787,N_9703);
or U10981 (N_10981,N_7834,N_9338);
nand U10982 (N_10982,N_7737,N_9901);
or U10983 (N_10983,N_8078,N_8629);
nor U10984 (N_10984,N_8815,N_9850);
xor U10985 (N_10985,N_9788,N_7576);
nor U10986 (N_10986,N_7823,N_9810);
and U10987 (N_10987,N_8296,N_9076);
nand U10988 (N_10988,N_7767,N_9248);
or U10989 (N_10989,N_7638,N_7662);
nor U10990 (N_10990,N_9213,N_9171);
or U10991 (N_10991,N_7798,N_7939);
xor U10992 (N_10992,N_9371,N_9694);
or U10993 (N_10993,N_9835,N_9693);
and U10994 (N_10994,N_9812,N_9432);
nor U10995 (N_10995,N_7804,N_8791);
nand U10996 (N_10996,N_8560,N_8987);
and U10997 (N_10997,N_9580,N_9165);
xnor U10998 (N_10998,N_7866,N_8191);
xnor U10999 (N_10999,N_7639,N_8194);
nor U11000 (N_11000,N_9643,N_8976);
nand U11001 (N_11001,N_8792,N_7553);
nand U11002 (N_11002,N_7920,N_9301);
or U11003 (N_11003,N_8887,N_7660);
xnor U11004 (N_11004,N_9387,N_8901);
nor U11005 (N_11005,N_8373,N_9630);
xnor U11006 (N_11006,N_9245,N_8420);
nand U11007 (N_11007,N_8797,N_7735);
and U11008 (N_11008,N_8085,N_8605);
nand U11009 (N_11009,N_8357,N_8509);
and U11010 (N_11010,N_9663,N_9480);
and U11011 (N_11011,N_8313,N_9401);
xnor U11012 (N_11012,N_9720,N_8843);
xnor U11013 (N_11013,N_8345,N_8595);
and U11014 (N_11014,N_9648,N_8212);
and U11015 (N_11015,N_8059,N_9060);
or U11016 (N_11016,N_9669,N_9154);
nand U11017 (N_11017,N_8899,N_7864);
xnor U11018 (N_11018,N_9830,N_8125);
and U11019 (N_11019,N_8020,N_9935);
nor U11020 (N_11020,N_9863,N_9435);
xor U11021 (N_11021,N_8582,N_7870);
and U11022 (N_11022,N_8186,N_8014);
nor U11023 (N_11023,N_7913,N_7930);
and U11024 (N_11024,N_7967,N_8389);
or U11025 (N_11025,N_9907,N_8794);
xnor U11026 (N_11026,N_7822,N_7772);
nor U11027 (N_11027,N_9831,N_9035);
nand U11028 (N_11028,N_9650,N_7687);
nor U11029 (N_11029,N_8913,N_9519);
nor U11030 (N_11030,N_9868,N_8034);
nor U11031 (N_11031,N_9404,N_8101);
nor U11032 (N_11032,N_9370,N_7940);
nor U11033 (N_11033,N_9688,N_8292);
or U11034 (N_11034,N_9017,N_7769);
xnor U11035 (N_11035,N_7515,N_8249);
and U11036 (N_11036,N_9313,N_9251);
or U11037 (N_11037,N_9377,N_9668);
nand U11038 (N_11038,N_7909,N_8795);
and U11039 (N_11039,N_7985,N_9180);
xor U11040 (N_11040,N_7713,N_8427);
nor U11041 (N_11041,N_9210,N_9764);
xor U11042 (N_11042,N_8431,N_9357);
xnor U11043 (N_11043,N_9517,N_8742);
xor U11044 (N_11044,N_8459,N_9051);
or U11045 (N_11045,N_8555,N_8950);
xor U11046 (N_11046,N_9369,N_9535);
or U11047 (N_11047,N_8231,N_9383);
or U11048 (N_11048,N_8705,N_7867);
nand U11049 (N_11049,N_8601,N_9290);
or U11050 (N_11050,N_8368,N_8408);
xnor U11051 (N_11051,N_9556,N_8991);
nor U11052 (N_11052,N_8840,N_8650);
nand U11053 (N_11053,N_7505,N_8970);
or U11054 (N_11054,N_8285,N_9136);
nor U11055 (N_11055,N_9043,N_7621);
or U11056 (N_11056,N_8469,N_9033);
nor U11057 (N_11057,N_9858,N_7611);
nor U11058 (N_11058,N_9612,N_9470);
nand U11059 (N_11059,N_9054,N_9614);
nand U11060 (N_11060,N_7995,N_8099);
and U11061 (N_11061,N_9146,N_8434);
nand U11062 (N_11062,N_7540,N_7525);
or U11063 (N_11063,N_9437,N_9123);
xor U11064 (N_11064,N_9342,N_9569);
or U11065 (N_11065,N_7739,N_8433);
or U11066 (N_11066,N_9679,N_9870);
nand U11067 (N_11067,N_7642,N_9458);
xnor U11068 (N_11068,N_7724,N_9904);
and U11069 (N_11069,N_9405,N_9302);
nand U11070 (N_11070,N_9316,N_8833);
nand U11071 (N_11071,N_8756,N_9201);
xnor U11072 (N_11072,N_7984,N_8502);
and U11073 (N_11073,N_9143,N_9391);
xor U11074 (N_11074,N_8062,N_8153);
nor U11075 (N_11075,N_7850,N_8302);
or U11076 (N_11076,N_7819,N_8393);
xnor U11077 (N_11077,N_7556,N_9071);
nor U11078 (N_11078,N_8026,N_8005);
or U11079 (N_11079,N_9384,N_7613);
and U11080 (N_11080,N_7543,N_9408);
or U11081 (N_11081,N_8008,N_9303);
xor U11082 (N_11082,N_8390,N_7878);
nor U11083 (N_11083,N_9996,N_9625);
nand U11084 (N_11084,N_9275,N_7596);
or U11085 (N_11085,N_8316,N_8848);
and U11086 (N_11086,N_8217,N_9860);
nor U11087 (N_11087,N_9501,N_9662);
nand U11088 (N_11088,N_7503,N_9908);
and U11089 (N_11089,N_9570,N_8332);
nor U11090 (N_11090,N_8281,N_9701);
or U11091 (N_11091,N_9728,N_9318);
nand U11092 (N_11092,N_9278,N_7905);
or U11093 (N_11093,N_9808,N_8254);
and U11094 (N_11094,N_7830,N_9447);
nand U11095 (N_11095,N_7615,N_9127);
xor U11096 (N_11096,N_8160,N_8350);
xnor U11097 (N_11097,N_8364,N_8483);
or U11098 (N_11098,N_9474,N_8371);
nor U11099 (N_11099,N_8358,N_8180);
and U11100 (N_11100,N_9492,N_8831);
xnor U11101 (N_11101,N_7591,N_7781);
and U11102 (N_11102,N_7535,N_8992);
and U11103 (N_11103,N_9624,N_9075);
or U11104 (N_11104,N_8378,N_9224);
nand U11105 (N_11105,N_9696,N_7817);
nor U11106 (N_11106,N_8485,N_9128);
and U11107 (N_11107,N_8721,N_7924);
nand U11108 (N_11108,N_8763,N_9364);
xnor U11109 (N_11109,N_8975,N_8243);
or U11110 (N_11110,N_9843,N_9587);
xnor U11111 (N_11111,N_8209,N_8645);
nor U11112 (N_11112,N_8968,N_8824);
nand U11113 (N_11113,N_9881,N_8093);
nor U11114 (N_11114,N_7758,N_8461);
or U11115 (N_11115,N_8934,N_9869);
xor U11116 (N_11116,N_9939,N_7816);
xnor U11117 (N_11117,N_9155,N_9877);
and U11118 (N_11118,N_7858,N_8942);
nor U11119 (N_11119,N_9953,N_7862);
and U11120 (N_11120,N_8061,N_7655);
xnor U11121 (N_11121,N_8799,N_8623);
nand U11122 (N_11122,N_9206,N_7974);
xnor U11123 (N_11123,N_8945,N_9115);
nor U11124 (N_11124,N_9132,N_9833);
and U11125 (N_11125,N_9211,N_8075);
nand U11126 (N_11126,N_9601,N_7608);
or U11127 (N_11127,N_9880,N_8464);
and U11128 (N_11128,N_9406,N_7567);
or U11129 (N_11129,N_8598,N_8896);
nand U11130 (N_11130,N_8669,N_9821);
and U11131 (N_11131,N_9976,N_7745);
or U11132 (N_11132,N_9745,N_9823);
nor U11133 (N_11133,N_8309,N_9018);
xnor U11134 (N_11134,N_7646,N_9848);
and U11135 (N_11135,N_8722,N_8151);
and U11136 (N_11136,N_8288,N_7821);
nand U11137 (N_11137,N_7579,N_8715);
and U11138 (N_11138,N_7695,N_9844);
or U11139 (N_11139,N_7991,N_8686);
xor U11140 (N_11140,N_9659,N_9056);
nor U11141 (N_11141,N_8369,N_8871);
nor U11142 (N_11142,N_8443,N_8809);
or U11143 (N_11143,N_7701,N_9040);
nand U11144 (N_11144,N_7845,N_9379);
nand U11145 (N_11145,N_9828,N_8086);
nand U11146 (N_11146,N_9736,N_9864);
xor U11147 (N_11147,N_8478,N_7549);
or U11148 (N_11148,N_8038,N_9258);
nor U11149 (N_11149,N_8272,N_9050);
and U11150 (N_11150,N_9011,N_8683);
xor U11151 (N_11151,N_9385,N_8446);
or U11152 (N_11152,N_7857,N_9003);
or U11153 (N_11153,N_8615,N_9236);
and U11154 (N_11154,N_9190,N_7890);
nor U11155 (N_11155,N_8874,N_8397);
xnor U11156 (N_11156,N_9977,N_8096);
or U11157 (N_11157,N_7521,N_7825);
and U11158 (N_11158,N_7802,N_7900);
xor U11159 (N_11159,N_9912,N_9678);
nand U11160 (N_11160,N_9015,N_8575);
nand U11161 (N_11161,N_8830,N_9859);
xor U11162 (N_11162,N_9750,N_8718);
xnor U11163 (N_11163,N_9037,N_8166);
xor U11164 (N_11164,N_9177,N_9965);
nor U11165 (N_11165,N_9305,N_9752);
or U11166 (N_11166,N_9324,N_8082);
and U11167 (N_11167,N_7792,N_9882);
xnor U11168 (N_11168,N_9315,N_7934);
nand U11169 (N_11169,N_9938,N_7559);
or U11170 (N_11170,N_9105,N_9707);
nor U11171 (N_11171,N_8277,N_7689);
nand U11172 (N_11172,N_8597,N_9602);
or U11173 (N_11173,N_8204,N_8139);
nor U11174 (N_11174,N_8111,N_9666);
nor U11175 (N_11175,N_8568,N_9872);
nand U11176 (N_11176,N_9913,N_9137);
and U11177 (N_11177,N_8806,N_8300);
xor U11178 (N_11178,N_9049,N_9362);
or U11179 (N_11179,N_9299,N_9294);
nor U11180 (N_11180,N_9887,N_8563);
nand U11181 (N_11181,N_9038,N_9936);
xor U11182 (N_11182,N_9252,N_8684);
and U11183 (N_11183,N_9328,N_9697);
nor U11184 (N_11184,N_9604,N_7552);
nand U11185 (N_11185,N_8394,N_9910);
nand U11186 (N_11186,N_9358,N_9735);
nor U11187 (N_11187,N_8001,N_9595);
and U11188 (N_11188,N_7951,N_8123);
xor U11189 (N_11189,N_9591,N_9103);
and U11190 (N_11190,N_9974,N_9512);
or U11191 (N_11191,N_7637,N_9260);
or U11192 (N_11192,N_8952,N_8532);
nand U11193 (N_11193,N_9922,N_8528);
and U11194 (N_11194,N_8223,N_8712);
nor U11195 (N_11195,N_8999,N_9925);
and U11196 (N_11196,N_8377,N_9993);
nor U11197 (N_11197,N_9134,N_7848);
nand U11198 (N_11198,N_8375,N_9657);
nor U11199 (N_11199,N_9148,N_8807);
nand U11200 (N_11200,N_8549,N_7961);
nand U11201 (N_11201,N_9096,N_9558);
xor U11202 (N_11202,N_9682,N_9271);
xor U11203 (N_11203,N_7791,N_8399);
or U11204 (N_11204,N_8362,N_8726);
nor U11205 (N_11205,N_9547,N_9692);
and U11206 (N_11206,N_8606,N_7513);
and U11207 (N_11207,N_7846,N_9846);
or U11208 (N_11208,N_9344,N_8336);
nor U11209 (N_11209,N_9801,N_7634);
nand U11210 (N_11210,N_9617,N_7949);
and U11211 (N_11211,N_9506,N_9884);
xnor U11212 (N_11212,N_7520,N_7558);
and U11213 (N_11213,N_9786,N_9582);
xnor U11214 (N_11214,N_9048,N_8982);
and U11215 (N_11215,N_7696,N_8037);
nand U11216 (N_11216,N_8178,N_9080);
nor U11217 (N_11217,N_8529,N_9467);
nand U11218 (N_11218,N_8352,N_9022);
and U11219 (N_11219,N_7663,N_9005);
and U11220 (N_11220,N_8337,N_8677);
xnor U11221 (N_11221,N_8890,N_7972);
or U11222 (N_11222,N_8200,N_7738);
and U11223 (N_11223,N_7979,N_8947);
nand U11224 (N_11224,N_7682,N_7647);
nor U11225 (N_11225,N_9053,N_8967);
or U11226 (N_11226,N_8503,N_8069);
nor U11227 (N_11227,N_7754,N_8102);
and U11228 (N_11228,N_9497,N_9151);
and U11229 (N_11229,N_9336,N_9756);
and U11230 (N_11230,N_7805,N_9980);
and U11231 (N_11231,N_9655,N_9815);
xor U11232 (N_11232,N_9681,N_8504);
xor U11233 (N_11233,N_9092,N_8639);
xnor U11234 (N_11234,N_9094,N_9596);
xnor U11235 (N_11235,N_9298,N_9429);
nor U11236 (N_11236,N_9873,N_8079);
nor U11237 (N_11237,N_9413,N_8384);
nand U11238 (N_11238,N_9428,N_7555);
nor U11239 (N_11239,N_8501,N_7813);
and U11240 (N_11240,N_7635,N_7502);
nand U11241 (N_11241,N_7942,N_8754);
or U11242 (N_11242,N_7572,N_8553);
xnor U11243 (N_11243,N_8625,N_7780);
nor U11244 (N_11244,N_9119,N_7625);
and U11245 (N_11245,N_9459,N_9195);
and U11246 (N_11246,N_8381,N_7702);
nand U11247 (N_11247,N_9393,N_8727);
nor U11248 (N_11248,N_8491,N_7658);
and U11249 (N_11249,N_8066,N_9182);
nor U11250 (N_11250,N_7714,N_9329);
nor U11251 (N_11251,N_7907,N_8202);
xor U11252 (N_11252,N_8430,N_9185);
xnor U11253 (N_11253,N_9387,N_8288);
nand U11254 (N_11254,N_7873,N_8832);
nor U11255 (N_11255,N_9744,N_7651);
nor U11256 (N_11256,N_8748,N_7981);
and U11257 (N_11257,N_9761,N_8824);
xnor U11258 (N_11258,N_8094,N_8994);
xnor U11259 (N_11259,N_9637,N_8102);
xor U11260 (N_11260,N_8931,N_9696);
xor U11261 (N_11261,N_8567,N_8281);
and U11262 (N_11262,N_9950,N_8867);
or U11263 (N_11263,N_7926,N_9995);
nand U11264 (N_11264,N_8777,N_9325);
and U11265 (N_11265,N_9353,N_9748);
and U11266 (N_11266,N_9827,N_9226);
nand U11267 (N_11267,N_9800,N_8141);
xor U11268 (N_11268,N_7560,N_7689);
xnor U11269 (N_11269,N_7810,N_9905);
xnor U11270 (N_11270,N_8269,N_8719);
xor U11271 (N_11271,N_8395,N_7935);
nor U11272 (N_11272,N_8409,N_9986);
nand U11273 (N_11273,N_8216,N_7733);
or U11274 (N_11274,N_7660,N_9867);
xor U11275 (N_11275,N_7786,N_8486);
xor U11276 (N_11276,N_8343,N_8598);
xor U11277 (N_11277,N_9359,N_7579);
nand U11278 (N_11278,N_9575,N_7503);
or U11279 (N_11279,N_9303,N_8539);
or U11280 (N_11280,N_9730,N_9227);
nand U11281 (N_11281,N_9034,N_8039);
nor U11282 (N_11282,N_8258,N_9735);
or U11283 (N_11283,N_7713,N_8231);
nor U11284 (N_11284,N_9931,N_9052);
or U11285 (N_11285,N_8932,N_9581);
xor U11286 (N_11286,N_8528,N_8452);
nor U11287 (N_11287,N_9645,N_8562);
or U11288 (N_11288,N_7884,N_9070);
and U11289 (N_11289,N_9895,N_8795);
xnor U11290 (N_11290,N_8120,N_9017);
and U11291 (N_11291,N_7739,N_9968);
and U11292 (N_11292,N_9139,N_9821);
or U11293 (N_11293,N_7928,N_8069);
nor U11294 (N_11294,N_7774,N_8510);
and U11295 (N_11295,N_8057,N_8162);
and U11296 (N_11296,N_9857,N_8999);
and U11297 (N_11297,N_8018,N_8769);
or U11298 (N_11298,N_7541,N_9413);
nand U11299 (N_11299,N_9390,N_9734);
or U11300 (N_11300,N_8785,N_7899);
xor U11301 (N_11301,N_8981,N_9465);
nand U11302 (N_11302,N_9269,N_9984);
xor U11303 (N_11303,N_9973,N_8220);
nor U11304 (N_11304,N_7712,N_8373);
nand U11305 (N_11305,N_9927,N_7858);
nor U11306 (N_11306,N_9788,N_8550);
nand U11307 (N_11307,N_9223,N_7661);
nand U11308 (N_11308,N_8238,N_8878);
xor U11309 (N_11309,N_9708,N_7890);
or U11310 (N_11310,N_8951,N_9368);
nor U11311 (N_11311,N_8284,N_8273);
xor U11312 (N_11312,N_7901,N_7612);
and U11313 (N_11313,N_9640,N_7627);
nor U11314 (N_11314,N_8012,N_7537);
nand U11315 (N_11315,N_9490,N_8474);
nor U11316 (N_11316,N_8055,N_7881);
or U11317 (N_11317,N_9159,N_8900);
xnor U11318 (N_11318,N_7625,N_8098);
or U11319 (N_11319,N_8000,N_9466);
and U11320 (N_11320,N_9492,N_8851);
nand U11321 (N_11321,N_8385,N_9325);
or U11322 (N_11322,N_9769,N_8800);
or U11323 (N_11323,N_8672,N_8945);
or U11324 (N_11324,N_8466,N_9644);
or U11325 (N_11325,N_9919,N_9134);
or U11326 (N_11326,N_8197,N_9844);
and U11327 (N_11327,N_8624,N_8225);
xnor U11328 (N_11328,N_9394,N_7588);
or U11329 (N_11329,N_9145,N_8703);
or U11330 (N_11330,N_9981,N_8280);
xor U11331 (N_11331,N_8492,N_9647);
and U11332 (N_11332,N_7513,N_8398);
nand U11333 (N_11333,N_9660,N_9873);
nand U11334 (N_11334,N_9954,N_9213);
and U11335 (N_11335,N_9587,N_7920);
or U11336 (N_11336,N_9423,N_8835);
nor U11337 (N_11337,N_7945,N_8483);
nand U11338 (N_11338,N_7997,N_8694);
or U11339 (N_11339,N_8853,N_8858);
and U11340 (N_11340,N_9597,N_9335);
xnor U11341 (N_11341,N_9057,N_8865);
or U11342 (N_11342,N_9230,N_8638);
and U11343 (N_11343,N_9389,N_8884);
nand U11344 (N_11344,N_8577,N_9822);
or U11345 (N_11345,N_8588,N_7934);
and U11346 (N_11346,N_9313,N_9991);
or U11347 (N_11347,N_8092,N_7709);
nor U11348 (N_11348,N_9684,N_8757);
nand U11349 (N_11349,N_9090,N_9835);
nor U11350 (N_11350,N_8427,N_9378);
xor U11351 (N_11351,N_8314,N_8296);
xor U11352 (N_11352,N_8997,N_9710);
nor U11353 (N_11353,N_9022,N_8895);
nand U11354 (N_11354,N_8710,N_7765);
and U11355 (N_11355,N_9697,N_8772);
nor U11356 (N_11356,N_9811,N_9092);
or U11357 (N_11357,N_8936,N_8599);
nand U11358 (N_11358,N_8291,N_7925);
nand U11359 (N_11359,N_7906,N_9321);
or U11360 (N_11360,N_8905,N_8281);
and U11361 (N_11361,N_9786,N_8315);
or U11362 (N_11362,N_8945,N_9734);
xor U11363 (N_11363,N_7516,N_9267);
xnor U11364 (N_11364,N_7918,N_8276);
and U11365 (N_11365,N_7645,N_9298);
nor U11366 (N_11366,N_8992,N_8697);
nor U11367 (N_11367,N_8408,N_8291);
or U11368 (N_11368,N_9620,N_8090);
nor U11369 (N_11369,N_8270,N_7955);
xnor U11370 (N_11370,N_7906,N_8336);
or U11371 (N_11371,N_8618,N_9395);
nor U11372 (N_11372,N_9842,N_7813);
xor U11373 (N_11373,N_9036,N_7999);
and U11374 (N_11374,N_9385,N_9561);
nand U11375 (N_11375,N_9319,N_8573);
and U11376 (N_11376,N_8736,N_9796);
nand U11377 (N_11377,N_7645,N_7985);
and U11378 (N_11378,N_8179,N_8188);
xnor U11379 (N_11379,N_9787,N_8268);
and U11380 (N_11380,N_9531,N_8979);
xor U11381 (N_11381,N_9094,N_7680);
or U11382 (N_11382,N_9176,N_9878);
and U11383 (N_11383,N_9829,N_9022);
and U11384 (N_11384,N_9983,N_7828);
or U11385 (N_11385,N_9176,N_9237);
and U11386 (N_11386,N_8108,N_9256);
nand U11387 (N_11387,N_8059,N_9967);
nor U11388 (N_11388,N_8787,N_8020);
nand U11389 (N_11389,N_8626,N_9234);
and U11390 (N_11390,N_9135,N_9741);
nand U11391 (N_11391,N_9026,N_8235);
nor U11392 (N_11392,N_8715,N_9203);
xor U11393 (N_11393,N_7945,N_9624);
nor U11394 (N_11394,N_9868,N_9180);
nand U11395 (N_11395,N_9829,N_9386);
nand U11396 (N_11396,N_8962,N_8013);
or U11397 (N_11397,N_9977,N_8703);
nand U11398 (N_11398,N_9118,N_8987);
nand U11399 (N_11399,N_8658,N_9220);
and U11400 (N_11400,N_9908,N_8302);
nor U11401 (N_11401,N_7919,N_9887);
nor U11402 (N_11402,N_7701,N_8077);
nor U11403 (N_11403,N_9556,N_8024);
or U11404 (N_11404,N_9995,N_9923);
nor U11405 (N_11405,N_7575,N_8530);
nor U11406 (N_11406,N_8963,N_8923);
nand U11407 (N_11407,N_7779,N_8365);
and U11408 (N_11408,N_9144,N_8290);
or U11409 (N_11409,N_9374,N_7599);
and U11410 (N_11410,N_8924,N_7899);
and U11411 (N_11411,N_8600,N_8961);
and U11412 (N_11412,N_8474,N_9869);
xnor U11413 (N_11413,N_8523,N_9721);
and U11414 (N_11414,N_9307,N_8222);
nor U11415 (N_11415,N_7660,N_8878);
xnor U11416 (N_11416,N_9639,N_8345);
xor U11417 (N_11417,N_8127,N_9391);
xnor U11418 (N_11418,N_9062,N_9767);
and U11419 (N_11419,N_9884,N_7575);
or U11420 (N_11420,N_8402,N_9330);
xnor U11421 (N_11421,N_8957,N_9287);
xnor U11422 (N_11422,N_8342,N_9077);
xnor U11423 (N_11423,N_7907,N_9639);
xor U11424 (N_11424,N_7952,N_9112);
or U11425 (N_11425,N_9904,N_8190);
nor U11426 (N_11426,N_9687,N_7511);
nor U11427 (N_11427,N_9324,N_7810);
nor U11428 (N_11428,N_7584,N_8477);
or U11429 (N_11429,N_9432,N_9180);
xor U11430 (N_11430,N_8992,N_9067);
xnor U11431 (N_11431,N_9183,N_9444);
nand U11432 (N_11432,N_9484,N_9089);
and U11433 (N_11433,N_8940,N_8945);
xnor U11434 (N_11434,N_9575,N_9400);
or U11435 (N_11435,N_8482,N_8116);
or U11436 (N_11436,N_9666,N_7723);
nor U11437 (N_11437,N_8404,N_8470);
nand U11438 (N_11438,N_9869,N_8758);
nand U11439 (N_11439,N_8323,N_9793);
nand U11440 (N_11440,N_9925,N_9782);
or U11441 (N_11441,N_9024,N_8706);
and U11442 (N_11442,N_7750,N_8566);
and U11443 (N_11443,N_8484,N_7896);
and U11444 (N_11444,N_8457,N_8967);
nand U11445 (N_11445,N_8382,N_9114);
xnor U11446 (N_11446,N_8206,N_9965);
or U11447 (N_11447,N_8650,N_9353);
or U11448 (N_11448,N_8043,N_7923);
nor U11449 (N_11449,N_9126,N_8329);
nand U11450 (N_11450,N_9430,N_8139);
xnor U11451 (N_11451,N_8344,N_7818);
nor U11452 (N_11452,N_8978,N_8929);
and U11453 (N_11453,N_8723,N_9593);
nor U11454 (N_11454,N_8388,N_7503);
nand U11455 (N_11455,N_9777,N_9020);
nor U11456 (N_11456,N_8046,N_7835);
or U11457 (N_11457,N_7589,N_9055);
or U11458 (N_11458,N_9859,N_7510);
or U11459 (N_11459,N_7786,N_7955);
nor U11460 (N_11460,N_8961,N_9060);
nand U11461 (N_11461,N_8982,N_8643);
or U11462 (N_11462,N_7597,N_8979);
or U11463 (N_11463,N_9623,N_9648);
nor U11464 (N_11464,N_8400,N_7928);
and U11465 (N_11465,N_8672,N_7870);
xnor U11466 (N_11466,N_9466,N_7501);
or U11467 (N_11467,N_8502,N_9868);
or U11468 (N_11468,N_9033,N_8227);
or U11469 (N_11469,N_8151,N_8915);
and U11470 (N_11470,N_9370,N_9972);
xor U11471 (N_11471,N_9160,N_9766);
xor U11472 (N_11472,N_9432,N_8167);
or U11473 (N_11473,N_8162,N_7638);
nor U11474 (N_11474,N_9277,N_8212);
or U11475 (N_11475,N_8492,N_8299);
nor U11476 (N_11476,N_8137,N_7883);
xor U11477 (N_11477,N_8965,N_9069);
and U11478 (N_11478,N_8153,N_7797);
and U11479 (N_11479,N_8829,N_7688);
and U11480 (N_11480,N_8662,N_8548);
or U11481 (N_11481,N_8223,N_8534);
and U11482 (N_11482,N_8483,N_9326);
xnor U11483 (N_11483,N_7535,N_8412);
and U11484 (N_11484,N_8202,N_9338);
xor U11485 (N_11485,N_9845,N_9859);
xor U11486 (N_11486,N_8798,N_8903);
xnor U11487 (N_11487,N_9384,N_9758);
nand U11488 (N_11488,N_8263,N_9502);
nor U11489 (N_11489,N_7750,N_8691);
and U11490 (N_11490,N_9871,N_9437);
and U11491 (N_11491,N_9104,N_8151);
or U11492 (N_11492,N_9587,N_9872);
and U11493 (N_11493,N_8495,N_7977);
nand U11494 (N_11494,N_9472,N_8555);
and U11495 (N_11495,N_9870,N_9247);
xnor U11496 (N_11496,N_9222,N_9372);
xor U11497 (N_11497,N_8975,N_8741);
nor U11498 (N_11498,N_9067,N_8872);
or U11499 (N_11499,N_9767,N_8603);
or U11500 (N_11500,N_8987,N_8610);
or U11501 (N_11501,N_9376,N_9104);
or U11502 (N_11502,N_8786,N_9634);
nor U11503 (N_11503,N_8378,N_7954);
nor U11504 (N_11504,N_9259,N_7566);
nand U11505 (N_11505,N_9315,N_9084);
nand U11506 (N_11506,N_9349,N_7928);
nand U11507 (N_11507,N_9646,N_8884);
nand U11508 (N_11508,N_7527,N_8098);
nand U11509 (N_11509,N_9478,N_8976);
nand U11510 (N_11510,N_9569,N_8360);
nor U11511 (N_11511,N_8974,N_7545);
xor U11512 (N_11512,N_8077,N_7923);
nand U11513 (N_11513,N_8007,N_8628);
and U11514 (N_11514,N_8592,N_8154);
and U11515 (N_11515,N_7547,N_9025);
xnor U11516 (N_11516,N_9658,N_9178);
xnor U11517 (N_11517,N_8908,N_9849);
or U11518 (N_11518,N_8834,N_8647);
and U11519 (N_11519,N_7981,N_9962);
nor U11520 (N_11520,N_7638,N_7539);
xnor U11521 (N_11521,N_7778,N_7915);
nand U11522 (N_11522,N_8342,N_8730);
nor U11523 (N_11523,N_8105,N_7521);
or U11524 (N_11524,N_9227,N_9676);
nor U11525 (N_11525,N_8977,N_9212);
and U11526 (N_11526,N_7926,N_9638);
xnor U11527 (N_11527,N_9440,N_9503);
and U11528 (N_11528,N_8230,N_9106);
nor U11529 (N_11529,N_8416,N_8793);
and U11530 (N_11530,N_8836,N_9109);
xor U11531 (N_11531,N_7814,N_8809);
and U11532 (N_11532,N_8869,N_9590);
xnor U11533 (N_11533,N_7854,N_9481);
nand U11534 (N_11534,N_8270,N_8788);
xor U11535 (N_11535,N_9815,N_8395);
xor U11536 (N_11536,N_8035,N_9491);
or U11537 (N_11537,N_8948,N_8748);
or U11538 (N_11538,N_8978,N_8185);
and U11539 (N_11539,N_9523,N_8670);
nand U11540 (N_11540,N_9778,N_8634);
xor U11541 (N_11541,N_9866,N_9303);
and U11542 (N_11542,N_7982,N_9470);
nand U11543 (N_11543,N_9774,N_8675);
nor U11544 (N_11544,N_8504,N_8914);
or U11545 (N_11545,N_9042,N_8660);
or U11546 (N_11546,N_8835,N_9172);
nand U11547 (N_11547,N_8311,N_8098);
xnor U11548 (N_11548,N_7797,N_9383);
nor U11549 (N_11549,N_9927,N_9478);
nor U11550 (N_11550,N_8652,N_9380);
xnor U11551 (N_11551,N_8817,N_9114);
nand U11552 (N_11552,N_9202,N_7731);
nor U11553 (N_11553,N_9468,N_9877);
and U11554 (N_11554,N_7849,N_8454);
nand U11555 (N_11555,N_9765,N_9268);
xnor U11556 (N_11556,N_8242,N_8900);
and U11557 (N_11557,N_9433,N_9263);
xnor U11558 (N_11558,N_8983,N_9628);
xnor U11559 (N_11559,N_7972,N_8309);
nand U11560 (N_11560,N_7528,N_7772);
nor U11561 (N_11561,N_8062,N_9585);
xor U11562 (N_11562,N_9897,N_9293);
nor U11563 (N_11563,N_9531,N_8805);
and U11564 (N_11564,N_7660,N_8340);
or U11565 (N_11565,N_9764,N_9717);
and U11566 (N_11566,N_7523,N_7945);
or U11567 (N_11567,N_9818,N_8960);
or U11568 (N_11568,N_9151,N_8744);
nor U11569 (N_11569,N_9705,N_8663);
and U11570 (N_11570,N_9438,N_8022);
nand U11571 (N_11571,N_9013,N_9344);
xnor U11572 (N_11572,N_8756,N_7732);
and U11573 (N_11573,N_9454,N_9814);
nand U11574 (N_11574,N_9349,N_9384);
xor U11575 (N_11575,N_8794,N_9560);
or U11576 (N_11576,N_9100,N_8781);
and U11577 (N_11577,N_9271,N_7874);
or U11578 (N_11578,N_9156,N_8005);
nand U11579 (N_11579,N_9036,N_9656);
xnor U11580 (N_11580,N_9393,N_8021);
xor U11581 (N_11581,N_7959,N_8970);
and U11582 (N_11582,N_9795,N_8898);
or U11583 (N_11583,N_8009,N_7730);
nor U11584 (N_11584,N_8361,N_8054);
nor U11585 (N_11585,N_7720,N_9056);
and U11586 (N_11586,N_8214,N_8795);
and U11587 (N_11587,N_9320,N_9936);
nor U11588 (N_11588,N_9680,N_8793);
xnor U11589 (N_11589,N_7661,N_8183);
or U11590 (N_11590,N_9488,N_8113);
and U11591 (N_11591,N_9515,N_9022);
and U11592 (N_11592,N_8677,N_9221);
or U11593 (N_11593,N_8512,N_9751);
xnor U11594 (N_11594,N_7817,N_9447);
and U11595 (N_11595,N_9231,N_7925);
nand U11596 (N_11596,N_9804,N_7916);
and U11597 (N_11597,N_8578,N_9818);
nand U11598 (N_11598,N_8731,N_9687);
xor U11599 (N_11599,N_9172,N_9118);
nand U11600 (N_11600,N_8842,N_8133);
nand U11601 (N_11601,N_9346,N_7821);
xor U11602 (N_11602,N_9199,N_7702);
xnor U11603 (N_11603,N_9042,N_7690);
nand U11604 (N_11604,N_9284,N_8634);
xnor U11605 (N_11605,N_8537,N_9644);
or U11606 (N_11606,N_9895,N_8589);
or U11607 (N_11607,N_9639,N_9244);
and U11608 (N_11608,N_8078,N_7632);
nand U11609 (N_11609,N_8948,N_9341);
nor U11610 (N_11610,N_7786,N_8643);
nor U11611 (N_11611,N_9916,N_7641);
nor U11612 (N_11612,N_9536,N_8274);
or U11613 (N_11613,N_9233,N_8916);
nor U11614 (N_11614,N_9883,N_9892);
or U11615 (N_11615,N_7738,N_9009);
and U11616 (N_11616,N_9269,N_7544);
nor U11617 (N_11617,N_9203,N_9505);
and U11618 (N_11618,N_7706,N_8843);
and U11619 (N_11619,N_8405,N_7948);
nand U11620 (N_11620,N_8242,N_9099);
or U11621 (N_11621,N_7953,N_7706);
xor U11622 (N_11622,N_9918,N_9532);
and U11623 (N_11623,N_7544,N_8495);
or U11624 (N_11624,N_8977,N_9080);
or U11625 (N_11625,N_9947,N_7866);
nand U11626 (N_11626,N_8172,N_9627);
nand U11627 (N_11627,N_8437,N_9522);
and U11628 (N_11628,N_9914,N_7702);
and U11629 (N_11629,N_7522,N_9119);
xnor U11630 (N_11630,N_8820,N_9013);
and U11631 (N_11631,N_8653,N_8470);
or U11632 (N_11632,N_7829,N_7976);
xnor U11633 (N_11633,N_8119,N_9270);
or U11634 (N_11634,N_9284,N_7542);
nand U11635 (N_11635,N_8993,N_8233);
nor U11636 (N_11636,N_9510,N_8773);
or U11637 (N_11637,N_9543,N_9050);
nor U11638 (N_11638,N_8515,N_9944);
nor U11639 (N_11639,N_8455,N_7866);
nor U11640 (N_11640,N_9917,N_9263);
xor U11641 (N_11641,N_9803,N_9146);
nor U11642 (N_11642,N_9149,N_8050);
nand U11643 (N_11643,N_9080,N_9637);
or U11644 (N_11644,N_8169,N_8456);
nand U11645 (N_11645,N_8904,N_9810);
or U11646 (N_11646,N_7674,N_9762);
or U11647 (N_11647,N_9862,N_8542);
and U11648 (N_11648,N_9169,N_9910);
xnor U11649 (N_11649,N_8425,N_8849);
and U11650 (N_11650,N_7624,N_9762);
xor U11651 (N_11651,N_8607,N_9535);
xor U11652 (N_11652,N_9147,N_8476);
nor U11653 (N_11653,N_9427,N_9160);
nor U11654 (N_11654,N_8712,N_8202);
or U11655 (N_11655,N_8004,N_9327);
nor U11656 (N_11656,N_9179,N_7864);
nor U11657 (N_11657,N_8128,N_9270);
nand U11658 (N_11658,N_8419,N_8469);
nor U11659 (N_11659,N_9575,N_9037);
xor U11660 (N_11660,N_9670,N_8037);
and U11661 (N_11661,N_7608,N_9145);
nor U11662 (N_11662,N_9819,N_9581);
and U11663 (N_11663,N_8171,N_8941);
nor U11664 (N_11664,N_7723,N_7765);
and U11665 (N_11665,N_9487,N_8814);
nand U11666 (N_11666,N_9439,N_9027);
nand U11667 (N_11667,N_8104,N_8698);
or U11668 (N_11668,N_8245,N_8224);
or U11669 (N_11669,N_8701,N_7822);
or U11670 (N_11670,N_9158,N_9090);
xor U11671 (N_11671,N_8260,N_8980);
nand U11672 (N_11672,N_9654,N_8405);
nor U11673 (N_11673,N_9151,N_8673);
nand U11674 (N_11674,N_9652,N_8321);
xor U11675 (N_11675,N_7591,N_8758);
and U11676 (N_11676,N_9566,N_8644);
or U11677 (N_11677,N_8234,N_9243);
xor U11678 (N_11678,N_8981,N_9250);
xnor U11679 (N_11679,N_8851,N_8452);
and U11680 (N_11680,N_8190,N_8489);
nor U11681 (N_11681,N_9453,N_7877);
or U11682 (N_11682,N_9920,N_9597);
nand U11683 (N_11683,N_9128,N_8053);
and U11684 (N_11684,N_8745,N_9812);
xor U11685 (N_11685,N_8679,N_8071);
and U11686 (N_11686,N_7968,N_9216);
xor U11687 (N_11687,N_7554,N_9549);
or U11688 (N_11688,N_9206,N_9621);
or U11689 (N_11689,N_8632,N_9994);
and U11690 (N_11690,N_7876,N_7849);
or U11691 (N_11691,N_9341,N_7914);
nand U11692 (N_11692,N_8447,N_9617);
nand U11693 (N_11693,N_9322,N_9184);
nor U11694 (N_11694,N_8165,N_9852);
or U11695 (N_11695,N_8861,N_8625);
xnor U11696 (N_11696,N_8652,N_8154);
or U11697 (N_11697,N_9062,N_7998);
or U11698 (N_11698,N_9008,N_7573);
xor U11699 (N_11699,N_8565,N_9069);
xnor U11700 (N_11700,N_9693,N_8594);
xnor U11701 (N_11701,N_9309,N_8254);
nor U11702 (N_11702,N_9620,N_9054);
nand U11703 (N_11703,N_8682,N_8421);
and U11704 (N_11704,N_9908,N_8076);
nand U11705 (N_11705,N_7658,N_9805);
and U11706 (N_11706,N_8527,N_8433);
nor U11707 (N_11707,N_9584,N_7693);
or U11708 (N_11708,N_9237,N_7783);
xor U11709 (N_11709,N_8870,N_8302);
nor U11710 (N_11710,N_9812,N_9255);
or U11711 (N_11711,N_9393,N_8140);
nor U11712 (N_11712,N_7980,N_9674);
and U11713 (N_11713,N_8005,N_9683);
nand U11714 (N_11714,N_8596,N_9888);
nor U11715 (N_11715,N_7966,N_9774);
xor U11716 (N_11716,N_8223,N_9724);
xor U11717 (N_11717,N_7894,N_8202);
or U11718 (N_11718,N_9408,N_9713);
and U11719 (N_11719,N_7674,N_7560);
or U11720 (N_11720,N_8368,N_8166);
nor U11721 (N_11721,N_8895,N_7665);
and U11722 (N_11722,N_7709,N_8028);
or U11723 (N_11723,N_9740,N_9352);
or U11724 (N_11724,N_7943,N_8312);
nor U11725 (N_11725,N_9590,N_8012);
or U11726 (N_11726,N_8236,N_8188);
and U11727 (N_11727,N_9430,N_8928);
and U11728 (N_11728,N_8482,N_7579);
or U11729 (N_11729,N_8512,N_7657);
nor U11730 (N_11730,N_8993,N_9143);
or U11731 (N_11731,N_9882,N_9305);
nor U11732 (N_11732,N_8514,N_9561);
and U11733 (N_11733,N_8311,N_8856);
nor U11734 (N_11734,N_8851,N_9912);
and U11735 (N_11735,N_9517,N_9306);
xor U11736 (N_11736,N_9647,N_7544);
xnor U11737 (N_11737,N_8467,N_8302);
and U11738 (N_11738,N_8679,N_8245);
xnor U11739 (N_11739,N_8176,N_8062);
or U11740 (N_11740,N_7650,N_8691);
nand U11741 (N_11741,N_9720,N_8237);
nand U11742 (N_11742,N_9070,N_9542);
and U11743 (N_11743,N_9479,N_7792);
or U11744 (N_11744,N_9567,N_8077);
or U11745 (N_11745,N_9278,N_7573);
or U11746 (N_11746,N_8099,N_9198);
xor U11747 (N_11747,N_7637,N_8216);
nor U11748 (N_11748,N_9562,N_8945);
xor U11749 (N_11749,N_9441,N_9264);
nand U11750 (N_11750,N_8522,N_8222);
xnor U11751 (N_11751,N_9989,N_8491);
and U11752 (N_11752,N_9033,N_8384);
or U11753 (N_11753,N_9968,N_9850);
and U11754 (N_11754,N_8850,N_7814);
or U11755 (N_11755,N_9149,N_9181);
nor U11756 (N_11756,N_7612,N_8968);
xnor U11757 (N_11757,N_9418,N_7860);
nor U11758 (N_11758,N_8946,N_9248);
or U11759 (N_11759,N_9380,N_9274);
nand U11760 (N_11760,N_8144,N_8393);
nand U11761 (N_11761,N_8982,N_9542);
or U11762 (N_11762,N_8650,N_7751);
and U11763 (N_11763,N_7993,N_8486);
and U11764 (N_11764,N_9464,N_7804);
nand U11765 (N_11765,N_7774,N_7986);
nor U11766 (N_11766,N_7508,N_9953);
nand U11767 (N_11767,N_9554,N_8955);
xor U11768 (N_11768,N_9986,N_9272);
xnor U11769 (N_11769,N_9345,N_8561);
nand U11770 (N_11770,N_8627,N_8704);
nor U11771 (N_11771,N_8579,N_8244);
nor U11772 (N_11772,N_8538,N_9985);
nor U11773 (N_11773,N_9510,N_8948);
or U11774 (N_11774,N_9057,N_8939);
and U11775 (N_11775,N_9863,N_9537);
nor U11776 (N_11776,N_8666,N_8642);
xor U11777 (N_11777,N_8491,N_7729);
or U11778 (N_11778,N_8386,N_8375);
nor U11779 (N_11779,N_8027,N_9086);
or U11780 (N_11780,N_9382,N_8939);
xnor U11781 (N_11781,N_9136,N_9879);
xor U11782 (N_11782,N_7963,N_9734);
and U11783 (N_11783,N_8962,N_9828);
nand U11784 (N_11784,N_9044,N_7800);
and U11785 (N_11785,N_9996,N_8471);
and U11786 (N_11786,N_8543,N_9178);
or U11787 (N_11787,N_8994,N_8362);
nor U11788 (N_11788,N_8136,N_8810);
xor U11789 (N_11789,N_8110,N_9598);
or U11790 (N_11790,N_7530,N_9776);
xor U11791 (N_11791,N_8336,N_8570);
nor U11792 (N_11792,N_8311,N_8702);
xnor U11793 (N_11793,N_7710,N_9669);
or U11794 (N_11794,N_8395,N_9803);
nor U11795 (N_11795,N_8696,N_8452);
nand U11796 (N_11796,N_9726,N_8845);
nand U11797 (N_11797,N_7560,N_8108);
nor U11798 (N_11798,N_8044,N_9070);
and U11799 (N_11799,N_8472,N_8054);
xnor U11800 (N_11800,N_9457,N_9451);
nor U11801 (N_11801,N_9113,N_9397);
or U11802 (N_11802,N_8405,N_9984);
xor U11803 (N_11803,N_7776,N_9506);
nand U11804 (N_11804,N_7907,N_8772);
and U11805 (N_11805,N_8518,N_8629);
and U11806 (N_11806,N_9253,N_9694);
or U11807 (N_11807,N_7993,N_9058);
nand U11808 (N_11808,N_8874,N_7529);
nand U11809 (N_11809,N_8592,N_7936);
or U11810 (N_11810,N_9955,N_8857);
and U11811 (N_11811,N_8202,N_9262);
nor U11812 (N_11812,N_9797,N_7580);
nor U11813 (N_11813,N_9213,N_8279);
xor U11814 (N_11814,N_8268,N_8184);
or U11815 (N_11815,N_9188,N_9226);
nand U11816 (N_11816,N_7911,N_8891);
and U11817 (N_11817,N_9107,N_8587);
xnor U11818 (N_11818,N_9226,N_9183);
and U11819 (N_11819,N_9398,N_9102);
nor U11820 (N_11820,N_9555,N_8702);
nand U11821 (N_11821,N_7506,N_9435);
nor U11822 (N_11822,N_7873,N_8130);
xnor U11823 (N_11823,N_8511,N_7948);
nor U11824 (N_11824,N_9783,N_9996);
and U11825 (N_11825,N_9558,N_8140);
nor U11826 (N_11826,N_8366,N_8145);
and U11827 (N_11827,N_9269,N_9933);
nor U11828 (N_11828,N_8684,N_8139);
and U11829 (N_11829,N_9981,N_8122);
and U11830 (N_11830,N_7626,N_9681);
nand U11831 (N_11831,N_8838,N_9981);
nor U11832 (N_11832,N_8547,N_8667);
xnor U11833 (N_11833,N_9002,N_9270);
nor U11834 (N_11834,N_8933,N_8436);
and U11835 (N_11835,N_8872,N_9093);
xnor U11836 (N_11836,N_9537,N_9023);
or U11837 (N_11837,N_7955,N_9830);
nand U11838 (N_11838,N_8589,N_9659);
nand U11839 (N_11839,N_9728,N_9434);
nor U11840 (N_11840,N_9571,N_9658);
nor U11841 (N_11841,N_8547,N_9006);
xnor U11842 (N_11842,N_7770,N_9849);
nand U11843 (N_11843,N_8894,N_8358);
nor U11844 (N_11844,N_8607,N_8231);
nor U11845 (N_11845,N_9792,N_8019);
or U11846 (N_11846,N_9711,N_8885);
xnor U11847 (N_11847,N_8439,N_8495);
xor U11848 (N_11848,N_7537,N_8785);
xnor U11849 (N_11849,N_7749,N_9642);
or U11850 (N_11850,N_8433,N_8756);
xor U11851 (N_11851,N_7885,N_9788);
nand U11852 (N_11852,N_9857,N_8677);
nand U11853 (N_11853,N_7862,N_7822);
xnor U11854 (N_11854,N_8805,N_7828);
and U11855 (N_11855,N_9650,N_8123);
or U11856 (N_11856,N_8840,N_8910);
nor U11857 (N_11857,N_8758,N_9029);
nand U11858 (N_11858,N_8703,N_9853);
nand U11859 (N_11859,N_7895,N_7558);
or U11860 (N_11860,N_9258,N_7765);
xor U11861 (N_11861,N_8098,N_8908);
nand U11862 (N_11862,N_7744,N_9564);
and U11863 (N_11863,N_8994,N_7738);
and U11864 (N_11864,N_8041,N_9563);
nor U11865 (N_11865,N_8494,N_9967);
nand U11866 (N_11866,N_9628,N_9706);
xnor U11867 (N_11867,N_8844,N_9218);
nand U11868 (N_11868,N_8374,N_8707);
xor U11869 (N_11869,N_9637,N_9349);
or U11870 (N_11870,N_7691,N_8898);
xor U11871 (N_11871,N_8695,N_7893);
xnor U11872 (N_11872,N_8211,N_9463);
nor U11873 (N_11873,N_9492,N_9488);
xor U11874 (N_11874,N_9722,N_9162);
or U11875 (N_11875,N_7546,N_9258);
xnor U11876 (N_11876,N_8598,N_9759);
nand U11877 (N_11877,N_9107,N_9247);
or U11878 (N_11878,N_7891,N_8061);
xor U11879 (N_11879,N_9604,N_8860);
nor U11880 (N_11880,N_8818,N_9672);
xor U11881 (N_11881,N_8210,N_8548);
nand U11882 (N_11882,N_8447,N_8513);
and U11883 (N_11883,N_9019,N_9263);
xor U11884 (N_11884,N_9620,N_7799);
nand U11885 (N_11885,N_9341,N_9839);
and U11886 (N_11886,N_8941,N_9831);
nand U11887 (N_11887,N_9829,N_7594);
and U11888 (N_11888,N_9984,N_9249);
xor U11889 (N_11889,N_8930,N_9388);
xnor U11890 (N_11890,N_8903,N_9713);
or U11891 (N_11891,N_7830,N_8108);
nor U11892 (N_11892,N_7962,N_8622);
nand U11893 (N_11893,N_9145,N_9670);
and U11894 (N_11894,N_9150,N_8032);
nor U11895 (N_11895,N_8880,N_9193);
and U11896 (N_11896,N_9552,N_8567);
and U11897 (N_11897,N_8277,N_8950);
or U11898 (N_11898,N_8723,N_7837);
or U11899 (N_11899,N_7726,N_8664);
and U11900 (N_11900,N_8326,N_7664);
and U11901 (N_11901,N_9118,N_9670);
nand U11902 (N_11902,N_9971,N_8591);
xnor U11903 (N_11903,N_9468,N_8290);
nor U11904 (N_11904,N_8623,N_9157);
and U11905 (N_11905,N_8621,N_9811);
nand U11906 (N_11906,N_8487,N_9804);
nand U11907 (N_11907,N_9921,N_8003);
and U11908 (N_11908,N_9531,N_9175);
xor U11909 (N_11909,N_9314,N_8079);
nand U11910 (N_11910,N_7800,N_7638);
nand U11911 (N_11911,N_7603,N_8373);
xor U11912 (N_11912,N_8900,N_7798);
nand U11913 (N_11913,N_9821,N_9005);
or U11914 (N_11914,N_9446,N_9022);
or U11915 (N_11915,N_8176,N_8719);
or U11916 (N_11916,N_8350,N_9236);
nor U11917 (N_11917,N_9585,N_8546);
nand U11918 (N_11918,N_9785,N_8983);
and U11919 (N_11919,N_9137,N_9893);
or U11920 (N_11920,N_8252,N_8334);
xor U11921 (N_11921,N_8662,N_8835);
xor U11922 (N_11922,N_9753,N_8807);
or U11923 (N_11923,N_8576,N_9667);
xor U11924 (N_11924,N_9027,N_7976);
nor U11925 (N_11925,N_9600,N_7954);
nand U11926 (N_11926,N_9814,N_8229);
nor U11927 (N_11927,N_9093,N_8348);
and U11928 (N_11928,N_8676,N_8546);
xnor U11929 (N_11929,N_9171,N_8540);
or U11930 (N_11930,N_9833,N_9523);
and U11931 (N_11931,N_8576,N_7624);
and U11932 (N_11932,N_9842,N_8702);
and U11933 (N_11933,N_9791,N_9877);
xnor U11934 (N_11934,N_8314,N_9435);
nand U11935 (N_11935,N_8302,N_7579);
or U11936 (N_11936,N_7648,N_7605);
or U11937 (N_11937,N_9719,N_9431);
or U11938 (N_11938,N_8925,N_7641);
or U11939 (N_11939,N_9680,N_7635);
xnor U11940 (N_11940,N_8062,N_7858);
or U11941 (N_11941,N_9114,N_7992);
nor U11942 (N_11942,N_9588,N_7927);
or U11943 (N_11943,N_9919,N_7991);
nor U11944 (N_11944,N_8805,N_9591);
or U11945 (N_11945,N_9032,N_8858);
and U11946 (N_11946,N_8147,N_8066);
or U11947 (N_11947,N_8842,N_9796);
or U11948 (N_11948,N_8386,N_8420);
or U11949 (N_11949,N_8193,N_7752);
and U11950 (N_11950,N_7550,N_9071);
nand U11951 (N_11951,N_9350,N_9688);
or U11952 (N_11952,N_7535,N_9930);
xnor U11953 (N_11953,N_8771,N_9129);
or U11954 (N_11954,N_7645,N_8927);
nand U11955 (N_11955,N_8375,N_8084);
xnor U11956 (N_11956,N_9774,N_8008);
nor U11957 (N_11957,N_9856,N_9448);
nor U11958 (N_11958,N_9753,N_9009);
nand U11959 (N_11959,N_9469,N_9334);
nand U11960 (N_11960,N_9401,N_8285);
nor U11961 (N_11961,N_7843,N_8288);
or U11962 (N_11962,N_7702,N_8386);
or U11963 (N_11963,N_7795,N_9491);
and U11964 (N_11964,N_8574,N_8923);
nand U11965 (N_11965,N_9459,N_9514);
and U11966 (N_11966,N_8522,N_7566);
nand U11967 (N_11967,N_9680,N_9411);
nand U11968 (N_11968,N_9982,N_8594);
nand U11969 (N_11969,N_8053,N_7840);
xor U11970 (N_11970,N_9990,N_7508);
xor U11971 (N_11971,N_7629,N_8839);
nand U11972 (N_11972,N_9720,N_8465);
and U11973 (N_11973,N_9840,N_8747);
nor U11974 (N_11974,N_9300,N_9234);
nand U11975 (N_11975,N_8481,N_9642);
nand U11976 (N_11976,N_8645,N_9394);
xnor U11977 (N_11977,N_7660,N_9271);
nor U11978 (N_11978,N_9037,N_7696);
nor U11979 (N_11979,N_7823,N_8953);
nor U11980 (N_11980,N_8779,N_8205);
nor U11981 (N_11981,N_8094,N_9024);
and U11982 (N_11982,N_8070,N_9297);
xnor U11983 (N_11983,N_7596,N_7939);
nor U11984 (N_11984,N_9398,N_9774);
nor U11985 (N_11985,N_8872,N_8338);
nor U11986 (N_11986,N_7806,N_9153);
and U11987 (N_11987,N_8054,N_7547);
nand U11988 (N_11988,N_9199,N_9275);
nand U11989 (N_11989,N_8112,N_9033);
nand U11990 (N_11990,N_9340,N_7849);
nand U11991 (N_11991,N_8705,N_9743);
nand U11992 (N_11992,N_9648,N_8639);
nand U11993 (N_11993,N_7794,N_7591);
xor U11994 (N_11994,N_7876,N_9727);
or U11995 (N_11995,N_9799,N_8102);
and U11996 (N_11996,N_9955,N_9985);
nor U11997 (N_11997,N_8675,N_9461);
or U11998 (N_11998,N_8318,N_9784);
nor U11999 (N_11999,N_8444,N_7842);
xnor U12000 (N_12000,N_7542,N_7711);
xnor U12001 (N_12001,N_8660,N_7905);
and U12002 (N_12002,N_7790,N_7732);
or U12003 (N_12003,N_8877,N_8796);
or U12004 (N_12004,N_9661,N_8682);
nor U12005 (N_12005,N_9590,N_8849);
nor U12006 (N_12006,N_9756,N_7633);
nor U12007 (N_12007,N_8936,N_8649);
and U12008 (N_12008,N_8513,N_8906);
nand U12009 (N_12009,N_8334,N_7516);
xnor U12010 (N_12010,N_7571,N_8519);
or U12011 (N_12011,N_8924,N_7962);
xor U12012 (N_12012,N_9136,N_8877);
nor U12013 (N_12013,N_9819,N_8132);
nor U12014 (N_12014,N_8172,N_8337);
nor U12015 (N_12015,N_8769,N_8141);
and U12016 (N_12016,N_8007,N_9716);
and U12017 (N_12017,N_7812,N_9898);
and U12018 (N_12018,N_8713,N_8156);
nand U12019 (N_12019,N_9142,N_9362);
nand U12020 (N_12020,N_9536,N_9867);
nand U12021 (N_12021,N_7730,N_9084);
nand U12022 (N_12022,N_8868,N_8287);
nor U12023 (N_12023,N_7656,N_9990);
nor U12024 (N_12024,N_9118,N_8428);
or U12025 (N_12025,N_9934,N_9856);
and U12026 (N_12026,N_8054,N_9256);
nand U12027 (N_12027,N_9642,N_8155);
nand U12028 (N_12028,N_9903,N_7529);
nor U12029 (N_12029,N_8272,N_9142);
or U12030 (N_12030,N_8240,N_7547);
or U12031 (N_12031,N_8101,N_7990);
nor U12032 (N_12032,N_7666,N_7645);
nor U12033 (N_12033,N_8776,N_9148);
or U12034 (N_12034,N_8116,N_7524);
nor U12035 (N_12035,N_8016,N_9896);
nor U12036 (N_12036,N_8270,N_7730);
nand U12037 (N_12037,N_9643,N_8029);
xnor U12038 (N_12038,N_8980,N_8602);
and U12039 (N_12039,N_9859,N_8279);
xor U12040 (N_12040,N_7565,N_7899);
xnor U12041 (N_12041,N_9169,N_9522);
xnor U12042 (N_12042,N_8064,N_9429);
nor U12043 (N_12043,N_8442,N_8628);
xnor U12044 (N_12044,N_7665,N_9285);
nand U12045 (N_12045,N_8441,N_8940);
nor U12046 (N_12046,N_9904,N_9227);
and U12047 (N_12047,N_8041,N_9003);
xor U12048 (N_12048,N_9267,N_9283);
or U12049 (N_12049,N_8124,N_9084);
nor U12050 (N_12050,N_8841,N_9215);
xnor U12051 (N_12051,N_7511,N_8442);
and U12052 (N_12052,N_8425,N_9912);
nor U12053 (N_12053,N_9425,N_8153);
xor U12054 (N_12054,N_7610,N_8866);
and U12055 (N_12055,N_8002,N_8583);
nor U12056 (N_12056,N_8535,N_8206);
or U12057 (N_12057,N_7800,N_9430);
and U12058 (N_12058,N_8251,N_8249);
or U12059 (N_12059,N_8132,N_7882);
xnor U12060 (N_12060,N_9578,N_9892);
and U12061 (N_12061,N_9143,N_9165);
and U12062 (N_12062,N_8561,N_7990);
or U12063 (N_12063,N_9622,N_9458);
nand U12064 (N_12064,N_7787,N_7600);
or U12065 (N_12065,N_8182,N_8205);
xor U12066 (N_12066,N_9630,N_9177);
nor U12067 (N_12067,N_8041,N_8540);
nand U12068 (N_12068,N_8920,N_8967);
xnor U12069 (N_12069,N_8455,N_9378);
nor U12070 (N_12070,N_8175,N_7719);
nor U12071 (N_12071,N_8900,N_8246);
nand U12072 (N_12072,N_9747,N_8976);
nand U12073 (N_12073,N_8083,N_9950);
nand U12074 (N_12074,N_8777,N_8510);
or U12075 (N_12075,N_7943,N_9421);
nand U12076 (N_12076,N_9572,N_7811);
xor U12077 (N_12077,N_7642,N_7623);
or U12078 (N_12078,N_8187,N_9134);
and U12079 (N_12079,N_7803,N_8902);
and U12080 (N_12080,N_9312,N_8792);
or U12081 (N_12081,N_8045,N_8653);
or U12082 (N_12082,N_9611,N_7865);
xnor U12083 (N_12083,N_7504,N_8299);
or U12084 (N_12084,N_9611,N_8295);
or U12085 (N_12085,N_7628,N_8103);
or U12086 (N_12086,N_8956,N_9027);
nand U12087 (N_12087,N_7841,N_9640);
nor U12088 (N_12088,N_9004,N_9593);
xnor U12089 (N_12089,N_9716,N_7682);
xor U12090 (N_12090,N_8387,N_8511);
and U12091 (N_12091,N_7851,N_8037);
xor U12092 (N_12092,N_8037,N_8758);
and U12093 (N_12093,N_8721,N_8154);
nor U12094 (N_12094,N_9817,N_8219);
nand U12095 (N_12095,N_9749,N_9674);
nand U12096 (N_12096,N_7532,N_7924);
nor U12097 (N_12097,N_9775,N_9834);
xor U12098 (N_12098,N_8043,N_9684);
nand U12099 (N_12099,N_9279,N_7640);
nor U12100 (N_12100,N_8401,N_8138);
or U12101 (N_12101,N_7921,N_7851);
or U12102 (N_12102,N_9412,N_8189);
or U12103 (N_12103,N_7796,N_7631);
nand U12104 (N_12104,N_8901,N_8047);
nand U12105 (N_12105,N_7809,N_8149);
xor U12106 (N_12106,N_7980,N_7831);
or U12107 (N_12107,N_9453,N_8430);
xnor U12108 (N_12108,N_8353,N_7634);
nor U12109 (N_12109,N_9249,N_8403);
or U12110 (N_12110,N_9729,N_7934);
and U12111 (N_12111,N_9721,N_7966);
nand U12112 (N_12112,N_8845,N_8294);
or U12113 (N_12113,N_9389,N_7750);
nor U12114 (N_12114,N_9749,N_9281);
and U12115 (N_12115,N_8021,N_8064);
and U12116 (N_12116,N_9323,N_9686);
or U12117 (N_12117,N_8518,N_9376);
and U12118 (N_12118,N_7590,N_9829);
or U12119 (N_12119,N_9511,N_9632);
xnor U12120 (N_12120,N_8145,N_7606);
xor U12121 (N_12121,N_9242,N_8809);
xnor U12122 (N_12122,N_9836,N_9187);
nor U12123 (N_12123,N_8744,N_9023);
or U12124 (N_12124,N_8118,N_9819);
or U12125 (N_12125,N_7536,N_8190);
xnor U12126 (N_12126,N_7680,N_9148);
nand U12127 (N_12127,N_9273,N_9893);
xnor U12128 (N_12128,N_8997,N_8372);
or U12129 (N_12129,N_9357,N_9825);
xor U12130 (N_12130,N_8029,N_8682);
nor U12131 (N_12131,N_9576,N_9323);
and U12132 (N_12132,N_7651,N_7917);
nor U12133 (N_12133,N_9506,N_9962);
nand U12134 (N_12134,N_8458,N_9529);
xor U12135 (N_12135,N_9038,N_9024);
and U12136 (N_12136,N_9564,N_9687);
or U12137 (N_12137,N_8058,N_9528);
xnor U12138 (N_12138,N_7939,N_8793);
nor U12139 (N_12139,N_8521,N_9920);
or U12140 (N_12140,N_9153,N_8937);
and U12141 (N_12141,N_9363,N_8811);
or U12142 (N_12142,N_9453,N_8392);
or U12143 (N_12143,N_8048,N_9928);
xnor U12144 (N_12144,N_9384,N_8200);
and U12145 (N_12145,N_9872,N_9896);
xor U12146 (N_12146,N_7658,N_9582);
xnor U12147 (N_12147,N_7660,N_8487);
nand U12148 (N_12148,N_8057,N_8260);
and U12149 (N_12149,N_8060,N_9917);
nand U12150 (N_12150,N_7954,N_9751);
xor U12151 (N_12151,N_8043,N_9061);
nand U12152 (N_12152,N_9300,N_9657);
xor U12153 (N_12153,N_9614,N_8563);
or U12154 (N_12154,N_9051,N_8382);
xnor U12155 (N_12155,N_9082,N_9298);
nand U12156 (N_12156,N_9387,N_8813);
and U12157 (N_12157,N_7957,N_8171);
and U12158 (N_12158,N_9337,N_7825);
and U12159 (N_12159,N_7638,N_9859);
nand U12160 (N_12160,N_9895,N_8069);
nand U12161 (N_12161,N_8341,N_8222);
and U12162 (N_12162,N_8272,N_9141);
or U12163 (N_12163,N_8398,N_9534);
xnor U12164 (N_12164,N_8624,N_9987);
nor U12165 (N_12165,N_8921,N_7503);
xor U12166 (N_12166,N_9884,N_8475);
nand U12167 (N_12167,N_9255,N_8100);
nand U12168 (N_12168,N_9548,N_8091);
and U12169 (N_12169,N_7892,N_9280);
and U12170 (N_12170,N_7518,N_8632);
or U12171 (N_12171,N_8882,N_8111);
nand U12172 (N_12172,N_8083,N_9642);
or U12173 (N_12173,N_9794,N_7760);
nand U12174 (N_12174,N_9841,N_8182);
and U12175 (N_12175,N_9035,N_8050);
nor U12176 (N_12176,N_8318,N_7523);
xnor U12177 (N_12177,N_7876,N_9189);
xor U12178 (N_12178,N_8137,N_7846);
nor U12179 (N_12179,N_9540,N_9734);
nand U12180 (N_12180,N_8063,N_8126);
xnor U12181 (N_12181,N_8713,N_9348);
or U12182 (N_12182,N_9135,N_9839);
xnor U12183 (N_12183,N_9476,N_8321);
or U12184 (N_12184,N_7592,N_8144);
and U12185 (N_12185,N_9094,N_9701);
xor U12186 (N_12186,N_9934,N_8875);
nand U12187 (N_12187,N_8704,N_9358);
and U12188 (N_12188,N_8129,N_9547);
or U12189 (N_12189,N_9604,N_9192);
and U12190 (N_12190,N_9298,N_8547);
xor U12191 (N_12191,N_9978,N_9725);
nand U12192 (N_12192,N_7559,N_7571);
xnor U12193 (N_12193,N_9718,N_9794);
or U12194 (N_12194,N_8634,N_7619);
xor U12195 (N_12195,N_9117,N_9079);
and U12196 (N_12196,N_8627,N_7891);
or U12197 (N_12197,N_8886,N_9489);
xor U12198 (N_12198,N_8980,N_7634);
xnor U12199 (N_12199,N_7513,N_7623);
and U12200 (N_12200,N_7504,N_8036);
nand U12201 (N_12201,N_8943,N_8625);
or U12202 (N_12202,N_8251,N_7648);
and U12203 (N_12203,N_8124,N_8421);
or U12204 (N_12204,N_9224,N_7618);
nand U12205 (N_12205,N_7569,N_8855);
nor U12206 (N_12206,N_9826,N_8437);
xor U12207 (N_12207,N_9199,N_9336);
or U12208 (N_12208,N_9120,N_8574);
nand U12209 (N_12209,N_8929,N_7873);
nand U12210 (N_12210,N_7597,N_8904);
nand U12211 (N_12211,N_9567,N_9626);
or U12212 (N_12212,N_8925,N_9005);
or U12213 (N_12213,N_8926,N_7790);
nor U12214 (N_12214,N_8114,N_8787);
nor U12215 (N_12215,N_8587,N_9650);
or U12216 (N_12216,N_9614,N_7831);
xnor U12217 (N_12217,N_9320,N_7725);
or U12218 (N_12218,N_8557,N_9545);
and U12219 (N_12219,N_9273,N_8921);
xor U12220 (N_12220,N_7938,N_8548);
and U12221 (N_12221,N_9725,N_7837);
nand U12222 (N_12222,N_8098,N_9832);
xor U12223 (N_12223,N_8369,N_7834);
nor U12224 (N_12224,N_8272,N_8836);
nor U12225 (N_12225,N_7528,N_8592);
or U12226 (N_12226,N_9966,N_8040);
xor U12227 (N_12227,N_8645,N_7976);
or U12228 (N_12228,N_9443,N_8866);
and U12229 (N_12229,N_7697,N_9512);
xor U12230 (N_12230,N_8814,N_8570);
nand U12231 (N_12231,N_7718,N_8850);
and U12232 (N_12232,N_8374,N_8603);
nand U12233 (N_12233,N_7599,N_9833);
nor U12234 (N_12234,N_9737,N_9940);
nor U12235 (N_12235,N_9486,N_9677);
or U12236 (N_12236,N_9255,N_8433);
nand U12237 (N_12237,N_9643,N_9255);
or U12238 (N_12238,N_9613,N_9606);
or U12239 (N_12239,N_7716,N_8561);
or U12240 (N_12240,N_9382,N_7870);
xor U12241 (N_12241,N_7706,N_8623);
and U12242 (N_12242,N_9950,N_9902);
and U12243 (N_12243,N_8892,N_9356);
and U12244 (N_12244,N_8577,N_8370);
xor U12245 (N_12245,N_8351,N_7893);
xnor U12246 (N_12246,N_8068,N_9128);
and U12247 (N_12247,N_8503,N_8230);
nor U12248 (N_12248,N_8561,N_9962);
or U12249 (N_12249,N_8200,N_8478);
nand U12250 (N_12250,N_8184,N_9586);
xor U12251 (N_12251,N_8278,N_8799);
nor U12252 (N_12252,N_7501,N_9185);
xor U12253 (N_12253,N_8148,N_7541);
nand U12254 (N_12254,N_8177,N_9352);
xor U12255 (N_12255,N_8299,N_8909);
nand U12256 (N_12256,N_8849,N_8789);
xor U12257 (N_12257,N_8443,N_9946);
or U12258 (N_12258,N_8624,N_9597);
nand U12259 (N_12259,N_7794,N_9966);
or U12260 (N_12260,N_9934,N_8158);
nand U12261 (N_12261,N_8605,N_7970);
xor U12262 (N_12262,N_9133,N_9963);
or U12263 (N_12263,N_8982,N_8901);
nor U12264 (N_12264,N_9955,N_8889);
nor U12265 (N_12265,N_9395,N_8334);
and U12266 (N_12266,N_9454,N_8464);
nor U12267 (N_12267,N_8427,N_9033);
xnor U12268 (N_12268,N_8530,N_9071);
nand U12269 (N_12269,N_9774,N_9189);
or U12270 (N_12270,N_8322,N_9154);
nor U12271 (N_12271,N_7721,N_9435);
and U12272 (N_12272,N_9416,N_9740);
nand U12273 (N_12273,N_8808,N_8931);
nor U12274 (N_12274,N_7899,N_8993);
and U12275 (N_12275,N_9160,N_8615);
or U12276 (N_12276,N_7559,N_8226);
and U12277 (N_12277,N_9384,N_9852);
xnor U12278 (N_12278,N_9774,N_8347);
nand U12279 (N_12279,N_8088,N_7609);
xor U12280 (N_12280,N_7520,N_9813);
or U12281 (N_12281,N_9212,N_8005);
or U12282 (N_12282,N_9622,N_7964);
nor U12283 (N_12283,N_9175,N_7559);
and U12284 (N_12284,N_9053,N_9962);
xor U12285 (N_12285,N_8744,N_9082);
xnor U12286 (N_12286,N_8841,N_7813);
nand U12287 (N_12287,N_7523,N_8995);
or U12288 (N_12288,N_9842,N_8259);
nand U12289 (N_12289,N_8750,N_9551);
nand U12290 (N_12290,N_9974,N_8520);
or U12291 (N_12291,N_9631,N_7664);
or U12292 (N_12292,N_8915,N_8207);
and U12293 (N_12293,N_8784,N_8036);
nor U12294 (N_12294,N_7907,N_9025);
nand U12295 (N_12295,N_9347,N_8161);
nand U12296 (N_12296,N_9186,N_7763);
nor U12297 (N_12297,N_7845,N_9186);
nand U12298 (N_12298,N_7821,N_8774);
xnor U12299 (N_12299,N_9442,N_8722);
nand U12300 (N_12300,N_8843,N_9548);
nand U12301 (N_12301,N_8899,N_7999);
xnor U12302 (N_12302,N_8031,N_8100);
and U12303 (N_12303,N_7731,N_7626);
and U12304 (N_12304,N_9185,N_9103);
nor U12305 (N_12305,N_8987,N_9388);
xor U12306 (N_12306,N_8706,N_9425);
xnor U12307 (N_12307,N_7676,N_9537);
nor U12308 (N_12308,N_8482,N_9439);
or U12309 (N_12309,N_9452,N_8801);
nor U12310 (N_12310,N_8370,N_9222);
xor U12311 (N_12311,N_8041,N_8480);
and U12312 (N_12312,N_9751,N_9452);
and U12313 (N_12313,N_7571,N_9015);
nor U12314 (N_12314,N_8752,N_7632);
nor U12315 (N_12315,N_9009,N_8951);
xor U12316 (N_12316,N_8522,N_9539);
xnor U12317 (N_12317,N_9811,N_9438);
nor U12318 (N_12318,N_9979,N_8438);
nand U12319 (N_12319,N_8772,N_9789);
nor U12320 (N_12320,N_8123,N_8936);
nor U12321 (N_12321,N_9009,N_9590);
and U12322 (N_12322,N_8740,N_8887);
nand U12323 (N_12323,N_8824,N_9262);
and U12324 (N_12324,N_8099,N_8398);
nand U12325 (N_12325,N_9520,N_8671);
and U12326 (N_12326,N_8157,N_9146);
nand U12327 (N_12327,N_9078,N_9810);
xnor U12328 (N_12328,N_8057,N_8817);
nand U12329 (N_12329,N_9529,N_9639);
nand U12330 (N_12330,N_7909,N_9429);
or U12331 (N_12331,N_8451,N_8803);
nor U12332 (N_12332,N_7909,N_9732);
or U12333 (N_12333,N_7800,N_7786);
xor U12334 (N_12334,N_8698,N_9622);
or U12335 (N_12335,N_8520,N_9100);
nor U12336 (N_12336,N_8040,N_8970);
nand U12337 (N_12337,N_8556,N_9222);
and U12338 (N_12338,N_9735,N_7518);
or U12339 (N_12339,N_8879,N_8129);
and U12340 (N_12340,N_8001,N_8046);
xor U12341 (N_12341,N_7566,N_9407);
and U12342 (N_12342,N_9607,N_8768);
nand U12343 (N_12343,N_9976,N_9634);
and U12344 (N_12344,N_9066,N_8198);
xnor U12345 (N_12345,N_8826,N_8060);
and U12346 (N_12346,N_8823,N_8305);
and U12347 (N_12347,N_8854,N_9865);
and U12348 (N_12348,N_7772,N_8038);
nor U12349 (N_12349,N_8834,N_8477);
nand U12350 (N_12350,N_8937,N_7773);
nor U12351 (N_12351,N_7638,N_8834);
xor U12352 (N_12352,N_8040,N_8793);
nand U12353 (N_12353,N_8001,N_9284);
and U12354 (N_12354,N_8449,N_9652);
nor U12355 (N_12355,N_9128,N_8669);
or U12356 (N_12356,N_9456,N_8891);
xor U12357 (N_12357,N_8283,N_8527);
nand U12358 (N_12358,N_7714,N_8851);
or U12359 (N_12359,N_9912,N_8083);
nor U12360 (N_12360,N_8259,N_9160);
or U12361 (N_12361,N_7604,N_8262);
xor U12362 (N_12362,N_8936,N_7617);
or U12363 (N_12363,N_8264,N_8286);
or U12364 (N_12364,N_7932,N_9626);
or U12365 (N_12365,N_8132,N_8300);
or U12366 (N_12366,N_8199,N_7530);
nand U12367 (N_12367,N_7900,N_8481);
and U12368 (N_12368,N_9624,N_8804);
nand U12369 (N_12369,N_9646,N_9023);
nor U12370 (N_12370,N_8566,N_7609);
xnor U12371 (N_12371,N_8552,N_9978);
and U12372 (N_12372,N_9364,N_8937);
nand U12373 (N_12373,N_8453,N_8691);
nand U12374 (N_12374,N_8005,N_7606);
nand U12375 (N_12375,N_8940,N_9157);
or U12376 (N_12376,N_8903,N_7823);
nand U12377 (N_12377,N_7945,N_9104);
nor U12378 (N_12378,N_9378,N_8969);
nor U12379 (N_12379,N_8978,N_8949);
or U12380 (N_12380,N_9449,N_9356);
nor U12381 (N_12381,N_7918,N_9781);
and U12382 (N_12382,N_9073,N_9636);
nor U12383 (N_12383,N_8247,N_8621);
or U12384 (N_12384,N_8454,N_7862);
nand U12385 (N_12385,N_7610,N_7763);
and U12386 (N_12386,N_9105,N_9950);
xnor U12387 (N_12387,N_7612,N_9630);
xnor U12388 (N_12388,N_9036,N_8267);
nand U12389 (N_12389,N_9891,N_9654);
nor U12390 (N_12390,N_9531,N_9595);
or U12391 (N_12391,N_7907,N_7731);
nand U12392 (N_12392,N_9517,N_8983);
nand U12393 (N_12393,N_9894,N_9963);
nor U12394 (N_12394,N_9309,N_8167);
and U12395 (N_12395,N_7655,N_8430);
or U12396 (N_12396,N_7601,N_9622);
nand U12397 (N_12397,N_8358,N_9986);
nor U12398 (N_12398,N_9364,N_7661);
xnor U12399 (N_12399,N_8376,N_8601);
nor U12400 (N_12400,N_9094,N_8645);
nand U12401 (N_12401,N_8608,N_8124);
or U12402 (N_12402,N_9699,N_9340);
nor U12403 (N_12403,N_8020,N_7722);
xor U12404 (N_12404,N_9919,N_8934);
xor U12405 (N_12405,N_9735,N_9823);
or U12406 (N_12406,N_9004,N_9788);
xor U12407 (N_12407,N_9943,N_9729);
or U12408 (N_12408,N_8340,N_8253);
and U12409 (N_12409,N_9997,N_8984);
and U12410 (N_12410,N_7986,N_7963);
and U12411 (N_12411,N_9744,N_8592);
nand U12412 (N_12412,N_8421,N_8474);
or U12413 (N_12413,N_9208,N_8166);
nor U12414 (N_12414,N_9459,N_9771);
nor U12415 (N_12415,N_8407,N_9257);
nor U12416 (N_12416,N_8466,N_8235);
and U12417 (N_12417,N_9836,N_9760);
nand U12418 (N_12418,N_8966,N_9532);
and U12419 (N_12419,N_7639,N_7539);
or U12420 (N_12420,N_9730,N_9684);
and U12421 (N_12421,N_8049,N_8118);
or U12422 (N_12422,N_7563,N_8447);
and U12423 (N_12423,N_9155,N_9303);
nand U12424 (N_12424,N_9568,N_9787);
xnor U12425 (N_12425,N_9437,N_8795);
and U12426 (N_12426,N_8539,N_9559);
xor U12427 (N_12427,N_7847,N_8026);
xor U12428 (N_12428,N_8896,N_9611);
or U12429 (N_12429,N_9100,N_8453);
nor U12430 (N_12430,N_7644,N_8793);
nor U12431 (N_12431,N_8047,N_9013);
xor U12432 (N_12432,N_8656,N_8266);
nand U12433 (N_12433,N_9609,N_9576);
nand U12434 (N_12434,N_9744,N_8195);
nand U12435 (N_12435,N_9434,N_8080);
xnor U12436 (N_12436,N_9627,N_9118);
or U12437 (N_12437,N_8612,N_8315);
xor U12438 (N_12438,N_8253,N_9919);
nor U12439 (N_12439,N_8063,N_9961);
or U12440 (N_12440,N_7635,N_7649);
xor U12441 (N_12441,N_9550,N_9736);
nand U12442 (N_12442,N_7634,N_9856);
or U12443 (N_12443,N_8972,N_9206);
nor U12444 (N_12444,N_7607,N_9800);
nand U12445 (N_12445,N_8534,N_8770);
nand U12446 (N_12446,N_8340,N_9521);
and U12447 (N_12447,N_8086,N_8788);
and U12448 (N_12448,N_7633,N_8773);
nor U12449 (N_12449,N_7504,N_8332);
nand U12450 (N_12450,N_9688,N_8691);
or U12451 (N_12451,N_8347,N_7733);
nand U12452 (N_12452,N_9896,N_9990);
or U12453 (N_12453,N_9559,N_7535);
xor U12454 (N_12454,N_9758,N_8518);
xor U12455 (N_12455,N_8927,N_8344);
or U12456 (N_12456,N_9982,N_9186);
xnor U12457 (N_12457,N_7885,N_7999);
nor U12458 (N_12458,N_9372,N_7618);
or U12459 (N_12459,N_7843,N_8133);
and U12460 (N_12460,N_9215,N_7718);
or U12461 (N_12461,N_7880,N_8187);
and U12462 (N_12462,N_9588,N_8962);
nand U12463 (N_12463,N_7513,N_9782);
or U12464 (N_12464,N_9320,N_7564);
nand U12465 (N_12465,N_9487,N_7646);
xor U12466 (N_12466,N_8180,N_9701);
and U12467 (N_12467,N_9595,N_7907);
xor U12468 (N_12468,N_7527,N_8318);
and U12469 (N_12469,N_8181,N_9798);
nand U12470 (N_12470,N_7612,N_9479);
nor U12471 (N_12471,N_8849,N_9272);
nand U12472 (N_12472,N_7966,N_9776);
xor U12473 (N_12473,N_7703,N_8528);
xor U12474 (N_12474,N_7910,N_7633);
and U12475 (N_12475,N_9360,N_8997);
nand U12476 (N_12476,N_9973,N_8550);
and U12477 (N_12477,N_8186,N_9887);
or U12478 (N_12478,N_8730,N_7520);
xor U12479 (N_12479,N_9164,N_8010);
nand U12480 (N_12480,N_9721,N_9976);
or U12481 (N_12481,N_7962,N_9876);
xnor U12482 (N_12482,N_8197,N_9939);
or U12483 (N_12483,N_7730,N_9838);
nand U12484 (N_12484,N_7536,N_9185);
nand U12485 (N_12485,N_9851,N_8633);
nand U12486 (N_12486,N_9482,N_9325);
nand U12487 (N_12487,N_8033,N_8910);
nor U12488 (N_12488,N_7550,N_8233);
nand U12489 (N_12489,N_9364,N_8230);
nand U12490 (N_12490,N_8365,N_9133);
or U12491 (N_12491,N_8230,N_9957);
nor U12492 (N_12492,N_8966,N_8162);
or U12493 (N_12493,N_8650,N_9425);
nor U12494 (N_12494,N_9050,N_9003);
or U12495 (N_12495,N_9925,N_9021);
xor U12496 (N_12496,N_9060,N_8648);
nor U12497 (N_12497,N_9952,N_9192);
nand U12498 (N_12498,N_9226,N_8124);
or U12499 (N_12499,N_8191,N_8814);
nor U12500 (N_12500,N_11155,N_10023);
nand U12501 (N_12501,N_10414,N_10848);
xor U12502 (N_12502,N_11133,N_12024);
nor U12503 (N_12503,N_10521,N_10867);
or U12504 (N_12504,N_10174,N_10100);
nand U12505 (N_12505,N_11860,N_11895);
nor U12506 (N_12506,N_11753,N_10253);
xor U12507 (N_12507,N_11379,N_11115);
or U12508 (N_12508,N_11444,N_11593);
and U12509 (N_12509,N_12127,N_11058);
and U12510 (N_12510,N_11701,N_11461);
or U12511 (N_12511,N_10643,N_12368);
or U12512 (N_12512,N_11838,N_11498);
nor U12513 (N_12513,N_10520,N_12421);
nand U12514 (N_12514,N_10494,N_10468);
nor U12515 (N_12515,N_11523,N_10540);
or U12516 (N_12516,N_11845,N_11198);
and U12517 (N_12517,N_10908,N_12443);
and U12518 (N_12518,N_12359,N_11485);
xor U12519 (N_12519,N_10961,N_11512);
and U12520 (N_12520,N_11104,N_11316);
and U12521 (N_12521,N_11026,N_10072);
xnor U12522 (N_12522,N_12075,N_10065);
nor U12523 (N_12523,N_10877,N_11965);
and U12524 (N_12524,N_12477,N_12398);
nand U12525 (N_12525,N_10423,N_11029);
or U12526 (N_12526,N_10478,N_12200);
and U12527 (N_12527,N_10706,N_11415);
or U12528 (N_12528,N_11466,N_12006);
xnor U12529 (N_12529,N_10671,N_10500);
or U12530 (N_12530,N_12470,N_10452);
xnor U12531 (N_12531,N_12099,N_10792);
nor U12532 (N_12532,N_10568,N_12390);
nor U12533 (N_12533,N_11399,N_11047);
xnor U12534 (N_12534,N_10497,N_11916);
nor U12535 (N_12535,N_10873,N_10167);
xor U12536 (N_12536,N_10129,N_11188);
nor U12537 (N_12537,N_12343,N_10831);
and U12538 (N_12538,N_12394,N_11468);
nand U12539 (N_12539,N_12197,N_11050);
or U12540 (N_12540,N_10888,N_10070);
xor U12541 (N_12541,N_11849,N_10721);
or U12542 (N_12542,N_11140,N_10110);
nand U12543 (N_12543,N_10524,N_12320);
nor U12544 (N_12544,N_10829,N_11728);
or U12545 (N_12545,N_12045,N_10291);
xnor U12546 (N_12546,N_10281,N_10959);
nor U12547 (N_12547,N_11241,N_11378);
nor U12548 (N_12548,N_12439,N_10410);
nor U12549 (N_12549,N_10240,N_10482);
and U12550 (N_12550,N_11550,N_10034);
xor U12551 (N_12551,N_11715,N_10418);
xor U12552 (N_12552,N_12466,N_12034);
nand U12553 (N_12553,N_11305,N_10089);
nor U12554 (N_12554,N_11724,N_10196);
xnor U12555 (N_12555,N_11108,N_12212);
xor U12556 (N_12556,N_12057,N_12152);
xor U12557 (N_12557,N_11835,N_11999);
xor U12558 (N_12558,N_10736,N_11095);
nor U12559 (N_12559,N_11689,N_11488);
xor U12560 (N_12560,N_11346,N_11322);
nand U12561 (N_12561,N_12358,N_11688);
and U12562 (N_12562,N_10631,N_11417);
and U12563 (N_12563,N_11056,N_11237);
or U12564 (N_12564,N_11479,N_11912);
nand U12565 (N_12565,N_10723,N_10910);
nor U12566 (N_12566,N_11165,N_11635);
or U12567 (N_12567,N_10224,N_11000);
xor U12568 (N_12568,N_10286,N_12108);
nand U12569 (N_12569,N_12076,N_10903);
nor U12570 (N_12570,N_10173,N_11214);
or U12571 (N_12571,N_10639,N_12277);
nor U12572 (N_12572,N_10632,N_12300);
or U12573 (N_12573,N_11362,N_11252);
nand U12574 (N_12574,N_12445,N_11347);
and U12575 (N_12575,N_10691,N_11159);
xnor U12576 (N_12576,N_10672,N_12220);
nand U12577 (N_12577,N_10475,N_12309);
or U12578 (N_12578,N_10162,N_10476);
and U12579 (N_12579,N_11310,N_11220);
and U12580 (N_12580,N_11424,N_10607);
and U12581 (N_12581,N_11385,N_10301);
xnor U12582 (N_12582,N_12077,N_10629);
xor U12583 (N_12583,N_10579,N_10298);
and U12584 (N_12584,N_10587,N_11693);
or U12585 (N_12585,N_12037,N_12064);
or U12586 (N_12586,N_12178,N_10597);
nor U12587 (N_12587,N_11117,N_12475);
or U12588 (N_12588,N_10765,N_10287);
nand U12589 (N_12589,N_11678,N_11568);
and U12590 (N_12590,N_12317,N_10821);
and U12591 (N_12591,N_10443,N_10726);
nand U12592 (N_12592,N_10337,N_10036);
xnor U12593 (N_12593,N_10472,N_11672);
or U12594 (N_12594,N_11492,N_10285);
and U12595 (N_12595,N_11869,N_10318);
xor U12596 (N_12596,N_12248,N_12216);
xnor U12597 (N_12597,N_11826,N_10803);
or U12598 (N_12598,N_10398,N_12088);
nand U12599 (N_12599,N_12464,N_11705);
nor U12600 (N_12600,N_12177,N_12459);
nand U12601 (N_12601,N_10202,N_10455);
xnor U12602 (N_12602,N_11010,N_10709);
and U12603 (N_12603,N_10391,N_10633);
and U12604 (N_12604,N_11832,N_11273);
or U12605 (N_12605,N_10514,N_11756);
nor U12606 (N_12606,N_11407,N_11991);
and U12607 (N_12607,N_10053,N_10615);
xor U12608 (N_12608,N_11719,N_11784);
and U12609 (N_12609,N_10471,N_11189);
xor U12610 (N_12610,N_10872,N_12314);
and U12611 (N_12611,N_12379,N_10113);
and U12612 (N_12612,N_12257,N_12245);
nor U12613 (N_12613,N_10772,N_11565);
nor U12614 (N_12614,N_10256,N_11878);
xnor U12615 (N_12615,N_12307,N_10499);
xnor U12616 (N_12616,N_11883,N_10662);
and U12617 (N_12617,N_12051,N_11011);
and U12618 (N_12618,N_11298,N_10433);
or U12619 (N_12619,N_12079,N_10866);
nor U12620 (N_12620,N_11994,N_11998);
and U12621 (N_12621,N_10536,N_10740);
or U12622 (N_12622,N_12308,N_10451);
nand U12623 (N_12623,N_11259,N_11797);
and U12624 (N_12624,N_11937,N_10095);
or U12625 (N_12625,N_11540,N_10506);
xor U12626 (N_12626,N_11277,N_11044);
xor U12627 (N_12627,N_10182,N_11266);
xnor U12628 (N_12628,N_10642,N_10421);
nor U12629 (N_12629,N_11004,N_10109);
xor U12630 (N_12630,N_10555,N_10751);
nor U12631 (N_12631,N_11588,N_12346);
xor U12632 (N_12632,N_10832,N_12080);
xor U12633 (N_12633,N_10128,N_12322);
nor U12634 (N_12634,N_11284,N_10450);
or U12635 (N_12635,N_10377,N_10355);
xor U12636 (N_12636,N_11100,N_11644);
nand U12637 (N_12637,N_11828,N_10952);
nor U12638 (N_12638,N_12162,N_10339);
or U12639 (N_12639,N_11702,N_10878);
xor U12640 (N_12640,N_11889,N_10766);
xnor U12641 (N_12641,N_11369,N_11027);
nor U12642 (N_12642,N_12053,N_10558);
xor U12643 (N_12643,N_10650,N_11008);
nand U12644 (N_12644,N_10134,N_10094);
nor U12645 (N_12645,N_11203,N_10950);
and U12646 (N_12646,N_11321,N_10796);
and U12647 (N_12647,N_11223,N_11146);
nor U12648 (N_12648,N_12066,N_12395);
nand U12649 (N_12649,N_11748,N_10327);
xor U12650 (N_12650,N_10243,N_12331);
and U12651 (N_12651,N_11939,N_11367);
and U12652 (N_12652,N_10120,N_12310);
xnor U12653 (N_12653,N_11830,N_10146);
nand U12654 (N_12654,N_10739,N_11254);
or U12655 (N_12655,N_11548,N_10170);
xor U12656 (N_12656,N_11616,N_11098);
or U12657 (N_12657,N_11012,N_10058);
and U12658 (N_12658,N_10016,N_12371);
xnor U12659 (N_12659,N_12411,N_10371);
or U12660 (N_12660,N_10933,N_12240);
nand U12661 (N_12661,N_12166,N_11422);
nand U12662 (N_12662,N_12402,N_12494);
and U12663 (N_12663,N_12260,N_11981);
or U12664 (N_12664,N_11038,N_10075);
nor U12665 (N_12665,N_12000,N_11506);
nand U12666 (N_12666,N_12446,N_11647);
or U12667 (N_12667,N_11920,N_10782);
and U12668 (N_12668,N_10229,N_10913);
nand U12669 (N_12669,N_10851,N_11013);
and U12670 (N_12670,N_12004,N_12087);
nand U12671 (N_12671,N_11018,N_12335);
and U12672 (N_12672,N_11571,N_10673);
nor U12673 (N_12673,N_11197,N_10649);
and U12674 (N_12674,N_12126,N_11881);
xor U12675 (N_12675,N_11914,N_11729);
nor U12676 (N_12676,N_10150,N_10336);
and U12677 (N_12677,N_11561,N_10352);
and U12678 (N_12678,N_12265,N_10080);
nand U12679 (N_12679,N_11410,N_12497);
nor U12680 (N_12680,N_11125,N_11544);
and U12681 (N_12681,N_11552,N_10039);
and U12682 (N_12682,N_10571,N_11216);
or U12683 (N_12683,N_11211,N_11674);
nand U12684 (N_12684,N_10530,N_10083);
nand U12685 (N_12685,N_10117,N_11199);
nor U12686 (N_12686,N_10144,N_12151);
or U12687 (N_12687,N_10131,N_12280);
nor U12688 (N_12688,N_12097,N_11128);
xnor U12689 (N_12689,N_10787,N_10988);
xnor U12690 (N_12690,N_12058,N_11037);
nand U12691 (N_12691,N_10984,N_11208);
or U12692 (N_12692,N_11196,N_10460);
and U12693 (N_12693,N_10600,N_11777);
or U12694 (N_12694,N_10618,N_12254);
nor U12695 (N_12695,N_10152,N_11345);
and U12696 (N_12696,N_11077,N_12128);
nor U12697 (N_12697,N_11687,N_10528);
nand U12698 (N_12698,N_10802,N_11755);
nor U12699 (N_12699,N_11969,N_10975);
nor U12700 (N_12700,N_12025,N_11185);
xnor U12701 (N_12701,N_11684,N_12154);
nor U12702 (N_12702,N_12067,N_11080);
xor U12703 (N_12703,N_10572,N_11781);
xor U12704 (N_12704,N_11767,N_11068);
xor U12705 (N_12705,N_10047,N_10955);
and U12706 (N_12706,N_10981,N_12454);
and U12707 (N_12707,N_12124,N_11853);
xnor U12708 (N_12708,N_10936,N_10546);
and U12709 (N_12709,N_11288,N_11726);
nor U12710 (N_12710,N_11820,N_10362);
or U12711 (N_12711,N_12388,N_12062);
and U12712 (N_12712,N_11886,N_11352);
nor U12713 (N_12713,N_12050,N_12451);
or U12714 (N_12714,N_10727,N_11441);
nand U12715 (N_12715,N_10771,N_11390);
nor U12716 (N_12716,N_10860,N_11107);
or U12717 (N_12717,N_10824,N_10960);
xnor U12718 (N_12718,N_11624,N_12341);
and U12719 (N_12719,N_11111,N_10680);
or U12720 (N_12720,N_10864,N_11792);
or U12721 (N_12721,N_10653,N_10003);
xnor U12722 (N_12722,N_10177,N_12195);
or U12723 (N_12723,N_10595,N_11015);
xnor U12724 (N_12724,N_11944,N_12206);
or U12725 (N_12725,N_12173,N_11537);
xnor U12726 (N_12726,N_12374,N_10998);
or U12727 (N_12727,N_10021,N_10176);
nand U12728 (N_12728,N_10325,N_12082);
xnor U12729 (N_12729,N_10416,N_12137);
nand U12730 (N_12730,N_11289,N_10805);
xor U12731 (N_12731,N_10799,N_11127);
nand U12732 (N_12732,N_11502,N_11081);
and U12733 (N_12733,N_10665,N_10891);
nand U12734 (N_12734,N_11679,N_11698);
and U12735 (N_12735,N_10332,N_12493);
nand U12736 (N_12736,N_10985,N_10508);
or U12737 (N_12737,N_11236,N_11727);
nand U12738 (N_12738,N_12488,N_11360);
nor U12739 (N_12739,N_11434,N_11594);
nand U12740 (N_12740,N_11180,N_11141);
and U12741 (N_12741,N_10326,N_10097);
or U12742 (N_12742,N_10213,N_12179);
nand U12743 (N_12743,N_10310,N_11609);
and U12744 (N_12744,N_11657,N_10742);
and U12745 (N_12745,N_10349,N_10221);
nor U12746 (N_12746,N_11151,N_11435);
and U12747 (N_12747,N_12301,N_11694);
xor U12748 (N_12748,N_10406,N_10348);
and U12749 (N_12749,N_10785,N_10601);
nand U12750 (N_12750,N_10092,N_10096);
xnor U12751 (N_12751,N_10823,N_11733);
nor U12752 (N_12752,N_12121,N_10931);
nand U12753 (N_12753,N_10188,N_10350);
or U12754 (N_12754,N_10901,N_11928);
xor U12755 (N_12755,N_11903,N_12263);
or U12756 (N_12756,N_12271,N_10598);
nand U12757 (N_12757,N_11480,N_11613);
or U12758 (N_12758,N_10522,N_11306);
xnor U12759 (N_12759,N_12040,N_10695);
nor U12760 (N_12760,N_11612,N_10390);
nand U12761 (N_12761,N_10809,N_10504);
or U12762 (N_12762,N_12396,N_11822);
and U12763 (N_12763,N_11737,N_12141);
or U12764 (N_12764,N_11618,N_10470);
nor U12765 (N_12765,N_11639,N_10214);
nor U12766 (N_12766,N_11952,N_11195);
and U12767 (N_12767,N_10532,N_11400);
nor U12768 (N_12768,N_11675,N_10011);
or U12769 (N_12769,N_11487,N_11516);
and U12770 (N_12770,N_11365,N_11072);
xnor U12771 (N_12771,N_12408,N_11167);
and U12772 (N_12772,N_11774,N_11597);
nand U12773 (N_12773,N_12242,N_12336);
and U12774 (N_12774,N_12274,N_10582);
xnor U12775 (N_12775,N_10543,N_12420);
nor U12776 (N_12776,N_12273,N_10741);
xor U12777 (N_12777,N_11780,N_11403);
and U12778 (N_12778,N_12223,N_11476);
nand U12779 (N_12779,N_10290,N_11414);
nor U12780 (N_12780,N_11619,N_10657);
nand U12781 (N_12781,N_10605,N_11730);
or U12782 (N_12782,N_10538,N_12354);
xnor U12783 (N_12783,N_10000,N_10289);
nor U12784 (N_12784,N_12019,N_12232);
nand U12785 (N_12785,N_11515,N_11779);
xor U12786 (N_12786,N_10263,N_10825);
nand U12787 (N_12787,N_10063,N_11874);
and U12788 (N_12788,N_10602,N_10667);
xnor U12789 (N_12789,N_11739,N_10820);
or U12790 (N_12790,N_12023,N_11655);
or U12791 (N_12791,N_12282,N_10446);
or U12792 (N_12792,N_12455,N_10502);
or U12793 (N_12793,N_11919,N_10028);
or U12794 (N_12794,N_10516,N_11174);
nand U12795 (N_12795,N_10485,N_10437);
or U12796 (N_12796,N_11086,N_12095);
and U12797 (N_12797,N_11228,N_10067);
and U12798 (N_12798,N_12284,N_10335);
xnor U12799 (N_12799,N_10160,N_12172);
xnor U12800 (N_12800,N_10217,N_10868);
and U12801 (N_12801,N_12204,N_10424);
or U12802 (N_12802,N_11328,N_11771);
nor U12803 (N_12803,N_11173,N_11268);
and U12804 (N_12804,N_10195,N_10885);
nand U12805 (N_12805,N_10486,N_11901);
or U12806 (N_12806,N_10135,N_11793);
and U12807 (N_12807,N_10774,N_11551);
and U12808 (N_12808,N_11930,N_11202);
and U12809 (N_12809,N_11484,N_12109);
nor U12810 (N_12810,N_10581,N_11610);
nand U12811 (N_12811,N_10231,N_12258);
xnor U12812 (N_12812,N_10123,N_12054);
xnor U12813 (N_12813,N_10505,N_11885);
or U12814 (N_12814,N_12430,N_10951);
xnor U12815 (N_12815,N_12083,N_11045);
and U12816 (N_12816,N_11136,N_11114);
xnor U12817 (N_12817,N_10139,N_11307);
xnor U12818 (N_12818,N_12068,N_11640);
xor U12819 (N_12819,N_10957,N_11314);
or U12820 (N_12820,N_11253,N_11430);
or U12821 (N_12821,N_10899,N_10790);
nor U12822 (N_12822,N_10022,N_10085);
nand U12823 (N_12823,N_12409,N_11723);
or U12824 (N_12824,N_10495,N_10140);
or U12825 (N_12825,N_10259,N_10190);
and U12826 (N_12826,N_11409,N_10839);
or U12827 (N_12827,N_10939,N_10778);
nand U12828 (N_12828,N_10840,N_12165);
xor U12829 (N_12829,N_10679,N_10200);
or U12830 (N_12830,N_12191,N_10019);
or U12831 (N_12831,N_10404,N_10165);
xnor U12832 (N_12832,N_10449,N_10013);
and U12833 (N_12833,N_11227,N_11564);
and U12834 (N_12834,N_12189,N_11162);
xor U12835 (N_12835,N_11384,N_11852);
and U12836 (N_12836,N_11255,N_11866);
nor U12837 (N_12837,N_10315,N_10842);
nand U12838 (N_12838,N_11245,N_11718);
nand U12839 (N_12839,N_10748,N_10225);
and U12840 (N_12840,N_11576,N_12246);
nor U12841 (N_12841,N_12462,N_12495);
xor U12842 (N_12842,N_11495,N_12298);
nand U12843 (N_12843,N_11170,N_11653);
nor U12844 (N_12844,N_10261,N_11156);
nand U12845 (N_12845,N_12442,N_11622);
nor U12846 (N_12846,N_10490,N_10941);
and U12847 (N_12847,N_10386,N_10590);
xor U12848 (N_12848,N_11311,N_10852);
and U12849 (N_12849,N_11789,N_10454);
nor U12850 (N_12850,N_11521,N_11926);
or U12851 (N_12851,N_11201,N_11582);
or U12852 (N_12852,N_10054,N_12176);
and U12853 (N_12853,N_11962,N_10242);
or U12854 (N_12854,N_10324,N_10970);
and U12855 (N_12855,N_10826,N_10252);
or U12856 (N_12856,N_10668,N_10991);
xnor U12857 (N_12857,N_10218,N_12171);
or U12858 (N_12858,N_10312,N_11121);
xor U12859 (N_12859,N_11749,N_11842);
xor U12860 (N_12860,N_11645,N_10007);
or U12861 (N_12861,N_11342,N_10853);
and U12862 (N_12862,N_10834,N_11317);
nand U12863 (N_12863,N_10453,N_11992);
and U12864 (N_12864,N_11530,N_11848);
and U12865 (N_12865,N_11925,N_12044);
and U12866 (N_12866,N_10719,N_12028);
or U12867 (N_12867,N_10978,N_10122);
xor U12868 (N_12868,N_11813,N_11017);
or U12869 (N_12869,N_12407,N_11932);
nor U12870 (N_12870,N_10645,N_11910);
nand U12871 (N_12871,N_12306,N_10353);
nor U12872 (N_12872,N_10258,N_10030);
nand U12873 (N_12873,N_12429,N_11534);
nand U12874 (N_12874,N_11039,N_12016);
and U12875 (N_12875,N_10277,N_12149);
nand U12876 (N_12876,N_11810,N_10690);
or U12877 (N_12877,N_10609,N_10702);
nor U12878 (N_12878,N_12366,N_12432);
nor U12879 (N_12879,N_11806,N_10479);
or U12880 (N_12880,N_11043,N_11088);
nand U12881 (N_12881,N_11865,N_12334);
or U12882 (N_12882,N_11945,N_12198);
and U12883 (N_12883,N_10967,N_12404);
nand U12884 (N_12884,N_10330,N_10375);
nor U12885 (N_12885,N_10576,N_10964);
and U12886 (N_12886,N_11335,N_11979);
xor U12887 (N_12887,N_10574,N_11032);
nand U12888 (N_12888,N_11176,N_10425);
and U12889 (N_12889,N_11898,N_10807);
nand U12890 (N_12890,N_11758,N_10725);
nor U12891 (N_12891,N_11851,N_11704);
nand U12892 (N_12892,N_12086,N_11595);
nor U12893 (N_12893,N_11711,N_10205);
nand U12894 (N_12894,N_11396,N_11833);
nand U12895 (N_12895,N_12303,N_11243);
and U12896 (N_12896,N_12030,N_12382);
and U12897 (N_12897,N_11145,N_10280);
nand U12898 (N_12898,N_10111,N_11264);
nor U12899 (N_12899,N_11683,N_12218);
or U12900 (N_12900,N_11531,N_11230);
nand U12901 (N_12901,N_12405,N_10535);
xor U12902 (N_12902,N_11831,N_12069);
or U12903 (N_12903,N_12499,N_10812);
xnor U12904 (N_12904,N_12412,N_10227);
nor U12905 (N_12905,N_11235,N_10930);
xor U12906 (N_12906,N_11073,N_11389);
and U12907 (N_12907,N_12210,N_11493);
and U12908 (N_12908,N_11605,N_10661);
and U12909 (N_12909,N_10886,N_10493);
and U12910 (N_12910,N_10971,N_11292);
or U12911 (N_12911,N_12196,N_10008);
or U12912 (N_12912,N_12315,N_11968);
and U12913 (N_12913,N_10808,N_12113);
nor U12914 (N_12914,N_11249,N_10026);
or U12915 (N_12915,N_11269,N_12281);
nor U12916 (N_12916,N_11517,N_10343);
and U12917 (N_12917,N_11248,N_12117);
and U12918 (N_12918,N_11099,N_11840);
nand U12919 (N_12919,N_11818,N_10363);
xor U12920 (N_12920,N_10064,N_10753);
nor U12921 (N_12921,N_10014,N_10874);
and U12922 (N_12922,N_11611,N_11160);
nor U12923 (N_12923,N_11929,N_11750);
nor U12924 (N_12924,N_10948,N_10760);
and U12925 (N_12925,N_12479,N_11168);
or U12926 (N_12926,N_10382,N_11329);
xor U12927 (N_12927,N_11261,N_10299);
xnor U12928 (N_12928,N_10005,N_10862);
xnor U12929 (N_12929,N_10338,N_12392);
nand U12930 (N_12930,N_11420,N_10237);
or U12931 (N_12931,N_11184,N_12125);
nor U12932 (N_12932,N_10038,N_10436);
and U12933 (N_12933,N_11313,N_11633);
or U12934 (N_12934,N_10688,N_10119);
xnor U12935 (N_12935,N_11035,N_12283);
nor U12936 (N_12936,N_12349,N_10551);
or U12937 (N_12937,N_10077,N_10800);
and U12938 (N_12938,N_10814,N_10518);
and U12939 (N_12939,N_12342,N_10015);
or U12940 (N_12940,N_12406,N_12249);
nand U12941 (N_12941,N_10399,N_11112);
nand U12942 (N_12942,N_11814,N_10447);
xnor U12943 (N_12943,N_12226,N_12410);
xnor U12944 (N_12944,N_11557,N_12202);
nand U12945 (N_12945,N_10488,N_10627);
and U12946 (N_12946,N_11083,N_12397);
xor U12947 (N_12947,N_10296,N_10513);
or U12948 (N_12948,N_11798,N_10223);
or U12949 (N_12949,N_12393,N_12375);
xnor U12950 (N_12950,N_10611,N_10062);
nor U12951 (N_12951,N_10898,N_11584);
nand U12952 (N_12952,N_10676,N_10033);
and U12953 (N_12953,N_12434,N_10917);
xor U12954 (N_12954,N_12001,N_12483);
xnor U12955 (N_12955,N_12188,N_11232);
nand U12956 (N_12956,N_11532,N_11631);
nand U12957 (N_12957,N_10902,N_11690);
or U12958 (N_12958,N_12175,N_11376);
nand U12959 (N_12959,N_11880,N_12463);
nor U12960 (N_12960,N_11258,N_12319);
nand U12961 (N_12961,N_12471,N_10798);
nor U12962 (N_12962,N_10239,N_10469);
nor U12963 (N_12963,N_11486,N_10278);
nor U12964 (N_12964,N_12444,N_11303);
nand U12965 (N_12965,N_12078,N_11129);
xnor U12966 (N_12966,N_10919,N_10703);
and U12967 (N_12967,N_10845,N_11786);
and U12968 (N_12968,N_10481,N_10457);
xor U12969 (N_12969,N_11953,N_11747);
nor U12970 (N_12970,N_10523,N_11995);
and U12971 (N_12971,N_11547,N_10857);
and U12972 (N_12972,N_11082,N_11955);
xnor U12973 (N_12973,N_10757,N_11087);
or U12974 (N_12974,N_12328,N_12187);
xor U12975 (N_12975,N_11442,N_11790);
and U12976 (N_12976,N_11134,N_10204);
xnor U12977 (N_12977,N_10344,N_11431);
or U12978 (N_12978,N_11796,N_11001);
or U12979 (N_12979,N_10735,N_11787);
xnor U12980 (N_12980,N_12116,N_11783);
nor U12981 (N_12981,N_11101,N_12452);
xnor U12982 (N_12982,N_10491,N_10145);
nand U12983 (N_12983,N_11902,N_12422);
nor U12984 (N_12984,N_11652,N_10704);
nand U12985 (N_12985,N_11106,N_12266);
nor U12986 (N_12986,N_10731,N_12160);
and U12987 (N_12987,N_10996,N_10103);
nor U12988 (N_12988,N_10730,N_11364);
or U12989 (N_12989,N_11332,N_10752);
or U12990 (N_12990,N_10619,N_11036);
or U12991 (N_12991,N_11319,N_11200);
xnor U12992 (N_12992,N_11391,N_11666);
or U12993 (N_12993,N_11935,N_11807);
or U12994 (N_12994,N_11872,N_10701);
or U12995 (N_12995,N_11918,N_10138);
nor U12996 (N_12996,N_12145,N_11710);
nand U12997 (N_12997,N_12238,N_10905);
nand U12998 (N_12998,N_11546,N_12474);
nand U12999 (N_12999,N_11413,N_11663);
or U13000 (N_13000,N_11425,N_12481);
nor U13001 (N_13001,N_10376,N_11028);
and U13002 (N_13002,N_12272,N_11857);
nand U13003 (N_13003,N_11559,N_10439);
nor U13004 (N_13004,N_11827,N_11630);
nor U13005 (N_13005,N_11716,N_10461);
nor U13006 (N_13006,N_10250,N_12143);
or U13007 (N_13007,N_12457,N_12377);
and U13008 (N_13008,N_12465,N_10945);
or U13009 (N_13009,N_12180,N_11281);
xnor U13010 (N_13010,N_10664,N_10958);
and U13011 (N_13011,N_10419,N_11648);
nor U13012 (N_13012,N_11875,N_11394);
or U13013 (N_13013,N_11344,N_11246);
nor U13014 (N_13014,N_12041,N_12456);
nor U13015 (N_13015,N_12056,N_10098);
xnor U13016 (N_13016,N_11966,N_11016);
or U13017 (N_13017,N_12098,N_11397);
nand U13018 (N_13018,N_11089,N_11302);
or U13019 (N_13019,N_10604,N_10401);
or U13020 (N_13020,N_11988,N_10463);
and U13021 (N_13021,N_11069,N_12168);
or U13022 (N_13022,N_12026,N_10300);
or U13023 (N_13023,N_10358,N_10309);
xor U13024 (N_13024,N_10801,N_11590);
and U13025 (N_13025,N_10329,N_11859);
xor U13026 (N_13026,N_10927,N_11731);
nand U13027 (N_13027,N_11300,N_10341);
nor U13028 (N_13028,N_11494,N_11229);
and U13029 (N_13029,N_11060,N_11250);
xor U13030 (N_13030,N_11971,N_12021);
xnor U13031 (N_13031,N_12440,N_10887);
nor U13032 (N_13032,N_10351,N_11144);
nand U13033 (N_13033,N_10010,N_10086);
xnor U13034 (N_13034,N_11242,N_11641);
nand U13035 (N_13035,N_10172,N_11408);
nand U13036 (N_13036,N_11061,N_10032);
xnor U13037 (N_13037,N_10394,N_11805);
and U13038 (N_13038,N_12476,N_10232);
nand U13039 (N_13039,N_11967,N_11118);
nand U13040 (N_13040,N_12033,N_12352);
or U13041 (N_13041,N_10669,N_10686);
and U13042 (N_13042,N_10552,N_11308);
and U13043 (N_13043,N_10271,N_11572);
xor U13044 (N_13044,N_10819,N_11393);
xnor U13045 (N_13045,N_10219,N_11183);
nand U13046 (N_13046,N_11518,N_12369);
nor U13047 (N_13047,N_10302,N_11153);
nand U13048 (N_13048,N_11163,N_10987);
and U13049 (N_13049,N_10194,N_11138);
nand U13050 (N_13050,N_11947,N_11556);
or U13051 (N_13051,N_11964,N_10179);
and U13052 (N_13052,N_11280,N_11186);
nor U13053 (N_13053,N_11251,N_10198);
nor U13054 (N_13054,N_12449,N_10187);
xnor U13055 (N_13055,N_10420,N_10512);
and U13056 (N_13056,N_11986,N_10562);
nor U13057 (N_13057,N_10046,N_10185);
nand U13058 (N_13058,N_11990,N_11583);
nand U13059 (N_13059,N_12262,N_10384);
nor U13060 (N_13060,N_11856,N_10817);
xor U13061 (N_13061,N_12059,N_11339);
and U13062 (N_13062,N_10681,N_11501);
xnor U13063 (N_13063,N_11513,N_10559);
and U13064 (N_13064,N_10746,N_10804);
and U13065 (N_13065,N_10159,N_12423);
and U13066 (N_13066,N_10603,N_11267);
or U13067 (N_13067,N_12122,N_11368);
nand U13068 (N_13068,N_11412,N_11536);
xnor U13069 (N_13069,N_11897,N_11987);
xor U13070 (N_13070,N_12092,N_10417);
and U13071 (N_13071,N_11941,N_10659);
nor U13072 (N_13072,N_11525,N_10265);
xor U13073 (N_13073,N_12381,N_11474);
and U13074 (N_13074,N_10136,N_10045);
xnor U13075 (N_13075,N_12047,N_11766);
and U13076 (N_13076,N_10379,N_12340);
and U13077 (N_13077,N_11664,N_12387);
and U13078 (N_13078,N_11464,N_12115);
and U13079 (N_13079,N_11950,N_12365);
or U13080 (N_13080,N_10870,N_12135);
xor U13081 (N_13081,N_11132,N_12046);
or U13082 (N_13082,N_12485,N_12362);
nand U13083 (N_13083,N_11071,N_11740);
nand U13084 (N_13084,N_11404,N_12299);
xnor U13085 (N_13085,N_11634,N_11218);
nor U13086 (N_13086,N_10319,N_11074);
xnor U13087 (N_13087,N_12461,N_11888);
and U13088 (N_13088,N_10636,N_11963);
nand U13089 (N_13089,N_10056,N_10477);
nand U13090 (N_13090,N_11324,N_11437);
or U13091 (N_13091,N_11057,N_10606);
nor U13092 (N_13092,N_12032,N_12247);
nand U13093 (N_13093,N_10938,N_11142);
or U13094 (N_13094,N_12304,N_11327);
or U13095 (N_13095,N_10986,N_12012);
nand U13096 (N_13096,N_11179,N_11921);
nor U13097 (N_13097,N_10126,N_10374);
and U13098 (N_13098,N_11497,N_11119);
and U13099 (N_13099,N_11383,N_11650);
xor U13100 (N_13100,N_10613,N_10308);
nand U13101 (N_13101,N_11421,N_10728);
nand U13102 (N_13102,N_12219,N_12294);
or U13103 (N_13103,N_10115,N_11542);
or U13104 (N_13104,N_11225,N_11019);
nor U13105 (N_13105,N_10282,N_10462);
xnor U13106 (N_13106,N_10369,N_11312);
and U13107 (N_13107,N_10793,N_10354);
xor U13108 (N_13108,N_11432,N_12424);
xor U13109 (N_13109,N_10548,N_10954);
nor U13110 (N_13110,N_10983,N_10169);
nand U13111 (N_13111,N_11465,N_10429);
nand U13112 (N_13112,N_10025,N_11846);
xnor U13113 (N_13113,N_12293,N_12373);
nand U13114 (N_13114,N_11959,N_10674);
or U13115 (N_13115,N_12385,N_11938);
nor U13116 (N_13116,N_10953,N_12438);
and U13117 (N_13117,N_11993,N_11006);
nor U13118 (N_13118,N_11470,N_10228);
nand U13119 (N_13119,N_10048,N_12170);
nor U13120 (N_13120,N_11560,N_10132);
nand U13121 (N_13121,N_12433,N_11110);
and U13122 (N_13122,N_11122,N_10614);
nand U13123 (N_13123,N_12261,N_10594);
and U13124 (N_13124,N_11735,N_10322);
xor U13125 (N_13125,N_10775,N_11528);
and U13126 (N_13126,N_11102,N_11014);
nand U13127 (N_13127,N_10539,N_10368);
nand U13128 (N_13128,N_11439,N_10212);
or U13129 (N_13129,N_10037,N_11206);
nor U13130 (N_13130,N_11263,N_11481);
and U13131 (N_13131,N_11182,N_11440);
and U13132 (N_13132,N_11854,N_10297);
xor U13133 (N_13133,N_11398,N_10810);
or U13134 (N_13134,N_11535,N_11699);
and U13135 (N_13135,N_11714,N_12091);
nand U13136 (N_13136,N_10199,N_10440);
nor U13137 (N_13137,N_10272,N_10737);
xnor U13138 (N_13138,N_12090,N_11773);
and U13139 (N_13139,N_12148,N_11040);
or U13140 (N_13140,N_10969,N_11894);
or U13141 (N_13141,N_11725,N_11181);
xnor U13142 (N_13142,N_11309,N_11778);
and U13143 (N_13143,N_12042,N_12049);
xnor U13144 (N_13144,N_11580,N_10722);
or U13145 (N_13145,N_10527,N_11983);
xor U13146 (N_13146,N_11529,N_10087);
xnor U13147 (N_13147,N_10052,N_11091);
and U13148 (N_13148,N_10178,N_12235);
or U13149 (N_13149,N_12129,N_11062);
and U13150 (N_13150,N_10906,N_11649);
xnor U13151 (N_13151,N_10155,N_10525);
xnor U13152 (N_13152,N_10141,N_11450);
nor U13153 (N_13153,N_12130,N_11052);
and U13154 (N_13154,N_11785,N_12017);
nor U13155 (N_13155,N_12185,N_10402);
xor U13156 (N_13156,N_11911,N_11913);
or U13157 (N_13157,N_12061,N_10161);
xor U13158 (N_13158,N_10876,N_11053);
and U13159 (N_13159,N_10544,N_10400);
nand U13160 (N_13160,N_10541,N_11685);
xnor U13161 (N_13161,N_11152,N_11761);
nor U13162 (N_13162,N_11712,N_11446);
or U13163 (N_13163,N_11627,N_11997);
or U13164 (N_13164,N_11333,N_10846);
xor U13165 (N_13165,N_10158,N_11262);
xor U13166 (N_13166,N_10677,N_12389);
nor U13167 (N_13167,N_11330,N_12435);
nand U13168 (N_13168,N_10397,N_10593);
or U13169 (N_13169,N_11638,N_10881);
or U13170 (N_13170,N_11489,N_10275);
nand U13171 (N_13171,N_10738,N_11116);
xor U13172 (N_13172,N_10101,N_11617);
and U13173 (N_13173,N_12351,N_12380);
and U13174 (N_13174,N_11763,N_11989);
nor U13175 (N_13175,N_10156,N_10473);
and U13176 (N_13176,N_12330,N_10806);
and U13177 (N_13177,N_12103,N_11504);
xor U13178 (N_13178,N_12250,N_10102);
nand U13179 (N_13179,N_11054,N_10623);
or U13180 (N_13180,N_10626,N_12278);
or U13181 (N_13181,N_10537,N_11591);
or U13182 (N_13182,N_10762,N_11667);
nor U13183 (N_13183,N_12230,N_11917);
and U13184 (N_13184,N_10533,N_10492);
nor U13185 (N_13185,N_11923,N_10884);
and U13186 (N_13186,N_11996,N_11387);
nor U13187 (N_13187,N_12448,N_10783);
and U13188 (N_13188,N_11337,N_10646);
or U13189 (N_13189,N_11975,N_12020);
or U13190 (N_13190,N_10779,N_11794);
xor U13191 (N_13191,N_10389,N_11658);
or U13192 (N_13192,N_11873,N_11769);
or U13193 (N_13193,N_10168,N_11570);
nand U13194 (N_13194,N_10018,N_11059);
or U13195 (N_13195,N_10578,N_10181);
nand U13196 (N_13196,N_12234,N_11802);
and U13197 (N_13197,N_12425,N_11503);
nand U13198 (N_13198,N_12428,N_10699);
or U13199 (N_13199,N_10550,N_10995);
or U13200 (N_13200,N_10251,N_11841);
or U13201 (N_13201,N_10307,N_11864);
nand U13202 (N_13202,N_11460,N_11762);
nand U13203 (N_13203,N_10480,N_10711);
nor U13204 (N_13204,N_12264,N_10584);
and U13205 (N_13205,N_11469,N_12181);
or U13206 (N_13206,N_11175,N_10640);
and U13207 (N_13207,N_12201,N_10118);
xor U13208 (N_13208,N_10255,N_12081);
nand U13209 (N_13209,N_10154,N_10922);
or U13210 (N_13210,N_11244,N_10434);
nor U13211 (N_13211,N_12207,N_10001);
xnor U13212 (N_13212,N_10108,N_11816);
or U13213 (N_13213,N_11418,N_10438);
nand U13214 (N_13214,N_10912,N_11172);
nor U13215 (N_13215,N_10426,N_10747);
or U13216 (N_13216,N_11867,N_11178);
nor U13217 (N_13217,N_11380,N_11219);
nor U13218 (N_13218,N_10393,N_11192);
nor U13219 (N_13219,N_10515,N_10896);
nor U13220 (N_13220,N_11585,N_11215);
nand U13221 (N_13221,N_10929,N_11187);
or U13222 (N_13222,N_10345,N_11428);
and U13223 (N_13223,N_10099,N_12236);
or U13224 (N_13224,N_10942,N_11686);
nand U13225 (N_13225,N_10260,N_10830);
and U13226 (N_13226,N_11003,N_11980);
and U13227 (N_13227,N_11351,N_12071);
nand U13228 (N_13228,N_11651,N_11021);
xnor U13229 (N_13229,N_10051,N_10153);
xnor U13230 (N_13230,N_11299,N_11934);
or U13231 (N_13231,N_10074,N_11297);
or U13232 (N_13232,N_10763,N_12490);
or U13233 (N_13233,N_12347,N_10427);
and U13234 (N_13234,N_10982,N_10445);
and U13235 (N_13235,N_11795,N_10180);
and U13236 (N_13236,N_12084,N_11765);
nand U13237 (N_13237,N_10002,N_11586);
xnor U13238 (N_13238,N_10777,N_12450);
or U13239 (N_13239,N_11668,N_11221);
or U13240 (N_13240,N_10586,N_12227);
or U13241 (N_13241,N_11850,N_11799);
or U13242 (N_13242,N_11957,N_11922);
xnor U13243 (N_13243,N_11217,N_11757);
nand U13244 (N_13244,N_10850,N_10569);
nor U13245 (N_13245,N_11320,N_10781);
xor U13246 (N_13246,N_12164,N_10836);
nor U13247 (N_13247,N_11348,N_11030);
and U13248 (N_13248,N_10624,N_10334);
and U13249 (N_13249,N_10407,N_10565);
nand U13250 (N_13250,N_11707,N_12043);
xnor U13251 (N_13251,N_11543,N_11363);
and U13252 (N_13252,N_10422,N_11909);
xor U13253 (N_13253,N_11373,N_11782);
or U13254 (N_13254,N_10784,N_12114);
and U13255 (N_13255,N_12367,N_12253);
nand U13256 (N_13256,N_11131,N_10313);
and U13257 (N_13257,N_11154,N_11477);
nor U13258 (N_13258,N_10321,N_12399);
nor U13259 (N_13259,N_12085,N_10926);
nor U13260 (N_13260,N_12478,N_11554);
nor U13261 (N_13261,N_12391,N_11887);
and U13262 (N_13262,N_11721,N_12208);
nand U13263 (N_13263,N_10789,N_12100);
nand U13264 (N_13264,N_11366,N_10192);
and U13265 (N_13265,N_10106,N_10459);
nand U13266 (N_13266,N_11751,N_11809);
and U13267 (N_13267,N_10222,N_10621);
nand U13268 (N_13268,N_11812,N_12120);
and U13269 (N_13269,N_10685,N_10648);
nor U13270 (N_13270,N_11563,N_11109);
nor U13271 (N_13271,N_12296,N_11065);
nor U13272 (N_13272,N_12400,N_10235);
or U13273 (N_13273,N_10822,N_10088);
nand U13274 (N_13274,N_11411,N_12018);
and U13275 (N_13275,N_12101,N_12159);
xor U13276 (N_13276,N_12332,N_11356);
nand U13277 (N_13277,N_10768,N_10889);
or U13278 (N_13278,N_11193,N_10127);
and U13279 (N_13279,N_11596,N_10588);
or U13280 (N_13280,N_10510,N_10432);
nor U13281 (N_13281,N_10163,N_10655);
or U13282 (N_13282,N_12311,N_10380);
xnor U13283 (N_13283,N_12106,N_10041);
xor U13284 (N_13284,N_11448,N_12318);
or U13285 (N_13285,N_11084,N_10915);
nand U13286 (N_13286,N_10284,N_11603);
nor U13287 (N_13287,N_10408,N_12498);
xor U13288 (N_13288,N_10316,N_11207);
xor U13289 (N_13289,N_12417,N_10055);
xor U13290 (N_13290,N_12286,N_10547);
xnor U13291 (N_13291,N_10698,N_10556);
or U13292 (N_13292,N_10684,N_10732);
nand U13293 (N_13293,N_11713,N_11304);
nand U13294 (N_13294,N_10892,N_12241);
nor U13295 (N_13295,N_12297,N_12403);
nor U13296 (N_13296,N_10017,N_11164);
nand U13297 (N_13297,N_10818,N_12138);
or U13298 (N_13298,N_12468,N_12229);
and U13299 (N_13299,N_10211,N_12372);
nand U13300 (N_13300,N_11355,N_12123);
xnor U13301 (N_13301,N_11113,N_12183);
and U13302 (N_13302,N_12144,N_10435);
nor U13303 (N_13303,N_10940,N_11372);
nor U13304 (N_13304,N_11738,N_10233);
nor U13305 (N_13305,N_11406,N_12146);
nor U13306 (N_13306,N_11843,N_10773);
nand U13307 (N_13307,N_10976,N_10043);
nor U13308 (N_13308,N_12473,N_12279);
xor U13309 (N_13309,N_12376,N_10755);
and U13310 (N_13310,N_10909,N_10246);
xor U13311 (N_13311,N_11628,N_10081);
and U13312 (N_13312,N_10564,N_10758);
nor U13313 (N_13313,N_11600,N_12224);
nand U13314 (N_13314,N_12142,N_11524);
nor U13315 (N_13315,N_12312,N_12111);
nor U13316 (N_13316,N_10776,N_11978);
nor U13317 (N_13317,N_10612,N_10184);
and U13318 (N_13318,N_11478,N_11205);
nor U13319 (N_13319,N_11906,N_10356);
or U13320 (N_13320,N_11499,N_12094);
and U13321 (N_13321,N_12039,N_12252);
and U13322 (N_13322,N_10591,N_10687);
nand U13323 (N_13323,N_10935,N_10531);
xnor U13324 (N_13324,N_12487,N_10894);
nand U13325 (N_13325,N_11904,N_12169);
or U13326 (N_13326,N_11670,N_10828);
and U13327 (N_13327,N_10795,N_11876);
or U13328 (N_13328,N_10616,N_12256);
and U13329 (N_13329,N_11671,N_12337);
nand U13330 (N_13330,N_11148,N_10143);
or U13331 (N_13331,N_11931,N_11078);
nand U13332 (N_13332,N_11323,N_11770);
or U13333 (N_13333,N_10268,N_12383);
and U13334 (N_13334,N_10236,N_10230);
nand U13335 (N_13335,N_10266,N_10932);
nor U13336 (N_13336,N_11042,N_11575);
and U13337 (N_13337,N_10644,N_11533);
and U13338 (N_13338,N_12131,N_11943);
nor U13339 (N_13339,N_10360,N_11419);
or U13340 (N_13340,N_10359,N_10811);
xor U13341 (N_13341,N_11659,N_11927);
nand U13342 (N_13342,N_12276,N_11009);
and U13343 (N_13343,N_10770,N_10678);
nor U13344 (N_13344,N_10718,N_10561);
nand U13345 (N_13345,N_10142,N_12437);
nand U13346 (N_13346,N_10720,N_10295);
and U13347 (N_13347,N_10331,N_10367);
and U13348 (N_13348,N_11291,N_12110);
xnor U13349 (N_13349,N_11287,N_10412);
xor U13350 (N_13350,N_12350,N_11985);
nand U13351 (N_13351,N_10880,N_10928);
nand U13352 (N_13352,N_11510,N_12013);
nor U13353 (N_13353,N_10164,N_10947);
nor U13354 (N_13354,N_10415,N_11462);
xor U13355 (N_13355,N_10079,N_11276);
and U13356 (N_13356,N_10378,N_12480);
nand U13357 (N_13357,N_11157,N_11958);
and U13358 (N_13358,N_10835,N_10317);
xor U13359 (N_13359,N_12364,N_11539);
or U13360 (N_13360,N_10756,N_11844);
or U13361 (N_13361,N_11381,N_11046);
and U13362 (N_13362,N_10583,N_12415);
nand U13363 (N_13363,N_12291,N_10764);
and U13364 (N_13364,N_12492,N_11815);
xnor U13365 (N_13365,N_11210,N_10666);
nor U13366 (N_13366,N_10914,N_12401);
or U13367 (N_13367,N_10361,N_10511);
or U13368 (N_13368,N_12011,N_10637);
or U13369 (N_13369,N_10883,N_10107);
xnor U13370 (N_13370,N_10871,N_11490);
xor U13371 (N_13371,N_10157,N_10467);
nor U13372 (N_13372,N_12386,N_11746);
and U13373 (N_13373,N_12031,N_12213);
nand U13374 (N_13374,N_12270,N_10381);
nor U13375 (N_13375,N_11891,N_12288);
nand U13376 (N_13376,N_10501,N_11388);
and U13377 (N_13377,N_11334,N_10916);
or U13378 (N_13378,N_10149,N_12305);
xnor U13379 (N_13379,N_11625,N_12093);
xnor U13380 (N_13380,N_10675,N_11285);
nor U13381 (N_13381,N_10897,N_11224);
or U13382 (N_13382,N_11491,N_10311);
nor U13383 (N_13383,N_12209,N_12027);
nor U13384 (N_13384,N_11942,N_10241);
nor U13385 (N_13385,N_12484,N_10980);
and U13386 (N_13386,N_11022,N_11438);
nand U13387 (N_13387,N_11374,N_11070);
or U13388 (N_13388,N_11423,N_10567);
or U13389 (N_13389,N_10946,N_11954);
or U13390 (N_13390,N_11656,N_11956);
nor U13391 (N_13391,N_11899,N_11169);
nor U13392 (N_13392,N_10713,N_10403);
xnor U13393 (N_13393,N_10697,N_12222);
xnor U13394 (N_13394,N_12089,N_11933);
nand U13395 (N_13395,N_11924,N_10847);
nor U13396 (N_13396,N_11341,N_10890);
nand U13397 (N_13397,N_10193,N_10570);
nand U13398 (N_13398,N_11507,N_11884);
and U13399 (N_13399,N_12194,N_11602);
and U13400 (N_13400,N_10733,N_10797);
or U13401 (N_13401,N_10040,N_12107);
or U13402 (N_13402,N_11282,N_11260);
nand U13403 (N_13403,N_11598,N_11336);
and U13404 (N_13404,N_12215,N_10274);
and U13405 (N_13405,N_11034,N_11676);
and U13406 (N_13406,N_11296,N_11680);
or U13407 (N_13407,N_10059,N_12313);
and U13408 (N_13408,N_12353,N_11075);
nor U13409 (N_13409,N_11452,N_12156);
or U13410 (N_13410,N_10049,N_11092);
and U13411 (N_13411,N_10734,N_10208);
nor U13412 (N_13412,N_11984,N_10956);
nor U13413 (N_13413,N_10105,N_10465);
nand U13414 (N_13414,N_11511,N_12038);
and U13415 (N_13415,N_12472,N_11265);
and U13416 (N_13416,N_10875,N_12255);
xnor U13417 (N_13417,N_12112,N_10992);
or U13418 (N_13418,N_11433,N_10431);
or U13419 (N_13419,N_10882,N_11661);
xnor U13420 (N_13420,N_11948,N_11982);
or U13421 (N_13421,N_10201,N_11692);
nor U13422 (N_13422,N_10288,N_12199);
or U13423 (N_13423,N_10340,N_12302);
nor U13424 (N_13424,N_10148,N_11977);
nor U13425 (N_13425,N_12102,N_10166);
xnor U13426 (N_13426,N_11824,N_10788);
nand U13427 (N_13427,N_11274,N_12186);
or U13428 (N_13428,N_10977,N_12015);
nor U13429 (N_13429,N_10305,N_11436);
or U13430 (N_13430,N_11213,N_10215);
nor U13431 (N_13431,N_10635,N_12356);
xor U13432 (N_13432,N_10428,N_12295);
and U13433 (N_13433,N_11601,N_11256);
or U13434 (N_13434,N_10444,N_12416);
nor U13435 (N_13435,N_10396,N_11861);
or U13436 (N_13436,N_10342,N_11278);
and U13437 (N_13437,N_10585,N_11821);
nor U13438 (N_13438,N_11871,N_11562);
xor U13439 (N_13439,N_10689,N_12285);
and U13440 (N_13440,N_10973,N_11722);
nor U13441 (N_13441,N_11623,N_10273);
nor U13442 (N_13442,N_10966,N_12489);
xnor U13443 (N_13443,N_10745,N_11147);
nand U13444 (N_13444,N_11177,N_11063);
and U13445 (N_13445,N_11343,N_12345);
xnor U13446 (N_13446,N_10294,N_11458);
nand U13447 (N_13447,N_10474,N_11161);
nor U13448 (N_13448,N_11457,N_12447);
and U13449 (N_13449,N_11896,N_11094);
nand U13450 (N_13450,N_11836,N_11545);
or U13451 (N_13451,N_11326,N_11555);
xor U13452 (N_13452,N_10395,N_10963);
nor U13453 (N_13453,N_10534,N_11454);
or U13454 (N_13454,N_11626,N_10843);
nand U13455 (N_13455,N_12361,N_10006);
xor U13456 (N_13456,N_11817,N_12190);
xnor U13457 (N_13457,N_10292,N_11754);
and U13458 (N_13458,N_10707,N_11031);
or U13459 (N_13459,N_11522,N_10608);
xnor U13460 (N_13460,N_10366,N_12008);
xor U13461 (N_13461,N_10767,N_12231);
or U13462 (N_13462,N_11041,N_10020);
and U13463 (N_13463,N_12329,N_12333);
and U13464 (N_13464,N_10151,N_10563);
nand U13465 (N_13465,N_12167,N_10071);
xnor U13466 (N_13466,N_10968,N_11717);
or U13467 (N_13467,N_10580,N_10206);
nand U13468 (N_13468,N_11837,N_12323);
nand U13469 (N_13469,N_10076,N_11811);
nor U13470 (N_13470,N_10245,N_11375);
or U13471 (N_13471,N_10589,N_10009);
nand U13472 (N_13472,N_11204,N_12161);
nand U13473 (N_13473,N_10306,N_10907);
nand U13474 (N_13474,N_10249,N_10244);
and U13475 (N_13475,N_10654,N_12150);
nor U13476 (N_13476,N_11272,N_10869);
xor U13477 (N_13477,N_12344,N_10060);
and U13478 (N_13478,N_10813,N_12243);
or U13479 (N_13479,N_11064,N_11700);
nand U13480 (N_13480,N_12192,N_12029);
xnor U13481 (N_13481,N_11271,N_10226);
or U13482 (N_13482,N_11976,N_11212);
xnor U13483 (N_13483,N_10496,N_10269);
nor U13484 (N_13484,N_11768,N_10112);
and U13485 (N_13485,N_11443,N_11496);
and U13486 (N_13486,N_12003,N_10849);
and U13487 (N_13487,N_11002,N_12275);
or U13488 (N_13488,N_12155,N_10487);
and U13489 (N_13489,N_10464,N_10858);
xnor U13490 (N_13490,N_10347,N_11970);
or U13491 (N_13491,N_10863,N_10879);
nand U13492 (N_13492,N_10692,N_12140);
nand U13493 (N_13493,N_12268,N_10124);
and U13494 (N_13494,N_10171,N_10373);
or U13495 (N_13495,N_11669,N_10090);
or U13496 (N_13496,N_11681,N_12022);
nand U13497 (N_13497,N_11338,N_10921);
or U13498 (N_13498,N_10372,N_10656);
nand U13499 (N_13499,N_11500,N_12431);
xor U13500 (N_13500,N_11429,N_11257);
and U13501 (N_13501,N_10628,N_10658);
and U13502 (N_13502,N_12132,N_10717);
or U13503 (N_13503,N_12414,N_11592);
or U13504 (N_13504,N_10780,N_11103);
nand U13505 (N_13505,N_10207,N_11472);
nor U13506 (N_13506,N_10365,N_10708);
nand U13507 (N_13507,N_10413,N_10549);
or U13508 (N_13508,N_11706,N_10769);
nor U13509 (N_13509,N_11577,N_10183);
and U13510 (N_13510,N_10854,N_11940);
xor U13511 (N_13511,N_10304,N_11775);
nor U13512 (N_13512,N_10710,N_10203);
or U13513 (N_13513,N_11574,N_10091);
and U13514 (N_13514,N_12486,N_11890);
nand U13515 (N_13515,N_11463,N_10387);
xnor U13516 (N_13516,N_12134,N_10385);
nand U13517 (N_13517,N_12072,N_10974);
nand U13518 (N_13518,N_11318,N_12163);
nor U13519 (N_13519,N_11171,N_10943);
and U13520 (N_13520,N_12413,N_10743);
nor U13521 (N_13521,N_11395,N_10137);
xnor U13522 (N_13522,N_12147,N_10042);
nor U13523 (N_13523,N_11703,N_10130);
or U13524 (N_13524,N_11067,N_11357);
or U13525 (N_13525,N_11033,N_10004);
xor U13526 (N_13526,N_11377,N_12014);
xnor U13527 (N_13527,N_11801,N_10303);
nand U13528 (N_13528,N_11800,N_12338);
or U13529 (N_13529,N_11240,N_11764);
or U13530 (N_13530,N_12269,N_10012);
nand U13531 (N_13531,N_10093,N_11025);
and U13532 (N_13532,N_10920,N_12096);
xor U13533 (N_13533,N_11558,N_11695);
or U13534 (N_13534,N_11416,N_11455);
xor U13535 (N_13535,N_11093,N_11862);
and U13536 (N_13536,N_10965,N_11606);
and U13537 (N_13537,N_11744,N_10147);
xor U13538 (N_13538,N_12496,N_12469);
or U13539 (N_13539,N_11549,N_11361);
nand U13540 (N_13540,N_11222,N_10270);
and U13541 (N_13541,N_11149,N_10694);
or U13542 (N_13542,N_10855,N_12239);
and U13543 (N_13543,N_11471,N_11520);
xor U13544 (N_13544,N_11951,N_11819);
nor U13545 (N_13545,N_10262,N_11823);
nor U13546 (N_13546,N_12326,N_10838);
and U13547 (N_13547,N_12104,N_10121);
and U13548 (N_13548,N_10911,N_11079);
and U13549 (N_13549,N_10786,N_11350);
or U13550 (N_13550,N_10517,N_11587);
nand U13551 (N_13551,N_12048,N_10293);
nand U13552 (N_13552,N_10264,N_10893);
nand U13553 (N_13553,N_11972,N_11607);
xor U13554 (N_13554,N_10856,N_12491);
or U13555 (N_13555,N_10507,N_10560);
xor U13556 (N_13556,N_10989,N_10029);
and U13557 (N_13557,N_11741,N_10557);
and U13558 (N_13558,N_11239,N_11120);
nand U13559 (N_13559,N_10693,N_11855);
nor U13560 (N_13560,N_12174,N_11286);
nor U13561 (N_13561,N_10682,N_11090);
and U13562 (N_13562,N_11742,N_10283);
and U13563 (N_13563,N_10553,N_11519);
or U13564 (N_13564,N_11007,N_12458);
and U13565 (N_13565,N_11581,N_11538);
nand U13566 (N_13566,N_10599,N_11126);
and U13567 (N_13567,N_10934,N_12193);
or U13568 (N_13568,N_11905,N_10276);
or U13569 (N_13569,N_11734,N_10638);
and U13570 (N_13570,N_11946,N_10700);
xor U13571 (N_13571,N_11961,N_11974);
nor U13572 (N_13572,N_10125,N_10458);
nor U13573 (N_13573,N_10705,N_12184);
xnor U13574 (N_13574,N_10652,N_12244);
or U13575 (N_13575,N_12427,N_10620);
nand U13576 (N_13576,N_12055,N_11233);
nor U13577 (N_13577,N_12237,N_10234);
nor U13578 (N_13578,N_10257,N_10254);
xnor U13579 (N_13579,N_11907,N_11708);
nor U13580 (N_13580,N_10456,N_12228);
and U13581 (N_13581,N_11791,N_12360);
or U13582 (N_13582,N_12357,N_11720);
nor U13583 (N_13583,N_12348,N_11402);
or U13584 (N_13584,N_11776,N_11697);
nand U13585 (N_13585,N_11759,N_11696);
or U13586 (N_13586,N_11829,N_11660);
or U13587 (N_13587,N_10575,N_11325);
or U13588 (N_13588,N_11915,N_10267);
nand U13589 (N_13589,N_10084,N_11279);
nand U13590 (N_13590,N_11055,N_11023);
or U13591 (N_13591,N_11139,N_10918);
and U13592 (N_13592,N_11405,N_10328);
nand U13593 (N_13593,N_11960,N_12289);
nor U13594 (N_13594,N_11005,N_12036);
or U13595 (N_13595,N_10972,N_11137);
xnor U13596 (N_13596,N_10683,N_10724);
xor U13597 (N_13597,N_12052,N_10069);
xnor U13598 (N_13598,N_11847,N_10509);
and U13599 (N_13599,N_11808,N_10073);
or U13600 (N_13600,N_10035,N_11353);
nor U13601 (N_13601,N_11076,N_11646);
nor U13602 (N_13602,N_11392,N_10383);
and U13603 (N_13603,N_12370,N_11451);
or U13604 (N_13604,N_10622,N_10066);
nor U13605 (N_13605,N_10744,N_11677);
xnor U13606 (N_13606,N_10392,N_11234);
and U13607 (N_13607,N_10430,N_10573);
nand U13608 (N_13608,N_11382,N_11447);
xor U13609 (N_13609,N_10542,N_11275);
or U13610 (N_13610,N_11135,N_11453);
nand U13611 (N_13611,N_12214,N_11578);
nor U13612 (N_13612,N_10050,N_10238);
and U13613 (N_13613,N_10904,N_10833);
or U13614 (N_13614,N_11637,N_11620);
xor U13615 (N_13615,N_11614,N_10815);
xnor U13616 (N_13616,N_12205,N_10895);
xnor U13617 (N_13617,N_11459,N_11231);
nor U13618 (N_13618,N_12363,N_12290);
xnor U13619 (N_13619,N_10197,N_11426);
nand U13620 (N_13620,N_10696,N_11893);
nor U13621 (N_13621,N_11709,N_11371);
or U13622 (N_13622,N_11370,N_11863);
or U13623 (N_13623,N_11541,N_11772);
nor U13624 (N_13624,N_11858,N_11482);
nor U13625 (N_13625,N_11509,N_11642);
or U13626 (N_13626,N_11673,N_11621);
nor U13627 (N_13627,N_10279,N_10448);
or U13628 (N_13628,N_11589,N_11354);
nand U13629 (N_13629,N_10364,N_11483);
nor U13630 (N_13630,N_10923,N_12005);
or U13631 (N_13631,N_11066,N_10827);
xor U13632 (N_13632,N_11209,N_10944);
xor U13633 (N_13633,N_10216,N_11654);
and U13634 (N_13634,N_10519,N_10554);
nor U13635 (N_13635,N_11270,N_10592);
nor U13636 (N_13636,N_11048,N_10949);
and U13637 (N_13637,N_11736,N_11804);
and U13638 (N_13638,N_10346,N_11553);
nor U13639 (N_13639,N_10175,N_12105);
and U13640 (N_13640,N_10663,N_10114);
or U13641 (N_13641,N_10333,N_10104);
nor U13642 (N_13642,N_12074,N_10924);
nor U13643 (N_13643,N_10651,N_10625);
or U13644 (N_13644,N_12467,N_10754);
xnor U13645 (N_13645,N_10411,N_10660);
and U13646 (N_13646,N_10082,N_11505);
nand U13647 (N_13647,N_12418,N_11579);
nor U13648 (N_13648,N_11879,N_11315);
nand U13649 (N_13649,N_11473,N_10630);
or U13650 (N_13650,N_11745,N_10357);
or U13651 (N_13651,N_11877,N_10994);
xor U13652 (N_13652,N_11105,N_11803);
nand U13653 (N_13653,N_12292,N_12211);
xor U13654 (N_13654,N_10647,N_10247);
xnor U13655 (N_13655,N_11024,N_11973);
nor U13656 (N_13656,N_11143,N_11615);
and U13657 (N_13657,N_10044,N_11445);
xor U13658 (N_13658,N_11882,N_10962);
nand U13659 (N_13659,N_11629,N_11158);
nor U13660 (N_13660,N_11456,N_10712);
nand U13661 (N_13661,N_10716,N_11514);
nand U13662 (N_13662,N_11340,N_11194);
nor U13663 (N_13663,N_11599,N_12259);
and U13664 (N_13664,N_12153,N_10670);
xor U13665 (N_13665,N_12136,N_10484);
xnor U13666 (N_13666,N_11247,N_10409);
xnor U13667 (N_13667,N_10993,N_12460);
nand U13668 (N_13668,N_12065,N_11839);
or U13669 (N_13669,N_11825,N_10210);
or U13670 (N_13670,N_11567,N_10634);
or U13671 (N_13671,N_10861,N_11085);
xor U13672 (N_13672,N_12327,N_10529);
nor U13673 (N_13673,N_11632,N_10837);
nor U13674 (N_13674,N_10186,N_12233);
xor U13675 (N_13675,N_11386,N_12063);
or U13676 (N_13676,N_11020,N_11892);
nand U13677 (N_13677,N_11096,N_11049);
nor U13678 (N_13678,N_10314,N_11051);
or U13679 (N_13679,N_12482,N_10189);
nand U13680 (N_13680,N_11124,N_12287);
nand U13681 (N_13681,N_12070,N_11752);
xnor U13682 (N_13682,N_10441,N_11604);
nand U13683 (N_13683,N_12324,N_10990);
xor U13684 (N_13684,N_12060,N_11662);
and U13685 (N_13685,N_12221,N_11569);
nor U13686 (N_13686,N_12139,N_11331);
and U13687 (N_13687,N_11401,N_12355);
and U13688 (N_13688,N_11643,N_11290);
xor U13689 (N_13689,N_10844,N_11949);
and U13690 (N_13690,N_11349,N_10078);
xnor U13691 (N_13691,N_12453,N_10498);
nand U13692 (N_13692,N_12251,N_11834);
or U13693 (N_13693,N_10191,N_10526);
and U13694 (N_13694,N_10405,N_11293);
nor U13695 (N_13695,N_10024,N_11150);
xor U13696 (N_13696,N_12316,N_12378);
or U13697 (N_13697,N_11743,N_11788);
xor U13698 (N_13698,N_12419,N_11123);
or U13699 (N_13699,N_12436,N_10865);
or U13700 (N_13700,N_12157,N_10209);
xor U13701 (N_13701,N_10900,N_12217);
and U13702 (N_13702,N_11358,N_11900);
or U13703 (N_13703,N_11665,N_10617);
nand U13704 (N_13704,N_10750,N_11283);
and U13705 (N_13705,N_11191,N_10442);
and U13706 (N_13706,N_10466,N_11908);
or U13707 (N_13707,N_12384,N_10715);
xor U13708 (N_13708,N_12426,N_12182);
xnor U13709 (N_13709,N_11190,N_10937);
nor U13710 (N_13710,N_11130,N_10841);
xnor U13711 (N_13711,N_12321,N_10999);
xnor U13712 (N_13712,N_12133,N_10388);
nand U13713 (N_13713,N_11475,N_10057);
nand U13714 (N_13714,N_10641,N_11294);
nand U13715 (N_13715,N_10794,N_11608);
xnor U13716 (N_13716,N_12007,N_10031);
and U13717 (N_13717,N_12002,N_10596);
xnor U13718 (N_13718,N_10791,N_10483);
or U13719 (N_13719,N_10068,N_11732);
and U13720 (N_13720,N_10816,N_11238);
nor U13721 (N_13721,N_12441,N_11868);
nand U13722 (N_13722,N_12339,N_11870);
nand U13723 (N_13723,N_12158,N_11508);
nor U13724 (N_13724,N_10859,N_11573);
or U13725 (N_13725,N_11097,N_11427);
nand U13726 (N_13726,N_10220,N_11226);
nand U13727 (N_13727,N_11359,N_10370);
and U13728 (N_13728,N_11760,N_10545);
or U13729 (N_13729,N_11467,N_12267);
nor U13730 (N_13730,N_10997,N_10320);
or U13731 (N_13731,N_10610,N_10925);
or U13732 (N_13732,N_11566,N_11691);
or U13733 (N_13733,N_10761,N_12225);
or U13734 (N_13734,N_10729,N_11936);
nand U13735 (N_13735,N_10503,N_10027);
nand U13736 (N_13736,N_12325,N_11636);
xnor U13737 (N_13737,N_11682,N_11166);
nand U13738 (N_13738,N_11301,N_12118);
or U13739 (N_13739,N_12203,N_10489);
nor U13740 (N_13740,N_10323,N_11526);
xnor U13741 (N_13741,N_12009,N_12010);
nor U13742 (N_13742,N_12073,N_10979);
or U13743 (N_13743,N_10749,N_12035);
nor U13744 (N_13744,N_10061,N_10116);
xnor U13745 (N_13745,N_11295,N_10759);
and U13746 (N_13746,N_10133,N_10566);
and U13747 (N_13747,N_10248,N_10714);
or U13748 (N_13748,N_11449,N_12119);
or U13749 (N_13749,N_11527,N_10577);
or U13750 (N_13750,N_11094,N_11846);
xor U13751 (N_13751,N_10441,N_11194);
xnor U13752 (N_13752,N_11416,N_11008);
and U13753 (N_13753,N_10360,N_11538);
nand U13754 (N_13754,N_11377,N_11703);
or U13755 (N_13755,N_12060,N_11385);
or U13756 (N_13756,N_10165,N_10569);
and U13757 (N_13757,N_11057,N_10102);
xnor U13758 (N_13758,N_10345,N_11665);
nand U13759 (N_13759,N_12219,N_11503);
or U13760 (N_13760,N_10654,N_10991);
or U13761 (N_13761,N_12306,N_10375);
nand U13762 (N_13762,N_10291,N_10389);
nor U13763 (N_13763,N_12118,N_12353);
xor U13764 (N_13764,N_12125,N_10617);
and U13765 (N_13765,N_10242,N_11513);
nand U13766 (N_13766,N_10219,N_10448);
nor U13767 (N_13767,N_11556,N_10607);
xor U13768 (N_13768,N_10878,N_10305);
nor U13769 (N_13769,N_10027,N_11211);
nand U13770 (N_13770,N_10248,N_11792);
or U13771 (N_13771,N_10384,N_10174);
nor U13772 (N_13772,N_11132,N_10021);
nand U13773 (N_13773,N_10423,N_11454);
xnor U13774 (N_13774,N_11257,N_10499);
nand U13775 (N_13775,N_10805,N_10523);
and U13776 (N_13776,N_10250,N_10820);
xor U13777 (N_13777,N_11187,N_12468);
nand U13778 (N_13778,N_12360,N_10997);
or U13779 (N_13779,N_12286,N_11943);
or U13780 (N_13780,N_11498,N_10649);
nand U13781 (N_13781,N_10292,N_10172);
nand U13782 (N_13782,N_11574,N_12352);
xnor U13783 (N_13783,N_11324,N_12129);
nor U13784 (N_13784,N_10487,N_10628);
xor U13785 (N_13785,N_10035,N_11617);
xnor U13786 (N_13786,N_11775,N_12476);
nand U13787 (N_13787,N_12380,N_12156);
nand U13788 (N_13788,N_10587,N_10294);
nor U13789 (N_13789,N_11617,N_11373);
xnor U13790 (N_13790,N_11374,N_10607);
nor U13791 (N_13791,N_11027,N_10011);
nor U13792 (N_13792,N_10969,N_10064);
and U13793 (N_13793,N_11793,N_10059);
and U13794 (N_13794,N_11542,N_10989);
nor U13795 (N_13795,N_11934,N_10529);
and U13796 (N_13796,N_11382,N_10953);
or U13797 (N_13797,N_10849,N_10250);
or U13798 (N_13798,N_10588,N_11432);
nand U13799 (N_13799,N_10345,N_11447);
nor U13800 (N_13800,N_11379,N_11079);
and U13801 (N_13801,N_12150,N_11814);
xor U13802 (N_13802,N_10929,N_10561);
xnor U13803 (N_13803,N_12356,N_10776);
and U13804 (N_13804,N_11306,N_10248);
nand U13805 (N_13805,N_11475,N_10079);
xor U13806 (N_13806,N_12321,N_10248);
and U13807 (N_13807,N_10497,N_10760);
nand U13808 (N_13808,N_10557,N_10427);
nand U13809 (N_13809,N_11429,N_10321);
nor U13810 (N_13810,N_12218,N_11957);
nand U13811 (N_13811,N_12299,N_10828);
nand U13812 (N_13812,N_12476,N_10423);
or U13813 (N_13813,N_10036,N_10834);
or U13814 (N_13814,N_10377,N_11777);
nor U13815 (N_13815,N_11646,N_11467);
and U13816 (N_13816,N_10824,N_11639);
and U13817 (N_13817,N_11624,N_11216);
nor U13818 (N_13818,N_12319,N_12296);
or U13819 (N_13819,N_11605,N_10758);
nand U13820 (N_13820,N_12452,N_10805);
nand U13821 (N_13821,N_11405,N_12392);
and U13822 (N_13822,N_12123,N_10183);
nor U13823 (N_13823,N_10408,N_11218);
xor U13824 (N_13824,N_10888,N_12236);
nand U13825 (N_13825,N_12419,N_11918);
nand U13826 (N_13826,N_10111,N_10604);
or U13827 (N_13827,N_11613,N_11909);
xor U13828 (N_13828,N_10936,N_10799);
nor U13829 (N_13829,N_10426,N_12295);
or U13830 (N_13830,N_10340,N_11135);
xor U13831 (N_13831,N_10169,N_12343);
xor U13832 (N_13832,N_11511,N_12258);
or U13833 (N_13833,N_10975,N_12066);
or U13834 (N_13834,N_11296,N_11887);
or U13835 (N_13835,N_11465,N_11880);
nor U13836 (N_13836,N_12328,N_11205);
nand U13837 (N_13837,N_10125,N_12244);
and U13838 (N_13838,N_12108,N_11179);
nand U13839 (N_13839,N_10788,N_10949);
xor U13840 (N_13840,N_12009,N_10448);
and U13841 (N_13841,N_12145,N_10061);
nand U13842 (N_13842,N_10145,N_10168);
xor U13843 (N_13843,N_11221,N_10947);
or U13844 (N_13844,N_11383,N_12406);
nor U13845 (N_13845,N_10385,N_11673);
nand U13846 (N_13846,N_12262,N_12092);
or U13847 (N_13847,N_10101,N_11913);
nor U13848 (N_13848,N_11264,N_10296);
nor U13849 (N_13849,N_11922,N_10215);
xnor U13850 (N_13850,N_12144,N_10075);
or U13851 (N_13851,N_11017,N_11204);
nor U13852 (N_13852,N_10047,N_11147);
nor U13853 (N_13853,N_12276,N_12478);
xnor U13854 (N_13854,N_12035,N_12240);
nand U13855 (N_13855,N_11981,N_11105);
or U13856 (N_13856,N_11950,N_10973);
and U13857 (N_13857,N_11955,N_11910);
nand U13858 (N_13858,N_10577,N_11560);
xor U13859 (N_13859,N_10013,N_10476);
or U13860 (N_13860,N_12424,N_11068);
and U13861 (N_13861,N_10735,N_12458);
or U13862 (N_13862,N_11157,N_12265);
or U13863 (N_13863,N_10443,N_10460);
xor U13864 (N_13864,N_10931,N_10659);
and U13865 (N_13865,N_11089,N_12135);
and U13866 (N_13866,N_12348,N_11970);
xnor U13867 (N_13867,N_11348,N_11158);
and U13868 (N_13868,N_10832,N_11164);
nand U13869 (N_13869,N_10189,N_11879);
or U13870 (N_13870,N_11772,N_11623);
or U13871 (N_13871,N_10059,N_11266);
nor U13872 (N_13872,N_10857,N_11176);
nand U13873 (N_13873,N_11114,N_11388);
and U13874 (N_13874,N_11750,N_11212);
and U13875 (N_13875,N_11445,N_10547);
and U13876 (N_13876,N_11009,N_10899);
or U13877 (N_13877,N_10100,N_10192);
xor U13878 (N_13878,N_11310,N_11179);
and U13879 (N_13879,N_11221,N_10022);
and U13880 (N_13880,N_10828,N_10385);
nand U13881 (N_13881,N_10828,N_12379);
nand U13882 (N_13882,N_10979,N_10209);
nor U13883 (N_13883,N_10270,N_11700);
nor U13884 (N_13884,N_12337,N_11067);
nor U13885 (N_13885,N_10423,N_11067);
and U13886 (N_13886,N_11212,N_10764);
or U13887 (N_13887,N_11875,N_11528);
xor U13888 (N_13888,N_11192,N_10803);
and U13889 (N_13889,N_12306,N_11656);
nor U13890 (N_13890,N_12125,N_12255);
or U13891 (N_13891,N_12453,N_10183);
nand U13892 (N_13892,N_12404,N_11213);
xor U13893 (N_13893,N_11088,N_11670);
nand U13894 (N_13894,N_12380,N_10275);
nand U13895 (N_13895,N_10882,N_11154);
and U13896 (N_13896,N_11258,N_12202);
or U13897 (N_13897,N_12013,N_11875);
and U13898 (N_13898,N_11289,N_12437);
and U13899 (N_13899,N_11592,N_12033);
and U13900 (N_13900,N_11960,N_12126);
or U13901 (N_13901,N_10503,N_11052);
or U13902 (N_13902,N_11111,N_11570);
and U13903 (N_13903,N_10158,N_10372);
or U13904 (N_13904,N_12470,N_12342);
xor U13905 (N_13905,N_11102,N_10226);
xor U13906 (N_13906,N_12389,N_11251);
xor U13907 (N_13907,N_11639,N_10987);
and U13908 (N_13908,N_10474,N_11529);
or U13909 (N_13909,N_10768,N_11396);
nand U13910 (N_13910,N_12349,N_12075);
or U13911 (N_13911,N_11335,N_12281);
xnor U13912 (N_13912,N_10144,N_11192);
nand U13913 (N_13913,N_10719,N_10085);
and U13914 (N_13914,N_10831,N_12166);
nor U13915 (N_13915,N_11976,N_11567);
or U13916 (N_13916,N_10699,N_10603);
xnor U13917 (N_13917,N_10648,N_12412);
or U13918 (N_13918,N_10885,N_12261);
and U13919 (N_13919,N_12442,N_11399);
nand U13920 (N_13920,N_11662,N_12316);
xnor U13921 (N_13921,N_12275,N_11141);
and U13922 (N_13922,N_12046,N_11066);
and U13923 (N_13923,N_11407,N_10676);
or U13924 (N_13924,N_11515,N_12239);
nor U13925 (N_13925,N_12055,N_12327);
and U13926 (N_13926,N_12338,N_11416);
nor U13927 (N_13927,N_11596,N_10580);
nand U13928 (N_13928,N_12369,N_11781);
xnor U13929 (N_13929,N_12206,N_11859);
nor U13930 (N_13930,N_12343,N_10277);
and U13931 (N_13931,N_11214,N_12451);
nor U13932 (N_13932,N_12317,N_12006);
xor U13933 (N_13933,N_12473,N_10213);
nand U13934 (N_13934,N_11384,N_10836);
nand U13935 (N_13935,N_10018,N_12368);
nand U13936 (N_13936,N_10623,N_10970);
nor U13937 (N_13937,N_10268,N_11477);
nand U13938 (N_13938,N_10253,N_11869);
or U13939 (N_13939,N_10860,N_10409);
or U13940 (N_13940,N_11005,N_11230);
nor U13941 (N_13941,N_12438,N_11214);
nor U13942 (N_13942,N_11582,N_10267);
nor U13943 (N_13943,N_12368,N_10687);
or U13944 (N_13944,N_10630,N_11104);
nand U13945 (N_13945,N_11375,N_12286);
xnor U13946 (N_13946,N_10581,N_11259);
nand U13947 (N_13947,N_11913,N_11375);
or U13948 (N_13948,N_10985,N_10788);
nand U13949 (N_13949,N_10366,N_11796);
xor U13950 (N_13950,N_12379,N_12298);
and U13951 (N_13951,N_10333,N_11246);
nor U13952 (N_13952,N_10616,N_11994);
nand U13953 (N_13953,N_10085,N_12132);
xor U13954 (N_13954,N_10975,N_10222);
xor U13955 (N_13955,N_12043,N_11509);
or U13956 (N_13956,N_10236,N_11874);
and U13957 (N_13957,N_11624,N_10473);
or U13958 (N_13958,N_11283,N_10481);
or U13959 (N_13959,N_11588,N_12357);
and U13960 (N_13960,N_11780,N_11583);
nand U13961 (N_13961,N_10151,N_11446);
or U13962 (N_13962,N_11303,N_10097);
and U13963 (N_13963,N_10881,N_12145);
nand U13964 (N_13964,N_11206,N_11637);
and U13965 (N_13965,N_11161,N_10094);
and U13966 (N_13966,N_11085,N_12101);
and U13967 (N_13967,N_11450,N_11954);
or U13968 (N_13968,N_10692,N_11730);
nand U13969 (N_13969,N_12135,N_10559);
nor U13970 (N_13970,N_11165,N_11877);
and U13971 (N_13971,N_11360,N_12117);
or U13972 (N_13972,N_10458,N_10016);
or U13973 (N_13973,N_11217,N_10976);
and U13974 (N_13974,N_10818,N_12379);
xnor U13975 (N_13975,N_11968,N_11886);
or U13976 (N_13976,N_12158,N_11795);
nor U13977 (N_13977,N_11116,N_11104);
nor U13978 (N_13978,N_11195,N_11831);
nor U13979 (N_13979,N_11954,N_11498);
nand U13980 (N_13980,N_11915,N_12120);
nand U13981 (N_13981,N_10720,N_12166);
nor U13982 (N_13982,N_12382,N_11470);
nand U13983 (N_13983,N_10317,N_12125);
and U13984 (N_13984,N_10694,N_10917);
and U13985 (N_13985,N_10212,N_10886);
and U13986 (N_13986,N_11291,N_11476);
or U13987 (N_13987,N_12184,N_11818);
nand U13988 (N_13988,N_10052,N_11664);
xnor U13989 (N_13989,N_11127,N_10244);
and U13990 (N_13990,N_11360,N_10119);
or U13991 (N_13991,N_10490,N_12251);
nand U13992 (N_13992,N_11240,N_11616);
nor U13993 (N_13993,N_11224,N_11070);
xor U13994 (N_13994,N_11695,N_12179);
nand U13995 (N_13995,N_10532,N_12220);
and U13996 (N_13996,N_12449,N_10672);
nand U13997 (N_13997,N_11015,N_10878);
xnor U13998 (N_13998,N_12356,N_11052);
nand U13999 (N_13999,N_10462,N_11285);
xor U14000 (N_14000,N_10489,N_11168);
or U14001 (N_14001,N_10705,N_11695);
nor U14002 (N_14002,N_12135,N_10988);
xnor U14003 (N_14003,N_11232,N_11377);
nand U14004 (N_14004,N_11824,N_11525);
xor U14005 (N_14005,N_11284,N_10721);
nor U14006 (N_14006,N_11139,N_11979);
nor U14007 (N_14007,N_10969,N_10194);
xnor U14008 (N_14008,N_10168,N_10077);
nor U14009 (N_14009,N_11259,N_11941);
xor U14010 (N_14010,N_12074,N_10168);
nand U14011 (N_14011,N_10710,N_10258);
and U14012 (N_14012,N_10152,N_12443);
xor U14013 (N_14013,N_11909,N_10675);
xnor U14014 (N_14014,N_11685,N_11035);
nand U14015 (N_14015,N_10922,N_12188);
nand U14016 (N_14016,N_11506,N_12281);
nor U14017 (N_14017,N_11648,N_12432);
or U14018 (N_14018,N_11426,N_11817);
nand U14019 (N_14019,N_10416,N_11917);
or U14020 (N_14020,N_10852,N_12158);
nand U14021 (N_14021,N_11875,N_12019);
and U14022 (N_14022,N_10276,N_12302);
nor U14023 (N_14023,N_10368,N_10894);
nor U14024 (N_14024,N_10474,N_11721);
nand U14025 (N_14025,N_11618,N_10086);
nand U14026 (N_14026,N_10006,N_11247);
or U14027 (N_14027,N_12154,N_10568);
and U14028 (N_14028,N_11896,N_11832);
and U14029 (N_14029,N_10850,N_11101);
xor U14030 (N_14030,N_10587,N_10708);
nor U14031 (N_14031,N_11316,N_10455);
and U14032 (N_14032,N_11883,N_12196);
or U14033 (N_14033,N_10379,N_10683);
and U14034 (N_14034,N_12392,N_11074);
or U14035 (N_14035,N_11367,N_10175);
or U14036 (N_14036,N_12428,N_10659);
nand U14037 (N_14037,N_12018,N_11719);
xor U14038 (N_14038,N_11591,N_11424);
nand U14039 (N_14039,N_12464,N_12185);
or U14040 (N_14040,N_11094,N_10591);
xor U14041 (N_14041,N_10406,N_10025);
or U14042 (N_14042,N_11724,N_10827);
and U14043 (N_14043,N_10533,N_11440);
and U14044 (N_14044,N_12223,N_10522);
nand U14045 (N_14045,N_12305,N_10056);
nand U14046 (N_14046,N_10867,N_11135);
or U14047 (N_14047,N_12088,N_11395);
or U14048 (N_14048,N_11472,N_10471);
nand U14049 (N_14049,N_12197,N_10386);
nor U14050 (N_14050,N_11443,N_10138);
and U14051 (N_14051,N_10569,N_12030);
and U14052 (N_14052,N_10960,N_11068);
nand U14053 (N_14053,N_12301,N_10842);
or U14054 (N_14054,N_11682,N_10883);
nand U14055 (N_14055,N_11984,N_11460);
xnor U14056 (N_14056,N_11213,N_10046);
and U14057 (N_14057,N_10797,N_10678);
xor U14058 (N_14058,N_11072,N_11778);
nor U14059 (N_14059,N_11208,N_10264);
or U14060 (N_14060,N_10784,N_10419);
nand U14061 (N_14061,N_10603,N_11076);
nor U14062 (N_14062,N_11950,N_10117);
or U14063 (N_14063,N_11932,N_10760);
or U14064 (N_14064,N_12001,N_10612);
xnor U14065 (N_14065,N_10049,N_11962);
and U14066 (N_14066,N_11504,N_12047);
nand U14067 (N_14067,N_10896,N_10370);
and U14068 (N_14068,N_10543,N_12051);
xor U14069 (N_14069,N_11748,N_10398);
or U14070 (N_14070,N_12282,N_11581);
or U14071 (N_14071,N_11144,N_11183);
and U14072 (N_14072,N_12473,N_10240);
nor U14073 (N_14073,N_10815,N_12298);
nand U14074 (N_14074,N_10527,N_11379);
or U14075 (N_14075,N_11143,N_10316);
xnor U14076 (N_14076,N_12024,N_10483);
nand U14077 (N_14077,N_10187,N_10020);
nand U14078 (N_14078,N_10144,N_12254);
nor U14079 (N_14079,N_11835,N_10082);
nor U14080 (N_14080,N_11133,N_11722);
xnor U14081 (N_14081,N_11251,N_10943);
xnor U14082 (N_14082,N_12205,N_11241);
or U14083 (N_14083,N_10975,N_10177);
nand U14084 (N_14084,N_12109,N_11476);
and U14085 (N_14085,N_12215,N_10726);
or U14086 (N_14086,N_10369,N_11924);
and U14087 (N_14087,N_11392,N_11398);
xnor U14088 (N_14088,N_11074,N_11951);
nand U14089 (N_14089,N_11396,N_10576);
nand U14090 (N_14090,N_12217,N_11832);
and U14091 (N_14091,N_10999,N_10652);
and U14092 (N_14092,N_11475,N_12163);
xnor U14093 (N_14093,N_12038,N_10552);
nand U14094 (N_14094,N_12152,N_11059);
xnor U14095 (N_14095,N_11160,N_12184);
and U14096 (N_14096,N_11925,N_12002);
xor U14097 (N_14097,N_11462,N_10863);
nand U14098 (N_14098,N_11120,N_12182);
or U14099 (N_14099,N_11997,N_11245);
or U14100 (N_14100,N_12377,N_12239);
nand U14101 (N_14101,N_11742,N_11028);
or U14102 (N_14102,N_11346,N_11394);
nor U14103 (N_14103,N_11598,N_10133);
xnor U14104 (N_14104,N_10087,N_11303);
or U14105 (N_14105,N_11619,N_12201);
nand U14106 (N_14106,N_10358,N_11351);
or U14107 (N_14107,N_11761,N_12321);
nand U14108 (N_14108,N_11745,N_12340);
or U14109 (N_14109,N_11426,N_12060);
and U14110 (N_14110,N_11832,N_11481);
and U14111 (N_14111,N_12035,N_11663);
or U14112 (N_14112,N_12090,N_10354);
nor U14113 (N_14113,N_11652,N_11198);
and U14114 (N_14114,N_12023,N_12134);
nor U14115 (N_14115,N_10229,N_12331);
and U14116 (N_14116,N_10144,N_10852);
nand U14117 (N_14117,N_10387,N_10150);
nor U14118 (N_14118,N_11874,N_10895);
or U14119 (N_14119,N_10504,N_11223);
or U14120 (N_14120,N_11288,N_11078);
or U14121 (N_14121,N_10405,N_12182);
and U14122 (N_14122,N_10367,N_11134);
xnor U14123 (N_14123,N_11152,N_11394);
or U14124 (N_14124,N_11392,N_11205);
xor U14125 (N_14125,N_12213,N_10105);
nand U14126 (N_14126,N_11461,N_12234);
nor U14127 (N_14127,N_11520,N_10019);
xnor U14128 (N_14128,N_11285,N_10909);
or U14129 (N_14129,N_11485,N_10248);
or U14130 (N_14130,N_10515,N_12080);
and U14131 (N_14131,N_10033,N_10476);
nand U14132 (N_14132,N_10982,N_11733);
or U14133 (N_14133,N_10886,N_10255);
nor U14134 (N_14134,N_12441,N_10850);
nand U14135 (N_14135,N_10682,N_11573);
nand U14136 (N_14136,N_12003,N_11688);
nor U14137 (N_14137,N_10757,N_11453);
xor U14138 (N_14138,N_10053,N_12068);
or U14139 (N_14139,N_11614,N_10466);
and U14140 (N_14140,N_12366,N_12333);
or U14141 (N_14141,N_10813,N_11036);
and U14142 (N_14142,N_10200,N_10193);
nor U14143 (N_14143,N_11909,N_11421);
and U14144 (N_14144,N_10050,N_10672);
or U14145 (N_14145,N_11675,N_10724);
or U14146 (N_14146,N_11152,N_12156);
and U14147 (N_14147,N_12176,N_10959);
and U14148 (N_14148,N_11726,N_12374);
or U14149 (N_14149,N_10491,N_10544);
and U14150 (N_14150,N_11148,N_10211);
and U14151 (N_14151,N_10322,N_10262);
or U14152 (N_14152,N_11780,N_11276);
and U14153 (N_14153,N_10112,N_10838);
nor U14154 (N_14154,N_12279,N_12042);
nand U14155 (N_14155,N_12340,N_11173);
nor U14156 (N_14156,N_10275,N_10745);
nand U14157 (N_14157,N_11855,N_12253);
and U14158 (N_14158,N_12059,N_11204);
nor U14159 (N_14159,N_12063,N_11348);
nor U14160 (N_14160,N_11614,N_10251);
and U14161 (N_14161,N_11261,N_11895);
or U14162 (N_14162,N_11329,N_11734);
nand U14163 (N_14163,N_11890,N_10952);
xnor U14164 (N_14164,N_11077,N_10318);
nor U14165 (N_14165,N_12404,N_11703);
nand U14166 (N_14166,N_10883,N_12135);
or U14167 (N_14167,N_10354,N_11231);
nor U14168 (N_14168,N_12045,N_11522);
or U14169 (N_14169,N_11394,N_11427);
and U14170 (N_14170,N_11847,N_11377);
and U14171 (N_14171,N_11877,N_11810);
nand U14172 (N_14172,N_10646,N_11780);
or U14173 (N_14173,N_12077,N_11456);
nor U14174 (N_14174,N_12006,N_11623);
or U14175 (N_14175,N_11649,N_11414);
nor U14176 (N_14176,N_11862,N_12227);
nor U14177 (N_14177,N_10393,N_10648);
or U14178 (N_14178,N_10192,N_10221);
or U14179 (N_14179,N_10742,N_11719);
and U14180 (N_14180,N_12123,N_10720);
nor U14181 (N_14181,N_11330,N_11666);
nand U14182 (N_14182,N_10942,N_10663);
nor U14183 (N_14183,N_10785,N_11181);
nor U14184 (N_14184,N_10329,N_10761);
nor U14185 (N_14185,N_11587,N_11134);
xnor U14186 (N_14186,N_10475,N_10266);
and U14187 (N_14187,N_11435,N_11792);
xnor U14188 (N_14188,N_10673,N_10778);
or U14189 (N_14189,N_11981,N_10749);
and U14190 (N_14190,N_10439,N_11316);
nand U14191 (N_14191,N_10325,N_11457);
nor U14192 (N_14192,N_10324,N_11591);
nor U14193 (N_14193,N_10686,N_12089);
nand U14194 (N_14194,N_11125,N_11441);
nor U14195 (N_14195,N_12439,N_11062);
and U14196 (N_14196,N_12477,N_10069);
nand U14197 (N_14197,N_11787,N_11387);
or U14198 (N_14198,N_10029,N_11813);
and U14199 (N_14199,N_10400,N_11838);
xnor U14200 (N_14200,N_10073,N_11008);
xor U14201 (N_14201,N_11485,N_11336);
xor U14202 (N_14202,N_11216,N_11825);
and U14203 (N_14203,N_12348,N_11800);
nand U14204 (N_14204,N_11435,N_11903);
nand U14205 (N_14205,N_10311,N_10200);
or U14206 (N_14206,N_10335,N_11636);
and U14207 (N_14207,N_11410,N_10294);
nor U14208 (N_14208,N_11010,N_11503);
nand U14209 (N_14209,N_11540,N_10444);
and U14210 (N_14210,N_10129,N_11474);
nand U14211 (N_14211,N_10926,N_12313);
xnor U14212 (N_14212,N_12108,N_11546);
xor U14213 (N_14213,N_11453,N_11824);
nor U14214 (N_14214,N_11100,N_11666);
xor U14215 (N_14215,N_11250,N_12305);
nor U14216 (N_14216,N_11150,N_10764);
xnor U14217 (N_14217,N_12461,N_11030);
nor U14218 (N_14218,N_11416,N_12080);
or U14219 (N_14219,N_12258,N_11930);
xor U14220 (N_14220,N_11298,N_12031);
or U14221 (N_14221,N_12130,N_11676);
or U14222 (N_14222,N_10180,N_11281);
nand U14223 (N_14223,N_11624,N_10091);
nor U14224 (N_14224,N_11789,N_10312);
or U14225 (N_14225,N_10485,N_10566);
nor U14226 (N_14226,N_12350,N_10372);
xnor U14227 (N_14227,N_10165,N_11031);
or U14228 (N_14228,N_11369,N_12059);
or U14229 (N_14229,N_10709,N_10344);
or U14230 (N_14230,N_10387,N_12415);
nand U14231 (N_14231,N_10341,N_12286);
or U14232 (N_14232,N_10560,N_10382);
nor U14233 (N_14233,N_11928,N_11986);
xor U14234 (N_14234,N_11552,N_11340);
xor U14235 (N_14235,N_10086,N_10323);
or U14236 (N_14236,N_10800,N_11786);
nor U14237 (N_14237,N_10943,N_11291);
or U14238 (N_14238,N_11806,N_11630);
xor U14239 (N_14239,N_11411,N_11679);
or U14240 (N_14240,N_10656,N_12471);
xor U14241 (N_14241,N_12071,N_10320);
nand U14242 (N_14242,N_10876,N_12481);
nor U14243 (N_14243,N_11501,N_12196);
or U14244 (N_14244,N_12221,N_10353);
nor U14245 (N_14245,N_11378,N_10845);
xor U14246 (N_14246,N_10422,N_11883);
or U14247 (N_14247,N_11341,N_11204);
nand U14248 (N_14248,N_11725,N_11462);
and U14249 (N_14249,N_11921,N_10983);
and U14250 (N_14250,N_12045,N_10171);
xor U14251 (N_14251,N_11200,N_11288);
nor U14252 (N_14252,N_11525,N_12397);
nand U14253 (N_14253,N_11911,N_11029);
xnor U14254 (N_14254,N_12493,N_11521);
nand U14255 (N_14255,N_11540,N_10840);
or U14256 (N_14256,N_12099,N_12296);
nand U14257 (N_14257,N_12036,N_10110);
and U14258 (N_14258,N_11939,N_10469);
and U14259 (N_14259,N_11313,N_11208);
nor U14260 (N_14260,N_10683,N_11387);
xnor U14261 (N_14261,N_12448,N_12482);
xnor U14262 (N_14262,N_10274,N_12475);
nand U14263 (N_14263,N_12386,N_12089);
xnor U14264 (N_14264,N_11658,N_10406);
nor U14265 (N_14265,N_11519,N_11217);
and U14266 (N_14266,N_10512,N_11739);
nand U14267 (N_14267,N_11163,N_12079);
and U14268 (N_14268,N_10648,N_11512);
xor U14269 (N_14269,N_10362,N_10000);
xnor U14270 (N_14270,N_10463,N_11887);
nand U14271 (N_14271,N_11763,N_10403);
nor U14272 (N_14272,N_11996,N_12343);
and U14273 (N_14273,N_11126,N_10537);
nand U14274 (N_14274,N_11212,N_11251);
and U14275 (N_14275,N_11493,N_10946);
nand U14276 (N_14276,N_12002,N_11975);
nand U14277 (N_14277,N_12434,N_12059);
xor U14278 (N_14278,N_10589,N_11334);
and U14279 (N_14279,N_11101,N_12328);
or U14280 (N_14280,N_10259,N_11626);
nor U14281 (N_14281,N_11458,N_10645);
or U14282 (N_14282,N_11208,N_10905);
and U14283 (N_14283,N_12053,N_11718);
or U14284 (N_14284,N_10827,N_12113);
xnor U14285 (N_14285,N_12060,N_10240);
nand U14286 (N_14286,N_11340,N_12155);
nor U14287 (N_14287,N_10899,N_10531);
or U14288 (N_14288,N_12185,N_10493);
nand U14289 (N_14289,N_11708,N_11614);
and U14290 (N_14290,N_11082,N_11481);
nand U14291 (N_14291,N_10097,N_10241);
and U14292 (N_14292,N_11939,N_10015);
xnor U14293 (N_14293,N_11513,N_11935);
nor U14294 (N_14294,N_10507,N_10546);
nand U14295 (N_14295,N_11403,N_12109);
xor U14296 (N_14296,N_12215,N_10107);
nor U14297 (N_14297,N_10947,N_12400);
xor U14298 (N_14298,N_11033,N_12134);
nor U14299 (N_14299,N_11910,N_10635);
xor U14300 (N_14300,N_10807,N_12042);
xor U14301 (N_14301,N_12285,N_10151);
nor U14302 (N_14302,N_12014,N_10522);
nand U14303 (N_14303,N_12161,N_12041);
nand U14304 (N_14304,N_10475,N_11841);
nand U14305 (N_14305,N_11394,N_11179);
nor U14306 (N_14306,N_11799,N_10862);
nor U14307 (N_14307,N_10295,N_10812);
xor U14308 (N_14308,N_12258,N_11213);
xor U14309 (N_14309,N_10804,N_11600);
and U14310 (N_14310,N_11352,N_10968);
nand U14311 (N_14311,N_10689,N_11333);
nand U14312 (N_14312,N_11993,N_11846);
nand U14313 (N_14313,N_12001,N_10472);
nor U14314 (N_14314,N_10322,N_11145);
nand U14315 (N_14315,N_10111,N_10980);
nand U14316 (N_14316,N_12390,N_11139);
nand U14317 (N_14317,N_10153,N_12125);
or U14318 (N_14318,N_11651,N_12424);
xnor U14319 (N_14319,N_10669,N_10343);
or U14320 (N_14320,N_10518,N_12024);
nand U14321 (N_14321,N_11608,N_12356);
xor U14322 (N_14322,N_11881,N_10819);
or U14323 (N_14323,N_11240,N_11428);
and U14324 (N_14324,N_10193,N_12197);
xnor U14325 (N_14325,N_10038,N_12195);
xor U14326 (N_14326,N_10466,N_12069);
xnor U14327 (N_14327,N_11717,N_10211);
nand U14328 (N_14328,N_10873,N_10401);
and U14329 (N_14329,N_11368,N_11772);
or U14330 (N_14330,N_11630,N_10734);
nor U14331 (N_14331,N_10387,N_11479);
or U14332 (N_14332,N_11270,N_11166);
nor U14333 (N_14333,N_11437,N_10050);
nor U14334 (N_14334,N_11117,N_10384);
xor U14335 (N_14335,N_11046,N_10310);
nor U14336 (N_14336,N_11580,N_12377);
xor U14337 (N_14337,N_10123,N_10048);
or U14338 (N_14338,N_11632,N_12057);
xor U14339 (N_14339,N_12382,N_10916);
or U14340 (N_14340,N_11234,N_10182);
xnor U14341 (N_14341,N_10256,N_11382);
or U14342 (N_14342,N_11351,N_11483);
nand U14343 (N_14343,N_12141,N_11050);
xnor U14344 (N_14344,N_11194,N_11572);
nor U14345 (N_14345,N_11377,N_11282);
nand U14346 (N_14346,N_11998,N_10734);
and U14347 (N_14347,N_11279,N_11499);
nand U14348 (N_14348,N_11116,N_11795);
and U14349 (N_14349,N_11435,N_10541);
nand U14350 (N_14350,N_12289,N_11136);
or U14351 (N_14351,N_10182,N_10647);
or U14352 (N_14352,N_11661,N_10049);
xnor U14353 (N_14353,N_12289,N_10372);
xor U14354 (N_14354,N_11225,N_10008);
nand U14355 (N_14355,N_10744,N_10945);
nor U14356 (N_14356,N_10461,N_12375);
nand U14357 (N_14357,N_10652,N_11321);
or U14358 (N_14358,N_11789,N_10712);
nor U14359 (N_14359,N_10256,N_10516);
nand U14360 (N_14360,N_11439,N_11698);
and U14361 (N_14361,N_11562,N_10251);
nor U14362 (N_14362,N_11097,N_12465);
xnor U14363 (N_14363,N_11277,N_10325);
nor U14364 (N_14364,N_11603,N_10057);
or U14365 (N_14365,N_11415,N_11438);
xor U14366 (N_14366,N_10820,N_10055);
and U14367 (N_14367,N_11505,N_10162);
and U14368 (N_14368,N_10935,N_10264);
xnor U14369 (N_14369,N_11956,N_11084);
and U14370 (N_14370,N_10638,N_11641);
or U14371 (N_14371,N_10999,N_11684);
and U14372 (N_14372,N_12390,N_10246);
or U14373 (N_14373,N_11723,N_12485);
or U14374 (N_14374,N_10210,N_10540);
nor U14375 (N_14375,N_11307,N_10375);
or U14376 (N_14376,N_11297,N_10088);
nor U14377 (N_14377,N_10391,N_12314);
xor U14378 (N_14378,N_11176,N_10884);
nand U14379 (N_14379,N_12417,N_11014);
nand U14380 (N_14380,N_12206,N_12441);
nand U14381 (N_14381,N_12116,N_11207);
or U14382 (N_14382,N_12292,N_10191);
or U14383 (N_14383,N_12452,N_10014);
nor U14384 (N_14384,N_12059,N_11880);
and U14385 (N_14385,N_10627,N_10117);
or U14386 (N_14386,N_10752,N_11237);
xor U14387 (N_14387,N_10450,N_10579);
nor U14388 (N_14388,N_12479,N_12315);
and U14389 (N_14389,N_11224,N_12288);
and U14390 (N_14390,N_10677,N_11442);
nand U14391 (N_14391,N_12276,N_12182);
nand U14392 (N_14392,N_11052,N_11706);
and U14393 (N_14393,N_10763,N_10944);
nand U14394 (N_14394,N_10541,N_11410);
xor U14395 (N_14395,N_12483,N_12270);
nor U14396 (N_14396,N_12095,N_12441);
xnor U14397 (N_14397,N_10090,N_10194);
nor U14398 (N_14398,N_10433,N_12499);
xor U14399 (N_14399,N_11170,N_10898);
nand U14400 (N_14400,N_11701,N_11784);
and U14401 (N_14401,N_10880,N_11430);
xor U14402 (N_14402,N_10038,N_10059);
or U14403 (N_14403,N_11921,N_12419);
xor U14404 (N_14404,N_10560,N_11765);
and U14405 (N_14405,N_10714,N_10092);
xnor U14406 (N_14406,N_10911,N_10180);
nor U14407 (N_14407,N_10900,N_10477);
or U14408 (N_14408,N_10736,N_10922);
nand U14409 (N_14409,N_10496,N_11604);
xor U14410 (N_14410,N_10645,N_10196);
and U14411 (N_14411,N_11423,N_11441);
nor U14412 (N_14412,N_10041,N_12151);
xnor U14413 (N_14413,N_12303,N_11084);
nand U14414 (N_14414,N_12307,N_11223);
nor U14415 (N_14415,N_10959,N_10201);
and U14416 (N_14416,N_11508,N_12231);
nand U14417 (N_14417,N_12268,N_11017);
xor U14418 (N_14418,N_11085,N_11707);
nand U14419 (N_14419,N_11765,N_11160);
or U14420 (N_14420,N_10438,N_11995);
and U14421 (N_14421,N_10727,N_10971);
and U14422 (N_14422,N_12161,N_12420);
or U14423 (N_14423,N_10203,N_11947);
xor U14424 (N_14424,N_10278,N_10042);
xnor U14425 (N_14425,N_10891,N_11235);
or U14426 (N_14426,N_11322,N_11439);
xnor U14427 (N_14427,N_10848,N_12332);
xnor U14428 (N_14428,N_10009,N_11609);
xor U14429 (N_14429,N_12009,N_11374);
xor U14430 (N_14430,N_11286,N_11792);
nand U14431 (N_14431,N_12134,N_12145);
nor U14432 (N_14432,N_11443,N_10427);
nor U14433 (N_14433,N_10484,N_10791);
nand U14434 (N_14434,N_10727,N_10981);
and U14435 (N_14435,N_10580,N_11602);
and U14436 (N_14436,N_12325,N_12467);
xor U14437 (N_14437,N_11530,N_11255);
nand U14438 (N_14438,N_10278,N_10195);
or U14439 (N_14439,N_10725,N_10751);
nand U14440 (N_14440,N_10470,N_10068);
nor U14441 (N_14441,N_11349,N_10511);
or U14442 (N_14442,N_10291,N_12049);
and U14443 (N_14443,N_10736,N_10111);
nor U14444 (N_14444,N_12400,N_11590);
nand U14445 (N_14445,N_10925,N_11007);
and U14446 (N_14446,N_10216,N_11855);
or U14447 (N_14447,N_11248,N_10702);
and U14448 (N_14448,N_11723,N_12298);
or U14449 (N_14449,N_11656,N_10045);
nor U14450 (N_14450,N_10835,N_12498);
nor U14451 (N_14451,N_10909,N_11502);
xor U14452 (N_14452,N_10365,N_12018);
xnor U14453 (N_14453,N_10457,N_12086);
nor U14454 (N_14454,N_11544,N_10884);
nand U14455 (N_14455,N_12485,N_11404);
nand U14456 (N_14456,N_10722,N_10610);
nand U14457 (N_14457,N_12292,N_12147);
or U14458 (N_14458,N_10993,N_10283);
nand U14459 (N_14459,N_12169,N_11235);
xnor U14460 (N_14460,N_10616,N_11549);
xnor U14461 (N_14461,N_11863,N_12062);
nand U14462 (N_14462,N_11201,N_10393);
nor U14463 (N_14463,N_11464,N_10465);
and U14464 (N_14464,N_11223,N_10493);
xor U14465 (N_14465,N_11108,N_10684);
and U14466 (N_14466,N_11938,N_11614);
and U14467 (N_14467,N_10710,N_12467);
nor U14468 (N_14468,N_11044,N_12383);
and U14469 (N_14469,N_10199,N_11104);
or U14470 (N_14470,N_12198,N_11739);
and U14471 (N_14471,N_10948,N_10027);
xnor U14472 (N_14472,N_10954,N_12402);
nor U14473 (N_14473,N_11421,N_10827);
xor U14474 (N_14474,N_11425,N_11688);
nor U14475 (N_14475,N_11324,N_12131);
and U14476 (N_14476,N_10803,N_11175);
or U14477 (N_14477,N_10698,N_10776);
and U14478 (N_14478,N_11015,N_11818);
xnor U14479 (N_14479,N_12195,N_11451);
and U14480 (N_14480,N_11907,N_12478);
nand U14481 (N_14481,N_12407,N_12450);
nand U14482 (N_14482,N_10522,N_12053);
nor U14483 (N_14483,N_10452,N_11149);
and U14484 (N_14484,N_11222,N_10411);
or U14485 (N_14485,N_10290,N_11273);
and U14486 (N_14486,N_11151,N_10024);
nor U14487 (N_14487,N_11924,N_10585);
nor U14488 (N_14488,N_10890,N_11918);
nor U14489 (N_14489,N_10492,N_10115);
xor U14490 (N_14490,N_11398,N_10120);
xnor U14491 (N_14491,N_11855,N_11367);
nand U14492 (N_14492,N_10817,N_11065);
nor U14493 (N_14493,N_11331,N_10249);
xor U14494 (N_14494,N_11891,N_11184);
or U14495 (N_14495,N_10884,N_12049);
nand U14496 (N_14496,N_11800,N_12496);
xor U14497 (N_14497,N_11240,N_12037);
nor U14498 (N_14498,N_10292,N_10232);
nor U14499 (N_14499,N_10542,N_11558);
nand U14500 (N_14500,N_11174,N_12284);
nand U14501 (N_14501,N_10194,N_11062);
or U14502 (N_14502,N_10172,N_11964);
and U14503 (N_14503,N_10406,N_12343);
xor U14504 (N_14504,N_10426,N_10477);
or U14505 (N_14505,N_11151,N_10308);
nand U14506 (N_14506,N_12487,N_11695);
xor U14507 (N_14507,N_11560,N_11457);
nor U14508 (N_14508,N_10229,N_12360);
or U14509 (N_14509,N_11943,N_10951);
and U14510 (N_14510,N_11784,N_12471);
xor U14511 (N_14511,N_10373,N_10372);
nand U14512 (N_14512,N_12265,N_10504);
nand U14513 (N_14513,N_12321,N_10446);
nor U14514 (N_14514,N_11486,N_11163);
or U14515 (N_14515,N_11914,N_11140);
xnor U14516 (N_14516,N_11987,N_10119);
nor U14517 (N_14517,N_11513,N_10268);
and U14518 (N_14518,N_11372,N_10138);
or U14519 (N_14519,N_11819,N_11258);
or U14520 (N_14520,N_12291,N_10978);
nor U14521 (N_14521,N_10759,N_12195);
or U14522 (N_14522,N_12343,N_12448);
nor U14523 (N_14523,N_10743,N_12112);
nor U14524 (N_14524,N_11844,N_11980);
nand U14525 (N_14525,N_11616,N_11842);
nor U14526 (N_14526,N_10511,N_12063);
and U14527 (N_14527,N_10283,N_10650);
nand U14528 (N_14528,N_11913,N_11395);
nand U14529 (N_14529,N_10364,N_12350);
and U14530 (N_14530,N_11318,N_11714);
nand U14531 (N_14531,N_10158,N_10265);
or U14532 (N_14532,N_10022,N_10370);
nor U14533 (N_14533,N_10623,N_10910);
nand U14534 (N_14534,N_12136,N_11448);
and U14535 (N_14535,N_10758,N_11018);
xor U14536 (N_14536,N_10739,N_10981);
and U14537 (N_14537,N_10877,N_10611);
nor U14538 (N_14538,N_11975,N_11515);
xnor U14539 (N_14539,N_10614,N_12448);
nor U14540 (N_14540,N_11255,N_10560);
nand U14541 (N_14541,N_11954,N_10557);
nand U14542 (N_14542,N_12153,N_10968);
xor U14543 (N_14543,N_10330,N_10928);
xor U14544 (N_14544,N_11544,N_12185);
nor U14545 (N_14545,N_10592,N_12442);
and U14546 (N_14546,N_12071,N_10369);
or U14547 (N_14547,N_12341,N_10050);
nand U14548 (N_14548,N_11876,N_12313);
or U14549 (N_14549,N_12119,N_11587);
nor U14550 (N_14550,N_10320,N_12012);
and U14551 (N_14551,N_12299,N_11997);
and U14552 (N_14552,N_11112,N_11039);
nor U14553 (N_14553,N_11282,N_11883);
or U14554 (N_14554,N_11368,N_11832);
nand U14555 (N_14555,N_12142,N_12249);
xor U14556 (N_14556,N_11812,N_12326);
or U14557 (N_14557,N_11142,N_10781);
xnor U14558 (N_14558,N_11782,N_11002);
xor U14559 (N_14559,N_11092,N_12461);
and U14560 (N_14560,N_10519,N_12396);
xnor U14561 (N_14561,N_10089,N_10531);
and U14562 (N_14562,N_11327,N_11601);
or U14563 (N_14563,N_11730,N_12476);
nand U14564 (N_14564,N_12110,N_10458);
nand U14565 (N_14565,N_10613,N_10662);
nor U14566 (N_14566,N_10631,N_12078);
nand U14567 (N_14567,N_10500,N_11950);
nor U14568 (N_14568,N_11774,N_10038);
nand U14569 (N_14569,N_11864,N_10462);
xor U14570 (N_14570,N_10320,N_10292);
and U14571 (N_14571,N_10259,N_10012);
xor U14572 (N_14572,N_12431,N_11640);
nor U14573 (N_14573,N_12169,N_12205);
and U14574 (N_14574,N_10918,N_11358);
xor U14575 (N_14575,N_10720,N_10199);
or U14576 (N_14576,N_12165,N_12323);
and U14577 (N_14577,N_11551,N_11594);
nor U14578 (N_14578,N_11967,N_12335);
nor U14579 (N_14579,N_10512,N_10443);
nor U14580 (N_14580,N_10413,N_11515);
nand U14581 (N_14581,N_10126,N_10426);
nor U14582 (N_14582,N_12161,N_10793);
xor U14583 (N_14583,N_11074,N_11950);
nand U14584 (N_14584,N_11058,N_11677);
xor U14585 (N_14585,N_11409,N_11625);
nor U14586 (N_14586,N_10727,N_10147);
or U14587 (N_14587,N_12493,N_12459);
and U14588 (N_14588,N_11702,N_12184);
and U14589 (N_14589,N_11666,N_11263);
nor U14590 (N_14590,N_12074,N_10392);
or U14591 (N_14591,N_10500,N_11098);
xnor U14592 (N_14592,N_11927,N_10523);
nor U14593 (N_14593,N_10690,N_12295);
or U14594 (N_14594,N_12051,N_12115);
nor U14595 (N_14595,N_11534,N_10142);
nor U14596 (N_14596,N_10441,N_10009);
or U14597 (N_14597,N_11095,N_11072);
nor U14598 (N_14598,N_11015,N_11613);
xor U14599 (N_14599,N_12030,N_11914);
and U14600 (N_14600,N_10530,N_10475);
nand U14601 (N_14601,N_10477,N_10576);
nor U14602 (N_14602,N_10707,N_10594);
and U14603 (N_14603,N_11578,N_11569);
xor U14604 (N_14604,N_12099,N_12199);
xnor U14605 (N_14605,N_12224,N_10013);
nor U14606 (N_14606,N_11410,N_10591);
or U14607 (N_14607,N_11545,N_10635);
and U14608 (N_14608,N_11625,N_10128);
xor U14609 (N_14609,N_10388,N_10865);
or U14610 (N_14610,N_10069,N_11771);
or U14611 (N_14611,N_10763,N_11496);
nand U14612 (N_14612,N_12184,N_10637);
or U14613 (N_14613,N_11642,N_11038);
xor U14614 (N_14614,N_11361,N_10079);
nor U14615 (N_14615,N_11938,N_11013);
nand U14616 (N_14616,N_12336,N_11440);
and U14617 (N_14617,N_12478,N_11718);
nor U14618 (N_14618,N_12123,N_10912);
and U14619 (N_14619,N_10111,N_10998);
nand U14620 (N_14620,N_11858,N_12336);
or U14621 (N_14621,N_12234,N_11787);
nand U14622 (N_14622,N_11054,N_11001);
xor U14623 (N_14623,N_11881,N_11388);
nand U14624 (N_14624,N_12283,N_10853);
xor U14625 (N_14625,N_11864,N_11585);
and U14626 (N_14626,N_11183,N_10145);
nand U14627 (N_14627,N_10022,N_11134);
or U14628 (N_14628,N_10394,N_11737);
nor U14629 (N_14629,N_11903,N_12222);
or U14630 (N_14630,N_11912,N_10558);
and U14631 (N_14631,N_11720,N_10429);
or U14632 (N_14632,N_10504,N_11354);
nand U14633 (N_14633,N_12388,N_11458);
nand U14634 (N_14634,N_11627,N_11250);
nand U14635 (N_14635,N_10563,N_10950);
nand U14636 (N_14636,N_11572,N_10358);
xnor U14637 (N_14637,N_11511,N_10810);
xor U14638 (N_14638,N_11640,N_12453);
xnor U14639 (N_14639,N_10918,N_10849);
nor U14640 (N_14640,N_10233,N_11828);
and U14641 (N_14641,N_11712,N_10054);
xnor U14642 (N_14642,N_11074,N_11073);
xnor U14643 (N_14643,N_12119,N_10342);
nand U14644 (N_14644,N_10505,N_12132);
and U14645 (N_14645,N_11366,N_11585);
and U14646 (N_14646,N_10413,N_11571);
nor U14647 (N_14647,N_10225,N_10755);
and U14648 (N_14648,N_12411,N_10143);
or U14649 (N_14649,N_10435,N_11309);
nand U14650 (N_14650,N_10165,N_11400);
or U14651 (N_14651,N_10758,N_11302);
and U14652 (N_14652,N_11244,N_12136);
xor U14653 (N_14653,N_12126,N_10572);
and U14654 (N_14654,N_10205,N_11513);
nand U14655 (N_14655,N_11590,N_12065);
or U14656 (N_14656,N_11106,N_10029);
nor U14657 (N_14657,N_11526,N_11597);
and U14658 (N_14658,N_11600,N_11438);
xnor U14659 (N_14659,N_12463,N_11438);
and U14660 (N_14660,N_11239,N_12013);
nor U14661 (N_14661,N_11998,N_12381);
nand U14662 (N_14662,N_12121,N_10217);
nor U14663 (N_14663,N_11944,N_11965);
nor U14664 (N_14664,N_11424,N_12242);
or U14665 (N_14665,N_11056,N_10969);
and U14666 (N_14666,N_10473,N_11641);
xnor U14667 (N_14667,N_10234,N_11168);
or U14668 (N_14668,N_10478,N_11411);
or U14669 (N_14669,N_10547,N_10334);
nand U14670 (N_14670,N_11567,N_10402);
nor U14671 (N_14671,N_12112,N_10720);
and U14672 (N_14672,N_11218,N_11921);
or U14673 (N_14673,N_11749,N_11186);
nor U14674 (N_14674,N_12304,N_12248);
and U14675 (N_14675,N_11511,N_11324);
and U14676 (N_14676,N_12174,N_12140);
xnor U14677 (N_14677,N_11319,N_10434);
and U14678 (N_14678,N_11161,N_12397);
or U14679 (N_14679,N_11664,N_10218);
and U14680 (N_14680,N_10181,N_12256);
and U14681 (N_14681,N_10840,N_12307);
nor U14682 (N_14682,N_12076,N_11599);
and U14683 (N_14683,N_11632,N_11606);
nand U14684 (N_14684,N_12311,N_10697);
and U14685 (N_14685,N_11706,N_11426);
nand U14686 (N_14686,N_11844,N_10608);
xnor U14687 (N_14687,N_11628,N_11800);
xor U14688 (N_14688,N_10940,N_10020);
nor U14689 (N_14689,N_11591,N_10796);
nand U14690 (N_14690,N_11707,N_10171);
xor U14691 (N_14691,N_11733,N_11965);
and U14692 (N_14692,N_10148,N_11445);
nor U14693 (N_14693,N_10110,N_11851);
and U14694 (N_14694,N_10799,N_11535);
nor U14695 (N_14695,N_11808,N_10759);
or U14696 (N_14696,N_10095,N_10426);
and U14697 (N_14697,N_10358,N_11131);
nand U14698 (N_14698,N_10113,N_10822);
and U14699 (N_14699,N_10526,N_10832);
nor U14700 (N_14700,N_11379,N_11444);
or U14701 (N_14701,N_11553,N_11477);
xnor U14702 (N_14702,N_11214,N_12380);
xor U14703 (N_14703,N_11085,N_10828);
xor U14704 (N_14704,N_11539,N_11843);
or U14705 (N_14705,N_11973,N_10244);
nor U14706 (N_14706,N_11356,N_10290);
and U14707 (N_14707,N_12203,N_10964);
and U14708 (N_14708,N_10184,N_10275);
and U14709 (N_14709,N_11840,N_12099);
xor U14710 (N_14710,N_11167,N_10360);
nand U14711 (N_14711,N_12362,N_12108);
or U14712 (N_14712,N_12362,N_12267);
nand U14713 (N_14713,N_10502,N_10490);
nand U14714 (N_14714,N_10103,N_11450);
nor U14715 (N_14715,N_11862,N_11999);
xor U14716 (N_14716,N_11347,N_11066);
or U14717 (N_14717,N_10895,N_12022);
and U14718 (N_14718,N_11342,N_10186);
nor U14719 (N_14719,N_10518,N_10964);
and U14720 (N_14720,N_10163,N_12159);
xor U14721 (N_14721,N_11857,N_11650);
and U14722 (N_14722,N_12370,N_11013);
and U14723 (N_14723,N_11976,N_11952);
nand U14724 (N_14724,N_12265,N_10288);
nor U14725 (N_14725,N_12346,N_10770);
nor U14726 (N_14726,N_10245,N_11976);
and U14727 (N_14727,N_10631,N_11883);
and U14728 (N_14728,N_10815,N_11644);
or U14729 (N_14729,N_11286,N_11595);
xor U14730 (N_14730,N_11319,N_10478);
nand U14731 (N_14731,N_12214,N_10784);
nand U14732 (N_14732,N_11290,N_10051);
nor U14733 (N_14733,N_10255,N_12124);
or U14734 (N_14734,N_12026,N_10074);
and U14735 (N_14735,N_10083,N_11313);
xnor U14736 (N_14736,N_12067,N_10034);
and U14737 (N_14737,N_11169,N_12180);
nand U14738 (N_14738,N_12461,N_10686);
or U14739 (N_14739,N_10324,N_11277);
nand U14740 (N_14740,N_10842,N_11323);
nor U14741 (N_14741,N_10372,N_12027);
nand U14742 (N_14742,N_12197,N_12094);
xnor U14743 (N_14743,N_11955,N_12146);
xnor U14744 (N_14744,N_10851,N_10628);
xnor U14745 (N_14745,N_11591,N_10745);
nand U14746 (N_14746,N_11728,N_11351);
xnor U14747 (N_14747,N_10447,N_10055);
nand U14748 (N_14748,N_10520,N_10362);
or U14749 (N_14749,N_10996,N_10066);
nand U14750 (N_14750,N_10753,N_11157);
nor U14751 (N_14751,N_11158,N_12368);
xnor U14752 (N_14752,N_11699,N_12476);
xnor U14753 (N_14753,N_12063,N_10482);
or U14754 (N_14754,N_11986,N_10534);
nor U14755 (N_14755,N_11579,N_11802);
nor U14756 (N_14756,N_10414,N_12451);
nand U14757 (N_14757,N_10572,N_10159);
and U14758 (N_14758,N_10758,N_10769);
nor U14759 (N_14759,N_10907,N_11607);
and U14760 (N_14760,N_10207,N_11609);
nor U14761 (N_14761,N_10547,N_10138);
and U14762 (N_14762,N_10216,N_10480);
xor U14763 (N_14763,N_11937,N_10427);
xor U14764 (N_14764,N_12428,N_11704);
nand U14765 (N_14765,N_10469,N_11708);
nand U14766 (N_14766,N_11725,N_12154);
and U14767 (N_14767,N_11641,N_11901);
nor U14768 (N_14768,N_11851,N_10626);
nand U14769 (N_14769,N_10223,N_11241);
or U14770 (N_14770,N_12463,N_12024);
or U14771 (N_14771,N_11182,N_10796);
nand U14772 (N_14772,N_12048,N_10969);
and U14773 (N_14773,N_11654,N_11854);
and U14774 (N_14774,N_11486,N_11465);
and U14775 (N_14775,N_12338,N_11764);
nand U14776 (N_14776,N_10611,N_12216);
and U14777 (N_14777,N_11653,N_10088);
and U14778 (N_14778,N_11445,N_10899);
nor U14779 (N_14779,N_12218,N_12242);
and U14780 (N_14780,N_10145,N_11940);
or U14781 (N_14781,N_10248,N_11116);
nand U14782 (N_14782,N_12315,N_11077);
or U14783 (N_14783,N_11864,N_11798);
nor U14784 (N_14784,N_10582,N_10854);
or U14785 (N_14785,N_10134,N_12117);
xnor U14786 (N_14786,N_11180,N_10631);
and U14787 (N_14787,N_10228,N_10058);
nor U14788 (N_14788,N_11558,N_11212);
and U14789 (N_14789,N_10795,N_11638);
xnor U14790 (N_14790,N_10885,N_10131);
or U14791 (N_14791,N_11486,N_12111);
or U14792 (N_14792,N_12021,N_10430);
or U14793 (N_14793,N_10669,N_10474);
xnor U14794 (N_14794,N_11431,N_11948);
nand U14795 (N_14795,N_10419,N_10706);
nor U14796 (N_14796,N_12027,N_11574);
and U14797 (N_14797,N_11971,N_12208);
xnor U14798 (N_14798,N_11943,N_12460);
xor U14799 (N_14799,N_10974,N_11684);
xor U14800 (N_14800,N_10696,N_12478);
and U14801 (N_14801,N_10568,N_12350);
xor U14802 (N_14802,N_12078,N_11985);
and U14803 (N_14803,N_11416,N_11466);
and U14804 (N_14804,N_10066,N_10685);
xnor U14805 (N_14805,N_11659,N_12445);
nand U14806 (N_14806,N_10369,N_10022);
xor U14807 (N_14807,N_10708,N_11847);
nor U14808 (N_14808,N_11618,N_10486);
nor U14809 (N_14809,N_10621,N_11653);
and U14810 (N_14810,N_11057,N_12368);
nand U14811 (N_14811,N_11259,N_10935);
xnor U14812 (N_14812,N_11134,N_11898);
and U14813 (N_14813,N_11189,N_12412);
nor U14814 (N_14814,N_11779,N_12196);
xnor U14815 (N_14815,N_11830,N_10030);
or U14816 (N_14816,N_11350,N_10374);
and U14817 (N_14817,N_11412,N_10392);
nor U14818 (N_14818,N_11655,N_12197);
or U14819 (N_14819,N_10881,N_11593);
nor U14820 (N_14820,N_11380,N_10625);
nor U14821 (N_14821,N_10093,N_10241);
or U14822 (N_14822,N_12301,N_11667);
xnor U14823 (N_14823,N_11879,N_10956);
xor U14824 (N_14824,N_11657,N_10920);
nor U14825 (N_14825,N_11396,N_10154);
or U14826 (N_14826,N_12295,N_11993);
and U14827 (N_14827,N_11011,N_10632);
xor U14828 (N_14828,N_11683,N_10666);
xor U14829 (N_14829,N_12495,N_10376);
nor U14830 (N_14830,N_12498,N_10502);
xnor U14831 (N_14831,N_11423,N_10531);
or U14832 (N_14832,N_11055,N_11315);
nor U14833 (N_14833,N_10578,N_11103);
nand U14834 (N_14834,N_11519,N_10501);
or U14835 (N_14835,N_10674,N_12128);
and U14836 (N_14836,N_10118,N_10870);
and U14837 (N_14837,N_10606,N_11560);
or U14838 (N_14838,N_10244,N_10686);
or U14839 (N_14839,N_11698,N_10501);
xnor U14840 (N_14840,N_11753,N_12387);
and U14841 (N_14841,N_10510,N_10158);
and U14842 (N_14842,N_11237,N_11607);
nand U14843 (N_14843,N_11800,N_12346);
nand U14844 (N_14844,N_11089,N_11291);
or U14845 (N_14845,N_12493,N_10287);
and U14846 (N_14846,N_11013,N_10509);
xor U14847 (N_14847,N_11695,N_10133);
or U14848 (N_14848,N_11625,N_12025);
nor U14849 (N_14849,N_11266,N_10300);
nand U14850 (N_14850,N_10371,N_10989);
xnor U14851 (N_14851,N_12314,N_10717);
or U14852 (N_14852,N_11156,N_11612);
xnor U14853 (N_14853,N_10377,N_11058);
or U14854 (N_14854,N_12297,N_10036);
and U14855 (N_14855,N_10241,N_11054);
nor U14856 (N_14856,N_12250,N_11000);
nor U14857 (N_14857,N_11513,N_11331);
xor U14858 (N_14858,N_10713,N_10940);
nor U14859 (N_14859,N_10548,N_10807);
nor U14860 (N_14860,N_11090,N_11561);
and U14861 (N_14861,N_10287,N_10377);
xnor U14862 (N_14862,N_10271,N_11809);
xor U14863 (N_14863,N_10779,N_10491);
xnor U14864 (N_14864,N_10031,N_10688);
and U14865 (N_14865,N_10780,N_12005);
xnor U14866 (N_14866,N_10544,N_11999);
nor U14867 (N_14867,N_11113,N_10942);
or U14868 (N_14868,N_11351,N_12182);
xor U14869 (N_14869,N_12083,N_11924);
xnor U14870 (N_14870,N_11586,N_12491);
xor U14871 (N_14871,N_12212,N_12331);
nand U14872 (N_14872,N_11763,N_10233);
nor U14873 (N_14873,N_10461,N_10066);
nor U14874 (N_14874,N_11923,N_10710);
and U14875 (N_14875,N_11090,N_10398);
or U14876 (N_14876,N_10471,N_10388);
nor U14877 (N_14877,N_11899,N_12383);
and U14878 (N_14878,N_10124,N_10331);
or U14879 (N_14879,N_11580,N_12048);
nand U14880 (N_14880,N_12203,N_10676);
xnor U14881 (N_14881,N_11063,N_11259);
or U14882 (N_14882,N_11576,N_12219);
and U14883 (N_14883,N_11258,N_11180);
nand U14884 (N_14884,N_11269,N_10269);
nand U14885 (N_14885,N_10733,N_10767);
nand U14886 (N_14886,N_11381,N_10275);
nand U14887 (N_14887,N_11718,N_12319);
xor U14888 (N_14888,N_11511,N_10570);
nand U14889 (N_14889,N_10550,N_12427);
nand U14890 (N_14890,N_11818,N_11196);
nand U14891 (N_14891,N_11476,N_10083);
or U14892 (N_14892,N_11585,N_11588);
and U14893 (N_14893,N_10817,N_12283);
nor U14894 (N_14894,N_11109,N_10915);
or U14895 (N_14895,N_11803,N_10425);
and U14896 (N_14896,N_11253,N_10971);
and U14897 (N_14897,N_12117,N_10230);
or U14898 (N_14898,N_11738,N_12102);
and U14899 (N_14899,N_11855,N_10636);
and U14900 (N_14900,N_10194,N_11822);
nand U14901 (N_14901,N_10389,N_11771);
nor U14902 (N_14902,N_10782,N_12493);
xnor U14903 (N_14903,N_11223,N_12493);
xnor U14904 (N_14904,N_10033,N_10470);
xnor U14905 (N_14905,N_12158,N_10452);
or U14906 (N_14906,N_11140,N_10955);
nand U14907 (N_14907,N_11071,N_11023);
and U14908 (N_14908,N_11801,N_11232);
and U14909 (N_14909,N_10003,N_10442);
nand U14910 (N_14910,N_10370,N_11444);
or U14911 (N_14911,N_12338,N_11789);
nor U14912 (N_14912,N_12387,N_11425);
and U14913 (N_14913,N_11293,N_10706);
nor U14914 (N_14914,N_11154,N_10780);
nor U14915 (N_14915,N_12260,N_12480);
and U14916 (N_14916,N_11434,N_11715);
or U14917 (N_14917,N_12252,N_11631);
xnor U14918 (N_14918,N_11105,N_11394);
nor U14919 (N_14919,N_11714,N_10210);
nor U14920 (N_14920,N_10612,N_11138);
nand U14921 (N_14921,N_12166,N_10247);
or U14922 (N_14922,N_10110,N_11784);
xnor U14923 (N_14923,N_12268,N_11000);
xor U14924 (N_14924,N_11504,N_12324);
and U14925 (N_14925,N_11874,N_11285);
nor U14926 (N_14926,N_10036,N_11712);
nand U14927 (N_14927,N_11013,N_11484);
xor U14928 (N_14928,N_10382,N_11163);
nand U14929 (N_14929,N_10476,N_10334);
nand U14930 (N_14930,N_11408,N_11977);
or U14931 (N_14931,N_11283,N_10244);
xnor U14932 (N_14932,N_10388,N_10015);
nor U14933 (N_14933,N_10354,N_11441);
or U14934 (N_14934,N_11081,N_10680);
xor U14935 (N_14935,N_11465,N_10623);
nor U14936 (N_14936,N_10103,N_11046);
and U14937 (N_14937,N_11203,N_12252);
nor U14938 (N_14938,N_10308,N_12269);
nor U14939 (N_14939,N_11154,N_11701);
nand U14940 (N_14940,N_10260,N_10656);
nor U14941 (N_14941,N_10871,N_11308);
xor U14942 (N_14942,N_10496,N_12117);
nor U14943 (N_14943,N_10074,N_11926);
nor U14944 (N_14944,N_10131,N_10827);
xnor U14945 (N_14945,N_10945,N_10503);
xor U14946 (N_14946,N_10474,N_10687);
xor U14947 (N_14947,N_12024,N_10298);
and U14948 (N_14948,N_10427,N_12241);
or U14949 (N_14949,N_10214,N_12252);
nor U14950 (N_14950,N_10487,N_11268);
or U14951 (N_14951,N_11638,N_10148);
and U14952 (N_14952,N_12460,N_12469);
and U14953 (N_14953,N_10726,N_10873);
or U14954 (N_14954,N_10376,N_11879);
nor U14955 (N_14955,N_10862,N_12207);
xnor U14956 (N_14956,N_10001,N_11011);
nand U14957 (N_14957,N_10338,N_11225);
xor U14958 (N_14958,N_11646,N_12008);
xnor U14959 (N_14959,N_12284,N_11746);
nand U14960 (N_14960,N_10091,N_11554);
nor U14961 (N_14961,N_12119,N_12022);
nor U14962 (N_14962,N_10623,N_11408);
nand U14963 (N_14963,N_11609,N_11320);
xnor U14964 (N_14964,N_11081,N_10293);
nor U14965 (N_14965,N_11215,N_10069);
xnor U14966 (N_14966,N_12078,N_11653);
nor U14967 (N_14967,N_10053,N_10928);
and U14968 (N_14968,N_11488,N_12129);
or U14969 (N_14969,N_10870,N_10415);
nand U14970 (N_14970,N_10007,N_10723);
and U14971 (N_14971,N_10767,N_10272);
xor U14972 (N_14972,N_12295,N_11378);
nand U14973 (N_14973,N_10325,N_11303);
and U14974 (N_14974,N_11263,N_10987);
nand U14975 (N_14975,N_12475,N_11676);
and U14976 (N_14976,N_11443,N_11225);
and U14977 (N_14977,N_11367,N_10275);
nor U14978 (N_14978,N_10420,N_12366);
and U14979 (N_14979,N_10515,N_11210);
and U14980 (N_14980,N_12489,N_11174);
xnor U14981 (N_14981,N_10537,N_11552);
nor U14982 (N_14982,N_12228,N_12152);
xnor U14983 (N_14983,N_10989,N_11651);
nor U14984 (N_14984,N_11301,N_10065);
nand U14985 (N_14985,N_12225,N_11064);
or U14986 (N_14986,N_10557,N_12288);
nor U14987 (N_14987,N_12337,N_12349);
xor U14988 (N_14988,N_12290,N_12319);
xor U14989 (N_14989,N_12251,N_11745);
or U14990 (N_14990,N_11686,N_11391);
and U14991 (N_14991,N_10259,N_10602);
and U14992 (N_14992,N_11133,N_10204);
xnor U14993 (N_14993,N_10913,N_11014);
nand U14994 (N_14994,N_11193,N_10360);
nor U14995 (N_14995,N_10243,N_10967);
nor U14996 (N_14996,N_11892,N_11767);
nand U14997 (N_14997,N_12109,N_11442);
or U14998 (N_14998,N_10016,N_11734);
nor U14999 (N_14999,N_10117,N_12442);
xor U15000 (N_15000,N_14073,N_13712);
nand U15001 (N_15001,N_14184,N_13189);
nor U15002 (N_15002,N_14898,N_13156);
xnor U15003 (N_15003,N_13181,N_13808);
nor U15004 (N_15004,N_13837,N_12634);
nand U15005 (N_15005,N_14534,N_14291);
nand U15006 (N_15006,N_14472,N_12756);
and U15007 (N_15007,N_12827,N_14607);
and U15008 (N_15008,N_13715,N_14144);
xor U15009 (N_15009,N_13240,N_13481);
and U15010 (N_15010,N_14127,N_14849);
nor U15011 (N_15011,N_13599,N_14005);
nor U15012 (N_15012,N_14589,N_14720);
nor U15013 (N_15013,N_13135,N_12943);
or U15014 (N_15014,N_14575,N_12895);
nor U15015 (N_15015,N_14738,N_12899);
nor U15016 (N_15016,N_13980,N_12721);
and U15017 (N_15017,N_12601,N_13755);
nor U15018 (N_15018,N_13816,N_13107);
nand U15019 (N_15019,N_13019,N_13640);
and U15020 (N_15020,N_13876,N_14043);
nor U15021 (N_15021,N_14775,N_13253);
xor U15022 (N_15022,N_14404,N_13138);
xor U15023 (N_15023,N_13539,N_13778);
xnor U15024 (N_15024,N_14927,N_12732);
xor U15025 (N_15025,N_13171,N_13942);
and U15026 (N_15026,N_14514,N_13681);
or U15027 (N_15027,N_13713,N_14094);
or U15028 (N_15028,N_14086,N_12906);
nor U15029 (N_15029,N_14429,N_14804);
xnor U15030 (N_15030,N_13070,N_12679);
or U15031 (N_15031,N_12521,N_12682);
and U15032 (N_15032,N_14106,N_13362);
xnor U15033 (N_15033,N_12954,N_14440);
and U15034 (N_15034,N_14822,N_14598);
xor U15035 (N_15035,N_14739,N_14956);
xnor U15036 (N_15036,N_13066,N_12700);
or U15037 (N_15037,N_13913,N_14207);
and U15038 (N_15038,N_14353,N_14177);
nand U15039 (N_15039,N_13044,N_13573);
or U15040 (N_15040,N_13245,N_13392);
nand U15041 (N_15041,N_13074,N_13443);
or U15042 (N_15042,N_13623,N_14085);
or U15043 (N_15043,N_14842,N_14277);
xor U15044 (N_15044,N_12828,N_12977);
or U15045 (N_15045,N_13215,N_12534);
xnor U15046 (N_15046,N_13738,N_13486);
xnor U15047 (N_15047,N_13807,N_12594);
and U15048 (N_15048,N_14134,N_13525);
nor U15049 (N_15049,N_13109,N_13519);
nor U15050 (N_15050,N_13055,N_13763);
nor U15051 (N_15051,N_14566,N_13062);
xnor U15052 (N_15052,N_12583,N_13842);
xor U15053 (N_15053,N_12597,N_14966);
and U15054 (N_15054,N_13923,N_13665);
and U15055 (N_15055,N_12595,N_13088);
nor U15056 (N_15056,N_14886,N_13933);
or U15057 (N_15057,N_13431,N_14868);
and U15058 (N_15058,N_14905,N_12872);
and U15059 (N_15059,N_14488,N_13436);
nor U15060 (N_15060,N_14345,N_14936);
nor U15061 (N_15061,N_14672,N_13534);
xnor U15062 (N_15062,N_12904,N_14707);
nor U15063 (N_15063,N_14046,N_12878);
nand U15064 (N_15064,N_13307,N_14202);
nand U15065 (N_15065,N_14585,N_13495);
nand U15066 (N_15066,N_13955,N_13321);
xor U15067 (N_15067,N_12946,N_13024);
and U15068 (N_15068,N_14968,N_14932);
xnor U15069 (N_15069,N_14253,N_13988);
or U15070 (N_15070,N_12739,N_14596);
nor U15071 (N_15071,N_13036,N_14301);
xnor U15072 (N_15072,N_14137,N_12754);
xor U15073 (N_15073,N_12608,N_13094);
or U15074 (N_15074,N_13317,N_12550);
nor U15075 (N_15075,N_14327,N_13375);
nor U15076 (N_15076,N_12777,N_13508);
nand U15077 (N_15077,N_13318,N_13149);
nor U15078 (N_15078,N_13590,N_12952);
xor U15079 (N_15079,N_13207,N_13475);
nor U15080 (N_15080,N_13790,N_14477);
nand U15081 (N_15081,N_13946,N_14881);
nor U15082 (N_15082,N_12549,N_14829);
xor U15083 (N_15083,N_13646,N_13717);
or U15084 (N_15084,N_13624,N_13775);
xnor U15085 (N_15085,N_14896,N_13878);
or U15086 (N_15086,N_14835,N_14568);
and U15087 (N_15087,N_13100,N_14728);
or U15088 (N_15088,N_13226,N_13006);
nor U15089 (N_15089,N_13602,N_12784);
or U15090 (N_15090,N_14119,N_14336);
nor U15091 (N_15091,N_12653,N_14518);
nor U15092 (N_15092,N_12651,N_14975);
nand U15093 (N_15093,N_12837,N_14870);
and U15094 (N_15094,N_14313,N_13448);
xor U15095 (N_15095,N_14104,N_13709);
and U15096 (N_15096,N_14805,N_14569);
and U15097 (N_15097,N_13160,N_12633);
nand U15098 (N_15098,N_13880,N_13735);
nand U15099 (N_15099,N_12706,N_14464);
nand U15100 (N_15100,N_14632,N_14764);
or U15101 (N_15101,N_13848,N_14325);
and U15102 (N_15102,N_12845,N_13956);
nand U15103 (N_15103,N_14729,N_14688);
xnor U15104 (N_15104,N_13246,N_12781);
nand U15105 (N_15105,N_13984,N_14330);
nor U15106 (N_15106,N_13881,N_14516);
nand U15107 (N_15107,N_14016,N_14690);
and U15108 (N_15108,N_12885,N_13161);
nor U15109 (N_15109,N_14268,N_14121);
nor U15110 (N_15110,N_12511,N_12888);
nand U15111 (N_15111,N_14480,N_14267);
xnor U15112 (N_15112,N_14957,N_14809);
and U15113 (N_15113,N_13982,N_14282);
nand U15114 (N_15114,N_13370,N_12585);
nor U15115 (N_15115,N_14733,N_12913);
or U15116 (N_15116,N_14722,N_13187);
nand U15117 (N_15117,N_13502,N_12935);
xnor U15118 (N_15118,N_13256,N_14639);
and U15119 (N_15119,N_12810,N_14546);
xor U15120 (N_15120,N_13708,N_14820);
and U15121 (N_15121,N_13470,N_14996);
nand U15122 (N_15122,N_14871,N_12570);
xnor U15123 (N_15123,N_13450,N_13991);
xnor U15124 (N_15124,N_14827,N_14597);
nor U15125 (N_15125,N_14387,N_12856);
nand U15126 (N_15126,N_13018,N_14080);
nor U15127 (N_15127,N_14053,N_14487);
or U15128 (N_15128,N_13582,N_13313);
xnor U15129 (N_15129,N_13934,N_12625);
and U15130 (N_15130,N_12582,N_12745);
nor U15131 (N_15131,N_14066,N_14882);
nand U15132 (N_15132,N_14269,N_14035);
and U15133 (N_15133,N_13581,N_13541);
nand U15134 (N_15134,N_14506,N_14993);
nor U15135 (N_15135,N_13858,N_14960);
nand U15136 (N_15136,N_13429,N_14679);
nor U15137 (N_15137,N_14825,N_14347);
and U15138 (N_15138,N_13061,N_13205);
xor U15139 (N_15139,N_13966,N_14232);
and U15140 (N_15140,N_12842,N_13437);
xor U15141 (N_15141,N_12751,N_14740);
xor U15142 (N_15142,N_13445,N_14060);
and U15143 (N_15143,N_13671,N_12799);
xor U15144 (N_15144,N_12510,N_13049);
nor U15145 (N_15145,N_14977,N_14941);
nand U15146 (N_15146,N_13041,N_12527);
nor U15147 (N_15147,N_13761,N_14236);
xor U15148 (N_15148,N_13521,N_12865);
and U15149 (N_15149,N_14348,N_14789);
or U15150 (N_15150,N_13585,N_12541);
and U15151 (N_15151,N_13556,N_13685);
xnor U15152 (N_15152,N_14608,N_14502);
nor U15153 (N_15153,N_12612,N_14390);
xor U15154 (N_15154,N_12978,N_12826);
or U15155 (N_15155,N_14640,N_14560);
nand U15156 (N_15156,N_14974,N_13554);
or U15157 (N_15157,N_13469,N_14408);
and U15158 (N_15158,N_14595,N_13907);
nand U15159 (N_15159,N_14479,N_13523);
or U15160 (N_15160,N_13059,N_14039);
or U15161 (N_15161,N_12726,N_14928);
or U15162 (N_15162,N_12795,N_13320);
nand U15163 (N_15163,N_13349,N_13103);
and U15164 (N_15164,N_14366,N_14492);
or U15165 (N_15165,N_13021,N_13089);
nand U15166 (N_15166,N_14337,N_13356);
and U15167 (N_15167,N_13048,N_14485);
and U15168 (N_15168,N_12602,N_12881);
nor U15169 (N_15169,N_13977,N_13015);
or U15170 (N_15170,N_12821,N_12868);
nand U15171 (N_15171,N_13308,N_13007);
xnor U15172 (N_15172,N_14671,N_13853);
or U15173 (N_15173,N_14208,N_13493);
and U15174 (N_15174,N_13310,N_13643);
and U15175 (N_15175,N_13672,N_13580);
nand U15176 (N_15176,N_14605,N_14675);
and U15177 (N_15177,N_13614,N_13434);
nor U15178 (N_15178,N_13522,N_13221);
and U15179 (N_15179,N_13082,N_13978);
nor U15180 (N_15180,N_14162,N_14055);
or U15181 (N_15181,N_14840,N_14493);
nand U15182 (N_15182,N_13770,N_13928);
xor U15183 (N_15183,N_13768,N_13260);
or U15184 (N_15184,N_14634,N_14624);
and U15185 (N_15185,N_13119,N_12723);
nand U15186 (N_15186,N_14403,N_14765);
and U15187 (N_15187,N_12686,N_12957);
or U15188 (N_15188,N_14792,N_14101);
nand U15189 (N_15189,N_13140,N_14475);
xor U15190 (N_15190,N_12643,N_12921);
and U15191 (N_15191,N_14258,N_13827);
nor U15192 (N_15192,N_12640,N_13458);
or U15193 (N_15193,N_12569,N_12728);
xnor U15194 (N_15194,N_13162,N_14854);
nor U15195 (N_15195,N_12814,N_13746);
xnor U15196 (N_15196,N_13121,N_13178);
or U15197 (N_15197,N_12623,N_14098);
xnor U15198 (N_15198,N_14581,N_13087);
xor U15199 (N_15199,N_14423,N_12849);
nor U15200 (N_15200,N_14368,N_13996);
nor U15201 (N_15201,N_14553,N_12769);
nor U15202 (N_15202,N_12554,N_14042);
and U15203 (N_15203,N_14287,N_12532);
xnor U15204 (N_15204,N_13306,N_12553);
nor U15205 (N_15205,N_14782,N_13097);
nand U15206 (N_15206,N_13824,N_14185);
and U15207 (N_15207,N_14445,N_13645);
or U15208 (N_15208,N_14242,N_12770);
and U15209 (N_15209,N_13455,N_14385);
and U15210 (N_15210,N_13981,N_13208);
nand U15211 (N_15211,N_12609,N_14572);
and U15212 (N_15212,N_13369,N_14548);
xor U15213 (N_15213,N_12563,N_13930);
or U15214 (N_15214,N_13417,N_13060);
or U15215 (N_15215,N_13249,N_13057);
nor U15216 (N_15216,N_13705,N_13845);
or U15217 (N_15217,N_14311,N_13504);
or U15218 (N_15218,N_12876,N_13673);
and U15219 (N_15219,N_14677,N_13424);
xnor U15220 (N_15220,N_13067,N_13091);
xor U15221 (N_15221,N_14384,N_13727);
nand U15222 (N_15222,N_13366,N_12650);
nand U15223 (N_15223,N_14401,N_14963);
nand U15224 (N_15224,N_14578,N_14685);
and U15225 (N_15225,N_13796,N_12871);
and U15226 (N_15226,N_14843,N_14939);
or U15227 (N_15227,N_13201,N_13284);
nor U15228 (N_15228,N_12681,N_13542);
and U15229 (N_15229,N_14525,N_13723);
and U15230 (N_15230,N_13740,N_13787);
or U15231 (N_15231,N_13127,N_14845);
xor U15232 (N_15232,N_13029,N_13315);
or U15233 (N_15233,N_14017,N_14419);
and U15234 (N_15234,N_14174,N_14248);
nor U15235 (N_15235,N_14441,N_13903);
nor U15236 (N_15236,N_14321,N_13346);
xor U15237 (N_15237,N_12956,N_13791);
nor U15238 (N_15238,N_14245,N_14997);
or U15239 (N_15239,N_13010,N_13871);
or U15240 (N_15240,N_14357,N_13304);
nor U15241 (N_15241,N_14083,N_12676);
or U15242 (N_15242,N_12970,N_13714);
and U15243 (N_15243,N_12808,N_13684);
and U15244 (N_15244,N_13028,N_13792);
or U15245 (N_15245,N_13446,N_12588);
nand U15246 (N_15246,N_13394,N_14826);
nor U15247 (N_15247,N_13077,N_14000);
nor U15248 (N_15248,N_14433,N_12517);
or U15249 (N_15249,N_14491,N_13471);
xor U15250 (N_15250,N_12704,N_13874);
nor U15251 (N_15251,N_14030,N_12546);
or U15252 (N_15252,N_14049,N_13002);
nand U15253 (N_15253,N_14618,N_14201);
or U15254 (N_15254,N_13551,N_13276);
or U15255 (N_15255,N_14784,N_13964);
nand U15256 (N_15256,N_14389,N_13479);
nand U15257 (N_15257,N_14079,N_14075);
and U15258 (N_15258,N_13299,N_13213);
nand U15259 (N_15259,N_13868,N_14584);
and U15260 (N_15260,N_14630,N_14413);
nor U15261 (N_15261,N_14527,N_13168);
xnor U15262 (N_15262,N_13997,N_12599);
nor U15263 (N_15263,N_13005,N_13258);
or U15264 (N_15264,N_12772,N_14355);
nor U15265 (N_15265,N_14743,N_14724);
nor U15266 (N_15266,N_14961,N_13707);
or U15267 (N_15267,N_13506,N_14734);
nand U15268 (N_15268,N_12657,N_13247);
nand U15269 (N_15269,N_14302,N_13562);
nand U15270 (N_15270,N_14887,N_14931);
or U15271 (N_15271,N_13352,N_13102);
xor U15272 (N_15272,N_14143,N_14594);
nand U15273 (N_15273,N_14367,N_12813);
nand U15274 (N_15274,N_14140,N_14539);
nor U15275 (N_15275,N_14542,N_12755);
nor U15276 (N_15276,N_13420,N_13179);
nand U15277 (N_15277,N_14278,N_14834);
xor U15278 (N_15278,N_13828,N_13209);
nor U15279 (N_15279,N_14863,N_12816);
xnor U15280 (N_15280,N_13090,N_14567);
and U15281 (N_15281,N_12938,N_14097);
xor U15282 (N_15282,N_13336,N_13578);
xnor U15283 (N_15283,N_12917,N_13721);
xor U15284 (N_15284,N_13527,N_14767);
or U15285 (N_15285,N_14266,N_13368);
or U15286 (N_15286,N_13850,N_13421);
and U15287 (N_15287,N_14217,N_13785);
nand U15288 (N_15288,N_13776,N_14274);
and U15289 (N_15289,N_13572,N_12961);
xnor U15290 (N_15290,N_13620,N_14836);
or U15291 (N_15291,N_13695,N_12874);
xor U15292 (N_15292,N_13012,N_12823);
and U15293 (N_15293,N_12836,N_13990);
nor U15294 (N_15294,N_14536,N_14785);
nand U15295 (N_15295,N_14744,N_14333);
nor U15296 (N_15296,N_13341,N_14293);
xnor U15297 (N_15297,N_14444,N_13425);
xor U15298 (N_15298,N_13638,N_14194);
nand U15299 (N_15299,N_12903,N_12819);
nor U15300 (N_15300,N_14806,N_14151);
nand U15301 (N_15301,N_14240,N_13043);
nand U15302 (N_15302,N_13490,N_13274);
nand U15303 (N_15303,N_13288,N_12565);
nor U15304 (N_15304,N_14796,N_14577);
xnor U15305 (N_15305,N_12984,N_14352);
or U15306 (N_15306,N_12670,N_12635);
xor U15307 (N_15307,N_14965,N_14591);
and U15308 (N_15308,N_12966,N_12782);
xnor U15309 (N_15309,N_12675,N_13969);
nand U15310 (N_15310,N_12998,N_13206);
nand U15311 (N_15311,N_13634,N_12951);
nor U15312 (N_15312,N_13388,N_13296);
and U15313 (N_15313,N_12668,N_14741);
nand U15314 (N_15314,N_14755,N_12844);
xnor U15315 (N_15315,N_14406,N_13217);
and U15316 (N_15316,N_12709,N_14727);
or U15317 (N_15317,N_12886,N_13548);
or U15318 (N_15318,N_12556,N_14793);
nand U15319 (N_15319,N_12516,N_12760);
nand U15320 (N_15320,N_14848,N_13952);
nor U15321 (N_15321,N_12815,N_13960);
or U15322 (N_15322,N_14486,N_13733);
nand U15323 (N_15323,N_12611,N_12501);
and U15324 (N_15324,N_14980,N_12829);
or U15325 (N_15325,N_12843,N_12729);
and U15326 (N_15326,N_12919,N_13657);
nor U15327 (N_15327,N_14521,N_13625);
or U15328 (N_15328,N_13322,N_13566);
or U15329 (N_15329,N_13945,N_14422);
and U15330 (N_15330,N_13937,N_13261);
and U15331 (N_15331,N_13574,N_14645);
and U15332 (N_15332,N_12765,N_12989);
and U15333 (N_15333,N_12860,N_13344);
xnor U15334 (N_15334,N_12900,N_13616);
or U15335 (N_15335,N_12524,N_13460);
xor U15336 (N_15336,N_14320,N_12735);
nand U15337 (N_15337,N_13153,N_13817);
nand U15338 (N_15338,N_13391,N_14821);
or U15339 (N_15339,N_14601,N_14658);
nand U15340 (N_15340,N_13718,N_13297);
and U15341 (N_15341,N_13766,N_12674);
nor U15342 (N_15342,N_13724,N_13563);
nor U15343 (N_15343,N_13901,N_14654);
or U15344 (N_15344,N_13697,N_13826);
nand U15345 (N_15345,N_13814,N_12936);
or U15346 (N_15346,N_14778,N_14118);
and U15347 (N_15347,N_14034,N_14716);
xnor U15348 (N_15348,N_13706,N_13414);
nor U15349 (N_15349,N_14620,N_13557);
and U15350 (N_15350,N_14100,N_14179);
or U15351 (N_15351,N_13216,N_13569);
and U15352 (N_15352,N_13503,N_13243);
and U15353 (N_15353,N_13423,N_13372);
and U15354 (N_15354,N_14289,N_14647);
or U15355 (N_15355,N_13360,N_13204);
and U15356 (N_15356,N_12867,N_13851);
nor U15357 (N_15357,N_12787,N_14978);
or U15358 (N_15358,N_14531,N_14702);
nor U15359 (N_15359,N_13642,N_13795);
xnor U15360 (N_15360,N_14431,N_14225);
nor U15361 (N_15361,N_13197,N_13759);
and U15362 (N_15362,N_12790,N_12548);
and U15363 (N_15363,N_13641,N_13540);
nand U15364 (N_15364,N_12560,N_13403);
nor U15365 (N_15365,N_13008,N_14081);
xor U15366 (N_15366,N_13799,N_14398);
or U15367 (N_15367,N_13914,N_14222);
xnor U15368 (N_15368,N_14467,N_12660);
xor U15369 (N_15369,N_14686,N_13176);
and U15370 (N_15370,N_13856,N_12536);
xnor U15371 (N_15371,N_13682,N_13658);
nor U15372 (N_15372,N_14633,N_14175);
and U15373 (N_15373,N_14196,N_13877);
or U15374 (N_15374,N_14522,N_12942);
xor U15375 (N_15375,N_13301,N_12622);
nor U15376 (N_15376,N_14582,N_12758);
nor U15377 (N_15377,N_14895,N_14211);
and U15378 (N_15378,N_12539,N_14865);
nand U15379 (N_15379,N_12776,N_13499);
and U15380 (N_15380,N_12547,N_14270);
and U15381 (N_15381,N_14169,N_14869);
nand U15382 (N_15382,N_12775,N_14517);
or U15383 (N_15383,N_14857,N_14948);
or U15384 (N_15384,N_14261,N_14994);
and U15385 (N_15385,N_14471,N_14470);
xnor U15386 (N_15386,N_13354,N_13038);
and U15387 (N_15387,N_13891,N_12927);
and U15388 (N_15388,N_13753,N_13374);
and U15389 (N_15389,N_12986,N_12805);
and U15390 (N_15390,N_14001,N_13225);
nand U15391 (N_15391,N_14761,N_12630);
or U15392 (N_15392,N_14923,N_14456);
and U15393 (N_15393,N_14197,N_14621);
nand U15394 (N_15394,N_14652,N_13804);
and U15395 (N_15395,N_14379,N_14354);
and U15396 (N_15396,N_13902,N_14953);
xnor U15397 (N_15397,N_14750,N_14603);
nand U15398 (N_15398,N_12944,N_12964);
or U15399 (N_15399,N_12576,N_13428);
nand U15400 (N_15400,N_14284,N_14942);
nor U15401 (N_15401,N_14280,N_13633);
nor U15402 (N_15402,N_14771,N_13269);
or U15403 (N_15403,N_12665,N_12981);
nand U15404 (N_15404,N_14713,N_13944);
nand U15405 (N_15405,N_14549,N_14565);
and U15406 (N_15406,N_12533,N_14275);
and U15407 (N_15407,N_13772,N_12901);
xor U15408 (N_15408,N_13741,N_13326);
xor U15409 (N_15409,N_14532,N_14847);
or U15410 (N_15410,N_14115,N_12680);
nand U15411 (N_15411,N_13841,N_13777);
xnor U15412 (N_15412,N_14984,N_13604);
and U15413 (N_15413,N_14797,N_14047);
or U15414 (N_15414,N_13133,N_14884);
or U15415 (N_15415,N_12786,N_14823);
or U15416 (N_15416,N_13251,N_13939);
or U15417 (N_15417,N_12544,N_13843);
xnor U15418 (N_15418,N_14123,N_14183);
and U15419 (N_15419,N_12531,N_13432);
nor U15420 (N_15420,N_13972,N_14204);
nand U15421 (N_15421,N_14428,N_14014);
nand U15422 (N_15422,N_14737,N_13295);
nor U15423 (N_15423,N_13917,N_13183);
nor U15424 (N_15424,N_14430,N_14970);
nor U15425 (N_15425,N_13520,N_13918);
or U15426 (N_15426,N_13611,N_13950);
nor U15427 (N_15427,N_13905,N_14851);
xnor U15428 (N_15428,N_14283,N_13789);
nand U15429 (N_15429,N_14766,N_13263);
and U15430 (N_15430,N_13679,N_14641);
nand U15431 (N_15431,N_14296,N_13603);
or U15432 (N_15432,N_13762,N_13806);
or U15433 (N_15433,N_14919,N_12789);
or U15434 (N_15434,N_13989,N_12694);
and U15435 (N_15435,N_14130,N_12962);
nand U15436 (N_15436,N_13266,N_12631);
xnor U15437 (N_15437,N_14526,N_13866);
or U15438 (N_15438,N_14816,N_13147);
xnor U15439 (N_15439,N_13512,N_14964);
nand U15440 (N_15440,N_13617,N_14171);
and U15441 (N_15441,N_13861,N_14341);
or U15442 (N_15442,N_13085,N_14853);
or U15443 (N_15443,N_13000,N_13017);
or U15444 (N_15444,N_14742,N_13919);
nand U15445 (N_15445,N_13302,N_14692);
xnor U15446 (N_15446,N_14650,N_14052);
xnor U15447 (N_15447,N_13080,N_14400);
and U15448 (N_15448,N_12822,N_13836);
nand U15449 (N_15449,N_14622,N_14375);
or U15450 (N_15450,N_13259,N_14704);
xor U15451 (N_15451,N_13750,N_13118);
nand U15452 (N_15452,N_14138,N_14719);
xnor U15453 (N_15453,N_14676,N_14091);
nand U15454 (N_15454,N_13922,N_13500);
or U15455 (N_15455,N_13154,N_14421);
or U15456 (N_15456,N_13340,N_14873);
nand U15457 (N_15457,N_13058,N_12526);
nor U15458 (N_15458,N_14051,N_14714);
and U15459 (N_15459,N_14831,N_14223);
and U15460 (N_15460,N_14959,N_13001);
nand U15461 (N_15461,N_14391,N_14880);
nor U15462 (N_15462,N_14382,N_13511);
and U15463 (N_15463,N_13860,N_12774);
xor U15464 (N_15464,N_12915,N_12696);
xnor U15465 (N_15465,N_13649,N_14399);
nor U15466 (N_15466,N_12930,N_13510);
or U15467 (N_15467,N_14180,N_14904);
and U15468 (N_15468,N_14316,N_14332);
and U15469 (N_15469,N_14856,N_14089);
or U15470 (N_15470,N_14528,N_13104);
nand U15471 (N_15471,N_13547,N_13351);
nand U15472 (N_15472,N_14044,N_13769);
xnor U15473 (N_15473,N_12830,N_13815);
xor U15474 (N_15474,N_12959,N_14219);
and U15475 (N_15475,N_13325,N_13889);
nor U15476 (N_15476,N_14288,N_13281);
and U15477 (N_15477,N_12863,N_12731);
nor U15478 (N_15478,N_14523,N_12642);
xnor U15479 (N_15479,N_14356,N_13892);
or U15480 (N_15480,N_13131,N_13254);
nand U15481 (N_15481,N_13968,N_14649);
nor U15482 (N_15482,N_14246,N_12991);
nand U15483 (N_15483,N_14988,N_14461);
and U15484 (N_15484,N_13887,N_14735);
and U15485 (N_15485,N_13821,N_14986);
or U15486 (N_15486,N_14718,N_13238);
and U15487 (N_15487,N_13378,N_13323);
xor U15488 (N_15488,N_13916,N_14371);
or U15489 (N_15489,N_13365,N_12649);
and U15490 (N_15490,N_13651,N_13331);
and U15491 (N_15491,N_13046,N_12708);
nor U15492 (N_15492,N_13289,N_13594);
and U15493 (N_15493,N_14732,N_14573);
and U15494 (N_15494,N_12687,N_14239);
and U15495 (N_15495,N_13014,N_13647);
nand U15496 (N_15496,N_13833,N_13275);
nand U15497 (N_15497,N_13742,N_12852);
nand U15498 (N_15498,N_13234,N_12551);
xor U15499 (N_15499,N_14450,N_13971);
nand U15500 (N_15500,N_14818,N_12841);
nor U15501 (N_15501,N_12949,N_14883);
or U15502 (N_15502,N_14125,N_13987);
or U15503 (N_15503,N_12727,N_13983);
nand U15504 (N_15504,N_14794,N_13380);
nor U15505 (N_15505,N_13128,N_14558);
and U15506 (N_15506,N_14770,N_14715);
nor U15507 (N_15507,N_13632,N_14411);
and U15508 (N_15508,N_13210,N_14373);
and U15509 (N_15509,N_14457,N_14260);
or U15510 (N_15510,N_13167,N_14272);
nand U15511 (N_15511,N_14551,N_14200);
or U15512 (N_15512,N_14310,N_13571);
nor U15513 (N_15513,N_14210,N_12506);
or U15514 (N_15514,N_14612,N_14407);
or U15515 (N_15515,N_13524,N_12697);
xor U15516 (N_15516,N_13600,N_14499);
or U15517 (N_15517,N_12923,N_14418);
and U15518 (N_15518,N_14338,N_14925);
or U15519 (N_15519,N_13567,N_13803);
and U15520 (N_15520,N_14380,N_14807);
and U15521 (N_15521,N_14946,N_14535);
and U15522 (N_15522,N_13098,N_12690);
nor U15523 (N_15523,N_13530,N_13400);
nand U15524 (N_15524,N_14420,N_13357);
nor U15525 (N_15525,N_12641,N_14078);
or U15526 (N_15526,N_13030,N_13533);
xnor U15527 (N_15527,N_14643,N_12990);
or U15528 (N_15528,N_12880,N_13045);
and U15529 (N_15529,N_13381,N_14076);
xnor U15530 (N_15530,N_13442,N_13319);
or U15531 (N_15531,N_13644,N_14547);
nor U15532 (N_15532,N_14828,N_13056);
and U15533 (N_15533,N_12911,N_13823);
xor U15534 (N_15534,N_13630,N_14082);
and U15535 (N_15535,N_13636,N_14150);
and U15536 (N_15536,N_12717,N_13973);
or U15537 (N_15537,N_13747,N_14859);
and U15538 (N_15538,N_13875,N_12948);
nor U15539 (N_15539,N_13053,N_13338);
xnor U15540 (N_15540,N_14007,N_14139);
nand U15541 (N_15541,N_12629,N_14908);
or U15542 (N_15542,N_14992,N_12934);
or U15543 (N_15543,N_12580,N_13531);
or U15544 (N_15544,N_13361,N_12792);
or U15545 (N_15545,N_14334,N_14917);
nor U15546 (N_15546,N_12924,N_14590);
nand U15547 (N_15547,N_12768,N_14096);
or U15548 (N_15548,N_13272,N_13975);
nor U15549 (N_15549,N_12514,N_12636);
nand U15550 (N_15550,N_12688,N_14298);
xnor U15551 (N_15551,N_14213,N_13328);
xnor U15552 (N_15552,N_13895,N_14815);
or U15553 (N_15553,N_13752,N_14777);
or U15554 (N_15554,N_14576,N_14160);
nor U15555 (N_15555,N_12577,N_14780);
xor U15556 (N_15556,N_12587,N_14902);
xnor U15557 (N_15557,N_12616,N_13265);
or U15558 (N_15558,N_13023,N_13229);
nand U15559 (N_15559,N_14036,N_14879);
nor U15560 (N_15560,N_13674,N_14700);
nor U15561 (N_15561,N_14152,N_13290);
xnor U15562 (N_15562,N_14074,N_13656);
nand U15563 (N_15563,N_14554,N_12566);
xnor U15564 (N_15564,N_13526,N_14746);
nor U15565 (N_15565,N_14799,N_14229);
xnor U15566 (N_15566,N_12940,N_13767);
nor U15567 (N_15567,N_12802,N_12932);
and U15568 (N_15568,N_13478,N_13165);
and U15569 (N_15569,N_14434,N_12647);
and U15570 (N_15570,N_12683,N_12596);
nor U15571 (N_15571,N_14305,N_14190);
xor U15572 (N_15572,N_14570,N_13662);
xor U15573 (N_15573,N_12764,N_13129);
nor U15574 (N_15574,N_13995,N_14303);
and U15575 (N_15575,N_14448,N_14803);
xor U15576 (N_15576,N_14319,N_14136);
and U15577 (N_15577,N_13257,N_12766);
nor U15578 (N_15578,N_14872,N_14442);
xnor U15579 (N_15579,N_14126,N_13188);
nand U15580 (N_15580,N_13899,N_14519);
or U15581 (N_15581,N_13373,N_14810);
nor U15582 (N_15582,N_13921,N_12907);
xnor U15583 (N_15583,N_13605,N_13139);
or U15584 (N_15584,N_13834,N_14580);
nor U15585 (N_15585,N_12887,N_12807);
nor U15586 (N_15586,N_12809,N_14971);
xnor U15587 (N_15587,N_14495,N_13722);
nand U15588 (N_15588,N_13575,N_14416);
or U15589 (N_15589,N_13359,N_14841);
nor U15590 (N_15590,N_13227,N_12581);
nor U15591 (N_15591,N_14008,N_14215);
xnor U15592 (N_15592,N_12983,N_14538);
or U15593 (N_15593,N_12733,N_13222);
and U15594 (N_15594,N_13925,N_13278);
or U15595 (N_15595,N_13819,N_14364);
and U15596 (N_15596,N_14157,N_12502);
nand U15597 (N_15597,N_12854,N_14726);
or U15598 (N_15598,N_14481,N_14682);
nand U15599 (N_15599,N_14962,N_14637);
xnor U15600 (N_15600,N_14571,N_14774);
xnor U15601 (N_15601,N_14556,N_12960);
nand U15602 (N_15602,N_13716,N_13389);
or U15603 (N_15603,N_13353,N_13904);
or U15604 (N_15604,N_12825,N_14669);
and U15605 (N_15605,N_12590,N_13332);
xor U15606 (N_15606,N_14292,N_13402);
and U15607 (N_15607,N_13552,N_12500);
nand U15608 (N_15608,N_14717,N_14920);
nand U15609 (N_15609,N_14439,N_12677);
and U15610 (N_15610,N_12976,N_14511);
and U15611 (N_15611,N_12645,N_12853);
xnor U15612 (N_15612,N_14393,N_13734);
and U15613 (N_15613,N_12788,N_14504);
or U15614 (N_15614,N_12503,N_14773);
nor U15615 (N_15615,N_13397,N_13517);
nand U15616 (N_15616,N_14132,N_13553);
and U15617 (N_15617,N_13985,N_13812);
and U15618 (N_15618,N_13404,N_14656);
or U15619 (N_15619,N_14402,N_13915);
and U15620 (N_15620,N_14344,N_13011);
nor U15621 (N_15621,N_14899,N_14752);
nor U15622 (N_15622,N_13339,N_14484);
nor U15623 (N_15623,N_14972,N_14824);
and U15624 (N_15624,N_14256,N_13099);
nand U15625 (N_15625,N_13537,N_13078);
nor U15626 (N_15626,N_13453,N_13760);
and U15627 (N_15627,N_13754,N_12713);
or U15628 (N_15628,N_13063,N_13025);
nand U15629 (N_15629,N_14876,N_13748);
or U15630 (N_15630,N_13084,N_14013);
nand U15631 (N_15631,N_13686,N_12757);
and U15632 (N_15632,N_12523,N_14252);
xor U15633 (N_15633,N_14263,N_12710);
or U15634 (N_15634,N_12965,N_13155);
xnor U15635 (N_15635,N_13854,N_13264);
and U15636 (N_15636,N_14698,N_13194);
nor U15637 (N_15637,N_14473,N_12812);
nand U15638 (N_15638,N_13186,N_14490);
xor U15639 (N_15639,N_13492,N_14619);
nand U15640 (N_15640,N_14660,N_13115);
nor U15641 (N_15641,N_14146,N_12507);
and U15642 (N_15642,N_13488,N_13454);
nand U15643 (N_15643,N_14543,N_13358);
xor U15644 (N_15644,N_13039,N_14850);
and U15645 (N_15645,N_14615,N_13701);
and U15646 (N_15646,N_14339,N_13680);
nand U15647 (N_15647,N_13954,N_13698);
xnor U15648 (N_15648,N_13773,N_12522);
xor U15649 (N_15649,N_14642,N_14004);
xor U15650 (N_15650,N_14955,N_14410);
and U15651 (N_15651,N_14234,N_14205);
or U15652 (N_15652,N_13009,N_14653);
or U15653 (N_15653,N_13598,N_12656);
xor U15654 (N_15654,N_13438,N_13241);
and U15655 (N_15655,N_12783,N_14022);
xnor U15656 (N_15656,N_14651,N_12567);
or U15657 (N_15657,N_13291,N_14530);
nor U15658 (N_15658,N_14041,N_12988);
xnor U15659 (N_15659,N_14930,N_14369);
xnor U15660 (N_15660,N_12691,N_14435);
and U15661 (N_15661,N_14214,N_14924);
xnor U15662 (N_15662,N_12664,N_12559);
and U15663 (N_15663,N_14616,N_14324);
xor U15664 (N_15664,N_13589,N_14754);
or U15665 (N_15665,N_14068,N_13233);
and U15666 (N_15666,N_13235,N_14867);
or U15667 (N_15667,N_13621,N_13166);
and U15668 (N_15668,N_14802,N_13668);
xnor U15669 (N_15669,N_12692,N_12833);
xor U15670 (N_15670,N_12562,N_14890);
xnor U15671 (N_15671,N_13449,N_12791);
or U15672 (N_15672,N_14417,N_13794);
nand U15673 (N_15673,N_12955,N_14875);
and U15674 (N_15674,N_13484,N_14164);
nand U15675 (N_15675,N_13050,N_14299);
or U15676 (N_15676,N_14760,N_14524);
nand U15677 (N_15677,N_14736,N_13677);
nor U15678 (N_15678,N_13141,N_13013);
and U15679 (N_15679,N_13465,N_14155);
nor U15680 (N_15680,N_13696,N_13071);
nand U15681 (N_15681,N_14967,N_13936);
nor U15682 (N_15682,N_13466,N_14788);
or U15683 (N_15683,N_13784,N_13736);
or U15684 (N_15684,N_14552,N_12971);
and U15685 (N_15685,N_14749,N_13654);
and U15686 (N_15686,N_12574,N_14203);
or U15687 (N_15687,N_13948,N_14113);
xnor U15688 (N_15688,N_12832,N_13963);
nand U15689 (N_15689,N_13890,N_14644);
xor U15690 (N_15690,N_14862,N_12579);
nand U15691 (N_15691,N_13003,N_12555);
or U15692 (N_15692,N_14926,N_13037);
nor U15693 (N_15693,N_12973,N_14309);
xnor U15694 (N_15694,N_13765,N_14588);
or U15695 (N_15695,N_14218,N_14635);
nor U15696 (N_15696,N_12741,N_13016);
nand U15697 (N_15697,N_14593,N_13883);
and U15698 (N_15698,N_14861,N_14623);
or U15699 (N_15699,N_13561,N_13386);
nor U15700 (N_15700,N_13214,N_13849);
xor U15701 (N_15701,N_14111,N_14592);
xor U15702 (N_15702,N_13408,N_13924);
or U15703 (N_15703,N_13678,N_12568);
and U15704 (N_15704,N_13474,N_13416);
xor U15705 (N_15705,N_14048,N_14885);
or U15706 (N_15706,N_12761,N_13335);
nor U15707 (N_15707,N_13054,N_13065);
and U15708 (N_15708,N_12619,N_12639);
and U15709 (N_15709,N_13626,N_13193);
and U15710 (N_15710,N_13664,N_14243);
xnor U15711 (N_15711,N_14864,N_12525);
xnor U15712 (N_15712,N_12909,N_13200);
or U15713 (N_15713,N_14259,N_14281);
nand U15714 (N_15714,N_13190,N_12763);
nor U15715 (N_15715,N_13756,N_14706);
or U15716 (N_15716,N_14072,N_13692);
xnor U15717 (N_15717,N_14909,N_13022);
and U15718 (N_15718,N_14024,N_12654);
nand U15719 (N_15719,N_14262,N_12801);
and U15720 (N_15720,N_14359,N_12627);
nor U15721 (N_15721,N_14855,N_12513);
xor U15722 (N_15722,N_13157,N_14317);
xnor U15723 (N_15723,N_14665,N_13271);
xnor U15724 (N_15724,N_12543,N_13979);
or U15725 (N_15725,N_14181,N_12509);
xor U15726 (N_15726,N_12620,N_12831);
and U15727 (N_15727,N_14501,N_13462);
and U15728 (N_15728,N_13818,N_12626);
and U15729 (N_15729,N_14163,N_12673);
nor U15730 (N_15730,N_13280,N_14340);
and U15731 (N_15731,N_14673,N_12606);
nand U15732 (N_15732,N_13086,N_14537);
nand U15733 (N_15733,N_14587,N_14579);
and U15734 (N_15734,N_14723,N_14757);
and U15735 (N_15735,N_13409,N_12658);
or U15736 (N_15736,N_14378,N_14206);
nor U15737 (N_15737,N_14077,N_13612);
nor U15738 (N_15738,N_13586,N_14405);
and U15739 (N_15739,N_13461,N_12767);
or U15740 (N_15740,N_12992,N_14561);
nand U15741 (N_15741,N_14124,N_12859);
and U15742 (N_15742,N_12811,N_14631);
and U15743 (N_15743,N_14129,N_13998);
nor U15744 (N_15744,N_12747,N_14695);
or U15745 (N_15745,N_13004,N_14602);
nand U15746 (N_15746,N_13652,N_13407);
and U15747 (N_15747,N_14228,N_14383);
nand U15748 (N_15748,N_13840,N_14730);
xnor U15749 (N_15749,N_12779,N_12504);
nor U15750 (N_15750,N_12987,N_12613);
nand U15751 (N_15751,N_13931,N_13545);
and U15752 (N_15752,N_13663,N_14376);
xnor U15753 (N_15753,N_12771,N_13123);
or U15754 (N_15754,N_12968,N_14696);
nor U15755 (N_15755,N_13075,N_14731);
nand U15756 (N_15756,N_13655,N_14981);
nor U15757 (N_15757,N_13184,N_14921);
nor U15758 (N_15758,N_13316,N_12896);
nand U15759 (N_15759,N_12712,N_13185);
nor U15760 (N_15760,N_13406,N_14817);
nor U15761 (N_15761,N_13689,N_12605);
or U15762 (N_15762,N_13513,N_13451);
nor U15763 (N_15763,N_13710,N_13095);
and U15764 (N_15764,N_12725,N_13852);
and U15765 (N_15765,N_13393,N_12618);
nor U15766 (N_15766,N_14787,N_14396);
and U15767 (N_15767,N_14989,N_14026);
nand U15768 (N_15768,N_13870,N_12646);
nor U15769 (N_15769,N_14331,N_13467);
xor U15770 (N_15770,N_12730,N_13609);
nand U15771 (N_15771,N_14438,N_13252);
and U15772 (N_15772,N_12752,N_12818);
and U15773 (N_15773,N_13330,N_12847);
xnor U15774 (N_15774,N_14613,N_13401);
xnor U15775 (N_15775,N_14762,N_13305);
nor U15776 (N_15776,N_14374,N_14933);
nor U15777 (N_15777,N_13528,N_12672);
nand U15778 (N_15778,N_13144,N_14306);
or U15779 (N_15779,N_13601,N_13026);
or U15780 (N_15780,N_13962,N_14691);
or U15781 (N_15781,N_12598,N_14693);
nand U15782 (N_15782,N_13150,N_12724);
xor U15783 (N_15783,N_12793,N_14069);
nand U15784 (N_15784,N_14209,N_12794);
xnor U15785 (N_15785,N_13800,N_14710);
nand U15786 (N_15786,N_13994,N_12667);
and U15787 (N_15787,N_14709,N_12610);
nand U15788 (N_15788,N_13106,N_14540);
or U15789 (N_15789,N_13110,N_13774);
xnor U15790 (N_15790,N_13218,N_14102);
nand U15791 (N_15791,N_13839,N_12603);
or U15792 (N_15792,N_13659,N_12893);
or U15793 (N_15793,N_13130,N_13124);
or U15794 (N_15794,N_13237,N_13419);
and U15795 (N_15795,N_14117,N_13405);
or U15796 (N_15796,N_12607,N_14342);
nand U15797 (N_15797,N_12850,N_14308);
xor U15798 (N_15798,N_12743,N_14469);
nor U15799 (N_15799,N_14460,N_14915);
xnor U15800 (N_15800,N_14628,N_14911);
xnor U15801 (N_15801,N_14610,N_12529);
or U15802 (N_15802,N_13838,N_14609);
nor U15803 (N_15803,N_13334,N_14498);
nor U15804 (N_15804,N_13811,N_14168);
xor U15805 (N_15805,N_13532,N_12950);
nor U15806 (N_15806,N_13830,N_12877);
or U15807 (N_15807,N_13314,N_14020);
and U15808 (N_15808,N_13287,N_13390);
or U15809 (N_15809,N_14414,N_14513);
xor U15810 (N_15810,N_14798,N_14018);
nor U15811 (N_15811,N_13953,N_14701);
and U15812 (N_15812,N_14227,N_13653);
nand U15813 (N_15813,N_14503,N_13427);
nand U15814 (N_15814,N_14889,N_14386);
and U15815 (N_15815,N_14037,N_12578);
nand U15816 (N_15816,N_13576,N_12928);
nand U15817 (N_15817,N_13262,N_12820);
or U15818 (N_15818,N_14800,N_14346);
xor U15819 (N_15819,N_12716,N_14172);
and U15820 (N_15820,N_14683,N_14092);
nor U15821 (N_15821,N_13615,N_13464);
nor U15822 (N_15822,N_14395,N_13606);
xnor U15823 (N_15823,N_12883,N_14254);
or U15824 (N_15824,N_14149,N_14600);
xor U15825 (N_15825,N_12520,N_14230);
and U15826 (N_15826,N_13516,N_13219);
or U15827 (N_15827,N_13377,N_14877);
and U15828 (N_15828,N_13584,N_13732);
nand U15829 (N_15829,N_14648,N_14038);
nand U15830 (N_15830,N_13846,N_14852);
xor U15831 (N_15831,N_12744,N_13908);
or U15832 (N_15832,N_14922,N_13592);
nand U15833 (N_15833,N_14779,N_13282);
nor U15834 (N_15834,N_12734,N_14178);
and U15835 (N_15835,N_13782,N_14860);
and U15836 (N_15836,N_13798,N_13999);
nor U15837 (N_15837,N_13105,N_14304);
nor U15838 (N_15838,N_13379,N_13228);
or U15839 (N_15839,N_13072,N_12974);
nor U15840 (N_15840,N_13726,N_12858);
nor U15841 (N_15841,N_12707,N_13932);
xor U15842 (N_15842,N_13476,N_13411);
nand U15843 (N_15843,N_12866,N_13081);
xnor U15844 (N_15844,N_14453,N_14655);
xnor U15845 (N_15845,N_12879,N_13294);
nor U15846 (N_15846,N_12855,N_13267);
nor U15847 (N_15847,N_13483,N_14661);
nor U15848 (N_15848,N_14141,N_13435);
xor U15849 (N_15849,N_12838,N_13730);
and U15850 (N_15850,N_13293,N_13337);
and U15851 (N_15851,N_13691,N_13224);
nor U15852 (N_15852,N_14758,N_13793);
and U15853 (N_15853,N_14286,N_14878);
nand U15854 (N_15854,N_14224,N_14314);
or U15855 (N_15855,N_14954,N_12851);
or U15856 (N_15856,N_13285,N_14465);
nand U15857 (N_15857,N_13494,N_13180);
nor U15858 (N_15858,N_13809,N_14424);
xnor U15859 (N_15859,N_13489,N_13951);
nand U15860 (N_15860,N_12720,N_13893);
nand U15861 (N_15861,N_13820,N_14002);
xnor U15862 (N_15862,N_13223,N_12920);
and U15863 (N_15863,N_14235,N_13093);
nand U15864 (N_15864,N_14508,N_14510);
xnor U15865 (N_15865,N_13096,N_13961);
nand U15866 (N_15866,N_14158,N_12515);
or U15867 (N_15867,N_14952,N_14220);
nor U15868 (N_15868,N_14323,N_14377);
or U15869 (N_15869,N_14257,N_13020);
or U15870 (N_15870,N_13108,N_14913);
xnor U15871 (N_15871,N_14216,N_12695);
nor U15872 (N_15872,N_12655,N_13993);
and U15873 (N_15873,N_13415,N_12803);
xor U15874 (N_15874,N_13244,N_12552);
and U15875 (N_15875,N_13970,N_14721);
nor U15876 (N_15876,N_13324,N_13941);
nor U15877 (N_15877,N_13220,N_12748);
or U15878 (N_15878,N_14033,N_14533);
nor U15879 (N_15879,N_12589,N_14891);
nand U15880 (N_15880,N_12894,N_14063);
and U15881 (N_15881,N_14496,N_12902);
nand U15882 (N_15882,N_12804,N_13885);
nand U15883 (N_15883,N_13859,N_14763);
or U15884 (N_15884,N_14858,N_13587);
nand U15885 (N_15885,N_12621,N_13441);
xnor U15886 (N_15886,N_13248,N_13142);
nand U15887 (N_15887,N_13145,N_13570);
or U15888 (N_15888,N_13042,N_14271);
or U15889 (N_15889,N_12796,N_12750);
and U15890 (N_15890,N_13396,N_13704);
or U15891 (N_15891,N_12685,N_14394);
and U15892 (N_15892,N_13863,N_13413);
or U15893 (N_15893,N_13473,N_12890);
nand U15894 (N_15894,N_14900,N_14599);
nor U15895 (N_15895,N_13940,N_12958);
nor U15896 (N_15896,N_13596,N_13595);
or U15897 (N_15897,N_14279,N_14918);
and U15898 (N_15898,N_12604,N_14003);
nand U15899 (N_15899,N_14520,N_14663);
nand U15900 (N_15900,N_14193,N_13588);
nand U15901 (N_15901,N_12519,N_14056);
nand U15902 (N_15902,N_12908,N_14935);
or U15903 (N_15903,N_13862,N_14786);
nor U15904 (N_15904,N_13051,N_14813);
or U15905 (N_15905,N_12918,N_14318);
xnor U15906 (N_15906,N_13327,N_13700);
nor U15907 (N_15907,N_13079,N_12703);
xor U15908 (N_15908,N_14659,N_14459);
xor U15909 (N_15909,N_12835,N_14409);
and U15910 (N_15910,N_13230,N_14745);
and U15911 (N_15911,N_14090,N_14938);
xor U15912 (N_15912,N_12749,N_13549);
and U15913 (N_15913,N_14795,N_14509);
xor U15914 (N_15914,N_14109,N_13618);
nor U15915 (N_15915,N_14425,N_13873);
nor U15916 (N_15916,N_14012,N_13992);
xor U15917 (N_15917,N_13675,N_13699);
nand U15918 (N_15918,N_14040,N_12600);
or U15919 (N_15919,N_13897,N_14892);
nand U15920 (N_15920,N_14910,N_12540);
or U15921 (N_15921,N_13591,N_12910);
or U15922 (N_15922,N_14358,N_13565);
and U15923 (N_15923,N_14010,N_13122);
xnor U15924 (N_15924,N_13810,N_13169);
nand U15925 (N_15925,N_12624,N_14057);
or U15926 (N_15926,N_13559,N_13236);
nand U15927 (N_15927,N_12678,N_14830);
xnor U15928 (N_15928,N_12995,N_14768);
nand U15929 (N_15929,N_12982,N_14748);
nand U15930 (N_15930,N_14611,N_14703);
or U15931 (N_15931,N_13311,N_13148);
nand U15932 (N_15932,N_14708,N_14153);
or U15933 (N_15933,N_14814,N_13544);
nor U15934 (N_15934,N_14846,N_14998);
nor U15935 (N_15935,N_12937,N_14238);
and U15936 (N_15936,N_13117,N_14617);
or U15937 (N_15937,N_13801,N_12884);
xnor U15938 (N_15938,N_14122,N_13783);
or U15939 (N_15939,N_13844,N_13593);
nand U15940 (N_15940,N_13771,N_13949);
nand U15941 (N_15941,N_13456,N_14711);
or U15942 (N_15942,N_12824,N_14273);
and U15943 (N_15943,N_12941,N_14195);
xor U15944 (N_15944,N_13440,N_12891);
nor U15945 (N_15945,N_13501,N_12785);
and U15946 (N_15946,N_12659,N_14247);
or U15947 (N_15947,N_13719,N_13927);
and U15948 (N_15948,N_13690,N_12914);
and U15949 (N_15949,N_13444,N_14999);
nand U15950 (N_15950,N_14783,N_13170);
nor U15951 (N_15951,N_14837,N_13345);
and U15952 (N_15952,N_13363,N_12963);
nor U15953 (N_15953,N_14067,N_13943);
and U15954 (N_15954,N_14983,N_14315);
and U15955 (N_15955,N_13751,N_12573);
and U15956 (N_15956,N_12797,N_13273);
xor U15957 (N_15957,N_13035,N_14145);
nor U15958 (N_15958,N_14427,N_13974);
or U15959 (N_15959,N_14388,N_14199);
nand U15960 (N_15960,N_12557,N_12905);
and U15961 (N_15961,N_13909,N_13430);
nand U15962 (N_15962,N_13515,N_14494);
nand U15963 (N_15963,N_14343,N_14363);
and U15964 (N_15964,N_12780,N_14545);
nor U15965 (N_15965,N_14985,N_13720);
and U15966 (N_15966,N_13032,N_13628);
and U15967 (N_15967,N_13535,N_13418);
xnor U15968 (N_15968,N_14626,N_13367);
nor U15969 (N_15969,N_14322,N_13976);
or U15970 (N_15970,N_14107,N_14294);
nand U15971 (N_15971,N_13622,N_14638);
nor U15972 (N_15972,N_13250,N_14165);
nor U15973 (N_15973,N_14023,N_12593);
nor U15974 (N_15974,N_13143,N_13371);
or U15975 (N_15975,N_13920,N_14351);
or U15976 (N_15976,N_14776,N_12889);
nand U15977 (N_15977,N_14135,N_14131);
nand U15978 (N_15978,N_13926,N_13509);
xor U15979 (N_15979,N_14170,N_14025);
nand U15980 (N_15980,N_12869,N_13459);
nor U15981 (N_15981,N_13579,N_13487);
xor U15982 (N_15982,N_13433,N_13670);
nand U15983 (N_15983,N_12689,N_12671);
nand U15984 (N_15984,N_14529,N_14027);
or U15985 (N_15985,N_13669,N_14173);
nand U15986 (N_15986,N_14251,N_14019);
xnor U15987 (N_15987,N_14226,N_12997);
or U15988 (N_15988,N_12738,N_12530);
or U15989 (N_15989,N_14329,N_14156);
and U15990 (N_15990,N_14751,N_14360);
or U15991 (N_15991,N_13558,N_14812);
and U15992 (N_15992,N_13052,N_12564);
xor U15993 (N_15993,N_14772,N_13745);
and U15994 (N_15994,N_13912,N_14032);
nand U15995 (N_15995,N_13113,N_12537);
xnor U15996 (N_15996,N_14976,N_13457);
nand U15997 (N_15997,N_14468,N_14466);
or U15998 (N_15998,N_12994,N_14105);
or U15999 (N_15999,N_13805,N_12538);
and U16000 (N_16000,N_13268,N_12545);
xor U16001 (N_16001,N_13758,N_14555);
nand U16002 (N_16002,N_13725,N_14372);
and U16003 (N_16003,N_13608,N_14604);
or U16004 (N_16004,N_12800,N_13957);
nor U16005 (N_16005,N_12933,N_13702);
xnor U16006 (N_16006,N_12669,N_14606);
and U16007 (N_16007,N_14894,N_13911);
nand U16008 (N_16008,N_13333,N_12719);
or U16009 (N_16009,N_14147,N_14426);
or U16010 (N_16010,N_12561,N_12979);
nor U16011 (N_16011,N_14791,N_14307);
or U16012 (N_16012,N_14990,N_13092);
xor U16013 (N_16013,N_13292,N_14801);
and U16014 (N_16014,N_14681,N_13610);
or U16015 (N_16015,N_14167,N_13731);
and U16016 (N_16016,N_13650,N_12558);
xor U16017 (N_16017,N_14064,N_13376);
xnor U16018 (N_16018,N_13744,N_13111);
xor U16019 (N_16019,N_13112,N_14678);
and U16020 (N_16020,N_13882,N_13518);
and U16021 (N_16021,N_14300,N_14563);
xor U16022 (N_16022,N_14680,N_14705);
nor U16023 (N_16023,N_14231,N_13384);
or U16024 (N_16024,N_13813,N_14550);
xnor U16025 (N_16025,N_14392,N_13303);
and U16026 (N_16026,N_14627,N_12985);
xor U16027 (N_16027,N_13069,N_13232);
nand U16028 (N_16028,N_14029,N_14350);
and U16029 (N_16029,N_14874,N_13779);
or U16030 (N_16030,N_13134,N_13426);
xor U16031 (N_16031,N_12661,N_14668);
and U16032 (N_16032,N_14666,N_14148);
nand U16033 (N_16033,N_13497,N_13536);
or U16034 (N_16034,N_14045,N_14697);
or U16035 (N_16035,N_14050,N_12926);
or U16036 (N_16036,N_14614,N_13757);
or U16037 (N_16037,N_12897,N_14478);
and U16038 (N_16038,N_13802,N_14781);
or U16039 (N_16039,N_12505,N_13152);
nand U16040 (N_16040,N_12939,N_14221);
nand U16041 (N_16041,N_12518,N_13900);
nor U16042 (N_16042,N_13382,N_14759);
or U16043 (N_16043,N_14839,N_13164);
xnor U16044 (N_16044,N_14906,N_13857);
xor U16045 (N_16045,N_14290,N_13896);
nor U16046 (N_16046,N_14093,N_13822);
nand U16047 (N_16047,N_14116,N_14945);
nor U16048 (N_16048,N_12839,N_14982);
xor U16049 (N_16049,N_13693,N_12898);
and U16050 (N_16050,N_14629,N_14212);
and U16051 (N_16051,N_12705,N_14451);
nor U16052 (N_16052,N_13872,N_13279);
nand U16053 (N_16053,N_13412,N_14071);
xnor U16054 (N_16054,N_14667,N_13703);
or U16055 (N_16055,N_12742,N_13832);
xor U16056 (N_16056,N_13211,N_14189);
xnor U16057 (N_16057,N_13158,N_12806);
xor U16058 (N_16058,N_13173,N_14969);
xnor U16059 (N_16059,N_13538,N_13855);
nor U16060 (N_16060,N_13781,N_13395);
or U16061 (N_16061,N_14437,N_14128);
nor U16062 (N_16062,N_13040,N_14059);
nor U16063 (N_16063,N_13083,N_12663);
or U16064 (N_16064,N_12929,N_14712);
nand U16065 (N_16065,N_14657,N_12591);
and U16066 (N_16066,N_13577,N_13385);
nor U16067 (N_16067,N_13938,N_13329);
xor U16068 (N_16068,N_13159,N_14255);
and U16069 (N_16069,N_14505,N_13879);
nor U16070 (N_16070,N_14973,N_12864);
and U16071 (N_16071,N_13383,N_14684);
nand U16072 (N_16072,N_14436,N_13047);
and U16073 (N_16073,N_14951,N_14361);
nand U16074 (N_16074,N_13076,N_12699);
and U16075 (N_16075,N_14811,N_13583);
xor U16076 (N_16076,N_14120,N_13174);
nand U16077 (N_16077,N_14062,N_14455);
and U16078 (N_16078,N_14893,N_13906);
nor U16079 (N_16079,N_14694,N_13597);
xnor U16080 (N_16080,N_14958,N_13136);
and U16081 (N_16081,N_14901,N_13073);
and U16082 (N_16082,N_14031,N_14095);
and U16083 (N_16083,N_13312,N_14159);
nand U16084 (N_16084,N_14866,N_13505);
nor U16085 (N_16085,N_14769,N_13203);
and U16086 (N_16086,N_14054,N_14191);
nor U16087 (N_16087,N_12662,N_14370);
and U16088 (N_16088,N_13348,N_13034);
nor U16089 (N_16089,N_12922,N_12848);
or U16090 (N_16090,N_14362,N_13347);
nor U16091 (N_16091,N_14934,N_14447);
nand U16092 (N_16092,N_12916,N_13212);
or U16093 (N_16093,N_13172,N_12773);
xor U16094 (N_16094,N_14625,N_13711);
or U16095 (N_16095,N_13192,N_14103);
nand U16096 (N_16096,N_14916,N_14912);
nand U16097 (N_16097,N_14264,N_12980);
nand U16098 (N_16098,N_14687,N_12512);
or U16099 (N_16099,N_14365,N_13639);
and U16100 (N_16100,N_13568,N_13888);
nand U16101 (N_16101,N_13350,N_13959);
nor U16102 (N_16102,N_14088,N_13146);
nand U16103 (N_16103,N_13182,N_13514);
or U16104 (N_16104,N_13231,N_13635);
nand U16105 (N_16105,N_13191,N_14265);
or U16106 (N_16106,N_12834,N_12953);
xnor U16107 (N_16107,N_14328,N_12945);
or U16108 (N_16108,N_14237,N_14832);
or U16109 (N_16109,N_14497,N_14907);
and U16110 (N_16110,N_13286,N_14326);
xnor U16111 (N_16111,N_14562,N_13867);
or U16112 (N_16112,N_13894,N_13101);
and U16113 (N_16113,N_13177,N_13398);
xnor U16114 (N_16114,N_12722,N_13546);
nand U16115 (N_16115,N_14670,N_14636);
or U16116 (N_16116,N_14198,N_13364);
nor U16117 (N_16117,N_12542,N_13831);
xnor U16118 (N_16118,N_13298,N_12614);
nor U16119 (N_16119,N_13472,N_12701);
or U16120 (N_16120,N_13764,N_13482);
or U16121 (N_16121,N_13242,N_12737);
nor U16122 (N_16122,N_13151,N_12882);
nand U16123 (N_16123,N_14142,N_14295);
xor U16124 (N_16124,N_13195,N_12993);
nor U16125 (N_16125,N_13163,N_13929);
or U16126 (N_16126,N_13739,N_14112);
and U16127 (N_16127,N_12873,N_14233);
nor U16128 (N_16128,N_13629,N_14747);
xor U16129 (N_16129,N_13343,N_12817);
nor U16130 (N_16130,N_14187,N_14463);
nand U16131 (N_16131,N_14452,N_12870);
or U16132 (N_16132,N_14192,N_13387);
nand U16133 (N_16133,N_13485,N_13543);
or U16134 (N_16134,N_12648,N_13447);
or U16135 (N_16135,N_13132,N_14446);
nor U16136 (N_16136,N_13342,N_14838);
nand U16137 (N_16137,N_14662,N_14084);
xnor U16138 (N_16138,N_14166,N_13491);
nor U16139 (N_16139,N_13780,N_13031);
or U16140 (N_16140,N_13198,N_12746);
and U16141 (N_16141,N_13965,N_13694);
nand U16142 (N_16142,N_13729,N_13967);
nand U16143 (N_16143,N_12857,N_12628);
xor U16144 (N_16144,N_13661,N_14108);
and U16145 (N_16145,N_13935,N_14087);
nor U16146 (N_16146,N_14476,N_13120);
and U16147 (N_16147,N_13277,N_14790);
xor U16148 (N_16148,N_13898,N_14949);
or U16149 (N_16149,N_12572,N_12778);
or U16150 (N_16150,N_14015,N_14586);
or U16151 (N_16151,N_14756,N_13463);
xnor U16152 (N_16152,N_14753,N_13560);
nand U16153 (N_16153,N_14250,N_13283);
nand U16154 (N_16154,N_13498,N_13825);
or U16155 (N_16155,N_12637,N_12912);
nand U16156 (N_16156,N_14154,N_12535);
or U16157 (N_16157,N_14161,N_13477);
xor U16158 (N_16158,N_13199,N_13439);
xor U16159 (N_16159,N_12975,N_13910);
or U16160 (N_16160,N_12711,N_13607);
and U16161 (N_16161,N_13743,N_14065);
and U16162 (N_16162,N_14244,N_14979);
or U16163 (N_16163,N_14544,N_14833);
xor U16164 (N_16164,N_14947,N_14689);
xnor U16165 (N_16165,N_13496,N_12693);
or U16166 (N_16166,N_13637,N_13835);
nand U16167 (N_16167,N_13027,N_14507);
and U16168 (N_16168,N_12892,N_14929);
nand U16169 (N_16169,N_12862,N_13737);
or U16170 (N_16170,N_13202,N_13788);
or U16171 (N_16171,N_14276,N_14483);
nand U16172 (N_16172,N_13114,N_14454);
nor U16173 (N_16173,N_14819,N_14099);
nor U16174 (N_16174,N_14249,N_13270);
nand U16175 (N_16175,N_12586,N_13529);
and U16176 (N_16176,N_14725,N_14009);
and U16177 (N_16177,N_13865,N_13958);
and U16178 (N_16178,N_14188,N_13886);
nor U16179 (N_16179,N_14397,N_14489);
nand U16180 (N_16180,N_12714,N_14449);
and U16181 (N_16181,N_14512,N_14335);
and U16182 (N_16182,N_14699,N_12584);
nand U16183 (N_16183,N_13829,N_12698);
and U16184 (N_16184,N_14011,N_13480);
and U16185 (N_16185,N_13786,N_13126);
xor U16186 (N_16186,N_12947,N_14186);
nand U16187 (N_16187,N_14541,N_12702);
nand U16188 (N_16188,N_13631,N_14950);
or U16189 (N_16189,N_14061,N_12740);
nand U16190 (N_16190,N_13239,N_14515);
and U16191 (N_16191,N_13300,N_14646);
or U16192 (N_16192,N_12592,N_13869);
nand U16193 (N_16193,N_13125,N_13688);
and U16194 (N_16194,N_13687,N_14462);
or U16195 (N_16195,N_13116,N_13468);
nor U16196 (N_16196,N_13555,N_13619);
nor U16197 (N_16197,N_12666,N_13196);
nand U16198 (N_16198,N_14482,N_14415);
nand U16199 (N_16199,N_12931,N_13255);
nand U16200 (N_16200,N_13068,N_14574);
nand U16201 (N_16201,N_14070,N_12617);
xor U16202 (N_16202,N_12996,N_13749);
xnor U16203 (N_16203,N_13033,N_14943);
or U16204 (N_16204,N_14443,N_14312);
xnor U16205 (N_16205,N_14557,N_13137);
or U16206 (N_16206,N_13728,N_14987);
nor U16207 (N_16207,N_14241,N_12753);
xnor U16208 (N_16208,N_14844,N_12798);
xor U16209 (N_16209,N_14559,N_12571);
nand U16210 (N_16210,N_14937,N_14297);
xnor U16211 (N_16211,N_12736,N_13683);
nor U16212 (N_16212,N_12969,N_14991);
xor U16213 (N_16213,N_12718,N_12632);
and U16214 (N_16214,N_14349,N_14944);
or U16215 (N_16215,N_12759,N_13175);
nor U16216 (N_16216,N_13422,N_12715);
xor U16217 (N_16217,N_13550,N_14432);
or U16218 (N_16218,N_12762,N_13667);
nor U16219 (N_16219,N_14564,N_14006);
nand U16220 (N_16220,N_13613,N_14458);
and U16221 (N_16221,N_14176,N_12644);
nand U16222 (N_16222,N_14808,N_13355);
nand U16223 (N_16223,N_12615,N_13309);
and U16224 (N_16224,N_14897,N_14500);
xor U16225 (N_16225,N_13986,N_13676);
nor U16226 (N_16226,N_14903,N_13666);
and U16227 (N_16227,N_14674,N_14381);
nand U16228 (N_16228,N_13410,N_13648);
or U16229 (N_16229,N_13064,N_14940);
or U16230 (N_16230,N_14021,N_12846);
nand U16231 (N_16231,N_14664,N_13507);
or U16232 (N_16232,N_12684,N_13884);
nand U16233 (N_16233,N_14182,N_14412);
nor U16234 (N_16234,N_12840,N_14133);
nor U16235 (N_16235,N_14114,N_13452);
and U16236 (N_16236,N_14028,N_14474);
nand U16237 (N_16237,N_13864,N_13399);
xnor U16238 (N_16238,N_12999,N_14914);
nand U16239 (N_16239,N_12638,N_13660);
nand U16240 (N_16240,N_14110,N_12967);
or U16241 (N_16241,N_13947,N_13847);
nor U16242 (N_16242,N_13627,N_12925);
nor U16243 (N_16243,N_12972,N_12528);
nor U16244 (N_16244,N_14888,N_14285);
xnor U16245 (N_16245,N_14058,N_13564);
or U16246 (N_16246,N_14583,N_13797);
or U16247 (N_16247,N_12508,N_12652);
xor U16248 (N_16248,N_14995,N_12575);
nor U16249 (N_16249,N_12875,N_12861);
xor U16250 (N_16250,N_13071,N_14489);
and U16251 (N_16251,N_13907,N_14493);
or U16252 (N_16252,N_14748,N_14498);
or U16253 (N_16253,N_14181,N_13968);
nand U16254 (N_16254,N_14908,N_13923);
xnor U16255 (N_16255,N_13719,N_14547);
nand U16256 (N_16256,N_13332,N_12511);
nand U16257 (N_16257,N_14325,N_13756);
nand U16258 (N_16258,N_13023,N_13953);
or U16259 (N_16259,N_13447,N_13476);
xnor U16260 (N_16260,N_13780,N_13018);
nand U16261 (N_16261,N_13393,N_14292);
xnor U16262 (N_16262,N_13488,N_13558);
and U16263 (N_16263,N_14687,N_12664);
nand U16264 (N_16264,N_14680,N_13406);
nand U16265 (N_16265,N_12915,N_12539);
and U16266 (N_16266,N_13697,N_14461);
nand U16267 (N_16267,N_13116,N_13532);
nor U16268 (N_16268,N_14375,N_14177);
xnor U16269 (N_16269,N_13657,N_13977);
nand U16270 (N_16270,N_12861,N_13954);
nand U16271 (N_16271,N_12673,N_13757);
and U16272 (N_16272,N_13901,N_14035);
or U16273 (N_16273,N_14618,N_12522);
or U16274 (N_16274,N_12848,N_13577);
xnor U16275 (N_16275,N_14237,N_13968);
nor U16276 (N_16276,N_14894,N_13364);
xor U16277 (N_16277,N_13585,N_14963);
nor U16278 (N_16278,N_14252,N_14009);
and U16279 (N_16279,N_12520,N_12657);
nor U16280 (N_16280,N_14192,N_14340);
xnor U16281 (N_16281,N_14956,N_14822);
nor U16282 (N_16282,N_12950,N_14343);
and U16283 (N_16283,N_14814,N_13648);
nor U16284 (N_16284,N_13503,N_14247);
nor U16285 (N_16285,N_13145,N_12554);
or U16286 (N_16286,N_14848,N_14405);
nor U16287 (N_16287,N_12555,N_14034);
and U16288 (N_16288,N_13396,N_14739);
and U16289 (N_16289,N_13265,N_12965);
or U16290 (N_16290,N_14519,N_12943);
nor U16291 (N_16291,N_14424,N_13409);
nor U16292 (N_16292,N_14045,N_12986);
xor U16293 (N_16293,N_13847,N_14392);
xor U16294 (N_16294,N_14550,N_14574);
nand U16295 (N_16295,N_13947,N_13655);
nand U16296 (N_16296,N_12896,N_14494);
nand U16297 (N_16297,N_14863,N_14677);
or U16298 (N_16298,N_13693,N_14454);
xor U16299 (N_16299,N_12567,N_13718);
or U16300 (N_16300,N_14296,N_13376);
or U16301 (N_16301,N_12843,N_13340);
xnor U16302 (N_16302,N_14244,N_13332);
nand U16303 (N_16303,N_14563,N_14617);
and U16304 (N_16304,N_13567,N_13260);
xnor U16305 (N_16305,N_12831,N_14280);
nand U16306 (N_16306,N_13238,N_14415);
nand U16307 (N_16307,N_13833,N_13539);
or U16308 (N_16308,N_12855,N_14819);
nand U16309 (N_16309,N_14091,N_13087);
and U16310 (N_16310,N_13593,N_14778);
nor U16311 (N_16311,N_14681,N_13698);
nand U16312 (N_16312,N_14542,N_14930);
and U16313 (N_16313,N_13357,N_14284);
nor U16314 (N_16314,N_13675,N_14679);
and U16315 (N_16315,N_14842,N_14746);
nor U16316 (N_16316,N_12800,N_13189);
nor U16317 (N_16317,N_13331,N_13028);
and U16318 (N_16318,N_13671,N_14166);
or U16319 (N_16319,N_14906,N_13136);
or U16320 (N_16320,N_14202,N_14852);
xnor U16321 (N_16321,N_13478,N_12774);
nor U16322 (N_16322,N_12728,N_14499);
nand U16323 (N_16323,N_13035,N_14996);
and U16324 (N_16324,N_14786,N_12721);
and U16325 (N_16325,N_14105,N_12851);
nor U16326 (N_16326,N_14001,N_14393);
and U16327 (N_16327,N_14423,N_13355);
xor U16328 (N_16328,N_13276,N_13178);
nand U16329 (N_16329,N_14925,N_13626);
nand U16330 (N_16330,N_14416,N_14462);
xor U16331 (N_16331,N_12824,N_13335);
xor U16332 (N_16332,N_14163,N_14934);
xnor U16333 (N_16333,N_14008,N_13032);
xor U16334 (N_16334,N_14536,N_14929);
or U16335 (N_16335,N_13211,N_12948);
nand U16336 (N_16336,N_12592,N_14776);
nand U16337 (N_16337,N_13913,N_13725);
nand U16338 (N_16338,N_14510,N_13912);
or U16339 (N_16339,N_13467,N_13919);
xor U16340 (N_16340,N_14228,N_12985);
and U16341 (N_16341,N_14046,N_13088);
xnor U16342 (N_16342,N_14716,N_12516);
xor U16343 (N_16343,N_14800,N_13360);
and U16344 (N_16344,N_13214,N_14812);
or U16345 (N_16345,N_14035,N_14195);
nand U16346 (N_16346,N_12957,N_13619);
nor U16347 (N_16347,N_13275,N_12509);
nor U16348 (N_16348,N_13854,N_13131);
nand U16349 (N_16349,N_13666,N_13772);
and U16350 (N_16350,N_13172,N_14195);
and U16351 (N_16351,N_13348,N_13836);
or U16352 (N_16352,N_12883,N_14992);
and U16353 (N_16353,N_12527,N_12600);
and U16354 (N_16354,N_14839,N_13992);
nand U16355 (N_16355,N_14040,N_14649);
nor U16356 (N_16356,N_14812,N_12571);
xor U16357 (N_16357,N_13555,N_12623);
xor U16358 (N_16358,N_12571,N_12747);
nor U16359 (N_16359,N_14804,N_13587);
nor U16360 (N_16360,N_14294,N_14543);
xnor U16361 (N_16361,N_12814,N_12823);
and U16362 (N_16362,N_13952,N_13547);
or U16363 (N_16363,N_13982,N_12563);
xnor U16364 (N_16364,N_13869,N_12767);
and U16365 (N_16365,N_12863,N_14895);
nand U16366 (N_16366,N_14736,N_13614);
nor U16367 (N_16367,N_13998,N_14290);
or U16368 (N_16368,N_12696,N_14830);
or U16369 (N_16369,N_12591,N_13541);
and U16370 (N_16370,N_13018,N_13822);
or U16371 (N_16371,N_14587,N_14113);
nor U16372 (N_16372,N_14497,N_14814);
xnor U16373 (N_16373,N_12973,N_14026);
nand U16374 (N_16374,N_14362,N_14799);
xnor U16375 (N_16375,N_13558,N_13546);
xor U16376 (N_16376,N_12553,N_14274);
nor U16377 (N_16377,N_12894,N_14270);
nor U16378 (N_16378,N_12567,N_13995);
nand U16379 (N_16379,N_14846,N_13871);
xor U16380 (N_16380,N_14563,N_14421);
and U16381 (N_16381,N_13941,N_14048);
nand U16382 (N_16382,N_14187,N_14589);
and U16383 (N_16383,N_12723,N_12847);
or U16384 (N_16384,N_14830,N_14413);
nand U16385 (N_16385,N_12872,N_12969);
xor U16386 (N_16386,N_13578,N_14746);
or U16387 (N_16387,N_14345,N_13631);
or U16388 (N_16388,N_14721,N_14199);
xor U16389 (N_16389,N_14823,N_12678);
nand U16390 (N_16390,N_12590,N_13367);
or U16391 (N_16391,N_14189,N_12916);
nand U16392 (N_16392,N_12543,N_12848);
and U16393 (N_16393,N_13300,N_13666);
nand U16394 (N_16394,N_12520,N_14948);
and U16395 (N_16395,N_14987,N_13294);
nor U16396 (N_16396,N_13543,N_13628);
nand U16397 (N_16397,N_14255,N_14083);
nand U16398 (N_16398,N_14438,N_12600);
nand U16399 (N_16399,N_14487,N_14515);
xnor U16400 (N_16400,N_14340,N_14876);
nand U16401 (N_16401,N_13921,N_13414);
nor U16402 (N_16402,N_14226,N_14416);
or U16403 (N_16403,N_12717,N_14326);
nor U16404 (N_16404,N_14169,N_12695);
nor U16405 (N_16405,N_14775,N_13169);
or U16406 (N_16406,N_14582,N_13209);
nand U16407 (N_16407,N_13553,N_13187);
and U16408 (N_16408,N_13775,N_13120);
nor U16409 (N_16409,N_13835,N_12798);
xnor U16410 (N_16410,N_14389,N_12736);
xnor U16411 (N_16411,N_14125,N_13268);
or U16412 (N_16412,N_13810,N_13045);
and U16413 (N_16413,N_14529,N_13781);
or U16414 (N_16414,N_13264,N_14372);
and U16415 (N_16415,N_14473,N_13197);
and U16416 (N_16416,N_14898,N_12547);
and U16417 (N_16417,N_13939,N_12686);
and U16418 (N_16418,N_14909,N_12887);
xnor U16419 (N_16419,N_13816,N_14689);
and U16420 (N_16420,N_14775,N_12920);
nand U16421 (N_16421,N_14040,N_13090);
and U16422 (N_16422,N_12747,N_14453);
nor U16423 (N_16423,N_12823,N_13465);
and U16424 (N_16424,N_13775,N_13534);
xnor U16425 (N_16425,N_14635,N_13427);
and U16426 (N_16426,N_13817,N_14492);
xnor U16427 (N_16427,N_13241,N_13767);
nand U16428 (N_16428,N_14056,N_13216);
nor U16429 (N_16429,N_14455,N_12656);
nor U16430 (N_16430,N_13553,N_12512);
nand U16431 (N_16431,N_13466,N_13979);
nor U16432 (N_16432,N_14857,N_14638);
and U16433 (N_16433,N_13191,N_14924);
and U16434 (N_16434,N_14577,N_14122);
and U16435 (N_16435,N_14190,N_13555);
xnor U16436 (N_16436,N_14324,N_13243);
or U16437 (N_16437,N_14588,N_13656);
nand U16438 (N_16438,N_13883,N_14401);
xor U16439 (N_16439,N_14314,N_14541);
or U16440 (N_16440,N_13325,N_14367);
xor U16441 (N_16441,N_14790,N_12501);
xnor U16442 (N_16442,N_12912,N_13503);
xor U16443 (N_16443,N_14005,N_14670);
nor U16444 (N_16444,N_14638,N_13928);
nand U16445 (N_16445,N_13591,N_13046);
and U16446 (N_16446,N_13260,N_14124);
nor U16447 (N_16447,N_14239,N_14106);
nor U16448 (N_16448,N_12522,N_13013);
nand U16449 (N_16449,N_12887,N_12754);
or U16450 (N_16450,N_13362,N_13975);
and U16451 (N_16451,N_12999,N_13984);
nand U16452 (N_16452,N_14890,N_13664);
xor U16453 (N_16453,N_14947,N_14172);
nor U16454 (N_16454,N_13626,N_12638);
nand U16455 (N_16455,N_13337,N_12790);
xnor U16456 (N_16456,N_13247,N_13281);
nand U16457 (N_16457,N_13487,N_13635);
nor U16458 (N_16458,N_13422,N_14936);
xnor U16459 (N_16459,N_13340,N_13025);
or U16460 (N_16460,N_13664,N_13023);
xnor U16461 (N_16461,N_14549,N_13843);
xnor U16462 (N_16462,N_14515,N_14882);
and U16463 (N_16463,N_12886,N_13580);
and U16464 (N_16464,N_14879,N_14520);
nand U16465 (N_16465,N_13438,N_13534);
xnor U16466 (N_16466,N_14907,N_13540);
and U16467 (N_16467,N_13075,N_14503);
xnor U16468 (N_16468,N_13641,N_14070);
and U16469 (N_16469,N_14297,N_13744);
xor U16470 (N_16470,N_13813,N_14847);
xor U16471 (N_16471,N_13441,N_12944);
and U16472 (N_16472,N_14170,N_13550);
and U16473 (N_16473,N_13008,N_13815);
nor U16474 (N_16474,N_13422,N_12894);
xnor U16475 (N_16475,N_14455,N_13172);
and U16476 (N_16476,N_13281,N_14543);
or U16477 (N_16477,N_14405,N_13295);
or U16478 (N_16478,N_12622,N_13429);
xnor U16479 (N_16479,N_14214,N_13940);
nor U16480 (N_16480,N_13009,N_12658);
and U16481 (N_16481,N_13243,N_14173);
nor U16482 (N_16482,N_14712,N_13787);
nor U16483 (N_16483,N_13291,N_14635);
xor U16484 (N_16484,N_13637,N_14012);
and U16485 (N_16485,N_12598,N_13638);
xnor U16486 (N_16486,N_12894,N_14244);
nand U16487 (N_16487,N_14145,N_13192);
and U16488 (N_16488,N_14051,N_13651);
xnor U16489 (N_16489,N_12917,N_14778);
nand U16490 (N_16490,N_13819,N_14512);
nand U16491 (N_16491,N_12719,N_14202);
or U16492 (N_16492,N_14053,N_13249);
xor U16493 (N_16493,N_13787,N_13223);
nand U16494 (N_16494,N_14817,N_14591);
nand U16495 (N_16495,N_13439,N_13284);
or U16496 (N_16496,N_13660,N_14950);
or U16497 (N_16497,N_14554,N_13031);
nor U16498 (N_16498,N_13189,N_14462);
xnor U16499 (N_16499,N_13675,N_14639);
nand U16500 (N_16500,N_12903,N_14900);
nor U16501 (N_16501,N_13628,N_12707);
nor U16502 (N_16502,N_14869,N_13487);
and U16503 (N_16503,N_12635,N_12707);
xnor U16504 (N_16504,N_13950,N_13120);
and U16505 (N_16505,N_12659,N_14580);
nand U16506 (N_16506,N_13718,N_14953);
nand U16507 (N_16507,N_13240,N_14608);
nor U16508 (N_16508,N_14053,N_13550);
nand U16509 (N_16509,N_13968,N_13985);
nor U16510 (N_16510,N_12502,N_13917);
nand U16511 (N_16511,N_12746,N_12733);
and U16512 (N_16512,N_13552,N_13534);
and U16513 (N_16513,N_13215,N_14848);
and U16514 (N_16514,N_14595,N_13997);
nor U16515 (N_16515,N_14525,N_14216);
and U16516 (N_16516,N_12642,N_14482);
nand U16517 (N_16517,N_14557,N_13902);
nor U16518 (N_16518,N_13772,N_13455);
xor U16519 (N_16519,N_14626,N_13949);
xor U16520 (N_16520,N_14882,N_13655);
xor U16521 (N_16521,N_13967,N_13865);
nand U16522 (N_16522,N_13633,N_14287);
nor U16523 (N_16523,N_13809,N_12769);
xor U16524 (N_16524,N_14854,N_12577);
nand U16525 (N_16525,N_14547,N_14695);
nand U16526 (N_16526,N_12518,N_13583);
and U16527 (N_16527,N_13317,N_13304);
nor U16528 (N_16528,N_13354,N_12538);
and U16529 (N_16529,N_13760,N_14290);
or U16530 (N_16530,N_12515,N_13039);
xor U16531 (N_16531,N_14912,N_13760);
nand U16532 (N_16532,N_13997,N_14015);
nor U16533 (N_16533,N_13693,N_12783);
and U16534 (N_16534,N_13482,N_13740);
or U16535 (N_16535,N_14601,N_13680);
or U16536 (N_16536,N_14475,N_12590);
nand U16537 (N_16537,N_13285,N_13873);
xor U16538 (N_16538,N_13672,N_12968);
nand U16539 (N_16539,N_12993,N_13014);
or U16540 (N_16540,N_14823,N_12552);
xnor U16541 (N_16541,N_14972,N_14962);
xor U16542 (N_16542,N_13343,N_14860);
and U16543 (N_16543,N_13729,N_14813);
nand U16544 (N_16544,N_14071,N_14126);
or U16545 (N_16545,N_14412,N_12887);
xnor U16546 (N_16546,N_12546,N_14714);
nand U16547 (N_16547,N_13507,N_14465);
nor U16548 (N_16548,N_13687,N_13273);
nand U16549 (N_16549,N_13456,N_12880);
nand U16550 (N_16550,N_14361,N_13310);
xor U16551 (N_16551,N_14451,N_13768);
and U16552 (N_16552,N_14675,N_13744);
nor U16553 (N_16553,N_13100,N_13077);
and U16554 (N_16554,N_14626,N_14220);
or U16555 (N_16555,N_12950,N_13705);
nor U16556 (N_16556,N_13473,N_12553);
or U16557 (N_16557,N_14388,N_13079);
and U16558 (N_16558,N_13049,N_12766);
and U16559 (N_16559,N_13574,N_12709);
nor U16560 (N_16560,N_14822,N_13907);
xor U16561 (N_16561,N_13706,N_13084);
and U16562 (N_16562,N_12944,N_14026);
and U16563 (N_16563,N_12952,N_14328);
nor U16564 (N_16564,N_13074,N_12594);
nand U16565 (N_16565,N_13643,N_13139);
or U16566 (N_16566,N_13664,N_13686);
or U16567 (N_16567,N_13580,N_12892);
or U16568 (N_16568,N_13372,N_14804);
or U16569 (N_16569,N_12946,N_13785);
xor U16570 (N_16570,N_14195,N_13665);
and U16571 (N_16571,N_13805,N_13240);
xnor U16572 (N_16572,N_13325,N_14701);
nand U16573 (N_16573,N_12612,N_14402);
and U16574 (N_16574,N_14225,N_14661);
xnor U16575 (N_16575,N_12819,N_13789);
and U16576 (N_16576,N_13841,N_12510);
nand U16577 (N_16577,N_12846,N_14391);
or U16578 (N_16578,N_14511,N_12580);
and U16579 (N_16579,N_13322,N_14866);
xnor U16580 (N_16580,N_14546,N_12986);
nand U16581 (N_16581,N_12820,N_14681);
xnor U16582 (N_16582,N_14040,N_13003);
xor U16583 (N_16583,N_14206,N_13887);
nand U16584 (N_16584,N_14486,N_12591);
and U16585 (N_16585,N_13217,N_12631);
or U16586 (N_16586,N_14484,N_12845);
or U16587 (N_16587,N_13165,N_12621);
and U16588 (N_16588,N_13873,N_14724);
nor U16589 (N_16589,N_14283,N_13703);
nor U16590 (N_16590,N_12521,N_12904);
nor U16591 (N_16591,N_13523,N_12984);
xnor U16592 (N_16592,N_14849,N_13005);
nand U16593 (N_16593,N_12864,N_13373);
nand U16594 (N_16594,N_14479,N_13553);
xnor U16595 (N_16595,N_12996,N_13191);
xnor U16596 (N_16596,N_14518,N_12518);
or U16597 (N_16597,N_14929,N_13944);
and U16598 (N_16598,N_14232,N_14817);
nor U16599 (N_16599,N_12950,N_14893);
and U16600 (N_16600,N_14932,N_14922);
or U16601 (N_16601,N_13285,N_13182);
nor U16602 (N_16602,N_12972,N_12865);
or U16603 (N_16603,N_14555,N_14621);
and U16604 (N_16604,N_12642,N_14765);
or U16605 (N_16605,N_14768,N_13864);
nor U16606 (N_16606,N_13661,N_14279);
and U16607 (N_16607,N_13951,N_12620);
or U16608 (N_16608,N_13936,N_14564);
and U16609 (N_16609,N_14495,N_12845);
or U16610 (N_16610,N_12960,N_14482);
nand U16611 (N_16611,N_14305,N_14701);
xor U16612 (N_16612,N_12514,N_14726);
xnor U16613 (N_16613,N_13048,N_12517);
xor U16614 (N_16614,N_13620,N_14821);
and U16615 (N_16615,N_14771,N_13596);
nor U16616 (N_16616,N_13234,N_14270);
and U16617 (N_16617,N_12987,N_14377);
nor U16618 (N_16618,N_14443,N_13723);
and U16619 (N_16619,N_14686,N_14738);
xor U16620 (N_16620,N_13948,N_12990);
or U16621 (N_16621,N_14286,N_14678);
and U16622 (N_16622,N_14620,N_13429);
or U16623 (N_16623,N_14339,N_13604);
or U16624 (N_16624,N_14938,N_12686);
nand U16625 (N_16625,N_14946,N_13270);
or U16626 (N_16626,N_12981,N_14447);
xor U16627 (N_16627,N_12521,N_13025);
nor U16628 (N_16628,N_14429,N_12905);
and U16629 (N_16629,N_12613,N_13639);
and U16630 (N_16630,N_12798,N_14909);
nand U16631 (N_16631,N_14498,N_13936);
nor U16632 (N_16632,N_14317,N_13218);
xor U16633 (N_16633,N_14290,N_14364);
nor U16634 (N_16634,N_14958,N_14185);
xnor U16635 (N_16635,N_14558,N_12839);
nand U16636 (N_16636,N_12572,N_13128);
nand U16637 (N_16637,N_14253,N_13769);
nor U16638 (N_16638,N_12624,N_14813);
nand U16639 (N_16639,N_14822,N_13046);
or U16640 (N_16640,N_13401,N_14450);
nor U16641 (N_16641,N_14370,N_12622);
and U16642 (N_16642,N_13360,N_14305);
nand U16643 (N_16643,N_13945,N_12787);
nand U16644 (N_16644,N_14299,N_13813);
xor U16645 (N_16645,N_12804,N_13142);
nor U16646 (N_16646,N_13388,N_14722);
nor U16647 (N_16647,N_13129,N_13748);
nor U16648 (N_16648,N_14862,N_13031);
nand U16649 (N_16649,N_14837,N_14725);
nand U16650 (N_16650,N_12737,N_13366);
and U16651 (N_16651,N_13883,N_14240);
xnor U16652 (N_16652,N_13797,N_14280);
and U16653 (N_16653,N_14131,N_14704);
or U16654 (N_16654,N_13216,N_12942);
and U16655 (N_16655,N_13510,N_12706);
xor U16656 (N_16656,N_12946,N_13082);
and U16657 (N_16657,N_13785,N_13315);
or U16658 (N_16658,N_12686,N_14781);
and U16659 (N_16659,N_13501,N_13083);
or U16660 (N_16660,N_12843,N_13475);
nor U16661 (N_16661,N_14265,N_14872);
nor U16662 (N_16662,N_14079,N_13636);
xor U16663 (N_16663,N_13179,N_14856);
and U16664 (N_16664,N_13348,N_12898);
and U16665 (N_16665,N_13256,N_13626);
and U16666 (N_16666,N_12793,N_14937);
nor U16667 (N_16667,N_13239,N_14208);
or U16668 (N_16668,N_13337,N_13099);
nand U16669 (N_16669,N_14423,N_13951);
nor U16670 (N_16670,N_14053,N_12870);
and U16671 (N_16671,N_12554,N_12935);
nor U16672 (N_16672,N_13848,N_14568);
or U16673 (N_16673,N_14136,N_13419);
or U16674 (N_16674,N_14031,N_12681);
nand U16675 (N_16675,N_12911,N_13765);
nand U16676 (N_16676,N_14181,N_12583);
and U16677 (N_16677,N_14064,N_14247);
nand U16678 (N_16678,N_13192,N_14298);
xnor U16679 (N_16679,N_14468,N_14121);
nand U16680 (N_16680,N_13191,N_12568);
nor U16681 (N_16681,N_13503,N_13370);
and U16682 (N_16682,N_14053,N_14453);
nor U16683 (N_16683,N_13907,N_13452);
and U16684 (N_16684,N_13559,N_14130);
xnor U16685 (N_16685,N_13937,N_14201);
nor U16686 (N_16686,N_13200,N_14076);
nor U16687 (N_16687,N_13349,N_14139);
xnor U16688 (N_16688,N_14733,N_12630);
or U16689 (N_16689,N_12896,N_14914);
and U16690 (N_16690,N_13034,N_12601);
nand U16691 (N_16691,N_13106,N_14906);
and U16692 (N_16692,N_14495,N_14975);
nor U16693 (N_16693,N_13248,N_14295);
or U16694 (N_16694,N_13331,N_14928);
nor U16695 (N_16695,N_13538,N_14404);
nor U16696 (N_16696,N_13472,N_13292);
nand U16697 (N_16697,N_13516,N_13795);
nor U16698 (N_16698,N_13786,N_14600);
and U16699 (N_16699,N_14978,N_13703);
or U16700 (N_16700,N_14437,N_14054);
xor U16701 (N_16701,N_14723,N_13761);
nand U16702 (N_16702,N_13164,N_14683);
nor U16703 (N_16703,N_12943,N_13212);
xor U16704 (N_16704,N_13350,N_13722);
xor U16705 (N_16705,N_14597,N_13184);
nor U16706 (N_16706,N_14915,N_12698);
nor U16707 (N_16707,N_12796,N_13825);
nor U16708 (N_16708,N_12519,N_14285);
and U16709 (N_16709,N_14309,N_14992);
xor U16710 (N_16710,N_12699,N_13953);
nand U16711 (N_16711,N_12621,N_14024);
xor U16712 (N_16712,N_13333,N_14532);
nand U16713 (N_16713,N_14477,N_14886);
or U16714 (N_16714,N_14958,N_14204);
xnor U16715 (N_16715,N_14030,N_13444);
nor U16716 (N_16716,N_14599,N_13115);
xnor U16717 (N_16717,N_12774,N_13839);
and U16718 (N_16718,N_14169,N_13101);
nand U16719 (N_16719,N_13340,N_13914);
and U16720 (N_16720,N_13575,N_12765);
xnor U16721 (N_16721,N_13815,N_13460);
and U16722 (N_16722,N_13523,N_14929);
and U16723 (N_16723,N_13606,N_13122);
nor U16724 (N_16724,N_13178,N_14361);
nand U16725 (N_16725,N_14306,N_12915);
nand U16726 (N_16726,N_14314,N_14152);
nand U16727 (N_16727,N_12695,N_13674);
and U16728 (N_16728,N_14509,N_13290);
xnor U16729 (N_16729,N_12672,N_14060);
nor U16730 (N_16730,N_13984,N_13729);
nand U16731 (N_16731,N_14707,N_12955);
xor U16732 (N_16732,N_12697,N_12891);
nand U16733 (N_16733,N_13752,N_14633);
nand U16734 (N_16734,N_12764,N_12814);
nor U16735 (N_16735,N_13577,N_12614);
or U16736 (N_16736,N_14478,N_13024);
nor U16737 (N_16737,N_14377,N_13780);
xnor U16738 (N_16738,N_13441,N_13421);
or U16739 (N_16739,N_13100,N_14821);
and U16740 (N_16740,N_14600,N_13473);
nor U16741 (N_16741,N_12578,N_14146);
nor U16742 (N_16742,N_13093,N_13427);
and U16743 (N_16743,N_12637,N_14126);
or U16744 (N_16744,N_13106,N_12825);
nand U16745 (N_16745,N_12730,N_14335);
nand U16746 (N_16746,N_13586,N_14762);
nor U16747 (N_16747,N_13014,N_13957);
xnor U16748 (N_16748,N_13187,N_14112);
or U16749 (N_16749,N_13222,N_14579);
nor U16750 (N_16750,N_14937,N_12760);
and U16751 (N_16751,N_14590,N_14676);
nand U16752 (N_16752,N_13601,N_14988);
nand U16753 (N_16753,N_13226,N_12576);
nor U16754 (N_16754,N_14810,N_14886);
and U16755 (N_16755,N_12624,N_13614);
nand U16756 (N_16756,N_13689,N_13462);
nand U16757 (N_16757,N_14467,N_13083);
nand U16758 (N_16758,N_13569,N_13702);
or U16759 (N_16759,N_14241,N_14686);
xor U16760 (N_16760,N_13249,N_13443);
or U16761 (N_16761,N_14558,N_14533);
or U16762 (N_16762,N_14437,N_14418);
or U16763 (N_16763,N_13948,N_13681);
nor U16764 (N_16764,N_13549,N_13081);
xor U16765 (N_16765,N_14807,N_13824);
xnor U16766 (N_16766,N_12553,N_13132);
xor U16767 (N_16767,N_12820,N_12800);
or U16768 (N_16768,N_14110,N_13064);
xor U16769 (N_16769,N_13436,N_12512);
and U16770 (N_16770,N_14529,N_13328);
nor U16771 (N_16771,N_14873,N_14491);
xnor U16772 (N_16772,N_14572,N_14148);
xor U16773 (N_16773,N_14886,N_14035);
nor U16774 (N_16774,N_14438,N_12818);
or U16775 (N_16775,N_14386,N_12576);
or U16776 (N_16776,N_12676,N_14118);
nor U16777 (N_16777,N_13364,N_13665);
or U16778 (N_16778,N_14344,N_13348);
nand U16779 (N_16779,N_13761,N_14414);
and U16780 (N_16780,N_13981,N_14901);
nor U16781 (N_16781,N_14546,N_14391);
nor U16782 (N_16782,N_14743,N_12838);
and U16783 (N_16783,N_12661,N_13666);
nor U16784 (N_16784,N_12660,N_13210);
and U16785 (N_16785,N_14178,N_12754);
nand U16786 (N_16786,N_13811,N_12563);
and U16787 (N_16787,N_14843,N_14842);
or U16788 (N_16788,N_13361,N_14383);
and U16789 (N_16789,N_14858,N_14451);
or U16790 (N_16790,N_14521,N_12742);
xor U16791 (N_16791,N_14245,N_13774);
and U16792 (N_16792,N_13474,N_14754);
nor U16793 (N_16793,N_14832,N_14969);
nand U16794 (N_16794,N_14126,N_13578);
nand U16795 (N_16795,N_14686,N_13716);
or U16796 (N_16796,N_13981,N_14795);
nand U16797 (N_16797,N_13438,N_12747);
xnor U16798 (N_16798,N_14514,N_13446);
or U16799 (N_16799,N_14613,N_13933);
xor U16800 (N_16800,N_14548,N_13008);
nand U16801 (N_16801,N_13420,N_14710);
nor U16802 (N_16802,N_14916,N_14214);
and U16803 (N_16803,N_12994,N_13700);
xnor U16804 (N_16804,N_13216,N_13437);
nor U16805 (N_16805,N_14913,N_13710);
or U16806 (N_16806,N_14101,N_14254);
xor U16807 (N_16807,N_14669,N_14988);
or U16808 (N_16808,N_14152,N_14463);
nor U16809 (N_16809,N_14688,N_13988);
or U16810 (N_16810,N_13088,N_13289);
or U16811 (N_16811,N_14444,N_13769);
nand U16812 (N_16812,N_13067,N_14459);
and U16813 (N_16813,N_14933,N_13551);
and U16814 (N_16814,N_14088,N_14888);
nor U16815 (N_16815,N_12834,N_13676);
or U16816 (N_16816,N_12786,N_12790);
or U16817 (N_16817,N_12508,N_14262);
or U16818 (N_16818,N_12957,N_12565);
and U16819 (N_16819,N_13147,N_13251);
xnor U16820 (N_16820,N_14813,N_13011);
xor U16821 (N_16821,N_13438,N_13488);
nand U16822 (N_16822,N_14980,N_14727);
nand U16823 (N_16823,N_13981,N_14702);
nor U16824 (N_16824,N_14918,N_13417);
or U16825 (N_16825,N_13498,N_12755);
nand U16826 (N_16826,N_13363,N_14381);
and U16827 (N_16827,N_14767,N_12910);
nor U16828 (N_16828,N_14379,N_13323);
nand U16829 (N_16829,N_12678,N_14315);
nor U16830 (N_16830,N_14618,N_12724);
nand U16831 (N_16831,N_13558,N_13318);
xnor U16832 (N_16832,N_13201,N_12683);
nor U16833 (N_16833,N_14765,N_13182);
and U16834 (N_16834,N_13399,N_13628);
or U16835 (N_16835,N_13069,N_14353);
or U16836 (N_16836,N_14788,N_14383);
or U16837 (N_16837,N_13335,N_13705);
and U16838 (N_16838,N_14130,N_12696);
nand U16839 (N_16839,N_14272,N_12588);
nand U16840 (N_16840,N_13692,N_13195);
or U16841 (N_16841,N_12745,N_14164);
nor U16842 (N_16842,N_14515,N_13545);
nor U16843 (N_16843,N_14161,N_13433);
or U16844 (N_16844,N_14615,N_13366);
nor U16845 (N_16845,N_14843,N_13220);
and U16846 (N_16846,N_14522,N_14276);
and U16847 (N_16847,N_14164,N_13104);
xnor U16848 (N_16848,N_13191,N_14625);
or U16849 (N_16849,N_14260,N_13148);
or U16850 (N_16850,N_13592,N_12747);
or U16851 (N_16851,N_14754,N_14013);
and U16852 (N_16852,N_13315,N_14237);
xnor U16853 (N_16853,N_13547,N_13476);
nand U16854 (N_16854,N_12841,N_13736);
xnor U16855 (N_16855,N_13179,N_12615);
or U16856 (N_16856,N_13283,N_14072);
nor U16857 (N_16857,N_13078,N_14383);
and U16858 (N_16858,N_14132,N_14807);
xnor U16859 (N_16859,N_13339,N_14347);
nor U16860 (N_16860,N_13738,N_12680);
or U16861 (N_16861,N_13810,N_12652);
nor U16862 (N_16862,N_14073,N_13186);
and U16863 (N_16863,N_12758,N_13531);
xnor U16864 (N_16864,N_14983,N_12785);
or U16865 (N_16865,N_14787,N_14496);
nor U16866 (N_16866,N_14182,N_13668);
xnor U16867 (N_16867,N_12956,N_14312);
and U16868 (N_16868,N_14626,N_13557);
or U16869 (N_16869,N_14281,N_13139);
and U16870 (N_16870,N_14890,N_13229);
or U16871 (N_16871,N_14946,N_14158);
and U16872 (N_16872,N_13920,N_12661);
or U16873 (N_16873,N_14330,N_14984);
nor U16874 (N_16874,N_13422,N_13566);
or U16875 (N_16875,N_12956,N_14813);
xor U16876 (N_16876,N_13273,N_14138);
nand U16877 (N_16877,N_14529,N_13784);
xnor U16878 (N_16878,N_14349,N_13705);
nand U16879 (N_16879,N_13394,N_13455);
and U16880 (N_16880,N_13254,N_13792);
xnor U16881 (N_16881,N_12797,N_13352);
nor U16882 (N_16882,N_14624,N_14036);
nor U16883 (N_16883,N_14517,N_12577);
and U16884 (N_16884,N_12713,N_12515);
nor U16885 (N_16885,N_14412,N_13527);
nand U16886 (N_16886,N_12935,N_14760);
nor U16887 (N_16887,N_14498,N_13866);
and U16888 (N_16888,N_14289,N_14655);
nor U16889 (N_16889,N_14698,N_13120);
or U16890 (N_16890,N_12703,N_13742);
and U16891 (N_16891,N_14223,N_14392);
or U16892 (N_16892,N_14871,N_13370);
nand U16893 (N_16893,N_13211,N_13856);
xor U16894 (N_16894,N_13994,N_14466);
nand U16895 (N_16895,N_13535,N_12981);
nor U16896 (N_16896,N_13858,N_14449);
and U16897 (N_16897,N_14995,N_14241);
or U16898 (N_16898,N_14667,N_13432);
nor U16899 (N_16899,N_12640,N_14998);
nor U16900 (N_16900,N_13424,N_12845);
or U16901 (N_16901,N_13448,N_14576);
and U16902 (N_16902,N_13348,N_14469);
xnor U16903 (N_16903,N_13314,N_13772);
or U16904 (N_16904,N_14796,N_12864);
or U16905 (N_16905,N_13752,N_14104);
nor U16906 (N_16906,N_12883,N_14972);
or U16907 (N_16907,N_13513,N_12628);
nand U16908 (N_16908,N_13501,N_13014);
nor U16909 (N_16909,N_12740,N_14788);
nand U16910 (N_16910,N_13780,N_14263);
and U16911 (N_16911,N_13292,N_12993);
or U16912 (N_16912,N_13405,N_13543);
and U16913 (N_16913,N_13122,N_12567);
xnor U16914 (N_16914,N_13598,N_14285);
nand U16915 (N_16915,N_14384,N_12944);
nand U16916 (N_16916,N_12500,N_14879);
and U16917 (N_16917,N_14545,N_13474);
nand U16918 (N_16918,N_14735,N_13624);
or U16919 (N_16919,N_12584,N_13969);
or U16920 (N_16920,N_13435,N_13716);
xnor U16921 (N_16921,N_12958,N_14159);
xor U16922 (N_16922,N_14287,N_14828);
nand U16923 (N_16923,N_13838,N_14604);
and U16924 (N_16924,N_12571,N_12977);
nand U16925 (N_16925,N_13377,N_12952);
and U16926 (N_16926,N_13203,N_14760);
xnor U16927 (N_16927,N_14694,N_14673);
or U16928 (N_16928,N_13602,N_12673);
nand U16929 (N_16929,N_13484,N_12503);
and U16930 (N_16930,N_14874,N_12616);
and U16931 (N_16931,N_13782,N_14950);
or U16932 (N_16932,N_13815,N_14663);
nor U16933 (N_16933,N_13932,N_14408);
nor U16934 (N_16934,N_12759,N_14019);
nor U16935 (N_16935,N_13852,N_13720);
nand U16936 (N_16936,N_13734,N_14205);
nor U16937 (N_16937,N_14833,N_14326);
nor U16938 (N_16938,N_14785,N_13214);
nor U16939 (N_16939,N_14536,N_14965);
or U16940 (N_16940,N_12526,N_13105);
nor U16941 (N_16941,N_13691,N_13022);
and U16942 (N_16942,N_14535,N_14747);
and U16943 (N_16943,N_13998,N_13520);
and U16944 (N_16944,N_12830,N_12501);
xor U16945 (N_16945,N_14620,N_13360);
xnor U16946 (N_16946,N_14882,N_14724);
xnor U16947 (N_16947,N_13301,N_13574);
nand U16948 (N_16948,N_13322,N_12883);
xnor U16949 (N_16949,N_14230,N_13507);
nand U16950 (N_16950,N_12565,N_13421);
and U16951 (N_16951,N_14775,N_14752);
nand U16952 (N_16952,N_14778,N_12546);
nor U16953 (N_16953,N_13039,N_12550);
and U16954 (N_16954,N_12667,N_14810);
nor U16955 (N_16955,N_13931,N_14981);
nor U16956 (N_16956,N_14522,N_12643);
nor U16957 (N_16957,N_14084,N_13391);
nand U16958 (N_16958,N_12674,N_13669);
and U16959 (N_16959,N_13548,N_13273);
and U16960 (N_16960,N_13830,N_14608);
and U16961 (N_16961,N_13705,N_12849);
nor U16962 (N_16962,N_14271,N_13624);
nor U16963 (N_16963,N_12865,N_13034);
nor U16964 (N_16964,N_12683,N_13007);
or U16965 (N_16965,N_14855,N_13319);
nand U16966 (N_16966,N_14237,N_12780);
and U16967 (N_16967,N_14969,N_13862);
nor U16968 (N_16968,N_14641,N_14596);
nor U16969 (N_16969,N_13759,N_13426);
nand U16970 (N_16970,N_12528,N_14705);
or U16971 (N_16971,N_14449,N_14955);
or U16972 (N_16972,N_14484,N_14882);
xor U16973 (N_16973,N_12720,N_14928);
nor U16974 (N_16974,N_14956,N_13630);
or U16975 (N_16975,N_13054,N_14815);
nor U16976 (N_16976,N_13447,N_12900);
and U16977 (N_16977,N_13077,N_12674);
nor U16978 (N_16978,N_13697,N_12811);
and U16979 (N_16979,N_13338,N_14225);
nand U16980 (N_16980,N_14828,N_13749);
nand U16981 (N_16981,N_13352,N_13510);
or U16982 (N_16982,N_12971,N_12502);
nand U16983 (N_16983,N_12616,N_13596);
xor U16984 (N_16984,N_13170,N_13975);
and U16985 (N_16985,N_13645,N_14129);
or U16986 (N_16986,N_14282,N_13341);
and U16987 (N_16987,N_13469,N_13909);
nor U16988 (N_16988,N_14314,N_13614);
or U16989 (N_16989,N_14929,N_14667);
xnor U16990 (N_16990,N_14275,N_14858);
and U16991 (N_16991,N_13575,N_13955);
xor U16992 (N_16992,N_13474,N_13457);
xor U16993 (N_16993,N_13790,N_13488);
or U16994 (N_16994,N_14522,N_12562);
or U16995 (N_16995,N_13147,N_14516);
nor U16996 (N_16996,N_14032,N_13399);
or U16997 (N_16997,N_13878,N_14966);
and U16998 (N_16998,N_14169,N_14662);
or U16999 (N_16999,N_13946,N_13406);
or U17000 (N_17000,N_13801,N_14990);
nand U17001 (N_17001,N_12873,N_14898);
nand U17002 (N_17002,N_14116,N_14030);
nor U17003 (N_17003,N_14365,N_12929);
nor U17004 (N_17004,N_12718,N_14966);
nor U17005 (N_17005,N_13335,N_13117);
and U17006 (N_17006,N_14364,N_12512);
or U17007 (N_17007,N_12966,N_13188);
or U17008 (N_17008,N_14035,N_14680);
nand U17009 (N_17009,N_14793,N_13090);
nand U17010 (N_17010,N_12846,N_14524);
and U17011 (N_17011,N_14561,N_14300);
nand U17012 (N_17012,N_13363,N_13940);
nor U17013 (N_17013,N_13243,N_13558);
nor U17014 (N_17014,N_14801,N_12767);
or U17015 (N_17015,N_14596,N_13760);
or U17016 (N_17016,N_14942,N_14159);
or U17017 (N_17017,N_12726,N_12916);
nor U17018 (N_17018,N_12921,N_13153);
nor U17019 (N_17019,N_12852,N_14306);
nand U17020 (N_17020,N_13230,N_12755);
xnor U17021 (N_17021,N_14687,N_14039);
and U17022 (N_17022,N_14838,N_14605);
nand U17023 (N_17023,N_14675,N_12743);
nand U17024 (N_17024,N_13974,N_12628);
nand U17025 (N_17025,N_13019,N_14595);
nor U17026 (N_17026,N_14008,N_12516);
or U17027 (N_17027,N_13052,N_13993);
or U17028 (N_17028,N_14481,N_12878);
xor U17029 (N_17029,N_14896,N_13088);
nand U17030 (N_17030,N_14395,N_14687);
nand U17031 (N_17031,N_14128,N_12984);
xnor U17032 (N_17032,N_13226,N_13897);
nor U17033 (N_17033,N_14328,N_12976);
nor U17034 (N_17034,N_13842,N_13752);
xor U17035 (N_17035,N_13267,N_13328);
xor U17036 (N_17036,N_13877,N_14817);
nor U17037 (N_17037,N_14164,N_12617);
or U17038 (N_17038,N_12935,N_13201);
or U17039 (N_17039,N_14015,N_14258);
nand U17040 (N_17040,N_12989,N_14238);
and U17041 (N_17041,N_14039,N_13309);
nor U17042 (N_17042,N_13563,N_13307);
nor U17043 (N_17043,N_14855,N_12831);
xnor U17044 (N_17044,N_12617,N_14489);
nor U17045 (N_17045,N_14620,N_14150);
and U17046 (N_17046,N_14607,N_12625);
or U17047 (N_17047,N_12500,N_14565);
or U17048 (N_17048,N_13339,N_13487);
xor U17049 (N_17049,N_14951,N_13764);
and U17050 (N_17050,N_12845,N_14092);
nor U17051 (N_17051,N_14950,N_14789);
or U17052 (N_17052,N_13238,N_14593);
nor U17053 (N_17053,N_13795,N_13396);
or U17054 (N_17054,N_14470,N_13959);
or U17055 (N_17055,N_13836,N_13521);
and U17056 (N_17056,N_12823,N_14977);
and U17057 (N_17057,N_14177,N_14539);
nand U17058 (N_17058,N_12977,N_12649);
and U17059 (N_17059,N_12565,N_14378);
xnor U17060 (N_17060,N_13466,N_14572);
nand U17061 (N_17061,N_13250,N_13291);
nand U17062 (N_17062,N_13714,N_14211);
nand U17063 (N_17063,N_14570,N_14721);
nand U17064 (N_17064,N_13535,N_14518);
nor U17065 (N_17065,N_13869,N_13369);
nand U17066 (N_17066,N_14723,N_14810);
and U17067 (N_17067,N_14652,N_14185);
xor U17068 (N_17068,N_13056,N_14026);
nand U17069 (N_17069,N_13540,N_12530);
and U17070 (N_17070,N_13918,N_13154);
xnor U17071 (N_17071,N_14658,N_14872);
nor U17072 (N_17072,N_12886,N_13634);
xor U17073 (N_17073,N_13424,N_14965);
xor U17074 (N_17074,N_14609,N_13759);
or U17075 (N_17075,N_14184,N_14786);
xnor U17076 (N_17076,N_13191,N_13336);
xor U17077 (N_17077,N_14216,N_14077);
or U17078 (N_17078,N_14716,N_14606);
xnor U17079 (N_17079,N_12828,N_13368);
or U17080 (N_17080,N_13246,N_14176);
nor U17081 (N_17081,N_13769,N_12770);
nor U17082 (N_17082,N_13541,N_12962);
nand U17083 (N_17083,N_12969,N_14458);
xor U17084 (N_17084,N_13729,N_12928);
xor U17085 (N_17085,N_13255,N_13795);
nor U17086 (N_17086,N_12807,N_12981);
xor U17087 (N_17087,N_13716,N_14673);
xnor U17088 (N_17088,N_13589,N_13037);
and U17089 (N_17089,N_13571,N_14502);
or U17090 (N_17090,N_13529,N_14371);
nor U17091 (N_17091,N_13032,N_12945);
nor U17092 (N_17092,N_12962,N_13805);
nor U17093 (N_17093,N_14892,N_14492);
or U17094 (N_17094,N_13489,N_13393);
xor U17095 (N_17095,N_12764,N_12938);
nor U17096 (N_17096,N_13425,N_12801);
or U17097 (N_17097,N_14688,N_13876);
xor U17098 (N_17098,N_13337,N_14247);
xnor U17099 (N_17099,N_14683,N_12515);
nor U17100 (N_17100,N_12613,N_13820);
or U17101 (N_17101,N_12577,N_13428);
nand U17102 (N_17102,N_13880,N_13107);
nand U17103 (N_17103,N_12739,N_14758);
nor U17104 (N_17104,N_13262,N_14952);
nor U17105 (N_17105,N_14315,N_13712);
nor U17106 (N_17106,N_12655,N_13999);
nand U17107 (N_17107,N_12605,N_12612);
and U17108 (N_17108,N_13765,N_13339);
nor U17109 (N_17109,N_14037,N_14185);
xnor U17110 (N_17110,N_14930,N_12686);
and U17111 (N_17111,N_13513,N_14521);
nor U17112 (N_17112,N_14495,N_14554);
xor U17113 (N_17113,N_14764,N_14995);
xor U17114 (N_17114,N_13154,N_13954);
or U17115 (N_17115,N_13316,N_14292);
nor U17116 (N_17116,N_14354,N_13818);
and U17117 (N_17117,N_13181,N_14835);
nand U17118 (N_17118,N_14844,N_12802);
nor U17119 (N_17119,N_14649,N_13451);
or U17120 (N_17120,N_14636,N_14501);
nand U17121 (N_17121,N_13424,N_12628);
or U17122 (N_17122,N_14899,N_13103);
nand U17123 (N_17123,N_14976,N_12924);
nor U17124 (N_17124,N_12573,N_14989);
xnor U17125 (N_17125,N_13310,N_14959);
xnor U17126 (N_17126,N_14758,N_13484);
and U17127 (N_17127,N_14370,N_12623);
and U17128 (N_17128,N_13798,N_14298);
xnor U17129 (N_17129,N_12841,N_12643);
xor U17130 (N_17130,N_14526,N_14710);
and U17131 (N_17131,N_14500,N_13727);
and U17132 (N_17132,N_13061,N_14422);
or U17133 (N_17133,N_14556,N_14176);
nor U17134 (N_17134,N_12511,N_14041);
nand U17135 (N_17135,N_12559,N_12867);
and U17136 (N_17136,N_14686,N_12977);
nor U17137 (N_17137,N_13440,N_13178);
xor U17138 (N_17138,N_12900,N_13912);
xnor U17139 (N_17139,N_13953,N_14996);
nor U17140 (N_17140,N_14094,N_13902);
xnor U17141 (N_17141,N_13660,N_12967);
xnor U17142 (N_17142,N_14304,N_13163);
xnor U17143 (N_17143,N_14728,N_14849);
nor U17144 (N_17144,N_13966,N_14996);
nand U17145 (N_17145,N_13767,N_14821);
xor U17146 (N_17146,N_14204,N_13741);
nand U17147 (N_17147,N_13054,N_13711);
nor U17148 (N_17148,N_12779,N_13443);
nor U17149 (N_17149,N_14769,N_14174);
xnor U17150 (N_17150,N_14403,N_13430);
or U17151 (N_17151,N_14105,N_13532);
nand U17152 (N_17152,N_13497,N_14059);
or U17153 (N_17153,N_14714,N_13096);
and U17154 (N_17154,N_13439,N_13869);
xnor U17155 (N_17155,N_13120,N_14298);
nand U17156 (N_17156,N_14884,N_12960);
or U17157 (N_17157,N_13322,N_13900);
nand U17158 (N_17158,N_14001,N_13751);
xnor U17159 (N_17159,N_14181,N_14492);
xnor U17160 (N_17160,N_14590,N_12669);
or U17161 (N_17161,N_13326,N_12651);
and U17162 (N_17162,N_13741,N_13750);
nor U17163 (N_17163,N_13962,N_14656);
and U17164 (N_17164,N_12688,N_13655);
nand U17165 (N_17165,N_14853,N_14295);
or U17166 (N_17166,N_13526,N_13143);
nor U17167 (N_17167,N_13268,N_14808);
and U17168 (N_17168,N_13055,N_13105);
nand U17169 (N_17169,N_14584,N_13117);
nand U17170 (N_17170,N_13295,N_13264);
xnor U17171 (N_17171,N_13838,N_12760);
or U17172 (N_17172,N_14299,N_14127);
xor U17173 (N_17173,N_13225,N_12983);
xor U17174 (N_17174,N_14262,N_14919);
or U17175 (N_17175,N_12539,N_12530);
xnor U17176 (N_17176,N_13169,N_13905);
or U17177 (N_17177,N_13801,N_13492);
and U17178 (N_17178,N_14346,N_13735);
or U17179 (N_17179,N_12682,N_13699);
or U17180 (N_17180,N_13728,N_14086);
and U17181 (N_17181,N_14794,N_14697);
nand U17182 (N_17182,N_14558,N_13817);
and U17183 (N_17183,N_13400,N_14315);
xnor U17184 (N_17184,N_13267,N_14132);
or U17185 (N_17185,N_14769,N_13166);
and U17186 (N_17186,N_12972,N_14672);
or U17187 (N_17187,N_13067,N_12595);
nor U17188 (N_17188,N_14571,N_12991);
nor U17189 (N_17189,N_13964,N_12624);
xnor U17190 (N_17190,N_14309,N_14170);
or U17191 (N_17191,N_14070,N_12732);
or U17192 (N_17192,N_13040,N_14911);
nand U17193 (N_17193,N_13196,N_14215);
or U17194 (N_17194,N_14632,N_12556);
nor U17195 (N_17195,N_14001,N_14064);
and U17196 (N_17196,N_13536,N_14108);
xnor U17197 (N_17197,N_13408,N_13804);
and U17198 (N_17198,N_14929,N_12541);
or U17199 (N_17199,N_14660,N_14412);
or U17200 (N_17200,N_13466,N_14089);
and U17201 (N_17201,N_12882,N_14264);
nor U17202 (N_17202,N_13952,N_13291);
and U17203 (N_17203,N_14061,N_13199);
and U17204 (N_17204,N_12824,N_12782);
nand U17205 (N_17205,N_13313,N_13279);
or U17206 (N_17206,N_13766,N_13007);
nand U17207 (N_17207,N_13295,N_14207);
and U17208 (N_17208,N_14724,N_13122);
xor U17209 (N_17209,N_12614,N_12608);
nor U17210 (N_17210,N_14068,N_14994);
nand U17211 (N_17211,N_14734,N_13305);
or U17212 (N_17212,N_12622,N_14148);
nor U17213 (N_17213,N_14876,N_13529);
nor U17214 (N_17214,N_13490,N_14201);
nand U17215 (N_17215,N_12680,N_12801);
nor U17216 (N_17216,N_14090,N_14069);
and U17217 (N_17217,N_13767,N_12800);
nand U17218 (N_17218,N_13043,N_13484);
or U17219 (N_17219,N_13603,N_13636);
and U17220 (N_17220,N_14971,N_14087);
nor U17221 (N_17221,N_14204,N_14955);
and U17222 (N_17222,N_14802,N_13542);
nor U17223 (N_17223,N_14259,N_14687);
or U17224 (N_17224,N_14005,N_14580);
xnor U17225 (N_17225,N_14630,N_13701);
xnor U17226 (N_17226,N_13492,N_13212);
nor U17227 (N_17227,N_12683,N_12561);
nor U17228 (N_17228,N_14268,N_13826);
nand U17229 (N_17229,N_14150,N_13009);
nand U17230 (N_17230,N_13545,N_14110);
nor U17231 (N_17231,N_13499,N_12852);
nor U17232 (N_17232,N_12822,N_13313);
nand U17233 (N_17233,N_13754,N_14766);
nand U17234 (N_17234,N_12729,N_14930);
xnor U17235 (N_17235,N_13511,N_13029);
nor U17236 (N_17236,N_14761,N_14769);
nand U17237 (N_17237,N_13412,N_13814);
or U17238 (N_17238,N_14758,N_14028);
xor U17239 (N_17239,N_13054,N_13471);
nand U17240 (N_17240,N_14653,N_12983);
nand U17241 (N_17241,N_13464,N_14635);
nand U17242 (N_17242,N_14842,N_13094);
nor U17243 (N_17243,N_13077,N_12858);
xnor U17244 (N_17244,N_12600,N_14680);
nand U17245 (N_17245,N_12664,N_13136);
and U17246 (N_17246,N_13123,N_14335);
xor U17247 (N_17247,N_14554,N_14299);
xor U17248 (N_17248,N_13911,N_12835);
and U17249 (N_17249,N_14782,N_14223);
xor U17250 (N_17250,N_14940,N_14375);
nor U17251 (N_17251,N_13835,N_14525);
nor U17252 (N_17252,N_13426,N_13906);
nand U17253 (N_17253,N_14522,N_13952);
and U17254 (N_17254,N_14383,N_13964);
xnor U17255 (N_17255,N_13617,N_14876);
and U17256 (N_17256,N_13178,N_14328);
xor U17257 (N_17257,N_14682,N_12634);
nor U17258 (N_17258,N_12559,N_14886);
nor U17259 (N_17259,N_13966,N_14294);
or U17260 (N_17260,N_13515,N_13611);
or U17261 (N_17261,N_14745,N_13503);
xnor U17262 (N_17262,N_14090,N_12781);
and U17263 (N_17263,N_14026,N_13316);
nand U17264 (N_17264,N_13613,N_13331);
and U17265 (N_17265,N_14923,N_13551);
xnor U17266 (N_17266,N_14002,N_12500);
or U17267 (N_17267,N_13309,N_14893);
xnor U17268 (N_17268,N_13624,N_14428);
and U17269 (N_17269,N_14240,N_14697);
and U17270 (N_17270,N_12759,N_13484);
or U17271 (N_17271,N_13567,N_13254);
nor U17272 (N_17272,N_14625,N_14302);
xor U17273 (N_17273,N_13349,N_14894);
xor U17274 (N_17274,N_12880,N_13111);
xor U17275 (N_17275,N_14418,N_14765);
and U17276 (N_17276,N_13179,N_14799);
nor U17277 (N_17277,N_14271,N_13207);
or U17278 (N_17278,N_13090,N_14184);
and U17279 (N_17279,N_12752,N_12608);
nand U17280 (N_17280,N_13457,N_12699);
nand U17281 (N_17281,N_13016,N_14995);
xor U17282 (N_17282,N_13322,N_14825);
nor U17283 (N_17283,N_14209,N_12717);
and U17284 (N_17284,N_13106,N_13637);
nor U17285 (N_17285,N_14497,N_14627);
or U17286 (N_17286,N_14658,N_12771);
xnor U17287 (N_17287,N_14729,N_12853);
or U17288 (N_17288,N_13998,N_12578);
nor U17289 (N_17289,N_12992,N_12716);
xnor U17290 (N_17290,N_14695,N_13949);
nand U17291 (N_17291,N_13790,N_14113);
and U17292 (N_17292,N_14703,N_13639);
xor U17293 (N_17293,N_14235,N_12953);
nand U17294 (N_17294,N_14505,N_14818);
nand U17295 (N_17295,N_12779,N_13637);
and U17296 (N_17296,N_12812,N_13871);
nand U17297 (N_17297,N_14996,N_12727);
and U17298 (N_17298,N_13508,N_14988);
and U17299 (N_17299,N_13802,N_13327);
and U17300 (N_17300,N_13257,N_14007);
xor U17301 (N_17301,N_13328,N_14089);
or U17302 (N_17302,N_13548,N_13898);
and U17303 (N_17303,N_14160,N_14884);
nand U17304 (N_17304,N_12907,N_13756);
and U17305 (N_17305,N_14164,N_14045);
xor U17306 (N_17306,N_13495,N_14273);
or U17307 (N_17307,N_13295,N_12681);
and U17308 (N_17308,N_14231,N_14093);
and U17309 (N_17309,N_14003,N_12835);
nand U17310 (N_17310,N_13154,N_13248);
nand U17311 (N_17311,N_14003,N_14659);
and U17312 (N_17312,N_12649,N_14585);
nor U17313 (N_17313,N_13872,N_14884);
nand U17314 (N_17314,N_14913,N_14298);
nand U17315 (N_17315,N_13340,N_14190);
xnor U17316 (N_17316,N_14120,N_14470);
xor U17317 (N_17317,N_12907,N_14821);
and U17318 (N_17318,N_14113,N_13919);
and U17319 (N_17319,N_13525,N_13985);
nand U17320 (N_17320,N_14369,N_14392);
or U17321 (N_17321,N_13836,N_14663);
and U17322 (N_17322,N_14062,N_12780);
xnor U17323 (N_17323,N_14969,N_12800);
nand U17324 (N_17324,N_13806,N_14659);
and U17325 (N_17325,N_12924,N_13598);
or U17326 (N_17326,N_14760,N_13742);
and U17327 (N_17327,N_14826,N_13315);
nand U17328 (N_17328,N_13027,N_12725);
or U17329 (N_17329,N_13104,N_13873);
nor U17330 (N_17330,N_14038,N_14362);
or U17331 (N_17331,N_13585,N_14249);
nand U17332 (N_17332,N_14355,N_13102);
or U17333 (N_17333,N_14969,N_12665);
nor U17334 (N_17334,N_14776,N_12744);
and U17335 (N_17335,N_14727,N_13524);
nor U17336 (N_17336,N_13244,N_13531);
xnor U17337 (N_17337,N_14188,N_14699);
and U17338 (N_17338,N_14549,N_13812);
or U17339 (N_17339,N_13363,N_13810);
nand U17340 (N_17340,N_14986,N_14768);
xnor U17341 (N_17341,N_14405,N_14253);
and U17342 (N_17342,N_14847,N_13829);
nor U17343 (N_17343,N_14207,N_14484);
nor U17344 (N_17344,N_14737,N_12503);
nor U17345 (N_17345,N_14907,N_14677);
xor U17346 (N_17346,N_12989,N_14268);
xor U17347 (N_17347,N_14713,N_14703);
xor U17348 (N_17348,N_14432,N_14530);
or U17349 (N_17349,N_12765,N_14888);
or U17350 (N_17350,N_13435,N_13836);
nand U17351 (N_17351,N_13593,N_14565);
and U17352 (N_17352,N_14136,N_14065);
nand U17353 (N_17353,N_13509,N_13355);
nand U17354 (N_17354,N_13082,N_13775);
and U17355 (N_17355,N_12606,N_13229);
or U17356 (N_17356,N_13521,N_14662);
nand U17357 (N_17357,N_13654,N_12766);
and U17358 (N_17358,N_13223,N_12710);
or U17359 (N_17359,N_14453,N_13217);
nor U17360 (N_17360,N_13307,N_14512);
or U17361 (N_17361,N_13113,N_13746);
nand U17362 (N_17362,N_13591,N_14382);
nand U17363 (N_17363,N_12848,N_13478);
nand U17364 (N_17364,N_13590,N_14869);
or U17365 (N_17365,N_13577,N_13542);
and U17366 (N_17366,N_13132,N_13989);
nor U17367 (N_17367,N_12806,N_13412);
xnor U17368 (N_17368,N_12945,N_14631);
xor U17369 (N_17369,N_14155,N_13547);
xnor U17370 (N_17370,N_13312,N_13061);
or U17371 (N_17371,N_13649,N_14523);
nand U17372 (N_17372,N_14510,N_14279);
nand U17373 (N_17373,N_14074,N_14314);
and U17374 (N_17374,N_14587,N_14693);
xnor U17375 (N_17375,N_14423,N_14332);
nor U17376 (N_17376,N_12658,N_14297);
and U17377 (N_17377,N_14443,N_14840);
nand U17378 (N_17378,N_13072,N_13981);
or U17379 (N_17379,N_12516,N_14048);
nand U17380 (N_17380,N_14772,N_14860);
nor U17381 (N_17381,N_14281,N_14626);
and U17382 (N_17382,N_13996,N_13357);
or U17383 (N_17383,N_14346,N_13183);
nand U17384 (N_17384,N_14874,N_14444);
or U17385 (N_17385,N_14074,N_12664);
and U17386 (N_17386,N_13462,N_13493);
nand U17387 (N_17387,N_14223,N_14935);
xor U17388 (N_17388,N_12933,N_13509);
xor U17389 (N_17389,N_13822,N_13888);
nor U17390 (N_17390,N_14851,N_13108);
xnor U17391 (N_17391,N_13129,N_13475);
nor U17392 (N_17392,N_14862,N_13043);
nand U17393 (N_17393,N_14752,N_14948);
and U17394 (N_17394,N_14130,N_14098);
xor U17395 (N_17395,N_13694,N_14690);
or U17396 (N_17396,N_14820,N_14341);
xnor U17397 (N_17397,N_14430,N_13274);
nor U17398 (N_17398,N_14059,N_13639);
nor U17399 (N_17399,N_14600,N_14873);
nand U17400 (N_17400,N_14557,N_12526);
or U17401 (N_17401,N_13909,N_12993);
nand U17402 (N_17402,N_13898,N_13144);
and U17403 (N_17403,N_12841,N_14980);
nand U17404 (N_17404,N_13703,N_12556);
or U17405 (N_17405,N_13718,N_14105);
xor U17406 (N_17406,N_14415,N_14530);
and U17407 (N_17407,N_13821,N_14145);
xnor U17408 (N_17408,N_13444,N_14710);
nor U17409 (N_17409,N_14864,N_13651);
nand U17410 (N_17410,N_14102,N_14407);
or U17411 (N_17411,N_13228,N_14489);
xor U17412 (N_17412,N_14794,N_14122);
xnor U17413 (N_17413,N_12695,N_14890);
xor U17414 (N_17414,N_13116,N_12764);
or U17415 (N_17415,N_14887,N_14538);
or U17416 (N_17416,N_14724,N_13657);
nor U17417 (N_17417,N_14459,N_14758);
and U17418 (N_17418,N_14846,N_13029);
nor U17419 (N_17419,N_14383,N_13331);
and U17420 (N_17420,N_13093,N_12820);
nor U17421 (N_17421,N_14294,N_14826);
and U17422 (N_17422,N_13153,N_14434);
and U17423 (N_17423,N_13543,N_12846);
nand U17424 (N_17424,N_13094,N_13890);
xnor U17425 (N_17425,N_14389,N_13248);
xnor U17426 (N_17426,N_14090,N_13735);
nor U17427 (N_17427,N_13692,N_12660);
and U17428 (N_17428,N_14078,N_13178);
nand U17429 (N_17429,N_13183,N_13408);
nor U17430 (N_17430,N_12793,N_12856);
nor U17431 (N_17431,N_12610,N_12594);
and U17432 (N_17432,N_12902,N_14395);
xnor U17433 (N_17433,N_13572,N_12888);
and U17434 (N_17434,N_12923,N_13650);
nor U17435 (N_17435,N_12857,N_14425);
xnor U17436 (N_17436,N_13701,N_12881);
xor U17437 (N_17437,N_13568,N_13220);
nor U17438 (N_17438,N_14396,N_14430);
and U17439 (N_17439,N_14911,N_14370);
nand U17440 (N_17440,N_13533,N_14461);
and U17441 (N_17441,N_13479,N_14008);
nand U17442 (N_17442,N_13450,N_13329);
and U17443 (N_17443,N_13220,N_12807);
and U17444 (N_17444,N_14521,N_12778);
nor U17445 (N_17445,N_13290,N_14532);
xor U17446 (N_17446,N_12722,N_14265);
or U17447 (N_17447,N_13528,N_13709);
and U17448 (N_17448,N_13932,N_14053);
or U17449 (N_17449,N_12798,N_14785);
xor U17450 (N_17450,N_14085,N_13310);
nand U17451 (N_17451,N_13891,N_14321);
nand U17452 (N_17452,N_12951,N_14918);
or U17453 (N_17453,N_13242,N_14096);
and U17454 (N_17454,N_14492,N_13335);
nand U17455 (N_17455,N_14995,N_13131);
and U17456 (N_17456,N_12651,N_14964);
nand U17457 (N_17457,N_13413,N_12800);
xnor U17458 (N_17458,N_13219,N_12738);
and U17459 (N_17459,N_13681,N_13264);
nand U17460 (N_17460,N_13063,N_14073);
nor U17461 (N_17461,N_14360,N_14959);
xor U17462 (N_17462,N_14299,N_13472);
xor U17463 (N_17463,N_12698,N_14866);
nand U17464 (N_17464,N_12703,N_14182);
xor U17465 (N_17465,N_13096,N_12741);
and U17466 (N_17466,N_14445,N_13656);
nor U17467 (N_17467,N_13473,N_14526);
or U17468 (N_17468,N_14182,N_14061);
nand U17469 (N_17469,N_13660,N_14966);
xor U17470 (N_17470,N_14065,N_13407);
and U17471 (N_17471,N_14052,N_13588);
nand U17472 (N_17472,N_14437,N_13335);
nand U17473 (N_17473,N_12752,N_14370);
or U17474 (N_17474,N_14810,N_13577);
and U17475 (N_17475,N_14064,N_13957);
xnor U17476 (N_17476,N_13844,N_12946);
or U17477 (N_17477,N_14803,N_14096);
nor U17478 (N_17478,N_13923,N_14978);
nor U17479 (N_17479,N_14704,N_14614);
or U17480 (N_17480,N_12854,N_13824);
nor U17481 (N_17481,N_13714,N_12500);
xnor U17482 (N_17482,N_13667,N_14251);
nand U17483 (N_17483,N_13157,N_14769);
or U17484 (N_17484,N_14940,N_13311);
and U17485 (N_17485,N_14608,N_13193);
xnor U17486 (N_17486,N_14022,N_12787);
or U17487 (N_17487,N_13230,N_14884);
or U17488 (N_17488,N_14402,N_13131);
and U17489 (N_17489,N_12523,N_13730);
or U17490 (N_17490,N_12660,N_13846);
or U17491 (N_17491,N_14730,N_13923);
or U17492 (N_17492,N_14706,N_13589);
or U17493 (N_17493,N_12964,N_14916);
nand U17494 (N_17494,N_13103,N_12659);
nand U17495 (N_17495,N_12634,N_14438);
xnor U17496 (N_17496,N_13933,N_14179);
nand U17497 (N_17497,N_14355,N_12719);
and U17498 (N_17498,N_14120,N_14843);
and U17499 (N_17499,N_13444,N_13827);
and U17500 (N_17500,N_16388,N_16159);
nor U17501 (N_17501,N_16113,N_17334);
and U17502 (N_17502,N_16542,N_15466);
and U17503 (N_17503,N_16746,N_17389);
or U17504 (N_17504,N_15549,N_16861);
and U17505 (N_17505,N_15231,N_15311);
nor U17506 (N_17506,N_17396,N_16638);
nor U17507 (N_17507,N_15998,N_15279);
xnor U17508 (N_17508,N_16312,N_16817);
nor U17509 (N_17509,N_17265,N_15253);
xnor U17510 (N_17510,N_16731,N_17108);
xor U17511 (N_17511,N_17069,N_15724);
or U17512 (N_17512,N_17315,N_17331);
nor U17513 (N_17513,N_16412,N_15923);
xor U17514 (N_17514,N_16450,N_17249);
nor U17515 (N_17515,N_17161,N_15778);
or U17516 (N_17516,N_15458,N_16441);
xnor U17517 (N_17517,N_15869,N_16714);
nand U17518 (N_17518,N_15830,N_15432);
or U17519 (N_17519,N_16551,N_16271);
and U17520 (N_17520,N_15944,N_17267);
and U17521 (N_17521,N_17157,N_15340);
or U17522 (N_17522,N_16032,N_16037);
nand U17523 (N_17523,N_15089,N_15605);
xor U17524 (N_17524,N_15134,N_15767);
or U17525 (N_17525,N_16524,N_16813);
nor U17526 (N_17526,N_15158,N_15259);
nand U17527 (N_17527,N_15962,N_16428);
and U17528 (N_17528,N_15516,N_15706);
xnor U17529 (N_17529,N_15063,N_15071);
and U17530 (N_17530,N_15648,N_17190);
xnor U17531 (N_17531,N_15272,N_16512);
and U17532 (N_17532,N_15807,N_17077);
nand U17533 (N_17533,N_16415,N_15856);
or U17534 (N_17534,N_16235,N_15121);
nand U17535 (N_17535,N_16144,N_17232);
nor U17536 (N_17536,N_15787,N_15203);
nor U17537 (N_17537,N_15591,N_16123);
xnor U17538 (N_17538,N_16955,N_16099);
xor U17539 (N_17539,N_16836,N_15192);
nand U17540 (N_17540,N_16419,N_16452);
and U17541 (N_17541,N_16921,N_15556);
xnor U17542 (N_17542,N_17115,N_15984);
and U17543 (N_17543,N_15740,N_17212);
nand U17544 (N_17544,N_16730,N_17063);
nor U17545 (N_17545,N_16248,N_15244);
xnor U17546 (N_17546,N_16100,N_15911);
and U17547 (N_17547,N_15209,N_15603);
nand U17548 (N_17548,N_16522,N_16360);
xnor U17549 (N_17549,N_15166,N_17263);
nor U17550 (N_17550,N_15617,N_17305);
nor U17551 (N_17551,N_16487,N_15622);
nor U17552 (N_17552,N_16437,N_15714);
nor U17553 (N_17553,N_16831,N_15827);
or U17554 (N_17554,N_16027,N_15333);
nor U17555 (N_17555,N_15111,N_17025);
nand U17556 (N_17556,N_16536,N_16461);
and U17557 (N_17557,N_16637,N_15927);
xnor U17558 (N_17558,N_17120,N_15201);
or U17559 (N_17559,N_17449,N_17175);
nor U17560 (N_17560,N_17406,N_16757);
and U17561 (N_17561,N_16747,N_15660);
nor U17562 (N_17562,N_15468,N_15914);
xnor U17563 (N_17563,N_15996,N_16752);
and U17564 (N_17564,N_16048,N_16626);
nand U17565 (N_17565,N_16076,N_16790);
xnor U17566 (N_17566,N_16614,N_15225);
or U17567 (N_17567,N_17193,N_15540);
nand U17568 (N_17568,N_16784,N_17083);
xnor U17569 (N_17569,N_15674,N_15289);
nor U17570 (N_17570,N_15337,N_15888);
or U17571 (N_17571,N_15080,N_15286);
nor U17572 (N_17572,N_16007,N_15119);
or U17573 (N_17573,N_16985,N_15183);
nand U17574 (N_17574,N_15173,N_17008);
or U17575 (N_17575,N_16339,N_15214);
and U17576 (N_17576,N_15169,N_15490);
nor U17577 (N_17577,N_17413,N_15314);
or U17578 (N_17578,N_15033,N_16655);
nand U17579 (N_17579,N_17234,N_15439);
and U17580 (N_17580,N_15663,N_16502);
or U17581 (N_17581,N_17252,N_15159);
nor U17582 (N_17582,N_16464,N_17089);
nand U17583 (N_17583,N_15789,N_16509);
nor U17584 (N_17584,N_16837,N_16128);
and U17585 (N_17585,N_15186,N_17274);
nor U17586 (N_17586,N_17095,N_17210);
nand U17587 (N_17587,N_16386,N_15946);
or U17588 (N_17588,N_16550,N_16807);
xor U17589 (N_17589,N_16012,N_16268);
xnor U17590 (N_17590,N_16265,N_15784);
nor U17591 (N_17591,N_16797,N_15939);
or U17592 (N_17592,N_16936,N_16965);
nor U17593 (N_17593,N_17477,N_16523);
xnor U17594 (N_17594,N_15631,N_15360);
xor U17595 (N_17595,N_15430,N_16920);
or U17596 (N_17596,N_15810,N_15051);
and U17597 (N_17597,N_17457,N_15167);
xnor U17598 (N_17598,N_17088,N_15970);
or U17599 (N_17599,N_15049,N_15363);
nor U17600 (N_17600,N_15711,N_16325);
nor U17601 (N_17601,N_16625,N_16697);
xor U17602 (N_17602,N_16309,N_17241);
nor U17603 (N_17603,N_16947,N_15278);
and U17604 (N_17604,N_15822,N_16600);
nand U17605 (N_17605,N_17408,N_15087);
nor U17606 (N_17606,N_16178,N_17174);
xnor U17607 (N_17607,N_16821,N_15846);
xor U17608 (N_17608,N_15851,N_15950);
xnor U17609 (N_17609,N_15759,N_15954);
or U17610 (N_17610,N_16355,N_16618);
and U17611 (N_17611,N_16408,N_15068);
xor U17612 (N_17612,N_17012,N_16979);
xnor U17613 (N_17613,N_16779,N_17309);
or U17614 (N_17614,N_17159,N_16071);
nand U17615 (N_17615,N_15451,N_16414);
xor U17616 (N_17616,N_16062,N_16395);
xor U17617 (N_17617,N_16809,N_16933);
or U17618 (N_17618,N_15669,N_15862);
or U17619 (N_17619,N_15814,N_15334);
nand U17620 (N_17620,N_16483,N_15771);
nand U17621 (N_17621,N_15366,N_17437);
nor U17622 (N_17622,N_16818,N_15568);
nand U17623 (N_17623,N_15084,N_17224);
xnor U17624 (N_17624,N_16025,N_15569);
nand U17625 (N_17625,N_15864,N_15424);
nand U17626 (N_17626,N_16376,N_16081);
or U17627 (N_17627,N_16950,N_15586);
xor U17628 (N_17628,N_17288,N_15057);
nand U17629 (N_17629,N_16663,N_16230);
nand U17630 (N_17630,N_15264,N_16763);
xor U17631 (N_17631,N_16303,N_15566);
nand U17632 (N_17632,N_17171,N_16195);
and U17633 (N_17633,N_16152,N_15298);
nand U17634 (N_17634,N_16801,N_16406);
xor U17635 (N_17635,N_17273,N_16892);
or U17636 (N_17636,N_16923,N_16770);
and U17637 (N_17637,N_16753,N_16744);
xor U17638 (N_17638,N_16343,N_17280);
or U17639 (N_17639,N_16451,N_15309);
xnor U17640 (N_17640,N_17292,N_17495);
nand U17641 (N_17641,N_15526,N_17092);
xnor U17642 (N_17642,N_16657,N_16151);
and U17643 (N_17643,N_15730,N_16847);
nor U17644 (N_17644,N_15429,N_15734);
xnor U17645 (N_17645,N_17164,N_16165);
nand U17646 (N_17646,N_15890,N_16276);
and U17647 (N_17647,N_15844,N_15092);
or U17648 (N_17648,N_15975,N_15554);
or U17649 (N_17649,N_15103,N_16702);
xor U17650 (N_17650,N_15721,N_16926);
nor U17651 (N_17651,N_17336,N_16842);
nand U17652 (N_17652,N_15713,N_15908);
nand U17653 (N_17653,N_16330,N_15551);
and U17654 (N_17654,N_16989,N_16260);
and U17655 (N_17655,N_17016,N_16768);
or U17656 (N_17656,N_15038,N_17376);
xnor U17657 (N_17657,N_16850,N_16196);
nand U17658 (N_17658,N_17483,N_15339);
nand U17659 (N_17659,N_15728,N_15130);
and U17660 (N_17660,N_15023,N_15933);
and U17661 (N_17661,N_15661,N_15606);
nand U17662 (N_17662,N_15188,N_15623);
xor U17663 (N_17663,N_16552,N_15376);
nor U17664 (N_17664,N_15821,N_15543);
nor U17665 (N_17665,N_15427,N_17319);
nand U17666 (N_17666,N_16410,N_17229);
nand U17667 (N_17667,N_16953,N_16934);
and U17668 (N_17668,N_15346,N_17145);
nand U17669 (N_17669,N_16392,N_16829);
xnor U17670 (N_17670,N_17140,N_15709);
nor U17671 (N_17671,N_17386,N_17259);
xnor U17672 (N_17672,N_17146,N_15578);
nor U17673 (N_17673,N_17141,N_15604);
and U17674 (N_17674,N_16290,N_17354);
xnor U17675 (N_17675,N_16073,N_17096);
xor U17676 (N_17676,N_16453,N_17478);
nor U17677 (N_17677,N_16578,N_17378);
and U17678 (N_17678,N_17446,N_15054);
nand U17679 (N_17679,N_17377,N_15283);
nor U17680 (N_17680,N_15282,N_17260);
or U17681 (N_17681,N_15003,N_15234);
nor U17682 (N_17682,N_15380,N_16438);
xnor U17683 (N_17683,N_16009,N_16036);
or U17684 (N_17684,N_15401,N_15959);
xnor U17685 (N_17685,N_16992,N_17294);
or U17686 (N_17686,N_15547,N_17430);
and U17687 (N_17687,N_15668,N_17411);
and U17688 (N_17688,N_15153,N_15753);
and U17689 (N_17689,N_15936,N_15992);
nor U17690 (N_17690,N_16340,N_16186);
xor U17691 (N_17691,N_15287,N_16171);
nor U17692 (N_17692,N_15383,N_15079);
xor U17693 (N_17693,N_15041,N_17407);
and U17694 (N_17694,N_15291,N_15277);
xnor U17695 (N_17695,N_16583,N_15562);
and U17696 (N_17696,N_16952,N_16532);
or U17697 (N_17697,N_16116,N_16828);
and U17698 (N_17698,N_16751,N_15780);
nor U17699 (N_17699,N_15132,N_15027);
xor U17700 (N_17700,N_16131,N_17189);
or U17701 (N_17701,N_15416,N_15075);
xnor U17702 (N_17702,N_15237,N_15756);
nor U17703 (N_17703,N_16232,N_16013);
xnor U17704 (N_17704,N_17176,N_16734);
xor U17705 (N_17705,N_15021,N_16822);
xor U17706 (N_17706,N_17126,N_16855);
nor U17707 (N_17707,N_16624,N_16398);
or U17708 (N_17708,N_16580,N_17087);
xnor U17709 (N_17709,N_15464,N_15522);
nor U17710 (N_17710,N_15945,N_17417);
xor U17711 (N_17711,N_15369,N_16463);
or U17712 (N_17712,N_15269,N_15300);
or U17713 (N_17713,N_16460,N_15115);
and U17714 (N_17714,N_15098,N_15645);
and U17715 (N_17715,N_15681,N_16827);
nor U17716 (N_17716,N_17065,N_16028);
nor U17717 (N_17717,N_16879,N_17187);
or U17718 (N_17718,N_15013,N_15723);
nand U17719 (N_17719,N_17492,N_16537);
or U17720 (N_17720,N_15917,N_15546);
or U17721 (N_17721,N_17110,N_16603);
nand U17722 (N_17722,N_16189,N_16244);
nand U17723 (N_17723,N_16191,N_16192);
nand U17724 (N_17724,N_15243,N_15726);
xnor U17725 (N_17725,N_15088,N_15099);
nor U17726 (N_17726,N_15128,N_16280);
or U17727 (N_17727,N_16002,N_15637);
or U17728 (N_17728,N_15976,N_15123);
xnor U17729 (N_17729,N_15431,N_15826);
xor U17730 (N_17730,N_17455,N_15532);
and U17731 (N_17731,N_16504,N_16860);
xnor U17732 (N_17732,N_15179,N_15215);
xnor U17733 (N_17733,N_15375,N_16440);
nand U17734 (N_17734,N_16984,N_15585);
xnor U17735 (N_17735,N_15861,N_16959);
xor U17736 (N_17736,N_15731,N_16117);
and U17737 (N_17737,N_15472,N_15988);
nor U17738 (N_17738,N_16940,N_16517);
xor U17739 (N_17739,N_17316,N_15628);
xor U17740 (N_17740,N_15572,N_17209);
nand U17741 (N_17741,N_16620,N_15797);
nand U17742 (N_17742,N_17067,N_16489);
nand U17743 (N_17743,N_15402,N_15717);
nor U17744 (N_17744,N_17447,N_16704);
and U17745 (N_17745,N_16685,N_16238);
and U17746 (N_17746,N_16038,N_16665);
nand U17747 (N_17747,N_16293,N_16890);
xnor U17748 (N_17748,N_16794,N_16957);
and U17749 (N_17749,N_16050,N_17036);
xor U17750 (N_17750,N_17081,N_17296);
nor U17751 (N_17751,N_15811,N_16215);
nand U17752 (N_17752,N_17277,N_15001);
xnor U17753 (N_17753,N_15804,N_15884);
or U17754 (N_17754,N_17424,N_15649);
xnor U17755 (N_17755,N_16511,N_15514);
nor U17756 (N_17756,N_17445,N_17398);
xnor U17757 (N_17757,N_16590,N_16249);
nand U17758 (N_17758,N_17432,N_17144);
and U17759 (N_17759,N_15155,N_15813);
and U17760 (N_17760,N_15794,N_15320);
nor U17761 (N_17761,N_15657,N_15961);
and U17762 (N_17762,N_15398,N_16815);
nor U17763 (N_17763,N_15228,N_17061);
nor U17764 (N_17764,N_16404,N_15437);
xor U17765 (N_17765,N_17243,N_16733);
nor U17766 (N_17766,N_16352,N_16227);
nand U17767 (N_17767,N_16683,N_15897);
or U17768 (N_17768,N_17481,N_16703);
nand U17769 (N_17769,N_17372,N_15284);
and U17770 (N_17770,N_15775,N_17245);
nor U17771 (N_17771,N_15446,N_16659);
xor U17772 (N_17772,N_15510,N_17484);
nor U17773 (N_17773,N_16986,N_16061);
xor U17774 (N_17774,N_16334,N_16868);
nand U17775 (N_17775,N_15639,N_16241);
nand U17776 (N_17776,N_15790,N_16636);
or U17777 (N_17777,N_15651,N_16572);
or U17778 (N_17778,N_16980,N_17248);
xor U17779 (N_17779,N_16592,N_16931);
xnor U17780 (N_17780,N_17099,N_17181);
xor U17781 (N_17781,N_16805,N_15247);
or U17782 (N_17782,N_15149,N_16876);
or U17783 (N_17783,N_16997,N_16493);
nor U17784 (N_17784,N_15871,N_16221);
xnor U17785 (N_17785,N_15671,N_16236);
nor U17786 (N_17786,N_16634,N_15619);
and U17787 (N_17787,N_17320,N_17299);
xor U17788 (N_17788,N_16998,N_15381);
nor U17789 (N_17789,N_16778,N_15608);
and U17790 (N_17790,N_17019,N_16561);
xnor U17791 (N_17791,N_17251,N_16254);
or U17792 (N_17792,N_17042,N_16381);
or U17793 (N_17793,N_15394,N_16729);
xor U17794 (N_17794,N_17058,N_16833);
nand U17795 (N_17795,N_15860,N_15417);
xor U17796 (N_17796,N_15438,N_16839);
nor U17797 (N_17797,N_15456,N_15067);
xor U17798 (N_17798,N_15716,N_16394);
xnor U17799 (N_17799,N_16399,N_17106);
nand U17800 (N_17800,N_17236,N_16172);
xnor U17801 (N_17801,N_15007,N_17202);
xor U17802 (N_17802,N_15015,N_15399);
nor U17803 (N_17803,N_15876,N_17031);
xor U17804 (N_17804,N_16677,N_15781);
and U17805 (N_17805,N_17488,N_16206);
or U17806 (N_17806,N_16396,N_15110);
or U17807 (N_17807,N_15178,N_17426);
nand U17808 (N_17808,N_16385,N_16246);
and U17809 (N_17809,N_16889,N_17246);
or U17810 (N_17810,N_16316,N_16362);
nand U17811 (N_17811,N_15539,N_17383);
or U17812 (N_17812,N_15990,N_17491);
and U17813 (N_17813,N_16516,N_16713);
or U17814 (N_17814,N_16257,N_15070);
or U17815 (N_17815,N_16401,N_15521);
nand U17816 (N_17816,N_16258,N_17313);
or U17817 (N_17817,N_15900,N_15332);
nor U17818 (N_17818,N_15364,N_16780);
xor U17819 (N_17819,N_15792,N_16764);
and U17820 (N_17820,N_15689,N_15727);
nand U17821 (N_17821,N_16595,N_15701);
xnor U17822 (N_17822,N_16198,N_15498);
nor U17823 (N_17823,N_16628,N_16084);
or U17824 (N_17824,N_15501,N_17184);
xor U17825 (N_17825,N_16885,N_15273);
nor U17826 (N_17826,N_17431,N_15989);
or U17827 (N_17827,N_17498,N_17211);
xor U17828 (N_17828,N_15517,N_16143);
or U17829 (N_17829,N_17205,N_16505);
nand U17830 (N_17830,N_17356,N_15573);
xnor U17831 (N_17831,N_15370,N_16905);
or U17832 (N_17832,N_16792,N_16650);
and U17833 (N_17833,N_17338,N_16211);
nor U17834 (N_17834,N_15545,N_16164);
xor U17835 (N_17835,N_17074,N_16534);
nor U17836 (N_17836,N_16444,N_16941);
nor U17837 (N_17837,N_15223,N_17045);
or U17838 (N_17838,N_16439,N_15597);
or U17839 (N_17839,N_16413,N_16278);
nor U17840 (N_17840,N_15896,N_16297);
or U17841 (N_17841,N_16688,N_15489);
and U17842 (N_17842,N_17476,N_16006);
or U17843 (N_17843,N_17297,N_16642);
and U17844 (N_17844,N_17068,N_15834);
nor U17845 (N_17845,N_16272,N_17361);
nand U17846 (N_17846,N_15020,N_16604);
or U17847 (N_17847,N_16155,N_15146);
and U17848 (N_17848,N_16181,N_16288);
xor U17849 (N_17849,N_17225,N_17400);
and U17850 (N_17850,N_16707,N_15331);
xor U17851 (N_17851,N_16194,N_15675);
and U17852 (N_17852,N_17073,N_16649);
or U17853 (N_17853,N_17179,N_16798);
nand U17854 (N_17854,N_16750,N_16000);
xnor U17855 (N_17855,N_16838,N_15969);
nand U17856 (N_17856,N_17071,N_15365);
nor U17857 (N_17857,N_17213,N_16954);
nor U17858 (N_17858,N_17156,N_16470);
nand U17859 (N_17859,N_16939,N_15191);
or U17860 (N_17860,N_15351,N_17394);
nand U17861 (N_17861,N_16893,N_16569);
xnor U17862 (N_17862,N_16462,N_17250);
xor U17863 (N_17863,N_17103,N_16443);
or U17864 (N_17864,N_16993,N_17183);
xnor U17865 (N_17865,N_16270,N_16044);
xor U17866 (N_17866,N_16031,N_15926);
xor U17867 (N_17867,N_16158,N_17423);
nor U17868 (N_17868,N_16422,N_15301);
nor U17869 (N_17869,N_17185,N_17276);
nand U17870 (N_17870,N_15891,N_16234);
and U17871 (N_17871,N_16156,N_15285);
or U17872 (N_17872,N_17167,N_15393);
xnor U17873 (N_17873,N_16996,N_16157);
nand U17874 (N_17874,N_15017,N_16279);
xor U17875 (N_17875,N_15587,N_15403);
nor U17876 (N_17876,N_17059,N_15863);
nand U17877 (N_17877,N_16387,N_16601);
nand U17878 (N_17878,N_16937,N_15066);
and U17879 (N_17879,N_15583,N_16786);
xor U17880 (N_17880,N_17456,N_15786);
xor U17881 (N_17881,N_16486,N_15904);
and U17882 (N_17882,N_15815,N_16354);
nor U17883 (N_17883,N_15582,N_15133);
nand U17884 (N_17884,N_17218,N_16035);
xor U17885 (N_17885,N_16029,N_15343);
xnor U17886 (N_17886,N_16812,N_17169);
xnor U17887 (N_17887,N_16264,N_15632);
or U17888 (N_17888,N_15518,N_15419);
or U17889 (N_17889,N_16286,N_16070);
or U17890 (N_17890,N_17295,N_15903);
and U17891 (N_17891,N_16901,N_16929);
nor U17892 (N_17892,N_17392,N_16558);
and U17893 (N_17893,N_16023,N_16327);
xnor U17894 (N_17894,N_16379,N_17186);
xor U17895 (N_17895,N_15349,N_16140);
xnor U17896 (N_17896,N_15595,N_16742);
and U17897 (N_17897,N_17034,N_16501);
nor U17898 (N_17898,N_15305,N_17390);
or U17899 (N_17899,N_17101,N_17370);
or U17900 (N_17900,N_17454,N_15208);
or U17901 (N_17901,N_16393,N_16546);
or U17902 (N_17902,N_16175,N_17384);
xor U17903 (N_17903,N_16758,N_15469);
and U17904 (N_17904,N_17147,N_17015);
nor U17905 (N_17905,N_17364,N_16120);
nand U17906 (N_17906,N_16067,N_16844);
nand U17907 (N_17907,N_16247,N_17009);
nor U17908 (N_17908,N_15249,N_15922);
nor U17909 (N_17909,N_17151,N_15136);
nor U17910 (N_17910,N_15306,N_15216);
xor U17911 (N_17911,N_15801,N_16689);
or U17912 (N_17912,N_15313,N_16425);
nor U17913 (N_17913,N_15042,N_16447);
or U17914 (N_17914,N_16220,N_15576);
nor U17915 (N_17915,N_15162,N_16167);
or U17916 (N_17916,N_16748,N_15101);
nand U17917 (N_17917,N_16307,N_17349);
xor U17918 (N_17918,N_15991,N_15492);
nand U17919 (N_17919,N_16964,N_16826);
xor U17920 (N_17920,N_15915,N_15388);
or U17921 (N_17921,N_15838,N_15978);
xor U17922 (N_17922,N_15602,N_16956);
or U17923 (N_17923,N_15808,N_16019);
nor U17924 (N_17924,N_15118,N_15327);
nor U17925 (N_17925,N_17123,N_16491);
nand U17926 (N_17926,N_16174,N_15009);
nand U17927 (N_17927,N_17168,N_15122);
and U17928 (N_17928,N_15615,N_15072);
xor U17929 (N_17929,N_16324,N_16124);
or U17930 (N_17930,N_17441,N_17165);
nor U17931 (N_17931,N_15144,N_15621);
and U17932 (N_17932,N_17271,N_15672);
xor U17933 (N_17933,N_17049,N_16130);
xor U17934 (N_17934,N_16856,N_15691);
xnor U17935 (N_17935,N_17075,N_17435);
nand U17936 (N_17936,N_15044,N_17052);
or U17937 (N_17937,N_16899,N_15507);
nor U17938 (N_17938,N_16357,N_17359);
or U17939 (N_17939,N_15584,N_16800);
nand U17940 (N_17940,N_16498,N_15131);
nand U17941 (N_17941,N_15267,N_16699);
nor U17942 (N_17942,N_15718,N_16865);
and U17943 (N_17943,N_17010,N_16864);
or U17944 (N_17944,N_15461,N_16342);
nand U17945 (N_17945,N_16176,N_15872);
or U17946 (N_17946,N_15949,N_16661);
nand U17947 (N_17947,N_15444,N_17300);
nand U17948 (N_17948,N_15528,N_16336);
or U17949 (N_17949,N_16743,N_15426);
and U17950 (N_17950,N_15534,N_17197);
nand U17951 (N_17951,N_15737,N_15770);
nor U17952 (N_17952,N_15414,N_16571);
xor U17953 (N_17953,N_15357,N_15952);
nand U17954 (N_17954,N_17467,N_16958);
and U17955 (N_17955,N_16991,N_17287);
xor U17956 (N_17956,N_16497,N_17029);
nor U17957 (N_17957,N_15077,N_16562);
xor U17958 (N_17958,N_15246,N_15942);
xnor U17959 (N_17959,N_15825,N_16673);
xnor U17960 (N_17960,N_17093,N_15238);
xor U17961 (N_17961,N_16466,N_17440);
and U17962 (N_17962,N_17085,N_15299);
xor U17963 (N_17963,N_15703,N_15448);
xor U17964 (N_17964,N_16251,N_15344);
and U17965 (N_17965,N_15853,N_17474);
or U17966 (N_17966,N_15684,N_17422);
or U17967 (N_17967,N_15390,N_15048);
nand U17968 (N_17968,N_16233,N_16052);
nor U17969 (N_17969,N_15116,N_16651);
xnor U17970 (N_17970,N_16640,N_15405);
or U17971 (N_17971,N_17125,N_17399);
xor U17972 (N_17972,N_15442,N_16331);
xor U17973 (N_17973,N_17013,N_15046);
and U17974 (N_17974,N_17040,N_16101);
or U17975 (N_17975,N_16848,N_15065);
and U17976 (N_17976,N_15537,N_15090);
nand U17977 (N_17977,N_17337,N_17253);
nor U17978 (N_17978,N_16135,N_15739);
or U17979 (N_17979,N_15694,N_15980);
nand U17980 (N_17980,N_16496,N_15204);
nor U17981 (N_17981,N_16318,N_15335);
nor U17982 (N_17982,N_16712,N_16843);
and U17983 (N_17983,N_16863,N_16105);
xnor U17984 (N_17984,N_16472,N_16180);
and U17985 (N_17985,N_15873,N_17262);
nor U17986 (N_17986,N_17054,N_17293);
or U17987 (N_17987,N_17072,N_16402);
nor U17988 (N_17988,N_16887,N_15124);
xnor U17989 (N_17989,N_15142,N_15019);
nor U17990 (N_17990,N_16667,N_16459);
nand U17991 (N_17991,N_15047,N_15704);
or U17992 (N_17992,N_16647,N_15934);
and U17993 (N_17993,N_15485,N_15145);
and U17994 (N_17994,N_15550,N_15773);
xor U17995 (N_17995,N_16298,N_16349);
or U17996 (N_17996,N_15290,N_16631);
or U17997 (N_17997,N_15607,N_15195);
xor U17998 (N_17998,N_15184,N_17358);
nand U17999 (N_17999,N_15774,N_16344);
nor U18000 (N_18000,N_15056,N_16633);
and U18001 (N_18001,N_17290,N_17256);
and U18002 (N_18002,N_16884,N_15303);
nand U18003 (N_18003,N_15212,N_16602);
or U18004 (N_18004,N_15034,N_17163);
xor U18005 (N_18005,N_16654,N_15754);
and U18006 (N_18006,N_15800,N_16894);
xor U18007 (N_18007,N_16161,N_15471);
nor U18008 (N_18008,N_15761,N_16597);
and U18009 (N_18009,N_15752,N_17155);
or U18010 (N_18010,N_17330,N_16974);
or U18011 (N_18011,N_15886,N_15744);
nand U18012 (N_18012,N_16341,N_15107);
nand U18013 (N_18013,N_16229,N_15168);
xor U18014 (N_18014,N_15028,N_15598);
or U18015 (N_18015,N_15920,N_15941);
or U18016 (N_18016,N_15475,N_16529);
and U18017 (N_18017,N_16075,N_16908);
or U18018 (N_18018,N_15652,N_16585);
nand U18019 (N_18019,N_16675,N_15638);
xor U18020 (N_18020,N_17237,N_15820);
and U18021 (N_18021,N_16237,N_15725);
or U18022 (N_18022,N_17343,N_16698);
nor U18023 (N_18023,N_15229,N_16645);
xnor U18024 (N_18024,N_15227,N_17475);
xnor U18025 (N_18025,N_15220,N_17434);
nor U18026 (N_18026,N_16201,N_15478);
or U18027 (N_18027,N_16914,N_16262);
xnor U18028 (N_18028,N_16648,N_16193);
and U18029 (N_18029,N_16304,N_15367);
and U18030 (N_18030,N_17128,N_15170);
xnor U18031 (N_18031,N_16912,N_15929);
nor U18032 (N_18032,N_16611,N_17291);
or U18033 (N_18033,N_16359,N_15533);
and U18034 (N_18034,N_16059,N_15338);
and U18035 (N_18035,N_15252,N_16994);
nor U18036 (N_18036,N_17001,N_16092);
or U18037 (N_18037,N_16811,N_15326);
and U18038 (N_18038,N_16560,N_15552);
nand U18039 (N_18039,N_15610,N_16300);
or U18040 (N_18040,N_16427,N_16066);
or U18041 (N_18041,N_15481,N_17464);
nand U18042 (N_18042,N_15487,N_15879);
nor U18043 (N_18043,N_16609,N_16126);
nor U18044 (N_18044,N_15509,N_16981);
nor U18045 (N_18045,N_15798,N_17166);
nor U18046 (N_18046,N_15329,N_15791);
and U18047 (N_18047,N_16185,N_16820);
nand U18048 (N_18048,N_16096,N_16458);
or U18049 (N_18049,N_16449,N_15086);
xor U18050 (N_18050,N_15199,N_16115);
and U18051 (N_18051,N_16374,N_16353);
nand U18052 (N_18052,N_15654,N_17460);
nor U18053 (N_18053,N_15589,N_16197);
nand U18054 (N_18054,N_17097,N_15708);
and U18055 (N_18055,N_16643,N_15483);
xor U18056 (N_18056,N_16814,N_15643);
xnor U18057 (N_18057,N_15105,N_16549);
xor U18058 (N_18058,N_15600,N_15973);
xor U18059 (N_18059,N_16356,N_16188);
xor U18060 (N_18060,N_16055,N_15176);
and U18061 (N_18061,N_15868,N_16499);
nand U18062 (N_18062,N_16781,N_16928);
and U18063 (N_18063,N_17057,N_16736);
nand U18064 (N_18064,N_15043,N_16245);
nor U18065 (N_18065,N_16103,N_16579);
nor U18066 (N_18066,N_17180,N_15935);
and U18067 (N_18067,N_16533,N_15785);
and U18068 (N_18068,N_16617,N_17381);
xnor U18069 (N_18069,N_16426,N_17289);
or U18070 (N_18070,N_15889,N_15924);
or U18071 (N_18071,N_16433,N_15143);
and U18072 (N_18072,N_15907,N_16320);
nand U18073 (N_18073,N_16005,N_15508);
or U18074 (N_18074,N_17321,N_16380);
nand U18075 (N_18075,N_17342,N_15180);
xnor U18076 (N_18076,N_17062,N_15010);
or U18077 (N_18077,N_16397,N_17385);
or U18078 (N_18078,N_16846,N_16544);
nand U18079 (N_18079,N_17149,N_16106);
and U18080 (N_18080,N_16769,N_15665);
nor U18081 (N_18081,N_16995,N_16141);
nor U18082 (N_18082,N_15139,N_17127);
nand U18083 (N_18083,N_16282,N_15196);
and U18084 (N_18084,N_16531,N_15211);
and U18085 (N_18085,N_15397,N_16599);
nor U18086 (N_18086,N_17285,N_17172);
xor U18087 (N_18087,N_16816,N_15722);
or U18088 (N_18088,N_17286,N_17402);
or U18089 (N_18089,N_16228,N_16373);
and U18090 (N_18090,N_15022,N_15477);
or U18091 (N_18091,N_17192,N_16796);
nor U18092 (N_18092,N_16719,N_15408);
and U18093 (N_18093,N_15467,N_15126);
and U18094 (N_18094,N_16840,N_15000);
and U18095 (N_18095,N_15995,N_16003);
xor U18096 (N_18096,N_16915,N_15656);
xor U18097 (N_18097,N_15404,N_16299);
and U18098 (N_18098,N_15542,N_16913);
and U18099 (N_18099,N_15330,N_15641);
nand U18100 (N_18100,N_16598,N_15336);
or U18101 (N_18101,N_17233,N_15696);
nor U18102 (N_18102,N_16372,N_17450);
xnor U18103 (N_18103,N_16375,N_17160);
and U18104 (N_18104,N_15497,N_16976);
nor U18105 (N_18105,N_15324,N_15407);
xnor U18106 (N_18106,N_17046,N_17047);
nand U18107 (N_18107,N_15384,N_17382);
nand U18108 (N_18108,N_16163,N_15050);
nor U18109 (N_18109,N_17223,N_16682);
or U18110 (N_18110,N_17324,N_16348);
nor U18111 (N_18111,N_15193,N_15640);
and U18112 (N_18112,N_16990,N_15200);
or U18113 (N_18113,N_16623,N_15899);
and U18114 (N_18114,N_15979,N_17347);
xor U18115 (N_18115,N_16097,N_15630);
nor U18116 (N_18116,N_16726,N_16338);
or U18117 (N_18117,N_17222,N_16506);
nor U18118 (N_18118,N_15560,N_16705);
nor U18119 (N_18119,N_15006,N_16001);
or U18120 (N_18120,N_16776,N_17242);
or U18121 (N_18121,N_15997,N_16240);
nor U18122 (N_18122,N_17269,N_16431);
xnor U18123 (N_18123,N_16527,N_15910);
nand U18124 (N_18124,N_15150,N_17451);
nand U18125 (N_18125,N_15292,N_15108);
xor U18126 (N_18126,N_15316,N_16434);
and U18127 (N_18127,N_15499,N_17462);
nand U18128 (N_18128,N_15294,N_16468);
or U18129 (N_18129,N_16557,N_15504);
and U18130 (N_18130,N_17107,N_17486);
and U18131 (N_18131,N_17111,N_16170);
xnor U18132 (N_18132,N_16063,N_15096);
nor U18133 (N_18133,N_17082,N_15677);
nor U18134 (N_18134,N_17104,N_16513);
or U18135 (N_18135,N_17133,N_15266);
xnor U18136 (N_18136,N_16277,N_15174);
nand U18137 (N_18137,N_16693,N_15008);
nor U18138 (N_18138,N_16306,N_15636);
or U18139 (N_18139,N_15601,N_15986);
nor U18140 (N_18140,N_17231,N_15081);
or U18141 (N_18141,N_16745,N_16891);
or U18142 (N_18142,N_15463,N_15745);
and U18143 (N_18143,N_15841,N_15769);
xnor U18144 (N_18144,N_16700,N_15304);
nand U18145 (N_18145,N_16266,N_16060);
and U18146 (N_18146,N_15913,N_17134);
nand U18147 (N_18147,N_16480,N_16718);
xor U18148 (N_18148,N_15114,N_15420);
xnor U18149 (N_18149,N_17469,N_17357);
or U18150 (N_18150,N_15928,N_17170);
or U18151 (N_18151,N_16573,N_15473);
and U18152 (N_18152,N_15957,N_17033);
and U18153 (N_18153,N_15406,N_16823);
and U18154 (N_18154,N_15902,N_16424);
or U18155 (N_18155,N_15493,N_16043);
and U18156 (N_18156,N_17458,N_17135);
and U18157 (N_18157,N_17219,N_15189);
and U18158 (N_18158,N_15315,N_16610);
nand U18159 (N_18159,N_17139,N_16948);
nand U18160 (N_18160,N_16724,N_16346);
nor U18161 (N_18161,N_15818,N_16026);
or U18162 (N_18162,N_17105,N_17270);
nand U18163 (N_18163,N_16202,N_15308);
xnor U18164 (N_18164,N_17203,N_15987);
nand U18165 (N_18165,N_15226,N_16350);
xnor U18166 (N_18166,N_16361,N_15037);
or U18167 (N_18167,N_15977,N_15919);
nor U18168 (N_18168,N_16390,N_17079);
nand U18169 (N_18169,N_16612,N_16938);
nor U18170 (N_18170,N_15317,N_16455);
or U18171 (N_18171,N_17112,N_16972);
xnor U18172 (N_18172,N_15207,N_17283);
and U18173 (N_18173,N_15854,N_15658);
nor U18174 (N_18174,N_16129,N_17078);
and U18175 (N_18175,N_16968,N_15956);
or U18176 (N_18176,N_16314,N_16479);
xnor U18177 (N_18177,N_15421,N_16109);
or U18178 (N_18178,N_17129,N_15755);
nand U18179 (N_18179,N_15750,N_15032);
or U18180 (N_18180,N_16973,N_17442);
and U18181 (N_18181,N_15719,N_17352);
nor U18182 (N_18182,N_15852,N_17162);
nand U18183 (N_18183,N_15881,N_17064);
xor U18184 (N_18184,N_15931,N_15647);
xor U18185 (N_18185,N_16051,N_15255);
or U18186 (N_18186,N_16436,N_16554);
xnor U18187 (N_18187,N_16409,N_16787);
xor U18188 (N_18188,N_16285,N_15930);
xor U18189 (N_18189,N_16619,N_16369);
and U18190 (N_18190,N_17208,N_16653);
and U18191 (N_18191,N_17226,N_16494);
nand U18192 (N_18192,N_16121,N_15161);
xnor U18193 (N_18193,N_16335,N_16679);
xor U18194 (N_18194,N_17038,N_15440);
nand U18195 (N_18195,N_15165,N_15036);
and U18196 (N_18196,N_16420,N_17275);
or U18197 (N_18197,N_16292,N_15297);
and U18198 (N_18198,N_17314,N_17403);
xnor U18199 (N_18199,N_15094,N_16319);
nand U18200 (N_18200,N_17055,N_16011);
nor U18201 (N_18201,N_16686,N_15422);
and U18202 (N_18202,N_16122,N_17326);
and U18203 (N_18203,N_15783,N_16715);
xnor U18204 (N_18204,N_15341,N_15635);
nor U18205 (N_18205,N_16252,N_15565);
nand U18206 (N_18206,N_15372,N_16738);
or U18207 (N_18207,N_17303,N_15757);
nor U18208 (N_18208,N_16421,N_17084);
nor U18209 (N_18209,N_17346,N_15548);
nor U18210 (N_18210,N_16717,N_15966);
xor U18211 (N_18211,N_15795,N_17340);
or U18212 (N_18212,N_15318,N_15793);
nand U18213 (N_18213,N_16605,N_17130);
or U18214 (N_18214,N_15396,N_16418);
xnor U18215 (N_18215,N_17306,N_17173);
and U18216 (N_18216,N_16187,N_16924);
and U18217 (N_18217,N_17217,N_16935);
and U18218 (N_18218,N_17247,N_15434);
or U18219 (N_18219,N_15348,N_16102);
xnor U18220 (N_18220,N_17216,N_16591);
nor U18221 (N_18221,N_15355,N_15806);
nand U18222 (N_18222,N_15251,N_15052);
and U18223 (N_18223,N_15127,N_16082);
or U18224 (N_18224,N_15395,N_15563);
or U18225 (N_18225,N_15222,N_16065);
and U18226 (N_18226,N_16795,N_15611);
and U18227 (N_18227,N_16875,N_16621);
or U18228 (N_18228,N_17221,N_16945);
nor U18229 (N_18229,N_15069,N_16883);
or U18230 (N_18230,N_15741,N_16485);
nand U18231 (N_18231,N_17136,N_17453);
xnor U18232 (N_18232,N_16173,N_16490);
nand U18233 (N_18233,N_16267,N_15570);
xnor U18234 (N_18234,N_16488,N_17416);
or U18235 (N_18235,N_15836,N_15480);
nor U18236 (N_18236,N_15371,N_16465);
nand U18237 (N_18237,N_15680,N_15894);
and U18238 (N_18238,N_16771,N_15310);
xor U18239 (N_18239,N_16112,N_15219);
and U18240 (N_18240,N_16365,N_15076);
nand U18241 (N_18241,N_15359,N_16004);
or U18242 (N_18242,N_15823,N_16377);
and U18243 (N_18243,N_16507,N_16056);
nand U18244 (N_18244,N_17070,N_16662);
nand U18245 (N_18245,N_17496,N_16918);
nand U18246 (N_18246,N_17206,N_16184);
nand U18247 (N_18247,N_15571,N_17182);
xor U18248 (N_18248,N_15425,N_16739);
or U18249 (N_18249,N_16095,N_15460);
xnor U18250 (N_18250,N_15932,N_15580);
nand U18251 (N_18251,N_15004,N_15379);
nor U18252 (N_18252,N_16323,N_15544);
and U18253 (N_18253,N_15218,N_16214);
and U18254 (N_18254,N_15002,N_16694);
nor U18255 (N_18255,N_16137,N_17215);
xnor U18256 (N_18256,N_16125,N_15024);
nand U18257 (N_18257,N_15525,N_16104);
nand U18258 (N_18258,N_16445,N_16204);
nand U18259 (N_18259,N_15221,N_15748);
xnor U18260 (N_18260,N_15590,N_15524);
or U18261 (N_18261,N_15882,N_17351);
nand U18262 (N_18262,N_16669,N_17004);
or U18263 (N_18263,N_17465,N_15307);
or U18264 (N_18264,N_15796,N_16806);
and U18265 (N_18265,N_16857,N_16589);
and U18266 (N_18266,N_16793,N_15985);
and U18267 (N_18267,N_16389,N_16302);
nor U18268 (N_18268,N_17195,N_17391);
nor U18269 (N_18269,N_15835,N_15151);
nand U18270 (N_18270,N_15644,N_15198);
nor U18271 (N_18271,N_16961,N_16224);
nand U18272 (N_18272,N_16039,N_16825);
or U18273 (N_18273,N_17348,N_17124);
nand U18274 (N_18274,N_16789,N_16146);
xor U18275 (N_18275,N_16111,N_15387);
nor U18276 (N_18276,N_16021,N_16089);
and U18277 (N_18277,N_17325,N_17368);
xor U18278 (N_18278,N_17405,N_16925);
or U18279 (N_18279,N_15867,N_16430);
and U18280 (N_18280,N_16017,N_15618);
nand U18281 (N_18281,N_16762,N_15257);
nor U18282 (N_18282,N_16761,N_17415);
and U18283 (N_18283,N_16457,N_15958);
xnor U18284 (N_18284,N_16832,N_17003);
nand U18285 (N_18285,N_17196,N_15523);
and U18286 (N_18286,N_15254,N_17086);
or U18287 (N_18287,N_16858,N_16741);
and U18288 (N_18288,N_16962,N_15236);
xnor U18289 (N_18289,N_16538,N_16723);
nand U18290 (N_18290,N_15536,N_15575);
and U18291 (N_18291,N_17345,N_15263);
xor U18292 (N_18292,N_15558,N_15682);
and U18293 (N_18293,N_16851,N_15058);
or U18294 (N_18294,N_15857,N_16970);
or U18295 (N_18295,N_16182,N_16966);
nor U18296 (N_18296,N_17037,N_15325);
nand U18297 (N_18297,N_17053,N_15520);
and U18298 (N_18298,N_17428,N_16727);
or U18299 (N_18299,N_15982,N_17002);
and U18300 (N_18300,N_15073,N_15901);
xor U18301 (N_18301,N_16584,N_15921);
and U18302 (N_18302,N_17191,N_16469);
xnor U18303 (N_18303,N_17118,N_17150);
and U18304 (N_18304,N_16596,N_15172);
xor U18305 (N_18305,N_16777,N_16337);
or U18306 (N_18306,N_16565,N_15655);
nor U18307 (N_18307,N_16949,N_15626);
xnor U18308 (N_18308,N_16930,N_16615);
nor U18309 (N_18309,N_16041,N_15206);
or U18310 (N_18310,N_15768,N_16008);
or U18311 (N_18311,N_15281,N_15673);
or U18312 (N_18312,N_15519,N_16256);
xnor U18313 (N_18313,N_17279,N_17393);
and U18314 (N_18314,N_15449,N_17367);
nand U18315 (N_18315,N_16830,N_15579);
nand U18316 (N_18316,N_16471,N_16416);
nand U18317 (N_18317,N_16367,N_15097);
nor U18318 (N_18318,N_15609,N_16364);
and U18319 (N_18319,N_16870,N_17482);
xnor U18320 (N_18320,N_16606,N_15061);
or U18321 (N_18321,N_17266,N_15612);
or U18322 (N_18322,N_17178,N_17032);
or U18323 (N_18323,N_17485,N_17235);
or U18324 (N_18324,N_15141,N_17201);
xnor U18325 (N_18325,N_16510,N_15574);
nor U18326 (N_18326,N_15382,N_16094);
nand U18327 (N_18327,N_17278,N_16684);
or U18328 (N_18328,N_16139,N_15553);
nand U18329 (N_18329,N_16110,N_17204);
xnor U18330 (N_18330,N_15345,N_15288);
nor U18331 (N_18331,N_15235,N_16681);
nor U18332 (N_18332,N_16514,N_16500);
nand U18333 (N_18333,N_17142,N_17420);
or U18334 (N_18334,N_15147,N_17494);
and U18335 (N_18335,N_15059,N_16326);
nor U18336 (N_18336,N_15599,N_15634);
xor U18337 (N_18337,N_15373,N_16058);
xor U18338 (N_18338,N_16911,N_15564);
nand U18339 (N_18339,N_15411,N_15577);
and U18340 (N_18340,N_17227,N_16190);
xor U18341 (N_18341,N_16835,N_16371);
and U18342 (N_18342,N_17353,N_15650);
nor U18343 (N_18343,N_15743,N_15848);
and U18344 (N_18344,N_15746,N_16305);
or U18345 (N_18345,N_16313,N_15486);
nor U18346 (N_18346,N_15697,N_16119);
nand U18347 (N_18347,N_17050,N_15840);
or U18348 (N_18348,N_15164,N_15060);
or U18349 (N_18349,N_17410,N_15210);
and U18350 (N_18350,N_16332,N_15156);
xor U18351 (N_18351,N_15940,N_15454);
or U18352 (N_18352,N_15265,N_15095);
nand U18353 (N_18353,N_15692,N_16301);
xor U18354 (N_18354,N_17060,N_16508);
xor U18355 (N_18355,N_15378,N_16239);
nand U18356 (N_18356,N_16243,N_15250);
and U18357 (N_18357,N_16896,N_15596);
and U18358 (N_18358,N_15715,N_15064);
and U18359 (N_18359,N_15453,N_16535);
nand U18360 (N_18360,N_15447,N_16088);
nor U18361 (N_18361,N_16015,N_16310);
and U18362 (N_18362,N_17264,N_16540);
or U18363 (N_18363,N_17090,N_17114);
or U18364 (N_18364,N_16725,N_16289);
nor U18365 (N_18365,N_15112,N_17281);
nor U18366 (N_18366,N_17094,N_16098);
or U18367 (N_18367,N_15455,N_16225);
xnor U18368 (N_18368,N_16695,N_16085);
or U18369 (N_18369,N_16200,N_15880);
nor U18370 (N_18370,N_16317,N_15465);
or U18371 (N_18371,N_15925,N_15014);
xnor U18372 (N_18372,N_15410,N_17312);
nand U18373 (N_18373,N_16072,N_15443);
nand U18374 (N_18374,N_15812,N_17024);
nand U18375 (N_18375,N_16093,N_16783);
or U18376 (N_18376,N_17199,N_15788);
and U18377 (N_18377,N_15906,N_16370);
and U18378 (N_18378,N_17244,N_17177);
nor U18379 (N_18379,N_15736,N_16287);
xor U18380 (N_18380,N_16975,N_16079);
and U18381 (N_18381,N_16563,N_16721);
and U18382 (N_18382,N_15968,N_15109);
or U18383 (N_18383,N_16217,N_15385);
and U18384 (N_18384,N_17339,N_15937);
nor U18385 (N_18385,N_17470,N_17298);
or U18386 (N_18386,N_15491,N_16519);
or U18387 (N_18387,N_15683,N_16904);
nor U18388 (N_18388,N_16575,N_17020);
nor U18389 (N_18389,N_16169,N_17048);
nor U18390 (N_18390,N_16086,N_16446);
and U18391 (N_18391,N_17459,N_15083);
nor U18392 (N_18392,N_16658,N_16919);
nor U18393 (N_18393,N_15620,N_15859);
nand U18394 (N_18394,N_15462,N_17200);
and U18395 (N_18395,N_16982,N_16692);
xnor U18396 (N_18396,N_15496,N_16147);
or U18397 (N_18397,N_16417,N_16261);
or U18398 (N_18398,N_16383,N_15005);
nor U18399 (N_18399,N_16859,N_15627);
xnor U18400 (N_18400,N_15883,N_16635);
and U18401 (N_18401,N_17327,N_15964);
or U18402 (N_18402,N_15678,N_17307);
and U18403 (N_18403,N_15135,N_16834);
or U18404 (N_18404,N_16142,N_15762);
or U18405 (N_18405,N_16588,N_15799);
xnor U18406 (N_18406,N_16114,N_15275);
xor U18407 (N_18407,N_16345,N_16068);
nand U18408 (N_18408,N_16576,N_16042);
or U18409 (N_18409,N_15817,N_17154);
nor U18410 (N_18410,N_17113,N_17006);
or U18411 (N_18411,N_17439,N_15738);
nor U18412 (N_18412,N_17117,N_17363);
nand U18413 (N_18413,N_15476,N_16090);
nand U18414 (N_18414,N_17018,N_15803);
and U18415 (N_18415,N_16138,N_15452);
nor U18416 (N_18416,N_16269,N_16582);
or U18417 (N_18417,N_16897,N_16046);
xor U18418 (N_18418,N_15106,N_15809);
or U18419 (N_18419,N_15031,N_15270);
or U18420 (N_18420,N_15555,N_15819);
and U18421 (N_18421,N_16378,N_15729);
and U18422 (N_18422,N_17395,N_16969);
and U18423 (N_18423,N_15892,N_16877);
xor U18424 (N_18424,N_16866,N_16322);
nor U18425 (N_18425,N_16646,N_16351);
xor U18426 (N_18426,N_17341,N_15233);
nand U18427 (N_18427,N_16521,N_16854);
xor U18428 (N_18428,N_16308,N_15177);
xor U18429 (N_18429,N_16802,N_17414);
and U18430 (N_18430,N_16951,N_17066);
or U18431 (N_18431,N_16907,N_15855);
nand U18432 (N_18432,N_15389,N_16932);
or U18433 (N_18433,N_15354,N_16363);
xnor U18434 (N_18434,N_16518,N_15513);
xnor U18435 (N_18435,N_17380,N_16545);
or U18436 (N_18436,N_17035,N_16477);
xnor U18437 (N_18437,N_15782,N_16690);
and U18438 (N_18438,N_16064,N_15011);
xor U18439 (N_18439,N_15506,N_17005);
xnor U18440 (N_18440,N_15163,N_17122);
or U18441 (N_18441,N_15874,N_15905);
nand U18442 (N_18442,N_16759,N_17433);
or U18443 (N_18443,N_16696,N_15831);
xor U18444 (N_18444,N_15592,N_15415);
xor U18445 (N_18445,N_16321,N_16680);
and U18446 (N_18446,N_15100,N_15039);
nand U18447 (N_18447,N_15895,N_16478);
and U18448 (N_18448,N_15642,N_15837);
xor U18449 (N_18449,N_15983,N_17369);
xor U18450 (N_18450,N_16391,N_15374);
or U18451 (N_18451,N_16149,N_16492);
nor U18452 (N_18452,N_17318,N_16607);
nand U18453 (N_18453,N_15423,N_16108);
or U18454 (N_18454,N_15720,N_16629);
xnor U18455 (N_18455,N_15776,N_15441);
nand U18456 (N_18456,N_16168,N_16212);
or U18457 (N_18457,N_16160,N_16503);
nand U18458 (N_18458,N_16382,N_17158);
and U18459 (N_18459,N_16701,N_16568);
or U18460 (N_18460,N_15450,N_15802);
xnor U18461 (N_18461,N_16691,N_16594);
xor U18462 (N_18462,N_17461,N_15625);
and U18463 (N_18463,N_16737,N_16040);
and U18464 (N_18464,N_17153,N_16944);
or U18465 (N_18465,N_15960,N_16018);
xor U18466 (N_18466,N_16862,N_15690);
nand U18467 (N_18467,N_16074,N_15847);
nor U18468 (N_18468,N_16153,N_15213);
or U18469 (N_18469,N_15845,N_16547);
nor U18470 (N_18470,N_15763,N_17007);
nand U18471 (N_18471,N_17419,N_16179);
and U18472 (N_18472,N_17429,N_15664);
xnor U18473 (N_18473,N_16788,N_17119);
nor U18474 (N_18474,N_16946,N_16710);
xnor U18475 (N_18475,N_15662,N_17387);
nor U18476 (N_18476,N_15353,N_16333);
nand U18477 (N_18477,N_16024,N_15241);
and U18478 (N_18478,N_16898,N_15040);
nor U18479 (N_18479,N_15505,N_15760);
nand U18480 (N_18480,N_17152,N_15700);
nand U18481 (N_18481,N_15160,N_16664);
xnor U18482 (N_18482,N_15772,N_15268);
xor U18483 (N_18483,N_16548,N_15120);
or U18484 (N_18484,N_16274,N_16528);
nand U18485 (N_18485,N_17043,N_15494);
nor U18486 (N_18486,N_17362,N_17056);
nand U18487 (N_18487,N_16671,N_16291);
and U18488 (N_18488,N_16735,N_16530);
nand U18489 (N_18489,N_15530,N_17023);
nand U18490 (N_18490,N_16740,N_16639);
nand U18491 (N_18491,N_15629,N_15953);
and U18492 (N_18492,N_16132,N_16872);
xnor U18493 (N_18493,N_16231,N_16539);
nor U18494 (N_18494,N_17466,N_16034);
and U18495 (N_18495,N_16627,N_17121);
xnor U18496 (N_18496,N_17268,N_16474);
nand U18497 (N_18497,N_16403,N_16886);
or U18498 (N_18498,N_17091,N_16049);
nor U18499 (N_18499,N_17418,N_15993);
and U18500 (N_18500,N_16641,N_15633);
and U18501 (N_18501,N_16294,N_17261);
nor U18502 (N_18502,N_16808,N_16559);
and U18503 (N_18503,N_16687,N_16283);
xnor U18504 (N_18504,N_16407,N_16987);
nand U18505 (N_18505,N_17328,N_15679);
nor U18506 (N_18506,N_15459,N_15016);
or U18507 (N_18507,N_17322,N_15676);
xor U18508 (N_18508,N_16902,N_16593);
nand U18509 (N_18509,N_16281,N_17444);
or U18510 (N_18510,N_16910,N_17332);
and U18511 (N_18511,N_15470,N_16022);
xor U18512 (N_18512,N_15274,N_15230);
nor U18513 (N_18513,N_16541,N_15280);
nor U18514 (N_18514,N_15239,N_16869);
or U18515 (N_18515,N_17468,N_16347);
xor U18516 (N_18516,N_16358,N_15436);
nor U18517 (N_18517,N_16054,N_15328);
or U18518 (N_18518,N_15764,N_16016);
xnor U18519 (N_18519,N_17448,N_17438);
and U18520 (N_18520,N_16775,N_15312);
xnor U18521 (N_18521,N_15302,N_16722);
and U18522 (N_18522,N_15839,N_17360);
and U18523 (N_18523,N_16118,N_15356);
nor U18524 (N_18524,N_16622,N_17022);
or U18525 (N_18525,N_15749,N_17302);
xnor U18526 (N_18526,N_15185,N_17350);
and U18527 (N_18527,N_15062,N_17230);
and U18528 (N_18528,N_15779,N_16136);
nand U18529 (N_18529,N_16916,N_17102);
and U18530 (N_18530,N_16328,N_16253);
nand U18531 (N_18531,N_15843,N_15347);
or U18532 (N_18532,N_16473,N_15154);
or U18533 (N_18533,N_17471,N_16525);
nor U18534 (N_18534,N_16162,N_16773);
xnor U18535 (N_18535,N_15698,N_16774);
xor U18536 (N_18536,N_16978,N_15742);
or U18537 (N_18537,N_16711,N_16967);
or U18538 (N_18538,N_16754,N_16014);
xnor U18539 (N_18539,N_15412,N_17284);
and U18540 (N_18540,N_16219,N_16145);
nor U18541 (N_18541,N_15951,N_16183);
xor U18542 (N_18542,N_15653,N_17489);
nand U18543 (N_18543,N_16922,N_17282);
and U18544 (N_18544,N_16177,N_15885);
nand U18545 (N_18545,N_16900,N_16960);
nor U18546 (N_18546,N_16942,N_16567);
nand U18547 (N_18547,N_16732,N_15194);
nand U18548 (N_18548,N_16845,N_15588);
xor U18549 (N_18549,N_17132,N_17452);
or U18550 (N_18550,N_17044,N_17311);
nand U18551 (N_18551,N_16429,N_17472);
xnor U18552 (N_18552,N_15148,N_16755);
xnor U18553 (N_18553,N_15488,N_16555);
or U18554 (N_18554,N_15512,N_15242);
xnor U18555 (N_18555,N_15368,N_16148);
nor U18556 (N_18556,N_16674,N_15457);
nor U18557 (N_18557,N_15409,N_15947);
xnor U18558 (N_18558,N_16709,N_15561);
and U18559 (N_18559,N_15567,N_17255);
xor U18560 (N_18560,N_16368,N_15104);
or U18561 (N_18561,N_15616,N_15025);
nor U18562 (N_18562,N_17473,N_15735);
or U18563 (N_18563,N_15495,N_15511);
xnor U18564 (N_18564,N_15140,N_16906);
xor U18565 (N_18565,N_16656,N_15030);
nand U18566 (N_18566,N_15295,N_15833);
nand U18567 (N_18567,N_15751,N_16405);
xnor U18568 (N_18568,N_15129,N_15938);
and U18569 (N_18569,N_15053,N_16284);
xor U18570 (N_18570,N_15624,N_16495);
nor U18571 (N_18571,N_15912,N_17490);
nor U18572 (N_18572,N_15893,N_15350);
xnor U18573 (N_18573,N_16873,N_16720);
nand U18574 (N_18574,N_15342,N_16672);
nor U18575 (N_18575,N_15688,N_15865);
nor U18576 (N_18576,N_15240,N_17116);
or U18577 (N_18577,N_16760,N_17379);
xnor U18578 (N_18578,N_16134,N_16423);
nor U18579 (N_18579,N_16630,N_17409);
nand U18580 (N_18580,N_16577,N_16083);
xor U18581 (N_18581,N_15386,N_16311);
or U18582 (N_18582,N_16329,N_17373);
xor U18583 (N_18583,N_15594,N_15029);
or U18584 (N_18584,N_16209,N_15256);
xnor U18585 (N_18585,N_16207,N_16448);
nor U18586 (N_18586,N_16250,N_15202);
xnor U18587 (N_18587,N_15358,N_15878);
nor U18588 (N_18588,N_17194,N_15994);
and U18589 (N_18589,N_16133,N_15113);
nand U18590 (N_18590,N_15321,N_17220);
and U18591 (N_18591,N_17344,N_16242);
or U18592 (N_18592,N_16484,N_16526);
nand U18593 (N_18593,N_15866,N_16366);
and U18594 (N_18594,N_16852,N_15018);
xor U18595 (N_18595,N_15593,N_16010);
nor U18596 (N_18596,N_16644,N_16078);
nand U18597 (N_18597,N_17051,N_15967);
and U18598 (N_18598,N_15093,N_16903);
nor U18599 (N_18599,N_16963,N_15918);
and U18600 (N_18600,N_16895,N_15916);
nand U18601 (N_18601,N_15190,N_16874);
nand U18602 (N_18602,N_17412,N_16223);
nor U18603 (N_18603,N_17014,N_16804);
xnor U18604 (N_18604,N_16030,N_15765);
and U18605 (N_18605,N_16666,N_16616);
nor U18606 (N_18606,N_16515,N_17098);
and U18607 (N_18607,N_17076,N_15026);
nor U18608 (N_18608,N_16553,N_16275);
nor U18609 (N_18609,N_16882,N_15646);
nand U18610 (N_18610,N_16668,N_17100);
nand U18611 (N_18611,N_16077,N_15527);
or U18612 (N_18612,N_15909,N_16315);
and U18613 (N_18613,N_16791,N_17207);
nand U18614 (N_18614,N_17436,N_15733);
xor U18615 (N_18615,N_17080,N_17365);
nand U18616 (N_18616,N_17371,N_16080);
and U18617 (N_18617,N_15428,N_16226);
nand U18618 (N_18618,N_16442,N_16799);
nand U18619 (N_18619,N_16150,N_17138);
nand U18620 (N_18620,N_16520,N_15850);
xor U18621 (N_18621,N_15963,N_15152);
nor U18622 (N_18622,N_15581,N_16782);
and U18623 (N_18623,N_16772,N_17109);
nor U18624 (N_18624,N_15082,N_15981);
and U18625 (N_18625,N_15666,N_16803);
nand U18626 (N_18626,N_16259,N_16199);
and U18627 (N_18627,N_16608,N_15535);
nand U18628 (N_18628,N_16045,N_15832);
nor U18629 (N_18629,N_15712,N_15687);
nand U18630 (N_18630,N_15157,N_15659);
and U18631 (N_18631,N_16435,N_16166);
and U18632 (N_18632,N_15391,N_17443);
or U18633 (N_18633,N_16218,N_16273);
and U18634 (N_18634,N_16205,N_15541);
xnor U18635 (N_18635,N_16853,N_15695);
or U18636 (N_18636,N_15777,N_15271);
or U18637 (N_18637,N_15531,N_17026);
nand U18638 (N_18638,N_16384,N_15732);
nor U18639 (N_18639,N_15171,N_17479);
nor U18640 (N_18640,N_15870,N_16570);
xor U18641 (N_18641,N_16154,N_16033);
and U18642 (N_18642,N_15529,N_15187);
nor U18643 (N_18643,N_15686,N_15999);
nand U18644 (N_18644,N_15699,N_15829);
xor U18645 (N_18645,N_15502,N_17131);
nand U18646 (N_18646,N_16020,N_16222);
nand U18647 (N_18647,N_15322,N_17228);
and U18648 (N_18648,N_15323,N_15828);
nor U18649 (N_18649,N_17021,N_17011);
nor U18650 (N_18650,N_15175,N_15613);
nor U18651 (N_18651,N_16632,N_16881);
xnor U18652 (N_18652,N_17366,N_16766);
nand U18653 (N_18653,N_15418,N_15045);
or U18654 (N_18654,N_17030,N_15117);
nor U18655 (N_18655,N_17143,N_15707);
and U18656 (N_18656,N_16053,N_17480);
nor U18657 (N_18657,N_15445,N_16047);
nor U18658 (N_18658,N_15137,N_16652);
nor U18659 (N_18659,N_15842,N_17254);
nor U18660 (N_18660,N_16456,N_15074);
xor U18661 (N_18661,N_15085,N_16810);
xor U18662 (N_18662,N_15559,N_17493);
nand U18663 (N_18663,N_16660,N_15413);
nor U18664 (N_18664,N_16057,N_15858);
nand U18665 (N_18665,N_15181,N_16476);
or U18666 (N_18666,N_15500,N_16867);
xnor U18667 (N_18667,N_15710,N_16091);
or U18668 (N_18668,N_16411,N_15877);
nor U18669 (N_18669,N_15245,N_15362);
or U18670 (N_18670,N_17304,N_17374);
or U18671 (N_18671,N_17375,N_15435);
and U18672 (N_18672,N_15705,N_17238);
or U18673 (N_18673,N_16482,N_15262);
or U18674 (N_18674,N_15685,N_16586);
nor U18675 (N_18675,N_15887,N_15538);
xor U18676 (N_18676,N_15078,N_15433);
nor U18677 (N_18677,N_17388,N_17329);
xor U18678 (N_18678,N_17487,N_17148);
xnor U18679 (N_18679,N_16255,N_15948);
xor U18680 (N_18680,N_15217,N_16127);
and U18681 (N_18681,N_17240,N_17301);
and U18682 (N_18682,N_15035,N_15474);
or U18683 (N_18683,N_16878,N_17497);
nor U18684 (N_18684,N_15702,N_17425);
or U18685 (N_18685,N_17188,N_17239);
xnor U18686 (N_18686,N_16676,N_15182);
xnor U18687 (N_18687,N_15747,N_17401);
nor U18688 (N_18688,N_16069,N_16841);
nor U18689 (N_18689,N_15971,N_15943);
xor U18690 (N_18690,N_16917,N_17323);
and U18691 (N_18691,N_15224,N_15012);
nand U18692 (N_18692,N_16785,N_16613);
nand U18693 (N_18693,N_15319,N_15955);
and U18694 (N_18694,N_17427,N_16880);
nor U18695 (N_18695,N_15125,N_17137);
nor U18696 (N_18696,N_15824,N_15392);
and U18697 (N_18697,N_15515,N_16670);
nor U18698 (N_18698,N_17027,N_15758);
or U18699 (N_18699,N_16756,N_17039);
xnor U18700 (N_18700,N_15296,N_15972);
or U18701 (N_18701,N_16203,N_16706);
or U18702 (N_18702,N_16210,N_16400);
nand U18703 (N_18703,N_17317,N_16767);
xor U18704 (N_18704,N_16988,N_15849);
and U18705 (N_18705,N_15482,N_16213);
xnor U18706 (N_18706,N_17421,N_15557);
nor U18707 (N_18707,N_15232,N_15503);
nand U18708 (N_18708,N_16749,N_16819);
xor U18709 (N_18709,N_17310,N_15974);
nand U18710 (N_18710,N_16467,N_17355);
nand U18711 (N_18711,N_15805,N_15091);
and U18712 (N_18712,N_16909,N_15261);
nand U18713 (N_18713,N_16581,N_16999);
xnor U18714 (N_18714,N_15138,N_17028);
xnor U18715 (N_18715,N_16263,N_15205);
nand U18716 (N_18716,N_16927,N_16871);
nor U18717 (N_18717,N_15352,N_15614);
xor U18718 (N_18718,N_17499,N_15816);
nand U18719 (N_18719,N_16295,N_16564);
and U18720 (N_18720,N_16556,N_17272);
xor U18721 (N_18721,N_16824,N_16708);
nand U18722 (N_18722,N_15484,N_15479);
xnor U18723 (N_18723,N_15875,N_16432);
nand U18724 (N_18724,N_15102,N_16977);
nor U18725 (N_18725,N_15766,N_17308);
or U18726 (N_18726,N_16765,N_16208);
xnor U18727 (N_18727,N_16454,N_17258);
or U18728 (N_18728,N_15293,N_17041);
or U18729 (N_18729,N_17397,N_16888);
or U18730 (N_18730,N_16943,N_15965);
and U18731 (N_18731,N_16475,N_16481);
or U18732 (N_18732,N_16543,N_15361);
and U18733 (N_18733,N_16983,N_17463);
or U18734 (N_18734,N_15670,N_16849);
nand U18735 (N_18735,N_16087,N_16566);
xor U18736 (N_18736,N_16971,N_15667);
or U18737 (N_18737,N_17017,N_16574);
nand U18738 (N_18738,N_15898,N_15693);
nor U18739 (N_18739,N_15377,N_16728);
and U18740 (N_18740,N_16216,N_15248);
xor U18741 (N_18741,N_15197,N_16678);
or U18742 (N_18742,N_17214,N_17335);
nor U18743 (N_18743,N_15258,N_16296);
xnor U18744 (N_18744,N_16107,N_16716);
nor U18745 (N_18745,N_15260,N_17257);
nand U18746 (N_18746,N_17404,N_17333);
nand U18747 (N_18747,N_17198,N_16587);
nand U18748 (N_18748,N_17000,N_15400);
nand U18749 (N_18749,N_15055,N_15276);
nand U18750 (N_18750,N_15741,N_16702);
nand U18751 (N_18751,N_17261,N_16478);
or U18752 (N_18752,N_15633,N_16072);
or U18753 (N_18753,N_16873,N_16918);
or U18754 (N_18754,N_16472,N_16615);
and U18755 (N_18755,N_15184,N_17330);
or U18756 (N_18756,N_15401,N_16706);
or U18757 (N_18757,N_15504,N_15374);
or U18758 (N_18758,N_15489,N_17495);
nand U18759 (N_18759,N_17103,N_15993);
nand U18760 (N_18760,N_16462,N_16477);
nor U18761 (N_18761,N_16797,N_16817);
or U18762 (N_18762,N_15373,N_15405);
xor U18763 (N_18763,N_17110,N_15194);
nor U18764 (N_18764,N_16628,N_17350);
and U18765 (N_18765,N_16321,N_16166);
xor U18766 (N_18766,N_15328,N_16343);
nand U18767 (N_18767,N_17365,N_17040);
nand U18768 (N_18768,N_15163,N_15677);
xor U18769 (N_18769,N_15061,N_17442);
or U18770 (N_18770,N_16385,N_15806);
nand U18771 (N_18771,N_16016,N_16696);
nor U18772 (N_18772,N_15297,N_15323);
nor U18773 (N_18773,N_15672,N_16490);
and U18774 (N_18774,N_15082,N_16510);
and U18775 (N_18775,N_15773,N_16807);
xor U18776 (N_18776,N_17412,N_15060);
nand U18777 (N_18777,N_16830,N_16817);
nor U18778 (N_18778,N_16140,N_17441);
and U18779 (N_18779,N_17445,N_16089);
xor U18780 (N_18780,N_17213,N_15508);
and U18781 (N_18781,N_17388,N_16355);
xnor U18782 (N_18782,N_16162,N_16749);
nand U18783 (N_18783,N_15538,N_16721);
xnor U18784 (N_18784,N_15872,N_17270);
nand U18785 (N_18785,N_16068,N_16108);
or U18786 (N_18786,N_15606,N_16137);
xnor U18787 (N_18787,N_15893,N_15595);
nand U18788 (N_18788,N_15030,N_15360);
xnor U18789 (N_18789,N_16181,N_15188);
nand U18790 (N_18790,N_17091,N_16699);
or U18791 (N_18791,N_16329,N_16489);
and U18792 (N_18792,N_16122,N_15247);
or U18793 (N_18793,N_15412,N_15548);
nand U18794 (N_18794,N_15971,N_16547);
or U18795 (N_18795,N_17321,N_15292);
nand U18796 (N_18796,N_17477,N_15630);
and U18797 (N_18797,N_15850,N_15696);
and U18798 (N_18798,N_17232,N_17300);
or U18799 (N_18799,N_16529,N_16595);
or U18800 (N_18800,N_15925,N_15909);
nand U18801 (N_18801,N_16199,N_15312);
or U18802 (N_18802,N_16759,N_15202);
or U18803 (N_18803,N_15246,N_15435);
xor U18804 (N_18804,N_15095,N_15564);
and U18805 (N_18805,N_17169,N_16024);
and U18806 (N_18806,N_15685,N_15325);
nor U18807 (N_18807,N_15671,N_16988);
nand U18808 (N_18808,N_16615,N_16876);
xor U18809 (N_18809,N_15136,N_16983);
nand U18810 (N_18810,N_15993,N_15718);
and U18811 (N_18811,N_17464,N_15258);
xnor U18812 (N_18812,N_15491,N_16266);
or U18813 (N_18813,N_16479,N_15638);
and U18814 (N_18814,N_15364,N_16199);
xor U18815 (N_18815,N_15081,N_15678);
and U18816 (N_18816,N_17056,N_16630);
xor U18817 (N_18817,N_17074,N_16305);
and U18818 (N_18818,N_16344,N_15348);
nand U18819 (N_18819,N_16527,N_15416);
nor U18820 (N_18820,N_15300,N_16267);
nor U18821 (N_18821,N_16767,N_16321);
xnor U18822 (N_18822,N_16856,N_16717);
and U18823 (N_18823,N_15045,N_16089);
nor U18824 (N_18824,N_15910,N_17091);
nor U18825 (N_18825,N_17315,N_15146);
and U18826 (N_18826,N_16445,N_17084);
xnor U18827 (N_18827,N_15691,N_16058);
nand U18828 (N_18828,N_15044,N_16476);
nor U18829 (N_18829,N_16502,N_16638);
and U18830 (N_18830,N_16990,N_15889);
and U18831 (N_18831,N_16582,N_16068);
and U18832 (N_18832,N_16980,N_15252);
xnor U18833 (N_18833,N_16577,N_15475);
nand U18834 (N_18834,N_15241,N_16982);
or U18835 (N_18835,N_15934,N_16183);
or U18836 (N_18836,N_15369,N_16646);
or U18837 (N_18837,N_15205,N_15184);
xnor U18838 (N_18838,N_16669,N_17183);
xnor U18839 (N_18839,N_15220,N_17123);
or U18840 (N_18840,N_15095,N_17448);
xor U18841 (N_18841,N_15310,N_15663);
and U18842 (N_18842,N_17317,N_15074);
xnor U18843 (N_18843,N_15396,N_15790);
xor U18844 (N_18844,N_17157,N_16311);
xnor U18845 (N_18845,N_17441,N_15489);
nand U18846 (N_18846,N_15399,N_16190);
and U18847 (N_18847,N_16292,N_15420);
and U18848 (N_18848,N_15304,N_16858);
nand U18849 (N_18849,N_16628,N_16064);
or U18850 (N_18850,N_17470,N_16578);
nor U18851 (N_18851,N_16693,N_15083);
nand U18852 (N_18852,N_17137,N_15248);
nand U18853 (N_18853,N_16741,N_16759);
xor U18854 (N_18854,N_16972,N_15894);
or U18855 (N_18855,N_17136,N_16470);
and U18856 (N_18856,N_15973,N_16068);
or U18857 (N_18857,N_16509,N_15022);
and U18858 (N_18858,N_16183,N_16936);
or U18859 (N_18859,N_17382,N_15978);
or U18860 (N_18860,N_15332,N_15177);
nand U18861 (N_18861,N_15150,N_15391);
or U18862 (N_18862,N_15527,N_17207);
and U18863 (N_18863,N_15492,N_15761);
nor U18864 (N_18864,N_16562,N_15804);
nor U18865 (N_18865,N_16198,N_15419);
xnor U18866 (N_18866,N_15209,N_16951);
nand U18867 (N_18867,N_15632,N_15996);
nand U18868 (N_18868,N_16085,N_16389);
and U18869 (N_18869,N_15731,N_15920);
and U18870 (N_18870,N_15009,N_16051);
nand U18871 (N_18871,N_15192,N_15717);
nand U18872 (N_18872,N_15181,N_15424);
or U18873 (N_18873,N_15672,N_17174);
or U18874 (N_18874,N_16334,N_17061);
xor U18875 (N_18875,N_17200,N_16385);
xor U18876 (N_18876,N_16075,N_15573);
nor U18877 (N_18877,N_15701,N_16850);
nor U18878 (N_18878,N_16823,N_16205);
or U18879 (N_18879,N_15244,N_15537);
nor U18880 (N_18880,N_17459,N_15506);
or U18881 (N_18881,N_16011,N_15767);
nor U18882 (N_18882,N_15919,N_16444);
nand U18883 (N_18883,N_16548,N_16591);
xor U18884 (N_18884,N_16797,N_15111);
nor U18885 (N_18885,N_15282,N_16737);
nand U18886 (N_18886,N_17437,N_16351);
and U18887 (N_18887,N_16099,N_15419);
or U18888 (N_18888,N_15978,N_15001);
xnor U18889 (N_18889,N_17184,N_17092);
nand U18890 (N_18890,N_17059,N_15098);
xor U18891 (N_18891,N_15690,N_17297);
and U18892 (N_18892,N_15731,N_16188);
or U18893 (N_18893,N_15069,N_16582);
nand U18894 (N_18894,N_15542,N_15032);
nand U18895 (N_18895,N_15654,N_15174);
xnor U18896 (N_18896,N_15406,N_15923);
xnor U18897 (N_18897,N_15431,N_17411);
and U18898 (N_18898,N_17266,N_15014);
and U18899 (N_18899,N_16895,N_16186);
xor U18900 (N_18900,N_15362,N_16303);
and U18901 (N_18901,N_17320,N_17097);
or U18902 (N_18902,N_15540,N_16378);
xor U18903 (N_18903,N_16019,N_15392);
xnor U18904 (N_18904,N_16509,N_16434);
xor U18905 (N_18905,N_15689,N_17105);
xnor U18906 (N_18906,N_17350,N_16245);
and U18907 (N_18907,N_16062,N_17033);
xnor U18908 (N_18908,N_15800,N_16787);
or U18909 (N_18909,N_15862,N_17341);
nand U18910 (N_18910,N_15751,N_15352);
and U18911 (N_18911,N_15159,N_17257);
and U18912 (N_18912,N_17159,N_16706);
nor U18913 (N_18913,N_17298,N_16137);
nor U18914 (N_18914,N_15370,N_17193);
nor U18915 (N_18915,N_15348,N_15998);
nor U18916 (N_18916,N_16984,N_16758);
nand U18917 (N_18917,N_15292,N_16124);
nand U18918 (N_18918,N_16719,N_15302);
and U18919 (N_18919,N_16090,N_16285);
or U18920 (N_18920,N_16713,N_16094);
or U18921 (N_18921,N_17371,N_15311);
and U18922 (N_18922,N_16109,N_15351);
and U18923 (N_18923,N_16699,N_16024);
nor U18924 (N_18924,N_17141,N_15505);
xnor U18925 (N_18925,N_16082,N_15919);
nand U18926 (N_18926,N_15214,N_16362);
or U18927 (N_18927,N_15493,N_17389);
and U18928 (N_18928,N_16399,N_16784);
and U18929 (N_18929,N_16678,N_17026);
xor U18930 (N_18930,N_16657,N_15474);
xor U18931 (N_18931,N_16197,N_15222);
or U18932 (N_18932,N_15311,N_16059);
nand U18933 (N_18933,N_15004,N_16797);
or U18934 (N_18934,N_15712,N_16422);
and U18935 (N_18935,N_15070,N_15437);
nor U18936 (N_18936,N_15500,N_16344);
or U18937 (N_18937,N_15765,N_15698);
nand U18938 (N_18938,N_16925,N_16864);
and U18939 (N_18939,N_15199,N_17032);
xnor U18940 (N_18940,N_15674,N_15920);
or U18941 (N_18941,N_16902,N_15349);
nand U18942 (N_18942,N_15039,N_16639);
nand U18943 (N_18943,N_17051,N_16166);
nor U18944 (N_18944,N_15063,N_16992);
xor U18945 (N_18945,N_17194,N_15972);
and U18946 (N_18946,N_16815,N_17463);
nor U18947 (N_18947,N_15175,N_16976);
nand U18948 (N_18948,N_16823,N_16411);
xor U18949 (N_18949,N_16431,N_16906);
or U18950 (N_18950,N_17339,N_16022);
nand U18951 (N_18951,N_16272,N_16810);
xor U18952 (N_18952,N_15068,N_15687);
xnor U18953 (N_18953,N_16309,N_15664);
nor U18954 (N_18954,N_16342,N_17306);
or U18955 (N_18955,N_15067,N_16064);
nand U18956 (N_18956,N_15958,N_15816);
xnor U18957 (N_18957,N_16983,N_16202);
nand U18958 (N_18958,N_15246,N_15057);
nand U18959 (N_18959,N_16630,N_15313);
xor U18960 (N_18960,N_16206,N_16900);
nand U18961 (N_18961,N_16483,N_15828);
and U18962 (N_18962,N_15179,N_15869);
nor U18963 (N_18963,N_17173,N_16361);
and U18964 (N_18964,N_15744,N_17311);
xnor U18965 (N_18965,N_16021,N_17443);
and U18966 (N_18966,N_16326,N_15647);
and U18967 (N_18967,N_15446,N_17405);
or U18968 (N_18968,N_16335,N_15084);
or U18969 (N_18969,N_16397,N_16573);
nand U18970 (N_18970,N_17440,N_17084);
or U18971 (N_18971,N_15166,N_16385);
and U18972 (N_18972,N_16237,N_17066);
and U18973 (N_18973,N_15145,N_17314);
and U18974 (N_18974,N_16375,N_15743);
nand U18975 (N_18975,N_15892,N_16069);
or U18976 (N_18976,N_17028,N_17460);
nor U18977 (N_18977,N_16715,N_16919);
nor U18978 (N_18978,N_16440,N_15514);
xor U18979 (N_18979,N_15946,N_16885);
xor U18980 (N_18980,N_17294,N_17054);
nor U18981 (N_18981,N_16750,N_15443);
or U18982 (N_18982,N_16401,N_15402);
nor U18983 (N_18983,N_16638,N_15829);
or U18984 (N_18984,N_17359,N_17154);
nor U18985 (N_18985,N_16693,N_17102);
or U18986 (N_18986,N_16871,N_15045);
and U18987 (N_18987,N_15719,N_16717);
or U18988 (N_18988,N_16804,N_15979);
nand U18989 (N_18989,N_16715,N_17289);
and U18990 (N_18990,N_17087,N_16090);
nand U18991 (N_18991,N_17474,N_15345);
or U18992 (N_18992,N_16896,N_16089);
and U18993 (N_18993,N_16204,N_15166);
and U18994 (N_18994,N_17253,N_15557);
and U18995 (N_18995,N_15905,N_15674);
nor U18996 (N_18996,N_16138,N_17176);
xnor U18997 (N_18997,N_15399,N_15681);
nor U18998 (N_18998,N_16816,N_15705);
nand U18999 (N_18999,N_15851,N_16714);
and U19000 (N_19000,N_16157,N_17186);
xor U19001 (N_19001,N_15152,N_16461);
nand U19002 (N_19002,N_16782,N_16346);
nor U19003 (N_19003,N_15894,N_16876);
nand U19004 (N_19004,N_17464,N_16479);
and U19005 (N_19005,N_15677,N_15867);
or U19006 (N_19006,N_16021,N_15532);
and U19007 (N_19007,N_17188,N_16051);
and U19008 (N_19008,N_16815,N_15201);
and U19009 (N_19009,N_15246,N_15271);
or U19010 (N_19010,N_15027,N_16027);
nor U19011 (N_19011,N_16935,N_16520);
nand U19012 (N_19012,N_17450,N_17038);
xnor U19013 (N_19013,N_16983,N_17034);
xnor U19014 (N_19014,N_17218,N_15334);
nor U19015 (N_19015,N_15131,N_15521);
nor U19016 (N_19016,N_17144,N_17270);
nand U19017 (N_19017,N_15762,N_15852);
nor U19018 (N_19018,N_17135,N_16008);
or U19019 (N_19019,N_16475,N_16373);
xor U19020 (N_19020,N_16744,N_16963);
nor U19021 (N_19021,N_15040,N_15271);
nor U19022 (N_19022,N_15008,N_15215);
nor U19023 (N_19023,N_16162,N_16343);
nor U19024 (N_19024,N_16778,N_16084);
xor U19025 (N_19025,N_15967,N_15666);
nand U19026 (N_19026,N_15525,N_17340);
nor U19027 (N_19027,N_16200,N_17176);
and U19028 (N_19028,N_17370,N_16238);
nor U19029 (N_19029,N_17167,N_16878);
or U19030 (N_19030,N_16253,N_16604);
nand U19031 (N_19031,N_16195,N_16900);
or U19032 (N_19032,N_16977,N_16965);
xor U19033 (N_19033,N_15487,N_16789);
nand U19034 (N_19034,N_16873,N_15838);
nand U19035 (N_19035,N_17228,N_15312);
xnor U19036 (N_19036,N_15877,N_16632);
and U19037 (N_19037,N_17427,N_16255);
xnor U19038 (N_19038,N_16867,N_16329);
or U19039 (N_19039,N_16654,N_15812);
nor U19040 (N_19040,N_15132,N_17239);
nor U19041 (N_19041,N_15535,N_15152);
nand U19042 (N_19042,N_15298,N_15427);
nor U19043 (N_19043,N_16271,N_17474);
or U19044 (N_19044,N_17049,N_17321);
nand U19045 (N_19045,N_16923,N_17249);
nand U19046 (N_19046,N_16654,N_16153);
or U19047 (N_19047,N_15672,N_15866);
or U19048 (N_19048,N_17400,N_15424);
xor U19049 (N_19049,N_15287,N_16352);
and U19050 (N_19050,N_17172,N_16269);
and U19051 (N_19051,N_17263,N_15451);
and U19052 (N_19052,N_15945,N_15083);
xnor U19053 (N_19053,N_15766,N_17116);
nand U19054 (N_19054,N_15769,N_15505);
nand U19055 (N_19055,N_17199,N_17448);
or U19056 (N_19056,N_16984,N_15126);
xnor U19057 (N_19057,N_17489,N_16299);
or U19058 (N_19058,N_15562,N_15932);
or U19059 (N_19059,N_15824,N_15285);
nand U19060 (N_19060,N_17102,N_16261);
nor U19061 (N_19061,N_16261,N_15114);
nor U19062 (N_19062,N_17257,N_15912);
and U19063 (N_19063,N_15455,N_15340);
or U19064 (N_19064,N_16190,N_16595);
or U19065 (N_19065,N_15508,N_16603);
nor U19066 (N_19066,N_15394,N_15836);
xnor U19067 (N_19067,N_15900,N_17212);
or U19068 (N_19068,N_15996,N_16591);
or U19069 (N_19069,N_15762,N_16612);
xnor U19070 (N_19070,N_15110,N_16774);
nor U19071 (N_19071,N_15223,N_16369);
nand U19072 (N_19072,N_17252,N_15339);
xnor U19073 (N_19073,N_15866,N_17394);
and U19074 (N_19074,N_15429,N_15113);
or U19075 (N_19075,N_17040,N_15725);
nor U19076 (N_19076,N_16662,N_16114);
and U19077 (N_19077,N_16191,N_15118);
nor U19078 (N_19078,N_16246,N_16520);
and U19079 (N_19079,N_16486,N_15426);
nor U19080 (N_19080,N_16357,N_15362);
xor U19081 (N_19081,N_15820,N_15327);
and U19082 (N_19082,N_15029,N_16180);
nand U19083 (N_19083,N_16867,N_17334);
nor U19084 (N_19084,N_16800,N_16792);
and U19085 (N_19085,N_17434,N_15083);
or U19086 (N_19086,N_15543,N_16976);
nand U19087 (N_19087,N_15033,N_16610);
and U19088 (N_19088,N_16535,N_15820);
nor U19089 (N_19089,N_17210,N_15961);
xnor U19090 (N_19090,N_15587,N_15156);
and U19091 (N_19091,N_16890,N_15056);
and U19092 (N_19092,N_15974,N_15197);
and U19093 (N_19093,N_16284,N_16681);
and U19094 (N_19094,N_16075,N_15241);
nor U19095 (N_19095,N_16533,N_15943);
nand U19096 (N_19096,N_17435,N_16643);
xor U19097 (N_19097,N_16057,N_16126);
nor U19098 (N_19098,N_16734,N_16012);
xor U19099 (N_19099,N_15978,N_17215);
and U19100 (N_19100,N_15663,N_16905);
and U19101 (N_19101,N_16515,N_17251);
or U19102 (N_19102,N_15494,N_15920);
nor U19103 (N_19103,N_15955,N_16133);
nor U19104 (N_19104,N_17455,N_16383);
nor U19105 (N_19105,N_16892,N_16183);
nor U19106 (N_19106,N_16313,N_17109);
nor U19107 (N_19107,N_16413,N_15787);
nand U19108 (N_19108,N_16870,N_16134);
nand U19109 (N_19109,N_17247,N_16753);
nand U19110 (N_19110,N_17234,N_15580);
and U19111 (N_19111,N_15550,N_16510);
or U19112 (N_19112,N_16708,N_17391);
nand U19113 (N_19113,N_15139,N_15639);
and U19114 (N_19114,N_16177,N_17354);
nand U19115 (N_19115,N_15100,N_16963);
nor U19116 (N_19116,N_15997,N_16995);
nor U19117 (N_19117,N_16674,N_17181);
or U19118 (N_19118,N_16309,N_15820);
or U19119 (N_19119,N_16739,N_15151);
xor U19120 (N_19120,N_15153,N_15122);
nand U19121 (N_19121,N_15621,N_16734);
nand U19122 (N_19122,N_16659,N_16568);
nor U19123 (N_19123,N_15437,N_16682);
nor U19124 (N_19124,N_15225,N_16020);
nor U19125 (N_19125,N_16274,N_17199);
and U19126 (N_19126,N_16048,N_17305);
xnor U19127 (N_19127,N_17303,N_15694);
or U19128 (N_19128,N_16296,N_15936);
nand U19129 (N_19129,N_15948,N_15426);
or U19130 (N_19130,N_16774,N_16691);
or U19131 (N_19131,N_15005,N_17448);
nor U19132 (N_19132,N_15491,N_17302);
xor U19133 (N_19133,N_16709,N_16256);
nand U19134 (N_19134,N_16578,N_15741);
and U19135 (N_19135,N_17312,N_16479);
or U19136 (N_19136,N_16469,N_15489);
and U19137 (N_19137,N_17385,N_16120);
nand U19138 (N_19138,N_15369,N_16074);
or U19139 (N_19139,N_16112,N_17085);
or U19140 (N_19140,N_15185,N_15003);
and U19141 (N_19141,N_15170,N_17058);
nor U19142 (N_19142,N_16054,N_15845);
or U19143 (N_19143,N_17163,N_16312);
xor U19144 (N_19144,N_16775,N_16553);
xnor U19145 (N_19145,N_15127,N_16224);
and U19146 (N_19146,N_15962,N_17256);
nor U19147 (N_19147,N_15806,N_16854);
or U19148 (N_19148,N_15230,N_16794);
xnor U19149 (N_19149,N_16529,N_16837);
nor U19150 (N_19150,N_15184,N_16382);
xnor U19151 (N_19151,N_16848,N_15079);
or U19152 (N_19152,N_16909,N_15571);
nand U19153 (N_19153,N_15384,N_15014);
or U19154 (N_19154,N_15163,N_17170);
or U19155 (N_19155,N_15741,N_17348);
nand U19156 (N_19156,N_16712,N_16948);
nor U19157 (N_19157,N_16973,N_16585);
nor U19158 (N_19158,N_15834,N_17132);
xor U19159 (N_19159,N_16577,N_15246);
or U19160 (N_19160,N_16513,N_15459);
nand U19161 (N_19161,N_17323,N_16863);
and U19162 (N_19162,N_15940,N_15244);
nor U19163 (N_19163,N_17447,N_15544);
nand U19164 (N_19164,N_15681,N_17484);
nor U19165 (N_19165,N_17136,N_15485);
or U19166 (N_19166,N_15116,N_16289);
or U19167 (N_19167,N_15932,N_15084);
nand U19168 (N_19168,N_16514,N_16847);
and U19169 (N_19169,N_15918,N_15194);
nand U19170 (N_19170,N_16535,N_15522);
and U19171 (N_19171,N_16135,N_16569);
xnor U19172 (N_19172,N_16314,N_17273);
or U19173 (N_19173,N_15813,N_16104);
xnor U19174 (N_19174,N_15819,N_16807);
and U19175 (N_19175,N_15196,N_16352);
nand U19176 (N_19176,N_16525,N_16895);
nand U19177 (N_19177,N_16796,N_17373);
xor U19178 (N_19178,N_16561,N_15326);
and U19179 (N_19179,N_16643,N_17046);
xor U19180 (N_19180,N_15891,N_15855);
nand U19181 (N_19181,N_15995,N_15845);
and U19182 (N_19182,N_15171,N_15620);
and U19183 (N_19183,N_15410,N_15990);
xor U19184 (N_19184,N_16672,N_16338);
xnor U19185 (N_19185,N_17195,N_16282);
nor U19186 (N_19186,N_15494,N_16887);
or U19187 (N_19187,N_16700,N_15583);
nand U19188 (N_19188,N_16069,N_15674);
nor U19189 (N_19189,N_16847,N_15142);
nor U19190 (N_19190,N_16700,N_16842);
and U19191 (N_19191,N_15303,N_16112);
nor U19192 (N_19192,N_15474,N_16525);
or U19193 (N_19193,N_17108,N_17423);
xnor U19194 (N_19194,N_15429,N_16075);
nand U19195 (N_19195,N_15405,N_16317);
and U19196 (N_19196,N_16425,N_16980);
or U19197 (N_19197,N_15155,N_15466);
nand U19198 (N_19198,N_15895,N_17381);
or U19199 (N_19199,N_16265,N_16423);
nand U19200 (N_19200,N_16752,N_16595);
nor U19201 (N_19201,N_17325,N_16190);
nor U19202 (N_19202,N_15526,N_15287);
xnor U19203 (N_19203,N_16188,N_16155);
nor U19204 (N_19204,N_16901,N_16443);
nor U19205 (N_19205,N_16800,N_17121);
nand U19206 (N_19206,N_15398,N_16894);
nor U19207 (N_19207,N_17252,N_15221);
nand U19208 (N_19208,N_17493,N_16734);
xnor U19209 (N_19209,N_15351,N_17094);
nand U19210 (N_19210,N_15376,N_16207);
nor U19211 (N_19211,N_15919,N_16586);
nor U19212 (N_19212,N_16958,N_17089);
and U19213 (N_19213,N_17397,N_16790);
or U19214 (N_19214,N_15053,N_15432);
and U19215 (N_19215,N_17350,N_16515);
nand U19216 (N_19216,N_15752,N_15700);
xnor U19217 (N_19217,N_16459,N_16745);
nor U19218 (N_19218,N_15005,N_16098);
and U19219 (N_19219,N_16832,N_16392);
or U19220 (N_19220,N_17170,N_16427);
xor U19221 (N_19221,N_17266,N_16018);
and U19222 (N_19222,N_15091,N_16920);
and U19223 (N_19223,N_15930,N_16823);
nand U19224 (N_19224,N_16768,N_17403);
and U19225 (N_19225,N_16527,N_16105);
xor U19226 (N_19226,N_16942,N_16655);
and U19227 (N_19227,N_17137,N_15245);
and U19228 (N_19228,N_16271,N_15560);
xnor U19229 (N_19229,N_16173,N_15200);
nand U19230 (N_19230,N_15945,N_15768);
and U19231 (N_19231,N_16133,N_15257);
xnor U19232 (N_19232,N_16594,N_17134);
or U19233 (N_19233,N_17130,N_16172);
xor U19234 (N_19234,N_16582,N_17410);
nand U19235 (N_19235,N_15144,N_16482);
nor U19236 (N_19236,N_16292,N_15955);
nor U19237 (N_19237,N_16656,N_16406);
nor U19238 (N_19238,N_16877,N_17198);
nor U19239 (N_19239,N_16119,N_15929);
or U19240 (N_19240,N_16705,N_15094);
nor U19241 (N_19241,N_16678,N_15342);
nor U19242 (N_19242,N_15261,N_16375);
and U19243 (N_19243,N_15303,N_15212);
and U19244 (N_19244,N_16452,N_16214);
nor U19245 (N_19245,N_16773,N_16562);
or U19246 (N_19246,N_16142,N_15813);
or U19247 (N_19247,N_16246,N_16322);
nor U19248 (N_19248,N_16262,N_16999);
nor U19249 (N_19249,N_15437,N_15375);
nand U19250 (N_19250,N_17305,N_17449);
nor U19251 (N_19251,N_15169,N_16221);
nand U19252 (N_19252,N_15786,N_15935);
nand U19253 (N_19253,N_16881,N_15522);
xor U19254 (N_19254,N_17071,N_17142);
nand U19255 (N_19255,N_15111,N_16042);
nand U19256 (N_19256,N_15836,N_16643);
nand U19257 (N_19257,N_16626,N_15485);
xnor U19258 (N_19258,N_15836,N_16617);
nand U19259 (N_19259,N_16807,N_15969);
nand U19260 (N_19260,N_16951,N_15772);
or U19261 (N_19261,N_17334,N_17432);
xor U19262 (N_19262,N_17399,N_15722);
or U19263 (N_19263,N_15552,N_17191);
or U19264 (N_19264,N_16928,N_17017);
and U19265 (N_19265,N_17090,N_15569);
nand U19266 (N_19266,N_16982,N_15773);
xnor U19267 (N_19267,N_16456,N_15147);
xnor U19268 (N_19268,N_15785,N_15953);
or U19269 (N_19269,N_17117,N_17025);
nand U19270 (N_19270,N_17247,N_16632);
nor U19271 (N_19271,N_15241,N_16734);
or U19272 (N_19272,N_16022,N_17325);
nor U19273 (N_19273,N_16436,N_15809);
nor U19274 (N_19274,N_15974,N_16184);
or U19275 (N_19275,N_16976,N_15813);
nand U19276 (N_19276,N_15034,N_16448);
and U19277 (N_19277,N_15373,N_15905);
nor U19278 (N_19278,N_17122,N_16956);
nor U19279 (N_19279,N_16574,N_17042);
nand U19280 (N_19280,N_16866,N_16775);
nor U19281 (N_19281,N_15627,N_16310);
nor U19282 (N_19282,N_15850,N_15271);
or U19283 (N_19283,N_16019,N_16030);
and U19284 (N_19284,N_15273,N_15490);
or U19285 (N_19285,N_17022,N_17328);
or U19286 (N_19286,N_16082,N_15219);
nor U19287 (N_19287,N_16530,N_15814);
xor U19288 (N_19288,N_17140,N_15443);
and U19289 (N_19289,N_15606,N_15063);
nor U19290 (N_19290,N_16990,N_15044);
and U19291 (N_19291,N_15880,N_16284);
nand U19292 (N_19292,N_15637,N_15638);
nand U19293 (N_19293,N_17234,N_15583);
nor U19294 (N_19294,N_16487,N_15991);
nor U19295 (N_19295,N_15812,N_15037);
and U19296 (N_19296,N_15457,N_17466);
xnor U19297 (N_19297,N_15469,N_15248);
nand U19298 (N_19298,N_16612,N_17261);
or U19299 (N_19299,N_16228,N_16274);
nor U19300 (N_19300,N_15845,N_15238);
nor U19301 (N_19301,N_15974,N_16356);
nand U19302 (N_19302,N_16915,N_15969);
or U19303 (N_19303,N_17425,N_16867);
or U19304 (N_19304,N_15039,N_16178);
and U19305 (N_19305,N_16680,N_16240);
or U19306 (N_19306,N_16771,N_17080);
xor U19307 (N_19307,N_16142,N_15461);
xor U19308 (N_19308,N_16937,N_16252);
nor U19309 (N_19309,N_15840,N_16850);
nor U19310 (N_19310,N_15826,N_16280);
or U19311 (N_19311,N_16157,N_16027);
xnor U19312 (N_19312,N_15142,N_15057);
xor U19313 (N_19313,N_16567,N_15612);
or U19314 (N_19314,N_16451,N_16122);
nand U19315 (N_19315,N_15562,N_16943);
or U19316 (N_19316,N_16861,N_17275);
xnor U19317 (N_19317,N_15198,N_15824);
nand U19318 (N_19318,N_16496,N_15894);
or U19319 (N_19319,N_16184,N_17037);
and U19320 (N_19320,N_15705,N_15701);
xor U19321 (N_19321,N_16161,N_17236);
nand U19322 (N_19322,N_16514,N_15990);
nor U19323 (N_19323,N_16770,N_17054);
nand U19324 (N_19324,N_17281,N_16797);
xor U19325 (N_19325,N_17054,N_17363);
or U19326 (N_19326,N_15218,N_17212);
or U19327 (N_19327,N_16541,N_17365);
or U19328 (N_19328,N_16653,N_15950);
nand U19329 (N_19329,N_15781,N_15139);
and U19330 (N_19330,N_17153,N_15287);
xor U19331 (N_19331,N_15633,N_15453);
or U19332 (N_19332,N_16519,N_15484);
or U19333 (N_19333,N_16144,N_15746);
nor U19334 (N_19334,N_16605,N_15087);
and U19335 (N_19335,N_17433,N_16924);
nor U19336 (N_19336,N_15346,N_15261);
nor U19337 (N_19337,N_15195,N_15120);
or U19338 (N_19338,N_15098,N_17311);
and U19339 (N_19339,N_15470,N_16196);
nor U19340 (N_19340,N_16485,N_16440);
nor U19341 (N_19341,N_16887,N_16698);
xnor U19342 (N_19342,N_15270,N_17157);
or U19343 (N_19343,N_16290,N_17284);
xnor U19344 (N_19344,N_15883,N_17239);
or U19345 (N_19345,N_15723,N_17310);
nor U19346 (N_19346,N_15062,N_15146);
nand U19347 (N_19347,N_15929,N_15124);
nand U19348 (N_19348,N_16541,N_16316);
xnor U19349 (N_19349,N_16831,N_16210);
xor U19350 (N_19350,N_15632,N_16378);
nand U19351 (N_19351,N_15239,N_17168);
nand U19352 (N_19352,N_16911,N_16578);
and U19353 (N_19353,N_16750,N_15441);
nand U19354 (N_19354,N_15271,N_16388);
nand U19355 (N_19355,N_15139,N_15653);
and U19356 (N_19356,N_16674,N_17435);
nand U19357 (N_19357,N_15049,N_15391);
xnor U19358 (N_19358,N_16511,N_16312);
or U19359 (N_19359,N_17012,N_15432);
nor U19360 (N_19360,N_17273,N_16713);
xnor U19361 (N_19361,N_15016,N_16480);
nor U19362 (N_19362,N_17375,N_16601);
or U19363 (N_19363,N_15524,N_15650);
or U19364 (N_19364,N_16128,N_17485);
nand U19365 (N_19365,N_15148,N_17172);
nand U19366 (N_19366,N_17088,N_16680);
nand U19367 (N_19367,N_16980,N_16228);
nor U19368 (N_19368,N_16001,N_16171);
or U19369 (N_19369,N_15173,N_16681);
xnor U19370 (N_19370,N_16176,N_16680);
nor U19371 (N_19371,N_17416,N_15365);
or U19372 (N_19372,N_15437,N_17254);
nor U19373 (N_19373,N_15442,N_17116);
or U19374 (N_19374,N_15082,N_16455);
or U19375 (N_19375,N_16602,N_15867);
xnor U19376 (N_19376,N_15850,N_15418);
or U19377 (N_19377,N_17006,N_15139);
or U19378 (N_19378,N_16398,N_16717);
or U19379 (N_19379,N_16149,N_16578);
or U19380 (N_19380,N_15299,N_16192);
xor U19381 (N_19381,N_16005,N_16567);
or U19382 (N_19382,N_16145,N_17031);
nor U19383 (N_19383,N_17073,N_17006);
xnor U19384 (N_19384,N_15317,N_16704);
nand U19385 (N_19385,N_16237,N_17058);
nor U19386 (N_19386,N_16832,N_15914);
or U19387 (N_19387,N_15881,N_15749);
nand U19388 (N_19388,N_16136,N_15491);
and U19389 (N_19389,N_17494,N_17320);
or U19390 (N_19390,N_15978,N_16043);
nand U19391 (N_19391,N_16584,N_15808);
nor U19392 (N_19392,N_16965,N_15562);
nand U19393 (N_19393,N_16841,N_15238);
nand U19394 (N_19394,N_15578,N_15177);
and U19395 (N_19395,N_17433,N_15270);
xor U19396 (N_19396,N_15341,N_16702);
xnor U19397 (N_19397,N_17431,N_16649);
nand U19398 (N_19398,N_16243,N_16714);
or U19399 (N_19399,N_17012,N_15734);
nor U19400 (N_19400,N_17444,N_15423);
xnor U19401 (N_19401,N_16056,N_15955);
xor U19402 (N_19402,N_17398,N_16123);
nor U19403 (N_19403,N_15293,N_15058);
and U19404 (N_19404,N_16136,N_16475);
and U19405 (N_19405,N_15540,N_16684);
nor U19406 (N_19406,N_15214,N_17136);
nand U19407 (N_19407,N_16786,N_16286);
nand U19408 (N_19408,N_15686,N_16751);
nor U19409 (N_19409,N_15804,N_17140);
xor U19410 (N_19410,N_15600,N_17141);
xor U19411 (N_19411,N_17413,N_16409);
nand U19412 (N_19412,N_15004,N_17402);
nor U19413 (N_19413,N_16641,N_17326);
or U19414 (N_19414,N_16949,N_15269);
and U19415 (N_19415,N_16693,N_16143);
nor U19416 (N_19416,N_15144,N_15616);
nand U19417 (N_19417,N_17149,N_17420);
xnor U19418 (N_19418,N_15644,N_16091);
and U19419 (N_19419,N_16222,N_15575);
nand U19420 (N_19420,N_15518,N_16631);
and U19421 (N_19421,N_17193,N_15480);
nand U19422 (N_19422,N_17477,N_17431);
or U19423 (N_19423,N_16950,N_15468);
nand U19424 (N_19424,N_15070,N_17151);
or U19425 (N_19425,N_16850,N_17289);
xnor U19426 (N_19426,N_17278,N_16074);
xor U19427 (N_19427,N_17148,N_15085);
xor U19428 (N_19428,N_15180,N_15445);
nand U19429 (N_19429,N_15511,N_16272);
and U19430 (N_19430,N_16027,N_16682);
and U19431 (N_19431,N_16723,N_17179);
xor U19432 (N_19432,N_16543,N_17245);
nor U19433 (N_19433,N_17126,N_15468);
nand U19434 (N_19434,N_16987,N_15983);
xor U19435 (N_19435,N_16748,N_16463);
or U19436 (N_19436,N_16360,N_15049);
nand U19437 (N_19437,N_16901,N_16503);
xnor U19438 (N_19438,N_15913,N_16100);
xnor U19439 (N_19439,N_15649,N_16993);
and U19440 (N_19440,N_16249,N_15755);
or U19441 (N_19441,N_15349,N_16372);
or U19442 (N_19442,N_16136,N_15437);
xor U19443 (N_19443,N_16445,N_15763);
xor U19444 (N_19444,N_15234,N_15294);
nand U19445 (N_19445,N_15921,N_15179);
xor U19446 (N_19446,N_15932,N_16026);
nand U19447 (N_19447,N_16679,N_16701);
nor U19448 (N_19448,N_16578,N_15120);
xor U19449 (N_19449,N_16136,N_16236);
nor U19450 (N_19450,N_17369,N_16132);
and U19451 (N_19451,N_16735,N_15301);
xor U19452 (N_19452,N_16284,N_15075);
xor U19453 (N_19453,N_15508,N_16919);
nand U19454 (N_19454,N_15025,N_17220);
xnor U19455 (N_19455,N_15183,N_17425);
nand U19456 (N_19456,N_16075,N_16530);
xnor U19457 (N_19457,N_16577,N_15630);
or U19458 (N_19458,N_17401,N_16523);
and U19459 (N_19459,N_15066,N_15413);
nand U19460 (N_19460,N_15037,N_17165);
nor U19461 (N_19461,N_16516,N_15990);
or U19462 (N_19462,N_16181,N_16384);
nor U19463 (N_19463,N_17394,N_16189);
and U19464 (N_19464,N_15259,N_15430);
xnor U19465 (N_19465,N_16364,N_15217);
and U19466 (N_19466,N_15504,N_17147);
nor U19467 (N_19467,N_16441,N_16566);
or U19468 (N_19468,N_15196,N_16358);
nand U19469 (N_19469,N_16660,N_16606);
or U19470 (N_19470,N_15950,N_17462);
nand U19471 (N_19471,N_15587,N_17117);
and U19472 (N_19472,N_16849,N_16761);
nor U19473 (N_19473,N_15743,N_17173);
xnor U19474 (N_19474,N_15495,N_15654);
and U19475 (N_19475,N_16467,N_16511);
nand U19476 (N_19476,N_15303,N_16525);
and U19477 (N_19477,N_16671,N_15275);
nand U19478 (N_19478,N_16475,N_16855);
xnor U19479 (N_19479,N_15358,N_15040);
nand U19480 (N_19480,N_16111,N_17107);
xnor U19481 (N_19481,N_16691,N_16676);
and U19482 (N_19482,N_15598,N_15038);
nand U19483 (N_19483,N_17451,N_16518);
nand U19484 (N_19484,N_16729,N_15741);
and U19485 (N_19485,N_15400,N_16762);
and U19486 (N_19486,N_15078,N_15108);
nor U19487 (N_19487,N_17329,N_15422);
nand U19488 (N_19488,N_15832,N_15520);
and U19489 (N_19489,N_16590,N_17279);
and U19490 (N_19490,N_15922,N_15687);
xor U19491 (N_19491,N_16532,N_15629);
or U19492 (N_19492,N_15562,N_16323);
and U19493 (N_19493,N_16204,N_16827);
xor U19494 (N_19494,N_17353,N_16055);
xnor U19495 (N_19495,N_15402,N_15812);
and U19496 (N_19496,N_16050,N_16758);
nor U19497 (N_19497,N_15591,N_17367);
nor U19498 (N_19498,N_17062,N_16149);
and U19499 (N_19499,N_16986,N_16488);
nand U19500 (N_19500,N_15658,N_17054);
and U19501 (N_19501,N_15993,N_16491);
and U19502 (N_19502,N_15474,N_15917);
nand U19503 (N_19503,N_16256,N_15750);
nor U19504 (N_19504,N_16839,N_16243);
and U19505 (N_19505,N_16059,N_16196);
nor U19506 (N_19506,N_15823,N_16048);
and U19507 (N_19507,N_15216,N_16242);
and U19508 (N_19508,N_15754,N_15787);
and U19509 (N_19509,N_15074,N_17428);
xnor U19510 (N_19510,N_16056,N_17221);
nor U19511 (N_19511,N_15891,N_15390);
or U19512 (N_19512,N_15091,N_16939);
nor U19513 (N_19513,N_15252,N_16673);
nand U19514 (N_19514,N_15499,N_15959);
nor U19515 (N_19515,N_17029,N_15007);
nand U19516 (N_19516,N_15328,N_15736);
or U19517 (N_19517,N_17225,N_15670);
nand U19518 (N_19518,N_15467,N_16962);
nand U19519 (N_19519,N_15359,N_17112);
and U19520 (N_19520,N_17074,N_16795);
xor U19521 (N_19521,N_17447,N_16637);
or U19522 (N_19522,N_16022,N_16356);
and U19523 (N_19523,N_15043,N_17305);
nand U19524 (N_19524,N_15201,N_16361);
nor U19525 (N_19525,N_16490,N_17433);
nor U19526 (N_19526,N_15990,N_16413);
xor U19527 (N_19527,N_16275,N_15770);
nand U19528 (N_19528,N_15159,N_16584);
nor U19529 (N_19529,N_16773,N_17314);
nand U19530 (N_19530,N_16468,N_17166);
nand U19531 (N_19531,N_16378,N_17417);
or U19532 (N_19532,N_15082,N_16263);
nor U19533 (N_19533,N_15686,N_16652);
nand U19534 (N_19534,N_15702,N_15929);
or U19535 (N_19535,N_16462,N_16139);
or U19536 (N_19536,N_16952,N_17022);
nor U19537 (N_19537,N_15661,N_16764);
nor U19538 (N_19538,N_16116,N_16016);
or U19539 (N_19539,N_16257,N_17429);
and U19540 (N_19540,N_17317,N_17173);
xnor U19541 (N_19541,N_16903,N_15450);
and U19542 (N_19542,N_16374,N_15484);
nand U19543 (N_19543,N_15350,N_15935);
xor U19544 (N_19544,N_16162,N_15270);
and U19545 (N_19545,N_16141,N_15841);
xor U19546 (N_19546,N_16564,N_16020);
and U19547 (N_19547,N_15617,N_16094);
and U19548 (N_19548,N_15798,N_16717);
xnor U19549 (N_19549,N_15785,N_15326);
xnor U19550 (N_19550,N_15560,N_16527);
xnor U19551 (N_19551,N_16615,N_15907);
nor U19552 (N_19552,N_17032,N_16333);
xor U19553 (N_19553,N_15733,N_17288);
nand U19554 (N_19554,N_15443,N_15050);
nand U19555 (N_19555,N_15924,N_15240);
or U19556 (N_19556,N_16370,N_17267);
nor U19557 (N_19557,N_17300,N_16292);
and U19558 (N_19558,N_15038,N_15713);
and U19559 (N_19559,N_15064,N_16715);
xnor U19560 (N_19560,N_16092,N_17463);
nor U19561 (N_19561,N_15264,N_15280);
nor U19562 (N_19562,N_16260,N_17067);
nand U19563 (N_19563,N_15666,N_16156);
nor U19564 (N_19564,N_16285,N_17329);
nand U19565 (N_19565,N_16071,N_15745);
nand U19566 (N_19566,N_17063,N_17147);
and U19567 (N_19567,N_15611,N_17408);
nor U19568 (N_19568,N_16425,N_16997);
or U19569 (N_19569,N_17286,N_15569);
xor U19570 (N_19570,N_17393,N_16192);
nand U19571 (N_19571,N_15640,N_15834);
nor U19572 (N_19572,N_16768,N_17030);
nand U19573 (N_19573,N_15119,N_16941);
and U19574 (N_19574,N_17007,N_17000);
or U19575 (N_19575,N_17044,N_16369);
or U19576 (N_19576,N_17461,N_16918);
or U19577 (N_19577,N_16059,N_15538);
or U19578 (N_19578,N_16774,N_16304);
nand U19579 (N_19579,N_15808,N_15300);
or U19580 (N_19580,N_16809,N_17229);
xor U19581 (N_19581,N_16396,N_16345);
nand U19582 (N_19582,N_17052,N_15222);
xnor U19583 (N_19583,N_15758,N_16826);
xor U19584 (N_19584,N_17303,N_16545);
nand U19585 (N_19585,N_16445,N_16744);
and U19586 (N_19586,N_17108,N_16933);
xnor U19587 (N_19587,N_15899,N_16458);
nand U19588 (N_19588,N_15160,N_15698);
xor U19589 (N_19589,N_15837,N_16771);
nand U19590 (N_19590,N_17193,N_17279);
xnor U19591 (N_19591,N_17319,N_17120);
or U19592 (N_19592,N_15251,N_17484);
nand U19593 (N_19593,N_16624,N_16328);
nand U19594 (N_19594,N_17411,N_15824);
and U19595 (N_19595,N_16596,N_15804);
nor U19596 (N_19596,N_15424,N_15571);
xor U19597 (N_19597,N_15925,N_17064);
nand U19598 (N_19598,N_15454,N_16808);
xnor U19599 (N_19599,N_15710,N_15237);
nand U19600 (N_19600,N_15393,N_15766);
nor U19601 (N_19601,N_15387,N_17334);
or U19602 (N_19602,N_17184,N_17109);
nor U19603 (N_19603,N_15580,N_17495);
and U19604 (N_19604,N_17336,N_17466);
nand U19605 (N_19605,N_17095,N_16049);
nand U19606 (N_19606,N_15039,N_16774);
or U19607 (N_19607,N_17218,N_16567);
xor U19608 (N_19608,N_15805,N_16257);
nand U19609 (N_19609,N_17162,N_16314);
and U19610 (N_19610,N_15700,N_15936);
nand U19611 (N_19611,N_15046,N_15522);
xor U19612 (N_19612,N_15128,N_15800);
xnor U19613 (N_19613,N_16339,N_15897);
xnor U19614 (N_19614,N_16048,N_15162);
nor U19615 (N_19615,N_16968,N_16649);
nor U19616 (N_19616,N_16430,N_16980);
or U19617 (N_19617,N_16607,N_16817);
nand U19618 (N_19618,N_17497,N_17459);
or U19619 (N_19619,N_16219,N_15400);
and U19620 (N_19620,N_16852,N_16423);
and U19621 (N_19621,N_16899,N_15371);
nand U19622 (N_19622,N_15720,N_17438);
or U19623 (N_19623,N_16203,N_16371);
xor U19624 (N_19624,N_15808,N_16673);
xor U19625 (N_19625,N_15380,N_15177);
and U19626 (N_19626,N_16665,N_15980);
and U19627 (N_19627,N_16639,N_15713);
nand U19628 (N_19628,N_16870,N_16055);
xor U19629 (N_19629,N_15170,N_16152);
nor U19630 (N_19630,N_17232,N_17184);
nor U19631 (N_19631,N_15591,N_16151);
or U19632 (N_19632,N_15188,N_17240);
nor U19633 (N_19633,N_15605,N_16544);
or U19634 (N_19634,N_16511,N_15469);
nor U19635 (N_19635,N_16187,N_15841);
xnor U19636 (N_19636,N_17019,N_15362);
xor U19637 (N_19637,N_15587,N_16747);
and U19638 (N_19638,N_16146,N_16936);
nor U19639 (N_19639,N_16948,N_17484);
nand U19640 (N_19640,N_17097,N_16152);
nor U19641 (N_19641,N_15528,N_15398);
nand U19642 (N_19642,N_16866,N_16354);
or U19643 (N_19643,N_15635,N_16690);
nand U19644 (N_19644,N_15869,N_16299);
and U19645 (N_19645,N_17061,N_16947);
and U19646 (N_19646,N_16332,N_17029);
and U19647 (N_19647,N_15473,N_16629);
or U19648 (N_19648,N_17419,N_16577);
and U19649 (N_19649,N_16523,N_15228);
nand U19650 (N_19650,N_15522,N_16542);
and U19651 (N_19651,N_15545,N_17323);
nand U19652 (N_19652,N_17402,N_16920);
xnor U19653 (N_19653,N_17420,N_15314);
and U19654 (N_19654,N_16844,N_17101);
xor U19655 (N_19655,N_16229,N_16284);
or U19656 (N_19656,N_17003,N_16039);
xor U19657 (N_19657,N_17116,N_16571);
nor U19658 (N_19658,N_15022,N_16364);
or U19659 (N_19659,N_15487,N_16783);
xnor U19660 (N_19660,N_16913,N_17103);
nand U19661 (N_19661,N_17033,N_16194);
xor U19662 (N_19662,N_16990,N_17428);
and U19663 (N_19663,N_17383,N_16672);
or U19664 (N_19664,N_16272,N_17415);
or U19665 (N_19665,N_15740,N_15239);
nor U19666 (N_19666,N_16381,N_17335);
nand U19667 (N_19667,N_16552,N_15911);
nor U19668 (N_19668,N_15130,N_16466);
and U19669 (N_19669,N_16307,N_15177);
xor U19670 (N_19670,N_15315,N_17479);
or U19671 (N_19671,N_15853,N_15176);
nor U19672 (N_19672,N_15471,N_15698);
nor U19673 (N_19673,N_17335,N_15816);
or U19674 (N_19674,N_17479,N_16271);
xnor U19675 (N_19675,N_17496,N_16274);
or U19676 (N_19676,N_16464,N_15798);
and U19677 (N_19677,N_15223,N_17210);
nand U19678 (N_19678,N_16283,N_15634);
nand U19679 (N_19679,N_16357,N_16278);
nand U19680 (N_19680,N_16700,N_15006);
nand U19681 (N_19681,N_15225,N_16118);
nand U19682 (N_19682,N_15512,N_17057);
xor U19683 (N_19683,N_17401,N_15447);
or U19684 (N_19684,N_15935,N_17028);
or U19685 (N_19685,N_17076,N_16877);
nand U19686 (N_19686,N_15028,N_15236);
or U19687 (N_19687,N_16582,N_15547);
or U19688 (N_19688,N_17174,N_15979);
xnor U19689 (N_19689,N_15391,N_15723);
nor U19690 (N_19690,N_17378,N_15808);
and U19691 (N_19691,N_16172,N_17278);
or U19692 (N_19692,N_16364,N_15842);
or U19693 (N_19693,N_15433,N_17196);
and U19694 (N_19694,N_16876,N_16830);
xor U19695 (N_19695,N_17292,N_16498);
nand U19696 (N_19696,N_16926,N_16819);
nand U19697 (N_19697,N_15834,N_16997);
and U19698 (N_19698,N_15608,N_16636);
nand U19699 (N_19699,N_15930,N_15239);
nor U19700 (N_19700,N_16056,N_17178);
nand U19701 (N_19701,N_15050,N_15805);
and U19702 (N_19702,N_15767,N_17366);
and U19703 (N_19703,N_17408,N_16587);
nand U19704 (N_19704,N_16196,N_17264);
xor U19705 (N_19705,N_16790,N_15766);
nor U19706 (N_19706,N_15338,N_16603);
and U19707 (N_19707,N_15532,N_16123);
xnor U19708 (N_19708,N_16042,N_16009);
nand U19709 (N_19709,N_16832,N_15155);
xor U19710 (N_19710,N_16089,N_15625);
and U19711 (N_19711,N_16428,N_16646);
and U19712 (N_19712,N_16026,N_17336);
and U19713 (N_19713,N_15975,N_15132);
xor U19714 (N_19714,N_16446,N_16318);
nor U19715 (N_19715,N_15827,N_17451);
and U19716 (N_19716,N_16829,N_16694);
and U19717 (N_19717,N_15588,N_16173);
and U19718 (N_19718,N_15221,N_16150);
nor U19719 (N_19719,N_15549,N_15073);
or U19720 (N_19720,N_15759,N_17486);
xnor U19721 (N_19721,N_15337,N_15063);
and U19722 (N_19722,N_17377,N_15638);
or U19723 (N_19723,N_16335,N_16297);
and U19724 (N_19724,N_17166,N_16461);
and U19725 (N_19725,N_16697,N_17131);
and U19726 (N_19726,N_16380,N_16919);
nand U19727 (N_19727,N_17111,N_17395);
nor U19728 (N_19728,N_17421,N_16872);
nand U19729 (N_19729,N_17106,N_17011);
or U19730 (N_19730,N_15418,N_17120);
nand U19731 (N_19731,N_16751,N_15284);
nor U19732 (N_19732,N_16235,N_16460);
and U19733 (N_19733,N_16543,N_16758);
xnor U19734 (N_19734,N_16839,N_17282);
or U19735 (N_19735,N_17318,N_16069);
nand U19736 (N_19736,N_16225,N_15854);
nand U19737 (N_19737,N_15846,N_16853);
and U19738 (N_19738,N_16082,N_16455);
and U19739 (N_19739,N_16897,N_16841);
xnor U19740 (N_19740,N_16672,N_15827);
and U19741 (N_19741,N_16870,N_16499);
xnor U19742 (N_19742,N_16229,N_16831);
or U19743 (N_19743,N_15259,N_16223);
or U19744 (N_19744,N_17468,N_16911);
nor U19745 (N_19745,N_16480,N_15739);
xnor U19746 (N_19746,N_16942,N_15350);
or U19747 (N_19747,N_15704,N_15436);
or U19748 (N_19748,N_17123,N_16589);
xnor U19749 (N_19749,N_16945,N_16883);
nand U19750 (N_19750,N_17011,N_15907);
nand U19751 (N_19751,N_15775,N_16534);
xor U19752 (N_19752,N_15552,N_16513);
and U19753 (N_19753,N_16397,N_17176);
or U19754 (N_19754,N_16417,N_15196);
xor U19755 (N_19755,N_16252,N_17410);
xor U19756 (N_19756,N_16051,N_16352);
and U19757 (N_19757,N_16263,N_17222);
and U19758 (N_19758,N_15379,N_17262);
or U19759 (N_19759,N_17191,N_15681);
and U19760 (N_19760,N_15179,N_15940);
or U19761 (N_19761,N_16418,N_16745);
nor U19762 (N_19762,N_15518,N_16640);
or U19763 (N_19763,N_16005,N_15076);
nand U19764 (N_19764,N_15703,N_16313);
xor U19765 (N_19765,N_16555,N_17464);
and U19766 (N_19766,N_16775,N_15260);
nor U19767 (N_19767,N_16323,N_15730);
nand U19768 (N_19768,N_15842,N_15560);
nor U19769 (N_19769,N_17395,N_15117);
and U19770 (N_19770,N_15706,N_15877);
and U19771 (N_19771,N_15647,N_15493);
nand U19772 (N_19772,N_16289,N_17365);
xor U19773 (N_19773,N_16148,N_17006);
and U19774 (N_19774,N_16788,N_17420);
nand U19775 (N_19775,N_17388,N_15921);
xor U19776 (N_19776,N_15881,N_16738);
xor U19777 (N_19777,N_15718,N_16684);
nand U19778 (N_19778,N_15552,N_16681);
nand U19779 (N_19779,N_17160,N_17356);
nor U19780 (N_19780,N_16785,N_15161);
nand U19781 (N_19781,N_16428,N_16569);
or U19782 (N_19782,N_16014,N_16959);
xnor U19783 (N_19783,N_15600,N_17238);
nand U19784 (N_19784,N_16695,N_16090);
or U19785 (N_19785,N_16459,N_15860);
or U19786 (N_19786,N_16991,N_16189);
nor U19787 (N_19787,N_17411,N_15987);
and U19788 (N_19788,N_16029,N_17061);
or U19789 (N_19789,N_16852,N_16097);
xor U19790 (N_19790,N_15949,N_15231);
or U19791 (N_19791,N_17494,N_16140);
xor U19792 (N_19792,N_17224,N_16353);
xnor U19793 (N_19793,N_17406,N_16383);
or U19794 (N_19794,N_15997,N_16112);
or U19795 (N_19795,N_15666,N_17488);
xor U19796 (N_19796,N_16812,N_16113);
xor U19797 (N_19797,N_17259,N_15001);
or U19798 (N_19798,N_15613,N_16358);
nor U19799 (N_19799,N_17222,N_16637);
xor U19800 (N_19800,N_16280,N_16087);
xnor U19801 (N_19801,N_15561,N_17024);
or U19802 (N_19802,N_17058,N_15953);
and U19803 (N_19803,N_16688,N_16599);
nand U19804 (N_19804,N_15826,N_15294);
and U19805 (N_19805,N_15316,N_17224);
and U19806 (N_19806,N_16108,N_16138);
and U19807 (N_19807,N_16161,N_17134);
and U19808 (N_19808,N_15962,N_15148);
or U19809 (N_19809,N_15754,N_15017);
nand U19810 (N_19810,N_17254,N_16018);
or U19811 (N_19811,N_17326,N_15961);
or U19812 (N_19812,N_15543,N_15139);
xor U19813 (N_19813,N_17259,N_15865);
nor U19814 (N_19814,N_17398,N_16147);
or U19815 (N_19815,N_16331,N_16538);
and U19816 (N_19816,N_15566,N_15433);
xnor U19817 (N_19817,N_16276,N_15965);
xor U19818 (N_19818,N_15097,N_16273);
and U19819 (N_19819,N_15763,N_17051);
or U19820 (N_19820,N_15396,N_15016);
nor U19821 (N_19821,N_15154,N_16688);
or U19822 (N_19822,N_17446,N_15635);
nand U19823 (N_19823,N_16957,N_16815);
xnor U19824 (N_19824,N_15488,N_16314);
and U19825 (N_19825,N_16600,N_15390);
or U19826 (N_19826,N_17393,N_15672);
nand U19827 (N_19827,N_17381,N_17118);
nand U19828 (N_19828,N_16428,N_16586);
or U19829 (N_19829,N_15442,N_15151);
and U19830 (N_19830,N_16587,N_15809);
nand U19831 (N_19831,N_16978,N_15846);
or U19832 (N_19832,N_17033,N_17040);
nand U19833 (N_19833,N_16905,N_15683);
or U19834 (N_19834,N_17177,N_17165);
or U19835 (N_19835,N_15082,N_15117);
or U19836 (N_19836,N_17461,N_17104);
or U19837 (N_19837,N_15605,N_15127);
nor U19838 (N_19838,N_15469,N_16282);
and U19839 (N_19839,N_15643,N_17491);
and U19840 (N_19840,N_15065,N_15926);
and U19841 (N_19841,N_16018,N_15697);
nand U19842 (N_19842,N_15954,N_15055);
or U19843 (N_19843,N_15697,N_15140);
and U19844 (N_19844,N_15467,N_17131);
and U19845 (N_19845,N_16647,N_16592);
or U19846 (N_19846,N_16946,N_16685);
nor U19847 (N_19847,N_16567,N_16339);
or U19848 (N_19848,N_15972,N_15994);
or U19849 (N_19849,N_16479,N_16581);
nor U19850 (N_19850,N_15115,N_15885);
nor U19851 (N_19851,N_15785,N_16668);
nor U19852 (N_19852,N_15469,N_16146);
nor U19853 (N_19853,N_16217,N_17034);
nor U19854 (N_19854,N_16695,N_16768);
and U19855 (N_19855,N_15355,N_16481);
nor U19856 (N_19856,N_15935,N_15627);
nor U19857 (N_19857,N_15991,N_17403);
nand U19858 (N_19858,N_16737,N_17446);
or U19859 (N_19859,N_16010,N_15950);
or U19860 (N_19860,N_16004,N_16897);
xnor U19861 (N_19861,N_17072,N_15808);
and U19862 (N_19862,N_15547,N_16039);
or U19863 (N_19863,N_15689,N_16175);
xor U19864 (N_19864,N_16648,N_17369);
nand U19865 (N_19865,N_16057,N_15778);
and U19866 (N_19866,N_16854,N_15927);
or U19867 (N_19867,N_16812,N_15630);
or U19868 (N_19868,N_15739,N_17396);
and U19869 (N_19869,N_17242,N_16039);
and U19870 (N_19870,N_17162,N_15137);
nor U19871 (N_19871,N_15600,N_17142);
nor U19872 (N_19872,N_16982,N_15150);
and U19873 (N_19873,N_17488,N_15326);
and U19874 (N_19874,N_15696,N_16836);
nor U19875 (N_19875,N_16296,N_16082);
and U19876 (N_19876,N_17069,N_15306);
nor U19877 (N_19877,N_17352,N_17185);
nand U19878 (N_19878,N_15724,N_16039);
nand U19879 (N_19879,N_15311,N_16850);
nor U19880 (N_19880,N_17168,N_16353);
nor U19881 (N_19881,N_16879,N_15425);
or U19882 (N_19882,N_17411,N_16018);
and U19883 (N_19883,N_16101,N_16921);
xor U19884 (N_19884,N_15599,N_16767);
xor U19885 (N_19885,N_17179,N_15248);
xor U19886 (N_19886,N_16177,N_16172);
nand U19887 (N_19887,N_16156,N_15806);
nor U19888 (N_19888,N_17028,N_15014);
nand U19889 (N_19889,N_16983,N_17249);
and U19890 (N_19890,N_17173,N_17463);
nor U19891 (N_19891,N_15432,N_15873);
nand U19892 (N_19892,N_16632,N_16288);
or U19893 (N_19893,N_16206,N_16257);
nand U19894 (N_19894,N_16057,N_15191);
nand U19895 (N_19895,N_15733,N_16577);
and U19896 (N_19896,N_15339,N_17041);
nor U19897 (N_19897,N_16452,N_16851);
or U19898 (N_19898,N_15570,N_15234);
and U19899 (N_19899,N_15495,N_15715);
and U19900 (N_19900,N_16301,N_15186);
nand U19901 (N_19901,N_15580,N_16025);
nand U19902 (N_19902,N_17493,N_16982);
nor U19903 (N_19903,N_16658,N_16394);
nand U19904 (N_19904,N_16224,N_17380);
xnor U19905 (N_19905,N_17032,N_15497);
and U19906 (N_19906,N_16714,N_16752);
xnor U19907 (N_19907,N_16791,N_15608);
and U19908 (N_19908,N_17093,N_15018);
or U19909 (N_19909,N_15610,N_17043);
xor U19910 (N_19910,N_16351,N_15241);
or U19911 (N_19911,N_15008,N_17020);
or U19912 (N_19912,N_15134,N_15369);
or U19913 (N_19913,N_17042,N_16741);
xnor U19914 (N_19914,N_16952,N_15327);
xor U19915 (N_19915,N_16334,N_16121);
xor U19916 (N_19916,N_15780,N_15942);
xor U19917 (N_19917,N_16992,N_15815);
nand U19918 (N_19918,N_15478,N_16222);
nor U19919 (N_19919,N_16825,N_17217);
nor U19920 (N_19920,N_16419,N_15761);
and U19921 (N_19921,N_15639,N_16227);
xor U19922 (N_19922,N_16804,N_16587);
or U19923 (N_19923,N_15616,N_17152);
nor U19924 (N_19924,N_16917,N_16250);
or U19925 (N_19925,N_15606,N_16666);
and U19926 (N_19926,N_16160,N_16316);
xnor U19927 (N_19927,N_16060,N_17022);
and U19928 (N_19928,N_16129,N_15495);
xor U19929 (N_19929,N_15770,N_15362);
xnor U19930 (N_19930,N_16763,N_16768);
nor U19931 (N_19931,N_16705,N_15288);
xnor U19932 (N_19932,N_16886,N_15103);
nor U19933 (N_19933,N_17154,N_16338);
and U19934 (N_19934,N_16937,N_15190);
and U19935 (N_19935,N_17480,N_15306);
nor U19936 (N_19936,N_16705,N_15727);
and U19937 (N_19937,N_15996,N_15412);
xor U19938 (N_19938,N_17369,N_16465);
nand U19939 (N_19939,N_16116,N_17347);
or U19940 (N_19940,N_16979,N_15222);
nand U19941 (N_19941,N_17403,N_17044);
xnor U19942 (N_19942,N_15891,N_16572);
and U19943 (N_19943,N_16928,N_17227);
or U19944 (N_19944,N_15842,N_16330);
nand U19945 (N_19945,N_16898,N_15432);
nand U19946 (N_19946,N_15369,N_15417);
or U19947 (N_19947,N_17315,N_17321);
or U19948 (N_19948,N_17442,N_16509);
or U19949 (N_19949,N_15476,N_17465);
or U19950 (N_19950,N_17488,N_16728);
nor U19951 (N_19951,N_17216,N_15863);
and U19952 (N_19952,N_15375,N_16448);
and U19953 (N_19953,N_16231,N_15311);
nor U19954 (N_19954,N_16235,N_16486);
nand U19955 (N_19955,N_17436,N_17367);
and U19956 (N_19956,N_17017,N_17415);
nor U19957 (N_19957,N_15690,N_16132);
or U19958 (N_19958,N_16904,N_15134);
or U19959 (N_19959,N_16906,N_17365);
nand U19960 (N_19960,N_17046,N_15599);
or U19961 (N_19961,N_16530,N_15764);
nand U19962 (N_19962,N_16843,N_17466);
and U19963 (N_19963,N_17382,N_17184);
and U19964 (N_19964,N_16535,N_15728);
xnor U19965 (N_19965,N_16376,N_16957);
nor U19966 (N_19966,N_17433,N_16106);
nand U19967 (N_19967,N_16463,N_15287);
and U19968 (N_19968,N_15520,N_17181);
nand U19969 (N_19969,N_16611,N_17261);
or U19970 (N_19970,N_16760,N_16833);
nand U19971 (N_19971,N_15396,N_15851);
and U19972 (N_19972,N_15355,N_16687);
xor U19973 (N_19973,N_17329,N_16812);
nand U19974 (N_19974,N_16097,N_16440);
nand U19975 (N_19975,N_16124,N_16885);
nand U19976 (N_19976,N_16267,N_17281);
nand U19977 (N_19977,N_16338,N_16295);
xnor U19978 (N_19978,N_17164,N_15181);
nand U19979 (N_19979,N_15413,N_16646);
and U19980 (N_19980,N_17327,N_16596);
xor U19981 (N_19981,N_15293,N_16268);
and U19982 (N_19982,N_16389,N_16873);
nor U19983 (N_19983,N_15060,N_16546);
nor U19984 (N_19984,N_16693,N_16313);
and U19985 (N_19985,N_15569,N_16470);
nor U19986 (N_19986,N_16194,N_16120);
and U19987 (N_19987,N_16667,N_15760);
or U19988 (N_19988,N_16360,N_16031);
nor U19989 (N_19989,N_16747,N_17010);
and U19990 (N_19990,N_15372,N_15104);
xor U19991 (N_19991,N_16439,N_17292);
and U19992 (N_19992,N_17418,N_16808);
nand U19993 (N_19993,N_15302,N_16577);
xnor U19994 (N_19994,N_17226,N_16827);
xor U19995 (N_19995,N_16398,N_15164);
xor U19996 (N_19996,N_17010,N_17447);
xnor U19997 (N_19997,N_17071,N_16515);
xnor U19998 (N_19998,N_17440,N_15830);
xnor U19999 (N_19999,N_15017,N_17142);
nand U20000 (N_20000,N_19396,N_18134);
xnor U20001 (N_20001,N_18486,N_19949);
and U20002 (N_20002,N_19023,N_18209);
nor U20003 (N_20003,N_18875,N_18837);
nand U20004 (N_20004,N_18353,N_17936);
and U20005 (N_20005,N_19835,N_19966);
nor U20006 (N_20006,N_19055,N_19323);
and U20007 (N_20007,N_18941,N_19439);
nand U20008 (N_20008,N_17883,N_19438);
nand U20009 (N_20009,N_18321,N_18064);
and U20010 (N_20010,N_17619,N_18729);
and U20011 (N_20011,N_17939,N_18653);
nor U20012 (N_20012,N_18590,N_19841);
xnor U20013 (N_20013,N_18559,N_19495);
xor U20014 (N_20014,N_19817,N_17555);
or U20015 (N_20015,N_18721,N_19540);
nand U20016 (N_20016,N_17801,N_17705);
nor U20017 (N_20017,N_19701,N_19277);
and U20018 (N_20018,N_19883,N_18476);
or U20019 (N_20019,N_19158,N_18635);
or U20020 (N_20020,N_18597,N_18129);
xnor U20021 (N_20021,N_18499,N_18539);
or U20022 (N_20022,N_19430,N_19991);
and U20023 (N_20023,N_17736,N_18211);
or U20024 (N_20024,N_19904,N_19785);
or U20025 (N_20025,N_19932,N_18581);
nor U20026 (N_20026,N_19382,N_19412);
xnor U20027 (N_20027,N_17903,N_19021);
nand U20028 (N_20028,N_17714,N_17972);
nor U20029 (N_20029,N_19106,N_19762);
and U20030 (N_20030,N_19857,N_19907);
or U20031 (N_20031,N_19369,N_19768);
or U20032 (N_20032,N_18423,N_19910);
and U20033 (N_20033,N_17851,N_17953);
xnor U20034 (N_20034,N_18548,N_19851);
xor U20035 (N_20035,N_18446,N_19291);
or U20036 (N_20036,N_19194,N_18582);
xnor U20037 (N_20037,N_18266,N_18143);
nor U20038 (N_20038,N_19811,N_17725);
and U20039 (N_20039,N_18177,N_18945);
nand U20040 (N_20040,N_18202,N_19088);
nor U20041 (N_20041,N_17968,N_19249);
xor U20042 (N_20042,N_17853,N_18487);
nor U20043 (N_20043,N_18053,N_19448);
nor U20044 (N_20044,N_18165,N_17734);
or U20045 (N_20045,N_19776,N_19180);
or U20046 (N_20046,N_19595,N_17647);
nand U20047 (N_20047,N_18869,N_18755);
nor U20048 (N_20048,N_18021,N_17676);
xor U20049 (N_20049,N_18550,N_19999);
nor U20050 (N_20050,N_19026,N_19225);
or U20051 (N_20051,N_18226,N_17803);
and U20052 (N_20052,N_19041,N_18271);
xnor U20053 (N_20053,N_19458,N_18455);
nor U20054 (N_20054,N_19507,N_18141);
nand U20055 (N_20055,N_18520,N_18528);
or U20056 (N_20056,N_18946,N_18010);
or U20057 (N_20057,N_18286,N_19905);
or U20058 (N_20058,N_18675,N_18799);
and U20059 (N_20059,N_17872,N_17909);
xor U20060 (N_20060,N_18359,N_19390);
or U20061 (N_20061,N_19693,N_19075);
or U20062 (N_20062,N_19102,N_19419);
nor U20063 (N_20063,N_18775,N_18648);
xnor U20064 (N_20064,N_19393,N_18467);
and U20065 (N_20065,N_19924,N_17686);
nand U20066 (N_20066,N_19029,N_19050);
and U20067 (N_20067,N_18567,N_19796);
nand U20068 (N_20068,N_18638,N_19282);
nor U20069 (N_20069,N_18504,N_18571);
xor U20070 (N_20070,N_19735,N_19141);
xnor U20071 (N_20071,N_18745,N_17822);
xor U20072 (N_20072,N_19349,N_19490);
or U20073 (N_20073,N_19379,N_17658);
nand U20074 (N_20074,N_17867,N_19053);
xor U20075 (N_20075,N_19696,N_19862);
and U20076 (N_20076,N_19231,N_19749);
nor U20077 (N_20077,N_19969,N_19128);
nand U20078 (N_20078,N_19274,N_19197);
and U20079 (N_20079,N_19228,N_18357);
xnor U20080 (N_20080,N_19046,N_19692);
nor U20081 (N_20081,N_17842,N_18480);
or U20082 (N_20082,N_19560,N_17528);
nand U20083 (N_20083,N_19486,N_18496);
xor U20084 (N_20084,N_19502,N_18771);
and U20085 (N_20085,N_19018,N_19844);
nand U20086 (N_20086,N_17825,N_19591);
nand U20087 (N_20087,N_19362,N_17958);
or U20088 (N_20088,N_17600,N_18676);
nor U20089 (N_20089,N_17761,N_18224);
and U20090 (N_20090,N_18599,N_19082);
or U20091 (N_20091,N_18050,N_19965);
nand U20092 (N_20092,N_19956,N_19901);
and U20093 (N_20093,N_17878,N_19188);
and U20094 (N_20094,N_19997,N_18960);
and U20095 (N_20095,N_18501,N_18909);
xnor U20096 (N_20096,N_19906,N_18629);
nor U20097 (N_20097,N_19415,N_18821);
nand U20098 (N_20098,N_17889,N_19518);
nor U20099 (N_20099,N_19056,N_18454);
nand U20100 (N_20100,N_18138,N_18984);
or U20101 (N_20101,N_19637,N_18944);
nor U20102 (N_20102,N_18898,N_18091);
nor U20103 (N_20103,N_18303,N_19004);
or U20104 (N_20104,N_19096,N_18565);
nand U20105 (N_20105,N_18131,N_18120);
nor U20106 (N_20106,N_19499,N_19423);
nand U20107 (N_20107,N_18758,N_18716);
or U20108 (N_20108,N_18937,N_17956);
xnor U20109 (N_20109,N_18623,N_18876);
and U20110 (N_20110,N_18324,N_19257);
nor U20111 (N_20111,N_17760,N_18686);
and U20112 (N_20112,N_18099,N_19121);
nand U20113 (N_20113,N_18412,N_19865);
and U20114 (N_20114,N_18166,N_19270);
nor U20115 (N_20115,N_18161,N_18116);
nand U20116 (N_20116,N_18636,N_17798);
and U20117 (N_20117,N_19480,N_18017);
nor U20118 (N_20118,N_19239,N_19162);
nand U20119 (N_20119,N_18335,N_18233);
nand U20120 (N_20120,N_18677,N_19112);
nand U20121 (N_20121,N_19936,N_18861);
nand U20122 (N_20122,N_18833,N_19359);
and U20123 (N_20123,N_18386,N_19453);
xor U20124 (N_20124,N_19047,N_18828);
and U20125 (N_20125,N_19947,N_18084);
and U20126 (N_20126,N_17911,N_17595);
nand U20127 (N_20127,N_18124,N_19827);
or U20128 (N_20128,N_18236,N_19977);
and U20129 (N_20129,N_19807,N_19243);
nand U20130 (N_20130,N_19996,N_19600);
xor U20131 (N_20131,N_18731,N_18052);
and U20132 (N_20132,N_18054,N_17787);
or U20133 (N_20133,N_19610,N_19957);
and U20134 (N_20134,N_19960,N_17532);
nand U20135 (N_20135,N_18664,N_17758);
and U20136 (N_20136,N_19424,N_18429);
or U20137 (N_20137,N_19979,N_18205);
nand U20138 (N_20138,N_17681,N_18525);
nand U20139 (N_20139,N_18179,N_19281);
nor U20140 (N_20140,N_18113,N_19131);
and U20141 (N_20141,N_18065,N_17777);
nor U20142 (N_20142,N_18047,N_18215);
or U20143 (N_20143,N_18870,N_18988);
or U20144 (N_20144,N_17844,N_19470);
and U20145 (N_20145,N_18155,N_19980);
nor U20146 (N_20146,N_18953,N_19392);
xnor U20147 (N_20147,N_19474,N_19992);
and U20148 (N_20148,N_19296,N_17654);
or U20149 (N_20149,N_18532,N_18261);
xor U20150 (N_20150,N_19466,N_17757);
or U20151 (N_20151,N_19034,N_17985);
and U20152 (N_20152,N_17567,N_19093);
xor U20153 (N_20153,N_18584,N_19802);
nor U20154 (N_20154,N_19090,N_17932);
nor U20155 (N_20155,N_19880,N_19210);
nand U20156 (N_20156,N_18048,N_17899);
xor U20157 (N_20157,N_17783,N_18100);
nor U20158 (N_20158,N_19577,N_18003);
nor U20159 (N_20159,N_19230,N_17662);
nand U20160 (N_20160,N_17680,N_18403);
or U20161 (N_20161,N_18829,N_19750);
xnor U20162 (N_20162,N_18690,N_18699);
nand U20163 (N_20163,N_18549,N_17922);
xnor U20164 (N_20164,N_19616,N_17652);
or U20165 (N_20165,N_17657,N_18368);
or U20166 (N_20166,N_18951,N_18045);
xor U20167 (N_20167,N_18297,N_19510);
nor U20168 (N_20168,N_18871,N_18471);
nor U20169 (N_20169,N_17625,N_17865);
or U20170 (N_20170,N_19397,N_18693);
and U20171 (N_20171,N_18231,N_18934);
and U20172 (N_20172,N_18826,N_19183);
nor U20173 (N_20173,N_18035,N_18092);
or U20174 (N_20174,N_19007,N_19437);
nand U20175 (N_20175,N_18268,N_19431);
or U20176 (N_20176,N_18254,N_19698);
or U20177 (N_20177,N_19298,N_19036);
nor U20178 (N_20178,N_18252,N_19982);
and U20179 (N_20179,N_19220,N_17963);
or U20180 (N_20180,N_17799,N_18272);
xor U20181 (N_20181,N_18601,N_19621);
xnor U20182 (N_20182,N_19516,N_18982);
and U20183 (N_20183,N_17523,N_17509);
xnor U20184 (N_20184,N_18665,N_19613);
and U20185 (N_20185,N_17781,N_17747);
or U20186 (N_20186,N_18557,N_18234);
or U20187 (N_20187,N_17768,N_17934);
xor U20188 (N_20188,N_18358,N_19729);
or U20189 (N_20189,N_18497,N_17780);
nand U20190 (N_20190,N_19655,N_17750);
and U20191 (N_20191,N_19297,N_19825);
nor U20192 (N_20192,N_18822,N_19712);
nor U20193 (N_20193,N_19653,N_19989);
nor U20194 (N_20194,N_19889,N_17898);
and U20195 (N_20195,N_19063,N_19142);
nand U20196 (N_20196,N_18634,N_19037);
nor U20197 (N_20197,N_18749,N_17916);
nand U20198 (N_20198,N_19011,N_19136);
and U20199 (N_20199,N_17887,N_17773);
nor U20200 (N_20200,N_18308,N_19867);
and U20201 (N_20201,N_17685,N_19689);
or U20202 (N_20202,N_17769,N_19363);
and U20203 (N_20203,N_19318,N_17752);
nand U20204 (N_20204,N_18466,N_19165);
xor U20205 (N_20205,N_18847,N_18872);
xnor U20206 (N_20206,N_19948,N_18023);
nand U20207 (N_20207,N_19548,N_18464);
nor U20208 (N_20208,N_19663,N_18865);
nor U20209 (N_20209,N_17581,N_18949);
xnor U20210 (N_20210,N_17744,N_18188);
nor U20211 (N_20211,N_18409,N_19464);
xnor U20212 (N_20212,N_18075,N_18442);
nor U20213 (N_20213,N_17827,N_17693);
and U20214 (N_20214,N_19832,N_17784);
xnor U20215 (N_20215,N_18850,N_19567);
xnor U20216 (N_20216,N_18685,N_17897);
and U20217 (N_20217,N_19624,N_18046);
or U20218 (N_20218,N_18614,N_17683);
nor U20219 (N_20219,N_18420,N_19280);
and U20220 (N_20220,N_18570,N_18517);
nand U20221 (N_20221,N_18733,N_18364);
or U20222 (N_20222,N_19308,N_18596);
nor U20223 (N_20223,N_19461,N_18316);
or U20224 (N_20224,N_19433,N_19067);
or U20225 (N_20225,N_19580,N_19273);
nand U20226 (N_20226,N_19787,N_18812);
xnor U20227 (N_20227,N_18132,N_19395);
nand U20228 (N_20228,N_18108,N_19923);
or U20229 (N_20229,N_19398,N_18313);
nor U20230 (N_20230,N_18203,N_19601);
and U20231 (N_20231,N_19452,N_17800);
nand U20232 (N_20232,N_19528,N_18873);
and U20233 (N_20233,N_18136,N_18877);
xor U20234 (N_20234,N_19682,N_18569);
xnor U20235 (N_20235,N_18394,N_18639);
nand U20236 (N_20236,N_19732,N_19734);
and U20237 (N_20237,N_19955,N_19240);
or U20238 (N_20238,N_18535,N_18462);
or U20239 (N_20239,N_17525,N_19761);
or U20240 (N_20240,N_18543,N_17863);
and U20241 (N_20241,N_18168,N_18798);
nand U20242 (N_20242,N_18106,N_17914);
nand U20243 (N_20243,N_17919,N_18456);
and U20244 (N_20244,N_19052,N_19048);
nand U20245 (N_20245,N_19019,N_18627);
and U20246 (N_20246,N_18818,N_17570);
and U20247 (N_20247,N_18621,N_17738);
xnor U20248 (N_20248,N_19607,N_19598);
xor U20249 (N_20249,N_18706,N_18808);
nand U20250 (N_20250,N_18175,N_18079);
or U20251 (N_20251,N_19976,N_18219);
nor U20252 (N_20252,N_18036,N_18253);
xnor U20253 (N_20253,N_19647,N_18162);
or U20254 (N_20254,N_18744,N_18383);
nand U20255 (N_20255,N_19890,N_18918);
and U20256 (N_20256,N_18836,N_19246);
nand U20257 (N_20257,N_19795,N_17650);
or U20258 (N_20258,N_18199,N_18698);
and U20259 (N_20259,N_19016,N_17874);
nand U20260 (N_20260,N_19632,N_19446);
xnor U20261 (N_20261,N_18576,N_18914);
or U20262 (N_20262,N_17824,N_18689);
nor U20263 (N_20263,N_19759,N_18327);
and U20264 (N_20264,N_18160,N_19385);
nand U20265 (N_20265,N_17712,N_19025);
or U20266 (N_20266,N_18326,N_19484);
nand U20267 (N_20267,N_18641,N_19557);
xnor U20268 (N_20268,N_18483,N_19990);
nand U20269 (N_20269,N_19138,N_18473);
and U20270 (N_20270,N_19893,N_18315);
and U20271 (N_20271,N_18555,N_17767);
nor U20272 (N_20272,N_18493,N_17518);
nand U20273 (N_20273,N_19833,N_19721);
nor U20274 (N_20274,N_19944,N_17500);
nor U20275 (N_20275,N_19185,N_17653);
or U20276 (N_20276,N_18007,N_18296);
nor U20277 (N_20277,N_17927,N_17710);
nor U20278 (N_20278,N_18238,N_18647);
and U20279 (N_20279,N_19572,N_18392);
xor U20280 (N_20280,N_18697,N_17537);
or U20281 (N_20281,N_17547,N_19354);
and U20282 (N_20282,N_17561,N_17735);
nor U20283 (N_20283,N_19937,N_19604);
nand U20284 (N_20284,N_19221,N_18938);
and U20285 (N_20285,N_19256,N_18411);
and U20286 (N_20286,N_17906,N_18391);
xor U20287 (N_20287,N_19603,N_19337);
nor U20288 (N_20288,N_18658,N_19677);
nor U20289 (N_20289,N_17794,N_18158);
nand U20290 (N_20290,N_19879,N_18849);
or U20291 (N_20291,N_18993,N_18086);
nor U20292 (N_20292,N_19706,N_18144);
nand U20293 (N_20293,N_18128,N_19711);
nand U20294 (N_20294,N_19266,N_18503);
nand U20295 (N_20295,N_19792,N_19513);
nand U20296 (N_20296,N_18593,N_17684);
nand U20297 (N_20297,N_17679,N_19312);
nand U20298 (N_20298,N_18484,N_19008);
xor U20299 (N_20299,N_19517,N_19565);
xor U20300 (N_20300,N_19953,N_17699);
nor U20301 (N_20301,N_18216,N_17539);
nand U20302 (N_20302,N_19497,N_18762);
nand U20303 (N_20303,N_18317,N_19463);
or U20304 (N_20304,N_18213,N_18961);
xor U20305 (N_20305,N_18246,N_19301);
or U20306 (N_20306,N_18996,N_19702);
or U20307 (N_20307,N_18970,N_17984);
xnor U20308 (N_20308,N_18974,N_17727);
and U20309 (N_20309,N_19163,N_18577);
or U20310 (N_20310,N_18591,N_18700);
or U20311 (N_20311,N_17704,N_18668);
xnor U20312 (N_20312,N_18150,N_18078);
nand U20313 (N_20313,N_18043,N_17772);
nand U20314 (N_20314,N_17622,N_19164);
nand U20315 (N_20315,N_19650,N_18458);
xnor U20316 (N_20316,N_17607,N_19127);
xor U20317 (N_20317,N_19235,N_17703);
and U20318 (N_20318,N_17568,N_19582);
and U20319 (N_20319,N_19330,N_19847);
or U20320 (N_20320,N_19781,N_18183);
nand U20321 (N_20321,N_17536,N_18221);
or U20322 (N_20322,N_18626,N_18475);
xor U20323 (N_20323,N_18972,N_18127);
nand U20324 (N_20324,N_17562,N_19739);
and U20325 (N_20325,N_19731,N_17740);
nor U20326 (N_20326,N_19837,N_19551);
nor U20327 (N_20327,N_18452,N_18580);
nor U20328 (N_20328,N_17741,N_19578);
xor U20329 (N_20329,N_18795,N_17908);
nor U20330 (N_20330,N_18190,N_18491);
or U20331 (N_20331,N_18310,N_17691);
xor U20332 (N_20332,N_19854,N_18044);
nand U20333 (N_20333,N_17942,N_18351);
or U20334 (N_20334,N_19987,N_18285);
nand U20335 (N_20335,N_19097,N_19355);
and U20336 (N_20336,N_18196,N_18575);
and U20337 (N_20337,N_18481,N_18145);
xnor U20338 (N_20338,N_18275,N_18025);
or U20339 (N_20339,N_19456,N_18217);
xor U20340 (N_20340,N_18172,N_19346);
nand U20341 (N_20341,N_19083,N_19079);
and U20342 (N_20342,N_18683,N_17791);
nand U20343 (N_20343,N_19814,N_19887);
nand U20344 (N_20344,N_18924,N_19175);
xnor U20345 (N_20345,N_18428,N_18232);
xor U20346 (N_20346,N_19681,N_19852);
nor U20347 (N_20347,N_17594,N_18192);
xnor U20348 (N_20348,N_18274,N_18478);
xor U20349 (N_20349,N_18650,N_18997);
and U20350 (N_20350,N_19631,N_18256);
or U20351 (N_20351,N_19575,N_19704);
or U20352 (N_20352,N_19813,N_19839);
and U20353 (N_20353,N_19483,N_17665);
or U20354 (N_20354,N_17690,N_19159);
nand U20355 (N_20355,N_17944,N_18752);
and U20356 (N_20356,N_17514,N_19917);
and U20357 (N_20357,N_18081,N_18193);
nand U20358 (N_20358,N_19413,N_19232);
xor U20359 (N_20359,N_18611,N_18425);
or U20360 (N_20360,N_19671,N_18319);
nand U20361 (N_20361,N_17632,N_19237);
nor U20362 (N_20362,N_17571,N_18374);
and U20363 (N_20363,N_19538,N_19238);
or U20364 (N_20364,N_19254,N_17764);
or U20365 (N_20365,N_18208,N_18556);
xnor U20366 (N_20366,N_18838,N_18606);
and U20367 (N_20367,N_19035,N_18076);
nand U20368 (N_20368,N_17621,N_18069);
or U20369 (N_20369,N_19658,N_19695);
nor U20370 (N_20370,N_19372,N_18171);
xor U20371 (N_20371,N_17976,N_19683);
and U20372 (N_20372,N_18255,N_18845);
xnor U20373 (N_20373,N_19933,N_18426);
nor U20374 (N_20374,N_19371,N_19771);
or U20375 (N_20375,N_19929,N_17847);
xnor U20376 (N_20376,N_19525,N_19199);
xnor U20377 (N_20377,N_17616,N_17876);
or U20378 (N_20378,N_18077,N_18016);
nor U20379 (N_20379,N_19328,N_19073);
xor U20380 (N_20380,N_17578,N_19251);
xor U20381 (N_20381,N_19092,N_18619);
nand U20382 (N_20382,N_18349,N_18149);
nand U20383 (N_20383,N_17795,N_17835);
and U20384 (N_20384,N_17651,N_18786);
nor U20385 (N_20385,N_18104,N_18402);
nand U20386 (N_20386,N_19533,N_19201);
nor U20387 (N_20387,N_19222,N_17510);
nand U20388 (N_20388,N_18059,N_18769);
nor U20389 (N_20389,N_18220,N_19039);
and U20390 (N_20390,N_19752,N_18718);
nand U20391 (N_20391,N_18547,N_18791);
nand U20392 (N_20392,N_19310,N_19515);
nor U20393 (N_20393,N_19680,N_18540);
or U20394 (N_20394,N_17614,N_18878);
nand U20395 (N_20395,N_18725,N_19375);
or U20396 (N_20396,N_18156,N_18325);
or U20397 (N_20397,N_19460,N_18692);
and U20398 (N_20398,N_18977,N_18336);
and U20399 (N_20399,N_19506,N_19592);
nor U20400 (N_20400,N_19845,N_19744);
and U20401 (N_20401,N_17587,N_18058);
and U20402 (N_20402,N_18856,N_18265);
nor U20403 (N_20403,N_17557,N_18019);
or U20404 (N_20404,N_17820,N_19491);
xor U20405 (N_20405,N_17974,N_17900);
nand U20406 (N_20406,N_19726,N_18612);
or U20407 (N_20407,N_18722,N_19736);
or U20408 (N_20408,N_18889,N_17950);
or U20409 (N_20409,N_18585,N_18770);
or U20410 (N_20410,N_18042,N_19182);
or U20411 (N_20411,N_17554,N_18470);
and U20412 (N_20412,N_18417,N_19728);
and U20413 (N_20413,N_17550,N_18527);
nand U20414 (N_20414,N_19676,N_17834);
or U20415 (N_20415,N_17765,N_18609);
or U20416 (N_20416,N_19236,N_19938);
and U20417 (N_20417,N_17648,N_18176);
or U20418 (N_20418,N_19267,N_17858);
or U20419 (N_20419,N_19125,N_17892);
nand U20420 (N_20420,N_19342,N_18737);
nand U20421 (N_20421,N_17678,N_18181);
xor U20422 (N_20422,N_17811,N_19585);
xnor U20423 (N_20423,N_18006,N_19263);
nor U20424 (N_20424,N_19898,N_19876);
nand U20425 (N_20425,N_19144,N_17638);
xor U20426 (N_20426,N_19897,N_18603);
nand U20427 (N_20427,N_19320,N_17655);
or U20428 (N_20428,N_19140,N_19118);
xnor U20429 (N_20429,N_18096,N_19786);
xnor U20430 (N_20430,N_19765,N_18250);
xnor U20431 (N_20431,N_18123,N_19512);
nor U20432 (N_20432,N_18682,N_17788);
or U20433 (N_20433,N_19022,N_17920);
nor U20434 (N_20434,N_18761,N_17885);
xnor U20435 (N_20435,N_18952,N_19198);
nor U20436 (N_20436,N_18735,N_19402);
xnor U20437 (N_20437,N_18257,N_19108);
xor U20438 (N_20438,N_19628,N_19511);
nand U20439 (N_20439,N_17633,N_18397);
nand U20440 (N_20440,N_18140,N_18242);
xor U20441 (N_20441,N_19849,N_17933);
and U20442 (N_20442,N_19756,N_19014);
and U20443 (N_20443,N_17831,N_19157);
nand U20444 (N_20444,N_19414,N_18788);
nor U20445 (N_20445,N_19935,N_19882);
xnor U20446 (N_20446,N_18897,N_19299);
xnor U20447 (N_20447,N_19559,N_17573);
or U20448 (N_20448,N_18995,N_19946);
nor U20449 (N_20449,N_19501,N_18142);
or U20450 (N_20450,N_17544,N_18090);
or U20451 (N_20451,N_19174,N_18276);
and U20452 (N_20452,N_18687,N_18029);
nand U20453 (N_20453,N_17626,N_18940);
and U20454 (N_20454,N_18978,N_18640);
or U20455 (N_20455,N_19531,N_18671);
or U20456 (N_20456,N_18578,N_18622);
nor U20457 (N_20457,N_19523,N_18508);
xor U20458 (N_20458,N_18151,N_18434);
xnor U20459 (N_20459,N_17879,N_18362);
nand U20460 (N_20460,N_18545,N_17864);
nand U20461 (N_20461,N_18874,N_19509);
nand U20462 (N_20462,N_17604,N_17507);
xnor U20463 (N_20463,N_19853,N_18976);
or U20464 (N_20464,N_19543,N_19068);
nor U20465 (N_20465,N_19838,N_19724);
nor U20466 (N_20466,N_19449,N_18920);
nand U20467 (N_20467,N_19091,N_18125);
and U20468 (N_20468,N_18290,N_18916);
or U20469 (N_20469,N_18477,N_17732);
xnor U20470 (N_20470,N_19360,N_19562);
nor U20471 (N_20471,N_18660,N_18943);
or U20472 (N_20472,N_19401,N_18115);
and U20473 (N_20473,N_19648,N_17960);
nand U20474 (N_20474,N_19115,N_19840);
or U20475 (N_20475,N_19766,N_19738);
or U20476 (N_20476,N_19196,N_19391);
xnor U20477 (N_20477,N_17702,N_17931);
or U20478 (N_20478,N_18200,N_18334);
or U20479 (N_20479,N_17511,N_17935);
xnor U20480 (N_20480,N_18933,N_18573);
or U20481 (N_20481,N_18880,N_18661);
xnor U20482 (N_20482,N_18345,N_18738);
xor U20483 (N_20483,N_18277,N_17610);
and U20484 (N_20484,N_17586,N_19815);
nand U20485 (N_20485,N_18249,N_18465);
or U20486 (N_20486,N_18009,N_18649);
or U20487 (N_20487,N_19477,N_17962);
xor U20488 (N_20488,N_19233,N_19444);
or U20489 (N_20489,N_17708,N_19836);
nand U20490 (N_20490,N_19149,N_19808);
or U20491 (N_20491,N_17771,N_17553);
or U20492 (N_20492,N_19903,N_18013);
nand U20493 (N_20493,N_17862,N_18506);
xnor U20494 (N_20494,N_18910,N_17793);
nor U20495 (N_20495,N_18247,N_19038);
nor U20496 (N_20496,N_17905,N_18381);
nand U20497 (N_20497,N_19454,N_18776);
xor U20498 (N_20498,N_18135,N_18824);
nand U20499 (N_20499,N_18363,N_18185);
xor U20500 (N_20500,N_17990,N_17964);
xor U20501 (N_20501,N_18989,N_19755);
or U20502 (N_20502,N_18057,N_19672);
nand U20503 (N_20503,N_17517,N_19877);
nor U20504 (N_20504,N_17928,N_19576);
xnor U20505 (N_20505,N_19856,N_17641);
xor U20506 (N_20506,N_17943,N_18212);
or U20507 (N_20507,N_19319,N_18337);
xnor U20508 (N_20508,N_17938,N_18842);
or U20509 (N_20509,N_18542,N_19451);
nor U20510 (N_20510,N_19745,N_19229);
xnor U20511 (N_20511,N_18890,N_19984);
nand U20512 (N_20512,N_19428,N_17718);
or U20513 (N_20513,N_19699,N_17875);
or U20514 (N_20514,N_18655,N_18028);
nor U20515 (N_20515,N_18588,N_18369);
xnor U20516 (N_20516,N_17924,N_18848);
nand U20517 (N_20517,N_17759,N_18892);
nor U20518 (N_20518,N_19153,N_18361);
and U20519 (N_20519,N_17877,N_18715);
nand U20520 (N_20520,N_18921,N_18169);
and U20521 (N_20521,N_17617,N_19450);
or U20522 (N_20522,N_19268,N_18544);
or U20523 (N_20523,N_17818,N_18121);
xnor U20524 (N_20524,N_18726,N_19919);
xor U20525 (N_20525,N_19304,N_18460);
and U20526 (N_20526,N_18062,N_19247);
and U20527 (N_20527,N_19057,N_19279);
or U20528 (N_20528,N_17672,N_18617);
and U20529 (N_20529,N_17521,N_17713);
nand U20530 (N_20530,N_18457,N_17873);
nand U20531 (N_20531,N_17808,N_18959);
xor U20532 (N_20532,N_18164,N_17722);
or U20533 (N_20533,N_18906,N_18210);
nor U20534 (N_20534,N_18302,N_18441);
xnor U20535 (N_20535,N_19272,N_18806);
xor U20536 (N_20536,N_19076,N_19058);
or U20537 (N_20537,N_18743,N_17513);
xor U20538 (N_20538,N_17564,N_19504);
nor U20539 (N_20539,N_18356,N_19252);
nand U20540 (N_20540,N_18522,N_17534);
or U20541 (N_20541,N_17698,N_19049);
xnor U20542 (N_20542,N_19060,N_18851);
and U20543 (N_20543,N_18939,N_18459);
xnor U20544 (N_20544,N_19920,N_18492);
nor U20545 (N_20545,N_19718,N_19561);
nand U20546 (N_20546,N_18839,N_19098);
and U20547 (N_20547,N_19794,N_18568);
xor U20548 (N_20548,N_17631,N_19044);
and U20549 (N_20549,N_18410,N_18002);
xnor U20550 (N_20550,N_19176,N_19555);
nand U20551 (N_20551,N_19714,N_19586);
nand U20552 (N_20552,N_19678,N_19553);
nand U20553 (N_20553,N_17574,N_17826);
nand U20554 (N_20554,N_19959,N_19061);
nand U20555 (N_20555,N_17749,N_19537);
xor U20556 (N_20556,N_18267,N_19657);
or U20557 (N_20557,N_18222,N_18507);
nand U20558 (N_20558,N_19978,N_18072);
and U20559 (N_20559,N_19974,N_18912);
nor U20560 (N_20560,N_18793,N_19260);
or U20561 (N_20561,N_18343,N_19574);
xor U20562 (N_20562,N_19485,N_17756);
and U20563 (N_20563,N_18804,N_17599);
xor U20564 (N_20564,N_19757,N_19894);
nor U20565 (N_20565,N_19380,N_18230);
or U20566 (N_20566,N_18620,N_18184);
xor U20567 (N_20567,N_19549,N_17664);
and U20568 (N_20568,N_18969,N_17526);
nand U20569 (N_20569,N_18524,N_18680);
or U20570 (N_20570,N_19488,N_19626);
nor U20571 (N_20571,N_19868,N_17975);
or U20572 (N_20572,N_17869,N_19001);
or U20573 (N_20573,N_18510,N_18347);
or U20574 (N_20574,N_18405,N_19322);
or U20575 (N_20575,N_19493,N_18957);
nand U20576 (N_20576,N_19383,N_19361);
nand U20577 (N_20577,N_17593,N_19130);
or U20578 (N_20578,N_19078,N_19244);
or U20579 (N_20579,N_19596,N_18862);
xnor U20580 (N_20580,N_18066,N_19192);
or U20581 (N_20581,N_18311,N_18797);
xnor U20582 (N_20582,N_19805,N_19986);
or U20583 (N_20583,N_19869,N_18366);
nand U20584 (N_20584,N_18884,N_17891);
nand U20585 (N_20585,N_18288,N_18186);
nand U20586 (N_20586,N_17527,N_18760);
xor U20587 (N_20587,N_19950,N_17669);
nand U20588 (N_20588,N_19527,N_18983);
xnor U20589 (N_20589,N_19740,N_17917);
or U20590 (N_20590,N_19881,N_18298);
xnor U20591 (N_20591,N_17577,N_19190);
nor U20592 (N_20592,N_19315,N_18846);
nand U20593 (N_20593,N_19764,N_17986);
xnor U20594 (N_20594,N_19309,N_17504);
xor U20595 (N_20595,N_18502,N_17694);
nand U20596 (N_20596,N_17785,N_18413);
xnor U20597 (N_20597,N_18679,N_18713);
or U20598 (N_20598,N_17980,N_19667);
xnor U20599 (N_20599,N_17910,N_18329);
xor U20600 (N_20600,N_18509,N_19223);
and U20601 (N_20601,N_19700,N_18586);
xor U20602 (N_20602,N_19307,N_18039);
or U20603 (N_20603,N_19200,N_18055);
nand U20604 (N_20604,N_19364,N_17821);
or U20605 (N_20605,N_17588,N_18061);
xnor U20606 (N_20606,N_18781,N_18270);
and U20607 (N_20607,N_18681,N_18225);
nor U20608 (N_20608,N_19614,N_19071);
xnor U20609 (N_20609,N_18170,N_18283);
xor U20610 (N_20610,N_18407,N_19666);
and U20611 (N_20611,N_19173,N_19816);
nor U20612 (N_20612,N_18538,N_18295);
and U20613 (N_20613,N_18739,N_19269);
and U20614 (N_20614,N_19120,N_19519);
and U20615 (N_20615,N_18756,N_19902);
nand U20616 (N_20616,N_17640,N_17753);
nor U20617 (N_20617,N_17629,N_19558);
and U20618 (N_20618,N_19045,N_19287);
and U20619 (N_20619,N_18073,N_19606);
or U20620 (N_20620,N_18322,N_18299);
or U20621 (N_20621,N_18024,N_19563);
and U20622 (N_20622,N_17731,N_19209);
xnor U20623 (N_20623,N_18421,N_18056);
and U20624 (N_20624,N_18439,N_19972);
and U20625 (N_20625,N_18696,N_19000);
or U20626 (N_20626,N_18854,N_19589);
nand U20627 (N_20627,N_18067,N_18783);
nor U20628 (N_20628,N_17841,N_18384);
xnor U20629 (N_20629,N_19215,N_19124);
nand U20630 (N_20630,N_17915,N_19147);
nor U20631 (N_20631,N_18757,N_18936);
xnor U20632 (N_20632,N_19760,N_19126);
or U20633 (N_20633,N_18333,N_17670);
or U20634 (N_20634,N_18643,N_19630);
and U20635 (N_20635,N_19258,N_18119);
nor U20636 (N_20636,N_17992,N_19072);
or U20637 (N_20637,N_18012,N_18103);
xor U20638 (N_20638,N_19089,N_17775);
or U20639 (N_20639,N_19546,N_18948);
nand U20640 (N_20640,N_18453,N_18998);
nor U20641 (N_20641,N_19564,N_17603);
nor U20642 (N_20642,N_18365,N_17804);
or U20643 (N_20643,N_19134,N_17812);
nor U20644 (N_20644,N_19394,N_19161);
nor U20645 (N_20645,N_18130,N_19387);
and U20646 (N_20646,N_17806,N_18947);
or U20647 (N_20647,N_19207,N_17782);
nor U20648 (N_20648,N_19416,N_18608);
nand U20649 (N_20649,N_17695,N_18490);
nand U20650 (N_20650,N_18049,N_19172);
nand U20651 (N_20651,N_19465,N_18985);
nor U20652 (N_20652,N_18536,N_19674);
xor U20653 (N_20653,N_18930,N_19971);
or U20654 (N_20654,N_18673,N_19915);
and U20655 (N_20655,N_18779,N_17659);
xor U20656 (N_20656,N_18840,N_19311);
or U20657 (N_20657,N_17815,N_19968);
and U20658 (N_20658,N_19030,N_17745);
nand U20659 (N_20659,N_18814,N_19733);
nor U20660 (N_20660,N_18642,N_17880);
nor U20661 (N_20661,N_18759,N_18235);
xor U20662 (N_20662,N_18885,N_19193);
nor U20663 (N_20663,N_18281,N_18973);
and U20664 (N_20664,N_18500,N_18448);
xnor U20665 (N_20665,N_19275,N_19489);
nand U20666 (N_20666,N_18197,N_19388);
or U20667 (N_20667,N_18163,N_18126);
xor U20668 (N_20668,N_17506,N_17997);
and U20669 (N_20669,N_19373,N_18282);
nand U20670 (N_20670,N_17682,N_18227);
nor U20671 (N_20671,N_17941,N_19803);
nand U20672 (N_20672,N_18907,N_18472);
xnor U20673 (N_20673,N_19099,N_19715);
and U20674 (N_20674,N_19656,N_19331);
xnor U20675 (N_20675,N_17560,N_18479);
and U20676 (N_20676,N_19262,N_17966);
nand U20677 (N_20677,N_19741,N_18723);
or U20678 (N_20678,N_18844,N_18292);
or U20679 (N_20679,N_19494,N_19292);
nand U20680 (N_20680,N_19169,N_19514);
nand U20681 (N_20681,N_19150,N_18001);
nor U20682 (N_20682,N_17717,N_19333);
and U20683 (N_20683,N_17819,N_19767);
xor U20684 (N_20684,N_18328,N_17623);
and U20685 (N_20685,N_19080,N_18741);
and U20686 (N_20686,N_18443,N_17709);
or U20687 (N_20687,N_19405,N_18832);
and U20688 (N_20688,N_17896,N_19922);
nand U20689 (N_20689,N_19661,N_17630);
nand U20690 (N_20690,N_18631,N_19443);
nor U20691 (N_20691,N_19788,N_17991);
nand U20692 (N_20692,N_18511,N_19583);
nor U20693 (N_20693,N_18109,N_19482);
or U20694 (N_20694,N_17529,N_19017);
xnor U20695 (N_20695,N_19476,N_19408);
and U20696 (N_20696,N_18962,N_18469);
or U20697 (N_20697,N_19107,N_17929);
or U20698 (N_20698,N_19863,N_19441);
nand U20699 (N_20699,N_18435,N_18427);
or U20700 (N_20700,N_17809,N_19440);
nor U20701 (N_20701,N_19104,N_19806);
xor U20702 (N_20702,N_19212,N_17618);
nor U20703 (N_20703,N_19469,N_19588);
xnor U20704 (N_20704,N_18223,N_17508);
nor U20705 (N_20705,N_18260,N_18494);
nand U20706 (N_20706,N_18782,N_19941);
xnor U20707 (N_20707,N_18157,N_18905);
nand U20708 (N_20708,N_19778,N_18037);
xor U20709 (N_20709,N_18809,N_18785);
nand U20710 (N_20710,N_18981,N_19028);
nor U20711 (N_20711,N_18098,N_18541);
nand U20712 (N_20712,N_17949,N_18917);
nand U20713 (N_20713,N_19539,N_19410);
or U20714 (N_20714,N_19707,N_19181);
nor U20715 (N_20715,N_17790,N_19885);
nor U20716 (N_20716,N_18923,N_19809);
or U20717 (N_20717,N_18750,N_19195);
and U20718 (N_20718,N_19900,N_18765);
nand U20719 (N_20719,N_17569,N_19399);
xor U20720 (N_20720,N_19675,N_19101);
and U20721 (N_20721,N_19264,N_17945);
or U20722 (N_20722,N_18008,N_19143);
nor U20723 (N_20723,N_18305,N_19316);
xor U20724 (N_20724,N_19952,N_17849);
nand U20725 (N_20725,N_18915,N_18153);
nand U20726 (N_20726,N_17838,N_19325);
nand U20727 (N_20727,N_18724,N_18882);
or U20728 (N_20728,N_19812,N_17559);
or U20729 (N_20729,N_19040,N_17840);
nand U20730 (N_20730,N_18746,N_18864);
and U20731 (N_20731,N_18041,N_19722);
or U20732 (N_20732,N_17692,N_19652);
or U20733 (N_20733,N_18958,N_19406);
nand U20734 (N_20734,N_18605,N_18736);
xnor U20735 (N_20735,N_18178,N_17994);
nor U20736 (N_20736,N_19973,N_18990);
or U20737 (N_20737,N_17546,N_18182);
or U20738 (N_20738,N_18422,N_17728);
and U20739 (N_20739,N_17754,N_17596);
nand U20740 (N_20740,N_19943,N_18005);
and U20741 (N_20741,N_18070,N_17688);
nor U20742 (N_20742,N_19368,N_17856);
nand U20743 (N_20743,N_19117,N_19524);
xnor U20744 (N_20744,N_19798,N_17558);
xnor U20745 (N_20745,N_18859,N_18340);
and U20746 (N_20746,N_17584,N_17726);
and U20747 (N_20747,N_17580,N_19685);
or U20748 (N_20748,N_18895,N_19926);
or U20749 (N_20749,N_18787,N_19995);
nor U20750 (N_20750,N_18780,N_19581);
nand U20751 (N_20751,N_18926,N_19975);
nor U20752 (N_20752,N_19166,N_19335);
nor U20753 (N_20753,N_17637,N_18688);
or U20754 (N_20754,N_19899,N_19300);
and U20755 (N_20755,N_19526,N_19178);
xor U20756 (N_20756,N_19293,N_18214);
or U20757 (N_20757,N_19462,N_18810);
nand U20758 (N_20758,N_17746,N_19800);
nand U20759 (N_20759,N_18925,N_18807);
nor U20760 (N_20760,N_17572,N_19148);
xnor U20761 (N_20761,N_17677,N_17971);
and U20762 (N_20762,N_17512,N_19521);
or U20763 (N_20763,N_18287,N_19646);
nor U20764 (N_20764,N_18600,N_17589);
or U20765 (N_20765,N_19250,N_19697);
or U20766 (N_20766,N_18618,N_19003);
nor U20767 (N_20767,N_18348,N_19404);
nand U20768 (N_20768,N_19289,N_17776);
nand U20769 (N_20769,N_19326,N_18264);
nand U20770 (N_20770,N_19226,N_19024);
nor U20771 (N_20771,N_19945,N_18887);
and U20772 (N_20772,N_18331,N_19145);
nor U20773 (N_20773,N_18816,N_17881);
xor U20774 (N_20774,N_17870,N_19302);
and U20775 (N_20775,N_18927,N_19859);
or U20776 (N_20776,N_18341,N_18060);
nand U20777 (N_20777,N_18908,N_18894);
or U20778 (N_20778,N_19659,N_18523);
or U20779 (N_20779,N_18237,N_19179);
xor U20780 (N_20780,N_17854,N_19691);
or U20781 (N_20781,N_19855,N_17837);
and U20782 (N_20782,N_17644,N_18521);
nor U20783 (N_20783,N_19891,N_19204);
and U20784 (N_20784,N_18717,N_19820);
nor U20785 (N_20785,N_19668,N_19763);
xnor U20786 (N_20786,N_19873,N_19187);
nor U20787 (N_20787,N_18684,N_18330);
and U20788 (N_20788,N_19860,N_18000);
and U20789 (N_20789,N_17832,N_18727);
nor U20790 (N_20790,N_19896,N_17959);
nor U20791 (N_20791,N_19871,N_18695);
and U20792 (N_20792,N_19643,N_19679);
nand U20793 (N_20793,N_18139,N_19569);
and U20794 (N_20794,N_18607,N_19620);
nand U20795 (N_20795,N_17860,N_18899);
xor U20796 (N_20796,N_19114,N_19612);
and U20797 (N_20797,N_19208,N_17597);
nor U20798 (N_20798,N_19609,N_18667);
xor U20799 (N_20799,N_19191,N_19791);
and U20800 (N_20800,N_19916,N_19964);
nor U20801 (N_20801,N_18245,N_17967);
nand U20802 (N_20802,N_18891,N_19069);
nor U20803 (N_20803,N_19753,N_19087);
and U20804 (N_20804,N_17982,N_17993);
xnor U20805 (N_20805,N_17766,N_18371);
xnor U20806 (N_20806,N_17639,N_19593);
and U20807 (N_20807,N_18904,N_19535);
nor U20808 (N_20808,N_17948,N_18154);
and U20809 (N_20809,N_18263,N_19227);
and U20810 (N_20810,N_18956,N_18338);
nor U20811 (N_20811,N_17998,N_19374);
or U20812 (N_20812,N_18244,N_17894);
or U20813 (N_20813,N_19219,N_19622);
and U20814 (N_20814,N_18594,N_18440);
nor U20815 (N_20815,N_17751,N_19160);
xnor U20816 (N_20816,N_19154,N_18445);
nand U20817 (N_20817,N_18097,N_19492);
and U20818 (N_20818,N_18415,N_19305);
nand U20819 (N_20819,N_18740,N_18033);
and U20820 (N_20820,N_19253,N_18777);
xnor U20821 (N_20821,N_17965,N_17807);
or U20822 (N_20822,N_17937,N_18867);
xnor U20823 (N_20823,N_19587,N_18307);
nor U20824 (N_20824,N_18602,N_18218);
and U20825 (N_20825,N_18881,N_18963);
or U20826 (N_20826,N_19345,N_19321);
xor U20827 (N_20827,N_19206,N_18147);
nor U20828 (N_20828,N_19343,N_19400);
and U20829 (N_20829,N_19290,N_17524);
or U20830 (N_20830,N_19411,N_19271);
nand U20831 (N_20831,N_19520,N_19888);
nand U20832 (N_20832,N_19005,N_19259);
xor U20833 (N_20833,N_18645,N_17913);
or U20834 (N_20834,N_17846,N_18291);
nor U20835 (N_20835,N_17947,N_18380);
xnor U20836 (N_20836,N_19084,N_19487);
or U20837 (N_20837,N_18015,N_19928);
nor U20838 (N_20838,N_19884,N_18817);
and U20839 (N_20839,N_19329,N_19822);
and U20840 (N_20840,N_17813,N_17789);
xor U20841 (N_20841,N_17545,N_17978);
xor U20842 (N_20842,N_19086,N_18312);
nor U20843 (N_20843,N_17689,N_19286);
or U20844 (N_20844,N_19110,N_19824);
or U20845 (N_20845,N_17520,N_17505);
xor U20846 (N_20846,N_19705,N_19967);
xnor U20847 (N_20847,N_17646,N_19338);
and U20848 (N_20848,N_17615,N_19042);
nand U20849 (N_20849,N_17829,N_19556);
nand U20850 (N_20850,N_19690,N_17954);
xnor U20851 (N_20851,N_19498,N_17871);
and U20852 (N_20852,N_17930,N_18074);
nand U20853 (N_20853,N_19717,N_17848);
nor U20854 (N_20854,N_17613,N_19202);
or U20855 (N_20855,N_19615,N_19545);
nand U20856 (N_20856,N_19623,N_19780);
xnor U20857 (N_20857,N_17805,N_19773);
xnor U20858 (N_20858,N_17723,N_19654);
and U20859 (N_20859,N_19177,N_18174);
and U20860 (N_20860,N_17720,N_19629);
and U20861 (N_20861,N_18841,N_18191);
and U20862 (N_20862,N_18694,N_19641);
nor U20863 (N_20863,N_19043,N_17823);
or U20864 (N_20864,N_19081,N_19934);
and U20865 (N_20865,N_19774,N_18355);
xnor U20866 (N_20866,N_18051,N_17828);
nand U20867 (N_20867,N_19983,N_18913);
xor U20868 (N_20868,N_18657,N_18444);
nand U20869 (N_20869,N_18574,N_18813);
nand U20870 (N_20870,N_17516,N_17656);
nand U20871 (N_20871,N_18301,N_18562);
nor U20872 (N_20872,N_17977,N_17861);
nand U20873 (N_20873,N_17850,N_18110);
nand U20874 (N_20874,N_18563,N_19077);
nand U20875 (N_20875,N_18825,N_18107);
or U20876 (N_20876,N_18111,N_19758);
nand U20877 (N_20877,N_19872,N_17778);
nand U20878 (N_20878,N_19306,N_18133);
nor U20879 (N_20879,N_19710,N_17739);
or U20880 (N_20880,N_19420,N_19366);
and U20881 (N_20881,N_18516,N_19878);
and U20882 (N_20882,N_18819,N_18866);
and U20883 (N_20883,N_17522,N_17810);
and U20884 (N_20884,N_18709,N_18763);
nand U20885 (N_20885,N_19065,N_18089);
nand U20886 (N_20886,N_18280,N_19829);
nand U20887 (N_20887,N_17895,N_18587);
or U20888 (N_20888,N_18625,N_19324);
or U20889 (N_20889,N_19843,N_17817);
or U20890 (N_20890,N_17608,N_17797);
nor U20891 (N_20891,N_17989,N_19314);
and U20892 (N_20892,N_18546,N_17548);
or U20893 (N_20893,N_18767,N_19032);
nor U20894 (N_20894,N_18346,N_19341);
xor U20895 (N_20895,N_19070,N_18774);
xnor U20896 (N_20896,N_18398,N_18662);
or U20897 (N_20897,N_17802,N_19720);
nand U20898 (N_20898,N_18967,N_18751);
or U20899 (N_20899,N_19417,N_17645);
nor U20900 (N_20900,N_18093,N_18014);
nor U20901 (N_20901,N_18707,N_19002);
nor U20902 (N_20902,N_18370,N_17628);
nand U20903 (N_20903,N_17531,N_17624);
xnor U20904 (N_20904,N_17836,N_18101);
nand U20905 (N_20905,N_19911,N_18032);
nand U20906 (N_20906,N_19716,N_19782);
nand U20907 (N_20907,N_19475,N_18855);
nand U20908 (N_20908,N_18942,N_19954);
xor U20909 (N_20909,N_19536,N_17970);
and U20910 (N_20910,N_19381,N_18040);
nor U20911 (N_20911,N_19703,N_19775);
nand U20912 (N_20912,N_17502,N_18883);
or U20913 (N_20913,N_19544,N_19719);
nor U20914 (N_20914,N_19100,N_18259);
or U20915 (N_20915,N_19031,N_18011);
xnor U20916 (N_20916,N_17620,N_18377);
and U20917 (N_20917,N_18595,N_19496);
or U20918 (N_20918,N_19834,N_19468);
nand U20919 (N_20919,N_18754,N_19547);
nand U20920 (N_20920,N_17855,N_19747);
xor U20921 (N_20921,N_19358,N_18248);
and U20922 (N_20922,N_19467,N_18360);
nor U20923 (N_20923,N_19818,N_19245);
or U20924 (N_20924,N_18071,N_18117);
nand U20925 (N_20925,N_19447,N_19831);
or U20926 (N_20926,N_17566,N_18632);
xor U20927 (N_20927,N_18644,N_17565);
and U20928 (N_20928,N_19033,N_19170);
xor U20929 (N_20929,N_18950,N_19985);
or U20930 (N_20930,N_19930,N_18390);
nand U20931 (N_20931,N_18919,N_19754);
nor U20932 (N_20932,N_19619,N_18332);
nand U20933 (N_20933,N_18589,N_18672);
nand U20934 (N_20934,N_19216,N_19951);
nor U20935 (N_20935,N_18615,N_18965);
or U20936 (N_20936,N_19530,N_18903);
nand U20937 (N_20937,N_17515,N_18703);
nand U20938 (N_20938,N_18669,N_19455);
xor U20939 (N_20939,N_19348,N_18314);
xnor U20940 (N_20940,N_18831,N_17779);
or U20941 (N_20941,N_17774,N_18495);
nor U20942 (N_20942,N_19224,N_19694);
nand U20943 (N_20943,N_17955,N_19573);
and U20944 (N_20944,N_19205,N_17859);
or U20945 (N_20945,N_19617,N_17715);
or U20946 (N_20946,N_18656,N_17673);
and U20947 (N_20947,N_19886,N_17845);
xor U20948 (N_20948,N_19409,N_19407);
nand U20949 (N_20949,N_17940,N_18986);
or U20950 (N_20950,N_19184,N_19062);
nor U20951 (N_20951,N_17716,N_18474);
xor U20952 (N_20952,N_19914,N_18551);
or U20953 (N_20953,N_17981,N_19522);
nor U20954 (N_20954,N_18118,N_18604);
and U20955 (N_20955,N_18461,N_19122);
xor U20956 (N_20956,N_18201,N_18404);
and U20957 (N_20957,N_19639,N_17866);
nor U20958 (N_20958,N_19870,N_17592);
or U20959 (N_20959,N_18323,N_19725);
or U20960 (N_20960,N_19542,N_19618);
xnor U20961 (N_20961,N_17979,N_19605);
or U20962 (N_20962,N_19434,N_18651);
or U20963 (N_20963,N_19429,N_19746);
nand U20964 (N_20964,N_19801,N_19064);
or U20965 (N_20965,N_19129,N_18262);
or U20966 (N_20966,N_18583,N_17575);
and U20967 (N_20967,N_19059,N_18344);
and U20968 (N_20968,N_18566,N_17951);
nand U20969 (N_20969,N_19211,N_18637);
or U20970 (N_20970,N_19295,N_17884);
or U20971 (N_20971,N_19810,N_18613);
nand U20972 (N_20972,N_17643,N_19344);
or U20973 (N_20973,N_18034,N_17996);
xnor U20974 (N_20974,N_19590,N_18624);
nor U20975 (N_20975,N_18436,N_17598);
and U20976 (N_20976,N_19939,N_18670);
and U20977 (N_20977,N_19790,N_19332);
nor U20978 (N_20978,N_18189,N_18537);
or U20979 (N_20979,N_19823,N_18269);
nand U20980 (N_20980,N_19895,N_18530);
and U20981 (N_20981,N_18954,N_18038);
nand U20982 (N_20982,N_18654,N_18388);
xor U20983 (N_20983,N_19500,N_17952);
and U20984 (N_20984,N_19594,N_19426);
xor U20985 (N_20985,N_19770,N_19051);
xor U20986 (N_20986,N_18610,N_19737);
xor U20987 (N_20987,N_17551,N_18004);
xor U20988 (N_20988,N_18027,N_19635);
or U20989 (N_20989,N_17582,N_17530);
nand U20990 (N_20990,N_19931,N_17995);
and U20991 (N_20991,N_19103,N_17742);
nand U20992 (N_20992,N_19597,N_17538);
or U20993 (N_20993,N_19772,N_19135);
and U20994 (N_20994,N_17668,N_18534);
xnor U20995 (N_20995,N_17890,N_19313);
nand U20996 (N_20996,N_19356,N_19242);
xor U20997 (N_20997,N_18796,N_19534);
xnor U20998 (N_20998,N_18431,N_19568);
nor U20999 (N_20999,N_19471,N_17602);
and U21000 (N_21000,N_19370,N_17667);
nor U21001 (N_21001,N_18734,N_19156);
nor U21002 (N_21002,N_19797,N_18714);
and U21003 (N_21003,N_18375,N_19789);
nand U21004 (N_21004,N_19473,N_18922);
nand U21005 (N_21005,N_19418,N_18396);
or U21006 (N_21006,N_19874,N_18418);
nand U21007 (N_21007,N_18827,N_17501);
nor U21008 (N_21008,N_19866,N_18558);
or U21009 (N_21009,N_17796,N_19687);
and U21010 (N_21010,N_18367,N_19294);
and U21011 (N_21011,N_18902,N_19958);
and U21012 (N_21012,N_19962,N_19132);
xnor U21013 (N_21013,N_19942,N_19111);
nand U21014 (N_21014,N_18419,N_18309);
xor U21015 (N_21015,N_19327,N_19074);
and U21016 (N_21016,N_17973,N_19427);
xor U21017 (N_21017,N_19783,N_19645);
xnor U21018 (N_21018,N_19686,N_18239);
and U21019 (N_21019,N_18350,N_17830);
and U21020 (N_21020,N_18278,N_19913);
nor U21021 (N_21021,N_19351,N_17674);
and U21022 (N_21022,N_18800,N_19625);
nand U21023 (N_21023,N_18379,N_19927);
nand U21024 (N_21024,N_18968,N_17661);
nand U21025 (N_21025,N_19970,N_19357);
nand U21026 (N_21026,N_18633,N_19445);
nand U21027 (N_21027,N_18994,N_17535);
nor U21028 (N_21028,N_19640,N_17957);
nand U21029 (N_21029,N_18803,N_18971);
xor U21030 (N_21030,N_18018,N_18893);
or U21031 (N_21031,N_19892,N_17707);
and U21032 (N_21032,N_17540,N_18195);
nand U21033 (N_21033,N_18955,N_17663);
nand U21034 (N_21034,N_18438,N_19119);
xor U21035 (N_21035,N_18728,N_17921);
nand U21036 (N_21036,N_19541,N_17868);
nand U21037 (N_21037,N_18691,N_18879);
and U21038 (N_21038,N_19532,N_17687);
and U21039 (N_21039,N_19864,N_18935);
nor U21040 (N_21040,N_19921,N_17711);
nand U21041 (N_21041,N_19133,N_18306);
or U21042 (N_21042,N_18485,N_18598);
or U21043 (N_21043,N_19642,N_18712);
and U21044 (N_21044,N_18180,N_18764);
and U21045 (N_21045,N_17634,N_18376);
xor U21046 (N_21046,N_17552,N_17926);
and U21047 (N_21047,N_19006,N_18243);
nor U21048 (N_21048,N_17737,N_18373);
nor U21049 (N_21049,N_19027,N_19340);
or U21050 (N_21050,N_19377,N_18742);
xor U21051 (N_21051,N_18646,N_18768);
and U21052 (N_21052,N_18284,N_19432);
and U21053 (N_21053,N_18784,N_17706);
and U21054 (N_21054,N_18766,N_18931);
xor U21055 (N_21055,N_18533,N_18519);
or U21056 (N_21056,N_19350,N_17576);
or U21057 (N_21057,N_18704,N_17843);
xor U21058 (N_21058,N_19529,N_19012);
or U21059 (N_21059,N_19777,N_19481);
nor U21060 (N_21060,N_18414,N_19662);
and U21061 (N_21061,N_19168,N_18901);
nand U21062 (N_21062,N_18730,N_18187);
nand U21063 (N_21063,N_18279,N_18082);
nand U21064 (N_21064,N_19505,N_17763);
nand U21065 (N_21065,N_18468,N_18561);
xnor U21066 (N_21066,N_18342,N_18241);
xnor U21067 (N_21067,N_18794,N_18152);
xor U21068 (N_21068,N_18719,N_18488);
or U21069 (N_21069,N_19727,N_19940);
xor U21070 (N_21070,N_18652,N_19627);
or U21071 (N_21071,N_18167,N_18251);
and U21072 (N_21072,N_18416,N_18159);
nor U21073 (N_21073,N_18289,N_18389);
or U21074 (N_21074,N_18747,N_18857);
or U21075 (N_21075,N_18858,N_17541);
or U21076 (N_21076,N_18991,N_19109);
or U21077 (N_21077,N_19850,N_17563);
or U21078 (N_21078,N_17839,N_19139);
xnor U21079 (N_21079,N_18835,N_18987);
nor U21080 (N_21080,N_18979,N_19599);
and U21081 (N_21081,N_18708,N_19566);
or U21082 (N_21082,N_19918,N_18401);
nor U21083 (N_21083,N_19688,N_18975);
nand U21084 (N_21084,N_17549,N_18339);
and U21085 (N_21085,N_19508,N_19425);
nand U21086 (N_21086,N_17987,N_19993);
or U21087 (N_21087,N_18228,N_19673);
nor U21088 (N_21088,N_18518,N_18240);
or U21089 (N_21089,N_18094,N_19010);
or U21090 (N_21090,N_18513,N_19095);
xor U21091 (N_21091,N_19709,N_18105);
nand U21092 (N_21092,N_18560,N_18823);
and U21093 (N_21093,N_18399,N_17743);
and U21094 (N_21094,N_18382,N_19819);
xnor U21095 (N_21095,N_18852,N_18408);
nor U21096 (N_21096,N_19636,N_18304);
nand U21097 (N_21097,N_19909,N_17606);
xnor U21098 (N_21098,N_17611,N_17912);
and U21099 (N_21099,N_17533,N_18896);
or U21100 (N_21100,N_18385,N_19998);
or U21101 (N_21101,N_18020,N_17893);
or U21102 (N_21102,N_18114,N_19317);
or U21103 (N_21103,N_19234,N_18929);
and U21104 (N_21104,N_18198,N_19020);
xor U21105 (N_21105,N_19821,N_18026);
xor U21106 (N_21106,N_18710,N_19861);
nor U21107 (N_21107,N_18112,N_19116);
xnor U21108 (N_21108,N_18860,N_19478);
xor U21109 (N_21109,N_19171,N_17591);
or U21110 (N_21110,N_18932,N_19217);
or U21111 (N_21111,N_19684,N_19842);
or U21112 (N_21112,N_19634,N_17697);
or U21113 (N_21113,N_18406,N_19769);
or U21114 (N_21114,N_19457,N_18063);
or U21115 (N_21115,N_18702,N_19846);
nor U21116 (N_21116,N_19751,N_18553);
or U21117 (N_21117,N_19384,N_18801);
nor U21118 (N_21118,N_17882,N_19123);
or U21119 (N_21119,N_18711,N_18449);
or U21120 (N_21120,N_18772,N_19830);
or U21121 (N_21121,N_19303,N_19276);
and U21122 (N_21122,N_17671,N_18705);
nand U21123 (N_21123,N_18853,N_19213);
nand U21124 (N_21124,N_18720,N_17701);
xnor U21125 (N_21125,N_17719,N_19611);
nand U21126 (N_21126,N_19389,N_17729);
xnor U21127 (N_21127,N_19283,N_17833);
and U21128 (N_21128,N_19278,N_17721);
or U21129 (N_21129,N_19151,N_19054);
nand U21130 (N_21130,N_18258,N_17923);
xor U21131 (N_21131,N_17696,N_19665);
or U21132 (N_21132,N_18789,N_19925);
nand U21133 (N_21133,N_18579,N_18430);
or U21134 (N_21134,N_19339,N_18505);
and U21135 (N_21135,N_18148,N_19137);
xor U21136 (N_21136,N_18294,N_18030);
or U21137 (N_21137,N_18531,N_18805);
or U21138 (N_21138,N_18352,N_17925);
and U21139 (N_21139,N_18843,N_19503);
nand U21140 (N_21140,N_19602,N_17635);
nand U21141 (N_21141,N_19186,N_19875);
or U21142 (N_21142,N_18678,N_19255);
and U21143 (N_21143,N_17786,N_19265);
nand U21144 (N_21144,N_17612,N_17585);
nand U21145 (N_21145,N_17649,N_18834);
nand U21146 (N_21146,N_18447,N_17730);
or U21147 (N_21147,N_19479,N_19723);
and U21148 (N_21148,N_18395,N_19664);
or U21149 (N_21149,N_19670,N_18820);
nor U21150 (N_21150,N_18432,N_18863);
or U21151 (N_21151,N_19708,N_17700);
xnor U21152 (N_21152,N_19608,N_18663);
and U21153 (N_21153,N_18088,N_18886);
and U21154 (N_21154,N_18437,N_17605);
xnor U21155 (N_21155,N_19353,N_17792);
xnor U21156 (N_21156,N_17609,N_17601);
nor U21157 (N_21157,N_17918,N_17503);
and U21158 (N_21158,N_17961,N_17946);
or U21159 (N_21159,N_17904,N_18630);
xnor U21160 (N_21160,N_18087,N_18393);
xnor U21161 (N_21161,N_19436,N_17556);
nand U21162 (N_21162,N_18273,N_18753);
xor U21163 (N_21163,N_19352,N_19713);
nand U21164 (N_21164,N_18964,N_18207);
nor U21165 (N_21165,N_18300,N_18628);
nand U21166 (N_21166,N_17816,N_18830);
and U21167 (N_21167,N_18552,N_18424);
nor U21168 (N_21168,N_19248,N_18526);
nand U21169 (N_21169,N_18372,N_19105);
nand U21170 (N_21170,N_19152,N_19113);
and U21171 (N_21171,N_18514,N_17901);
nor U21172 (N_21172,N_18802,N_18748);
and U21173 (N_21173,N_18815,N_19908);
or U21174 (N_21174,N_19403,N_19378);
nor U21175 (N_21175,N_19442,N_18146);
nand U21176 (N_21176,N_18592,N_19644);
or U21177 (N_21177,N_18433,N_19743);
or U21178 (N_21178,N_17660,N_18911);
nand U21179 (N_21179,N_19285,N_18701);
nor U21180 (N_21180,N_19828,N_18450);
nor U21181 (N_21181,N_17675,N_18095);
and U21182 (N_21182,N_17755,N_17543);
xnor U21183 (N_21183,N_17642,N_19218);
nand U21184 (N_21184,N_17907,N_17999);
nand U21185 (N_21185,N_18318,N_19799);
and U21186 (N_21186,N_19633,N_18482);
xor U21187 (N_21187,N_18378,N_18031);
xor U21188 (N_21188,N_17542,N_17902);
xor U21189 (N_21189,N_19552,N_18102);
or U21190 (N_21190,N_19826,N_18928);
nand U21191 (N_21191,N_19085,N_18778);
or U21192 (N_21192,N_18792,N_17983);
nand U21193 (N_21193,N_19550,N_19961);
nand U21194 (N_21194,N_19241,N_18194);
nor U21195 (N_21195,N_19214,N_18387);
or U21196 (N_21196,N_19963,N_19638);
or U21197 (N_21197,N_19421,N_19146);
xnor U21198 (N_21198,N_19793,N_19804);
or U21199 (N_21199,N_19334,N_19336);
xor U21200 (N_21200,N_19094,N_19013);
xor U21201 (N_21201,N_19435,N_19988);
and U21202 (N_21202,N_19015,N_17733);
or U21203 (N_21203,N_19994,N_17762);
xor U21204 (N_21204,N_17988,N_19742);
xnor U21205 (N_21205,N_18999,N_17814);
nand U21206 (N_21206,N_18992,N_18229);
nor U21207 (N_21207,N_18354,N_18888);
nand U21208 (N_21208,N_17519,N_17969);
xnor U21209 (N_21209,N_19981,N_19579);
nor U21210 (N_21210,N_18790,N_17852);
or U21211 (N_21211,N_18173,N_18572);
nand U21212 (N_21212,N_19288,N_18868);
and U21213 (N_21213,N_19651,N_18085);
nand U21214 (N_21214,N_19284,N_17666);
nand U21215 (N_21215,N_17748,N_19386);
nand U21216 (N_21216,N_18515,N_18068);
xnor U21217 (N_21217,N_19203,N_17627);
and U21218 (N_21218,N_17590,N_18320);
nand U21219 (N_21219,N_18293,N_19472);
and U21220 (N_21220,N_18489,N_19066);
or U21221 (N_21221,N_19660,N_18554);
xnor U21222 (N_21222,N_19912,N_18674);
and U21223 (N_21223,N_19848,N_18206);
and U21224 (N_21224,N_19009,N_18204);
xor U21225 (N_21225,N_19554,N_19422);
and U21226 (N_21226,N_18564,N_19779);
nand U21227 (N_21227,N_19571,N_17583);
nor U21228 (N_21228,N_19189,N_19730);
nor U21229 (N_21229,N_18980,N_19365);
or U21230 (N_21230,N_17886,N_18512);
xnor U21231 (N_21231,N_18463,N_17888);
nand U21232 (N_21232,N_18137,N_18451);
and U21233 (N_21233,N_19261,N_19570);
or U21234 (N_21234,N_18498,N_18400);
xnor U21235 (N_21235,N_19155,N_19376);
nand U21236 (N_21236,N_18659,N_19784);
nand U21237 (N_21237,N_18966,N_17724);
xnor U21238 (N_21238,N_19858,N_18666);
xnor U21239 (N_21239,N_17857,N_18616);
xor U21240 (N_21240,N_19584,N_17579);
xor U21241 (N_21241,N_19459,N_18811);
and U21242 (N_21242,N_19649,N_19748);
xnor U21243 (N_21243,N_18022,N_18083);
and U21244 (N_21244,N_19669,N_19347);
or U21245 (N_21245,N_18529,N_19167);
and U21246 (N_21246,N_18900,N_18080);
nand U21247 (N_21247,N_18122,N_17636);
xor U21248 (N_21248,N_18732,N_17770);
or U21249 (N_21249,N_18773,N_19367);
or U21250 (N_21250,N_18254,N_19735);
xor U21251 (N_21251,N_19101,N_19529);
xor U21252 (N_21252,N_18304,N_18030);
xnor U21253 (N_21253,N_18216,N_17952);
or U21254 (N_21254,N_19981,N_19761);
nor U21255 (N_21255,N_19076,N_17756);
nor U21256 (N_21256,N_17956,N_17756);
and U21257 (N_21257,N_18757,N_18932);
nor U21258 (N_21258,N_19275,N_17604);
nor U21259 (N_21259,N_19328,N_18720);
and U21260 (N_21260,N_18133,N_19189);
or U21261 (N_21261,N_18485,N_17530);
nand U21262 (N_21262,N_17984,N_19208);
xor U21263 (N_21263,N_19027,N_18152);
and U21264 (N_21264,N_17734,N_18789);
or U21265 (N_21265,N_18935,N_19035);
nand U21266 (N_21266,N_17861,N_19821);
and U21267 (N_21267,N_19640,N_18690);
nand U21268 (N_21268,N_19264,N_19413);
nand U21269 (N_21269,N_18205,N_19558);
and U21270 (N_21270,N_18846,N_18968);
xnor U21271 (N_21271,N_17928,N_18730);
and U21272 (N_21272,N_19571,N_18452);
nor U21273 (N_21273,N_18349,N_17648);
or U21274 (N_21274,N_18051,N_18264);
or U21275 (N_21275,N_19570,N_19482);
xor U21276 (N_21276,N_19257,N_18641);
and U21277 (N_21277,N_19104,N_19979);
nand U21278 (N_21278,N_18545,N_18009);
xor U21279 (N_21279,N_19583,N_19687);
nor U21280 (N_21280,N_18639,N_19991);
xor U21281 (N_21281,N_19334,N_19129);
and U21282 (N_21282,N_18609,N_18877);
nor U21283 (N_21283,N_19327,N_17531);
or U21284 (N_21284,N_19483,N_19272);
xor U21285 (N_21285,N_19535,N_18637);
nor U21286 (N_21286,N_18177,N_17697);
nand U21287 (N_21287,N_18402,N_19015);
and U21288 (N_21288,N_17509,N_18884);
nor U21289 (N_21289,N_18018,N_17912);
and U21290 (N_21290,N_18247,N_18553);
or U21291 (N_21291,N_17603,N_18553);
and U21292 (N_21292,N_18807,N_18520);
nor U21293 (N_21293,N_19496,N_17855);
nor U21294 (N_21294,N_19277,N_17779);
and U21295 (N_21295,N_19667,N_19090);
nand U21296 (N_21296,N_18571,N_18484);
nor U21297 (N_21297,N_18399,N_17990);
and U21298 (N_21298,N_19393,N_19855);
and U21299 (N_21299,N_18855,N_19187);
xor U21300 (N_21300,N_17944,N_18395);
or U21301 (N_21301,N_19913,N_19896);
or U21302 (N_21302,N_18281,N_19458);
nand U21303 (N_21303,N_18242,N_19009);
nand U21304 (N_21304,N_17945,N_19623);
nor U21305 (N_21305,N_18291,N_19164);
nor U21306 (N_21306,N_18152,N_19365);
and U21307 (N_21307,N_19647,N_17998);
nand U21308 (N_21308,N_17971,N_18555);
xnor U21309 (N_21309,N_18797,N_19100);
nand U21310 (N_21310,N_19478,N_19786);
xor U21311 (N_21311,N_17981,N_18697);
nand U21312 (N_21312,N_18355,N_19869);
nand U21313 (N_21313,N_19025,N_17988);
and U21314 (N_21314,N_19793,N_18798);
nor U21315 (N_21315,N_19820,N_18817);
xor U21316 (N_21316,N_17739,N_18849);
xor U21317 (N_21317,N_18574,N_18758);
or U21318 (N_21318,N_17766,N_18563);
nor U21319 (N_21319,N_18649,N_18318);
nor U21320 (N_21320,N_17875,N_18693);
xor U21321 (N_21321,N_18918,N_17813);
xor U21322 (N_21322,N_18473,N_18388);
nand U21323 (N_21323,N_18773,N_19298);
and U21324 (N_21324,N_18118,N_19530);
or U21325 (N_21325,N_19201,N_18509);
or U21326 (N_21326,N_17783,N_18942);
and U21327 (N_21327,N_17716,N_19929);
nor U21328 (N_21328,N_19667,N_17932);
and U21329 (N_21329,N_18083,N_19181);
nor U21330 (N_21330,N_18463,N_18619);
or U21331 (N_21331,N_17566,N_18643);
nand U21332 (N_21332,N_18924,N_17653);
xor U21333 (N_21333,N_19218,N_19163);
xor U21334 (N_21334,N_17896,N_18774);
nor U21335 (N_21335,N_18839,N_18334);
and U21336 (N_21336,N_18442,N_19283);
and U21337 (N_21337,N_19578,N_19020);
nor U21338 (N_21338,N_18219,N_18657);
xnor U21339 (N_21339,N_18980,N_17787);
or U21340 (N_21340,N_18653,N_17775);
xnor U21341 (N_21341,N_19697,N_17754);
or U21342 (N_21342,N_18184,N_19140);
nand U21343 (N_21343,N_19584,N_18502);
nand U21344 (N_21344,N_19859,N_17895);
or U21345 (N_21345,N_19118,N_17947);
and U21346 (N_21346,N_19737,N_19560);
nand U21347 (N_21347,N_18183,N_19569);
nand U21348 (N_21348,N_19607,N_19117);
and U21349 (N_21349,N_18808,N_18068);
nor U21350 (N_21350,N_17829,N_18302);
nand U21351 (N_21351,N_18182,N_19425);
xor U21352 (N_21352,N_19970,N_17794);
nor U21353 (N_21353,N_18112,N_18515);
or U21354 (N_21354,N_17910,N_18262);
xor U21355 (N_21355,N_19671,N_19293);
nand U21356 (N_21356,N_19374,N_18577);
or U21357 (N_21357,N_19358,N_18010);
nand U21358 (N_21358,N_19934,N_19156);
and U21359 (N_21359,N_19950,N_18434);
and U21360 (N_21360,N_17873,N_17819);
nand U21361 (N_21361,N_18976,N_19925);
nand U21362 (N_21362,N_18370,N_19141);
xor U21363 (N_21363,N_18027,N_18359);
and U21364 (N_21364,N_18800,N_19969);
or U21365 (N_21365,N_17876,N_19223);
nand U21366 (N_21366,N_18899,N_19652);
xnor U21367 (N_21367,N_19314,N_18940);
and U21368 (N_21368,N_17651,N_19441);
nand U21369 (N_21369,N_18925,N_18900);
and U21370 (N_21370,N_17574,N_18358);
nand U21371 (N_21371,N_18815,N_18759);
and U21372 (N_21372,N_18035,N_19325);
xor U21373 (N_21373,N_19072,N_19532);
nor U21374 (N_21374,N_19984,N_19942);
and U21375 (N_21375,N_17884,N_19873);
or U21376 (N_21376,N_19628,N_19516);
and U21377 (N_21377,N_17905,N_17864);
nor U21378 (N_21378,N_17748,N_19637);
or U21379 (N_21379,N_19202,N_18845);
nor U21380 (N_21380,N_19941,N_18958);
or U21381 (N_21381,N_17839,N_19141);
or U21382 (N_21382,N_19003,N_18820);
nand U21383 (N_21383,N_19690,N_18240);
nor U21384 (N_21384,N_19819,N_18372);
xnor U21385 (N_21385,N_18766,N_19436);
xor U21386 (N_21386,N_19523,N_19063);
nand U21387 (N_21387,N_19585,N_18972);
nor U21388 (N_21388,N_18959,N_19628);
or U21389 (N_21389,N_18097,N_19298);
nor U21390 (N_21390,N_19960,N_18154);
nor U21391 (N_21391,N_19861,N_19787);
or U21392 (N_21392,N_17934,N_18729);
or U21393 (N_21393,N_19210,N_18312);
nand U21394 (N_21394,N_18241,N_18264);
xor U21395 (N_21395,N_19276,N_18140);
xnor U21396 (N_21396,N_19917,N_18425);
and U21397 (N_21397,N_17664,N_19338);
and U21398 (N_21398,N_17847,N_19533);
nor U21399 (N_21399,N_19120,N_18292);
or U21400 (N_21400,N_19450,N_17764);
nor U21401 (N_21401,N_18158,N_18469);
and U21402 (N_21402,N_18086,N_19692);
nand U21403 (N_21403,N_17955,N_18996);
nand U21404 (N_21404,N_19065,N_19882);
nand U21405 (N_21405,N_18067,N_18220);
and U21406 (N_21406,N_18840,N_18352);
and U21407 (N_21407,N_18244,N_17699);
and U21408 (N_21408,N_19937,N_18756);
or U21409 (N_21409,N_19622,N_18131);
and U21410 (N_21410,N_19364,N_19432);
and U21411 (N_21411,N_19475,N_18342);
nor U21412 (N_21412,N_17866,N_19102);
or U21413 (N_21413,N_19236,N_19092);
and U21414 (N_21414,N_19501,N_17718);
xor U21415 (N_21415,N_18306,N_19271);
nand U21416 (N_21416,N_19447,N_17512);
xnor U21417 (N_21417,N_18538,N_19712);
nor U21418 (N_21418,N_19010,N_19977);
nand U21419 (N_21419,N_19454,N_19608);
or U21420 (N_21420,N_17519,N_17708);
or U21421 (N_21421,N_18994,N_18744);
or U21422 (N_21422,N_19127,N_19740);
xor U21423 (N_21423,N_19292,N_18316);
or U21424 (N_21424,N_17972,N_18838);
and U21425 (N_21425,N_18797,N_17596);
and U21426 (N_21426,N_19873,N_19673);
nor U21427 (N_21427,N_18488,N_19422);
or U21428 (N_21428,N_18169,N_19207);
and U21429 (N_21429,N_18168,N_18323);
nor U21430 (N_21430,N_19560,N_18351);
xnor U21431 (N_21431,N_17847,N_18380);
nand U21432 (N_21432,N_18767,N_18580);
xnor U21433 (N_21433,N_17920,N_19930);
and U21434 (N_21434,N_18297,N_18541);
or U21435 (N_21435,N_18476,N_18693);
or U21436 (N_21436,N_17630,N_18776);
xor U21437 (N_21437,N_18419,N_18195);
xnor U21438 (N_21438,N_19293,N_19049);
nand U21439 (N_21439,N_18672,N_19911);
and U21440 (N_21440,N_17756,N_18320);
and U21441 (N_21441,N_18906,N_18484);
or U21442 (N_21442,N_17600,N_19257);
and U21443 (N_21443,N_17833,N_18461);
nor U21444 (N_21444,N_19656,N_17965);
xor U21445 (N_21445,N_18382,N_18848);
nand U21446 (N_21446,N_19371,N_18369);
xor U21447 (N_21447,N_18066,N_19991);
xor U21448 (N_21448,N_18463,N_18656);
nor U21449 (N_21449,N_19864,N_18278);
xor U21450 (N_21450,N_18565,N_18930);
xnor U21451 (N_21451,N_18977,N_17920);
or U21452 (N_21452,N_19032,N_19072);
nand U21453 (N_21453,N_19564,N_18355);
or U21454 (N_21454,N_18754,N_17831);
or U21455 (N_21455,N_18172,N_18376);
nand U21456 (N_21456,N_19895,N_18585);
and U21457 (N_21457,N_19357,N_18247);
or U21458 (N_21458,N_19899,N_18601);
xnor U21459 (N_21459,N_17633,N_19790);
nand U21460 (N_21460,N_17725,N_17734);
xor U21461 (N_21461,N_17625,N_18508);
or U21462 (N_21462,N_18189,N_18252);
xnor U21463 (N_21463,N_19671,N_19460);
or U21464 (N_21464,N_17809,N_18661);
nor U21465 (N_21465,N_19586,N_18389);
and U21466 (N_21466,N_18657,N_19637);
and U21467 (N_21467,N_18655,N_17589);
nand U21468 (N_21468,N_18648,N_19018);
nor U21469 (N_21469,N_17659,N_19658);
xor U21470 (N_21470,N_19165,N_18635);
or U21471 (N_21471,N_19680,N_18276);
nor U21472 (N_21472,N_19436,N_17696);
and U21473 (N_21473,N_19831,N_17639);
xor U21474 (N_21474,N_19706,N_19293);
nand U21475 (N_21475,N_19451,N_17958);
and U21476 (N_21476,N_18782,N_18323);
and U21477 (N_21477,N_19603,N_19102);
nor U21478 (N_21478,N_19147,N_18515);
and U21479 (N_21479,N_18707,N_19757);
or U21480 (N_21480,N_18927,N_19684);
xor U21481 (N_21481,N_18365,N_18800);
xor U21482 (N_21482,N_18790,N_18346);
nor U21483 (N_21483,N_18899,N_18512);
nor U21484 (N_21484,N_18892,N_19324);
and U21485 (N_21485,N_17798,N_19359);
nor U21486 (N_21486,N_17961,N_18112);
or U21487 (N_21487,N_19810,N_19496);
xnor U21488 (N_21488,N_19183,N_18651);
or U21489 (N_21489,N_18080,N_19057);
xnor U21490 (N_21490,N_18394,N_18665);
nand U21491 (N_21491,N_18619,N_18151);
or U21492 (N_21492,N_18700,N_18881);
xor U21493 (N_21493,N_19076,N_18277);
and U21494 (N_21494,N_19526,N_18368);
nor U21495 (N_21495,N_19008,N_19341);
xnor U21496 (N_21496,N_18273,N_17825);
nand U21497 (N_21497,N_17668,N_18969);
xor U21498 (N_21498,N_18835,N_19530);
and U21499 (N_21499,N_17588,N_19215);
or U21500 (N_21500,N_19142,N_18823);
nand U21501 (N_21501,N_17938,N_19492);
or U21502 (N_21502,N_18999,N_19523);
and U21503 (N_21503,N_19869,N_18142);
nor U21504 (N_21504,N_19539,N_18395);
nand U21505 (N_21505,N_17711,N_18195);
xor U21506 (N_21506,N_17538,N_18460);
xnor U21507 (N_21507,N_19608,N_18083);
nor U21508 (N_21508,N_17754,N_17624);
xor U21509 (N_21509,N_19367,N_17915);
xor U21510 (N_21510,N_19774,N_17750);
nand U21511 (N_21511,N_17818,N_17588);
xor U21512 (N_21512,N_19980,N_17830);
nand U21513 (N_21513,N_18153,N_19182);
nor U21514 (N_21514,N_19561,N_19686);
nor U21515 (N_21515,N_17814,N_17509);
or U21516 (N_21516,N_18932,N_18939);
nor U21517 (N_21517,N_18327,N_19494);
and U21518 (N_21518,N_19479,N_18770);
xnor U21519 (N_21519,N_18684,N_19720);
xnor U21520 (N_21520,N_18590,N_18342);
or U21521 (N_21521,N_19333,N_18167);
nand U21522 (N_21522,N_19047,N_19139);
xnor U21523 (N_21523,N_18784,N_18464);
xor U21524 (N_21524,N_19638,N_19618);
nand U21525 (N_21525,N_19036,N_18664);
xor U21526 (N_21526,N_18918,N_19614);
or U21527 (N_21527,N_19048,N_18986);
or U21528 (N_21528,N_18031,N_17975);
or U21529 (N_21529,N_17534,N_17644);
or U21530 (N_21530,N_18010,N_19802);
and U21531 (N_21531,N_18307,N_18339);
and U21532 (N_21532,N_18010,N_17715);
xnor U21533 (N_21533,N_19153,N_18968);
nand U21534 (N_21534,N_18353,N_19313);
nor U21535 (N_21535,N_17673,N_19863);
nand U21536 (N_21536,N_18233,N_19475);
xnor U21537 (N_21537,N_19618,N_18333);
nor U21538 (N_21538,N_19466,N_19409);
xnor U21539 (N_21539,N_19336,N_18492);
xnor U21540 (N_21540,N_18225,N_18457);
nand U21541 (N_21541,N_19508,N_19075);
nor U21542 (N_21542,N_19257,N_18116);
xor U21543 (N_21543,N_17834,N_19473);
nand U21544 (N_21544,N_18251,N_19929);
xor U21545 (N_21545,N_18920,N_19885);
nand U21546 (N_21546,N_19494,N_18735);
and U21547 (N_21547,N_19439,N_17651);
and U21548 (N_21548,N_18552,N_19079);
xor U21549 (N_21549,N_18319,N_17888);
nand U21550 (N_21550,N_18059,N_18720);
xor U21551 (N_21551,N_19806,N_19116);
nand U21552 (N_21552,N_19805,N_19101);
and U21553 (N_21553,N_18913,N_19838);
or U21554 (N_21554,N_19481,N_19539);
nand U21555 (N_21555,N_18855,N_18065);
nor U21556 (N_21556,N_19366,N_17811);
and U21557 (N_21557,N_17915,N_19626);
nand U21558 (N_21558,N_19964,N_18480);
nand U21559 (N_21559,N_17625,N_19217);
nor U21560 (N_21560,N_19604,N_18886);
and U21561 (N_21561,N_19222,N_18585);
or U21562 (N_21562,N_19927,N_18626);
or U21563 (N_21563,N_19198,N_18794);
nand U21564 (N_21564,N_19305,N_17700);
nor U21565 (N_21565,N_19107,N_18863);
nand U21566 (N_21566,N_18849,N_17526);
nand U21567 (N_21567,N_17866,N_18046);
and U21568 (N_21568,N_18702,N_19642);
nor U21569 (N_21569,N_18013,N_18054);
and U21570 (N_21570,N_18462,N_19528);
xnor U21571 (N_21571,N_17581,N_17682);
or U21572 (N_21572,N_19046,N_18814);
nand U21573 (N_21573,N_19607,N_18506);
xor U21574 (N_21574,N_18392,N_19264);
xor U21575 (N_21575,N_18843,N_19084);
or U21576 (N_21576,N_19480,N_18845);
nand U21577 (N_21577,N_17921,N_19767);
or U21578 (N_21578,N_18098,N_19487);
nand U21579 (N_21579,N_19087,N_19212);
nor U21580 (N_21580,N_18326,N_17986);
nor U21581 (N_21581,N_17984,N_19996);
nor U21582 (N_21582,N_17978,N_17987);
and U21583 (N_21583,N_19583,N_19298);
nor U21584 (N_21584,N_19408,N_19074);
nor U21585 (N_21585,N_19391,N_18232);
nand U21586 (N_21586,N_19694,N_19317);
nor U21587 (N_21587,N_17686,N_19126);
nor U21588 (N_21588,N_17922,N_17643);
nand U21589 (N_21589,N_18099,N_19777);
nand U21590 (N_21590,N_19818,N_19379);
nor U21591 (N_21591,N_19846,N_19903);
and U21592 (N_21592,N_19358,N_18429);
nand U21593 (N_21593,N_18910,N_19936);
xor U21594 (N_21594,N_19210,N_18826);
xnor U21595 (N_21595,N_19044,N_18895);
and U21596 (N_21596,N_19444,N_18102);
nand U21597 (N_21597,N_18162,N_17814);
nor U21598 (N_21598,N_18366,N_19708);
nor U21599 (N_21599,N_19801,N_18548);
and U21600 (N_21600,N_18977,N_19814);
and U21601 (N_21601,N_18149,N_19909);
and U21602 (N_21602,N_17775,N_18985);
nand U21603 (N_21603,N_18199,N_19388);
nor U21604 (N_21604,N_17674,N_17986);
and U21605 (N_21605,N_17933,N_19517);
nor U21606 (N_21606,N_17887,N_19224);
nor U21607 (N_21607,N_19810,N_17959);
and U21608 (N_21608,N_19467,N_19820);
nand U21609 (N_21609,N_19266,N_17795);
nand U21610 (N_21610,N_19804,N_18096);
or U21611 (N_21611,N_17627,N_17784);
or U21612 (N_21612,N_18544,N_17689);
xor U21613 (N_21613,N_18221,N_19699);
nand U21614 (N_21614,N_18243,N_18458);
nand U21615 (N_21615,N_18088,N_19504);
and U21616 (N_21616,N_18602,N_19350);
nor U21617 (N_21617,N_18217,N_17515);
nand U21618 (N_21618,N_18321,N_18801);
or U21619 (N_21619,N_19914,N_19260);
nand U21620 (N_21620,N_19648,N_19116);
xnor U21621 (N_21621,N_18253,N_18882);
and U21622 (N_21622,N_19521,N_19790);
nand U21623 (N_21623,N_18643,N_18351);
nand U21624 (N_21624,N_18961,N_19672);
nand U21625 (N_21625,N_19127,N_18057);
or U21626 (N_21626,N_19618,N_18925);
nand U21627 (N_21627,N_19551,N_18021);
nand U21628 (N_21628,N_19389,N_17977);
or U21629 (N_21629,N_19130,N_19635);
or U21630 (N_21630,N_19793,N_17971);
and U21631 (N_21631,N_19380,N_19076);
nand U21632 (N_21632,N_19211,N_18350);
xor U21633 (N_21633,N_19716,N_19948);
nor U21634 (N_21634,N_18142,N_19358);
or U21635 (N_21635,N_18338,N_18118);
and U21636 (N_21636,N_17709,N_18035);
and U21637 (N_21637,N_18907,N_17956);
nor U21638 (N_21638,N_19211,N_17937);
xnor U21639 (N_21639,N_18108,N_19303);
nand U21640 (N_21640,N_17971,N_19227);
xnor U21641 (N_21641,N_19636,N_18515);
xnor U21642 (N_21642,N_17538,N_19473);
nor U21643 (N_21643,N_18192,N_19630);
nand U21644 (N_21644,N_18126,N_17979);
and U21645 (N_21645,N_18746,N_19411);
and U21646 (N_21646,N_18841,N_18380);
and U21647 (N_21647,N_17879,N_19859);
xnor U21648 (N_21648,N_18956,N_19256);
xor U21649 (N_21649,N_19539,N_19613);
nand U21650 (N_21650,N_19555,N_18426);
or U21651 (N_21651,N_19429,N_18268);
or U21652 (N_21652,N_17709,N_18430);
or U21653 (N_21653,N_19138,N_18142);
nor U21654 (N_21654,N_18089,N_18903);
xor U21655 (N_21655,N_19095,N_17510);
xnor U21656 (N_21656,N_17680,N_18504);
and U21657 (N_21657,N_18430,N_19509);
and U21658 (N_21658,N_17501,N_19450);
xor U21659 (N_21659,N_19435,N_19323);
xor U21660 (N_21660,N_17965,N_19661);
nor U21661 (N_21661,N_18120,N_17530);
nor U21662 (N_21662,N_19865,N_19312);
nor U21663 (N_21663,N_18346,N_18218);
xor U21664 (N_21664,N_18231,N_17559);
or U21665 (N_21665,N_18798,N_17663);
and U21666 (N_21666,N_19525,N_19942);
or U21667 (N_21667,N_17655,N_19611);
xor U21668 (N_21668,N_19657,N_19219);
nor U21669 (N_21669,N_18021,N_19774);
nand U21670 (N_21670,N_18802,N_17568);
xor U21671 (N_21671,N_17611,N_17865);
xnor U21672 (N_21672,N_17948,N_19123);
and U21673 (N_21673,N_18738,N_17915);
xor U21674 (N_21674,N_19199,N_18439);
and U21675 (N_21675,N_17972,N_19013);
or U21676 (N_21676,N_17717,N_19169);
xor U21677 (N_21677,N_19739,N_18397);
or U21678 (N_21678,N_19285,N_19983);
and U21679 (N_21679,N_19389,N_19290);
xor U21680 (N_21680,N_17803,N_18197);
xor U21681 (N_21681,N_19943,N_19956);
or U21682 (N_21682,N_18917,N_19031);
or U21683 (N_21683,N_18115,N_17803);
and U21684 (N_21684,N_19194,N_17974);
nor U21685 (N_21685,N_19316,N_19804);
nor U21686 (N_21686,N_17609,N_19956);
and U21687 (N_21687,N_19919,N_18671);
and U21688 (N_21688,N_18679,N_19122);
and U21689 (N_21689,N_18137,N_18323);
xor U21690 (N_21690,N_19195,N_18297);
or U21691 (N_21691,N_18414,N_19367);
or U21692 (N_21692,N_18083,N_19092);
nor U21693 (N_21693,N_18005,N_17523);
or U21694 (N_21694,N_19462,N_19518);
xnor U21695 (N_21695,N_19226,N_18821);
xor U21696 (N_21696,N_18060,N_17864);
nor U21697 (N_21697,N_18800,N_19721);
or U21698 (N_21698,N_18628,N_18032);
nor U21699 (N_21699,N_19516,N_18396);
or U21700 (N_21700,N_18171,N_17753);
and U21701 (N_21701,N_19988,N_18420);
nor U21702 (N_21702,N_19727,N_18476);
nor U21703 (N_21703,N_18185,N_18638);
nand U21704 (N_21704,N_19248,N_19049);
xor U21705 (N_21705,N_19400,N_18353);
nand U21706 (N_21706,N_19111,N_17757);
and U21707 (N_21707,N_17714,N_17891);
and U21708 (N_21708,N_19839,N_17803);
xnor U21709 (N_21709,N_19152,N_18937);
or U21710 (N_21710,N_17518,N_19217);
or U21711 (N_21711,N_18581,N_17756);
nand U21712 (N_21712,N_19847,N_17519);
or U21713 (N_21713,N_18654,N_18950);
xnor U21714 (N_21714,N_18952,N_19548);
and U21715 (N_21715,N_19347,N_19979);
and U21716 (N_21716,N_18658,N_19229);
and U21717 (N_21717,N_19203,N_18544);
nor U21718 (N_21718,N_19817,N_19183);
or U21719 (N_21719,N_18521,N_19238);
nor U21720 (N_21720,N_19930,N_18009);
or U21721 (N_21721,N_17542,N_18124);
xor U21722 (N_21722,N_18152,N_19686);
nor U21723 (N_21723,N_18770,N_19565);
nor U21724 (N_21724,N_17892,N_19326);
and U21725 (N_21725,N_18567,N_17597);
xor U21726 (N_21726,N_18223,N_18848);
xor U21727 (N_21727,N_17667,N_19963);
and U21728 (N_21728,N_19920,N_18292);
nor U21729 (N_21729,N_18073,N_18121);
xnor U21730 (N_21730,N_19819,N_19327);
nand U21731 (N_21731,N_18980,N_19006);
and U21732 (N_21732,N_18605,N_19432);
xnor U21733 (N_21733,N_18751,N_18400);
nand U21734 (N_21734,N_18176,N_19902);
nor U21735 (N_21735,N_17612,N_18374);
xor U21736 (N_21736,N_19263,N_19630);
and U21737 (N_21737,N_19625,N_17817);
and U21738 (N_21738,N_18781,N_17559);
nor U21739 (N_21739,N_19649,N_19001);
and U21740 (N_21740,N_18521,N_17753);
xnor U21741 (N_21741,N_17901,N_18953);
xnor U21742 (N_21742,N_18883,N_18892);
nor U21743 (N_21743,N_18069,N_18546);
nand U21744 (N_21744,N_18455,N_19386);
xor U21745 (N_21745,N_19021,N_19259);
xnor U21746 (N_21746,N_17808,N_18155);
xor U21747 (N_21747,N_19633,N_18118);
xnor U21748 (N_21748,N_17608,N_19628);
nor U21749 (N_21749,N_19461,N_19392);
nand U21750 (N_21750,N_19283,N_19209);
xor U21751 (N_21751,N_17704,N_18528);
or U21752 (N_21752,N_18722,N_17535);
and U21753 (N_21753,N_19588,N_19474);
and U21754 (N_21754,N_19644,N_19965);
and U21755 (N_21755,N_19696,N_19645);
and U21756 (N_21756,N_18813,N_19290);
nand U21757 (N_21757,N_19021,N_18498);
nor U21758 (N_21758,N_17533,N_18041);
nor U21759 (N_21759,N_19798,N_19776);
nand U21760 (N_21760,N_18236,N_18422);
nor U21761 (N_21761,N_18050,N_18022);
xor U21762 (N_21762,N_19310,N_19464);
or U21763 (N_21763,N_19771,N_17807);
or U21764 (N_21764,N_18401,N_18485);
and U21765 (N_21765,N_18937,N_18989);
or U21766 (N_21766,N_19073,N_18917);
nor U21767 (N_21767,N_18855,N_18761);
nand U21768 (N_21768,N_19836,N_17689);
nor U21769 (N_21769,N_19293,N_18814);
or U21770 (N_21770,N_18393,N_17634);
nor U21771 (N_21771,N_19278,N_17711);
nor U21772 (N_21772,N_18927,N_17890);
and U21773 (N_21773,N_18878,N_17563);
xor U21774 (N_21774,N_18606,N_19632);
and U21775 (N_21775,N_18918,N_17862);
nand U21776 (N_21776,N_19641,N_17867);
nand U21777 (N_21777,N_19734,N_19219);
or U21778 (N_21778,N_19662,N_18036);
nor U21779 (N_21779,N_18043,N_19569);
nor U21780 (N_21780,N_19829,N_19719);
nor U21781 (N_21781,N_18473,N_19347);
and U21782 (N_21782,N_18234,N_19343);
nand U21783 (N_21783,N_18857,N_19422);
or U21784 (N_21784,N_19173,N_18370);
nand U21785 (N_21785,N_19483,N_17692);
nor U21786 (N_21786,N_17672,N_19652);
xor U21787 (N_21787,N_19550,N_19917);
nand U21788 (N_21788,N_18268,N_18839);
nor U21789 (N_21789,N_19751,N_19103);
nand U21790 (N_21790,N_17852,N_18457);
nand U21791 (N_21791,N_18377,N_18537);
nand U21792 (N_21792,N_19160,N_19480);
nand U21793 (N_21793,N_18137,N_18174);
nor U21794 (N_21794,N_19199,N_18772);
and U21795 (N_21795,N_19991,N_19709);
or U21796 (N_21796,N_18445,N_17678);
nand U21797 (N_21797,N_19217,N_18491);
or U21798 (N_21798,N_19034,N_18812);
nor U21799 (N_21799,N_17731,N_19464);
nor U21800 (N_21800,N_18997,N_18922);
nor U21801 (N_21801,N_18136,N_18182);
xnor U21802 (N_21802,N_18490,N_19142);
or U21803 (N_21803,N_19574,N_18419);
xnor U21804 (N_21804,N_18996,N_18887);
nand U21805 (N_21805,N_18417,N_18952);
xnor U21806 (N_21806,N_18179,N_17556);
xnor U21807 (N_21807,N_18229,N_19001);
xor U21808 (N_21808,N_17790,N_18511);
or U21809 (N_21809,N_19695,N_17686);
and U21810 (N_21810,N_19598,N_18433);
or U21811 (N_21811,N_18474,N_19620);
or U21812 (N_21812,N_18864,N_19479);
nor U21813 (N_21813,N_18305,N_19051);
or U21814 (N_21814,N_18983,N_19252);
or U21815 (N_21815,N_17693,N_19551);
and U21816 (N_21816,N_18472,N_18260);
xor U21817 (N_21817,N_18191,N_18261);
and U21818 (N_21818,N_19000,N_17519);
nor U21819 (N_21819,N_19943,N_19892);
or U21820 (N_21820,N_19393,N_17502);
and U21821 (N_21821,N_18761,N_19733);
and U21822 (N_21822,N_18502,N_18559);
and U21823 (N_21823,N_19867,N_17564);
nor U21824 (N_21824,N_18336,N_17874);
nor U21825 (N_21825,N_18332,N_18966);
nor U21826 (N_21826,N_19309,N_18450);
nor U21827 (N_21827,N_18808,N_19767);
or U21828 (N_21828,N_19320,N_19864);
and U21829 (N_21829,N_18196,N_19142);
xor U21830 (N_21830,N_19577,N_19693);
nand U21831 (N_21831,N_18389,N_18976);
xor U21832 (N_21832,N_18023,N_18079);
nand U21833 (N_21833,N_17876,N_18152);
and U21834 (N_21834,N_18718,N_19750);
nand U21835 (N_21835,N_17556,N_18557);
xor U21836 (N_21836,N_19639,N_17824);
and U21837 (N_21837,N_19304,N_17916);
or U21838 (N_21838,N_18779,N_19191);
or U21839 (N_21839,N_19173,N_19865);
or U21840 (N_21840,N_17690,N_19603);
or U21841 (N_21841,N_18764,N_18391);
nor U21842 (N_21842,N_17770,N_18337);
nand U21843 (N_21843,N_19105,N_19168);
and U21844 (N_21844,N_19176,N_19133);
nor U21845 (N_21845,N_17692,N_19551);
and U21846 (N_21846,N_18041,N_18225);
or U21847 (N_21847,N_17504,N_18938);
or U21848 (N_21848,N_18549,N_19818);
and U21849 (N_21849,N_17711,N_18018);
nor U21850 (N_21850,N_18326,N_18180);
nor U21851 (N_21851,N_19299,N_19000);
nand U21852 (N_21852,N_17838,N_19293);
and U21853 (N_21853,N_18534,N_18040);
xnor U21854 (N_21854,N_18040,N_17854);
xor U21855 (N_21855,N_17825,N_18384);
nand U21856 (N_21856,N_18568,N_18423);
nand U21857 (N_21857,N_17827,N_19198);
and U21858 (N_21858,N_19256,N_19130);
and U21859 (N_21859,N_18116,N_17587);
xnor U21860 (N_21860,N_18422,N_19049);
nor U21861 (N_21861,N_19742,N_18213);
and U21862 (N_21862,N_18616,N_17959);
and U21863 (N_21863,N_17727,N_18711);
xor U21864 (N_21864,N_19827,N_19072);
nor U21865 (N_21865,N_19895,N_19221);
nand U21866 (N_21866,N_18436,N_18650);
and U21867 (N_21867,N_19714,N_17967);
or U21868 (N_21868,N_17850,N_18259);
nor U21869 (N_21869,N_18823,N_18656);
nor U21870 (N_21870,N_19385,N_19995);
nand U21871 (N_21871,N_18928,N_19889);
nor U21872 (N_21872,N_19959,N_19644);
nor U21873 (N_21873,N_19952,N_18772);
nand U21874 (N_21874,N_19857,N_17912);
nor U21875 (N_21875,N_17561,N_18436);
nand U21876 (N_21876,N_17892,N_19628);
xor U21877 (N_21877,N_19358,N_18645);
xnor U21878 (N_21878,N_18484,N_19748);
nand U21879 (N_21879,N_18447,N_19141);
nor U21880 (N_21880,N_19237,N_19246);
or U21881 (N_21881,N_19879,N_19321);
xnor U21882 (N_21882,N_17587,N_19556);
nand U21883 (N_21883,N_17874,N_17637);
xor U21884 (N_21884,N_18883,N_18919);
or U21885 (N_21885,N_17685,N_18432);
nor U21886 (N_21886,N_17902,N_18213);
nand U21887 (N_21887,N_19551,N_17785);
xnor U21888 (N_21888,N_19328,N_18329);
nor U21889 (N_21889,N_17564,N_19190);
or U21890 (N_21890,N_19531,N_18791);
xor U21891 (N_21891,N_18077,N_19269);
or U21892 (N_21892,N_17612,N_19099);
nor U21893 (N_21893,N_18718,N_18062);
nor U21894 (N_21894,N_17961,N_17509);
or U21895 (N_21895,N_19061,N_19281);
or U21896 (N_21896,N_19725,N_18441);
nor U21897 (N_21897,N_19157,N_18111);
nand U21898 (N_21898,N_18273,N_19931);
or U21899 (N_21899,N_18525,N_18335);
xnor U21900 (N_21900,N_19152,N_17732);
or U21901 (N_21901,N_19755,N_17672);
and U21902 (N_21902,N_17597,N_18668);
xor U21903 (N_21903,N_19448,N_19305);
nor U21904 (N_21904,N_17941,N_19545);
xnor U21905 (N_21905,N_19925,N_17821);
xor U21906 (N_21906,N_17657,N_18567);
nor U21907 (N_21907,N_18188,N_18955);
xnor U21908 (N_21908,N_19640,N_19008);
or U21909 (N_21909,N_18019,N_18798);
nand U21910 (N_21910,N_19492,N_18414);
nand U21911 (N_21911,N_17905,N_19159);
and U21912 (N_21912,N_18468,N_19623);
nor U21913 (N_21913,N_17963,N_17997);
or U21914 (N_21914,N_17827,N_18260);
xnor U21915 (N_21915,N_19348,N_18817);
nand U21916 (N_21916,N_19982,N_19347);
or U21917 (N_21917,N_18714,N_18575);
or U21918 (N_21918,N_18778,N_18303);
or U21919 (N_21919,N_19463,N_17845);
or U21920 (N_21920,N_19915,N_18137);
xor U21921 (N_21921,N_19216,N_17818);
and U21922 (N_21922,N_18114,N_18547);
and U21923 (N_21923,N_17622,N_17691);
nor U21924 (N_21924,N_19359,N_17724);
nor U21925 (N_21925,N_19661,N_19819);
nand U21926 (N_21926,N_19106,N_19522);
nor U21927 (N_21927,N_19587,N_18745);
xor U21928 (N_21928,N_18124,N_18383);
or U21929 (N_21929,N_17853,N_18067);
xor U21930 (N_21930,N_18265,N_19069);
nor U21931 (N_21931,N_17909,N_18225);
or U21932 (N_21932,N_18356,N_17874);
xor U21933 (N_21933,N_18915,N_19526);
or U21934 (N_21934,N_17827,N_18299);
nor U21935 (N_21935,N_18453,N_18619);
or U21936 (N_21936,N_19625,N_17644);
xor U21937 (N_21937,N_18235,N_19927);
xnor U21938 (N_21938,N_18317,N_17745);
nand U21939 (N_21939,N_18842,N_18038);
nor U21940 (N_21940,N_17643,N_17801);
nand U21941 (N_21941,N_17508,N_17712);
and U21942 (N_21942,N_19171,N_18202);
nor U21943 (N_21943,N_18048,N_18151);
nor U21944 (N_21944,N_18393,N_18192);
or U21945 (N_21945,N_18481,N_18139);
nor U21946 (N_21946,N_19407,N_17584);
nor U21947 (N_21947,N_19061,N_18499);
xor U21948 (N_21948,N_18965,N_18246);
nor U21949 (N_21949,N_19671,N_18961);
or U21950 (N_21950,N_18063,N_19293);
and U21951 (N_21951,N_17507,N_19045);
or U21952 (N_21952,N_17716,N_17575);
nor U21953 (N_21953,N_18319,N_18798);
and U21954 (N_21954,N_17684,N_17999);
xnor U21955 (N_21955,N_19222,N_18784);
xnor U21956 (N_21956,N_18044,N_18643);
or U21957 (N_21957,N_17903,N_18648);
nand U21958 (N_21958,N_17959,N_19545);
or U21959 (N_21959,N_18387,N_18314);
nor U21960 (N_21960,N_17801,N_18596);
or U21961 (N_21961,N_18701,N_18594);
nor U21962 (N_21962,N_18922,N_19099);
or U21963 (N_21963,N_19502,N_17545);
nor U21964 (N_21964,N_19295,N_18748);
and U21965 (N_21965,N_19683,N_18625);
and U21966 (N_21966,N_19965,N_19894);
or U21967 (N_21967,N_19492,N_18773);
and U21968 (N_21968,N_18939,N_17771);
xor U21969 (N_21969,N_19423,N_19590);
xnor U21970 (N_21970,N_19851,N_19675);
and U21971 (N_21971,N_18573,N_19052);
xor U21972 (N_21972,N_18054,N_18296);
xnor U21973 (N_21973,N_19644,N_18564);
nand U21974 (N_21974,N_17507,N_18694);
xnor U21975 (N_21975,N_19029,N_18993);
xnor U21976 (N_21976,N_19744,N_19375);
xor U21977 (N_21977,N_17953,N_18826);
or U21978 (N_21978,N_17633,N_19886);
or U21979 (N_21979,N_18900,N_19433);
or U21980 (N_21980,N_18400,N_18654);
or U21981 (N_21981,N_18055,N_17583);
nor U21982 (N_21982,N_19140,N_19711);
or U21983 (N_21983,N_18785,N_18384);
nor U21984 (N_21984,N_19699,N_18499);
nand U21985 (N_21985,N_18161,N_18975);
nand U21986 (N_21986,N_19017,N_19515);
or U21987 (N_21987,N_19754,N_19953);
nand U21988 (N_21988,N_17857,N_17820);
and U21989 (N_21989,N_19943,N_19514);
and U21990 (N_21990,N_19409,N_19963);
or U21991 (N_21991,N_18769,N_18260);
or U21992 (N_21992,N_17780,N_17569);
and U21993 (N_21993,N_18212,N_19040);
nor U21994 (N_21994,N_19503,N_19763);
or U21995 (N_21995,N_18840,N_18298);
nand U21996 (N_21996,N_18916,N_19927);
nor U21997 (N_21997,N_18855,N_18099);
and U21998 (N_21998,N_19050,N_19319);
nor U21999 (N_21999,N_18418,N_19057);
nor U22000 (N_22000,N_19388,N_18041);
nand U22001 (N_22001,N_17786,N_19005);
or U22002 (N_22002,N_19735,N_19522);
or U22003 (N_22003,N_19814,N_17945);
or U22004 (N_22004,N_19455,N_18930);
and U22005 (N_22005,N_19537,N_18478);
and U22006 (N_22006,N_18869,N_17662);
xor U22007 (N_22007,N_18602,N_18439);
and U22008 (N_22008,N_18062,N_18082);
nor U22009 (N_22009,N_18775,N_18945);
and U22010 (N_22010,N_18020,N_19355);
nor U22011 (N_22011,N_19183,N_17598);
nand U22012 (N_22012,N_19791,N_18083);
and U22013 (N_22013,N_18065,N_18841);
xor U22014 (N_22014,N_17745,N_18820);
nor U22015 (N_22015,N_18183,N_19323);
or U22016 (N_22016,N_17599,N_18109);
nand U22017 (N_22017,N_18794,N_17517);
or U22018 (N_22018,N_19889,N_19800);
nand U22019 (N_22019,N_17917,N_18670);
or U22020 (N_22020,N_17677,N_18075);
or U22021 (N_22021,N_18043,N_19752);
nor U22022 (N_22022,N_19225,N_17648);
xnor U22023 (N_22023,N_19031,N_18227);
xor U22024 (N_22024,N_17836,N_19853);
nand U22025 (N_22025,N_17578,N_17846);
or U22026 (N_22026,N_18511,N_19880);
and U22027 (N_22027,N_19579,N_17809);
and U22028 (N_22028,N_19425,N_19387);
nor U22029 (N_22029,N_17612,N_18756);
xor U22030 (N_22030,N_18245,N_17840);
xor U22031 (N_22031,N_17683,N_18531);
and U22032 (N_22032,N_19748,N_18435);
nand U22033 (N_22033,N_19591,N_17858);
xor U22034 (N_22034,N_17582,N_19140);
nor U22035 (N_22035,N_19131,N_19238);
or U22036 (N_22036,N_19204,N_18329);
nor U22037 (N_22037,N_18805,N_18192);
xnor U22038 (N_22038,N_19237,N_19085);
xor U22039 (N_22039,N_19190,N_19534);
nor U22040 (N_22040,N_19642,N_19447);
nor U22041 (N_22041,N_17648,N_18956);
nand U22042 (N_22042,N_17704,N_17738);
nand U22043 (N_22043,N_18370,N_19122);
xnor U22044 (N_22044,N_18679,N_17646);
and U22045 (N_22045,N_17952,N_17813);
and U22046 (N_22046,N_18518,N_19624);
xnor U22047 (N_22047,N_19643,N_19453);
nand U22048 (N_22048,N_17618,N_18017);
and U22049 (N_22049,N_19739,N_17724);
xor U22050 (N_22050,N_18174,N_18492);
nor U22051 (N_22051,N_19165,N_18059);
xnor U22052 (N_22052,N_18688,N_19571);
and U22053 (N_22053,N_18615,N_19524);
xor U22054 (N_22054,N_19994,N_17959);
nand U22055 (N_22055,N_19818,N_18764);
nor U22056 (N_22056,N_18517,N_18385);
nor U22057 (N_22057,N_18729,N_18238);
xnor U22058 (N_22058,N_19782,N_18619);
nor U22059 (N_22059,N_19625,N_18149);
nor U22060 (N_22060,N_19371,N_18527);
nor U22061 (N_22061,N_18893,N_18736);
or U22062 (N_22062,N_18181,N_19082);
and U22063 (N_22063,N_19674,N_17533);
xor U22064 (N_22064,N_19777,N_18016);
nand U22065 (N_22065,N_18894,N_18531);
or U22066 (N_22066,N_19443,N_18670);
and U22067 (N_22067,N_19833,N_17963);
or U22068 (N_22068,N_17978,N_19814);
nor U22069 (N_22069,N_19503,N_19958);
or U22070 (N_22070,N_18495,N_19333);
or U22071 (N_22071,N_19788,N_17779);
nand U22072 (N_22072,N_17561,N_19594);
nor U22073 (N_22073,N_19406,N_19977);
and U22074 (N_22074,N_18042,N_19633);
and U22075 (N_22075,N_17598,N_18800);
nor U22076 (N_22076,N_19979,N_19450);
and U22077 (N_22077,N_17748,N_18527);
nor U22078 (N_22078,N_19871,N_18464);
or U22079 (N_22079,N_17608,N_19808);
nand U22080 (N_22080,N_18412,N_17744);
or U22081 (N_22081,N_18641,N_19498);
and U22082 (N_22082,N_18817,N_19750);
nand U22083 (N_22083,N_19762,N_19467);
nor U22084 (N_22084,N_18094,N_18323);
nand U22085 (N_22085,N_19874,N_18307);
and U22086 (N_22086,N_19852,N_17647);
nor U22087 (N_22087,N_18674,N_19420);
and U22088 (N_22088,N_18014,N_18002);
and U22089 (N_22089,N_19804,N_19740);
nand U22090 (N_22090,N_19067,N_19914);
or U22091 (N_22091,N_18831,N_18655);
nand U22092 (N_22092,N_19434,N_17782);
nor U22093 (N_22093,N_19160,N_18967);
and U22094 (N_22094,N_19899,N_18070);
nand U22095 (N_22095,N_19730,N_18435);
nand U22096 (N_22096,N_18361,N_18339);
xnor U22097 (N_22097,N_19649,N_18082);
nor U22098 (N_22098,N_19690,N_18561);
xor U22099 (N_22099,N_18937,N_17737);
nand U22100 (N_22100,N_18228,N_17673);
nand U22101 (N_22101,N_19825,N_17909);
and U22102 (N_22102,N_18413,N_18701);
nand U22103 (N_22103,N_18858,N_18988);
or U22104 (N_22104,N_18025,N_19319);
and U22105 (N_22105,N_19359,N_18645);
or U22106 (N_22106,N_18594,N_19812);
nand U22107 (N_22107,N_18949,N_18483);
nor U22108 (N_22108,N_19277,N_19431);
and U22109 (N_22109,N_17989,N_17616);
xor U22110 (N_22110,N_18933,N_18449);
nand U22111 (N_22111,N_18569,N_19576);
xnor U22112 (N_22112,N_19783,N_18587);
and U22113 (N_22113,N_19963,N_19580);
or U22114 (N_22114,N_19802,N_18814);
and U22115 (N_22115,N_19929,N_17920);
xor U22116 (N_22116,N_17562,N_19677);
or U22117 (N_22117,N_19414,N_19658);
nand U22118 (N_22118,N_17687,N_18794);
xor U22119 (N_22119,N_18546,N_19583);
or U22120 (N_22120,N_17566,N_19142);
xor U22121 (N_22121,N_18600,N_19885);
or U22122 (N_22122,N_19004,N_19340);
xor U22123 (N_22123,N_19638,N_18626);
nand U22124 (N_22124,N_18005,N_17679);
and U22125 (N_22125,N_18464,N_18837);
nand U22126 (N_22126,N_18962,N_18810);
or U22127 (N_22127,N_18173,N_18658);
nor U22128 (N_22128,N_18806,N_18526);
nor U22129 (N_22129,N_18516,N_17580);
xnor U22130 (N_22130,N_17791,N_17758);
nor U22131 (N_22131,N_17943,N_18625);
or U22132 (N_22132,N_19240,N_19180);
and U22133 (N_22133,N_17512,N_18191);
and U22134 (N_22134,N_17719,N_18626);
and U22135 (N_22135,N_18667,N_19411);
nand U22136 (N_22136,N_19508,N_17796);
nand U22137 (N_22137,N_18967,N_17622);
xnor U22138 (N_22138,N_18972,N_18442);
and U22139 (N_22139,N_17558,N_17547);
xnor U22140 (N_22140,N_19432,N_19806);
xor U22141 (N_22141,N_18517,N_17524);
and U22142 (N_22142,N_18044,N_18564);
nor U22143 (N_22143,N_17865,N_19644);
or U22144 (N_22144,N_19918,N_19023);
xor U22145 (N_22145,N_17591,N_17604);
nor U22146 (N_22146,N_19645,N_19512);
xor U22147 (N_22147,N_18617,N_18540);
nand U22148 (N_22148,N_18482,N_18911);
nor U22149 (N_22149,N_19556,N_17698);
or U22150 (N_22150,N_19269,N_18303);
and U22151 (N_22151,N_18130,N_19981);
and U22152 (N_22152,N_19371,N_18705);
and U22153 (N_22153,N_19560,N_18847);
nor U22154 (N_22154,N_17519,N_18937);
nand U22155 (N_22155,N_18391,N_18626);
and U22156 (N_22156,N_19828,N_18624);
and U22157 (N_22157,N_18998,N_17612);
nor U22158 (N_22158,N_18584,N_17731);
and U22159 (N_22159,N_17529,N_18031);
nor U22160 (N_22160,N_19875,N_18145);
nand U22161 (N_22161,N_17992,N_18128);
nor U22162 (N_22162,N_19629,N_19741);
xnor U22163 (N_22163,N_19502,N_18548);
xor U22164 (N_22164,N_18769,N_19384);
and U22165 (N_22165,N_17642,N_19798);
or U22166 (N_22166,N_17680,N_18011);
or U22167 (N_22167,N_19869,N_18286);
nor U22168 (N_22168,N_19701,N_18543);
nand U22169 (N_22169,N_18339,N_19416);
or U22170 (N_22170,N_19999,N_17832);
or U22171 (N_22171,N_19207,N_18179);
nor U22172 (N_22172,N_19436,N_19779);
or U22173 (N_22173,N_17863,N_19202);
xor U22174 (N_22174,N_17578,N_19760);
xor U22175 (N_22175,N_17964,N_19851);
xnor U22176 (N_22176,N_19987,N_18997);
nand U22177 (N_22177,N_18472,N_18632);
nor U22178 (N_22178,N_19934,N_19958);
nor U22179 (N_22179,N_17535,N_19016);
nor U22180 (N_22180,N_18423,N_19780);
and U22181 (N_22181,N_19775,N_19714);
nor U22182 (N_22182,N_19857,N_19804);
xnor U22183 (N_22183,N_18927,N_19526);
xor U22184 (N_22184,N_17777,N_19438);
or U22185 (N_22185,N_19618,N_18994);
and U22186 (N_22186,N_18370,N_18576);
nor U22187 (N_22187,N_18239,N_19853);
or U22188 (N_22188,N_18386,N_19826);
nor U22189 (N_22189,N_19718,N_19575);
nor U22190 (N_22190,N_19793,N_18175);
xnor U22191 (N_22191,N_18422,N_18872);
xor U22192 (N_22192,N_18260,N_19541);
and U22193 (N_22193,N_17700,N_18011);
or U22194 (N_22194,N_18948,N_18937);
and U22195 (N_22195,N_17929,N_18544);
or U22196 (N_22196,N_18898,N_18232);
nor U22197 (N_22197,N_19289,N_18990);
xor U22198 (N_22198,N_19834,N_19015);
nand U22199 (N_22199,N_17612,N_17511);
and U22200 (N_22200,N_18146,N_18813);
or U22201 (N_22201,N_18535,N_19259);
and U22202 (N_22202,N_19213,N_18243);
and U22203 (N_22203,N_18631,N_19184);
nor U22204 (N_22204,N_19417,N_17680);
xor U22205 (N_22205,N_19599,N_19953);
nand U22206 (N_22206,N_19531,N_19541);
nor U22207 (N_22207,N_17790,N_17850);
and U22208 (N_22208,N_17807,N_17920);
xor U22209 (N_22209,N_17538,N_19759);
nor U22210 (N_22210,N_18079,N_18792);
and U22211 (N_22211,N_17698,N_18323);
xor U22212 (N_22212,N_18329,N_19131);
and U22213 (N_22213,N_18904,N_17753);
nand U22214 (N_22214,N_17868,N_18857);
and U22215 (N_22215,N_17960,N_19582);
xor U22216 (N_22216,N_18475,N_19732);
and U22217 (N_22217,N_18264,N_18533);
xor U22218 (N_22218,N_18306,N_17999);
or U22219 (N_22219,N_18052,N_19019);
or U22220 (N_22220,N_18902,N_18978);
and U22221 (N_22221,N_19271,N_17965);
and U22222 (N_22222,N_18048,N_19503);
or U22223 (N_22223,N_19828,N_19185);
or U22224 (N_22224,N_19086,N_17733);
nand U22225 (N_22225,N_19590,N_18309);
or U22226 (N_22226,N_17653,N_18971);
nor U22227 (N_22227,N_19622,N_18305);
or U22228 (N_22228,N_18243,N_18936);
and U22229 (N_22229,N_19446,N_17842);
or U22230 (N_22230,N_18881,N_17641);
xor U22231 (N_22231,N_19589,N_18293);
xor U22232 (N_22232,N_19712,N_18847);
xor U22233 (N_22233,N_19771,N_18425);
xor U22234 (N_22234,N_18909,N_18418);
nand U22235 (N_22235,N_19694,N_18539);
or U22236 (N_22236,N_17994,N_19369);
nand U22237 (N_22237,N_18631,N_18932);
nand U22238 (N_22238,N_19845,N_17635);
xor U22239 (N_22239,N_19824,N_18612);
or U22240 (N_22240,N_19858,N_17871);
nand U22241 (N_22241,N_17756,N_18177);
and U22242 (N_22242,N_18790,N_19464);
xnor U22243 (N_22243,N_18854,N_19335);
xnor U22244 (N_22244,N_17879,N_19723);
nor U22245 (N_22245,N_19138,N_17715);
nor U22246 (N_22246,N_18162,N_19421);
nor U22247 (N_22247,N_19227,N_19787);
or U22248 (N_22248,N_18072,N_19083);
nor U22249 (N_22249,N_19043,N_19590);
nand U22250 (N_22250,N_18348,N_18674);
nor U22251 (N_22251,N_18941,N_19642);
xor U22252 (N_22252,N_19862,N_19091);
and U22253 (N_22253,N_18730,N_18536);
or U22254 (N_22254,N_19432,N_19555);
xnor U22255 (N_22255,N_18101,N_19503);
xnor U22256 (N_22256,N_17643,N_19144);
xnor U22257 (N_22257,N_19819,N_19711);
or U22258 (N_22258,N_19488,N_19107);
nand U22259 (N_22259,N_19186,N_18718);
and U22260 (N_22260,N_18512,N_19545);
nor U22261 (N_22261,N_19718,N_19797);
nor U22262 (N_22262,N_19664,N_17525);
xor U22263 (N_22263,N_19472,N_17917);
and U22264 (N_22264,N_18069,N_18841);
nand U22265 (N_22265,N_18833,N_19009);
and U22266 (N_22266,N_19631,N_18973);
nand U22267 (N_22267,N_17672,N_18491);
and U22268 (N_22268,N_17877,N_18518);
nand U22269 (N_22269,N_18284,N_19838);
nor U22270 (N_22270,N_19717,N_17590);
nor U22271 (N_22271,N_19939,N_19663);
xor U22272 (N_22272,N_19206,N_18544);
xnor U22273 (N_22273,N_19510,N_17855);
and U22274 (N_22274,N_19315,N_19038);
nor U22275 (N_22275,N_18811,N_19645);
or U22276 (N_22276,N_17932,N_17651);
or U22277 (N_22277,N_19434,N_18466);
nor U22278 (N_22278,N_17667,N_19095);
or U22279 (N_22279,N_18937,N_19573);
and U22280 (N_22280,N_17987,N_19368);
nor U22281 (N_22281,N_18227,N_18956);
or U22282 (N_22282,N_18616,N_17651);
and U22283 (N_22283,N_19124,N_17518);
nand U22284 (N_22284,N_18504,N_18985);
nand U22285 (N_22285,N_18346,N_19937);
and U22286 (N_22286,N_18252,N_17988);
nor U22287 (N_22287,N_19869,N_19999);
and U22288 (N_22288,N_18145,N_19287);
nand U22289 (N_22289,N_18367,N_19348);
xor U22290 (N_22290,N_18274,N_17944);
nor U22291 (N_22291,N_18916,N_19514);
and U22292 (N_22292,N_17634,N_19006);
nand U22293 (N_22293,N_18173,N_18977);
and U22294 (N_22294,N_17633,N_19526);
nor U22295 (N_22295,N_18556,N_18940);
or U22296 (N_22296,N_17596,N_18141);
or U22297 (N_22297,N_19611,N_19225);
and U22298 (N_22298,N_18484,N_19173);
xor U22299 (N_22299,N_19943,N_19750);
nand U22300 (N_22300,N_18274,N_18205);
and U22301 (N_22301,N_17911,N_19606);
xnor U22302 (N_22302,N_18987,N_17638);
nor U22303 (N_22303,N_17741,N_19555);
nor U22304 (N_22304,N_19030,N_17879);
nand U22305 (N_22305,N_18940,N_19969);
nand U22306 (N_22306,N_18972,N_19636);
nor U22307 (N_22307,N_19035,N_19746);
xor U22308 (N_22308,N_18662,N_17801);
or U22309 (N_22309,N_17848,N_18878);
nand U22310 (N_22310,N_17912,N_17559);
and U22311 (N_22311,N_19071,N_17512);
and U22312 (N_22312,N_18315,N_18823);
nand U22313 (N_22313,N_19540,N_17624);
or U22314 (N_22314,N_17880,N_19901);
and U22315 (N_22315,N_19509,N_19468);
or U22316 (N_22316,N_19016,N_19019);
and U22317 (N_22317,N_19211,N_17961);
nor U22318 (N_22318,N_17911,N_19738);
and U22319 (N_22319,N_18788,N_17889);
xnor U22320 (N_22320,N_19962,N_17682);
nand U22321 (N_22321,N_18468,N_17611);
xnor U22322 (N_22322,N_19653,N_17824);
or U22323 (N_22323,N_19555,N_18439);
or U22324 (N_22324,N_17874,N_18682);
xnor U22325 (N_22325,N_18542,N_18300);
or U22326 (N_22326,N_18854,N_17683);
nor U22327 (N_22327,N_18038,N_17597);
or U22328 (N_22328,N_19496,N_19675);
xor U22329 (N_22329,N_18077,N_18903);
nor U22330 (N_22330,N_19895,N_19268);
and U22331 (N_22331,N_17703,N_18082);
nand U22332 (N_22332,N_19660,N_18370);
nor U22333 (N_22333,N_17738,N_19369);
and U22334 (N_22334,N_17667,N_18361);
or U22335 (N_22335,N_19186,N_18920);
nand U22336 (N_22336,N_19029,N_19263);
xor U22337 (N_22337,N_19387,N_18388);
and U22338 (N_22338,N_18198,N_19657);
and U22339 (N_22339,N_18330,N_19083);
xnor U22340 (N_22340,N_19883,N_18468);
nand U22341 (N_22341,N_19208,N_17882);
xnor U22342 (N_22342,N_17530,N_18017);
and U22343 (N_22343,N_17564,N_19964);
nand U22344 (N_22344,N_17819,N_17744);
nand U22345 (N_22345,N_18135,N_19016);
and U22346 (N_22346,N_17969,N_19033);
nand U22347 (N_22347,N_19717,N_18878);
or U22348 (N_22348,N_18417,N_19527);
nand U22349 (N_22349,N_18181,N_19930);
nand U22350 (N_22350,N_19878,N_18042);
or U22351 (N_22351,N_19547,N_19739);
xnor U22352 (N_22352,N_18516,N_19433);
nor U22353 (N_22353,N_19536,N_18898);
or U22354 (N_22354,N_19454,N_19664);
or U22355 (N_22355,N_19834,N_19199);
and U22356 (N_22356,N_19155,N_18438);
nand U22357 (N_22357,N_18058,N_19305);
and U22358 (N_22358,N_19752,N_19890);
nor U22359 (N_22359,N_19674,N_17813);
nor U22360 (N_22360,N_19287,N_18216);
nor U22361 (N_22361,N_19203,N_19652);
xnor U22362 (N_22362,N_17660,N_17809);
nor U22363 (N_22363,N_17947,N_19467);
and U22364 (N_22364,N_18005,N_18796);
or U22365 (N_22365,N_19075,N_19864);
or U22366 (N_22366,N_17680,N_19781);
or U22367 (N_22367,N_18215,N_18233);
xor U22368 (N_22368,N_17795,N_19251);
nor U22369 (N_22369,N_19874,N_19947);
xor U22370 (N_22370,N_18714,N_18015);
nand U22371 (N_22371,N_18849,N_17929);
xnor U22372 (N_22372,N_18659,N_19576);
xnor U22373 (N_22373,N_18235,N_18762);
or U22374 (N_22374,N_17966,N_18891);
and U22375 (N_22375,N_19643,N_19965);
xor U22376 (N_22376,N_19021,N_18330);
and U22377 (N_22377,N_19479,N_18409);
nor U22378 (N_22378,N_17941,N_17544);
xor U22379 (N_22379,N_19308,N_18725);
nand U22380 (N_22380,N_19264,N_19238);
nor U22381 (N_22381,N_18990,N_19759);
nand U22382 (N_22382,N_19065,N_18241);
and U22383 (N_22383,N_18494,N_19747);
and U22384 (N_22384,N_19619,N_17529);
nor U22385 (N_22385,N_18726,N_17929);
nand U22386 (N_22386,N_18182,N_18756);
nor U22387 (N_22387,N_18154,N_17576);
nand U22388 (N_22388,N_19541,N_18851);
and U22389 (N_22389,N_17863,N_19815);
nor U22390 (N_22390,N_18100,N_19415);
nor U22391 (N_22391,N_18795,N_19886);
or U22392 (N_22392,N_19125,N_18521);
xor U22393 (N_22393,N_19352,N_19593);
nor U22394 (N_22394,N_18120,N_19537);
nor U22395 (N_22395,N_18877,N_18510);
and U22396 (N_22396,N_19893,N_19023);
and U22397 (N_22397,N_18621,N_18319);
xnor U22398 (N_22398,N_18469,N_18475);
nor U22399 (N_22399,N_17925,N_19236);
and U22400 (N_22400,N_19565,N_18087);
xor U22401 (N_22401,N_19601,N_19490);
xor U22402 (N_22402,N_18395,N_18599);
xor U22403 (N_22403,N_18195,N_18906);
xnor U22404 (N_22404,N_18316,N_19278);
and U22405 (N_22405,N_19472,N_19792);
xor U22406 (N_22406,N_19111,N_19997);
and U22407 (N_22407,N_19160,N_18437);
or U22408 (N_22408,N_18948,N_19202);
and U22409 (N_22409,N_18661,N_19469);
nor U22410 (N_22410,N_19224,N_18456);
and U22411 (N_22411,N_18707,N_18891);
and U22412 (N_22412,N_18606,N_18815);
xor U22413 (N_22413,N_19686,N_17852);
xor U22414 (N_22414,N_18298,N_18357);
nand U22415 (N_22415,N_19626,N_19737);
nor U22416 (N_22416,N_18357,N_18315);
and U22417 (N_22417,N_18727,N_19451);
or U22418 (N_22418,N_18512,N_19128);
nor U22419 (N_22419,N_19312,N_18742);
nand U22420 (N_22420,N_18285,N_19479);
xnor U22421 (N_22421,N_19464,N_17689);
nor U22422 (N_22422,N_18685,N_19519);
nor U22423 (N_22423,N_19756,N_17934);
xor U22424 (N_22424,N_18045,N_17974);
nor U22425 (N_22425,N_19846,N_18047);
xor U22426 (N_22426,N_19748,N_18321);
nand U22427 (N_22427,N_18051,N_19705);
or U22428 (N_22428,N_18181,N_19457);
and U22429 (N_22429,N_18931,N_18241);
and U22430 (N_22430,N_19488,N_18283);
or U22431 (N_22431,N_19484,N_19768);
or U22432 (N_22432,N_18429,N_17806);
xor U22433 (N_22433,N_18212,N_17989);
or U22434 (N_22434,N_17522,N_17961);
nand U22435 (N_22435,N_18307,N_17761);
nor U22436 (N_22436,N_18576,N_19932);
nor U22437 (N_22437,N_18892,N_18299);
and U22438 (N_22438,N_18591,N_17634);
xor U22439 (N_22439,N_19624,N_19525);
nor U22440 (N_22440,N_17893,N_19716);
or U22441 (N_22441,N_18610,N_19651);
nand U22442 (N_22442,N_19598,N_19830);
nor U22443 (N_22443,N_18396,N_19720);
nor U22444 (N_22444,N_19981,N_19493);
nor U22445 (N_22445,N_17802,N_17919);
nand U22446 (N_22446,N_17940,N_19799);
nand U22447 (N_22447,N_17652,N_18588);
or U22448 (N_22448,N_17791,N_19218);
or U22449 (N_22449,N_18995,N_17717);
and U22450 (N_22450,N_19101,N_19273);
and U22451 (N_22451,N_18649,N_19500);
or U22452 (N_22452,N_17599,N_18478);
and U22453 (N_22453,N_19523,N_17806);
xor U22454 (N_22454,N_18264,N_18153);
nand U22455 (N_22455,N_17967,N_17568);
and U22456 (N_22456,N_19897,N_18550);
or U22457 (N_22457,N_17659,N_19534);
or U22458 (N_22458,N_17968,N_18576);
nand U22459 (N_22459,N_18414,N_17584);
nor U22460 (N_22460,N_18138,N_19250);
nand U22461 (N_22461,N_19580,N_19233);
nand U22462 (N_22462,N_18880,N_17998);
or U22463 (N_22463,N_18107,N_19144);
and U22464 (N_22464,N_18626,N_19473);
xnor U22465 (N_22465,N_19020,N_18727);
or U22466 (N_22466,N_18465,N_17593);
or U22467 (N_22467,N_18546,N_18322);
xor U22468 (N_22468,N_19595,N_19925);
or U22469 (N_22469,N_18725,N_19167);
or U22470 (N_22470,N_19072,N_18618);
nor U22471 (N_22471,N_17683,N_19629);
or U22472 (N_22472,N_18832,N_18008);
or U22473 (N_22473,N_19527,N_18955);
nand U22474 (N_22474,N_18277,N_18067);
xnor U22475 (N_22475,N_19581,N_19020);
and U22476 (N_22476,N_18505,N_18934);
nand U22477 (N_22477,N_18644,N_18465);
or U22478 (N_22478,N_18548,N_19608);
nor U22479 (N_22479,N_18721,N_17543);
nor U22480 (N_22480,N_19408,N_17757);
nor U22481 (N_22481,N_17573,N_19367);
xnor U22482 (N_22482,N_19461,N_18867);
nand U22483 (N_22483,N_19473,N_19566);
or U22484 (N_22484,N_19176,N_19432);
or U22485 (N_22485,N_19682,N_19293);
xor U22486 (N_22486,N_18050,N_17597);
xor U22487 (N_22487,N_19744,N_17747);
nor U22488 (N_22488,N_18672,N_19046);
xor U22489 (N_22489,N_17524,N_18666);
or U22490 (N_22490,N_17777,N_19230);
and U22491 (N_22491,N_19559,N_18419);
and U22492 (N_22492,N_18325,N_18582);
and U22493 (N_22493,N_17829,N_17600);
nor U22494 (N_22494,N_17750,N_18329);
nor U22495 (N_22495,N_18498,N_18088);
nand U22496 (N_22496,N_18924,N_17736);
xnor U22497 (N_22497,N_17916,N_19941);
nor U22498 (N_22498,N_18842,N_18016);
nand U22499 (N_22499,N_19562,N_19960);
and U22500 (N_22500,N_21768,N_20410);
nor U22501 (N_22501,N_21801,N_21035);
or U22502 (N_22502,N_22123,N_20113);
nand U22503 (N_22503,N_20852,N_21157);
nor U22504 (N_22504,N_21477,N_20195);
or U22505 (N_22505,N_21616,N_20418);
nor U22506 (N_22506,N_21694,N_20180);
and U22507 (N_22507,N_21502,N_21970);
nor U22508 (N_22508,N_20109,N_20601);
xnor U22509 (N_22509,N_21987,N_21865);
or U22510 (N_22510,N_20786,N_21274);
nor U22511 (N_22511,N_20815,N_21332);
nor U22512 (N_22512,N_22332,N_21193);
or U22513 (N_22513,N_21137,N_20117);
xnor U22514 (N_22514,N_22219,N_20803);
and U22515 (N_22515,N_22242,N_20271);
nand U22516 (N_22516,N_21837,N_20255);
xnor U22517 (N_22517,N_20773,N_21037);
nor U22518 (N_22518,N_22241,N_20179);
or U22519 (N_22519,N_20997,N_21109);
xnor U22520 (N_22520,N_20343,N_21379);
nand U22521 (N_22521,N_21203,N_20915);
nor U22522 (N_22522,N_20533,N_22309);
xor U22523 (N_22523,N_21878,N_20867);
xor U22524 (N_22524,N_21337,N_21160);
or U22525 (N_22525,N_22213,N_21481);
and U22526 (N_22526,N_21453,N_20840);
nor U22527 (N_22527,N_20051,N_21336);
nor U22528 (N_22528,N_22279,N_21155);
nor U22529 (N_22529,N_20686,N_20695);
xnor U22530 (N_22530,N_21682,N_22128);
nand U22531 (N_22531,N_21738,N_20282);
and U22532 (N_22532,N_22196,N_21102);
nand U22533 (N_22533,N_20459,N_22456);
or U22534 (N_22534,N_21787,N_21285);
and U22535 (N_22535,N_22016,N_20505);
nand U22536 (N_22536,N_20743,N_21630);
and U22537 (N_22537,N_20835,N_21334);
xnor U22538 (N_22538,N_20037,N_21357);
and U22539 (N_22539,N_21222,N_21911);
nand U22540 (N_22540,N_21556,N_21007);
nor U22541 (N_22541,N_21542,N_22311);
nor U22542 (N_22542,N_22084,N_21942);
and U22543 (N_22543,N_20754,N_21255);
and U22544 (N_22544,N_22064,N_20643);
and U22545 (N_22545,N_21955,N_20536);
xor U22546 (N_22546,N_20245,N_20402);
xnor U22547 (N_22547,N_22207,N_20281);
nand U22548 (N_22548,N_21309,N_20588);
nand U22549 (N_22549,N_20989,N_20640);
nor U22550 (N_22550,N_21218,N_21093);
and U22551 (N_22551,N_21894,N_20224);
or U22552 (N_22552,N_20912,N_21087);
nand U22553 (N_22553,N_20242,N_22139);
or U22554 (N_22554,N_21692,N_20041);
xor U22555 (N_22555,N_20913,N_21647);
and U22556 (N_22556,N_21472,N_22007);
and U22557 (N_22557,N_20470,N_20373);
nand U22558 (N_22558,N_21963,N_20603);
xor U22559 (N_22559,N_20995,N_20991);
and U22560 (N_22560,N_20190,N_21289);
or U22561 (N_22561,N_20589,N_21983);
xnor U22562 (N_22562,N_20518,N_20009);
nand U22563 (N_22563,N_20352,N_21219);
nor U22564 (N_22564,N_21816,N_20246);
xor U22565 (N_22565,N_22440,N_20682);
nor U22566 (N_22566,N_20199,N_21235);
or U22567 (N_22567,N_20286,N_20710);
nand U22568 (N_22568,N_22075,N_20371);
nor U22569 (N_22569,N_22347,N_21762);
xor U22570 (N_22570,N_20907,N_21301);
nand U22571 (N_22571,N_22203,N_22237);
xor U22572 (N_22572,N_20326,N_21423);
nand U22573 (N_22573,N_20759,N_20049);
and U22574 (N_22574,N_21493,N_22074);
xor U22575 (N_22575,N_20765,N_20755);
nand U22576 (N_22576,N_22336,N_21018);
nand U22577 (N_22577,N_22323,N_21809);
and U22578 (N_22578,N_22466,N_21425);
nor U22579 (N_22579,N_20114,N_20504);
xor U22580 (N_22580,N_21943,N_21592);
or U22581 (N_22581,N_20723,N_20737);
xnor U22582 (N_22582,N_22149,N_20706);
nor U22583 (N_22583,N_21376,N_21196);
or U22584 (N_22584,N_21550,N_21587);
nor U22585 (N_22585,N_20095,N_20705);
and U22586 (N_22586,N_20489,N_20283);
or U22587 (N_22587,N_21088,N_20426);
or U22588 (N_22588,N_20464,N_22005);
nor U22589 (N_22589,N_20217,N_21695);
and U22590 (N_22590,N_22288,N_20893);
and U22591 (N_22591,N_20253,N_20374);
nor U22592 (N_22592,N_21934,N_21780);
and U22593 (N_22593,N_21112,N_20314);
nor U22594 (N_22594,N_22246,N_22226);
and U22595 (N_22595,N_20138,N_21818);
xnor U22596 (N_22596,N_22021,N_20626);
nand U22597 (N_22597,N_20628,N_21342);
or U22598 (N_22598,N_21628,N_22027);
nor U22599 (N_22599,N_21115,N_20007);
and U22600 (N_22600,N_21622,N_21217);
nand U22601 (N_22601,N_20622,N_22432);
nor U22602 (N_22602,N_20690,N_20455);
nor U22603 (N_22603,N_21709,N_21824);
nor U22604 (N_22604,N_20456,N_21779);
or U22605 (N_22605,N_21514,N_21030);
xor U22606 (N_22606,N_21494,N_20667);
nand U22607 (N_22607,N_22099,N_22201);
or U22608 (N_22608,N_21988,N_20977);
nor U22609 (N_22609,N_20508,N_20671);
or U22610 (N_22610,N_20918,N_20808);
or U22611 (N_22611,N_21677,N_21230);
and U22612 (N_22612,N_20409,N_21914);
xor U22613 (N_22613,N_22085,N_21887);
nor U22614 (N_22614,N_20430,N_20218);
nand U22615 (N_22615,N_20724,N_21060);
nand U22616 (N_22616,N_21169,N_22434);
xnor U22617 (N_22617,N_20053,N_21406);
nor U22618 (N_22618,N_20862,N_20019);
nor U22619 (N_22619,N_21004,N_20036);
xnor U22620 (N_22620,N_21864,N_20099);
and U22621 (N_22621,N_21516,N_22164);
xor U22622 (N_22622,N_21827,N_20482);
nand U22623 (N_22623,N_21318,N_21449);
and U22624 (N_22624,N_21908,N_20787);
nor U22625 (N_22625,N_22061,N_21131);
or U22626 (N_22626,N_20760,N_20770);
and U22627 (N_22627,N_21426,N_21774);
nor U22628 (N_22628,N_20944,N_20161);
and U22629 (N_22629,N_20685,N_20244);
xor U22630 (N_22630,N_20540,N_21295);
nor U22631 (N_22631,N_21765,N_22256);
and U22632 (N_22632,N_20527,N_21001);
or U22633 (N_22633,N_22211,N_22025);
xnor U22634 (N_22634,N_21948,N_22119);
xnor U22635 (N_22635,N_20390,N_20318);
and U22636 (N_22636,N_20549,N_21106);
xnor U22637 (N_22637,N_21547,N_20300);
or U22638 (N_22638,N_20919,N_21886);
nand U22639 (N_22639,N_22182,N_20845);
xnor U22640 (N_22640,N_21447,N_20794);
nor U22641 (N_22641,N_21436,N_22244);
and U22642 (N_22642,N_21796,N_21909);
nand U22643 (N_22643,N_20085,N_20726);
xor U22644 (N_22644,N_21511,N_22282);
nand U22645 (N_22645,N_22298,N_20309);
xor U22646 (N_22646,N_20216,N_22438);
nor U22647 (N_22647,N_22103,N_20783);
nand U22648 (N_22648,N_20250,N_20621);
nand U22649 (N_22649,N_20015,N_21811);
nand U22650 (N_22650,N_21287,N_21640);
and U22651 (N_22651,N_21052,N_20288);
or U22652 (N_22652,N_21536,N_22316);
xor U22653 (N_22653,N_20156,N_21851);
or U22654 (N_22654,N_22055,N_21933);
or U22655 (N_22655,N_21889,N_21114);
or U22656 (N_22656,N_21476,N_20499);
and U22657 (N_22657,N_22006,N_21050);
nand U22658 (N_22658,N_21445,N_20872);
or U22659 (N_22659,N_21444,N_22072);
xnor U22660 (N_22660,N_20564,N_21896);
xnor U22661 (N_22661,N_22215,N_20477);
xnor U22662 (N_22662,N_22014,N_20078);
and U22663 (N_22663,N_21140,N_21183);
xor U22664 (N_22664,N_20057,N_21746);
nand U22665 (N_22665,N_20132,N_21194);
and U22666 (N_22666,N_20481,N_20939);
and U22667 (N_22667,N_20859,N_20964);
and U22668 (N_22668,N_20292,N_22138);
nand U22669 (N_22669,N_21526,N_20897);
nor U22670 (N_22670,N_21068,N_20709);
xor U22671 (N_22671,N_20994,N_21280);
nor U22672 (N_22672,N_21058,N_22469);
nand U22673 (N_22673,N_22190,N_21316);
xnor U22674 (N_22674,N_20362,N_21797);
xor U22675 (N_22675,N_20970,N_20774);
xnor U22676 (N_22676,N_22093,N_21282);
and U22677 (N_22677,N_20507,N_20359);
nand U22678 (N_22678,N_22429,N_20045);
or U22679 (N_22679,N_21741,N_21186);
nor U22680 (N_22680,N_22296,N_20437);
nand U22681 (N_22681,N_20637,N_21517);
xnor U22682 (N_22682,N_21856,N_22461);
nand U22683 (N_22683,N_20833,N_21105);
nor U22684 (N_22684,N_20559,N_21044);
nand U22685 (N_22685,N_20448,N_22041);
xnor U22686 (N_22686,N_21043,N_20302);
nor U22687 (N_22687,N_20008,N_20384);
and U22688 (N_22688,N_20097,N_21191);
or U22689 (N_22689,N_21825,N_20098);
and U22690 (N_22690,N_21240,N_22161);
nand U22691 (N_22691,N_21339,N_20503);
nor U22692 (N_22692,N_21498,N_20818);
or U22693 (N_22693,N_21712,N_21792);
and U22694 (N_22694,N_22388,N_21271);
and U22695 (N_22695,N_21129,N_21515);
or U22696 (N_22696,N_22329,N_20162);
nor U22697 (N_22697,N_21854,N_20451);
nand U22698 (N_22698,N_22338,N_22216);
nor U22699 (N_22699,N_21045,N_21591);
or U22700 (N_22700,N_21957,N_21932);
or U22701 (N_22701,N_21788,N_21852);
and U22702 (N_22702,N_22303,N_21653);
nand U22703 (N_22703,N_22422,N_21099);
xnor U22704 (N_22704,N_22158,N_20752);
and U22705 (N_22705,N_21149,N_21294);
or U22706 (N_22706,N_20853,N_20945);
or U22707 (N_22707,N_20553,N_20379);
or U22708 (N_22708,N_21504,N_21321);
and U22709 (N_22709,N_22283,N_21973);
xor U22710 (N_22710,N_20822,N_21945);
and U22711 (N_22711,N_20609,N_22319);
nor U22712 (N_22712,N_21072,N_22271);
xnor U22713 (N_22713,N_21220,N_20050);
or U22714 (N_22714,N_20229,N_20896);
nor U22715 (N_22715,N_20812,N_20836);
or U22716 (N_22716,N_22108,N_20149);
nor U22717 (N_22717,N_21808,N_21693);
nor U22718 (N_22718,N_22094,N_20443);
and U22719 (N_22719,N_21995,N_21588);
nand U22720 (N_22720,N_21228,N_20804);
nor U22721 (N_22721,N_21944,N_20651);
nor U22722 (N_22722,N_20150,N_21234);
xnor U22723 (N_22723,N_21884,N_21179);
xor U22724 (N_22724,N_21659,N_22322);
or U22725 (N_22725,N_20625,N_21171);
or U22726 (N_22726,N_20535,N_20018);
xor U22727 (N_22727,N_20920,N_20164);
and U22728 (N_22728,N_20142,N_21118);
or U22729 (N_22729,N_20399,N_20328);
nor U22730 (N_22730,N_20335,N_21090);
or U22731 (N_22731,N_20882,N_21290);
and U22732 (N_22732,N_21688,N_20337);
and U22733 (N_22733,N_20979,N_20642);
or U22734 (N_22734,N_22386,N_21200);
nand U22735 (N_22735,N_21078,N_20004);
nand U22736 (N_22736,N_21159,N_22290);
xor U22737 (N_22737,N_21019,N_20675);
or U22738 (N_22738,N_20345,N_20986);
nor U22739 (N_22739,N_21690,N_20073);
or U22740 (N_22740,N_22494,N_22328);
nor U22741 (N_22741,N_20147,N_21315);
and U22742 (N_22742,N_20312,N_20060);
nand U22743 (N_22743,N_21008,N_21313);
nor U22744 (N_22744,N_21325,N_20821);
xnor U22745 (N_22745,N_21360,N_20899);
or U22746 (N_22746,N_20076,N_20412);
xor U22747 (N_22747,N_20629,N_21980);
nand U22748 (N_22748,N_20084,N_20116);
or U22749 (N_22749,N_20093,N_21091);
and U22750 (N_22750,N_21654,N_20171);
or U22751 (N_22751,N_21966,N_21362);
or U22752 (N_22752,N_21836,N_21717);
and U22753 (N_22753,N_21495,N_21507);
and U22754 (N_22754,N_21446,N_21976);
and U22755 (N_22755,N_21789,N_22496);
or U22756 (N_22756,N_20475,N_20360);
nor U22757 (N_22757,N_22384,N_21311);
nor U22758 (N_22758,N_20140,N_22491);
and U22759 (N_22759,N_22333,N_21919);
and U22760 (N_22760,N_20168,N_20198);
and U22761 (N_22761,N_20059,N_20886);
xnor U22762 (N_22762,N_20157,N_20181);
nand U22763 (N_22763,N_20988,N_21113);
or U22764 (N_22764,N_21241,N_22208);
or U22765 (N_22765,N_20120,N_21522);
or U22766 (N_22766,N_20397,N_21278);
or U22767 (N_22767,N_22160,N_21519);
and U22768 (N_22768,N_21602,N_22417);
or U22769 (N_22769,N_20696,N_21211);
nor U22770 (N_22770,N_20809,N_20110);
nor U22771 (N_22771,N_21960,N_22243);
or U22772 (N_22772,N_21405,N_21916);
nor U22773 (N_22773,N_20514,N_21177);
nor U22774 (N_22774,N_20405,N_21303);
nor U22775 (N_22775,N_20884,N_21664);
or U22776 (N_22776,N_20347,N_20056);
or U22777 (N_22777,N_20829,N_21513);
nand U22778 (N_22778,N_21915,N_20781);
xor U22779 (N_22779,N_20903,N_21197);
nand U22780 (N_22780,N_22273,N_21882);
or U22781 (N_22781,N_21707,N_20584);
and U22782 (N_22782,N_21804,N_20513);
or U22783 (N_22783,N_20673,N_22212);
nor U22784 (N_22784,N_21949,N_22487);
nand U22785 (N_22785,N_22472,N_20129);
and U22786 (N_22786,N_20052,N_22033);
xor U22787 (N_22787,N_20606,N_22231);
xnor U22788 (N_22788,N_21040,N_22086);
nand U22789 (N_22789,N_21572,N_20728);
nand U22790 (N_22790,N_22034,N_20252);
nor U22791 (N_22791,N_21668,N_20233);
nor U22792 (N_22792,N_20515,N_21488);
and U22793 (N_22793,N_21126,N_21400);
nor U22794 (N_22794,N_21898,N_20516);
or U22795 (N_22795,N_20294,N_21953);
nand U22796 (N_22796,N_21273,N_21799);
nor U22797 (N_22797,N_21902,N_21431);
nor U22798 (N_22798,N_20058,N_20376);
or U22799 (N_22799,N_20869,N_22066);
nor U22800 (N_22800,N_20998,N_20074);
nor U22801 (N_22801,N_21028,N_21633);
or U22802 (N_22802,N_20207,N_20943);
or U22803 (N_22803,N_20555,N_21681);
and U22804 (N_22804,N_21680,N_21739);
nand U22805 (N_22805,N_20256,N_20429);
nor U22806 (N_22806,N_20068,N_21501);
and U22807 (N_22807,N_21358,N_20580);
nor U22808 (N_22808,N_21039,N_21086);
xor U22809 (N_22809,N_21466,N_20123);
xnor U22810 (N_22810,N_20700,N_22098);
nor U22811 (N_22811,N_20856,N_21356);
and U22812 (N_22812,N_22156,N_20756);
or U22813 (N_22813,N_22077,N_21540);
and U22814 (N_22814,N_21951,N_20526);
nand U22815 (N_22815,N_20725,N_20389);
or U22816 (N_22816,N_21393,N_21691);
xor U22817 (N_22817,N_20289,N_20023);
and U22818 (N_22818,N_20296,N_21785);
or U22819 (N_22819,N_21706,N_20226);
nor U22820 (N_22820,N_22399,N_20954);
nand U22821 (N_22821,N_20131,N_22143);
nand U22822 (N_22822,N_22278,N_22425);
nor U22823 (N_22823,N_20623,N_21564);
and U22824 (N_22824,N_20054,N_20635);
and U22825 (N_22825,N_20571,N_21333);
or U22826 (N_22826,N_22299,N_20680);
xnor U22827 (N_22827,N_20934,N_20687);
nand U22828 (N_22828,N_21868,N_22162);
nor U22829 (N_22829,N_20485,N_20802);
xor U22830 (N_22830,N_21010,N_22439);
and U22831 (N_22831,N_22222,N_22307);
nor U22832 (N_22832,N_21270,N_20452);
nor U22833 (N_22833,N_21998,N_21512);
and U22834 (N_22834,N_20987,N_21736);
nor U22835 (N_22835,N_21450,N_21428);
xnor U22836 (N_22836,N_22046,N_20428);
xnor U22837 (N_22837,N_21604,N_20611);
or U22838 (N_22838,N_20153,N_21246);
and U22839 (N_22839,N_21139,N_21745);
and U22840 (N_22840,N_21631,N_22266);
nand U22841 (N_22841,N_20031,N_20519);
nand U22842 (N_22842,N_22415,N_22154);
nor U22843 (N_22843,N_22252,N_20599);
and U22844 (N_22844,N_22489,N_20320);
nand U22845 (N_22845,N_22267,N_21958);
xnor U22846 (N_22846,N_22492,N_20938);
xor U22847 (N_22847,N_21097,N_22441);
and U22848 (N_22848,N_21831,N_21355);
nor U22849 (N_22849,N_20187,N_20435);
nor U22850 (N_22850,N_21154,N_21243);
and U22851 (N_22851,N_20735,N_22248);
nor U22852 (N_22852,N_20024,N_20581);
or U22853 (N_22853,N_21952,N_20354);
nand U22854 (N_22854,N_20895,N_20119);
xnor U22855 (N_22855,N_21569,N_20220);
nand U22856 (N_22856,N_22305,N_21705);
nand U22857 (N_22857,N_22214,N_20742);
nand U22858 (N_22858,N_21221,N_20324);
and U22859 (N_22859,N_22010,N_22452);
and U22860 (N_22860,N_21407,N_21857);
xnor U22861 (N_22861,N_22285,N_21317);
nor U22862 (N_22862,N_20194,N_21394);
or U22863 (N_22863,N_20063,N_20096);
xor U22864 (N_22864,N_20957,N_22331);
nor U22865 (N_22865,N_22312,N_20796);
nand U22866 (N_22866,N_21065,N_20105);
or U22867 (N_22867,N_20666,N_20849);
or U22868 (N_22868,N_21648,N_21991);
nor U22869 (N_22869,N_20883,N_21763);
and U22870 (N_22870,N_20414,N_21761);
and U22871 (N_22871,N_20887,N_21267);
and U22872 (N_22872,N_20670,N_20841);
and U22873 (N_22873,N_21467,N_21213);
nand U22874 (N_22874,N_21208,N_21686);
or U22875 (N_22875,N_21665,N_21810);
nand U22876 (N_22876,N_20958,N_21192);
nand U22877 (N_22877,N_22277,N_20016);
nor U22878 (N_22878,N_21275,N_21924);
and U22879 (N_22879,N_21083,N_20222);
nand U22880 (N_22880,N_20243,N_21667);
nor U22881 (N_22881,N_20453,N_21245);
nand U22882 (N_22882,N_22169,N_20871);
nand U22883 (N_22883,N_21612,N_20424);
xor U22884 (N_22884,N_21263,N_20863);
nor U22885 (N_22885,N_21474,N_22166);
nand U22886 (N_22886,N_20971,N_21624);
nand U22887 (N_22887,N_21594,N_21875);
xnor U22888 (N_22888,N_21331,N_20740);
or U22889 (N_22889,N_20419,N_20614);
nand U22890 (N_22890,N_22327,N_20681);
xnor U22891 (N_22891,N_22374,N_21229);
or U22892 (N_22892,N_20922,N_21098);
and U22893 (N_22893,N_22258,N_22498);
nand U22894 (N_22894,N_20088,N_21568);
nand U22895 (N_22895,N_20319,N_21092);
or U22896 (N_22896,N_20619,N_22484);
or U22897 (N_22897,N_21253,N_22454);
and U22898 (N_22898,N_21735,N_20751);
and U22899 (N_22899,N_21080,N_21020);
nor U22900 (N_22900,N_21181,N_22462);
nor U22901 (N_22901,N_22102,N_21702);
nor U22902 (N_22902,N_20657,N_21757);
xor U22903 (N_22903,N_20502,N_21666);
and U22904 (N_22904,N_21462,N_21926);
nand U22905 (N_22905,N_20631,N_21299);
nor U22906 (N_22906,N_21657,N_20279);
nand U22907 (N_22907,N_21907,N_22050);
and U22908 (N_22908,N_21254,N_20231);
nor U22909 (N_22909,N_20573,N_21150);
nor U22910 (N_22910,N_20738,N_22039);
or U22911 (N_22911,N_22057,N_21893);
or U22912 (N_22912,N_21658,N_22120);
and U22913 (N_22913,N_20228,N_20043);
or U22914 (N_22914,N_21642,N_20102);
or U22915 (N_22915,N_21800,N_20368);
and U22916 (N_22916,N_21881,N_20684);
or U22917 (N_22917,N_20427,N_21180);
xnor U22918 (N_22918,N_21188,N_21417);
nand U22919 (N_22919,N_21152,N_22192);
and U22920 (N_22920,N_20947,N_21390);
nand U22921 (N_22921,N_20258,N_22340);
xnor U22922 (N_22922,N_22470,N_21863);
or U22923 (N_22923,N_20425,N_21589);
nand U22924 (N_22924,N_22205,N_21034);
nor U22925 (N_22925,N_22089,N_21729);
xor U22926 (N_22926,N_21125,N_20590);
or U22927 (N_22927,N_21326,N_21500);
or U22928 (N_22928,N_21017,N_21482);
nand U22929 (N_22929,N_20612,N_20870);
nor U22930 (N_22930,N_20366,N_21162);
nor U22931 (N_22931,N_21912,N_21012);
nand U22932 (N_22932,N_22381,N_20472);
or U22933 (N_22933,N_20664,N_22315);
xnor U22934 (N_22934,N_22037,N_20926);
and U22935 (N_22935,N_20607,N_21764);
or U22936 (N_22936,N_21369,N_20811);
and U22937 (N_22937,N_21720,N_21530);
nor U22938 (N_22938,N_20185,N_21670);
nand U22939 (N_22939,N_21669,N_21448);
nor U22940 (N_22940,N_22326,N_21343);
or U22941 (N_22941,N_22485,N_21610);
nor U22942 (N_22942,N_20177,N_20627);
nor U22943 (N_22943,N_20145,N_22030);
nor U22944 (N_22944,N_20984,N_22132);
nand U22945 (N_22945,N_21031,N_21936);
nor U22946 (N_22946,N_21110,N_22349);
and U22947 (N_22947,N_20949,N_21967);
and U22948 (N_22948,N_20904,N_21901);
and U22949 (N_22949,N_21861,N_21575);
nand U22950 (N_22950,N_20188,N_21554);
and U22951 (N_22951,N_22183,N_22024);
nand U22952 (N_22952,N_22351,N_20107);
nand U22953 (N_22953,N_21307,N_20163);
and U22954 (N_22954,N_20771,N_22180);
or U22955 (N_22955,N_20081,N_21121);
or U22956 (N_22956,N_20062,N_22097);
nand U22957 (N_22957,N_22369,N_22223);
nand U22958 (N_22958,N_22082,N_21024);
nor U22959 (N_22959,N_21615,N_21079);
and U22960 (N_22960,N_21580,N_21605);
xor U22961 (N_22961,N_20510,N_22393);
and U22962 (N_22962,N_22379,N_20261);
or U22963 (N_22963,N_22435,N_22382);
nand U22964 (N_22964,N_22136,N_21509);
nand U22965 (N_22965,N_20757,N_20511);
and U22966 (N_22966,N_20386,N_22269);
xnor U22967 (N_22967,N_20247,N_20950);
nor U22968 (N_22968,N_21470,N_21921);
nor U22969 (N_22969,N_21869,N_21750);
and U22970 (N_22970,N_20227,N_20476);
or U22971 (N_22971,N_22090,N_20933);
nor U22972 (N_22972,N_20674,N_20520);
or U22973 (N_22973,N_21259,N_21850);
or U22974 (N_22974,N_20285,N_20763);
xor U22975 (N_22975,N_20531,N_22181);
and U22976 (N_22976,N_21608,N_21899);
nand U22977 (N_22977,N_22083,N_22483);
nor U22978 (N_22978,N_20239,N_20259);
or U22979 (N_22979,N_20493,N_22481);
nand U22980 (N_22980,N_20509,N_21158);
xnor U22981 (N_22981,N_22165,N_20963);
and U22982 (N_22982,N_21085,N_20273);
xnor U22983 (N_22983,N_21650,N_21742);
xor U22984 (N_22984,N_21204,N_22359);
and U22985 (N_22985,N_20931,N_21016);
or U22986 (N_22986,N_20800,N_22076);
or U22987 (N_22987,N_20557,N_21918);
or U22988 (N_22988,N_20878,N_22051);
nor U22989 (N_22989,N_21528,N_20965);
nor U22990 (N_22990,N_21728,N_22352);
xor U22991 (N_22991,N_21523,N_20322);
nor U22992 (N_22992,N_20436,N_21871);
and U22993 (N_22993,N_21485,N_21535);
xor U22994 (N_22994,N_22345,N_20544);
and U22995 (N_22995,N_22253,N_21561);
nor U22996 (N_22996,N_20972,N_21541);
and U22997 (N_22997,N_20235,N_20383);
and U22998 (N_22998,N_20423,N_21141);
nor U22999 (N_22999,N_22360,N_20914);
or U23000 (N_23000,N_21128,N_20290);
nor U23001 (N_23001,N_21286,N_22247);
xor U23002 (N_23002,N_20329,N_20567);
or U23003 (N_23003,N_21329,N_21619);
nand U23004 (N_23004,N_21418,N_20075);
nand U23005 (N_23005,N_20466,N_20025);
nor U23006 (N_23006,N_22346,N_22317);
nor U23007 (N_23007,N_21821,N_20183);
nand U23008 (N_23008,N_20167,N_21258);
and U23009 (N_23009,N_21974,N_20370);
nor U23010 (N_23010,N_22175,N_21938);
xnor U23011 (N_23011,N_21860,N_20134);
nand U23012 (N_23012,N_22060,N_20197);
or U23013 (N_23013,N_20730,N_22047);
xor U23014 (N_23014,N_20122,N_22117);
and U23015 (N_23015,N_22421,N_21011);
or U23016 (N_23016,N_20813,N_20395);
nor U23017 (N_23017,N_20942,N_22125);
xor U23018 (N_23018,N_20624,N_20638);
nor U23019 (N_23019,N_20141,N_22199);
nor U23020 (N_23020,N_21276,N_21798);
or U23021 (N_23021,N_21617,N_21661);
or U23022 (N_23022,N_20316,N_22071);
and U23023 (N_23023,N_21009,N_22091);
nand U23024 (N_23024,N_21176,N_21490);
xor U23025 (N_23025,N_22363,N_22176);
and U23026 (N_23026,N_20708,N_21782);
xnor U23027 (N_23027,N_21826,N_22420);
nor U23028 (N_23028,N_20556,N_20441);
xnor U23029 (N_23029,N_21817,N_21747);
and U23030 (N_23030,N_21338,N_20574);
xor U23031 (N_23031,N_22163,N_21056);
nor U23032 (N_23032,N_20020,N_21929);
or U23033 (N_23033,N_20035,N_21636);
or U23034 (N_23034,N_21127,N_21231);
xnor U23035 (N_23035,N_20980,N_20387);
nand U23036 (N_23036,N_22092,N_22455);
nand U23037 (N_23037,N_21135,N_22320);
xnor U23038 (N_23038,N_22294,N_22095);
or U23039 (N_23039,N_22357,N_21855);
xor U23040 (N_23040,N_21537,N_21582);
or U23041 (N_23041,N_20034,N_22257);
xnor U23042 (N_23042,N_22043,N_21460);
nand U23043 (N_23043,N_21730,N_22453);
nor U23044 (N_23044,N_20065,N_20659);
or U23045 (N_23045,N_20001,N_20061);
nand U23046 (N_23046,N_20750,N_22054);
xnor U23047 (N_23047,N_22459,N_22339);
or U23048 (N_23048,N_22121,N_20275);
or U23049 (N_23049,N_21441,N_20850);
nor U23050 (N_23050,N_21940,N_21382);
nand U23051 (N_23051,N_20468,N_21662);
xor U23052 (N_23052,N_21433,N_20780);
nor U23053 (N_23053,N_20240,N_21845);
nand U23054 (N_23054,N_21473,N_20669);
xor U23055 (N_23055,N_21409,N_20033);
nor U23056 (N_23056,N_20003,N_21454);
nand U23057 (N_23057,N_20653,N_21835);
or U23058 (N_23058,N_20948,N_21496);
and U23059 (N_23059,N_22159,N_21373);
and U23060 (N_23060,N_22184,N_21041);
nor U23061 (N_23061,N_21293,N_21471);
or U23062 (N_23062,N_20828,N_21754);
or U23063 (N_23063,N_22022,N_20576);
or U23064 (N_23064,N_20421,N_21880);
or U23065 (N_23065,N_20694,N_22414);
nor U23066 (N_23066,N_20413,N_22449);
nand U23067 (N_23067,N_20866,N_20940);
nand U23068 (N_23068,N_21212,N_21236);
and U23069 (N_23069,N_20982,N_20824);
nand U23070 (N_23070,N_21252,N_22284);
xor U23071 (N_23071,N_20665,N_21145);
nor U23072 (N_23072,N_20814,N_21146);
nor U23073 (N_23073,N_22234,N_22146);
and U23074 (N_23074,N_20407,N_21443);
nand U23075 (N_23075,N_22073,N_21248);
and U23076 (N_23076,N_22001,N_21609);
nor U23077 (N_23077,N_20342,N_21885);
and U23078 (N_23078,N_21451,N_21546);
nor U23079 (N_23079,N_21344,N_21993);
xnor U23080 (N_23080,N_21377,N_22080);
or U23081 (N_23081,N_21368,N_22088);
nand U23082 (N_23082,N_21698,N_21941);
nand U23083 (N_23083,N_21876,N_20166);
and U23084 (N_23084,N_22350,N_22144);
nand U23085 (N_23085,N_20369,N_20039);
xor U23086 (N_23086,N_20269,N_21385);
or U23087 (N_23087,N_22155,N_20234);
nor U23088 (N_23088,N_21296,N_20215);
nor U23089 (N_23089,N_21770,N_20325);
or U23090 (N_23090,N_20720,N_21363);
xor U23091 (N_23091,N_20064,N_21756);
and U23092 (N_23092,N_20909,N_22259);
and U23093 (N_23093,N_22000,N_22306);
nand U23094 (N_23094,N_20960,N_20471);
nand U23095 (N_23095,N_20565,N_20563);
nand U23096 (N_23096,N_20568,N_22118);
xnor U23097 (N_23097,N_21256,N_21320);
xor U23098 (N_23098,N_20363,N_22488);
xor U23099 (N_23099,N_21718,N_21237);
nand U23100 (N_23100,N_22126,N_20586);
nand U23101 (N_23101,N_20906,N_21820);
or U23102 (N_23102,N_22035,N_20610);
xor U23103 (N_23103,N_21366,N_21000);
nand U23104 (N_23104,N_21434,N_20501);
nand U23105 (N_23105,N_20582,N_20767);
nand U23106 (N_23106,N_20721,N_22334);
nand U23107 (N_23107,N_20873,N_22291);
nor U23108 (N_23108,N_21063,N_22437);
and U23109 (N_23109,N_20952,N_20332);
nor U23110 (N_23110,N_21215,N_21905);
nor U23111 (N_23111,N_20301,N_22238);
and U23112 (N_23112,N_21552,N_21675);
nand U23113 (N_23113,N_21689,N_20600);
xnor U23114 (N_23114,N_22191,N_21478);
nor U23115 (N_23115,N_21773,N_20956);
or U23116 (N_23116,N_22371,N_22368);
and U23117 (N_23117,N_22008,N_21853);
nand U23118 (N_23118,N_21025,N_21383);
and U23119 (N_23119,N_21365,N_20701);
nor U23120 (N_23120,N_21722,N_20978);
and U23121 (N_23121,N_22134,N_22408);
nor U23122 (N_23122,N_20570,N_20077);
nor U23123 (N_23123,N_20898,N_20858);
or U23124 (N_23124,N_20173,N_20839);
xnor U23125 (N_23125,N_22375,N_21674);
and U23126 (N_23126,N_20500,N_21716);
and U23127 (N_23127,N_20592,N_21656);
nor U23128 (N_23128,N_22141,N_22113);
or U23129 (N_23129,N_21607,N_21913);
xor U23130 (N_23130,N_20011,N_22302);
and U23131 (N_23131,N_22362,N_20356);
or U23132 (N_23132,N_21981,N_20676);
xor U23133 (N_23133,N_21671,N_20434);
xnor U23134 (N_23134,N_21961,N_21767);
nor U23135 (N_23135,N_20241,N_21205);
xnor U23136 (N_23136,N_21806,N_20985);
nand U23137 (N_23137,N_21904,N_21027);
nand U23138 (N_23138,N_22321,N_20561);
nor U23139 (N_23139,N_22036,N_21053);
and U23140 (N_23140,N_21210,N_21758);
or U23141 (N_23141,N_21984,N_21897);
nor U23142 (N_23142,N_20784,N_21364);
nand U23143 (N_23143,N_21209,N_22049);
and U23144 (N_23144,N_20154,N_21330);
nand U23145 (N_23145,N_20512,N_20826);
nand U23146 (N_23146,N_20254,N_20083);
nand U23147 (N_23147,N_20716,N_20875);
and U23148 (N_23148,N_22018,N_21769);
nor U23149 (N_23149,N_21463,N_21538);
xor U23150 (N_23150,N_21378,N_21581);
and U23151 (N_23151,N_20474,N_21566);
nor U23152 (N_23152,N_21927,N_20506);
nor U23153 (N_23153,N_20308,N_22400);
and U23154 (N_23154,N_20894,N_22272);
xnor U23155 (N_23155,N_21148,N_20733);
and U23156 (N_23156,N_22402,N_21094);
or U23157 (N_23157,N_21283,N_20479);
or U23158 (N_23158,N_21432,N_21062);
and U23159 (N_23159,N_20311,N_20223);
nor U23160 (N_23160,N_22474,N_21081);
xor U23161 (N_23161,N_22465,N_21895);
xnor U23162 (N_23162,N_21752,N_22067);
and U23163 (N_23163,N_20966,N_22101);
and U23164 (N_23164,N_22372,N_22418);
nor U23165 (N_23165,N_20213,N_20346);
and U23166 (N_23166,N_20293,N_20917);
xor U23167 (N_23167,N_21822,N_21807);
and U23168 (N_23168,N_21892,N_21663);
or U23169 (N_23169,N_21288,N_21725);
or U23170 (N_23170,N_22228,N_21573);
and U23171 (N_23171,N_22416,N_21392);
xnor U23172 (N_23172,N_20480,N_21786);
and U23173 (N_23173,N_21819,N_20248);
xnor U23174 (N_23174,N_20633,N_20983);
nand U23175 (N_23175,N_22127,N_20608);
nand U23176 (N_23176,N_20729,N_21802);
and U23177 (N_23177,N_20923,N_20650);
and U23178 (N_23178,N_21638,N_21651);
nand U23179 (N_23179,N_20572,N_21070);
nand U23180 (N_23180,N_20593,N_21557);
or U23181 (N_23181,N_21888,N_21147);
nor U23182 (N_23182,N_21601,N_21543);
nand U23183 (N_23183,N_20048,N_20543);
and U23184 (N_23184,N_20837,N_22068);
or U23185 (N_23185,N_20927,N_20072);
or U23186 (N_23186,N_21322,N_21634);
nor U23187 (N_23187,N_21866,N_21046);
nand U23188 (N_23188,N_21075,N_20127);
nor U23189 (N_23189,N_20365,N_21082);
or U23190 (N_23190,N_21185,N_20449);
nor U23191 (N_23191,N_20272,N_21175);
or U23192 (N_23192,N_21429,N_21989);
and U23193 (N_23193,N_20203,N_21521);
xor U23194 (N_23194,N_20375,N_20736);
nand U23195 (N_23195,N_22364,N_20587);
nand U23196 (N_23196,N_22318,N_21372);
xnor U23197 (N_23197,N_20617,N_20406);
and U23198 (N_23198,N_20495,N_20225);
nand U23199 (N_23199,N_20487,N_20021);
nor U23200 (N_23200,N_20645,N_21743);
nand U23201 (N_23201,N_20692,N_22356);
xnor U23202 (N_23202,N_22056,N_21959);
or U23203 (N_23203,N_20274,N_21348);
nor U23204 (N_23204,N_20046,N_20753);
nor U23205 (N_23205,N_22142,N_21401);
xor U23206 (N_23206,N_21910,N_20172);
or U23207 (N_23207,N_20277,N_20398);
or U23208 (N_23208,N_22063,N_21047);
or U23209 (N_23209,N_21996,N_21759);
nand U23210 (N_23210,N_22087,N_21161);
xor U23211 (N_23211,N_20126,N_21266);
or U23212 (N_23212,N_21384,N_20848);
nor U23213 (N_23213,N_20026,N_22115);
nor U23214 (N_23214,N_22314,N_21104);
nor U23215 (N_23215,N_20355,N_20178);
xnor U23216 (N_23216,N_20394,N_20758);
or U23217 (N_23217,N_20598,N_22264);
xor U23218 (N_23218,N_20295,N_20200);
nand U23219 (N_23219,N_21051,N_22275);
or U23220 (N_23220,N_21599,N_20646);
or U23221 (N_23221,N_21968,N_22195);
and U23222 (N_23222,N_20558,N_20490);
and U23223 (N_23223,N_21833,N_20941);
or U23224 (N_23224,N_21071,N_20974);
and U23225 (N_23225,N_21142,N_21840);
nor U23226 (N_23226,N_20577,N_22262);
nand U23227 (N_23227,N_21655,N_22245);
xnor U23228 (N_23228,N_21388,N_22444);
or U23229 (N_23229,N_21397,N_21842);
xor U23230 (N_23230,N_20440,N_20491);
nand U23231 (N_23231,N_21794,N_21903);
xor U23232 (N_23232,N_21111,N_22229);
and U23233 (N_23233,N_21260,N_21458);
nand U23234 (N_23234,N_21437,N_20496);
and U23235 (N_23235,N_21464,N_22482);
nand U23236 (N_23236,N_20569,N_22059);
and U23237 (N_23237,N_22137,N_20438);
and U23238 (N_23238,N_22153,N_20137);
nor U23239 (N_23239,N_22450,N_22499);
xor U23240 (N_23240,N_20842,N_21107);
or U23241 (N_23241,N_22287,N_22020);
or U23242 (N_23242,N_22194,N_21077);
nand U23243 (N_23243,N_21165,N_21975);
xor U23244 (N_23244,N_20400,N_22204);
nor U23245 (N_23245,N_22308,N_22286);
and U23246 (N_23246,N_22017,N_20597);
and U23247 (N_23247,N_22401,N_20890);
and U23248 (N_23248,N_22497,N_20778);
xor U23249 (N_23249,N_22404,N_21074);
and U23250 (N_23250,N_21710,N_21947);
nand U23251 (N_23251,N_21922,N_21781);
nor U23252 (N_23252,N_20091,N_20125);
xnor U23253 (N_23253,N_22009,N_22174);
xor U23254 (N_23254,N_21928,N_21354);
nand U23255 (N_23255,N_21678,N_20575);
or U23256 (N_23256,N_21262,N_21803);
and U23257 (N_23257,N_20660,N_21562);
nand U23258 (N_23258,N_22254,N_22265);
or U23259 (N_23259,N_22168,N_20251);
nor U23260 (N_23260,N_22457,N_20932);
xor U23261 (N_23261,N_20844,N_22343);
and U23262 (N_23262,N_20731,N_21595);
xor U23263 (N_23263,N_22032,N_21297);
xor U23264 (N_23264,N_20522,N_21867);
or U23265 (N_23265,N_21497,N_21224);
xor U23266 (N_23266,N_20315,N_20422);
nor U23267 (N_23267,N_21719,N_20017);
nand U23268 (N_23268,N_21122,N_20266);
nor U23269 (N_23269,N_20953,N_21603);
nand U23270 (N_23270,N_21772,N_20539);
or U23271 (N_23271,N_22433,N_20268);
or U23272 (N_23272,N_22427,N_20930);
or U23273 (N_23273,N_21351,N_20854);
or U23274 (N_23274,N_22045,N_20469);
nand U23275 (N_23275,N_20816,N_21214);
or U23276 (N_23276,N_22377,N_20566);
or U23277 (N_23277,N_21873,N_21032);
and U23278 (N_23278,N_20946,N_21304);
or U23279 (N_23279,N_21347,N_22413);
nand U23280 (N_23280,N_21784,N_20392);
and U23281 (N_23281,N_20679,N_20658);
xor U23282 (N_23282,N_20196,N_20652);
xnor U23283 (N_23283,N_22129,N_20381);
xor U23284 (N_23284,N_20718,N_20578);
and U23285 (N_23285,N_20420,N_22140);
nand U23286 (N_23286,N_22240,N_22394);
xor U23287 (N_23287,N_20212,N_20317);
and U23288 (N_23288,N_20079,N_22387);
nor U23289 (N_23289,N_20595,N_20662);
xor U23290 (N_23290,N_21151,N_20776);
xnor U23291 (N_23291,N_22002,N_20892);
nand U23292 (N_23292,N_20417,N_20094);
and U23293 (N_23293,N_20935,N_21626);
and U23294 (N_23294,N_22411,N_20560);
or U23295 (N_23295,N_22335,N_21570);
nor U23296 (N_23296,N_21997,N_21697);
or U23297 (N_23297,N_21832,N_21906);
xnor U23298 (N_23298,N_20022,N_20851);
nor U23299 (N_23299,N_20792,N_20267);
xor U23300 (N_23300,N_21199,N_21503);
or U23301 (N_23301,N_22383,N_20101);
or U23302 (N_23302,N_20367,N_20210);
or U23303 (N_23303,N_21300,N_22013);
xnor U23304 (N_23304,N_20703,N_22116);
xnor U23305 (N_23305,N_22423,N_20276);
nor U23306 (N_23306,N_22185,N_21133);
nor U23307 (N_23307,N_21173,N_20372);
or U23308 (N_23308,N_21900,N_20924);
or U23309 (N_23309,N_21830,N_22152);
nand U23310 (N_23310,N_20976,N_22109);
nor U23311 (N_23311,N_20298,N_20432);
and U23312 (N_23312,N_20029,N_20916);
nand U23313 (N_23313,N_20005,N_20121);
nand U23314 (N_23314,N_21103,N_22385);
or U23315 (N_23315,N_22111,N_20801);
or U23316 (N_23316,N_22031,N_20361);
and U23317 (N_23317,N_21969,N_20937);
and U23318 (N_23318,N_21487,N_21683);
nor U23319 (N_23319,N_21491,N_20182);
nor U23320 (N_23320,N_21265,N_21715);
or U23321 (N_23321,N_22397,N_21226);
nor U23322 (N_23322,N_21563,N_20214);
or U23323 (N_23323,N_22424,N_21123);
or U23324 (N_23324,N_21558,N_20905);
nand U23325 (N_23325,N_22062,N_21734);
nand U23326 (N_23326,N_20151,N_22430);
xnor U23327 (N_23327,N_22232,N_21042);
nor U23328 (N_23328,N_21006,N_21101);
or U23329 (N_23329,N_21328,N_21057);
nand U23330 (N_23330,N_20378,N_20739);
nor U23331 (N_23331,N_20827,N_22167);
xnor U23332 (N_23332,N_21277,N_20663);
xnor U23333 (N_23333,N_21048,N_22490);
or U23334 (N_23334,N_21954,N_20688);
xor U23335 (N_23335,N_20111,N_22220);
or U23336 (N_23336,N_21962,N_22366);
nand U23337 (N_23337,N_21415,N_20713);
or U23338 (N_23338,N_20331,N_20146);
xor U23339 (N_23339,N_20656,N_22324);
or U23340 (N_23340,N_21755,N_21163);
nor U23341 (N_23341,N_21791,N_21422);
or U23342 (N_23342,N_21410,N_21917);
nor U23343 (N_23343,N_20284,N_20955);
or U23344 (N_23344,N_21069,N_20401);
nand U23345 (N_23345,N_21251,N_22405);
xnor U23346 (N_23346,N_20602,N_20152);
xnor U23347 (N_23347,N_22239,N_21021);
nand U23348 (N_23348,N_21858,N_20461);
nor U23349 (N_23349,N_20541,N_20678);
nor U23350 (N_23350,N_21760,N_20962);
nor U23351 (N_23351,N_20462,N_21054);
or U23352 (N_23352,N_22187,N_20494);
xnor U23353 (N_23353,N_20969,N_21416);
nor U23354 (N_23354,N_21189,N_21396);
nor U23355 (N_23355,N_21812,N_22249);
or U23356 (N_23356,N_21727,N_21775);
nand U23357 (N_23357,N_22354,N_22358);
or U23358 (N_23358,N_20820,N_21015);
nor U23359 (N_23359,N_21778,N_22106);
xor U23360 (N_23360,N_21244,N_21660);
or U23361 (N_23361,N_20585,N_20175);
or U23362 (N_23362,N_20902,N_20785);
xor U23363 (N_23363,N_20596,N_20170);
and U23364 (N_23364,N_22476,N_21269);
xor U23365 (N_23365,N_20825,N_21777);
or U23366 (N_23366,N_20691,N_22003);
and U23367 (N_23367,N_20699,N_20348);
nand U23368 (N_23368,N_21144,N_21598);
or U23369 (N_23369,N_20880,N_20358);
nand U23370 (N_23370,N_22260,N_21323);
nand U23371 (N_23371,N_21849,N_22304);
nand U23372 (N_23372,N_21033,N_20169);
nor U23373 (N_23373,N_21308,N_20069);
nor U23374 (N_23374,N_20087,N_21153);
or U23375 (N_23375,N_21749,N_21925);
xnor U23376 (N_23376,N_20865,N_21402);
xor U23377 (N_23377,N_21468,N_20551);
and U23378 (N_23378,N_20265,N_21076);
nand U23379 (N_23379,N_22147,N_20613);
and U23380 (N_23380,N_20351,N_21585);
xor U23381 (N_23381,N_21279,N_20761);
xor U23382 (N_23382,N_22281,N_21838);
or U23383 (N_23383,N_20634,N_21859);
nand U23384 (N_23384,N_21232,N_21687);
nor U23385 (N_23385,N_21411,N_21751);
and U23386 (N_23386,N_21371,N_21284);
nor U23387 (N_23387,N_21946,N_21699);
or U23388 (N_23388,N_21314,N_20433);
xor U23389 (N_23389,N_22289,N_21479);
xnor U23390 (N_23390,N_21672,N_22446);
or U23391 (N_23391,N_20385,N_21469);
nand U23392 (N_23392,N_21527,N_21136);
xor U23393 (N_23393,N_20089,N_21935);
and U23394 (N_23394,N_21089,N_21386);
xor U23395 (N_23395,N_22270,N_21923);
nand U23396 (N_23396,N_20881,N_22150);
nand U23397 (N_23397,N_21525,N_20698);
xor U23398 (N_23398,N_20155,N_21744);
nand U23399 (N_23399,N_20693,N_21843);
nand U23400 (N_23400,N_20287,N_22297);
xnor U23401 (N_23401,N_20082,N_22255);
and U23402 (N_23402,N_20620,N_21257);
and U23403 (N_23403,N_20545,N_21982);
nand U23404 (N_23404,N_21979,N_21883);
and U23405 (N_23405,N_20497,N_22475);
or U23406 (N_23406,N_20530,N_20762);
or U23407 (N_23407,N_22148,N_21937);
and U23408 (N_23408,N_20910,N_22410);
xnor U23409 (N_23409,N_20860,N_21520);
nor U23410 (N_23410,N_22100,N_20534);
xnor U23411 (N_23411,N_22236,N_22188);
nand U23412 (N_23412,N_21370,N_22495);
or U23413 (N_23413,N_20403,N_22467);
nand U23414 (N_23414,N_20135,N_21026);
or U23415 (N_23415,N_20744,N_22268);
nand U23416 (N_23416,N_20855,N_21753);
nor U23417 (N_23417,N_22019,N_20364);
nor U23418 (N_23418,N_20768,N_21635);
nand U23419 (N_23419,N_20748,N_20030);
nand U23420 (N_23420,N_21964,N_21335);
nand U23421 (N_23421,N_20936,N_21584);
nor U23422 (N_23422,N_21499,N_21096);
and U23423 (N_23423,N_20353,N_22473);
and U23424 (N_23424,N_20857,N_20711);
xnor U23425 (N_23425,N_21732,N_20819);
nand U23426 (N_23426,N_20133,N_21184);
and U23427 (N_23427,N_21452,N_21002);
xor U23428 (N_23428,N_21067,N_21119);
nand U23429 (N_23429,N_22380,N_20636);
xnor U23430 (N_23430,N_21703,N_20090);
and U23431 (N_23431,N_21641,N_20864);
xnor U23432 (N_23432,N_22052,N_21644);
or U23433 (N_23433,N_21931,N_20310);
nor U23434 (N_23434,N_21327,N_21247);
xor U23435 (N_23435,N_21920,N_20262);
and U23436 (N_23436,N_22251,N_21120);
or U23437 (N_23437,N_20038,N_20103);
nor U23438 (N_23438,N_20843,N_20174);
and U23439 (N_23439,N_21305,N_21156);
nand U23440 (N_23440,N_21367,N_22028);
nor U23441 (N_23441,N_22445,N_21389);
nor U23442 (N_23442,N_21629,N_21518);
and U23443 (N_23443,N_21413,N_21733);
and U23444 (N_23444,N_22078,N_22210);
xnor U23445 (N_23445,N_21724,N_20306);
xnor U23446 (N_23446,N_21533,N_20615);
and U23447 (N_23447,N_21776,N_22341);
xor U23448 (N_23448,N_22447,N_20847);
nand U23449 (N_23449,N_22392,N_21586);
or U23450 (N_23450,N_20350,N_21701);
and U23451 (N_23451,N_20523,N_22295);
xor U23452 (N_23452,N_21977,N_20605);
and U23453 (N_23453,N_21625,N_20925);
and U23454 (N_23454,N_20874,N_20632);
and U23455 (N_23455,N_20000,N_22173);
nor U23456 (N_23456,N_21242,N_20130);
nand U23457 (N_23457,N_20299,N_22151);
nor U23458 (N_23458,N_22412,N_20442);
nand U23459 (N_23459,N_22145,N_22274);
or U23460 (N_23460,N_21108,N_20552);
nor U23461 (N_23461,N_20689,N_20165);
xor U23462 (N_23462,N_20307,N_20388);
nor U23463 (N_23463,N_22403,N_20447);
nand U23464 (N_23464,N_21381,N_22114);
nand U23465 (N_23465,N_21618,N_20291);
xnor U23466 (N_23466,N_21870,N_20832);
nand U23467 (N_23467,N_20745,N_22233);
or U23468 (N_23468,N_20715,N_21890);
nand U23469 (N_23469,N_22337,N_22200);
nor U23470 (N_23470,N_21435,N_21345);
nand U23471 (N_23471,N_22486,N_22448);
or U23472 (N_23472,N_20112,N_21532);
and U23473 (N_23473,N_20221,N_21646);
or U23474 (N_23474,N_20439,N_20981);
xor U23475 (N_23475,N_20330,N_21555);
xor U23476 (N_23476,N_20704,N_21480);
and U23477 (N_23477,N_20654,N_20831);
and U23478 (N_23478,N_21167,N_20450);
nor U23479 (N_23479,N_22451,N_21992);
and U23480 (N_23480,N_20999,N_22361);
nor U23481 (N_23481,N_21238,N_20793);
or U23482 (N_23482,N_21593,N_21559);
nor U23483 (N_23483,N_22428,N_21534);
and U23484 (N_23484,N_21198,N_20782);
nand U23485 (N_23485,N_22065,N_20086);
and U23486 (N_23486,N_21408,N_21823);
xor U23487 (N_23487,N_21891,N_20313);
nand U23488 (N_23488,N_20928,N_21548);
xor U23489 (N_23489,N_22131,N_20529);
nor U23490 (N_23490,N_22348,N_21748);
xor U23491 (N_23491,N_21461,N_21551);
or U23492 (N_23492,N_20648,N_21201);
nor U23493 (N_23493,N_20467,N_22179);
xnor U23494 (N_23494,N_22398,N_21403);
xnor U23495 (N_23495,N_22107,N_21560);
nor U23496 (N_23496,N_20579,N_20528);
xor U23497 (N_23497,N_22171,N_20550);
xnor U23498 (N_23498,N_21038,N_21164);
nor U23499 (N_23499,N_20128,N_22012);
nor U23500 (N_23500,N_22189,N_21359);
nor U23501 (N_23501,N_20649,N_22464);
and U23502 (N_23502,N_21319,N_20377);
xor U23503 (N_23503,N_21239,N_22198);
nand U23504 (N_23504,N_22458,N_21737);
or U23505 (N_23505,N_20677,N_22390);
xnor U23506 (N_23506,N_20473,N_20830);
and U23507 (N_23507,N_22250,N_21576);
and U23508 (N_23508,N_21395,N_21614);
nor U23509 (N_23509,N_21639,N_20486);
nor U23510 (N_23510,N_20717,N_20975);
xor U23511 (N_23511,N_20525,N_20341);
xnor U23512 (N_23512,N_21207,N_21100);
nor U23513 (N_23513,N_21985,N_21505);
or U23514 (N_23514,N_21649,N_20444);
xor U23515 (N_23515,N_21029,N_20159);
nor U23516 (N_23516,N_20719,N_20012);
nand U23517 (N_23517,N_20136,N_20888);
nand U23518 (N_23518,N_21465,N_21685);
nand U23519 (N_23519,N_20416,N_22070);
nor U23520 (N_23520,N_21524,N_21206);
xnor U23521 (N_23521,N_21567,N_20323);
xor U23522 (N_23522,N_20184,N_20206);
or U23523 (N_23523,N_21055,N_20463);
and U23524 (N_23524,N_21579,N_22378);
xor U23525 (N_23525,N_22300,N_20344);
nor U23526 (N_23526,N_22172,N_21847);
nand U23527 (N_23527,N_20108,N_21623);
xnor U23528 (N_23528,N_21250,N_21404);
and U23529 (N_23529,N_21578,N_21783);
or U23530 (N_23530,N_21731,N_20734);
nor U23531 (N_23531,N_22079,N_20321);
nand U23532 (N_23532,N_21965,N_21583);
nor U23533 (N_23533,N_21349,N_21475);
nor U23534 (N_23534,N_20201,N_21877);
nor U23535 (N_23535,N_21828,N_21095);
nand U23536 (N_23536,N_21352,N_20807);
nor U23537 (N_23537,N_20014,N_22313);
nand U23538 (N_23538,N_21600,N_21442);
and U23539 (N_23539,N_20879,N_21341);
and U23540 (N_23540,N_22436,N_20238);
or U23541 (N_23541,N_20334,N_21430);
xor U23542 (N_23542,N_22069,N_20993);
or U23543 (N_23543,N_20148,N_21421);
nand U23544 (N_23544,N_21972,N_20013);
or U23545 (N_23545,N_21627,N_20192);
nand U23546 (N_23546,N_21312,N_21387);
and U23547 (N_23547,N_22040,N_20788);
nand U23548 (N_23548,N_20547,N_20124);
nor U23549 (N_23549,N_20193,N_20404);
nand U23550 (N_23550,N_21740,N_21848);
xnor U23551 (N_23551,N_21841,N_22053);
xor U23552 (N_23552,N_21005,N_20118);
xor U23553 (N_23553,N_22395,N_21066);
or U23554 (N_23554,N_21419,N_22407);
nand U23555 (N_23555,N_22221,N_20779);
nor U23556 (N_23556,N_20304,N_20891);
or U23557 (N_23557,N_21264,N_21143);
and U23558 (N_23558,N_21874,N_20460);
nor U23559 (N_23559,N_22206,N_20040);
nor U23560 (N_23560,N_21166,N_20817);
nor U23561 (N_23561,N_21673,N_22479);
nand U23562 (N_23562,N_20877,N_20204);
and U23563 (N_23563,N_22235,N_22370);
xnor U23564 (N_23564,N_22419,N_22373);
and U23565 (N_23565,N_20209,N_21064);
or U23566 (N_23566,N_20722,N_20047);
or U23567 (N_23567,N_20806,N_20010);
nor U23568 (N_23568,N_21834,N_22342);
or U23569 (N_23569,N_20080,N_21340);
nand U23570 (N_23570,N_21544,N_21439);
nand U23571 (N_23571,N_21489,N_22042);
nand U23572 (N_23572,N_20236,N_20160);
and U23573 (N_23573,N_21306,N_20445);
nand U23574 (N_23574,N_21872,N_21721);
or U23575 (N_23575,N_20458,N_21223);
or U23576 (N_23576,N_21459,N_20661);
nand U23577 (N_23577,N_20219,N_20789);
nand U23578 (N_23578,N_20746,N_21414);
nor U23579 (N_23579,N_20604,N_21815);
nor U23580 (N_23580,N_22225,N_21420);
and U23581 (N_23581,N_20303,N_21723);
and U23582 (N_23582,N_22325,N_22276);
nor U23583 (N_23583,N_21846,N_21134);
xnor U23584 (N_23584,N_22104,N_20042);
xor U23585 (N_23585,N_21291,N_22442);
and U23586 (N_23586,N_21506,N_22355);
nand U23587 (N_23587,N_22443,N_21281);
xor U23588 (N_23588,N_21073,N_21061);
or U23589 (N_23589,N_20297,N_20929);
nand U23590 (N_23590,N_21261,N_21684);
and U23591 (N_23591,N_20532,N_20823);
nor U23592 (N_23592,N_22493,N_21814);
and U23593 (N_23593,N_20655,N_21713);
nand U23594 (N_23594,N_21956,N_20264);
nand U23595 (N_23595,N_22178,N_20548);
and U23596 (N_23596,N_20683,N_20562);
xnor U23597 (N_23597,N_21170,N_21292);
nor U23598 (N_23598,N_20260,N_22426);
nor U23599 (N_23599,N_22048,N_22081);
or U23600 (N_23600,N_20846,N_20712);
xor U23601 (N_23601,N_22230,N_21531);
nor U23602 (N_23602,N_21182,N_20799);
nor U23603 (N_23603,N_21795,N_20521);
and U23604 (N_23604,N_22193,N_22391);
and U23605 (N_23605,N_20071,N_21529);
and U23606 (N_23606,N_21375,N_22468);
nor U23607 (N_23607,N_20992,N_22029);
nor U23608 (N_23608,N_21726,N_21225);
xnor U23609 (N_23609,N_20868,N_20901);
nand U23610 (N_23610,N_22026,N_20208);
nand U23611 (N_23611,N_21399,N_20270);
and U23612 (N_23612,N_21172,N_20524);
nand U23613 (N_23613,N_21844,N_22477);
or U23614 (N_23614,N_21168,N_21839);
nand U23615 (N_23615,N_20106,N_21457);
and U23616 (N_23616,N_20775,N_20492);
xnor U23617 (N_23617,N_21003,N_22376);
nor U23618 (N_23618,N_20885,N_20280);
and U23619 (N_23619,N_22209,N_21298);
and U23620 (N_23620,N_20484,N_20115);
nor U23621 (N_23621,N_21398,N_20498);
nand U23622 (N_23622,N_21202,N_21138);
nor U23623 (N_23623,N_20205,N_20340);
nand U23624 (N_23624,N_21324,N_22170);
xnor U23625 (N_23625,N_21132,N_21711);
xor U23626 (N_23626,N_21766,N_22310);
or U23627 (N_23627,N_20092,N_21380);
or U23628 (N_23628,N_20594,N_21455);
or U23629 (N_23629,N_22478,N_22058);
or U23630 (N_23630,N_20382,N_21374);
nor U23631 (N_23631,N_20911,N_20191);
xnor U23632 (N_23632,N_22396,N_21704);
xor U23633 (N_23633,N_21216,N_22330);
nand U23634 (N_23634,N_21492,N_21412);
nand U23635 (N_23635,N_21805,N_20189);
or U23636 (N_23636,N_20876,N_22197);
nor U23637 (N_23637,N_21268,N_22263);
and U23638 (N_23638,N_20707,N_22280);
xnor U23639 (N_23639,N_20838,N_21014);
and U23640 (N_23640,N_21606,N_22044);
xor U23641 (N_23641,N_21227,N_22261);
or U23642 (N_23642,N_20158,N_20702);
nand U23643 (N_23643,N_21549,N_20672);
and U23644 (N_23644,N_20668,N_21059);
and U23645 (N_23645,N_21620,N_22463);
and U23646 (N_23646,N_20790,N_21879);
and U23647 (N_23647,N_20791,N_20554);
or U23648 (N_23648,N_20431,N_21611);
nor U23649 (N_23649,N_21621,N_21714);
and U23650 (N_23650,N_20805,N_20889);
xor U23651 (N_23651,N_20211,N_21700);
nand U23652 (N_23652,N_20232,N_21440);
nor U23653 (N_23653,N_21679,N_21272);
nor U23654 (N_23654,N_21438,N_21427);
nand U23655 (N_23655,N_21233,N_22112);
or U23656 (N_23656,N_21310,N_21178);
or U23657 (N_23657,N_20741,N_20380);
and U23658 (N_23658,N_21013,N_21484);
and U23659 (N_23659,N_22353,N_21950);
and U23660 (N_23660,N_22157,N_20630);
xnor U23661 (N_23661,N_22202,N_21771);
and U23662 (N_23662,N_20961,N_20066);
xnor U23663 (N_23663,N_21613,N_20810);
nor U23664 (N_23664,N_22096,N_21930);
or U23665 (N_23665,N_22480,N_20100);
nor U23666 (N_23666,N_20349,N_20028);
nor U23667 (N_23667,N_22186,N_20446);
nor U23668 (N_23668,N_21084,N_21130);
and U23669 (N_23669,N_20144,N_20454);
xor U23670 (N_23670,N_21939,N_21553);
nor U23671 (N_23671,N_21645,N_21353);
xor U23672 (N_23672,N_21346,N_21676);
xnor U23673 (N_23673,N_20202,N_21632);
nor U23674 (N_23674,N_20772,N_21049);
nor U23675 (N_23675,N_20070,N_21596);
or U23676 (N_23676,N_21708,N_20732);
xor U23677 (N_23677,N_22301,N_22038);
nor U23678 (N_23678,N_21302,N_20967);
or U23679 (N_23679,N_21483,N_20795);
nor U23680 (N_23680,N_20488,N_20697);
and U23681 (N_23681,N_20415,N_20263);
xor U23682 (N_23682,N_22406,N_22409);
and U23683 (N_23683,N_21813,N_22105);
nor U23684 (N_23684,N_20465,N_20616);
xnor U23685 (N_23685,N_21023,N_20764);
xnor U23686 (N_23686,N_20339,N_21539);
nor U23687 (N_23687,N_22217,N_20333);
nand U23688 (N_23688,N_21124,N_21187);
and U23689 (N_23689,N_21862,N_21994);
nor U23690 (N_23690,N_20639,N_20338);
or U23691 (N_23691,N_20968,N_20861);
and U23692 (N_23692,N_21117,N_22293);
and U23693 (N_23693,N_20006,N_21456);
and U23694 (N_23694,N_21652,N_20305);
nor U23695 (N_23695,N_20391,N_21990);
nor U23696 (N_23696,N_20908,N_22124);
nand U23697 (N_23697,N_20408,N_20591);
xor U23698 (N_23698,N_22227,N_21545);
nand U23699 (N_23699,N_20769,N_20411);
nand U23700 (N_23700,N_20834,N_20396);
xnor U23701 (N_23701,N_20002,N_21022);
nand U23702 (N_23702,N_20537,N_20641);
nand U23703 (N_23703,N_20749,N_21565);
nor U23704 (N_23704,N_21643,N_20067);
nand U23705 (N_23705,N_22133,N_22431);
or U23706 (N_23706,N_20973,N_20921);
nand U23707 (N_23707,N_21577,N_21971);
or U23708 (N_23708,N_21195,N_20278);
or U23709 (N_23709,N_21793,N_21829);
nand U23710 (N_23710,N_22122,N_21571);
xor U23711 (N_23711,N_20032,N_21510);
or U23712 (N_23712,N_20044,N_21174);
nor U23713 (N_23713,N_20766,N_20257);
nor U23714 (N_23714,N_20951,N_21590);
and U23715 (N_23715,N_20230,N_20457);
and U23716 (N_23716,N_22218,N_21637);
nand U23717 (N_23717,N_20357,N_20237);
xor U23718 (N_23718,N_21597,N_20336);
or U23719 (N_23719,N_21350,N_22365);
and U23720 (N_23720,N_21116,N_20583);
nor U23721 (N_23721,N_22344,N_21424);
xor U23722 (N_23722,N_20798,N_20727);
or U23723 (N_23723,N_20618,N_22130);
nand U23724 (N_23724,N_20996,N_21696);
xor U23725 (N_23725,N_21036,N_21508);
nand U23726 (N_23726,N_21249,N_20900);
or U23727 (N_23727,N_20797,N_21790);
xnor U23728 (N_23728,N_20538,N_20055);
or U23729 (N_23729,N_22015,N_22471);
nand U23730 (N_23730,N_20249,N_20478);
xnor U23731 (N_23731,N_20517,N_22011);
or U23732 (N_23732,N_22004,N_20186);
xor U23733 (N_23733,N_22224,N_20542);
nor U23734 (N_23734,N_20027,N_20327);
nor U23735 (N_23735,N_21391,N_22460);
or U23736 (N_23736,N_22023,N_21486);
and U23737 (N_23737,N_20393,N_20714);
and U23738 (N_23738,N_21978,N_20104);
nand U23739 (N_23739,N_22177,N_20647);
or U23740 (N_23740,N_22135,N_20777);
xor U23741 (N_23741,N_20143,N_22367);
or U23742 (N_23742,N_22110,N_22292);
nand U23743 (N_23743,N_20959,N_20747);
and U23744 (N_23744,N_21574,N_21999);
or U23745 (N_23745,N_20139,N_20990);
nand U23746 (N_23746,N_21190,N_20644);
xor U23747 (N_23747,N_20483,N_21986);
nor U23748 (N_23748,N_20546,N_21361);
xor U23749 (N_23749,N_22389,N_20176);
nor U23750 (N_23750,N_21912,N_21444);
nand U23751 (N_23751,N_21362,N_21887);
or U23752 (N_23752,N_21097,N_22437);
nand U23753 (N_23753,N_21374,N_20944);
xor U23754 (N_23754,N_20294,N_22381);
or U23755 (N_23755,N_20347,N_22249);
nor U23756 (N_23756,N_21757,N_21586);
nor U23757 (N_23757,N_22308,N_21276);
nor U23758 (N_23758,N_20405,N_20410);
and U23759 (N_23759,N_20057,N_21249);
or U23760 (N_23760,N_22298,N_21215);
or U23761 (N_23761,N_21723,N_21807);
nor U23762 (N_23762,N_21318,N_20659);
nand U23763 (N_23763,N_20742,N_21478);
or U23764 (N_23764,N_21085,N_21184);
nor U23765 (N_23765,N_21605,N_21868);
or U23766 (N_23766,N_20333,N_22413);
xnor U23767 (N_23767,N_22184,N_20686);
nand U23768 (N_23768,N_21091,N_20167);
nand U23769 (N_23769,N_20579,N_21552);
nor U23770 (N_23770,N_20509,N_20170);
and U23771 (N_23771,N_20484,N_20352);
nor U23772 (N_23772,N_22248,N_21144);
and U23773 (N_23773,N_21356,N_20797);
xor U23774 (N_23774,N_21420,N_21814);
or U23775 (N_23775,N_20864,N_20361);
or U23776 (N_23776,N_20227,N_21249);
xor U23777 (N_23777,N_21675,N_21008);
and U23778 (N_23778,N_21554,N_20752);
xor U23779 (N_23779,N_20912,N_20762);
nor U23780 (N_23780,N_21388,N_21387);
and U23781 (N_23781,N_22298,N_22172);
or U23782 (N_23782,N_21937,N_20021);
nor U23783 (N_23783,N_21635,N_20636);
and U23784 (N_23784,N_21946,N_20274);
or U23785 (N_23785,N_21016,N_22479);
and U23786 (N_23786,N_22472,N_20220);
xnor U23787 (N_23787,N_21291,N_20981);
xnor U23788 (N_23788,N_22086,N_20797);
nor U23789 (N_23789,N_22398,N_20662);
xor U23790 (N_23790,N_21051,N_20051);
xnor U23791 (N_23791,N_20338,N_21753);
xnor U23792 (N_23792,N_20630,N_20137);
and U23793 (N_23793,N_21101,N_20657);
or U23794 (N_23794,N_22449,N_20342);
xnor U23795 (N_23795,N_20139,N_21597);
nor U23796 (N_23796,N_21646,N_22026);
and U23797 (N_23797,N_20440,N_20002);
or U23798 (N_23798,N_21008,N_20239);
nor U23799 (N_23799,N_22272,N_21882);
and U23800 (N_23800,N_20715,N_21782);
nand U23801 (N_23801,N_21919,N_21616);
or U23802 (N_23802,N_22136,N_21951);
or U23803 (N_23803,N_21993,N_20804);
xor U23804 (N_23804,N_20636,N_21159);
and U23805 (N_23805,N_20207,N_21485);
nor U23806 (N_23806,N_20316,N_20158);
or U23807 (N_23807,N_21594,N_20364);
and U23808 (N_23808,N_20453,N_20196);
and U23809 (N_23809,N_21026,N_21234);
xnor U23810 (N_23810,N_22323,N_22076);
xnor U23811 (N_23811,N_22428,N_22231);
nand U23812 (N_23812,N_22336,N_22346);
xor U23813 (N_23813,N_20063,N_22059);
xor U23814 (N_23814,N_20033,N_20011);
xnor U23815 (N_23815,N_21949,N_22184);
xor U23816 (N_23816,N_20335,N_20149);
or U23817 (N_23817,N_21471,N_20694);
nor U23818 (N_23818,N_21287,N_22453);
or U23819 (N_23819,N_21656,N_22007);
nand U23820 (N_23820,N_21058,N_20521);
nand U23821 (N_23821,N_20382,N_20320);
and U23822 (N_23822,N_21520,N_21461);
and U23823 (N_23823,N_20791,N_21106);
xnor U23824 (N_23824,N_21864,N_20677);
or U23825 (N_23825,N_20357,N_21668);
nand U23826 (N_23826,N_21395,N_20399);
xnor U23827 (N_23827,N_21533,N_21977);
xnor U23828 (N_23828,N_22403,N_21583);
nand U23829 (N_23829,N_20244,N_21128);
and U23830 (N_23830,N_22316,N_20319);
nor U23831 (N_23831,N_20552,N_22271);
xnor U23832 (N_23832,N_21429,N_22057);
and U23833 (N_23833,N_21186,N_21264);
or U23834 (N_23834,N_20569,N_20653);
or U23835 (N_23835,N_20299,N_21047);
and U23836 (N_23836,N_21806,N_22088);
xnor U23837 (N_23837,N_20614,N_22135);
or U23838 (N_23838,N_20423,N_21905);
or U23839 (N_23839,N_21061,N_21838);
nor U23840 (N_23840,N_22093,N_22023);
and U23841 (N_23841,N_20409,N_20175);
or U23842 (N_23842,N_20192,N_20626);
and U23843 (N_23843,N_21848,N_22170);
xor U23844 (N_23844,N_21925,N_21553);
xnor U23845 (N_23845,N_21097,N_20004);
nor U23846 (N_23846,N_20434,N_22252);
nand U23847 (N_23847,N_20260,N_20283);
and U23848 (N_23848,N_21169,N_22427);
xor U23849 (N_23849,N_21248,N_20490);
or U23850 (N_23850,N_21574,N_21095);
nor U23851 (N_23851,N_22329,N_21499);
nand U23852 (N_23852,N_20806,N_22290);
and U23853 (N_23853,N_21755,N_22255);
nor U23854 (N_23854,N_22445,N_21062);
xnor U23855 (N_23855,N_20101,N_21887);
nand U23856 (N_23856,N_21816,N_21623);
or U23857 (N_23857,N_20733,N_20126);
nor U23858 (N_23858,N_20781,N_21393);
xnor U23859 (N_23859,N_20529,N_22282);
nor U23860 (N_23860,N_21695,N_20239);
or U23861 (N_23861,N_21890,N_21680);
or U23862 (N_23862,N_21738,N_20922);
nand U23863 (N_23863,N_22362,N_21591);
nand U23864 (N_23864,N_20996,N_21444);
nand U23865 (N_23865,N_22430,N_21600);
nand U23866 (N_23866,N_22442,N_20652);
and U23867 (N_23867,N_21064,N_21531);
or U23868 (N_23868,N_21519,N_20718);
and U23869 (N_23869,N_22336,N_21711);
and U23870 (N_23870,N_21067,N_22045);
nor U23871 (N_23871,N_22184,N_22388);
and U23872 (N_23872,N_21656,N_20770);
and U23873 (N_23873,N_20486,N_20170);
xnor U23874 (N_23874,N_20860,N_20383);
or U23875 (N_23875,N_22137,N_20520);
nor U23876 (N_23876,N_22315,N_22068);
and U23877 (N_23877,N_20304,N_21449);
or U23878 (N_23878,N_20250,N_21318);
and U23879 (N_23879,N_20756,N_22279);
nor U23880 (N_23880,N_20877,N_20061);
nand U23881 (N_23881,N_20394,N_20283);
and U23882 (N_23882,N_20304,N_21640);
nand U23883 (N_23883,N_22209,N_22293);
nor U23884 (N_23884,N_22338,N_21120);
and U23885 (N_23885,N_21165,N_21629);
and U23886 (N_23886,N_22007,N_20430);
nand U23887 (N_23887,N_21912,N_21865);
xnor U23888 (N_23888,N_21538,N_21785);
nand U23889 (N_23889,N_22463,N_20962);
xnor U23890 (N_23890,N_20115,N_20980);
or U23891 (N_23891,N_21120,N_22367);
nand U23892 (N_23892,N_21090,N_20844);
nand U23893 (N_23893,N_21907,N_20689);
xnor U23894 (N_23894,N_21454,N_21610);
or U23895 (N_23895,N_20653,N_21049);
or U23896 (N_23896,N_21467,N_22227);
or U23897 (N_23897,N_22427,N_21401);
xor U23898 (N_23898,N_22210,N_20489);
nand U23899 (N_23899,N_22466,N_21119);
or U23900 (N_23900,N_22274,N_20001);
or U23901 (N_23901,N_22258,N_21045);
nor U23902 (N_23902,N_21764,N_22095);
nand U23903 (N_23903,N_21585,N_22290);
nand U23904 (N_23904,N_20396,N_22149);
nor U23905 (N_23905,N_20009,N_20169);
nand U23906 (N_23906,N_22130,N_20931);
nand U23907 (N_23907,N_21992,N_20880);
nor U23908 (N_23908,N_22479,N_21024);
nand U23909 (N_23909,N_22233,N_20412);
nand U23910 (N_23910,N_20059,N_20765);
or U23911 (N_23911,N_21778,N_21096);
xnor U23912 (N_23912,N_21270,N_20521);
nor U23913 (N_23913,N_20758,N_20383);
and U23914 (N_23914,N_21673,N_21526);
and U23915 (N_23915,N_20578,N_20922);
and U23916 (N_23916,N_20136,N_21662);
xnor U23917 (N_23917,N_20630,N_22067);
and U23918 (N_23918,N_20401,N_20559);
or U23919 (N_23919,N_22426,N_21753);
nor U23920 (N_23920,N_22438,N_21921);
and U23921 (N_23921,N_22369,N_21210);
xnor U23922 (N_23922,N_20153,N_20867);
nand U23923 (N_23923,N_22138,N_20401);
nand U23924 (N_23924,N_21004,N_20558);
nor U23925 (N_23925,N_20974,N_20100);
nor U23926 (N_23926,N_20525,N_20238);
xnor U23927 (N_23927,N_21755,N_20691);
or U23928 (N_23928,N_20248,N_20116);
and U23929 (N_23929,N_21905,N_20515);
and U23930 (N_23930,N_21055,N_21308);
and U23931 (N_23931,N_21948,N_20981);
or U23932 (N_23932,N_20657,N_22179);
and U23933 (N_23933,N_20181,N_21313);
nand U23934 (N_23934,N_20479,N_21492);
and U23935 (N_23935,N_21595,N_20199);
or U23936 (N_23936,N_21910,N_21260);
nand U23937 (N_23937,N_21106,N_20783);
and U23938 (N_23938,N_21369,N_20466);
nor U23939 (N_23939,N_20191,N_22458);
xor U23940 (N_23940,N_20783,N_20093);
and U23941 (N_23941,N_20095,N_22064);
and U23942 (N_23942,N_20971,N_20508);
xnor U23943 (N_23943,N_21206,N_21595);
or U23944 (N_23944,N_21272,N_20212);
nor U23945 (N_23945,N_22008,N_20661);
xor U23946 (N_23946,N_22178,N_22081);
and U23947 (N_23947,N_20686,N_20425);
or U23948 (N_23948,N_22149,N_20229);
or U23949 (N_23949,N_20643,N_20815);
and U23950 (N_23950,N_20205,N_21820);
or U23951 (N_23951,N_20157,N_21346);
nor U23952 (N_23952,N_22284,N_21181);
or U23953 (N_23953,N_20612,N_21004);
nand U23954 (N_23954,N_21621,N_21826);
and U23955 (N_23955,N_20397,N_21343);
or U23956 (N_23956,N_21174,N_22426);
nand U23957 (N_23957,N_20805,N_22315);
nand U23958 (N_23958,N_21215,N_20718);
nor U23959 (N_23959,N_21531,N_20321);
nor U23960 (N_23960,N_21144,N_20070);
xnor U23961 (N_23961,N_20248,N_22278);
nor U23962 (N_23962,N_20135,N_22031);
nor U23963 (N_23963,N_22464,N_21520);
nor U23964 (N_23964,N_21083,N_21309);
xor U23965 (N_23965,N_21230,N_22327);
and U23966 (N_23966,N_20862,N_22284);
and U23967 (N_23967,N_20322,N_21957);
nand U23968 (N_23968,N_20221,N_21567);
and U23969 (N_23969,N_20032,N_21941);
or U23970 (N_23970,N_21701,N_20081);
nor U23971 (N_23971,N_21009,N_21670);
nor U23972 (N_23972,N_21872,N_21233);
or U23973 (N_23973,N_21574,N_21018);
xor U23974 (N_23974,N_22324,N_20867);
and U23975 (N_23975,N_21038,N_21386);
or U23976 (N_23976,N_21813,N_21774);
or U23977 (N_23977,N_22193,N_20265);
nand U23978 (N_23978,N_20405,N_20500);
nor U23979 (N_23979,N_21008,N_20110);
nand U23980 (N_23980,N_20111,N_21241);
and U23981 (N_23981,N_20493,N_21109);
or U23982 (N_23982,N_20940,N_21649);
or U23983 (N_23983,N_21892,N_20145);
nor U23984 (N_23984,N_21145,N_22077);
nand U23985 (N_23985,N_21637,N_20237);
nor U23986 (N_23986,N_21386,N_22480);
nor U23987 (N_23987,N_20962,N_21008);
or U23988 (N_23988,N_21112,N_20167);
nand U23989 (N_23989,N_20135,N_22372);
or U23990 (N_23990,N_22285,N_22108);
and U23991 (N_23991,N_21169,N_21425);
xor U23992 (N_23992,N_21512,N_20734);
or U23993 (N_23993,N_21485,N_21659);
or U23994 (N_23994,N_21175,N_22323);
or U23995 (N_23995,N_21253,N_21714);
nand U23996 (N_23996,N_20897,N_22020);
nor U23997 (N_23997,N_22344,N_20762);
or U23998 (N_23998,N_21672,N_21612);
xor U23999 (N_23999,N_20289,N_20838);
or U24000 (N_24000,N_21738,N_22409);
nand U24001 (N_24001,N_21920,N_21421);
nand U24002 (N_24002,N_20132,N_22341);
or U24003 (N_24003,N_20954,N_21361);
and U24004 (N_24004,N_20037,N_21568);
and U24005 (N_24005,N_22167,N_22335);
or U24006 (N_24006,N_20760,N_21087);
or U24007 (N_24007,N_20891,N_21455);
nand U24008 (N_24008,N_20349,N_21659);
and U24009 (N_24009,N_20500,N_20711);
nand U24010 (N_24010,N_22443,N_22078);
or U24011 (N_24011,N_20424,N_22227);
or U24012 (N_24012,N_21605,N_20677);
and U24013 (N_24013,N_22294,N_21906);
and U24014 (N_24014,N_21075,N_21548);
or U24015 (N_24015,N_20071,N_21649);
xor U24016 (N_24016,N_20577,N_21620);
nand U24017 (N_24017,N_22497,N_20141);
or U24018 (N_24018,N_21784,N_20017);
or U24019 (N_24019,N_20217,N_21733);
nor U24020 (N_24020,N_21219,N_22463);
and U24021 (N_24021,N_21200,N_22197);
nor U24022 (N_24022,N_21422,N_22170);
nor U24023 (N_24023,N_20264,N_21544);
nand U24024 (N_24024,N_20130,N_20942);
nor U24025 (N_24025,N_21536,N_21503);
and U24026 (N_24026,N_21415,N_22352);
nand U24027 (N_24027,N_20771,N_22342);
and U24028 (N_24028,N_20787,N_21297);
nand U24029 (N_24029,N_20579,N_20017);
and U24030 (N_24030,N_20731,N_22297);
and U24031 (N_24031,N_21813,N_21976);
nand U24032 (N_24032,N_20493,N_20741);
and U24033 (N_24033,N_20834,N_22342);
xor U24034 (N_24034,N_21800,N_21355);
xnor U24035 (N_24035,N_20387,N_21440);
and U24036 (N_24036,N_21611,N_21078);
and U24037 (N_24037,N_22431,N_22274);
nor U24038 (N_24038,N_21043,N_20625);
xor U24039 (N_24039,N_21732,N_22193);
and U24040 (N_24040,N_22234,N_22299);
xnor U24041 (N_24041,N_20937,N_21032);
or U24042 (N_24042,N_21703,N_21166);
xor U24043 (N_24043,N_20838,N_21895);
or U24044 (N_24044,N_22252,N_20672);
or U24045 (N_24045,N_21090,N_20656);
nand U24046 (N_24046,N_21044,N_21707);
nand U24047 (N_24047,N_21511,N_20336);
nor U24048 (N_24048,N_20648,N_21227);
xnor U24049 (N_24049,N_20691,N_22345);
nand U24050 (N_24050,N_20076,N_21569);
nor U24051 (N_24051,N_21946,N_20630);
or U24052 (N_24052,N_21427,N_21509);
and U24053 (N_24053,N_21032,N_22130);
nand U24054 (N_24054,N_21933,N_22175);
xnor U24055 (N_24055,N_21964,N_20567);
xor U24056 (N_24056,N_21971,N_21966);
nand U24057 (N_24057,N_20019,N_21649);
nand U24058 (N_24058,N_20720,N_21721);
xor U24059 (N_24059,N_21182,N_22400);
and U24060 (N_24060,N_20441,N_21410);
nor U24061 (N_24061,N_21773,N_21276);
and U24062 (N_24062,N_20133,N_21087);
or U24063 (N_24063,N_20711,N_20607);
xor U24064 (N_24064,N_20503,N_21982);
and U24065 (N_24065,N_21674,N_20135);
or U24066 (N_24066,N_20705,N_22020);
nand U24067 (N_24067,N_21671,N_20431);
and U24068 (N_24068,N_21104,N_20604);
nor U24069 (N_24069,N_21812,N_20303);
or U24070 (N_24070,N_21620,N_22391);
nand U24071 (N_24071,N_21357,N_22132);
nor U24072 (N_24072,N_21843,N_21821);
nor U24073 (N_24073,N_22480,N_20231);
nor U24074 (N_24074,N_20962,N_22159);
and U24075 (N_24075,N_22020,N_20606);
xnor U24076 (N_24076,N_20907,N_21982);
and U24077 (N_24077,N_20453,N_21573);
xor U24078 (N_24078,N_20801,N_22018);
xnor U24079 (N_24079,N_22284,N_21069);
xnor U24080 (N_24080,N_21775,N_21866);
and U24081 (N_24081,N_20320,N_21965);
xor U24082 (N_24082,N_22297,N_21437);
or U24083 (N_24083,N_20868,N_21148);
and U24084 (N_24084,N_21708,N_21950);
or U24085 (N_24085,N_20155,N_21665);
or U24086 (N_24086,N_21879,N_20416);
nand U24087 (N_24087,N_20959,N_21500);
xnor U24088 (N_24088,N_22207,N_22131);
nand U24089 (N_24089,N_21066,N_21968);
xor U24090 (N_24090,N_21983,N_22310);
xnor U24091 (N_24091,N_21307,N_21723);
nor U24092 (N_24092,N_20507,N_20280);
xor U24093 (N_24093,N_21648,N_22449);
nand U24094 (N_24094,N_21155,N_22272);
or U24095 (N_24095,N_20569,N_20585);
xnor U24096 (N_24096,N_21785,N_20562);
and U24097 (N_24097,N_21237,N_20890);
nand U24098 (N_24098,N_20250,N_20141);
nand U24099 (N_24099,N_22406,N_21653);
xor U24100 (N_24100,N_20289,N_20807);
xor U24101 (N_24101,N_22337,N_21076);
nor U24102 (N_24102,N_20535,N_20318);
nor U24103 (N_24103,N_21396,N_22355);
or U24104 (N_24104,N_21387,N_21276);
nand U24105 (N_24105,N_20154,N_20148);
xnor U24106 (N_24106,N_20318,N_20691);
or U24107 (N_24107,N_20414,N_21383);
nor U24108 (N_24108,N_21143,N_22491);
and U24109 (N_24109,N_20869,N_20617);
or U24110 (N_24110,N_20636,N_22307);
nor U24111 (N_24111,N_21111,N_20613);
or U24112 (N_24112,N_21472,N_20450);
or U24113 (N_24113,N_22248,N_21542);
nor U24114 (N_24114,N_21228,N_20566);
nand U24115 (N_24115,N_22179,N_20664);
nand U24116 (N_24116,N_20366,N_20113);
or U24117 (N_24117,N_21156,N_21078);
nor U24118 (N_24118,N_21000,N_21421);
xnor U24119 (N_24119,N_21243,N_22229);
nor U24120 (N_24120,N_22403,N_20221);
nand U24121 (N_24121,N_21857,N_22129);
and U24122 (N_24122,N_21035,N_21713);
nand U24123 (N_24123,N_22045,N_21659);
nand U24124 (N_24124,N_20519,N_20668);
nand U24125 (N_24125,N_22075,N_20332);
nor U24126 (N_24126,N_22360,N_21888);
nand U24127 (N_24127,N_20464,N_21770);
nor U24128 (N_24128,N_21906,N_20553);
nor U24129 (N_24129,N_20510,N_22242);
xor U24130 (N_24130,N_21776,N_21905);
nand U24131 (N_24131,N_21521,N_22018);
or U24132 (N_24132,N_21554,N_22321);
xor U24133 (N_24133,N_20249,N_20776);
and U24134 (N_24134,N_20433,N_20197);
nand U24135 (N_24135,N_20780,N_20944);
xor U24136 (N_24136,N_20163,N_21044);
or U24137 (N_24137,N_21277,N_20493);
and U24138 (N_24138,N_20901,N_22354);
xor U24139 (N_24139,N_21814,N_21146);
nand U24140 (N_24140,N_21112,N_22214);
xor U24141 (N_24141,N_20099,N_21615);
nor U24142 (N_24142,N_20095,N_22380);
nand U24143 (N_24143,N_21695,N_20975);
and U24144 (N_24144,N_20356,N_20949);
and U24145 (N_24145,N_21967,N_22433);
nand U24146 (N_24146,N_21317,N_21710);
nand U24147 (N_24147,N_20459,N_21499);
nand U24148 (N_24148,N_20827,N_21207);
nor U24149 (N_24149,N_20793,N_21056);
xor U24150 (N_24150,N_20772,N_21752);
xor U24151 (N_24151,N_20780,N_21012);
or U24152 (N_24152,N_21397,N_20429);
and U24153 (N_24153,N_21692,N_21959);
xor U24154 (N_24154,N_22123,N_22352);
nor U24155 (N_24155,N_21226,N_21489);
or U24156 (N_24156,N_21451,N_22417);
nor U24157 (N_24157,N_20999,N_20064);
or U24158 (N_24158,N_21571,N_21632);
nand U24159 (N_24159,N_20071,N_20245);
or U24160 (N_24160,N_20063,N_20773);
nand U24161 (N_24161,N_22043,N_21662);
or U24162 (N_24162,N_20861,N_22255);
xor U24163 (N_24163,N_21234,N_22343);
nor U24164 (N_24164,N_22394,N_21042);
nand U24165 (N_24165,N_21756,N_21415);
and U24166 (N_24166,N_20169,N_21734);
xnor U24167 (N_24167,N_20840,N_22282);
and U24168 (N_24168,N_20842,N_21788);
nor U24169 (N_24169,N_21611,N_22491);
or U24170 (N_24170,N_20700,N_22390);
or U24171 (N_24171,N_21281,N_20207);
or U24172 (N_24172,N_20092,N_21661);
or U24173 (N_24173,N_20751,N_20720);
nand U24174 (N_24174,N_22314,N_22083);
or U24175 (N_24175,N_21561,N_20638);
or U24176 (N_24176,N_20113,N_21548);
or U24177 (N_24177,N_21325,N_20295);
nor U24178 (N_24178,N_21303,N_20706);
nor U24179 (N_24179,N_21931,N_21661);
xor U24180 (N_24180,N_21320,N_20001);
nor U24181 (N_24181,N_22173,N_20468);
or U24182 (N_24182,N_21191,N_21804);
nor U24183 (N_24183,N_20124,N_20049);
nor U24184 (N_24184,N_20307,N_20806);
or U24185 (N_24185,N_22157,N_21246);
and U24186 (N_24186,N_21596,N_20865);
xor U24187 (N_24187,N_21488,N_21016);
nand U24188 (N_24188,N_20187,N_21763);
or U24189 (N_24189,N_21890,N_22408);
nand U24190 (N_24190,N_22200,N_20685);
and U24191 (N_24191,N_21791,N_22443);
or U24192 (N_24192,N_21087,N_20009);
or U24193 (N_24193,N_21500,N_20730);
xnor U24194 (N_24194,N_20547,N_20536);
nor U24195 (N_24195,N_20561,N_21330);
nand U24196 (N_24196,N_20287,N_22177);
nand U24197 (N_24197,N_20551,N_21576);
and U24198 (N_24198,N_20442,N_21306);
nand U24199 (N_24199,N_20086,N_21794);
and U24200 (N_24200,N_20190,N_22115);
nand U24201 (N_24201,N_20325,N_20805);
nand U24202 (N_24202,N_22487,N_22105);
nor U24203 (N_24203,N_20746,N_21800);
and U24204 (N_24204,N_20523,N_20425);
or U24205 (N_24205,N_21690,N_22432);
and U24206 (N_24206,N_20099,N_20639);
xor U24207 (N_24207,N_20467,N_20125);
and U24208 (N_24208,N_20893,N_21845);
or U24209 (N_24209,N_20602,N_21131);
nor U24210 (N_24210,N_20928,N_21887);
or U24211 (N_24211,N_20979,N_21303);
or U24212 (N_24212,N_21533,N_22345);
nand U24213 (N_24213,N_21759,N_21750);
xnor U24214 (N_24214,N_21795,N_21025);
or U24215 (N_24215,N_21253,N_20328);
nand U24216 (N_24216,N_21707,N_21106);
nand U24217 (N_24217,N_21872,N_20099);
or U24218 (N_24218,N_21327,N_20554);
nor U24219 (N_24219,N_21460,N_21665);
nor U24220 (N_24220,N_21617,N_20868);
nand U24221 (N_24221,N_20988,N_22066);
and U24222 (N_24222,N_21263,N_20357);
xor U24223 (N_24223,N_22370,N_20542);
nor U24224 (N_24224,N_21329,N_21059);
or U24225 (N_24225,N_21062,N_20396);
and U24226 (N_24226,N_21770,N_20814);
or U24227 (N_24227,N_20137,N_21869);
or U24228 (N_24228,N_20360,N_20327);
or U24229 (N_24229,N_20908,N_21431);
and U24230 (N_24230,N_20185,N_21893);
nor U24231 (N_24231,N_21860,N_21486);
nor U24232 (N_24232,N_21558,N_21944);
or U24233 (N_24233,N_21976,N_20885);
xnor U24234 (N_24234,N_21092,N_20950);
or U24235 (N_24235,N_21761,N_21162);
and U24236 (N_24236,N_21757,N_21961);
xnor U24237 (N_24237,N_20026,N_21424);
or U24238 (N_24238,N_22458,N_20299);
nor U24239 (N_24239,N_20303,N_21939);
xnor U24240 (N_24240,N_20988,N_20883);
nor U24241 (N_24241,N_20573,N_21901);
nor U24242 (N_24242,N_20752,N_21513);
nor U24243 (N_24243,N_21004,N_21469);
nor U24244 (N_24244,N_20179,N_21932);
xnor U24245 (N_24245,N_22015,N_20857);
nand U24246 (N_24246,N_21027,N_21918);
nor U24247 (N_24247,N_21963,N_22098);
and U24248 (N_24248,N_21301,N_20340);
xnor U24249 (N_24249,N_22052,N_20601);
nor U24250 (N_24250,N_22212,N_21997);
nand U24251 (N_24251,N_20143,N_20262);
xnor U24252 (N_24252,N_22399,N_22340);
nor U24253 (N_24253,N_20267,N_21780);
nor U24254 (N_24254,N_22247,N_20919);
xnor U24255 (N_24255,N_20324,N_20450);
and U24256 (N_24256,N_22415,N_22124);
nand U24257 (N_24257,N_20297,N_21966);
nor U24258 (N_24258,N_21169,N_20827);
and U24259 (N_24259,N_21801,N_20595);
or U24260 (N_24260,N_22138,N_21202);
and U24261 (N_24261,N_21199,N_21294);
nor U24262 (N_24262,N_21203,N_21166);
nor U24263 (N_24263,N_20777,N_20250);
nand U24264 (N_24264,N_20499,N_22328);
xnor U24265 (N_24265,N_20194,N_20514);
and U24266 (N_24266,N_21924,N_22415);
nor U24267 (N_24267,N_21651,N_20588);
or U24268 (N_24268,N_20458,N_20814);
nor U24269 (N_24269,N_21467,N_20482);
and U24270 (N_24270,N_20462,N_21754);
xor U24271 (N_24271,N_22385,N_20265);
or U24272 (N_24272,N_20675,N_20870);
or U24273 (N_24273,N_20242,N_22480);
xor U24274 (N_24274,N_21094,N_21500);
nand U24275 (N_24275,N_21608,N_20234);
nand U24276 (N_24276,N_21864,N_20156);
nand U24277 (N_24277,N_20312,N_20204);
nor U24278 (N_24278,N_21637,N_20668);
nand U24279 (N_24279,N_20883,N_21162);
nor U24280 (N_24280,N_21611,N_21813);
or U24281 (N_24281,N_21212,N_21042);
nand U24282 (N_24282,N_20674,N_22393);
xnor U24283 (N_24283,N_21883,N_21173);
nor U24284 (N_24284,N_21639,N_22383);
nor U24285 (N_24285,N_21953,N_21098);
xor U24286 (N_24286,N_20171,N_21923);
or U24287 (N_24287,N_22102,N_22062);
nand U24288 (N_24288,N_21168,N_20451);
and U24289 (N_24289,N_21581,N_20142);
nor U24290 (N_24290,N_22450,N_20119);
or U24291 (N_24291,N_20373,N_21510);
and U24292 (N_24292,N_22378,N_20020);
nor U24293 (N_24293,N_21208,N_21415);
and U24294 (N_24294,N_22138,N_22192);
nor U24295 (N_24295,N_22474,N_20238);
and U24296 (N_24296,N_20031,N_20943);
nor U24297 (N_24297,N_20723,N_20624);
and U24298 (N_24298,N_22065,N_21096);
and U24299 (N_24299,N_21248,N_22057);
nor U24300 (N_24300,N_21696,N_20492);
nand U24301 (N_24301,N_21126,N_20304);
or U24302 (N_24302,N_20033,N_21657);
xor U24303 (N_24303,N_21892,N_21375);
nor U24304 (N_24304,N_22168,N_22459);
xor U24305 (N_24305,N_20810,N_21601);
or U24306 (N_24306,N_20769,N_20472);
nand U24307 (N_24307,N_21790,N_21919);
or U24308 (N_24308,N_21245,N_22274);
nor U24309 (N_24309,N_20137,N_20721);
xor U24310 (N_24310,N_21813,N_22178);
and U24311 (N_24311,N_20249,N_21053);
nand U24312 (N_24312,N_20549,N_21355);
and U24313 (N_24313,N_20909,N_20789);
xor U24314 (N_24314,N_20538,N_21386);
xnor U24315 (N_24315,N_20648,N_21862);
nor U24316 (N_24316,N_20028,N_22018);
nand U24317 (N_24317,N_21403,N_21488);
nand U24318 (N_24318,N_21921,N_21168);
nor U24319 (N_24319,N_20327,N_20826);
and U24320 (N_24320,N_21819,N_22407);
or U24321 (N_24321,N_20178,N_20068);
xor U24322 (N_24322,N_20039,N_22265);
or U24323 (N_24323,N_21579,N_21945);
or U24324 (N_24324,N_21077,N_21372);
nand U24325 (N_24325,N_20778,N_20659);
xnor U24326 (N_24326,N_22426,N_21778);
nor U24327 (N_24327,N_20939,N_20648);
xor U24328 (N_24328,N_21157,N_22305);
nand U24329 (N_24329,N_21806,N_20519);
and U24330 (N_24330,N_20921,N_21437);
xnor U24331 (N_24331,N_21872,N_22305);
nand U24332 (N_24332,N_20305,N_20408);
or U24333 (N_24333,N_21536,N_20111);
nor U24334 (N_24334,N_21396,N_20371);
xnor U24335 (N_24335,N_21867,N_20881);
nand U24336 (N_24336,N_21440,N_21217);
nand U24337 (N_24337,N_21742,N_22060);
and U24338 (N_24338,N_22334,N_20177);
nand U24339 (N_24339,N_20546,N_21463);
nand U24340 (N_24340,N_21053,N_21400);
xnor U24341 (N_24341,N_22371,N_21781);
and U24342 (N_24342,N_21901,N_21308);
or U24343 (N_24343,N_21752,N_20469);
and U24344 (N_24344,N_21600,N_21439);
xnor U24345 (N_24345,N_20581,N_21933);
xnor U24346 (N_24346,N_22328,N_20690);
or U24347 (N_24347,N_20814,N_20865);
xnor U24348 (N_24348,N_21936,N_21350);
and U24349 (N_24349,N_21119,N_22366);
and U24350 (N_24350,N_21415,N_21015);
nor U24351 (N_24351,N_20162,N_21048);
xor U24352 (N_24352,N_21039,N_21234);
and U24353 (N_24353,N_21539,N_20423);
and U24354 (N_24354,N_21660,N_22362);
and U24355 (N_24355,N_21142,N_22394);
or U24356 (N_24356,N_21184,N_21639);
or U24357 (N_24357,N_20988,N_20447);
nor U24358 (N_24358,N_21455,N_22365);
or U24359 (N_24359,N_21584,N_20371);
nor U24360 (N_24360,N_22007,N_20704);
and U24361 (N_24361,N_21664,N_20709);
or U24362 (N_24362,N_21608,N_21327);
xor U24363 (N_24363,N_21561,N_20959);
or U24364 (N_24364,N_22122,N_20525);
nand U24365 (N_24365,N_21306,N_21323);
nand U24366 (N_24366,N_20788,N_21495);
and U24367 (N_24367,N_21943,N_21460);
and U24368 (N_24368,N_20364,N_20871);
and U24369 (N_24369,N_22221,N_20837);
xor U24370 (N_24370,N_21208,N_20100);
or U24371 (N_24371,N_21489,N_20428);
or U24372 (N_24372,N_20561,N_21194);
and U24373 (N_24373,N_20500,N_21568);
nand U24374 (N_24374,N_20497,N_21153);
nand U24375 (N_24375,N_20400,N_20402);
and U24376 (N_24376,N_20801,N_20212);
xnor U24377 (N_24377,N_20959,N_21795);
or U24378 (N_24378,N_20618,N_21824);
nand U24379 (N_24379,N_20561,N_20007);
and U24380 (N_24380,N_22415,N_21041);
xor U24381 (N_24381,N_21183,N_21757);
or U24382 (N_24382,N_21653,N_21916);
nand U24383 (N_24383,N_20991,N_20150);
nand U24384 (N_24384,N_20797,N_21698);
nor U24385 (N_24385,N_20537,N_21343);
nand U24386 (N_24386,N_22367,N_21422);
nand U24387 (N_24387,N_21715,N_21782);
nand U24388 (N_24388,N_21140,N_20975);
xor U24389 (N_24389,N_22399,N_21596);
nor U24390 (N_24390,N_21414,N_20460);
xnor U24391 (N_24391,N_21491,N_21299);
nor U24392 (N_24392,N_22194,N_20146);
xor U24393 (N_24393,N_21923,N_21872);
nand U24394 (N_24394,N_20718,N_21665);
and U24395 (N_24395,N_21314,N_22336);
xnor U24396 (N_24396,N_21375,N_20325);
xor U24397 (N_24397,N_21795,N_22058);
and U24398 (N_24398,N_20349,N_22297);
nor U24399 (N_24399,N_21781,N_20297);
nand U24400 (N_24400,N_21178,N_22378);
nand U24401 (N_24401,N_22292,N_21998);
or U24402 (N_24402,N_21024,N_21484);
xnor U24403 (N_24403,N_20827,N_21354);
xor U24404 (N_24404,N_21308,N_20903);
and U24405 (N_24405,N_21141,N_20337);
nand U24406 (N_24406,N_20529,N_20031);
or U24407 (N_24407,N_21547,N_20431);
and U24408 (N_24408,N_20942,N_20197);
and U24409 (N_24409,N_22083,N_21652);
nand U24410 (N_24410,N_22409,N_20998);
and U24411 (N_24411,N_20545,N_22308);
nor U24412 (N_24412,N_22122,N_20316);
nor U24413 (N_24413,N_20754,N_20147);
nand U24414 (N_24414,N_20561,N_20594);
or U24415 (N_24415,N_20651,N_21576);
xnor U24416 (N_24416,N_21653,N_21299);
and U24417 (N_24417,N_21605,N_20004);
xnor U24418 (N_24418,N_22469,N_21748);
nor U24419 (N_24419,N_22409,N_21120);
and U24420 (N_24420,N_22208,N_22248);
nand U24421 (N_24421,N_22168,N_21930);
nand U24422 (N_24422,N_20731,N_20216);
xnor U24423 (N_24423,N_20096,N_21089);
nor U24424 (N_24424,N_21028,N_21241);
xnor U24425 (N_24425,N_20676,N_21317);
or U24426 (N_24426,N_20850,N_22069);
xor U24427 (N_24427,N_22199,N_20179);
xnor U24428 (N_24428,N_22477,N_20530);
xnor U24429 (N_24429,N_21822,N_21909);
and U24430 (N_24430,N_20980,N_20877);
and U24431 (N_24431,N_20440,N_20526);
xnor U24432 (N_24432,N_20260,N_20332);
xor U24433 (N_24433,N_20383,N_21065);
and U24434 (N_24434,N_21535,N_22379);
nor U24435 (N_24435,N_20184,N_20059);
nand U24436 (N_24436,N_21174,N_21282);
nand U24437 (N_24437,N_21541,N_20266);
nor U24438 (N_24438,N_21076,N_20855);
and U24439 (N_24439,N_22019,N_20708);
nor U24440 (N_24440,N_21498,N_21386);
or U24441 (N_24441,N_22419,N_20000);
and U24442 (N_24442,N_20289,N_21789);
xnor U24443 (N_24443,N_22132,N_21771);
nand U24444 (N_24444,N_20097,N_21576);
or U24445 (N_24445,N_20941,N_20187);
nand U24446 (N_24446,N_22067,N_22445);
xnor U24447 (N_24447,N_20442,N_21192);
nand U24448 (N_24448,N_22206,N_20609);
xnor U24449 (N_24449,N_20124,N_20998);
nand U24450 (N_24450,N_20610,N_21735);
and U24451 (N_24451,N_21014,N_20733);
nor U24452 (N_24452,N_21114,N_22366);
xnor U24453 (N_24453,N_20600,N_20086);
and U24454 (N_24454,N_20511,N_21789);
or U24455 (N_24455,N_20620,N_21754);
xor U24456 (N_24456,N_20924,N_21915);
nor U24457 (N_24457,N_21616,N_21788);
nor U24458 (N_24458,N_21188,N_22028);
and U24459 (N_24459,N_21782,N_20962);
nand U24460 (N_24460,N_20685,N_22498);
and U24461 (N_24461,N_20672,N_20038);
xnor U24462 (N_24462,N_21459,N_21354);
and U24463 (N_24463,N_22179,N_22460);
nand U24464 (N_24464,N_21469,N_20101);
and U24465 (N_24465,N_21335,N_20590);
xor U24466 (N_24466,N_21710,N_21354);
nor U24467 (N_24467,N_21159,N_21359);
and U24468 (N_24468,N_20136,N_22216);
nor U24469 (N_24469,N_20030,N_21320);
nand U24470 (N_24470,N_22090,N_21283);
nand U24471 (N_24471,N_21478,N_20732);
xnor U24472 (N_24472,N_20627,N_21278);
nand U24473 (N_24473,N_21501,N_21311);
xnor U24474 (N_24474,N_21901,N_21060);
xor U24475 (N_24475,N_22114,N_21462);
nand U24476 (N_24476,N_20290,N_20536);
or U24477 (N_24477,N_20218,N_20277);
or U24478 (N_24478,N_20123,N_20856);
xnor U24479 (N_24479,N_22119,N_20407);
and U24480 (N_24480,N_21288,N_21312);
nand U24481 (N_24481,N_20392,N_20027);
nand U24482 (N_24482,N_20264,N_20114);
nor U24483 (N_24483,N_21547,N_21135);
or U24484 (N_24484,N_20231,N_20403);
nor U24485 (N_24485,N_20127,N_20820);
xnor U24486 (N_24486,N_21115,N_21683);
nor U24487 (N_24487,N_21109,N_22102);
xor U24488 (N_24488,N_21430,N_21782);
xor U24489 (N_24489,N_22056,N_20188);
nor U24490 (N_24490,N_21041,N_20836);
nand U24491 (N_24491,N_22230,N_21324);
and U24492 (N_24492,N_22041,N_21810);
xor U24493 (N_24493,N_20244,N_21733);
xnor U24494 (N_24494,N_20105,N_20496);
nor U24495 (N_24495,N_21623,N_21328);
nand U24496 (N_24496,N_21550,N_20062);
and U24497 (N_24497,N_20269,N_20249);
or U24498 (N_24498,N_20794,N_21698);
or U24499 (N_24499,N_21865,N_21125);
nand U24500 (N_24500,N_21602,N_22259);
or U24501 (N_24501,N_20385,N_21854);
nand U24502 (N_24502,N_21451,N_22328);
xnor U24503 (N_24503,N_20432,N_21904);
or U24504 (N_24504,N_21410,N_22467);
or U24505 (N_24505,N_20181,N_21704);
nand U24506 (N_24506,N_20777,N_21689);
xnor U24507 (N_24507,N_22349,N_21267);
nor U24508 (N_24508,N_21242,N_20284);
nand U24509 (N_24509,N_22468,N_21691);
nor U24510 (N_24510,N_22269,N_20152);
or U24511 (N_24511,N_20680,N_20633);
nand U24512 (N_24512,N_21399,N_20383);
and U24513 (N_24513,N_20617,N_20469);
nor U24514 (N_24514,N_20242,N_20123);
xor U24515 (N_24515,N_21686,N_21992);
or U24516 (N_24516,N_21337,N_21856);
xnor U24517 (N_24517,N_22095,N_21346);
or U24518 (N_24518,N_22319,N_21641);
or U24519 (N_24519,N_21643,N_22334);
and U24520 (N_24520,N_21121,N_20523);
nand U24521 (N_24521,N_20217,N_20507);
nand U24522 (N_24522,N_20118,N_22040);
or U24523 (N_24523,N_22474,N_21651);
nand U24524 (N_24524,N_20542,N_20402);
nor U24525 (N_24525,N_21280,N_20672);
nand U24526 (N_24526,N_20030,N_20738);
nor U24527 (N_24527,N_20592,N_21196);
or U24528 (N_24528,N_21456,N_21116);
or U24529 (N_24529,N_22112,N_21231);
or U24530 (N_24530,N_20023,N_21255);
and U24531 (N_24531,N_20506,N_21171);
nand U24532 (N_24532,N_21974,N_20217);
or U24533 (N_24533,N_22428,N_20180);
xor U24534 (N_24534,N_21133,N_20606);
nand U24535 (N_24535,N_21119,N_20466);
and U24536 (N_24536,N_21136,N_20626);
and U24537 (N_24537,N_22418,N_20093);
and U24538 (N_24538,N_20100,N_20468);
xnor U24539 (N_24539,N_20496,N_20407);
xor U24540 (N_24540,N_22182,N_22152);
xnor U24541 (N_24541,N_21798,N_21414);
nand U24542 (N_24542,N_22049,N_20659);
or U24543 (N_24543,N_20217,N_20649);
and U24544 (N_24544,N_21893,N_21775);
and U24545 (N_24545,N_21602,N_22496);
or U24546 (N_24546,N_20975,N_20718);
or U24547 (N_24547,N_21604,N_21220);
nor U24548 (N_24548,N_20427,N_21908);
nor U24549 (N_24549,N_21557,N_21585);
or U24550 (N_24550,N_21503,N_22128);
nor U24551 (N_24551,N_22441,N_21970);
and U24552 (N_24552,N_21912,N_22405);
and U24553 (N_24553,N_21111,N_20040);
and U24554 (N_24554,N_22048,N_22456);
or U24555 (N_24555,N_21767,N_21785);
xnor U24556 (N_24556,N_21788,N_20923);
and U24557 (N_24557,N_20888,N_21050);
xnor U24558 (N_24558,N_20701,N_21409);
nand U24559 (N_24559,N_22073,N_20408);
and U24560 (N_24560,N_21976,N_21283);
and U24561 (N_24561,N_21640,N_21660);
nor U24562 (N_24562,N_20383,N_22020);
nand U24563 (N_24563,N_20455,N_22297);
nand U24564 (N_24564,N_22057,N_21389);
and U24565 (N_24565,N_21864,N_21715);
or U24566 (N_24566,N_22105,N_21566);
or U24567 (N_24567,N_20250,N_21352);
and U24568 (N_24568,N_20327,N_21025);
xnor U24569 (N_24569,N_21231,N_21639);
or U24570 (N_24570,N_21726,N_20017);
xor U24571 (N_24571,N_20574,N_20820);
xor U24572 (N_24572,N_21691,N_21950);
or U24573 (N_24573,N_20312,N_20785);
nor U24574 (N_24574,N_22232,N_21500);
nand U24575 (N_24575,N_21446,N_21357);
or U24576 (N_24576,N_21091,N_20838);
nand U24577 (N_24577,N_22167,N_20484);
and U24578 (N_24578,N_20211,N_20154);
nand U24579 (N_24579,N_21518,N_21946);
nor U24580 (N_24580,N_20773,N_21222);
xnor U24581 (N_24581,N_21173,N_20159);
and U24582 (N_24582,N_21037,N_21936);
nand U24583 (N_24583,N_21337,N_21518);
xor U24584 (N_24584,N_20367,N_21473);
or U24585 (N_24585,N_21799,N_21286);
nor U24586 (N_24586,N_20544,N_20549);
and U24587 (N_24587,N_21032,N_21928);
and U24588 (N_24588,N_20979,N_21706);
nor U24589 (N_24589,N_20407,N_20103);
xor U24590 (N_24590,N_21993,N_21136);
nand U24591 (N_24591,N_20985,N_21475);
nor U24592 (N_24592,N_21341,N_22041);
xnor U24593 (N_24593,N_21531,N_20133);
nand U24594 (N_24594,N_22000,N_22312);
and U24595 (N_24595,N_20031,N_20269);
or U24596 (N_24596,N_22174,N_22206);
or U24597 (N_24597,N_21602,N_21397);
or U24598 (N_24598,N_20832,N_21718);
xnor U24599 (N_24599,N_20632,N_20552);
xor U24600 (N_24600,N_21860,N_20744);
nand U24601 (N_24601,N_20016,N_22399);
or U24602 (N_24602,N_21137,N_22496);
or U24603 (N_24603,N_21747,N_22296);
or U24604 (N_24604,N_20903,N_21637);
and U24605 (N_24605,N_20400,N_22241);
and U24606 (N_24606,N_20367,N_20643);
xnor U24607 (N_24607,N_20707,N_20329);
or U24608 (N_24608,N_21668,N_20980);
xor U24609 (N_24609,N_21892,N_22422);
or U24610 (N_24610,N_21364,N_21957);
nor U24611 (N_24611,N_21868,N_20193);
nand U24612 (N_24612,N_20911,N_21997);
xor U24613 (N_24613,N_21018,N_20367);
xor U24614 (N_24614,N_20847,N_21175);
or U24615 (N_24615,N_20464,N_20030);
nor U24616 (N_24616,N_20119,N_22211);
and U24617 (N_24617,N_21629,N_21149);
nand U24618 (N_24618,N_22364,N_21960);
xor U24619 (N_24619,N_22395,N_20735);
xor U24620 (N_24620,N_20890,N_20614);
xor U24621 (N_24621,N_21704,N_21514);
and U24622 (N_24622,N_20553,N_21802);
xnor U24623 (N_24623,N_21367,N_21490);
and U24624 (N_24624,N_21646,N_20444);
xnor U24625 (N_24625,N_20350,N_21549);
xor U24626 (N_24626,N_20448,N_22185);
and U24627 (N_24627,N_21454,N_21490);
and U24628 (N_24628,N_20171,N_21768);
nor U24629 (N_24629,N_22050,N_21389);
nand U24630 (N_24630,N_20950,N_20003);
nand U24631 (N_24631,N_21554,N_20197);
nand U24632 (N_24632,N_22350,N_22241);
nand U24633 (N_24633,N_21953,N_20438);
and U24634 (N_24634,N_21178,N_21986);
or U24635 (N_24635,N_20563,N_21045);
xnor U24636 (N_24636,N_22127,N_21174);
and U24637 (N_24637,N_20454,N_20927);
nor U24638 (N_24638,N_20120,N_20602);
and U24639 (N_24639,N_20482,N_21401);
and U24640 (N_24640,N_21166,N_20946);
nand U24641 (N_24641,N_20056,N_20462);
and U24642 (N_24642,N_22494,N_20687);
or U24643 (N_24643,N_21939,N_21760);
and U24644 (N_24644,N_20983,N_21933);
nand U24645 (N_24645,N_21355,N_20195);
nor U24646 (N_24646,N_21124,N_21902);
or U24647 (N_24647,N_21754,N_20955);
or U24648 (N_24648,N_20721,N_20343);
nand U24649 (N_24649,N_20808,N_20700);
nor U24650 (N_24650,N_20729,N_20756);
and U24651 (N_24651,N_21159,N_21437);
and U24652 (N_24652,N_20201,N_21337);
xnor U24653 (N_24653,N_20327,N_21450);
and U24654 (N_24654,N_22133,N_20615);
xnor U24655 (N_24655,N_21010,N_22465);
xnor U24656 (N_24656,N_21536,N_22233);
nand U24657 (N_24657,N_22181,N_21279);
nor U24658 (N_24658,N_21920,N_22361);
or U24659 (N_24659,N_20635,N_21024);
nand U24660 (N_24660,N_21580,N_22332);
or U24661 (N_24661,N_21208,N_20368);
and U24662 (N_24662,N_22228,N_21065);
xor U24663 (N_24663,N_22199,N_20370);
xnor U24664 (N_24664,N_20965,N_21455);
and U24665 (N_24665,N_22044,N_22376);
nor U24666 (N_24666,N_21206,N_20412);
xor U24667 (N_24667,N_20881,N_20834);
nor U24668 (N_24668,N_20748,N_20006);
and U24669 (N_24669,N_20358,N_22382);
xor U24670 (N_24670,N_21690,N_20110);
and U24671 (N_24671,N_21666,N_20189);
nand U24672 (N_24672,N_20436,N_22119);
xor U24673 (N_24673,N_21403,N_20532);
and U24674 (N_24674,N_21162,N_21508);
nand U24675 (N_24675,N_20934,N_21881);
or U24676 (N_24676,N_20861,N_20642);
nor U24677 (N_24677,N_20058,N_20618);
nand U24678 (N_24678,N_21377,N_20230);
nand U24679 (N_24679,N_21143,N_20444);
nand U24680 (N_24680,N_21901,N_21838);
nor U24681 (N_24681,N_21184,N_20790);
nand U24682 (N_24682,N_21947,N_21576);
or U24683 (N_24683,N_20373,N_21346);
or U24684 (N_24684,N_20674,N_21371);
xnor U24685 (N_24685,N_20503,N_20817);
and U24686 (N_24686,N_21531,N_20678);
nand U24687 (N_24687,N_21571,N_20807);
nand U24688 (N_24688,N_22127,N_21845);
or U24689 (N_24689,N_22165,N_22049);
xor U24690 (N_24690,N_21476,N_21955);
nand U24691 (N_24691,N_20619,N_21833);
or U24692 (N_24692,N_21042,N_20265);
or U24693 (N_24693,N_20243,N_22409);
or U24694 (N_24694,N_22442,N_22065);
or U24695 (N_24695,N_20972,N_20211);
and U24696 (N_24696,N_22265,N_20859);
nor U24697 (N_24697,N_22278,N_21484);
xnor U24698 (N_24698,N_20196,N_22210);
xor U24699 (N_24699,N_20981,N_22047);
or U24700 (N_24700,N_20061,N_20716);
or U24701 (N_24701,N_20511,N_21599);
nand U24702 (N_24702,N_21838,N_21695);
xor U24703 (N_24703,N_21050,N_21971);
nand U24704 (N_24704,N_20242,N_20826);
nor U24705 (N_24705,N_21661,N_21131);
or U24706 (N_24706,N_21457,N_21645);
and U24707 (N_24707,N_20870,N_22146);
and U24708 (N_24708,N_20634,N_21828);
nand U24709 (N_24709,N_22111,N_21123);
nor U24710 (N_24710,N_21383,N_20520);
nor U24711 (N_24711,N_21386,N_20769);
and U24712 (N_24712,N_21990,N_20558);
nor U24713 (N_24713,N_21919,N_20072);
or U24714 (N_24714,N_20341,N_20794);
xnor U24715 (N_24715,N_22221,N_21306);
nor U24716 (N_24716,N_20231,N_20156);
xnor U24717 (N_24717,N_20343,N_22380);
or U24718 (N_24718,N_21010,N_20816);
nand U24719 (N_24719,N_21258,N_22390);
and U24720 (N_24720,N_21495,N_20612);
xor U24721 (N_24721,N_21764,N_21083);
xnor U24722 (N_24722,N_22164,N_20717);
nor U24723 (N_24723,N_20783,N_21524);
and U24724 (N_24724,N_21375,N_21544);
nor U24725 (N_24725,N_21630,N_21196);
xor U24726 (N_24726,N_20774,N_20254);
nor U24727 (N_24727,N_20713,N_20318);
or U24728 (N_24728,N_20699,N_21333);
nor U24729 (N_24729,N_22283,N_20846);
and U24730 (N_24730,N_20338,N_20183);
xnor U24731 (N_24731,N_21955,N_20350);
nand U24732 (N_24732,N_21922,N_21513);
xor U24733 (N_24733,N_20252,N_21257);
and U24734 (N_24734,N_20389,N_21008);
and U24735 (N_24735,N_20861,N_20871);
nor U24736 (N_24736,N_21499,N_20322);
or U24737 (N_24737,N_20066,N_22304);
nand U24738 (N_24738,N_20845,N_21108);
nor U24739 (N_24739,N_21276,N_22125);
or U24740 (N_24740,N_22106,N_21274);
nor U24741 (N_24741,N_20455,N_21476);
nor U24742 (N_24742,N_21324,N_22488);
and U24743 (N_24743,N_20346,N_20766);
and U24744 (N_24744,N_20982,N_21832);
or U24745 (N_24745,N_22123,N_20302);
nor U24746 (N_24746,N_20461,N_22475);
xor U24747 (N_24747,N_20978,N_22246);
or U24748 (N_24748,N_20388,N_22336);
xor U24749 (N_24749,N_20595,N_21277);
and U24750 (N_24750,N_22214,N_22277);
and U24751 (N_24751,N_20574,N_21796);
or U24752 (N_24752,N_22141,N_21657);
and U24753 (N_24753,N_21286,N_22323);
nand U24754 (N_24754,N_22261,N_21241);
nand U24755 (N_24755,N_21291,N_21408);
or U24756 (N_24756,N_20491,N_22168);
and U24757 (N_24757,N_21664,N_20225);
nand U24758 (N_24758,N_21293,N_20500);
nor U24759 (N_24759,N_21891,N_20758);
and U24760 (N_24760,N_20275,N_22211);
and U24761 (N_24761,N_20056,N_20220);
nand U24762 (N_24762,N_21883,N_21985);
nand U24763 (N_24763,N_22089,N_20469);
nor U24764 (N_24764,N_22105,N_20112);
nand U24765 (N_24765,N_21408,N_21466);
nor U24766 (N_24766,N_20665,N_22288);
and U24767 (N_24767,N_20163,N_21596);
xor U24768 (N_24768,N_20398,N_20087);
nand U24769 (N_24769,N_20208,N_20852);
xor U24770 (N_24770,N_21215,N_21433);
or U24771 (N_24771,N_20104,N_21782);
nand U24772 (N_24772,N_20802,N_21820);
and U24773 (N_24773,N_20851,N_22474);
and U24774 (N_24774,N_20327,N_20512);
nor U24775 (N_24775,N_21114,N_22063);
xor U24776 (N_24776,N_21116,N_21601);
xor U24777 (N_24777,N_20824,N_20653);
xor U24778 (N_24778,N_20154,N_20429);
xor U24779 (N_24779,N_20773,N_20865);
xnor U24780 (N_24780,N_22403,N_22073);
and U24781 (N_24781,N_22236,N_20571);
xor U24782 (N_24782,N_20355,N_21944);
or U24783 (N_24783,N_20274,N_20405);
xor U24784 (N_24784,N_20731,N_21313);
nor U24785 (N_24785,N_21956,N_21996);
and U24786 (N_24786,N_21751,N_21069);
xor U24787 (N_24787,N_20869,N_20077);
or U24788 (N_24788,N_20742,N_20593);
and U24789 (N_24789,N_20106,N_22057);
nor U24790 (N_24790,N_20913,N_22249);
or U24791 (N_24791,N_21175,N_20287);
and U24792 (N_24792,N_22280,N_22428);
nand U24793 (N_24793,N_21650,N_20112);
xnor U24794 (N_24794,N_20368,N_21653);
or U24795 (N_24795,N_21825,N_20427);
xnor U24796 (N_24796,N_20795,N_22424);
or U24797 (N_24797,N_20678,N_21641);
and U24798 (N_24798,N_20040,N_22214);
nor U24799 (N_24799,N_22043,N_22224);
and U24800 (N_24800,N_21164,N_22328);
xnor U24801 (N_24801,N_20633,N_20911);
xnor U24802 (N_24802,N_22187,N_20236);
or U24803 (N_24803,N_22096,N_22198);
nand U24804 (N_24804,N_22388,N_20054);
or U24805 (N_24805,N_20989,N_21345);
or U24806 (N_24806,N_20262,N_20114);
and U24807 (N_24807,N_20190,N_21811);
nand U24808 (N_24808,N_21769,N_20335);
nand U24809 (N_24809,N_21647,N_21188);
xnor U24810 (N_24810,N_21663,N_20902);
and U24811 (N_24811,N_22224,N_20317);
or U24812 (N_24812,N_21381,N_22117);
xor U24813 (N_24813,N_20237,N_21023);
nand U24814 (N_24814,N_20768,N_20117);
nand U24815 (N_24815,N_22371,N_21546);
nor U24816 (N_24816,N_21269,N_21426);
nand U24817 (N_24817,N_21287,N_20293);
and U24818 (N_24818,N_21887,N_22111);
and U24819 (N_24819,N_20225,N_20842);
xnor U24820 (N_24820,N_20258,N_22417);
and U24821 (N_24821,N_20081,N_20020);
nor U24822 (N_24822,N_20648,N_20400);
nor U24823 (N_24823,N_20089,N_21060);
nand U24824 (N_24824,N_22270,N_20192);
nand U24825 (N_24825,N_22176,N_21684);
xor U24826 (N_24826,N_20499,N_20468);
xor U24827 (N_24827,N_21220,N_22259);
or U24828 (N_24828,N_20671,N_20554);
nor U24829 (N_24829,N_21517,N_20885);
xor U24830 (N_24830,N_20807,N_22045);
nand U24831 (N_24831,N_20225,N_21244);
nor U24832 (N_24832,N_20507,N_22391);
nor U24833 (N_24833,N_21731,N_21544);
nor U24834 (N_24834,N_21587,N_22091);
xnor U24835 (N_24835,N_22398,N_20122);
nor U24836 (N_24836,N_20846,N_21227);
or U24837 (N_24837,N_20129,N_21647);
nand U24838 (N_24838,N_21322,N_21658);
nor U24839 (N_24839,N_20780,N_22159);
nand U24840 (N_24840,N_20921,N_21793);
nand U24841 (N_24841,N_22479,N_21416);
nand U24842 (N_24842,N_21849,N_22336);
nor U24843 (N_24843,N_20518,N_20725);
xnor U24844 (N_24844,N_22323,N_21007);
nand U24845 (N_24845,N_21991,N_20309);
and U24846 (N_24846,N_22383,N_21872);
xor U24847 (N_24847,N_21116,N_21824);
or U24848 (N_24848,N_20080,N_22418);
xnor U24849 (N_24849,N_20864,N_22135);
xor U24850 (N_24850,N_21838,N_21519);
xnor U24851 (N_24851,N_21710,N_20032);
xnor U24852 (N_24852,N_21838,N_20563);
nand U24853 (N_24853,N_20634,N_21107);
nor U24854 (N_24854,N_22417,N_20527);
xnor U24855 (N_24855,N_22216,N_22229);
nand U24856 (N_24856,N_21893,N_21836);
xnor U24857 (N_24857,N_20301,N_20664);
nor U24858 (N_24858,N_21577,N_22036);
xnor U24859 (N_24859,N_21117,N_22073);
or U24860 (N_24860,N_22414,N_22330);
nand U24861 (N_24861,N_20586,N_21552);
or U24862 (N_24862,N_20084,N_20203);
and U24863 (N_24863,N_21623,N_21621);
and U24864 (N_24864,N_20233,N_20491);
nand U24865 (N_24865,N_22007,N_21190);
xor U24866 (N_24866,N_20939,N_22253);
nor U24867 (N_24867,N_22438,N_20240);
and U24868 (N_24868,N_22075,N_20432);
and U24869 (N_24869,N_22221,N_21436);
nor U24870 (N_24870,N_21634,N_20070);
or U24871 (N_24871,N_22448,N_21270);
nor U24872 (N_24872,N_20559,N_21004);
xnor U24873 (N_24873,N_20769,N_21120);
nor U24874 (N_24874,N_21187,N_20640);
xor U24875 (N_24875,N_21370,N_22063);
or U24876 (N_24876,N_21866,N_22011);
xnor U24877 (N_24877,N_20338,N_20559);
nand U24878 (N_24878,N_20127,N_21532);
xor U24879 (N_24879,N_21905,N_21551);
nor U24880 (N_24880,N_21812,N_21713);
or U24881 (N_24881,N_20848,N_22409);
nor U24882 (N_24882,N_21591,N_20889);
or U24883 (N_24883,N_20488,N_22452);
nand U24884 (N_24884,N_20060,N_20541);
nand U24885 (N_24885,N_20404,N_21947);
nor U24886 (N_24886,N_21213,N_21547);
xnor U24887 (N_24887,N_20968,N_22431);
or U24888 (N_24888,N_20155,N_21886);
xnor U24889 (N_24889,N_21137,N_21990);
nor U24890 (N_24890,N_21867,N_21712);
nand U24891 (N_24891,N_20180,N_20621);
or U24892 (N_24892,N_21961,N_20597);
and U24893 (N_24893,N_20081,N_21139);
xnor U24894 (N_24894,N_21249,N_21917);
and U24895 (N_24895,N_21619,N_22323);
and U24896 (N_24896,N_20002,N_21281);
nand U24897 (N_24897,N_22111,N_21476);
and U24898 (N_24898,N_20477,N_21591);
nand U24899 (N_24899,N_21285,N_21464);
xnor U24900 (N_24900,N_20778,N_22454);
or U24901 (N_24901,N_22497,N_20469);
and U24902 (N_24902,N_22296,N_20184);
nand U24903 (N_24903,N_22113,N_21485);
nand U24904 (N_24904,N_22056,N_22440);
nor U24905 (N_24905,N_21770,N_22284);
nand U24906 (N_24906,N_21510,N_20671);
nor U24907 (N_24907,N_20930,N_20711);
nor U24908 (N_24908,N_21017,N_20347);
and U24909 (N_24909,N_22467,N_20950);
nand U24910 (N_24910,N_20364,N_20404);
and U24911 (N_24911,N_20908,N_21051);
and U24912 (N_24912,N_20644,N_21763);
nor U24913 (N_24913,N_21773,N_20464);
or U24914 (N_24914,N_20807,N_20473);
and U24915 (N_24915,N_21008,N_21759);
xnor U24916 (N_24916,N_21504,N_22392);
nor U24917 (N_24917,N_22162,N_22128);
xnor U24918 (N_24918,N_21568,N_21004);
or U24919 (N_24919,N_20155,N_20370);
or U24920 (N_24920,N_20703,N_22297);
nor U24921 (N_24921,N_21610,N_20984);
nor U24922 (N_24922,N_21109,N_21627);
xnor U24923 (N_24923,N_20367,N_21074);
and U24924 (N_24924,N_20417,N_21780);
and U24925 (N_24925,N_21149,N_21320);
nor U24926 (N_24926,N_21014,N_20190);
nor U24927 (N_24927,N_20581,N_20749);
nor U24928 (N_24928,N_21813,N_21466);
or U24929 (N_24929,N_21700,N_20915);
xnor U24930 (N_24930,N_21040,N_21890);
xor U24931 (N_24931,N_21546,N_20659);
and U24932 (N_24932,N_20227,N_20164);
xor U24933 (N_24933,N_21563,N_22386);
nand U24934 (N_24934,N_21283,N_20341);
or U24935 (N_24935,N_21962,N_21926);
xnor U24936 (N_24936,N_21889,N_22097);
or U24937 (N_24937,N_20558,N_20087);
nand U24938 (N_24938,N_21697,N_22057);
or U24939 (N_24939,N_20834,N_21553);
and U24940 (N_24940,N_20039,N_21023);
or U24941 (N_24941,N_21941,N_21258);
xor U24942 (N_24942,N_21116,N_21642);
nand U24943 (N_24943,N_21321,N_21172);
nor U24944 (N_24944,N_22327,N_21949);
xnor U24945 (N_24945,N_21225,N_20668);
nand U24946 (N_24946,N_21761,N_21711);
xnor U24947 (N_24947,N_20537,N_21139);
nor U24948 (N_24948,N_20926,N_21264);
nor U24949 (N_24949,N_20705,N_22071);
and U24950 (N_24950,N_21311,N_22167);
or U24951 (N_24951,N_20207,N_22458);
or U24952 (N_24952,N_21911,N_21395);
or U24953 (N_24953,N_20636,N_21046);
or U24954 (N_24954,N_21450,N_20132);
xor U24955 (N_24955,N_22079,N_21211);
nand U24956 (N_24956,N_22397,N_21886);
xnor U24957 (N_24957,N_21324,N_22324);
xor U24958 (N_24958,N_20673,N_20904);
or U24959 (N_24959,N_20043,N_21624);
nand U24960 (N_24960,N_20177,N_22355);
and U24961 (N_24961,N_20246,N_21058);
nand U24962 (N_24962,N_22145,N_21244);
nor U24963 (N_24963,N_20056,N_21353);
or U24964 (N_24964,N_20316,N_20335);
nor U24965 (N_24965,N_22270,N_21110);
or U24966 (N_24966,N_21748,N_21321);
and U24967 (N_24967,N_22150,N_21707);
or U24968 (N_24968,N_20040,N_21059);
xor U24969 (N_24969,N_20238,N_20808);
nand U24970 (N_24970,N_21472,N_21585);
nand U24971 (N_24971,N_20581,N_22354);
nand U24972 (N_24972,N_20067,N_20028);
nor U24973 (N_24973,N_21205,N_21140);
xor U24974 (N_24974,N_21849,N_20706);
or U24975 (N_24975,N_22347,N_21200);
or U24976 (N_24976,N_21769,N_21658);
xor U24977 (N_24977,N_20266,N_21801);
or U24978 (N_24978,N_20462,N_21331);
nand U24979 (N_24979,N_20114,N_21778);
nand U24980 (N_24980,N_20786,N_21969);
and U24981 (N_24981,N_22211,N_21267);
nand U24982 (N_24982,N_20456,N_22092);
and U24983 (N_24983,N_21472,N_20447);
and U24984 (N_24984,N_20450,N_20093);
xor U24985 (N_24985,N_22198,N_21752);
and U24986 (N_24986,N_20490,N_20150);
and U24987 (N_24987,N_21139,N_21622);
nand U24988 (N_24988,N_22280,N_20739);
nand U24989 (N_24989,N_21077,N_20131);
and U24990 (N_24990,N_21608,N_20960);
and U24991 (N_24991,N_21805,N_22224);
or U24992 (N_24992,N_20987,N_22391);
or U24993 (N_24993,N_20063,N_20105);
xnor U24994 (N_24994,N_20274,N_20892);
nand U24995 (N_24995,N_22046,N_21101);
or U24996 (N_24996,N_20383,N_21428);
or U24997 (N_24997,N_20402,N_20552);
or U24998 (N_24998,N_20579,N_21674);
or U24999 (N_24999,N_20746,N_20702);
xor UO_0 (O_0,N_23492,N_23712);
xor UO_1 (O_1,N_22624,N_24065);
nor UO_2 (O_2,N_22746,N_23840);
nor UO_3 (O_3,N_24410,N_24292);
nor UO_4 (O_4,N_22994,N_24342);
nand UO_5 (O_5,N_22832,N_24205);
nor UO_6 (O_6,N_24710,N_22776);
and UO_7 (O_7,N_23613,N_24334);
or UO_8 (O_8,N_24793,N_23841);
and UO_9 (O_9,N_23667,N_22739);
or UO_10 (O_10,N_22753,N_23851);
or UO_11 (O_11,N_24878,N_24084);
or UO_12 (O_12,N_23450,N_24687);
and UO_13 (O_13,N_23551,N_23186);
xnor UO_14 (O_14,N_24962,N_24233);
nor UO_15 (O_15,N_24328,N_24248);
or UO_16 (O_16,N_22825,N_24970);
and UO_17 (O_17,N_24847,N_24034);
nand UO_18 (O_18,N_23955,N_24387);
nand UO_19 (O_19,N_24693,N_23499);
and UO_20 (O_20,N_23574,N_24299);
nor UO_21 (O_21,N_23232,N_22563);
nor UO_22 (O_22,N_23860,N_23548);
nand UO_23 (O_23,N_22916,N_23692);
and UO_24 (O_24,N_23282,N_23292);
or UO_25 (O_25,N_22521,N_24455);
nor UO_26 (O_26,N_24296,N_23979);
and UO_27 (O_27,N_22951,N_23188);
xor UO_28 (O_28,N_23842,N_22608);
xnor UO_29 (O_29,N_24649,N_23890);
nor UO_30 (O_30,N_23046,N_23828);
xor UO_31 (O_31,N_24005,N_24415);
nor UO_32 (O_32,N_24626,N_23318);
or UO_33 (O_33,N_24131,N_24185);
or UO_34 (O_34,N_23415,N_24460);
xnor UO_35 (O_35,N_24484,N_23988);
nor UO_36 (O_36,N_24853,N_23123);
nand UO_37 (O_37,N_24953,N_24020);
and UO_38 (O_38,N_24950,N_24492);
xor UO_39 (O_39,N_24906,N_23220);
xor UO_40 (O_40,N_22715,N_23767);
or UO_41 (O_41,N_24673,N_23383);
nor UO_42 (O_42,N_23049,N_23036);
nand UO_43 (O_43,N_22571,N_23482);
nand UO_44 (O_44,N_24527,N_22684);
nand UO_45 (O_45,N_23367,N_23958);
nand UO_46 (O_46,N_23020,N_24664);
and UO_47 (O_47,N_24766,N_24832);
or UO_48 (O_48,N_23946,N_24452);
xnor UO_49 (O_49,N_24273,N_24801);
xnor UO_50 (O_50,N_24163,N_23069);
xor UO_51 (O_51,N_22815,N_24930);
nor UO_52 (O_52,N_23016,N_22955);
nor UO_53 (O_53,N_22950,N_23187);
and UO_54 (O_54,N_22724,N_23353);
or UO_55 (O_55,N_23698,N_22827);
or UO_56 (O_56,N_23006,N_22519);
or UO_57 (O_57,N_24554,N_23409);
xnor UO_58 (O_58,N_22700,N_23075);
xnor UO_59 (O_59,N_23550,N_24317);
and UO_60 (O_60,N_24029,N_22819);
nor UO_61 (O_61,N_23330,N_24946);
and UO_62 (O_62,N_23470,N_24378);
nand UO_63 (O_63,N_23831,N_22796);
nor UO_64 (O_64,N_23673,N_22918);
nand UO_65 (O_65,N_22799,N_24918);
xnor UO_66 (O_66,N_23724,N_24954);
nand UO_67 (O_67,N_24340,N_24486);
and UO_68 (O_68,N_23182,N_22524);
nand UO_69 (O_69,N_23010,N_23568);
or UO_70 (O_70,N_24301,N_22894);
or UO_71 (O_71,N_24106,N_22784);
or UO_72 (O_72,N_24456,N_24718);
nand UO_73 (O_73,N_24618,N_22716);
nor UO_74 (O_74,N_22549,N_23636);
nand UO_75 (O_75,N_23910,N_22623);
and UO_76 (O_76,N_24570,N_22937);
or UO_77 (O_77,N_24272,N_23356);
and UO_78 (O_78,N_23795,N_24725);
nand UO_79 (O_79,N_23179,N_22869);
or UO_80 (O_80,N_24507,N_23242);
xor UO_81 (O_81,N_23430,N_24174);
nor UO_82 (O_82,N_23294,N_22628);
and UO_83 (O_83,N_24015,N_23661);
and UO_84 (O_84,N_23452,N_23818);
nand UO_85 (O_85,N_23271,N_24971);
or UO_86 (O_86,N_24081,N_24894);
and UO_87 (O_87,N_23813,N_24829);
nor UO_88 (O_88,N_24391,N_24311);
or UO_89 (O_89,N_22942,N_24482);
nor UO_90 (O_90,N_24468,N_24841);
or UO_91 (O_91,N_23653,N_23302);
and UO_92 (O_92,N_24158,N_23100);
nand UO_93 (O_93,N_22604,N_24382);
and UO_94 (O_94,N_23687,N_24908);
nand UO_95 (O_95,N_24435,N_23996);
or UO_96 (O_96,N_23956,N_23536);
nand UO_97 (O_97,N_24063,N_24436);
xnor UO_98 (O_98,N_23638,N_23730);
nor UO_99 (O_99,N_22903,N_23151);
and UO_100 (O_100,N_24432,N_23843);
and UO_101 (O_101,N_24344,N_24668);
and UO_102 (O_102,N_24910,N_24790);
or UO_103 (O_103,N_24975,N_23615);
nand UO_104 (O_104,N_22899,N_22779);
nor UO_105 (O_105,N_23906,N_24912);
xor UO_106 (O_106,N_22652,N_24497);
xor UO_107 (O_107,N_22809,N_24598);
xor UO_108 (O_108,N_23226,N_23697);
xor UO_109 (O_109,N_23559,N_24815);
and UO_110 (O_110,N_23835,N_24651);
nor UO_111 (O_111,N_23396,N_23354);
or UO_112 (O_112,N_23923,N_24602);
nor UO_113 (O_113,N_24009,N_24306);
nor UO_114 (O_114,N_24698,N_24500);
or UO_115 (O_115,N_24249,N_22817);
xnor UO_116 (O_116,N_24574,N_24103);
nand UO_117 (O_117,N_23774,N_23889);
xor UO_118 (O_118,N_24810,N_23796);
nor UO_119 (O_119,N_24412,N_24526);
nand UO_120 (O_120,N_22653,N_24275);
nand UO_121 (O_121,N_24111,N_24543);
xor UO_122 (O_122,N_23364,N_24449);
xnor UO_123 (O_123,N_23980,N_24068);
nor UO_124 (O_124,N_22971,N_23598);
and UO_125 (O_125,N_24733,N_24818);
nand UO_126 (O_126,N_23096,N_23408);
or UO_127 (O_127,N_22944,N_24771);
and UO_128 (O_128,N_23095,N_22760);
or UO_129 (O_129,N_23454,N_23917);
or UO_130 (O_130,N_24162,N_23051);
nand UO_131 (O_131,N_23891,N_24866);
or UO_132 (O_132,N_24367,N_22725);
nand UO_133 (O_133,N_23718,N_22742);
and UO_134 (O_134,N_23554,N_22929);
nand UO_135 (O_135,N_24268,N_22706);
nand UO_136 (O_136,N_24914,N_24924);
and UO_137 (O_137,N_24965,N_24506);
xor UO_138 (O_138,N_23210,N_24529);
nor UO_139 (O_139,N_23899,N_23264);
and UO_140 (O_140,N_24680,N_22601);
and UO_141 (O_141,N_22861,N_22925);
or UO_142 (O_142,N_23862,N_23021);
nor UO_143 (O_143,N_24764,N_23658);
nor UO_144 (O_144,N_24206,N_24514);
or UO_145 (O_145,N_24872,N_24699);
nor UO_146 (O_146,N_24294,N_23954);
or UO_147 (O_147,N_22849,N_24090);
or UO_148 (O_148,N_24259,N_24026);
xnor UO_149 (O_149,N_23513,N_22786);
nand UO_150 (O_150,N_23789,N_23883);
and UO_151 (O_151,N_23147,N_23714);
nand UO_152 (O_152,N_23875,N_22660);
or UO_153 (O_153,N_22647,N_24587);
and UO_154 (O_154,N_22898,N_22693);
nor UO_155 (O_155,N_23004,N_22514);
nor UO_156 (O_156,N_24134,N_24011);
xnor UO_157 (O_157,N_23245,N_24010);
xor UO_158 (O_158,N_22738,N_23237);
nor UO_159 (O_159,N_22666,N_24984);
and UO_160 (O_160,N_23394,N_23043);
nand UO_161 (O_161,N_22758,N_22854);
nor UO_162 (O_162,N_24321,N_24731);
xnor UO_163 (O_163,N_24339,N_22682);
nor UO_164 (O_164,N_23366,N_22677);
nor UO_165 (O_165,N_24440,N_24280);
and UO_166 (O_166,N_23908,N_24614);
nor UO_167 (O_167,N_22941,N_22713);
or UO_168 (O_168,N_24051,N_24697);
xnor UO_169 (O_169,N_24551,N_23558);
or UO_170 (O_170,N_24235,N_23710);
nand UO_171 (O_171,N_23553,N_23539);
and UO_172 (O_172,N_24018,N_23083);
and UO_173 (O_173,N_24461,N_22909);
xor UO_174 (O_174,N_24610,N_23463);
nor UO_175 (O_175,N_24003,N_23001);
and UO_176 (O_176,N_23876,N_22516);
xor UO_177 (O_177,N_24628,N_23416);
and UO_178 (O_178,N_23864,N_24776);
xnor UO_179 (O_179,N_24428,N_23543);
or UO_180 (O_180,N_23298,N_24159);
nor UO_181 (O_181,N_23628,N_23249);
and UO_182 (O_182,N_24365,N_24967);
or UO_183 (O_183,N_23017,N_23892);
nand UO_184 (O_184,N_24851,N_24336);
and UO_185 (O_185,N_22881,N_22954);
or UO_186 (O_186,N_23252,N_24004);
or UO_187 (O_187,N_24524,N_24871);
and UO_188 (O_188,N_22818,N_24149);
xor UO_189 (O_189,N_24980,N_24139);
xor UO_190 (O_190,N_23235,N_23530);
or UO_191 (O_191,N_24288,N_24190);
xor UO_192 (O_192,N_24549,N_23717);
nand UO_193 (O_193,N_24295,N_24330);
and UO_194 (O_194,N_24166,N_24438);
and UO_195 (O_195,N_23832,N_24744);
and UO_196 (O_196,N_22530,N_22676);
nand UO_197 (O_197,N_24545,N_24209);
nand UO_198 (O_198,N_24404,N_22748);
or UO_199 (O_199,N_23500,N_23120);
nand UO_200 (O_200,N_23678,N_22730);
xor UO_201 (O_201,N_23517,N_23392);
nor UO_202 (O_202,N_24147,N_24510);
or UO_203 (O_203,N_22871,N_24244);
nor UO_204 (O_204,N_22741,N_23327);
xnor UO_205 (O_205,N_23878,N_23750);
nand UO_206 (O_206,N_24012,N_22625);
or UO_207 (O_207,N_23672,N_23594);
or UO_208 (O_208,N_22593,N_24320);
xnor UO_209 (O_209,N_24183,N_24070);
xor UO_210 (O_210,N_23372,N_23116);
or UO_211 (O_211,N_24476,N_23675);
nor UO_212 (O_212,N_24993,N_23005);
or UO_213 (O_213,N_23531,N_23597);
or UO_214 (O_214,N_24552,N_23674);
nor UO_215 (O_215,N_23960,N_24937);
nand UO_216 (O_216,N_22680,N_23206);
nand UO_217 (O_217,N_24769,N_24932);
nor UO_218 (O_218,N_23321,N_24740);
nor UO_219 (O_219,N_24297,N_23097);
nand UO_220 (O_220,N_23900,N_23184);
nand UO_221 (O_221,N_22559,N_23305);
or UO_222 (O_222,N_23549,N_24243);
and UO_223 (O_223,N_24944,N_23039);
or UO_224 (O_224,N_23494,N_24966);
or UO_225 (O_225,N_23985,N_23177);
and UO_226 (O_226,N_23007,N_24172);
nand UO_227 (O_227,N_23625,N_24114);
and UO_228 (O_228,N_24487,N_22695);
or UO_229 (O_229,N_24493,N_23113);
nand UO_230 (O_230,N_23324,N_23379);
and UO_231 (O_231,N_23309,N_24623);
and UO_232 (O_232,N_23312,N_22597);
nand UO_233 (O_233,N_22502,N_24033);
nor UO_234 (O_234,N_22931,N_22936);
nor UO_235 (O_235,N_24751,N_22627);
nor UO_236 (O_236,N_22651,N_23865);
and UO_237 (O_237,N_23180,N_24176);
or UO_238 (O_238,N_24566,N_23257);
xor UO_239 (O_239,N_22997,N_23018);
nor UO_240 (O_240,N_22568,N_23991);
and UO_241 (O_241,N_23404,N_23150);
nor UO_242 (O_242,N_24092,N_23616);
or UO_243 (O_243,N_24671,N_23681);
or UO_244 (O_244,N_22875,N_23711);
xor UO_245 (O_245,N_24200,N_22777);
and UO_246 (O_246,N_22823,N_24027);
nor UO_247 (O_247,N_24694,N_23243);
or UO_248 (O_248,N_24054,N_22736);
nor UO_249 (O_249,N_22787,N_22639);
and UO_250 (O_250,N_23526,N_23871);
nand UO_251 (O_251,N_24153,N_24126);
nor UO_252 (O_252,N_22643,N_24262);
nor UO_253 (O_253,N_24416,N_24409);
or UO_254 (O_254,N_23125,N_24640);
nor UO_255 (O_255,N_23199,N_23939);
nand UO_256 (O_256,N_23694,N_23193);
nand UO_257 (O_257,N_23516,N_24379);
nand UO_258 (O_258,N_23212,N_23350);
and UO_259 (O_259,N_23152,N_23262);
nor UO_260 (O_260,N_23325,N_23501);
xor UO_261 (O_261,N_23734,N_24022);
and UO_262 (O_262,N_23916,N_23407);
nand UO_263 (O_263,N_23968,N_23927);
nand UO_264 (O_264,N_22681,N_24555);
nor UO_265 (O_265,N_23399,N_23617);
nor UO_266 (O_266,N_23427,N_23439);
nor UO_267 (O_267,N_23093,N_23304);
nor UO_268 (O_268,N_24977,N_24471);
or UO_269 (O_269,N_22719,N_22782);
nor UO_270 (O_270,N_22511,N_24044);
or UO_271 (O_271,N_24858,N_23168);
and UO_272 (O_272,N_24741,N_23491);
nand UO_273 (O_273,N_23291,N_24078);
nand UO_274 (O_274,N_22995,N_23112);
or UO_275 (O_275,N_23374,N_22607);
nor UO_276 (O_276,N_22634,N_24028);
or UO_277 (O_277,N_22833,N_23592);
or UO_278 (O_278,N_23902,N_23907);
or UO_279 (O_279,N_23317,N_23849);
xor UO_280 (O_280,N_23316,N_23942);
or UO_281 (O_281,N_22655,N_23745);
and UO_282 (O_282,N_23601,N_22862);
or UO_283 (O_283,N_23190,N_23082);
nand UO_284 (O_284,N_23753,N_24654);
and UO_285 (O_285,N_24855,N_24323);
or UO_286 (O_286,N_24040,N_23713);
nand UO_287 (O_287,N_23708,N_24304);
or UO_288 (O_288,N_24904,N_23014);
and UO_289 (O_289,N_23920,N_23783);
nor UO_290 (O_290,N_23510,N_23401);
or UO_291 (O_291,N_24319,N_23873);
nand UO_292 (O_292,N_24141,N_24036);
xor UO_293 (O_293,N_24783,N_22709);
or UO_294 (O_294,N_23512,N_22856);
nor UO_295 (O_295,N_22829,N_24913);
and UO_296 (O_296,N_23128,N_23192);
and UO_297 (O_297,N_22554,N_22866);
and UO_298 (O_298,N_24861,N_23341);
xnor UO_299 (O_299,N_23369,N_24477);
or UO_300 (O_300,N_22923,N_23640);
xor UO_301 (O_301,N_23222,N_23857);
or UO_302 (O_302,N_24341,N_22900);
xor UO_303 (O_303,N_23820,N_23664);
nand UO_304 (O_304,N_24223,N_22541);
nor UO_305 (O_305,N_24059,N_23062);
xor UO_306 (O_306,N_23445,N_24948);
nor UO_307 (O_307,N_24720,N_22814);
nor UO_308 (O_308,N_24997,N_23729);
xnor UO_309 (O_309,N_23848,N_22707);
or UO_310 (O_310,N_24825,N_23975);
and UO_311 (O_311,N_24348,N_23025);
nor UO_312 (O_312,N_23138,N_24509);
xnor UO_313 (O_313,N_24021,N_22588);
nand UO_314 (O_314,N_24934,N_22671);
nand UO_315 (O_315,N_23461,N_24363);
nand UO_316 (O_316,N_24228,N_23555);
and UO_317 (O_317,N_24260,N_23802);
xor UO_318 (O_318,N_23397,N_23576);
xor UO_319 (O_319,N_24531,N_23898);
nor UO_320 (O_320,N_24658,N_24122);
or UO_321 (O_321,N_23952,N_23108);
nor UO_322 (O_322,N_24263,N_24931);
nor UO_323 (O_323,N_23738,N_22662);
nand UO_324 (O_324,N_23869,N_22512);
or UO_325 (O_325,N_23219,N_23578);
and UO_326 (O_326,N_24096,N_22689);
nor UO_327 (O_327,N_24098,N_23685);
and UO_328 (O_328,N_24105,N_23178);
or UO_329 (O_329,N_23599,N_22921);
nor UO_330 (O_330,N_23080,N_22828);
and UO_331 (O_331,N_24737,N_22522);
nand UO_332 (O_332,N_24384,N_23903);
and UO_333 (O_333,N_23476,N_24433);
or UO_334 (O_334,N_23066,N_22976);
xor UO_335 (O_335,N_24253,N_24580);
nand UO_336 (O_336,N_24151,N_23444);
xor UO_337 (O_337,N_22617,N_22538);
nand UO_338 (O_338,N_24857,N_24723);
and UO_339 (O_339,N_22812,N_23989);
or UO_340 (O_340,N_23011,N_23153);
and UO_341 (O_341,N_22904,N_23921);
nand UO_342 (O_342,N_24662,N_24480);
and UO_343 (O_343,N_23238,N_22913);
nand UO_344 (O_344,N_24071,N_24921);
nor UO_345 (O_345,N_23825,N_23442);
or UO_346 (O_346,N_22972,N_24437);
or UO_347 (O_347,N_23816,N_24875);
nor UO_348 (O_348,N_24466,N_24030);
or UO_349 (O_349,N_22845,N_24298);
nand UO_350 (O_350,N_24544,N_24983);
nor UO_351 (O_351,N_23853,N_23131);
xor UO_352 (O_352,N_24095,N_23514);
and UO_353 (O_353,N_24761,N_23469);
xnor UO_354 (O_354,N_24760,N_23782);
and UO_355 (O_355,N_23425,N_24586);
and UO_356 (O_356,N_23498,N_24981);
nor UO_357 (O_357,N_23159,N_23218);
and UO_358 (O_358,N_23935,N_24085);
nand UO_359 (O_359,N_23326,N_23217);
nand UO_360 (O_360,N_24255,N_24862);
or UO_361 (O_361,N_24057,N_24406);
nor UO_362 (O_362,N_23197,N_23258);
xor UO_363 (O_363,N_22555,N_23301);
nor UO_364 (O_364,N_24191,N_24947);
nand UO_365 (O_365,N_24358,N_24901);
and UO_366 (O_366,N_23196,N_24985);
xor UO_367 (O_367,N_22963,N_24164);
nand UO_368 (O_368,N_23034,N_23807);
xnor UO_369 (O_369,N_24631,N_23544);
and UO_370 (O_370,N_23725,N_23641);
nand UO_371 (O_371,N_24375,N_22934);
and UO_372 (O_372,N_24584,N_24712);
and UO_373 (O_373,N_23142,N_24770);
nor UO_374 (O_374,N_22956,N_22551);
and UO_375 (O_375,N_22629,N_23583);
and UO_376 (O_376,N_23763,N_24778);
or UO_377 (O_377,N_24882,N_22831);
nand UO_378 (O_378,N_22768,N_22859);
xor UO_379 (O_379,N_24951,N_23297);
xnor UO_380 (O_380,N_24329,N_23272);
and UO_381 (O_381,N_23135,N_23457);
nor UO_382 (O_382,N_23183,N_23817);
and UO_383 (O_383,N_24806,N_22910);
xnor UO_384 (O_384,N_24831,N_24709);
or UO_385 (O_385,N_24665,N_22642);
xnor UO_386 (O_386,N_23505,N_24032);
nor UO_387 (O_387,N_22860,N_22970);
nor UO_388 (O_388,N_23788,N_22883);
and UO_389 (O_389,N_23969,N_24808);
nor UO_390 (O_390,N_23146,N_23044);
nand UO_391 (O_391,N_22844,N_24067);
nand UO_392 (O_392,N_24061,N_24113);
xnor UO_393 (O_393,N_23114,N_23518);
xor UO_394 (O_394,N_24881,N_23768);
or UO_395 (O_395,N_22714,N_22864);
xnor UO_396 (O_396,N_22975,N_23339);
nor UO_397 (O_397,N_23981,N_24474);
and UO_398 (O_398,N_24360,N_24335);
or UO_399 (O_399,N_24419,N_23458);
or UO_400 (O_400,N_23581,N_23124);
or UO_401 (O_401,N_23524,N_23023);
nor UO_402 (O_402,N_23451,N_23837);
and UO_403 (O_403,N_23269,N_22544);
and UO_404 (O_404,N_24705,N_23419);
nor UO_405 (O_405,N_22838,N_23705);
nor UO_406 (O_406,N_22774,N_24516);
and UO_407 (O_407,N_22945,N_24728);
nor UO_408 (O_408,N_23293,N_24923);
nor UO_409 (O_409,N_24603,N_23937);
nand UO_410 (O_410,N_22657,N_23680);
xor UO_411 (O_411,N_23926,N_23215);
or UO_412 (O_412,N_23570,N_23983);
xnor UO_413 (O_413,N_23683,N_24638);
or UO_414 (O_414,N_24883,N_23446);
nand UO_415 (O_415,N_23277,N_24772);
or UO_416 (O_416,N_24314,N_24874);
or UO_417 (O_417,N_22990,N_23701);
xnor UO_418 (O_418,N_22508,N_23970);
nor UO_419 (O_419,N_23794,N_23965);
nand UO_420 (O_420,N_24650,N_23154);
xor UO_421 (O_421,N_24792,N_23776);
nand UO_422 (O_422,N_23090,N_24635);
nand UO_423 (O_423,N_23744,N_24383);
nor UO_424 (O_424,N_24830,N_24564);
xnor UO_425 (O_425,N_24371,N_23588);
nor UO_426 (O_426,N_24605,N_23362);
xnor UO_427 (O_427,N_23977,N_22775);
nand UO_428 (O_428,N_22816,N_23976);
or UO_429 (O_429,N_23126,N_24525);
nand UO_430 (O_430,N_23585,N_24014);
nand UO_431 (O_431,N_23803,N_22843);
nor UO_432 (O_432,N_22535,N_22743);
nand UO_433 (O_433,N_23929,N_23208);
nor UO_434 (O_434,N_24613,N_24848);
xnor UO_435 (O_435,N_24667,N_23723);
xor UO_436 (O_436,N_24124,N_22801);
or UO_437 (O_437,N_22744,N_24522);
nand UO_438 (O_438,N_23122,N_24499);
nor UO_439 (O_439,N_22791,N_23241);
nor UO_440 (O_440,N_24047,N_22576);
nand UO_441 (O_441,N_23812,N_24748);
or UO_442 (O_442,N_24743,N_22594);
nand UO_443 (O_443,N_23614,N_23239);
or UO_444 (O_444,N_22747,N_24809);
nand UO_445 (O_445,N_24077,N_22612);
xnor UO_446 (O_446,N_24802,N_24788);
xor UO_447 (O_447,N_23659,N_24805);
nor UO_448 (O_448,N_22578,N_24916);
xnor UO_449 (O_449,N_22581,N_23938);
or UO_450 (O_450,N_23185,N_22586);
or UO_451 (O_451,N_23338,N_24824);
or UO_452 (O_452,N_23391,N_23345);
and UO_453 (O_453,N_24089,N_24094);
nor UO_454 (O_454,N_23541,N_24583);
xor UO_455 (O_455,N_24957,N_24178);
nand UO_456 (O_456,N_23104,N_23978);
nand UO_457 (O_457,N_24624,N_23329);
nand UO_458 (O_458,N_22811,N_23055);
and UO_459 (O_459,N_23897,N_23609);
or UO_460 (O_460,N_23663,N_24821);
or UO_461 (O_461,N_23565,N_24491);
xnor UO_462 (O_462,N_24989,N_23884);
or UO_463 (O_463,N_24612,N_24042);
and UO_464 (O_464,N_24424,N_23024);
nor UO_465 (O_465,N_23236,N_23944);
nand UO_466 (O_466,N_24579,N_22691);
nand UO_467 (O_467,N_24119,N_24445);
nor UO_468 (O_468,N_24565,N_22606);
xnor UO_469 (O_469,N_22723,N_23281);
nor UO_470 (O_470,N_24053,N_23911);
xnor UO_471 (O_471,N_23191,N_23751);
and UO_472 (O_472,N_24987,N_23048);
nor UO_473 (O_473,N_23176,N_24834);
xor UO_474 (O_474,N_23562,N_24394);
xor UO_475 (O_475,N_22754,N_24247);
or UO_476 (O_476,N_22729,N_24961);
xor UO_477 (O_477,N_22509,N_24893);
xnor UO_478 (O_478,N_23384,N_22579);
or UO_479 (O_479,N_23230,N_22901);
nor UO_480 (O_480,N_23194,N_24896);
nor UO_481 (O_481,N_24535,N_24305);
nor UO_482 (O_482,N_23342,N_23933);
or UO_483 (O_483,N_23785,N_23901);
xnor UO_484 (O_484,N_23564,N_24735);
and UO_485 (O_485,N_23644,N_23047);
nor UO_486 (O_486,N_23145,N_24611);
nand UO_487 (O_487,N_23880,N_23480);
nand UO_488 (O_488,N_24142,N_24481);
and UO_489 (O_489,N_23520,N_23612);
or UO_490 (O_490,N_24239,N_24843);
nand UO_491 (O_491,N_24179,N_23462);
xnor UO_492 (O_492,N_23618,N_24050);
xor UO_493 (O_493,N_24575,N_24282);
nand UO_494 (O_494,N_24657,N_24316);
nand UO_495 (O_495,N_22745,N_23861);
nor UO_496 (O_496,N_24828,N_24350);
xnor UO_497 (O_497,N_24541,N_22531);
nand UO_498 (O_498,N_23662,N_24659);
or UO_499 (O_499,N_22826,N_22885);
nand UO_500 (O_500,N_24447,N_23027);
xnor UO_501 (O_501,N_22546,N_23448);
or UO_502 (O_502,N_24726,N_23696);
and UO_503 (O_503,N_23732,N_23829);
nand UO_504 (O_504,N_23266,N_23834);
nand UO_505 (O_505,N_22722,N_23706);
and UO_506 (O_506,N_24269,N_24216);
nor UO_507 (O_507,N_23268,N_24257);
nand UO_508 (O_508,N_23308,N_24800);
nand UO_509 (O_509,N_23421,N_23037);
xnor UO_510 (O_510,N_23456,N_23821);
and UO_511 (O_511,N_23695,N_24368);
xor UO_512 (O_512,N_23885,N_24261);
or UO_513 (O_513,N_24569,N_24711);
and UO_514 (O_514,N_22765,N_24513);
xnor UO_515 (O_515,N_24146,N_22839);
xor UO_516 (O_516,N_23997,N_23117);
nor UO_517 (O_517,N_24642,N_22840);
nor UO_518 (O_518,N_23879,N_23200);
xor UO_519 (O_519,N_23797,N_24121);
nor UO_520 (O_520,N_22896,N_24212);
and UO_521 (O_521,N_24006,N_22592);
nand UO_522 (O_522,N_24986,N_24669);
nor UO_523 (O_523,N_24519,N_22892);
and UO_524 (O_524,N_23166,N_23072);
nand UO_525 (O_525,N_22939,N_24230);
nand UO_526 (O_526,N_23351,N_24300);
and UO_527 (O_527,N_23622,N_22922);
and UO_528 (O_528,N_24465,N_23627);
and UO_529 (O_529,N_23158,N_24707);
xnor UO_530 (O_530,N_23856,N_23387);
nand UO_531 (O_531,N_24045,N_24585);
nand UO_532 (O_532,N_22649,N_23233);
nor UO_533 (O_533,N_24643,N_23987);
xnor UO_534 (O_534,N_22943,N_24264);
and UO_535 (O_535,N_24945,N_24462);
and UO_536 (O_536,N_23743,N_22542);
xor UO_537 (O_537,N_24530,N_24289);
or UO_538 (O_538,N_24639,N_23042);
nand UO_539 (O_539,N_23483,N_24877);
and UO_540 (O_540,N_23525,N_24104);
nand UO_541 (O_541,N_24303,N_23503);
nor UO_542 (O_542,N_24738,N_22577);
and UO_543 (O_543,N_24351,N_22973);
or UO_544 (O_544,N_23134,N_23836);
nand UO_545 (O_545,N_24154,N_23671);
nand UO_546 (O_546,N_24418,N_23443);
xnor UO_547 (O_547,N_24083,N_24074);
nor UO_548 (O_548,N_22905,N_24198);
nand UO_549 (O_549,N_23056,N_23582);
nand UO_550 (O_550,N_24352,N_24889);
or UO_551 (O_551,N_23250,N_22558);
xor UO_552 (O_552,N_24789,N_24689);
or UO_553 (O_553,N_24779,N_22947);
or UO_554 (O_554,N_22533,N_24349);
or UO_555 (O_555,N_24992,N_24102);
nor UO_556 (O_556,N_23846,N_23566);
and UO_557 (O_557,N_24414,N_22857);
nor UO_558 (O_558,N_24187,N_23563);
nand UO_559 (O_559,N_24137,N_23914);
or UO_560 (O_560,N_23950,N_22969);
or UO_561 (O_561,N_23495,N_23635);
xnor UO_562 (O_562,N_24256,N_24762);
and UO_563 (O_563,N_24736,N_23781);
and UO_564 (O_564,N_24508,N_23079);
or UO_565 (O_565,N_22705,N_23299);
nand UO_566 (O_566,N_23728,N_23775);
or UO_567 (O_567,N_24700,N_24803);
and UO_568 (O_568,N_24488,N_24854);
and UO_569 (O_569,N_22992,N_23913);
or UO_570 (O_570,N_24540,N_24169);
nand UO_571 (O_571,N_24326,N_24859);
xnor UO_572 (O_572,N_23793,N_23943);
nor UO_573 (O_573,N_23111,N_24559);
nor UO_574 (O_574,N_24150,N_24286);
nand UO_575 (O_575,N_22622,N_24274);
nand UO_576 (O_576,N_23088,N_23381);
nand UO_577 (O_577,N_23932,N_24080);
or UO_578 (O_578,N_23646,N_24998);
xnor UO_579 (O_579,N_24281,N_22813);
and UO_580 (O_580,N_24648,N_23839);
xor UO_581 (O_581,N_24308,N_24390);
nand UO_582 (O_582,N_22590,N_23465);
nand UO_583 (O_583,N_23253,N_23267);
nand UO_584 (O_584,N_24956,N_23058);
or UO_585 (O_585,N_22763,N_23343);
nand UO_586 (O_586,N_23752,N_24988);
nor UO_587 (O_587,N_22635,N_23528);
xnor UO_588 (O_588,N_22600,N_22526);
xor UO_589 (O_589,N_23984,N_24767);
nand UO_590 (O_590,N_24160,N_24891);
and UO_591 (O_591,N_24537,N_22987);
or UO_592 (O_592,N_23357,N_23893);
or UO_593 (O_593,N_24785,N_22886);
or UO_594 (O_594,N_23827,N_22895);
and UO_595 (O_595,N_24777,N_22888);
and UO_596 (O_596,N_24227,N_23521);
nor UO_597 (O_597,N_23808,N_22670);
or UO_598 (O_598,N_24696,N_22890);
xnor UO_599 (O_599,N_24679,N_24926);
nand UO_600 (O_600,N_24454,N_22983);
xnor UO_601 (O_601,N_24116,N_24632);
and UO_602 (O_602,N_22851,N_24222);
nor UO_603 (O_603,N_23604,N_24224);
nand UO_604 (O_604,N_23067,N_22686);
nand UO_605 (O_605,N_24332,N_24072);
nand UO_606 (O_606,N_24899,N_22548);
and UO_607 (O_607,N_24393,N_23561);
nor UO_608 (O_608,N_22636,N_24678);
nor UO_609 (O_609,N_22683,N_24849);
nand UO_610 (O_610,N_24458,N_24746);
xnor UO_611 (O_611,N_23248,N_23596);
nand UO_612 (O_612,N_24627,N_23279);
nand UO_613 (O_613,N_23930,N_22615);
nor UO_614 (O_614,N_24043,N_24086);
and UO_615 (O_615,N_23886,N_23414);
or UO_616 (O_616,N_24266,N_24220);
xor UO_617 (O_617,N_23497,N_22726);
nor UO_618 (O_618,N_23519,N_24836);
nand UO_619 (O_619,N_24389,N_22620);
nor UO_620 (O_620,N_24396,N_23998);
xor UO_621 (O_621,N_22953,N_23633);
and UO_622 (O_622,N_22986,N_23009);
nor UO_623 (O_623,N_24429,N_24653);
or UO_624 (O_624,N_24346,N_24101);
xnor UO_625 (O_625,N_24182,N_22685);
nand UO_626 (O_626,N_23670,N_22834);
and UO_627 (O_627,N_24546,N_24608);
nor UO_628 (O_628,N_24817,N_22661);
nor UO_629 (O_629,N_22610,N_23511);
and UO_630 (O_630,N_23136,N_23804);
nor UO_631 (O_631,N_24443,N_23852);
or UO_632 (O_632,N_23974,N_23721);
nor UO_633 (O_633,N_23668,N_24372);
and UO_634 (O_634,N_23468,N_24241);
xnor UO_635 (O_635,N_22560,N_23679);
and UO_636 (O_636,N_24181,N_23105);
or UO_637 (O_637,N_22659,N_23809);
nor UO_638 (O_638,N_22868,N_24234);
nor UO_639 (O_639,N_22699,N_22794);
nand UO_640 (O_640,N_23484,N_23580);
and UO_641 (O_641,N_24100,N_24380);
xnor UO_642 (O_642,N_23737,N_23144);
or UO_643 (O_643,N_23995,N_23420);
and UO_644 (O_644,N_23283,N_23621);
nand UO_645 (O_645,N_22880,N_24943);
and UO_646 (O_646,N_22561,N_23571);
and UO_647 (O_647,N_24333,N_24338);
nor UO_648 (O_648,N_24568,N_24278);
nor UO_649 (O_649,N_22556,N_22752);
or UO_650 (O_650,N_22795,N_23888);
and UO_651 (O_651,N_23866,N_23493);
xor UO_652 (O_652,N_23089,N_22500);
nand UO_653 (O_653,N_24604,N_23590);
nor UO_654 (O_654,N_23863,N_24813);
or UO_655 (O_655,N_23755,N_24976);
nand UO_656 (O_656,N_24719,N_24536);
or UO_657 (O_657,N_24727,N_24732);
or UO_658 (O_658,N_24754,N_24502);
xnor UO_659 (O_659,N_23263,N_24617);
nand UO_660 (O_660,N_24097,N_22751);
xor UO_661 (O_661,N_23799,N_23211);
nand UO_662 (O_662,N_23091,N_24884);
or UO_663 (O_663,N_24959,N_23322);
nand UO_664 (O_664,N_24964,N_23478);
or UO_665 (O_665,N_23967,N_22529);
and UO_666 (O_666,N_24277,N_23361);
nor UO_667 (O_667,N_23972,N_23038);
nor UO_668 (O_668,N_23205,N_23490);
nand UO_669 (O_669,N_23447,N_24933);
and UO_670 (O_670,N_24629,N_23650);
and UO_671 (O_671,N_22720,N_24990);
and UO_672 (O_672,N_24318,N_24796);
nor UO_673 (O_673,N_23805,N_23572);
and UO_674 (O_674,N_23085,N_24799);
xnor UO_675 (O_675,N_23141,N_23216);
nand UO_676 (O_676,N_24794,N_23669);
xor UO_677 (O_677,N_24717,N_22988);
or UO_678 (O_678,N_24523,N_24165);
nand UO_679 (O_679,N_23964,N_23819);
and UO_680 (O_680,N_23260,N_24129);
nor UO_681 (O_681,N_23377,N_24844);
or UO_682 (O_682,N_24215,N_22879);
xor UO_683 (O_683,N_24749,N_23121);
or UO_684 (O_684,N_23426,N_22528);
xor UO_685 (O_685,N_22948,N_24708);
nor UO_686 (O_686,N_23754,N_23422);
nand UO_687 (O_687,N_24692,N_23527);
nand UO_688 (O_688,N_23380,N_24345);
nor UO_689 (O_689,N_23393,N_24619);
nand UO_690 (O_690,N_24902,N_23823);
nand UO_691 (O_691,N_23736,N_24293);
xnor UO_692 (O_692,N_23546,N_23660);
xor UO_693 (O_693,N_23847,N_23071);
nand UO_694 (O_694,N_24684,N_23052);
xor UO_695 (O_695,N_23240,N_22547);
and UO_696 (O_696,N_22762,N_24807);
or UO_697 (O_697,N_23406,N_23560);
nand UO_698 (O_698,N_23949,N_22598);
nor UO_699 (O_699,N_24448,N_22757);
or UO_700 (O_700,N_24685,N_23174);
xor UO_701 (O_701,N_24974,N_23961);
nor UO_702 (O_702,N_23896,N_23731);
and UO_703 (O_703,N_24145,N_22573);
xnor UO_704 (O_704,N_24217,N_24173);
nor UO_705 (O_705,N_24343,N_22805);
xnor UO_706 (O_706,N_22718,N_24539);
xor UO_707 (O_707,N_23157,N_24528);
and UO_708 (O_708,N_24473,N_23682);
or UO_709 (O_709,N_22701,N_23081);
nor UO_710 (O_710,N_24691,N_24402);
xor UO_711 (O_711,N_24238,N_24279);
nor UO_712 (O_712,N_22756,N_22842);
nor UO_713 (O_713,N_23854,N_23344);
nor UO_714 (O_714,N_22806,N_23791);
xnor UO_715 (O_715,N_23398,N_24052);
or UO_716 (O_716,N_22940,N_23373);
and UO_717 (O_717,N_22915,N_22979);
nor UO_718 (O_718,N_23137,N_23909);
nor UO_719 (O_719,N_22991,N_24939);
nand UO_720 (O_720,N_22584,N_23244);
and UO_721 (O_721,N_23905,N_23912);
xor UO_722 (O_722,N_23684,N_22638);
and UO_723 (O_723,N_23784,N_24475);
nand UO_724 (O_724,N_24819,N_24327);
nor UO_725 (O_725,N_23538,N_24676);
or UO_726 (O_726,N_23704,N_23534);
xor UO_727 (O_727,N_22687,N_23225);
xor UO_728 (O_728,N_23485,N_22599);
and UO_729 (O_729,N_22873,N_22674);
and UO_730 (O_730,N_24533,N_24787);
nand UO_731 (O_731,N_24716,N_22872);
and UO_732 (O_732,N_23285,N_23547);
xnor UO_733 (O_733,N_24837,N_22836);
nand UO_734 (O_734,N_24271,N_23296);
nor UO_735 (O_735,N_23798,N_24398);
nand UO_736 (O_736,N_24309,N_22766);
nor UO_737 (O_737,N_24532,N_23221);
nand UO_738 (O_738,N_24576,N_22637);
nand UO_739 (O_739,N_22632,N_23792);
or UO_740 (O_740,N_22648,N_24571);
or UO_741 (O_741,N_24686,N_23855);
or UO_742 (O_742,N_24804,N_24869);
nand UO_743 (O_743,N_22755,N_24184);
nand UO_744 (O_744,N_23022,N_24864);
or UO_745 (O_745,N_24838,N_23365);
and UO_746 (O_746,N_23579,N_24747);
and UO_747 (O_747,N_24225,N_22968);
nor UO_748 (O_748,N_24582,N_24860);
nor UO_749 (O_749,N_22999,N_23337);
and UO_750 (O_750,N_22621,N_23195);
xnor UO_751 (O_751,N_23504,N_22534);
and UO_752 (O_752,N_23477,N_23274);
nor UO_753 (O_753,N_23947,N_23602);
xnor UO_754 (O_754,N_22710,N_22804);
and UO_755 (O_755,N_22785,N_23639);
and UO_756 (O_756,N_24550,N_22717);
nor UO_757 (O_757,N_23306,N_24503);
or UO_758 (O_758,N_24324,N_22630);
and UO_759 (O_759,N_24088,N_24845);
and UO_760 (O_760,N_23428,N_23620);
or UO_761 (O_761,N_22589,N_22552);
xnor UO_762 (O_762,N_24763,N_24463);
nor UO_763 (O_763,N_22769,N_22863);
and UO_764 (O_764,N_22767,N_23400);
nand UO_765 (O_765,N_23739,N_23403);
nand UO_766 (O_766,N_23002,N_24202);
or UO_767 (O_767,N_22870,N_24759);
xor UO_768 (O_768,N_22735,N_22626);
or UO_769 (O_769,N_23487,N_24195);
or UO_770 (O_770,N_23720,N_24865);
nand UO_771 (O_771,N_24558,N_22602);
nor UO_772 (O_772,N_24739,N_23655);
and UO_773 (O_773,N_23320,N_22704);
xnor UO_774 (O_774,N_23319,N_24867);
nor UO_775 (O_775,N_22780,N_23787);
and UO_776 (O_776,N_24963,N_23676);
nor UO_777 (O_777,N_24521,N_24093);
nand UO_778 (O_778,N_23288,N_23273);
nand UO_779 (O_779,N_24594,N_23270);
nor UO_780 (O_780,N_24670,N_24325);
xor UO_781 (O_781,N_23756,N_24494);
xnor UO_782 (O_782,N_24213,N_22957);
nand UO_783 (O_783,N_24929,N_22800);
or UO_784 (O_784,N_23109,N_24464);
nand UO_785 (O_785,N_23552,N_24287);
and UO_786 (O_786,N_24556,N_24600);
and UO_787 (O_787,N_22708,N_22938);
nand UO_788 (O_788,N_24915,N_22668);
nor UO_789 (O_789,N_22536,N_23328);
xnor UO_790 (O_790,N_23719,N_22570);
and UO_791 (O_791,N_24373,N_24196);
or UO_792 (O_792,N_22789,N_23603);
nand UO_793 (O_793,N_24969,N_22613);
or UO_794 (O_794,N_23838,N_23348);
or UO_795 (O_795,N_24683,N_22678);
nand UO_796 (O_796,N_23375,N_22540);
or UO_797 (O_797,N_24016,N_23169);
or UO_798 (O_798,N_24087,N_23352);
nor UO_799 (O_799,N_22930,N_23189);
or UO_800 (O_800,N_24616,N_24577);
nand UO_801 (O_801,N_23261,N_22633);
nor UO_802 (O_802,N_23246,N_24470);
nand UO_803 (O_803,N_23076,N_23204);
or UO_804 (O_804,N_24826,N_22820);
xnor UO_805 (O_805,N_24405,N_22958);
and UO_806 (O_806,N_23060,N_24177);
nor UO_807 (O_807,N_23234,N_24722);
nor UO_808 (O_808,N_22852,N_24505);
nand UO_809 (O_809,N_23535,N_22650);
nor UO_810 (O_810,N_22619,N_22980);
and UO_811 (O_811,N_23030,N_22932);
nor UO_812 (O_812,N_24315,N_24958);
and UO_813 (O_813,N_24310,N_23915);
and UO_814 (O_814,N_23632,N_22525);
or UO_815 (O_815,N_23778,N_24408);
or UO_816 (O_816,N_23413,N_23313);
nand UO_817 (O_817,N_24978,N_24755);
nor UO_818 (O_818,N_23003,N_24660);
nor UO_819 (O_819,N_23496,N_23388);
nor UO_820 (O_820,N_24008,N_24750);
and UO_821 (O_821,N_24562,N_24636);
and UO_822 (O_822,N_23440,N_22848);
and UO_823 (O_823,N_23790,N_24907);
nor UO_824 (O_824,N_23690,N_23486);
nand UO_825 (O_825,N_23254,N_22609);
xnor UO_826 (O_826,N_22884,N_23600);
or UO_827 (O_827,N_24362,N_22537);
and UO_828 (O_828,N_23665,N_24439);
xnor UO_829 (O_829,N_22977,N_22702);
xnor UO_830 (O_830,N_22750,N_23464);
or UO_831 (O_831,N_24633,N_23858);
and UO_832 (O_832,N_22675,N_23904);
nand UO_833 (O_833,N_24548,N_24991);
nor UO_834 (O_834,N_24666,N_24900);
xnor UO_835 (O_835,N_23749,N_24768);
xnor UO_836 (O_836,N_23101,N_24251);
or UO_837 (O_837,N_22965,N_22961);
nor UO_838 (O_838,N_24125,N_24479);
xnor UO_839 (O_839,N_24041,N_24112);
and UO_840 (O_840,N_22572,N_24148);
and UO_841 (O_841,N_24240,N_22949);
or UO_842 (O_842,N_23033,N_23709);
and UO_843 (O_843,N_24017,N_22837);
nor UO_844 (O_844,N_23132,N_22867);
nor UO_845 (O_845,N_22911,N_23149);
nor UO_846 (O_846,N_22732,N_23438);
and UO_847 (O_847,N_24835,N_24811);
and UO_848 (O_848,N_23606,N_22821);
nand UO_849 (O_849,N_23231,N_23508);
and UO_850 (O_850,N_24942,N_24982);
xnor UO_851 (O_851,N_24688,N_22543);
xor UO_852 (O_852,N_23059,N_23368);
nor UO_853 (O_853,N_24784,N_24156);
xnor UO_854 (O_854,N_24695,N_24905);
and UO_855 (O_855,N_24781,N_24056);
and UO_856 (O_856,N_22565,N_23311);
xnor UO_857 (O_857,N_22761,N_24444);
or UO_858 (O_858,N_23143,N_24553);
nor UO_859 (O_859,N_23800,N_23573);
xor UO_860 (O_860,N_23762,N_23417);
xor UO_861 (O_861,N_23163,N_24450);
nor UO_862 (O_862,N_24968,N_24703);
nor UO_863 (O_863,N_23702,N_24180);
nor UO_864 (O_864,N_24203,N_24542);
xnor UO_865 (O_865,N_24927,N_23507);
nand UO_866 (O_866,N_23700,N_23973);
and UO_867 (O_867,N_24242,N_24385);
nand UO_868 (O_868,N_23441,N_23041);
and UO_869 (O_869,N_24538,N_22733);
and UO_870 (O_870,N_23133,N_24563);
and UO_871 (O_871,N_22656,N_22974);
nand UO_872 (O_872,N_23061,N_24208);
nor UO_873 (O_873,N_22778,N_24589);
xnor UO_874 (O_874,N_22790,N_24019);
nand UO_875 (O_875,N_24935,N_24399);
nor UO_876 (O_876,N_22964,N_24557);
and UO_877 (O_877,N_22587,N_22539);
nand UO_878 (O_878,N_22989,N_24037);
xor UO_879 (O_879,N_23489,N_23716);
and UO_880 (O_880,N_24928,N_23872);
or UO_881 (O_881,N_23874,N_23881);
or UO_882 (O_882,N_24400,N_24702);
xor UO_883 (O_883,N_22503,N_24742);
nand UO_884 (O_884,N_24211,N_22960);
xnor UO_885 (O_885,N_22505,N_24979);
nor UO_886 (O_886,N_24386,N_23651);
nand UO_887 (O_887,N_23488,N_24724);
or UO_888 (O_888,N_23586,N_24331);
xnor UO_889 (O_889,N_23963,N_23877);
nor UO_890 (O_890,N_24312,N_24229);
and UO_891 (O_891,N_24285,N_24138);
and UO_892 (O_892,N_23103,N_23280);
nor UO_893 (O_893,N_24823,N_22698);
xor UO_894 (O_894,N_23385,N_23050);
nor UO_895 (O_895,N_24024,N_24842);
nand UO_896 (O_896,N_23202,N_24001);
xor UO_897 (O_897,N_23411,N_23170);
and UO_898 (O_898,N_24420,N_23363);
xor UO_899 (O_899,N_24955,N_22672);
nor UO_900 (O_900,N_22616,N_23247);
and UO_901 (O_901,N_23953,N_23371);
xnor UO_902 (O_902,N_24591,N_24069);
or UO_903 (O_903,N_23346,N_24133);
or UO_904 (O_904,N_23637,N_23811);
nand UO_905 (O_905,N_23722,N_22764);
and UO_906 (O_906,N_23256,N_23332);
nor UO_907 (O_907,N_23649,N_23110);
nand UO_908 (O_908,N_23810,N_22569);
nor UO_909 (O_909,N_23429,N_23748);
nand UO_910 (O_910,N_23370,N_23314);
nor UO_911 (O_911,N_24606,N_22850);
and UO_912 (O_912,N_23691,N_23515);
nor UO_913 (O_913,N_23919,N_24107);
or UO_914 (O_914,N_24886,N_23181);
xnor UO_915 (O_915,N_23035,N_24451);
and UO_916 (O_916,N_23165,N_23626);
nor UO_917 (O_917,N_24547,N_24713);
nand UO_918 (O_918,N_24221,N_23127);
xor UO_919 (O_919,N_23654,N_23472);
nor UO_920 (O_920,N_23648,N_23040);
nor UO_921 (O_921,N_23951,N_22917);
nor UO_922 (O_922,N_24035,N_23223);
and UO_923 (O_923,N_23286,N_23276);
nand UO_924 (O_924,N_23334,N_24903);
nand UO_925 (O_925,N_24245,N_24283);
or UO_926 (O_926,N_22679,N_22696);
xnor UO_927 (O_927,N_23589,N_23766);
or UO_928 (O_928,N_22824,N_23801);
xor UO_929 (O_929,N_24411,N_22605);
nand UO_930 (O_930,N_23460,N_24058);
or UO_931 (O_931,N_23203,N_23207);
nor UO_932 (O_932,N_22566,N_23063);
or UO_933 (O_933,N_23735,N_23358);
xor UO_934 (O_934,N_23436,N_22721);
or UO_935 (O_935,N_23000,N_24322);
nor UO_936 (O_936,N_24890,N_24630);
or UO_937 (O_937,N_23053,N_24715);
xnor UO_938 (O_938,N_22993,N_23026);
nor UO_939 (O_939,N_22527,N_24607);
nand UO_940 (O_940,N_23015,N_23870);
nor UO_941 (O_941,N_23982,N_23814);
or UO_942 (O_942,N_23971,N_22697);
and UO_943 (O_943,N_23506,N_23540);
nand UO_944 (O_944,N_23431,N_24073);
or UO_945 (O_945,N_23376,N_22663);
nand UO_946 (O_946,N_22959,N_23948);
or UO_947 (O_947,N_23255,N_24188);
and UO_948 (O_948,N_23340,N_24876);
nand UO_949 (O_949,N_22966,N_22712);
or UO_950 (O_950,N_23070,N_23742);
and UO_951 (O_951,N_22822,N_24302);
and UO_952 (O_952,N_24403,N_24675);
nor UO_953 (O_953,N_24417,N_24560);
nor UO_954 (O_954,N_22553,N_23994);
or UO_955 (O_955,N_24573,N_23962);
nor UO_956 (O_956,N_24118,N_23733);
and UO_957 (O_957,N_24681,N_23459);
and UO_958 (O_958,N_24110,N_23529);
xnor UO_959 (O_959,N_24588,N_23251);
nor UO_960 (O_960,N_24392,N_22771);
nor UO_961 (O_961,N_22515,N_23850);
nor UO_962 (O_962,N_23424,N_23378);
xor UO_963 (O_963,N_24467,N_24189);
and UO_964 (O_964,N_22889,N_24140);
nor UO_965 (O_965,N_23209,N_23412);
or UO_966 (O_966,N_24721,N_24214);
or UO_967 (O_967,N_24284,N_23068);
xor UO_968 (O_968,N_22847,N_23064);
and UO_969 (O_969,N_23605,N_24290);
nor UO_970 (O_970,N_24850,N_24846);
or UO_971 (O_971,N_24431,N_22640);
and UO_972 (O_972,N_22740,N_22906);
nor UO_973 (O_973,N_24595,N_24127);
or UO_974 (O_974,N_23959,N_24395);
xor UO_975 (O_975,N_23642,N_23924);
xor UO_976 (O_976,N_23455,N_22783);
xnor UO_977 (O_977,N_22919,N_22727);
or UO_978 (O_978,N_23502,N_23130);
or UO_979 (O_979,N_23115,N_23140);
or UO_980 (O_980,N_24366,N_24397);
xor UO_981 (O_981,N_24258,N_24661);
xor UO_982 (O_982,N_24511,N_22518);
and UO_983 (O_983,N_23777,N_24109);
xor UO_984 (O_984,N_24441,N_23936);
nand UO_985 (O_985,N_22575,N_23747);
and UO_986 (O_986,N_23726,N_22501);
xor UO_987 (O_987,N_23523,N_22759);
nor UO_988 (O_988,N_24232,N_24960);
xnor UO_989 (O_989,N_24620,N_24002);
and UO_990 (O_990,N_24895,N_23008);
xnor UO_991 (O_991,N_24952,N_24922);
xor UO_992 (O_992,N_23432,N_24870);
xor UO_993 (O_993,N_24634,N_23992);
nor UO_994 (O_994,N_24641,N_23867);
or UO_995 (O_995,N_22924,N_24046);
or UO_996 (O_996,N_24425,N_24364);
or UO_997 (O_997,N_22952,N_24534);
nand UO_998 (O_998,N_24887,N_24897);
nand UO_999 (O_999,N_24136,N_24677);
and UO_1000 (O_1000,N_24936,N_24646);
xor UO_1001 (O_1001,N_24898,N_24376);
and UO_1002 (O_1002,N_23434,N_23645);
or UO_1003 (O_1003,N_24816,N_24204);
nand UO_1004 (O_1004,N_23467,N_23707);
nand UO_1005 (O_1005,N_23925,N_23290);
or UO_1006 (O_1006,N_23931,N_24757);
nand UO_1007 (O_1007,N_24814,N_22658);
nand UO_1008 (O_1008,N_23471,N_23656);
nor UO_1009 (O_1009,N_24885,N_22567);
xnor UO_1010 (O_1010,N_24082,N_22855);
and UO_1011 (O_1011,N_22878,N_23331);
xor UO_1012 (O_1012,N_23278,N_24730);
nor UO_1013 (O_1013,N_23643,N_23759);
and UO_1014 (O_1014,N_24413,N_22846);
nor UO_1015 (O_1015,N_22692,N_23833);
nor UO_1016 (O_1016,N_22582,N_22580);
or UO_1017 (O_1017,N_24496,N_24656);
xor UO_1018 (O_1018,N_23610,N_24512);
or UO_1019 (O_1019,N_23928,N_22967);
nand UO_1020 (O_1020,N_24193,N_23102);
nor UO_1021 (O_1021,N_23537,N_23466);
nor UO_1022 (O_1022,N_22876,N_23522);
nor UO_1023 (O_1023,N_23779,N_23757);
or UO_1024 (O_1024,N_22920,N_22982);
or UO_1025 (O_1025,N_22902,N_23845);
or UO_1026 (O_1026,N_22749,N_24210);
or UO_1027 (O_1027,N_24123,N_23386);
or UO_1028 (O_1028,N_24820,N_23623);
nor UO_1029 (O_1029,N_22893,N_24357);
or UO_1030 (O_1030,N_23054,N_24758);
or UO_1031 (O_1031,N_23689,N_24459);
nor UO_1032 (O_1032,N_24347,N_24973);
nand UO_1033 (O_1033,N_23688,N_24115);
or UO_1034 (O_1034,N_22772,N_23830);
nor UO_1035 (O_1035,N_22853,N_24999);
nand UO_1036 (O_1036,N_24672,N_22891);
nand UO_1037 (O_1037,N_24773,N_22703);
and UO_1038 (O_1038,N_23619,N_22887);
xor UO_1039 (O_1039,N_24422,N_23359);
nor UO_1040 (O_1040,N_24430,N_24199);
or UO_1041 (O_1041,N_23822,N_22946);
or UO_1042 (O_1042,N_23945,N_24055);
xor UO_1043 (O_1043,N_23587,N_24049);
xnor UO_1044 (O_1044,N_24197,N_23577);
nor UO_1045 (O_1045,N_23275,N_23310);
xnor UO_1046 (O_1046,N_24013,N_24120);
nand UO_1047 (O_1047,N_22803,N_24621);
and UO_1048 (O_1048,N_24873,N_24782);
nor UO_1049 (O_1049,N_24194,N_22882);
xor UO_1050 (O_1050,N_24157,N_22646);
xnor UO_1051 (O_1051,N_24337,N_23557);
or UO_1052 (O_1052,N_23815,N_24572);
nor UO_1053 (O_1053,N_24917,N_23161);
xor UO_1054 (O_1054,N_24252,N_22808);
nor UO_1055 (O_1055,N_22506,N_24270);
nand UO_1056 (O_1056,N_24972,N_24795);
xor UO_1057 (O_1057,N_24353,N_24827);
or UO_1058 (O_1058,N_23355,N_24170);
xor UO_1059 (O_1059,N_22654,N_22841);
and UO_1060 (O_1060,N_22557,N_24434);
or UO_1061 (O_1061,N_23824,N_22510);
xnor UO_1062 (O_1062,N_23214,N_24472);
nor UO_1063 (O_1063,N_24909,N_24593);
nand UO_1064 (O_1064,N_24128,N_24517);
xor UO_1065 (O_1065,N_22981,N_24601);
nand UO_1066 (O_1066,N_23677,N_23453);
and UO_1067 (O_1067,N_24062,N_24919);
nor UO_1068 (O_1068,N_24007,N_22611);
or UO_1069 (O_1069,N_22585,N_23086);
or UO_1070 (O_1070,N_23084,N_22797);
nor UO_1071 (O_1071,N_23227,N_24108);
nor UO_1072 (O_1072,N_24048,N_24879);
or UO_1073 (O_1073,N_23773,N_24226);
and UO_1074 (O_1074,N_23418,N_23336);
nand UO_1075 (O_1075,N_23287,N_23479);
nand UO_1076 (O_1076,N_23032,N_23941);
nand UO_1077 (O_1077,N_22935,N_24254);
nor UO_1078 (O_1078,N_24192,N_23295);
nand UO_1079 (O_1079,N_22908,N_24797);
xnor UO_1080 (O_1080,N_24775,N_23073);
nand UO_1081 (O_1081,N_23761,N_24765);
and UO_1082 (O_1082,N_23382,N_22513);
nor UO_1083 (O_1083,N_22770,N_24231);
or UO_1084 (O_1084,N_24786,N_23475);
or UO_1085 (O_1085,N_22865,N_22781);
nand UO_1086 (O_1086,N_24031,N_22665);
and UO_1087 (O_1087,N_23940,N_22907);
nand UO_1088 (O_1088,N_24427,N_24155);
and UO_1089 (O_1089,N_23993,N_24291);
xnor UO_1090 (O_1090,N_24246,N_23307);
and UO_1091 (O_1091,N_24745,N_23647);
nor UO_1092 (O_1092,N_24622,N_24099);
or UO_1093 (O_1093,N_24401,N_23634);
nand UO_1094 (O_1094,N_22912,N_24752);
xor UO_1095 (O_1095,N_23630,N_24426);
nand UO_1096 (O_1096,N_23347,N_23029);
or UO_1097 (O_1097,N_23410,N_24798);
or UO_1098 (O_1098,N_22962,N_23569);
nor UO_1099 (O_1099,N_23099,N_24791);
nand UO_1100 (O_1100,N_22504,N_24734);
nor UO_1101 (O_1101,N_22641,N_24920);
and UO_1102 (O_1102,N_23740,N_24704);
and UO_1103 (O_1103,N_24201,N_23591);
nor UO_1104 (O_1104,N_24489,N_23160);
and UO_1105 (O_1105,N_24483,N_24354);
xor UO_1106 (O_1106,N_23532,N_24888);
xor UO_1107 (O_1107,N_23167,N_24079);
nand UO_1108 (O_1108,N_23657,N_22810);
xnor UO_1109 (O_1109,N_24504,N_23284);
xor UO_1110 (O_1110,N_23213,N_24949);
or UO_1111 (O_1111,N_24250,N_23162);
nor UO_1112 (O_1112,N_24361,N_23201);
or UO_1113 (O_1113,N_23065,N_24498);
xnor UO_1114 (O_1114,N_24453,N_23156);
or UO_1115 (O_1115,N_22877,N_23423);
nand UO_1116 (O_1116,N_23435,N_23031);
and UO_1117 (O_1117,N_23198,N_22933);
and UO_1118 (O_1118,N_24596,N_24706);
and UO_1119 (O_1119,N_24812,N_22664);
or UO_1120 (O_1120,N_24637,N_23390);
and UO_1121 (O_1121,N_23556,N_23769);
xnor UO_1122 (O_1122,N_23693,N_23259);
nor UO_1123 (O_1123,N_22667,N_22545);
xnor UO_1124 (O_1124,N_24518,N_24276);
nor UO_1125 (O_1125,N_23106,N_23300);
nand UO_1126 (O_1126,N_22737,N_24446);
nor UO_1127 (O_1127,N_24590,N_24421);
nand UO_1128 (O_1128,N_22603,N_22614);
nor UO_1129 (O_1129,N_24313,N_22858);
nand UO_1130 (O_1130,N_23019,N_24167);
and UO_1131 (O_1131,N_24025,N_22792);
xnor UO_1132 (O_1132,N_24714,N_22728);
nor UO_1133 (O_1133,N_23918,N_24856);
and UO_1134 (O_1134,N_24023,N_22985);
and UO_1135 (O_1135,N_23699,N_24645);
nand UO_1136 (O_1136,N_22996,N_22835);
nand UO_1137 (O_1137,N_23957,N_24469);
nor UO_1138 (O_1138,N_23882,N_23402);
nand UO_1139 (O_1139,N_23844,N_24940);
or UO_1140 (O_1140,N_22631,N_24780);
and UO_1141 (O_1141,N_23013,N_24219);
nor UO_1142 (O_1142,N_24265,N_24064);
or UO_1143 (O_1143,N_22595,N_23289);
nor UO_1144 (O_1144,N_24407,N_24038);
and UO_1145 (O_1145,N_23652,N_22644);
or UO_1146 (O_1146,N_24171,N_23155);
and UO_1147 (O_1147,N_22550,N_24561);
and UO_1148 (O_1148,N_23045,N_24822);
and UO_1149 (O_1149,N_22523,N_23265);
nand UO_1150 (O_1150,N_23922,N_23741);
xor UO_1151 (O_1151,N_23094,N_23012);
nor UO_1152 (O_1152,N_22926,N_23764);
nand UO_1153 (O_1153,N_23575,N_22731);
or UO_1154 (O_1154,N_24490,N_24690);
nand UO_1155 (O_1155,N_23595,N_24066);
nor UO_1156 (O_1156,N_23760,N_24355);
or UO_1157 (O_1157,N_23567,N_22998);
nand UO_1158 (O_1158,N_24652,N_23481);
xnor UO_1159 (O_1159,N_23765,N_23077);
or UO_1160 (O_1160,N_22517,N_23826);
and UO_1161 (O_1161,N_24370,N_24423);
nand UO_1162 (O_1162,N_23686,N_23228);
nand UO_1163 (O_1163,N_23990,N_24161);
or UO_1164 (O_1164,N_22798,N_24609);
xor UO_1165 (O_1165,N_22583,N_23323);
nor UO_1166 (O_1166,N_24381,N_23078);
nor UO_1167 (O_1167,N_24144,N_24663);
xnor UO_1168 (O_1168,N_23474,N_24039);
xnor UO_1169 (O_1169,N_23360,N_24117);
and UO_1170 (O_1170,N_23405,N_22564);
or UO_1171 (O_1171,N_22562,N_22788);
or UO_1172 (O_1172,N_24674,N_24369);
nor UO_1173 (O_1173,N_23780,N_22734);
nor UO_1174 (O_1174,N_23074,N_22532);
nor UO_1175 (O_1175,N_24880,N_23119);
nor UO_1176 (O_1176,N_23129,N_23887);
or UO_1177 (O_1177,N_24868,N_22574);
nand UO_1178 (O_1178,N_23746,N_22618);
nor UO_1179 (O_1179,N_22830,N_24852);
nor UO_1180 (O_1180,N_23349,N_24938);
or UO_1181 (O_1181,N_23607,N_23164);
and UO_1182 (O_1182,N_23107,N_23758);
xnor UO_1183 (O_1183,N_23148,N_22874);
xnor UO_1184 (O_1184,N_22984,N_24091);
or UO_1185 (O_1185,N_24774,N_23999);
and UO_1186 (O_1186,N_24501,N_24237);
nand UO_1187 (O_1187,N_22645,N_24756);
xnor UO_1188 (O_1188,N_23593,N_24996);
and UO_1189 (O_1189,N_24267,N_23786);
nor UO_1190 (O_1190,N_24485,N_23303);
and UO_1191 (O_1191,N_23771,N_23868);
xnor UO_1192 (O_1192,N_23666,N_23172);
nand UO_1193 (O_1193,N_24307,N_22711);
and UO_1194 (O_1194,N_22773,N_24647);
nand UO_1195 (O_1195,N_22978,N_23542);
and UO_1196 (O_1196,N_24892,N_22673);
nand UO_1197 (O_1197,N_23171,N_23139);
xor UO_1198 (O_1198,N_24567,N_24130);
nand UO_1199 (O_1199,N_23118,N_24374);
and UO_1200 (O_1200,N_23173,N_24388);
nand UO_1201 (O_1201,N_24000,N_22694);
nor UO_1202 (O_1202,N_24075,N_22914);
xor UO_1203 (O_1203,N_22927,N_23473);
xor UO_1204 (O_1204,N_24592,N_22669);
and UO_1205 (O_1205,N_24701,N_24236);
nor UO_1206 (O_1206,N_23092,N_22520);
or UO_1207 (O_1207,N_23703,N_23584);
nor UO_1208 (O_1208,N_23098,N_23229);
nand UO_1209 (O_1209,N_24644,N_24060);
or UO_1210 (O_1210,N_23772,N_24753);
or UO_1211 (O_1211,N_24186,N_23986);
and UO_1212 (O_1212,N_24218,N_24833);
nand UO_1213 (O_1213,N_24925,N_24175);
and UO_1214 (O_1214,N_22802,N_24478);
xnor UO_1215 (O_1215,N_23437,N_23966);
or UO_1216 (O_1216,N_24356,N_24076);
nor UO_1217 (O_1217,N_22928,N_23608);
nor UO_1218 (O_1218,N_23859,N_24457);
nor UO_1219 (O_1219,N_24911,N_24168);
or UO_1220 (O_1220,N_24615,N_22591);
nand UO_1221 (O_1221,N_24495,N_23533);
nor UO_1222 (O_1222,N_24597,N_23631);
xor UO_1223 (O_1223,N_23433,N_23629);
and UO_1224 (O_1224,N_22507,N_24143);
nand UO_1225 (O_1225,N_24135,N_23895);
xnor UO_1226 (O_1226,N_24377,N_23770);
nor UO_1227 (O_1227,N_23449,N_24359);
xnor UO_1228 (O_1228,N_24729,N_24442);
nand UO_1229 (O_1229,N_23028,N_24207);
nand UO_1230 (O_1230,N_23894,N_24152);
nor UO_1231 (O_1231,N_24625,N_23389);
nand UO_1232 (O_1232,N_24839,N_23175);
xnor UO_1233 (O_1233,N_23315,N_22688);
and UO_1234 (O_1234,N_23395,N_22596);
or UO_1235 (O_1235,N_24995,N_23611);
nand UO_1236 (O_1236,N_23545,N_22690);
or UO_1237 (O_1237,N_24994,N_24581);
nand UO_1238 (O_1238,N_22807,N_23727);
nand UO_1239 (O_1239,N_24655,N_23335);
xnor UO_1240 (O_1240,N_24863,N_24578);
nor UO_1241 (O_1241,N_24132,N_24599);
and UO_1242 (O_1242,N_22897,N_23715);
nand UO_1243 (O_1243,N_24682,N_23624);
nand UO_1244 (O_1244,N_23224,N_23509);
or UO_1245 (O_1245,N_23934,N_23087);
nor UO_1246 (O_1246,N_23333,N_23806);
xnor UO_1247 (O_1247,N_24520,N_23057);
and UO_1248 (O_1248,N_22793,N_24515);
and UO_1249 (O_1249,N_24840,N_24941);
xor UO_1250 (O_1250,N_22605,N_23962);
nor UO_1251 (O_1251,N_23857,N_23178);
xor UO_1252 (O_1252,N_23475,N_22858);
nand UO_1253 (O_1253,N_22693,N_22563);
or UO_1254 (O_1254,N_22960,N_23854);
nor UO_1255 (O_1255,N_23563,N_24788);
xor UO_1256 (O_1256,N_22834,N_23044);
nor UO_1257 (O_1257,N_24785,N_23137);
nor UO_1258 (O_1258,N_24124,N_22547);
nand UO_1259 (O_1259,N_22659,N_24472);
nor UO_1260 (O_1260,N_23508,N_24354);
or UO_1261 (O_1261,N_23220,N_22881);
nand UO_1262 (O_1262,N_23248,N_22772);
or UO_1263 (O_1263,N_23526,N_24883);
or UO_1264 (O_1264,N_24383,N_24877);
xnor UO_1265 (O_1265,N_24277,N_22737);
and UO_1266 (O_1266,N_22952,N_24339);
and UO_1267 (O_1267,N_24000,N_23324);
and UO_1268 (O_1268,N_23597,N_24513);
xor UO_1269 (O_1269,N_22835,N_24524);
or UO_1270 (O_1270,N_24615,N_22848);
or UO_1271 (O_1271,N_23152,N_23117);
nor UO_1272 (O_1272,N_23243,N_22585);
nand UO_1273 (O_1273,N_24854,N_23446);
xnor UO_1274 (O_1274,N_24382,N_23817);
nor UO_1275 (O_1275,N_24904,N_23959);
or UO_1276 (O_1276,N_24104,N_24853);
xnor UO_1277 (O_1277,N_24007,N_23029);
nand UO_1278 (O_1278,N_23043,N_23963);
nand UO_1279 (O_1279,N_23378,N_23649);
or UO_1280 (O_1280,N_22932,N_23414);
nand UO_1281 (O_1281,N_24961,N_24717);
and UO_1282 (O_1282,N_22617,N_23736);
xnor UO_1283 (O_1283,N_22874,N_24180);
nor UO_1284 (O_1284,N_22771,N_24877);
nand UO_1285 (O_1285,N_23948,N_24700);
xnor UO_1286 (O_1286,N_22875,N_24191);
and UO_1287 (O_1287,N_22610,N_24604);
xnor UO_1288 (O_1288,N_24698,N_24962);
xor UO_1289 (O_1289,N_24063,N_24772);
nand UO_1290 (O_1290,N_24909,N_23400);
and UO_1291 (O_1291,N_22654,N_23789);
nand UO_1292 (O_1292,N_23817,N_23942);
or UO_1293 (O_1293,N_23637,N_22815);
nor UO_1294 (O_1294,N_23808,N_24699);
nor UO_1295 (O_1295,N_24479,N_24679);
xnor UO_1296 (O_1296,N_22909,N_22576);
nand UO_1297 (O_1297,N_22937,N_24333);
and UO_1298 (O_1298,N_23477,N_23013);
nand UO_1299 (O_1299,N_24270,N_23096);
nor UO_1300 (O_1300,N_24715,N_24707);
and UO_1301 (O_1301,N_23210,N_24829);
nor UO_1302 (O_1302,N_24302,N_24862);
nor UO_1303 (O_1303,N_24649,N_23539);
nor UO_1304 (O_1304,N_23307,N_22907);
or UO_1305 (O_1305,N_23331,N_23427);
nor UO_1306 (O_1306,N_22835,N_23044);
nor UO_1307 (O_1307,N_24256,N_24494);
nor UO_1308 (O_1308,N_24282,N_23654);
and UO_1309 (O_1309,N_23314,N_22645);
nor UO_1310 (O_1310,N_22627,N_24463);
and UO_1311 (O_1311,N_23120,N_24205);
or UO_1312 (O_1312,N_24890,N_22875);
xnor UO_1313 (O_1313,N_24940,N_22647);
xnor UO_1314 (O_1314,N_23637,N_22881);
nor UO_1315 (O_1315,N_24615,N_23510);
xor UO_1316 (O_1316,N_22890,N_24576);
and UO_1317 (O_1317,N_24465,N_24085);
nand UO_1318 (O_1318,N_22797,N_23675);
xnor UO_1319 (O_1319,N_24646,N_23846);
and UO_1320 (O_1320,N_22904,N_23778);
or UO_1321 (O_1321,N_24181,N_24800);
or UO_1322 (O_1322,N_22772,N_23837);
and UO_1323 (O_1323,N_23515,N_24495);
nor UO_1324 (O_1324,N_24924,N_23930);
and UO_1325 (O_1325,N_23207,N_23918);
nand UO_1326 (O_1326,N_24808,N_24515);
or UO_1327 (O_1327,N_22662,N_23728);
xnor UO_1328 (O_1328,N_23150,N_23521);
xor UO_1329 (O_1329,N_24097,N_24084);
xnor UO_1330 (O_1330,N_24721,N_24483);
nand UO_1331 (O_1331,N_23374,N_23770);
or UO_1332 (O_1332,N_23164,N_24296);
and UO_1333 (O_1333,N_24221,N_24919);
and UO_1334 (O_1334,N_22999,N_23564);
nor UO_1335 (O_1335,N_24202,N_23502);
nand UO_1336 (O_1336,N_24249,N_22608);
nor UO_1337 (O_1337,N_22807,N_22960);
or UO_1338 (O_1338,N_23805,N_24360);
nor UO_1339 (O_1339,N_24720,N_23022);
xor UO_1340 (O_1340,N_24375,N_23058);
xnor UO_1341 (O_1341,N_24584,N_22765);
and UO_1342 (O_1342,N_24245,N_23999);
nor UO_1343 (O_1343,N_24007,N_22995);
xnor UO_1344 (O_1344,N_24796,N_23294);
and UO_1345 (O_1345,N_22929,N_24983);
nand UO_1346 (O_1346,N_24027,N_24911);
and UO_1347 (O_1347,N_23852,N_23799);
nand UO_1348 (O_1348,N_24524,N_24111);
nor UO_1349 (O_1349,N_23986,N_23206);
or UO_1350 (O_1350,N_23338,N_24347);
nand UO_1351 (O_1351,N_23922,N_24908);
or UO_1352 (O_1352,N_24120,N_24409);
xnor UO_1353 (O_1353,N_22951,N_22728);
xnor UO_1354 (O_1354,N_23737,N_23137);
xnor UO_1355 (O_1355,N_23704,N_24031);
xor UO_1356 (O_1356,N_23594,N_22561);
xor UO_1357 (O_1357,N_23650,N_22897);
xnor UO_1358 (O_1358,N_24420,N_23264);
nand UO_1359 (O_1359,N_24314,N_23024);
nand UO_1360 (O_1360,N_22500,N_24689);
xnor UO_1361 (O_1361,N_23014,N_23262);
or UO_1362 (O_1362,N_24456,N_24307);
nand UO_1363 (O_1363,N_24651,N_24997);
or UO_1364 (O_1364,N_24597,N_23770);
and UO_1365 (O_1365,N_22665,N_23902);
nor UO_1366 (O_1366,N_23796,N_23517);
xnor UO_1367 (O_1367,N_23352,N_23082);
or UO_1368 (O_1368,N_24264,N_23362);
and UO_1369 (O_1369,N_22690,N_22982);
or UO_1370 (O_1370,N_22577,N_22732);
xor UO_1371 (O_1371,N_22721,N_23305);
and UO_1372 (O_1372,N_22781,N_23259);
nand UO_1373 (O_1373,N_23258,N_24376);
nand UO_1374 (O_1374,N_24963,N_22940);
and UO_1375 (O_1375,N_22745,N_24353);
nand UO_1376 (O_1376,N_24169,N_22995);
xor UO_1377 (O_1377,N_24911,N_23413);
or UO_1378 (O_1378,N_23573,N_23810);
nor UO_1379 (O_1379,N_23449,N_22902);
or UO_1380 (O_1380,N_24122,N_24555);
nor UO_1381 (O_1381,N_23913,N_22823);
or UO_1382 (O_1382,N_23469,N_24677);
or UO_1383 (O_1383,N_23307,N_23911);
or UO_1384 (O_1384,N_23560,N_24991);
nor UO_1385 (O_1385,N_23224,N_23358);
nand UO_1386 (O_1386,N_22977,N_24268);
nand UO_1387 (O_1387,N_24157,N_22676);
nor UO_1388 (O_1388,N_24533,N_22781);
and UO_1389 (O_1389,N_23436,N_23113);
nor UO_1390 (O_1390,N_22662,N_24471);
nand UO_1391 (O_1391,N_23883,N_24272);
nand UO_1392 (O_1392,N_24408,N_22716);
nand UO_1393 (O_1393,N_23880,N_24347);
and UO_1394 (O_1394,N_24837,N_23506);
nor UO_1395 (O_1395,N_23509,N_24589);
and UO_1396 (O_1396,N_22713,N_23125);
nor UO_1397 (O_1397,N_22507,N_23243);
xnor UO_1398 (O_1398,N_24522,N_23900);
nand UO_1399 (O_1399,N_24700,N_24012);
nor UO_1400 (O_1400,N_23512,N_23688);
nor UO_1401 (O_1401,N_24582,N_24402);
or UO_1402 (O_1402,N_24926,N_23472);
and UO_1403 (O_1403,N_23111,N_24072);
or UO_1404 (O_1404,N_23106,N_24500);
or UO_1405 (O_1405,N_24265,N_23795);
or UO_1406 (O_1406,N_23571,N_23867);
xor UO_1407 (O_1407,N_22856,N_24452);
and UO_1408 (O_1408,N_24587,N_23729);
nor UO_1409 (O_1409,N_23327,N_23264);
and UO_1410 (O_1410,N_23234,N_24396);
and UO_1411 (O_1411,N_23955,N_23256);
nor UO_1412 (O_1412,N_24494,N_23373);
xnor UO_1413 (O_1413,N_22687,N_23861);
nor UO_1414 (O_1414,N_24267,N_23969);
nand UO_1415 (O_1415,N_24533,N_24152);
nand UO_1416 (O_1416,N_23548,N_24601);
nor UO_1417 (O_1417,N_23278,N_23225);
or UO_1418 (O_1418,N_24391,N_22630);
xor UO_1419 (O_1419,N_24389,N_23488);
nand UO_1420 (O_1420,N_23226,N_23957);
nor UO_1421 (O_1421,N_22780,N_23945);
xor UO_1422 (O_1422,N_22825,N_22902);
xnor UO_1423 (O_1423,N_23861,N_22967);
nor UO_1424 (O_1424,N_22794,N_24390);
nand UO_1425 (O_1425,N_23106,N_22929);
and UO_1426 (O_1426,N_24328,N_23620);
nand UO_1427 (O_1427,N_23443,N_24426);
and UO_1428 (O_1428,N_24078,N_24505);
and UO_1429 (O_1429,N_22781,N_24436);
or UO_1430 (O_1430,N_22527,N_23950);
nor UO_1431 (O_1431,N_24566,N_23565);
and UO_1432 (O_1432,N_22591,N_22532);
nand UO_1433 (O_1433,N_24701,N_23845);
nand UO_1434 (O_1434,N_23711,N_24883);
nor UO_1435 (O_1435,N_24572,N_24409);
or UO_1436 (O_1436,N_24905,N_22902);
or UO_1437 (O_1437,N_24603,N_24918);
nand UO_1438 (O_1438,N_22812,N_22760);
or UO_1439 (O_1439,N_23089,N_23646);
nor UO_1440 (O_1440,N_22787,N_24811);
nand UO_1441 (O_1441,N_22558,N_22754);
nand UO_1442 (O_1442,N_23221,N_23565);
or UO_1443 (O_1443,N_23422,N_22788);
xnor UO_1444 (O_1444,N_22752,N_24115);
xnor UO_1445 (O_1445,N_22985,N_24452);
xnor UO_1446 (O_1446,N_23794,N_22849);
nand UO_1447 (O_1447,N_24590,N_23305);
and UO_1448 (O_1448,N_24964,N_23424);
or UO_1449 (O_1449,N_24606,N_24027);
and UO_1450 (O_1450,N_23724,N_22592);
nor UO_1451 (O_1451,N_24076,N_24892);
nand UO_1452 (O_1452,N_24852,N_22561);
or UO_1453 (O_1453,N_24447,N_23915);
nand UO_1454 (O_1454,N_23151,N_24134);
nand UO_1455 (O_1455,N_22522,N_24191);
nand UO_1456 (O_1456,N_23684,N_24871);
nand UO_1457 (O_1457,N_23945,N_24294);
nand UO_1458 (O_1458,N_24503,N_23971);
nor UO_1459 (O_1459,N_24546,N_23729);
nor UO_1460 (O_1460,N_23683,N_24321);
xor UO_1461 (O_1461,N_24908,N_22784);
xnor UO_1462 (O_1462,N_23844,N_23767);
and UO_1463 (O_1463,N_24338,N_22917);
or UO_1464 (O_1464,N_23699,N_23025);
nor UO_1465 (O_1465,N_23970,N_22636);
xnor UO_1466 (O_1466,N_22520,N_23046);
or UO_1467 (O_1467,N_24789,N_24054);
or UO_1468 (O_1468,N_23742,N_22589);
nor UO_1469 (O_1469,N_24785,N_23083);
or UO_1470 (O_1470,N_23277,N_24339);
nand UO_1471 (O_1471,N_23148,N_23482);
nor UO_1472 (O_1472,N_23043,N_24448);
xor UO_1473 (O_1473,N_22658,N_24132);
or UO_1474 (O_1474,N_24629,N_23153);
and UO_1475 (O_1475,N_24707,N_23707);
nand UO_1476 (O_1476,N_23957,N_23430);
nor UO_1477 (O_1477,N_22834,N_23879);
xnor UO_1478 (O_1478,N_23657,N_23108);
or UO_1479 (O_1479,N_23661,N_23897);
nor UO_1480 (O_1480,N_22743,N_23626);
or UO_1481 (O_1481,N_24153,N_22704);
nor UO_1482 (O_1482,N_23153,N_23045);
xnor UO_1483 (O_1483,N_24822,N_24969);
and UO_1484 (O_1484,N_22797,N_23354);
or UO_1485 (O_1485,N_22539,N_24308);
xnor UO_1486 (O_1486,N_23484,N_24700);
nand UO_1487 (O_1487,N_23831,N_23129);
and UO_1488 (O_1488,N_24895,N_23770);
or UO_1489 (O_1489,N_23732,N_23721);
or UO_1490 (O_1490,N_23860,N_24204);
and UO_1491 (O_1491,N_22806,N_24675);
nand UO_1492 (O_1492,N_23594,N_23116);
xor UO_1493 (O_1493,N_24096,N_24984);
xnor UO_1494 (O_1494,N_24415,N_24587);
xor UO_1495 (O_1495,N_23007,N_24431);
nand UO_1496 (O_1496,N_24331,N_23931);
xor UO_1497 (O_1497,N_22704,N_22530);
nand UO_1498 (O_1498,N_23850,N_24064);
nand UO_1499 (O_1499,N_24029,N_24228);
nor UO_1500 (O_1500,N_24457,N_23643);
or UO_1501 (O_1501,N_24404,N_23381);
and UO_1502 (O_1502,N_24471,N_24973);
and UO_1503 (O_1503,N_23987,N_23761);
xnor UO_1504 (O_1504,N_24592,N_24812);
xnor UO_1505 (O_1505,N_24637,N_23663);
or UO_1506 (O_1506,N_23401,N_23837);
nor UO_1507 (O_1507,N_22613,N_24137);
and UO_1508 (O_1508,N_22804,N_23551);
and UO_1509 (O_1509,N_24405,N_24564);
nor UO_1510 (O_1510,N_22627,N_24855);
or UO_1511 (O_1511,N_22720,N_22961);
or UO_1512 (O_1512,N_23966,N_24198);
nor UO_1513 (O_1513,N_23576,N_23985);
nor UO_1514 (O_1514,N_24271,N_24173);
nand UO_1515 (O_1515,N_24420,N_23169);
or UO_1516 (O_1516,N_23537,N_23736);
xnor UO_1517 (O_1517,N_23775,N_23633);
or UO_1518 (O_1518,N_24597,N_24782);
xnor UO_1519 (O_1519,N_22559,N_24886);
or UO_1520 (O_1520,N_24155,N_24503);
xor UO_1521 (O_1521,N_24606,N_23525);
or UO_1522 (O_1522,N_24997,N_24146);
nor UO_1523 (O_1523,N_22938,N_24078);
nand UO_1524 (O_1524,N_24849,N_23057);
nor UO_1525 (O_1525,N_22627,N_24154);
and UO_1526 (O_1526,N_23355,N_23061);
or UO_1527 (O_1527,N_23496,N_23336);
nor UO_1528 (O_1528,N_23308,N_23791);
or UO_1529 (O_1529,N_23475,N_23792);
nor UO_1530 (O_1530,N_23247,N_23084);
or UO_1531 (O_1531,N_23157,N_24248);
nor UO_1532 (O_1532,N_24110,N_24797);
xor UO_1533 (O_1533,N_23142,N_24960);
and UO_1534 (O_1534,N_24578,N_22859);
xor UO_1535 (O_1535,N_24847,N_23304);
nand UO_1536 (O_1536,N_24563,N_24234);
xor UO_1537 (O_1537,N_24171,N_23588);
and UO_1538 (O_1538,N_23183,N_22803);
and UO_1539 (O_1539,N_24711,N_23828);
or UO_1540 (O_1540,N_24224,N_23314);
nand UO_1541 (O_1541,N_22872,N_24094);
or UO_1542 (O_1542,N_24784,N_23397);
nor UO_1543 (O_1543,N_23647,N_23076);
xor UO_1544 (O_1544,N_23530,N_23478);
or UO_1545 (O_1545,N_24083,N_24906);
and UO_1546 (O_1546,N_23610,N_23401);
and UO_1547 (O_1547,N_23727,N_24383);
or UO_1548 (O_1548,N_22718,N_22568);
and UO_1549 (O_1549,N_23138,N_24439);
xnor UO_1550 (O_1550,N_23337,N_23014);
xnor UO_1551 (O_1551,N_23589,N_24871);
or UO_1552 (O_1552,N_24423,N_23867);
or UO_1553 (O_1553,N_24517,N_24035);
xnor UO_1554 (O_1554,N_22531,N_24332);
and UO_1555 (O_1555,N_23527,N_23001);
and UO_1556 (O_1556,N_24840,N_22673);
or UO_1557 (O_1557,N_24388,N_23520);
and UO_1558 (O_1558,N_24491,N_24265);
nand UO_1559 (O_1559,N_22540,N_23732);
and UO_1560 (O_1560,N_23740,N_24986);
nor UO_1561 (O_1561,N_23065,N_23884);
nor UO_1562 (O_1562,N_24182,N_23028);
or UO_1563 (O_1563,N_24563,N_24068);
xnor UO_1564 (O_1564,N_23557,N_23386);
nor UO_1565 (O_1565,N_24277,N_24576);
and UO_1566 (O_1566,N_23120,N_23050);
and UO_1567 (O_1567,N_24972,N_24898);
and UO_1568 (O_1568,N_23559,N_22795);
nand UO_1569 (O_1569,N_23903,N_23593);
nor UO_1570 (O_1570,N_24326,N_23269);
xnor UO_1571 (O_1571,N_24596,N_24300);
or UO_1572 (O_1572,N_23876,N_24592);
nand UO_1573 (O_1573,N_22731,N_23462);
nor UO_1574 (O_1574,N_23160,N_24513);
nand UO_1575 (O_1575,N_23632,N_22738);
xnor UO_1576 (O_1576,N_24274,N_24849);
or UO_1577 (O_1577,N_24411,N_24867);
nand UO_1578 (O_1578,N_22939,N_22822);
or UO_1579 (O_1579,N_23275,N_24900);
nand UO_1580 (O_1580,N_22825,N_22566);
or UO_1581 (O_1581,N_24126,N_22500);
and UO_1582 (O_1582,N_24534,N_24348);
nand UO_1583 (O_1583,N_24439,N_23926);
and UO_1584 (O_1584,N_22708,N_23712);
nand UO_1585 (O_1585,N_24586,N_23700);
and UO_1586 (O_1586,N_24339,N_23062);
and UO_1587 (O_1587,N_23931,N_22530);
and UO_1588 (O_1588,N_24629,N_22968);
or UO_1589 (O_1589,N_23714,N_22768);
nor UO_1590 (O_1590,N_22870,N_23323);
nand UO_1591 (O_1591,N_24158,N_23879);
xnor UO_1592 (O_1592,N_24467,N_22627);
or UO_1593 (O_1593,N_24668,N_22651);
or UO_1594 (O_1594,N_23739,N_22619);
nand UO_1595 (O_1595,N_24189,N_24239);
or UO_1596 (O_1596,N_24322,N_22700);
nand UO_1597 (O_1597,N_22657,N_23460);
or UO_1598 (O_1598,N_23533,N_24459);
or UO_1599 (O_1599,N_24444,N_24063);
nand UO_1600 (O_1600,N_23238,N_23750);
nand UO_1601 (O_1601,N_24581,N_24811);
xor UO_1602 (O_1602,N_23916,N_22568);
and UO_1603 (O_1603,N_24815,N_24334);
and UO_1604 (O_1604,N_23432,N_24469);
nor UO_1605 (O_1605,N_24482,N_24696);
or UO_1606 (O_1606,N_23582,N_23386);
nand UO_1607 (O_1607,N_23568,N_22785);
xnor UO_1608 (O_1608,N_23204,N_23125);
and UO_1609 (O_1609,N_24585,N_24245);
and UO_1610 (O_1610,N_24352,N_24644);
or UO_1611 (O_1611,N_24621,N_24977);
nor UO_1612 (O_1612,N_23953,N_23113);
nor UO_1613 (O_1613,N_24877,N_23056);
xnor UO_1614 (O_1614,N_24490,N_24341);
or UO_1615 (O_1615,N_23331,N_24992);
or UO_1616 (O_1616,N_23394,N_22996);
xor UO_1617 (O_1617,N_24064,N_23221);
nand UO_1618 (O_1618,N_23081,N_24431);
nor UO_1619 (O_1619,N_24452,N_22501);
xnor UO_1620 (O_1620,N_22908,N_24037);
and UO_1621 (O_1621,N_24394,N_23307);
nand UO_1622 (O_1622,N_23411,N_23307);
xnor UO_1623 (O_1623,N_24118,N_23535);
or UO_1624 (O_1624,N_23008,N_24567);
and UO_1625 (O_1625,N_23700,N_23112);
or UO_1626 (O_1626,N_23272,N_24561);
nor UO_1627 (O_1627,N_24946,N_24986);
xor UO_1628 (O_1628,N_23138,N_24814);
and UO_1629 (O_1629,N_23574,N_24218);
nor UO_1630 (O_1630,N_23720,N_22563);
or UO_1631 (O_1631,N_23463,N_24495);
xnor UO_1632 (O_1632,N_23583,N_24082);
and UO_1633 (O_1633,N_23206,N_23500);
nor UO_1634 (O_1634,N_24294,N_24533);
nand UO_1635 (O_1635,N_24882,N_24942);
nor UO_1636 (O_1636,N_23817,N_24018);
nor UO_1637 (O_1637,N_24332,N_24842);
and UO_1638 (O_1638,N_23269,N_24028);
nand UO_1639 (O_1639,N_22735,N_23757);
xnor UO_1640 (O_1640,N_23521,N_23237);
nor UO_1641 (O_1641,N_24131,N_22832);
and UO_1642 (O_1642,N_22755,N_22848);
nor UO_1643 (O_1643,N_23946,N_24566);
and UO_1644 (O_1644,N_24676,N_24291);
or UO_1645 (O_1645,N_22880,N_22601);
or UO_1646 (O_1646,N_24144,N_24975);
xnor UO_1647 (O_1647,N_22721,N_23953);
or UO_1648 (O_1648,N_23548,N_22792);
nand UO_1649 (O_1649,N_22519,N_23723);
nand UO_1650 (O_1650,N_24724,N_23545);
nand UO_1651 (O_1651,N_24155,N_24701);
nor UO_1652 (O_1652,N_23819,N_23099);
and UO_1653 (O_1653,N_22748,N_22575);
xor UO_1654 (O_1654,N_23603,N_22600);
nor UO_1655 (O_1655,N_23306,N_23166);
nand UO_1656 (O_1656,N_23822,N_22735);
or UO_1657 (O_1657,N_22789,N_22939);
nor UO_1658 (O_1658,N_24803,N_24936);
nand UO_1659 (O_1659,N_24872,N_24486);
nand UO_1660 (O_1660,N_23576,N_24991);
nor UO_1661 (O_1661,N_22961,N_23568);
nor UO_1662 (O_1662,N_23426,N_23691);
or UO_1663 (O_1663,N_22559,N_22994);
nand UO_1664 (O_1664,N_22720,N_24253);
nor UO_1665 (O_1665,N_23754,N_22575);
and UO_1666 (O_1666,N_24987,N_24538);
nand UO_1667 (O_1667,N_24188,N_23454);
and UO_1668 (O_1668,N_24892,N_24277);
or UO_1669 (O_1669,N_24083,N_24519);
xnor UO_1670 (O_1670,N_24689,N_24803);
nor UO_1671 (O_1671,N_22955,N_24999);
nand UO_1672 (O_1672,N_23128,N_24852);
nand UO_1673 (O_1673,N_23793,N_22662);
xor UO_1674 (O_1674,N_24873,N_23120);
nand UO_1675 (O_1675,N_24355,N_24683);
and UO_1676 (O_1676,N_24440,N_23584);
or UO_1677 (O_1677,N_23990,N_24736);
and UO_1678 (O_1678,N_23368,N_22968);
nor UO_1679 (O_1679,N_23223,N_22817);
nor UO_1680 (O_1680,N_24293,N_24160);
nand UO_1681 (O_1681,N_23363,N_24325);
and UO_1682 (O_1682,N_23307,N_23268);
nand UO_1683 (O_1683,N_23903,N_22968);
xnor UO_1684 (O_1684,N_24228,N_23985);
nand UO_1685 (O_1685,N_24735,N_24834);
nor UO_1686 (O_1686,N_22629,N_23446);
xnor UO_1687 (O_1687,N_24479,N_24039);
nor UO_1688 (O_1688,N_22817,N_24995);
or UO_1689 (O_1689,N_24914,N_24430);
nor UO_1690 (O_1690,N_24239,N_23680);
and UO_1691 (O_1691,N_24325,N_24145);
nor UO_1692 (O_1692,N_23386,N_23083);
and UO_1693 (O_1693,N_24620,N_22755);
nor UO_1694 (O_1694,N_22521,N_24876);
or UO_1695 (O_1695,N_24145,N_23655);
xor UO_1696 (O_1696,N_22639,N_24740);
xnor UO_1697 (O_1697,N_23402,N_24884);
xor UO_1698 (O_1698,N_23224,N_22693);
nor UO_1699 (O_1699,N_23227,N_23737);
xnor UO_1700 (O_1700,N_24308,N_24521);
xnor UO_1701 (O_1701,N_24115,N_23659);
nand UO_1702 (O_1702,N_22537,N_24071);
nor UO_1703 (O_1703,N_22770,N_24639);
xnor UO_1704 (O_1704,N_24492,N_24646);
xor UO_1705 (O_1705,N_23535,N_24512);
and UO_1706 (O_1706,N_23061,N_22884);
nand UO_1707 (O_1707,N_23025,N_23575);
or UO_1708 (O_1708,N_24770,N_23817);
and UO_1709 (O_1709,N_23619,N_22784);
xnor UO_1710 (O_1710,N_23331,N_24254);
xnor UO_1711 (O_1711,N_24204,N_24567);
nor UO_1712 (O_1712,N_23647,N_22961);
nor UO_1713 (O_1713,N_22840,N_23725);
nand UO_1714 (O_1714,N_24196,N_22997);
nor UO_1715 (O_1715,N_24669,N_24416);
xnor UO_1716 (O_1716,N_22798,N_24227);
nand UO_1717 (O_1717,N_22827,N_24502);
nor UO_1718 (O_1718,N_24161,N_23208);
and UO_1719 (O_1719,N_23170,N_24654);
and UO_1720 (O_1720,N_23888,N_22994);
xor UO_1721 (O_1721,N_23521,N_23558);
or UO_1722 (O_1722,N_22632,N_22645);
xnor UO_1723 (O_1723,N_23924,N_23193);
nand UO_1724 (O_1724,N_23741,N_23074);
nand UO_1725 (O_1725,N_24685,N_24161);
xnor UO_1726 (O_1726,N_23568,N_23479);
nand UO_1727 (O_1727,N_23171,N_24866);
nand UO_1728 (O_1728,N_23359,N_24846);
nor UO_1729 (O_1729,N_22800,N_23678);
and UO_1730 (O_1730,N_24182,N_24373);
nand UO_1731 (O_1731,N_23532,N_24962);
and UO_1732 (O_1732,N_23782,N_24111);
and UO_1733 (O_1733,N_24499,N_22945);
nor UO_1734 (O_1734,N_24171,N_24068);
nand UO_1735 (O_1735,N_24886,N_23177);
nor UO_1736 (O_1736,N_24649,N_22830);
and UO_1737 (O_1737,N_24081,N_24132);
nand UO_1738 (O_1738,N_22989,N_23572);
nor UO_1739 (O_1739,N_24890,N_24819);
nand UO_1740 (O_1740,N_23379,N_24625);
and UO_1741 (O_1741,N_23777,N_22844);
and UO_1742 (O_1742,N_24256,N_24962);
or UO_1743 (O_1743,N_22860,N_24618);
and UO_1744 (O_1744,N_23003,N_22742);
xnor UO_1745 (O_1745,N_23108,N_24912);
nor UO_1746 (O_1746,N_24560,N_24952);
or UO_1747 (O_1747,N_24964,N_24725);
nor UO_1748 (O_1748,N_23782,N_23761);
xor UO_1749 (O_1749,N_23617,N_24909);
nor UO_1750 (O_1750,N_22935,N_22668);
xnor UO_1751 (O_1751,N_22906,N_23844);
and UO_1752 (O_1752,N_24230,N_24053);
xnor UO_1753 (O_1753,N_23444,N_24326);
xor UO_1754 (O_1754,N_23448,N_23158);
nor UO_1755 (O_1755,N_23250,N_22615);
nand UO_1756 (O_1756,N_23097,N_24315);
nor UO_1757 (O_1757,N_22945,N_23194);
xnor UO_1758 (O_1758,N_24366,N_24942);
nor UO_1759 (O_1759,N_23459,N_24905);
and UO_1760 (O_1760,N_23887,N_24671);
or UO_1761 (O_1761,N_24543,N_24590);
or UO_1762 (O_1762,N_24349,N_23034);
or UO_1763 (O_1763,N_23576,N_22837);
nand UO_1764 (O_1764,N_23381,N_23113);
nor UO_1765 (O_1765,N_24939,N_23456);
and UO_1766 (O_1766,N_23693,N_24083);
nand UO_1767 (O_1767,N_23251,N_22715);
or UO_1768 (O_1768,N_22636,N_24607);
nand UO_1769 (O_1769,N_24339,N_24359);
or UO_1770 (O_1770,N_23076,N_22668);
or UO_1771 (O_1771,N_23130,N_24033);
and UO_1772 (O_1772,N_24705,N_24834);
nor UO_1773 (O_1773,N_24228,N_23465);
and UO_1774 (O_1774,N_23503,N_23695);
and UO_1775 (O_1775,N_23593,N_24998);
or UO_1776 (O_1776,N_23617,N_24870);
and UO_1777 (O_1777,N_23216,N_24203);
xor UO_1778 (O_1778,N_24208,N_23747);
nor UO_1779 (O_1779,N_23153,N_24324);
xnor UO_1780 (O_1780,N_23167,N_23170);
and UO_1781 (O_1781,N_22736,N_24798);
and UO_1782 (O_1782,N_23046,N_24046);
and UO_1783 (O_1783,N_24598,N_24273);
nor UO_1784 (O_1784,N_22766,N_24561);
nor UO_1785 (O_1785,N_23443,N_24797);
xor UO_1786 (O_1786,N_22643,N_23498);
nor UO_1787 (O_1787,N_23146,N_24862);
and UO_1788 (O_1788,N_24693,N_24117);
nand UO_1789 (O_1789,N_23480,N_24642);
or UO_1790 (O_1790,N_24759,N_22813);
and UO_1791 (O_1791,N_24170,N_23327);
and UO_1792 (O_1792,N_22987,N_23095);
nand UO_1793 (O_1793,N_24817,N_24733);
xor UO_1794 (O_1794,N_22919,N_24023);
nand UO_1795 (O_1795,N_24290,N_23163);
or UO_1796 (O_1796,N_22521,N_24483);
and UO_1797 (O_1797,N_23159,N_24872);
and UO_1798 (O_1798,N_24256,N_24464);
nand UO_1799 (O_1799,N_23557,N_22912);
xnor UO_1800 (O_1800,N_22944,N_23171);
or UO_1801 (O_1801,N_24654,N_22833);
and UO_1802 (O_1802,N_23563,N_22877);
xor UO_1803 (O_1803,N_22545,N_23118);
or UO_1804 (O_1804,N_22825,N_22612);
xor UO_1805 (O_1805,N_23521,N_23086);
xor UO_1806 (O_1806,N_24656,N_22999);
nand UO_1807 (O_1807,N_23159,N_24325);
or UO_1808 (O_1808,N_23555,N_24633);
xor UO_1809 (O_1809,N_23291,N_22679);
and UO_1810 (O_1810,N_22915,N_23374);
nor UO_1811 (O_1811,N_23897,N_24918);
xnor UO_1812 (O_1812,N_24582,N_23882);
nand UO_1813 (O_1813,N_23857,N_24990);
and UO_1814 (O_1814,N_24323,N_22865);
nor UO_1815 (O_1815,N_23495,N_23393);
nor UO_1816 (O_1816,N_24607,N_24633);
nor UO_1817 (O_1817,N_23654,N_23777);
or UO_1818 (O_1818,N_23920,N_24623);
and UO_1819 (O_1819,N_24091,N_24910);
or UO_1820 (O_1820,N_23054,N_24824);
or UO_1821 (O_1821,N_23635,N_22737);
nand UO_1822 (O_1822,N_24788,N_23994);
nor UO_1823 (O_1823,N_23542,N_24935);
nand UO_1824 (O_1824,N_24761,N_22548);
or UO_1825 (O_1825,N_24816,N_23635);
nand UO_1826 (O_1826,N_24172,N_24595);
and UO_1827 (O_1827,N_24722,N_22897);
xnor UO_1828 (O_1828,N_23980,N_22787);
nor UO_1829 (O_1829,N_24257,N_23091);
or UO_1830 (O_1830,N_23192,N_24025);
nor UO_1831 (O_1831,N_23780,N_24382);
nand UO_1832 (O_1832,N_23176,N_23957);
and UO_1833 (O_1833,N_22530,N_24054);
and UO_1834 (O_1834,N_24424,N_23031);
nor UO_1835 (O_1835,N_22529,N_23413);
nand UO_1836 (O_1836,N_24791,N_23293);
or UO_1837 (O_1837,N_24210,N_24590);
and UO_1838 (O_1838,N_23615,N_24844);
nor UO_1839 (O_1839,N_23594,N_22881);
and UO_1840 (O_1840,N_22804,N_23376);
and UO_1841 (O_1841,N_24898,N_24785);
nand UO_1842 (O_1842,N_22538,N_24130);
or UO_1843 (O_1843,N_23212,N_23032);
and UO_1844 (O_1844,N_23761,N_24771);
nand UO_1845 (O_1845,N_24176,N_22752);
or UO_1846 (O_1846,N_22824,N_23046);
nor UO_1847 (O_1847,N_24981,N_22520);
or UO_1848 (O_1848,N_23453,N_24209);
xor UO_1849 (O_1849,N_22554,N_23590);
nor UO_1850 (O_1850,N_23117,N_24351);
or UO_1851 (O_1851,N_23506,N_23255);
and UO_1852 (O_1852,N_22671,N_23275);
nand UO_1853 (O_1853,N_22601,N_24384);
xnor UO_1854 (O_1854,N_23033,N_23080);
xnor UO_1855 (O_1855,N_24285,N_22980);
xor UO_1856 (O_1856,N_22943,N_24967);
nand UO_1857 (O_1857,N_24429,N_23680);
nand UO_1858 (O_1858,N_23098,N_22824);
and UO_1859 (O_1859,N_22636,N_24414);
nand UO_1860 (O_1860,N_23972,N_24275);
or UO_1861 (O_1861,N_24508,N_24147);
and UO_1862 (O_1862,N_23687,N_23807);
xor UO_1863 (O_1863,N_22858,N_23084);
or UO_1864 (O_1864,N_23607,N_24826);
nand UO_1865 (O_1865,N_22689,N_24762);
and UO_1866 (O_1866,N_24599,N_23432);
or UO_1867 (O_1867,N_24267,N_22528);
or UO_1868 (O_1868,N_24197,N_23321);
and UO_1869 (O_1869,N_23969,N_23010);
nand UO_1870 (O_1870,N_24530,N_23976);
or UO_1871 (O_1871,N_24115,N_23825);
nor UO_1872 (O_1872,N_22738,N_22771);
and UO_1873 (O_1873,N_23541,N_23780);
xor UO_1874 (O_1874,N_24984,N_22926);
nand UO_1875 (O_1875,N_24271,N_23079);
or UO_1876 (O_1876,N_22884,N_24503);
xor UO_1877 (O_1877,N_23267,N_22990);
nand UO_1878 (O_1878,N_22513,N_23160);
nand UO_1879 (O_1879,N_24475,N_24673);
nor UO_1880 (O_1880,N_24426,N_22576);
xor UO_1881 (O_1881,N_22924,N_22648);
xor UO_1882 (O_1882,N_23974,N_24668);
nand UO_1883 (O_1883,N_23087,N_22630);
nand UO_1884 (O_1884,N_24547,N_22767);
nor UO_1885 (O_1885,N_24248,N_23355);
xor UO_1886 (O_1886,N_24889,N_24517);
nand UO_1887 (O_1887,N_22725,N_23238);
nand UO_1888 (O_1888,N_24603,N_24989);
and UO_1889 (O_1889,N_23501,N_22660);
nand UO_1890 (O_1890,N_22802,N_24737);
and UO_1891 (O_1891,N_23437,N_22822);
nand UO_1892 (O_1892,N_23051,N_22674);
nand UO_1893 (O_1893,N_24894,N_23489);
nand UO_1894 (O_1894,N_22552,N_22976);
nand UO_1895 (O_1895,N_24502,N_24234);
nor UO_1896 (O_1896,N_23715,N_23992);
and UO_1897 (O_1897,N_22783,N_23860);
and UO_1898 (O_1898,N_22718,N_22905);
nor UO_1899 (O_1899,N_24640,N_24949);
and UO_1900 (O_1900,N_22671,N_24574);
nand UO_1901 (O_1901,N_22998,N_23086);
or UO_1902 (O_1902,N_24645,N_23411);
and UO_1903 (O_1903,N_24210,N_24336);
xnor UO_1904 (O_1904,N_24989,N_24016);
and UO_1905 (O_1905,N_23114,N_23911);
and UO_1906 (O_1906,N_23637,N_22668);
nand UO_1907 (O_1907,N_24375,N_23488);
nor UO_1908 (O_1908,N_22713,N_24653);
or UO_1909 (O_1909,N_23719,N_24988);
nor UO_1910 (O_1910,N_23115,N_23409);
nand UO_1911 (O_1911,N_23145,N_24033);
and UO_1912 (O_1912,N_23549,N_24189);
or UO_1913 (O_1913,N_23853,N_23425);
nor UO_1914 (O_1914,N_24664,N_24059);
nor UO_1915 (O_1915,N_23784,N_24250);
xnor UO_1916 (O_1916,N_23695,N_24123);
and UO_1917 (O_1917,N_24966,N_24812);
nor UO_1918 (O_1918,N_23522,N_24232);
nand UO_1919 (O_1919,N_24825,N_23778);
or UO_1920 (O_1920,N_23233,N_24674);
nand UO_1921 (O_1921,N_23685,N_23326);
or UO_1922 (O_1922,N_22988,N_23307);
nor UO_1923 (O_1923,N_23387,N_24086);
nor UO_1924 (O_1924,N_23057,N_23752);
or UO_1925 (O_1925,N_23293,N_23031);
xnor UO_1926 (O_1926,N_22545,N_24738);
xor UO_1927 (O_1927,N_24255,N_22958);
nor UO_1928 (O_1928,N_22837,N_24910);
xnor UO_1929 (O_1929,N_23411,N_22892);
nor UO_1930 (O_1930,N_24114,N_22525);
nand UO_1931 (O_1931,N_23162,N_23599);
or UO_1932 (O_1932,N_23713,N_24749);
nand UO_1933 (O_1933,N_23333,N_22929);
and UO_1934 (O_1934,N_23581,N_23328);
and UO_1935 (O_1935,N_23479,N_22721);
and UO_1936 (O_1936,N_22666,N_23086);
xor UO_1937 (O_1937,N_23499,N_24431);
xor UO_1938 (O_1938,N_22920,N_24074);
xor UO_1939 (O_1939,N_23142,N_23119);
nor UO_1940 (O_1940,N_23762,N_22575);
and UO_1941 (O_1941,N_22989,N_24166);
xor UO_1942 (O_1942,N_22544,N_22726);
or UO_1943 (O_1943,N_24292,N_22530);
nor UO_1944 (O_1944,N_22759,N_24847);
or UO_1945 (O_1945,N_24554,N_24758);
xor UO_1946 (O_1946,N_24204,N_23012);
nand UO_1947 (O_1947,N_23270,N_24119);
and UO_1948 (O_1948,N_23771,N_24365);
or UO_1949 (O_1949,N_24032,N_23574);
or UO_1950 (O_1950,N_24986,N_24470);
nor UO_1951 (O_1951,N_22930,N_22524);
nor UO_1952 (O_1952,N_23348,N_22504);
xnor UO_1953 (O_1953,N_24569,N_23794);
nand UO_1954 (O_1954,N_24550,N_24415);
or UO_1955 (O_1955,N_23992,N_24806);
or UO_1956 (O_1956,N_24105,N_23941);
and UO_1957 (O_1957,N_24076,N_22632);
and UO_1958 (O_1958,N_23770,N_23609);
and UO_1959 (O_1959,N_23912,N_23240);
and UO_1960 (O_1960,N_23065,N_22781);
xor UO_1961 (O_1961,N_22620,N_24020);
and UO_1962 (O_1962,N_24066,N_22920);
nor UO_1963 (O_1963,N_24890,N_24206);
xor UO_1964 (O_1964,N_23837,N_22892);
and UO_1965 (O_1965,N_24483,N_24028);
or UO_1966 (O_1966,N_23605,N_24276);
nor UO_1967 (O_1967,N_24403,N_24682);
nor UO_1968 (O_1968,N_23587,N_24432);
and UO_1969 (O_1969,N_23700,N_23708);
nor UO_1970 (O_1970,N_24190,N_24376);
and UO_1971 (O_1971,N_24856,N_24702);
xnor UO_1972 (O_1972,N_23920,N_22554);
or UO_1973 (O_1973,N_23165,N_23580);
nor UO_1974 (O_1974,N_24605,N_23563);
or UO_1975 (O_1975,N_24955,N_22574);
and UO_1976 (O_1976,N_23087,N_23755);
nor UO_1977 (O_1977,N_23612,N_23580);
nor UO_1978 (O_1978,N_24218,N_23966);
nor UO_1979 (O_1979,N_24494,N_22916);
nor UO_1980 (O_1980,N_24371,N_24167);
nand UO_1981 (O_1981,N_23872,N_23277);
nor UO_1982 (O_1982,N_22613,N_23483);
nor UO_1983 (O_1983,N_23675,N_23851);
nand UO_1984 (O_1984,N_22935,N_24690);
nor UO_1985 (O_1985,N_23948,N_24554);
nand UO_1986 (O_1986,N_23259,N_22808);
or UO_1987 (O_1987,N_23503,N_24198);
and UO_1988 (O_1988,N_23076,N_24630);
or UO_1989 (O_1989,N_24347,N_23334);
nand UO_1990 (O_1990,N_24751,N_23551);
xor UO_1991 (O_1991,N_23762,N_22694);
or UO_1992 (O_1992,N_23331,N_24354);
nor UO_1993 (O_1993,N_24976,N_24947);
nand UO_1994 (O_1994,N_24511,N_24694);
nor UO_1995 (O_1995,N_23570,N_22597);
nand UO_1996 (O_1996,N_23532,N_24334);
nor UO_1997 (O_1997,N_24215,N_23673);
nand UO_1998 (O_1998,N_22518,N_24356);
or UO_1999 (O_1999,N_24986,N_24200);
and UO_2000 (O_2000,N_23634,N_24386);
xnor UO_2001 (O_2001,N_24393,N_22760);
nor UO_2002 (O_2002,N_24805,N_24017);
and UO_2003 (O_2003,N_22811,N_22547);
nor UO_2004 (O_2004,N_24518,N_23767);
nand UO_2005 (O_2005,N_23490,N_24497);
nor UO_2006 (O_2006,N_24998,N_22906);
nor UO_2007 (O_2007,N_23113,N_24217);
or UO_2008 (O_2008,N_24910,N_24469);
xnor UO_2009 (O_2009,N_23817,N_23650);
and UO_2010 (O_2010,N_22800,N_22934);
or UO_2011 (O_2011,N_23078,N_23056);
nand UO_2012 (O_2012,N_24479,N_23567);
and UO_2013 (O_2013,N_23191,N_23123);
nand UO_2014 (O_2014,N_23460,N_24478);
xor UO_2015 (O_2015,N_23371,N_24617);
or UO_2016 (O_2016,N_24945,N_23365);
and UO_2017 (O_2017,N_22689,N_23748);
nand UO_2018 (O_2018,N_23027,N_23252);
or UO_2019 (O_2019,N_24841,N_23674);
nand UO_2020 (O_2020,N_24900,N_24753);
nor UO_2021 (O_2021,N_24221,N_24955);
nand UO_2022 (O_2022,N_24690,N_22697);
nand UO_2023 (O_2023,N_24022,N_22668);
xnor UO_2024 (O_2024,N_23283,N_23278);
nand UO_2025 (O_2025,N_22592,N_24586);
nand UO_2026 (O_2026,N_23544,N_23741);
or UO_2027 (O_2027,N_23517,N_22910);
xnor UO_2028 (O_2028,N_24005,N_24279);
and UO_2029 (O_2029,N_23324,N_23241);
xor UO_2030 (O_2030,N_24796,N_24399);
or UO_2031 (O_2031,N_24540,N_23848);
nand UO_2032 (O_2032,N_23242,N_24285);
nand UO_2033 (O_2033,N_22797,N_22501);
or UO_2034 (O_2034,N_24448,N_24672);
nor UO_2035 (O_2035,N_24572,N_24329);
and UO_2036 (O_2036,N_23633,N_22859);
nor UO_2037 (O_2037,N_24399,N_22914);
xor UO_2038 (O_2038,N_23739,N_24101);
nor UO_2039 (O_2039,N_24874,N_23877);
or UO_2040 (O_2040,N_23807,N_22824);
xnor UO_2041 (O_2041,N_23366,N_23169);
or UO_2042 (O_2042,N_23223,N_23367);
or UO_2043 (O_2043,N_24717,N_22853);
xnor UO_2044 (O_2044,N_24147,N_23405);
nor UO_2045 (O_2045,N_24302,N_22662);
nand UO_2046 (O_2046,N_24768,N_23747);
and UO_2047 (O_2047,N_23794,N_23212);
nor UO_2048 (O_2048,N_24531,N_23880);
nand UO_2049 (O_2049,N_24801,N_23388);
or UO_2050 (O_2050,N_24765,N_23888);
or UO_2051 (O_2051,N_23711,N_23505);
nand UO_2052 (O_2052,N_23188,N_23192);
nand UO_2053 (O_2053,N_24097,N_22696);
xor UO_2054 (O_2054,N_24373,N_23122);
nor UO_2055 (O_2055,N_23510,N_22819);
nor UO_2056 (O_2056,N_23542,N_23570);
nand UO_2057 (O_2057,N_22653,N_22830);
or UO_2058 (O_2058,N_22530,N_23590);
and UO_2059 (O_2059,N_23147,N_23071);
and UO_2060 (O_2060,N_23389,N_22993);
and UO_2061 (O_2061,N_23284,N_24455);
nand UO_2062 (O_2062,N_24015,N_22544);
nand UO_2063 (O_2063,N_22726,N_22909);
xnor UO_2064 (O_2064,N_22795,N_23782);
nand UO_2065 (O_2065,N_24158,N_24230);
nor UO_2066 (O_2066,N_23574,N_23193);
and UO_2067 (O_2067,N_24854,N_24981);
nand UO_2068 (O_2068,N_22931,N_24096);
and UO_2069 (O_2069,N_22673,N_24930);
xnor UO_2070 (O_2070,N_23267,N_23395);
nand UO_2071 (O_2071,N_23090,N_24160);
nand UO_2072 (O_2072,N_24601,N_24903);
and UO_2073 (O_2073,N_23792,N_23073);
and UO_2074 (O_2074,N_23651,N_22513);
or UO_2075 (O_2075,N_23260,N_24748);
nand UO_2076 (O_2076,N_24064,N_22717);
nand UO_2077 (O_2077,N_24622,N_22966);
nand UO_2078 (O_2078,N_22744,N_23198);
nand UO_2079 (O_2079,N_22902,N_24450);
and UO_2080 (O_2080,N_24568,N_24986);
xor UO_2081 (O_2081,N_24016,N_23503);
xnor UO_2082 (O_2082,N_23663,N_22914);
nor UO_2083 (O_2083,N_24330,N_24556);
or UO_2084 (O_2084,N_23971,N_24204);
xnor UO_2085 (O_2085,N_22793,N_23500);
and UO_2086 (O_2086,N_23587,N_23628);
or UO_2087 (O_2087,N_24352,N_23700);
or UO_2088 (O_2088,N_24798,N_23039);
nand UO_2089 (O_2089,N_23081,N_24087);
xor UO_2090 (O_2090,N_23768,N_23610);
xor UO_2091 (O_2091,N_23629,N_24335);
nand UO_2092 (O_2092,N_23720,N_24566);
nand UO_2093 (O_2093,N_23812,N_24437);
nor UO_2094 (O_2094,N_23749,N_24120);
xnor UO_2095 (O_2095,N_23727,N_24512);
xnor UO_2096 (O_2096,N_23692,N_24526);
nor UO_2097 (O_2097,N_22576,N_23913);
xnor UO_2098 (O_2098,N_23768,N_22977);
nor UO_2099 (O_2099,N_24404,N_23404);
and UO_2100 (O_2100,N_23149,N_24050);
or UO_2101 (O_2101,N_23810,N_24827);
or UO_2102 (O_2102,N_23140,N_23549);
xor UO_2103 (O_2103,N_22656,N_24569);
nand UO_2104 (O_2104,N_22625,N_24471);
or UO_2105 (O_2105,N_23141,N_23777);
nand UO_2106 (O_2106,N_24870,N_23493);
nand UO_2107 (O_2107,N_24745,N_24561);
nand UO_2108 (O_2108,N_24149,N_22812);
or UO_2109 (O_2109,N_23570,N_23451);
nor UO_2110 (O_2110,N_24051,N_24187);
nand UO_2111 (O_2111,N_23292,N_24696);
or UO_2112 (O_2112,N_24014,N_22591);
or UO_2113 (O_2113,N_24828,N_24580);
and UO_2114 (O_2114,N_23189,N_24242);
xor UO_2115 (O_2115,N_22665,N_22659);
nand UO_2116 (O_2116,N_24037,N_22636);
xor UO_2117 (O_2117,N_24004,N_23530);
and UO_2118 (O_2118,N_22563,N_24348);
or UO_2119 (O_2119,N_24293,N_24225);
and UO_2120 (O_2120,N_22772,N_24254);
nor UO_2121 (O_2121,N_24963,N_24697);
and UO_2122 (O_2122,N_24429,N_22918);
and UO_2123 (O_2123,N_22632,N_22770);
xor UO_2124 (O_2124,N_24816,N_24872);
xor UO_2125 (O_2125,N_23215,N_24858);
xor UO_2126 (O_2126,N_23222,N_24723);
nor UO_2127 (O_2127,N_24035,N_22561);
and UO_2128 (O_2128,N_22762,N_23551);
xor UO_2129 (O_2129,N_23618,N_22729);
nand UO_2130 (O_2130,N_23194,N_22588);
nor UO_2131 (O_2131,N_23207,N_22564);
nand UO_2132 (O_2132,N_23560,N_23072);
xnor UO_2133 (O_2133,N_24204,N_23807);
xor UO_2134 (O_2134,N_24945,N_22579);
nand UO_2135 (O_2135,N_23002,N_23313);
or UO_2136 (O_2136,N_22837,N_23493);
xor UO_2137 (O_2137,N_24879,N_24975);
and UO_2138 (O_2138,N_24432,N_24664);
nand UO_2139 (O_2139,N_23727,N_22503);
nor UO_2140 (O_2140,N_23140,N_22926);
nor UO_2141 (O_2141,N_24796,N_22983);
nand UO_2142 (O_2142,N_23612,N_24847);
nand UO_2143 (O_2143,N_23582,N_22641);
nor UO_2144 (O_2144,N_23339,N_24403);
nand UO_2145 (O_2145,N_24839,N_23807);
nand UO_2146 (O_2146,N_24666,N_24117);
xnor UO_2147 (O_2147,N_24812,N_22788);
xnor UO_2148 (O_2148,N_24660,N_22848);
nand UO_2149 (O_2149,N_24597,N_24045);
or UO_2150 (O_2150,N_22944,N_22698);
and UO_2151 (O_2151,N_23967,N_23653);
nor UO_2152 (O_2152,N_24748,N_23775);
or UO_2153 (O_2153,N_24895,N_23717);
xnor UO_2154 (O_2154,N_24119,N_23574);
nor UO_2155 (O_2155,N_24678,N_23271);
nor UO_2156 (O_2156,N_22598,N_22653);
nand UO_2157 (O_2157,N_24653,N_23525);
xnor UO_2158 (O_2158,N_23242,N_24139);
and UO_2159 (O_2159,N_22536,N_24175);
or UO_2160 (O_2160,N_24095,N_22692);
nand UO_2161 (O_2161,N_23241,N_22670);
nand UO_2162 (O_2162,N_24090,N_24867);
or UO_2163 (O_2163,N_22556,N_23377);
nor UO_2164 (O_2164,N_23820,N_24514);
and UO_2165 (O_2165,N_24721,N_23389);
nor UO_2166 (O_2166,N_24607,N_22522);
or UO_2167 (O_2167,N_22659,N_23789);
nand UO_2168 (O_2168,N_24662,N_24529);
and UO_2169 (O_2169,N_24166,N_23645);
nor UO_2170 (O_2170,N_22647,N_24282);
nand UO_2171 (O_2171,N_23764,N_22503);
or UO_2172 (O_2172,N_22616,N_24127);
and UO_2173 (O_2173,N_23236,N_23146);
xnor UO_2174 (O_2174,N_23001,N_23721);
nor UO_2175 (O_2175,N_22871,N_23342);
xnor UO_2176 (O_2176,N_22921,N_22729);
xor UO_2177 (O_2177,N_23541,N_23392);
and UO_2178 (O_2178,N_22935,N_23782);
nand UO_2179 (O_2179,N_24209,N_23775);
nand UO_2180 (O_2180,N_23005,N_23869);
or UO_2181 (O_2181,N_24958,N_24680);
xnor UO_2182 (O_2182,N_23078,N_24059);
xnor UO_2183 (O_2183,N_23185,N_23428);
nand UO_2184 (O_2184,N_23559,N_22770);
and UO_2185 (O_2185,N_23104,N_24774);
and UO_2186 (O_2186,N_24113,N_23736);
nand UO_2187 (O_2187,N_22815,N_24741);
nand UO_2188 (O_2188,N_24463,N_24013);
xor UO_2189 (O_2189,N_24861,N_24449);
nor UO_2190 (O_2190,N_24577,N_22830);
or UO_2191 (O_2191,N_22740,N_22704);
and UO_2192 (O_2192,N_23616,N_24954);
or UO_2193 (O_2193,N_24234,N_22511);
and UO_2194 (O_2194,N_23589,N_23868);
nor UO_2195 (O_2195,N_22779,N_22519);
nand UO_2196 (O_2196,N_22753,N_24966);
and UO_2197 (O_2197,N_24223,N_24365);
xor UO_2198 (O_2198,N_23414,N_24703);
nor UO_2199 (O_2199,N_23530,N_22903);
nor UO_2200 (O_2200,N_23078,N_23346);
xor UO_2201 (O_2201,N_23141,N_23102);
xor UO_2202 (O_2202,N_23607,N_22957);
and UO_2203 (O_2203,N_24129,N_22930);
and UO_2204 (O_2204,N_24957,N_22541);
xnor UO_2205 (O_2205,N_23198,N_24233);
xnor UO_2206 (O_2206,N_23639,N_23141);
xnor UO_2207 (O_2207,N_24300,N_22636);
nor UO_2208 (O_2208,N_24306,N_24973);
or UO_2209 (O_2209,N_24111,N_23807);
nand UO_2210 (O_2210,N_23741,N_24687);
and UO_2211 (O_2211,N_23536,N_23791);
or UO_2212 (O_2212,N_22549,N_23441);
nand UO_2213 (O_2213,N_23461,N_23674);
and UO_2214 (O_2214,N_24681,N_23117);
xnor UO_2215 (O_2215,N_24518,N_23766);
xnor UO_2216 (O_2216,N_23705,N_22811);
nand UO_2217 (O_2217,N_23747,N_22800);
nand UO_2218 (O_2218,N_22965,N_23033);
or UO_2219 (O_2219,N_23014,N_23850);
nor UO_2220 (O_2220,N_22690,N_24079);
nand UO_2221 (O_2221,N_23318,N_24889);
nand UO_2222 (O_2222,N_24068,N_22677);
and UO_2223 (O_2223,N_24727,N_22625);
xor UO_2224 (O_2224,N_23791,N_24810);
xor UO_2225 (O_2225,N_24364,N_24208);
or UO_2226 (O_2226,N_23792,N_23820);
xor UO_2227 (O_2227,N_23883,N_24270);
xor UO_2228 (O_2228,N_22780,N_24850);
or UO_2229 (O_2229,N_23929,N_24895);
xor UO_2230 (O_2230,N_24638,N_23149);
or UO_2231 (O_2231,N_23540,N_24003);
nand UO_2232 (O_2232,N_24084,N_24396);
and UO_2233 (O_2233,N_24634,N_24482);
or UO_2234 (O_2234,N_23648,N_24751);
nand UO_2235 (O_2235,N_23294,N_24887);
nand UO_2236 (O_2236,N_23519,N_23971);
and UO_2237 (O_2237,N_24928,N_23659);
nor UO_2238 (O_2238,N_22764,N_24231);
and UO_2239 (O_2239,N_23396,N_24634);
and UO_2240 (O_2240,N_22812,N_24473);
and UO_2241 (O_2241,N_24485,N_23809);
or UO_2242 (O_2242,N_24076,N_24687);
and UO_2243 (O_2243,N_24071,N_23316);
nor UO_2244 (O_2244,N_22537,N_22906);
nor UO_2245 (O_2245,N_24084,N_24432);
nor UO_2246 (O_2246,N_23235,N_24619);
xnor UO_2247 (O_2247,N_23120,N_23144);
and UO_2248 (O_2248,N_23095,N_22941);
nand UO_2249 (O_2249,N_23671,N_23892);
nand UO_2250 (O_2250,N_24637,N_24523);
and UO_2251 (O_2251,N_23760,N_24334);
nand UO_2252 (O_2252,N_22637,N_24169);
nand UO_2253 (O_2253,N_23550,N_24348);
and UO_2254 (O_2254,N_22699,N_22941);
or UO_2255 (O_2255,N_23717,N_22507);
nand UO_2256 (O_2256,N_24632,N_23283);
nor UO_2257 (O_2257,N_23073,N_22595);
nor UO_2258 (O_2258,N_24297,N_24324);
xnor UO_2259 (O_2259,N_23463,N_24386);
or UO_2260 (O_2260,N_23386,N_24664);
nand UO_2261 (O_2261,N_24100,N_23988);
nand UO_2262 (O_2262,N_23677,N_22830);
nor UO_2263 (O_2263,N_24377,N_24454);
nor UO_2264 (O_2264,N_23925,N_23407);
nand UO_2265 (O_2265,N_23308,N_23253);
nor UO_2266 (O_2266,N_24633,N_22502);
or UO_2267 (O_2267,N_22740,N_24956);
xnor UO_2268 (O_2268,N_23107,N_23241);
and UO_2269 (O_2269,N_24573,N_23370);
or UO_2270 (O_2270,N_22898,N_22890);
nor UO_2271 (O_2271,N_22580,N_23741);
nor UO_2272 (O_2272,N_23902,N_24016);
or UO_2273 (O_2273,N_23284,N_23645);
nor UO_2274 (O_2274,N_22993,N_24392);
or UO_2275 (O_2275,N_22813,N_24966);
and UO_2276 (O_2276,N_23316,N_24058);
nand UO_2277 (O_2277,N_24081,N_24158);
nand UO_2278 (O_2278,N_22718,N_22714);
or UO_2279 (O_2279,N_23134,N_23873);
nor UO_2280 (O_2280,N_22741,N_24217);
xnor UO_2281 (O_2281,N_24016,N_23605);
nor UO_2282 (O_2282,N_22917,N_24700);
xnor UO_2283 (O_2283,N_24773,N_23623);
or UO_2284 (O_2284,N_23336,N_22608);
or UO_2285 (O_2285,N_24416,N_22993);
nor UO_2286 (O_2286,N_24811,N_24438);
nand UO_2287 (O_2287,N_23820,N_24695);
nor UO_2288 (O_2288,N_24548,N_23120);
nor UO_2289 (O_2289,N_22941,N_24195);
or UO_2290 (O_2290,N_24217,N_23310);
nand UO_2291 (O_2291,N_22742,N_24220);
or UO_2292 (O_2292,N_22788,N_23748);
and UO_2293 (O_2293,N_24148,N_23176);
and UO_2294 (O_2294,N_23781,N_22968);
nand UO_2295 (O_2295,N_23161,N_24985);
nand UO_2296 (O_2296,N_24234,N_23785);
or UO_2297 (O_2297,N_23173,N_23764);
nor UO_2298 (O_2298,N_23450,N_24203);
nand UO_2299 (O_2299,N_23061,N_22704);
nand UO_2300 (O_2300,N_22994,N_23024);
and UO_2301 (O_2301,N_23256,N_24918);
and UO_2302 (O_2302,N_23990,N_23635);
xnor UO_2303 (O_2303,N_23443,N_24125);
or UO_2304 (O_2304,N_24921,N_24997);
nor UO_2305 (O_2305,N_23025,N_23731);
nor UO_2306 (O_2306,N_24803,N_23910);
or UO_2307 (O_2307,N_23080,N_24653);
xnor UO_2308 (O_2308,N_24709,N_24013);
nand UO_2309 (O_2309,N_24414,N_24261);
nor UO_2310 (O_2310,N_23210,N_23266);
nor UO_2311 (O_2311,N_24183,N_22556);
nand UO_2312 (O_2312,N_23397,N_23654);
nor UO_2313 (O_2313,N_22921,N_22786);
and UO_2314 (O_2314,N_24753,N_23258);
xor UO_2315 (O_2315,N_24425,N_23773);
nand UO_2316 (O_2316,N_22737,N_22572);
nand UO_2317 (O_2317,N_24544,N_23722);
or UO_2318 (O_2318,N_23793,N_23726);
and UO_2319 (O_2319,N_24206,N_24545);
xnor UO_2320 (O_2320,N_24804,N_23932);
or UO_2321 (O_2321,N_24262,N_23804);
nand UO_2322 (O_2322,N_22851,N_24711);
nor UO_2323 (O_2323,N_24527,N_24384);
or UO_2324 (O_2324,N_24782,N_23396);
or UO_2325 (O_2325,N_23276,N_23287);
nor UO_2326 (O_2326,N_23174,N_22774);
and UO_2327 (O_2327,N_24672,N_24089);
xor UO_2328 (O_2328,N_24977,N_24675);
nand UO_2329 (O_2329,N_23306,N_24922);
nor UO_2330 (O_2330,N_23566,N_24842);
nand UO_2331 (O_2331,N_23954,N_24565);
nor UO_2332 (O_2332,N_23367,N_23189);
nor UO_2333 (O_2333,N_24389,N_24950);
xnor UO_2334 (O_2334,N_22816,N_23939);
nand UO_2335 (O_2335,N_23869,N_23902);
xor UO_2336 (O_2336,N_24549,N_24623);
and UO_2337 (O_2337,N_23641,N_23188);
or UO_2338 (O_2338,N_24434,N_24789);
xor UO_2339 (O_2339,N_24717,N_22903);
nand UO_2340 (O_2340,N_22603,N_24064);
and UO_2341 (O_2341,N_23819,N_24391);
nor UO_2342 (O_2342,N_24150,N_23490);
xnor UO_2343 (O_2343,N_24584,N_24513);
and UO_2344 (O_2344,N_24322,N_24376);
nor UO_2345 (O_2345,N_24126,N_22919);
and UO_2346 (O_2346,N_24445,N_23794);
and UO_2347 (O_2347,N_23334,N_23006);
nand UO_2348 (O_2348,N_24162,N_24776);
and UO_2349 (O_2349,N_22683,N_22970);
nand UO_2350 (O_2350,N_24384,N_24557);
or UO_2351 (O_2351,N_22671,N_23404);
xnor UO_2352 (O_2352,N_22906,N_24761);
and UO_2353 (O_2353,N_24263,N_22826);
and UO_2354 (O_2354,N_24818,N_24965);
or UO_2355 (O_2355,N_24061,N_24521);
and UO_2356 (O_2356,N_22663,N_22634);
and UO_2357 (O_2357,N_24702,N_24766);
or UO_2358 (O_2358,N_22502,N_22693);
xor UO_2359 (O_2359,N_23391,N_22979);
or UO_2360 (O_2360,N_23250,N_23607);
and UO_2361 (O_2361,N_23056,N_23896);
nand UO_2362 (O_2362,N_24963,N_23816);
nand UO_2363 (O_2363,N_23299,N_23699);
nor UO_2364 (O_2364,N_24335,N_23486);
xor UO_2365 (O_2365,N_23825,N_23451);
nand UO_2366 (O_2366,N_23734,N_23718);
and UO_2367 (O_2367,N_24098,N_23478);
xnor UO_2368 (O_2368,N_24211,N_24537);
nand UO_2369 (O_2369,N_22631,N_23497);
xnor UO_2370 (O_2370,N_23662,N_23554);
and UO_2371 (O_2371,N_23291,N_22626);
nand UO_2372 (O_2372,N_24316,N_24669);
nand UO_2373 (O_2373,N_24665,N_24506);
nor UO_2374 (O_2374,N_24223,N_23884);
and UO_2375 (O_2375,N_22889,N_24477);
and UO_2376 (O_2376,N_23027,N_24734);
nor UO_2377 (O_2377,N_23624,N_24209);
and UO_2378 (O_2378,N_24221,N_24262);
and UO_2379 (O_2379,N_23663,N_23899);
xor UO_2380 (O_2380,N_24496,N_24664);
and UO_2381 (O_2381,N_24222,N_24610);
and UO_2382 (O_2382,N_24480,N_23398);
nor UO_2383 (O_2383,N_23333,N_22766);
nand UO_2384 (O_2384,N_24852,N_23541);
or UO_2385 (O_2385,N_22713,N_22538);
nand UO_2386 (O_2386,N_24531,N_23108);
xnor UO_2387 (O_2387,N_23152,N_22600);
and UO_2388 (O_2388,N_23919,N_23807);
xnor UO_2389 (O_2389,N_24451,N_22726);
nor UO_2390 (O_2390,N_23921,N_23680);
and UO_2391 (O_2391,N_22561,N_23021);
nor UO_2392 (O_2392,N_22572,N_23650);
nor UO_2393 (O_2393,N_22804,N_23897);
xor UO_2394 (O_2394,N_24554,N_23552);
nand UO_2395 (O_2395,N_23705,N_24234);
xor UO_2396 (O_2396,N_23629,N_23458);
xnor UO_2397 (O_2397,N_23857,N_22842);
nand UO_2398 (O_2398,N_22762,N_22889);
nand UO_2399 (O_2399,N_24853,N_23862);
xor UO_2400 (O_2400,N_24978,N_24460);
nand UO_2401 (O_2401,N_22575,N_23575);
xnor UO_2402 (O_2402,N_23951,N_22906);
nor UO_2403 (O_2403,N_24438,N_22547);
and UO_2404 (O_2404,N_23507,N_22796);
and UO_2405 (O_2405,N_24625,N_24226);
nor UO_2406 (O_2406,N_23778,N_22827);
nor UO_2407 (O_2407,N_23415,N_22683);
nand UO_2408 (O_2408,N_22912,N_24615);
or UO_2409 (O_2409,N_24898,N_23682);
nor UO_2410 (O_2410,N_23781,N_24143);
and UO_2411 (O_2411,N_23767,N_24147);
nor UO_2412 (O_2412,N_23184,N_24154);
nand UO_2413 (O_2413,N_22689,N_22648);
xnor UO_2414 (O_2414,N_22830,N_22546);
or UO_2415 (O_2415,N_23111,N_24537);
or UO_2416 (O_2416,N_24230,N_23616);
nand UO_2417 (O_2417,N_23991,N_23994);
nor UO_2418 (O_2418,N_23368,N_23616);
nand UO_2419 (O_2419,N_23024,N_23258);
or UO_2420 (O_2420,N_23314,N_24478);
or UO_2421 (O_2421,N_24389,N_23392);
xnor UO_2422 (O_2422,N_23973,N_23050);
xor UO_2423 (O_2423,N_23100,N_23660);
and UO_2424 (O_2424,N_23154,N_23804);
nor UO_2425 (O_2425,N_23458,N_23069);
nor UO_2426 (O_2426,N_22756,N_24948);
nand UO_2427 (O_2427,N_24318,N_24182);
nand UO_2428 (O_2428,N_23669,N_24839);
and UO_2429 (O_2429,N_23984,N_24183);
nor UO_2430 (O_2430,N_24637,N_24879);
nand UO_2431 (O_2431,N_23767,N_24996);
nor UO_2432 (O_2432,N_24354,N_22865);
nand UO_2433 (O_2433,N_23512,N_23164);
nor UO_2434 (O_2434,N_22937,N_23236);
nand UO_2435 (O_2435,N_23210,N_24035);
or UO_2436 (O_2436,N_23139,N_24498);
or UO_2437 (O_2437,N_24248,N_24643);
or UO_2438 (O_2438,N_24813,N_24043);
nor UO_2439 (O_2439,N_23413,N_24505);
and UO_2440 (O_2440,N_22685,N_24266);
and UO_2441 (O_2441,N_22507,N_24201);
nor UO_2442 (O_2442,N_22857,N_24483);
xor UO_2443 (O_2443,N_23195,N_24503);
nor UO_2444 (O_2444,N_24647,N_24255);
and UO_2445 (O_2445,N_23326,N_23076);
and UO_2446 (O_2446,N_23883,N_22973);
and UO_2447 (O_2447,N_23211,N_23897);
xnor UO_2448 (O_2448,N_23466,N_24681);
nor UO_2449 (O_2449,N_23454,N_23517);
nor UO_2450 (O_2450,N_24091,N_23720);
and UO_2451 (O_2451,N_24369,N_23478);
and UO_2452 (O_2452,N_24224,N_23037);
nand UO_2453 (O_2453,N_22985,N_23859);
nor UO_2454 (O_2454,N_24370,N_22626);
nand UO_2455 (O_2455,N_24871,N_23815);
nor UO_2456 (O_2456,N_23119,N_24360);
xnor UO_2457 (O_2457,N_24789,N_23503);
or UO_2458 (O_2458,N_22860,N_22924);
or UO_2459 (O_2459,N_23730,N_24249);
nor UO_2460 (O_2460,N_22535,N_24332);
nor UO_2461 (O_2461,N_24380,N_24055);
and UO_2462 (O_2462,N_24263,N_24636);
nor UO_2463 (O_2463,N_24547,N_23789);
xnor UO_2464 (O_2464,N_23479,N_23223);
nand UO_2465 (O_2465,N_23416,N_24144);
and UO_2466 (O_2466,N_24600,N_24652);
or UO_2467 (O_2467,N_23105,N_23596);
and UO_2468 (O_2468,N_24319,N_22613);
nand UO_2469 (O_2469,N_23698,N_22598);
nor UO_2470 (O_2470,N_24463,N_22739);
xnor UO_2471 (O_2471,N_23736,N_22890);
nor UO_2472 (O_2472,N_23383,N_24650);
xor UO_2473 (O_2473,N_23907,N_23353);
or UO_2474 (O_2474,N_23595,N_23130);
and UO_2475 (O_2475,N_22906,N_24637);
or UO_2476 (O_2476,N_24420,N_23405);
nand UO_2477 (O_2477,N_24714,N_23066);
xnor UO_2478 (O_2478,N_24980,N_23236);
nand UO_2479 (O_2479,N_23944,N_22837);
or UO_2480 (O_2480,N_24090,N_24737);
nand UO_2481 (O_2481,N_24124,N_23497);
or UO_2482 (O_2482,N_22713,N_24796);
or UO_2483 (O_2483,N_24591,N_24065);
nor UO_2484 (O_2484,N_24739,N_23595);
xnor UO_2485 (O_2485,N_22962,N_24978);
nand UO_2486 (O_2486,N_24881,N_23808);
xnor UO_2487 (O_2487,N_24142,N_22517);
xnor UO_2488 (O_2488,N_22631,N_24848);
xor UO_2489 (O_2489,N_24349,N_22715);
or UO_2490 (O_2490,N_24114,N_23176);
and UO_2491 (O_2491,N_23197,N_23647);
or UO_2492 (O_2492,N_24245,N_24410);
or UO_2493 (O_2493,N_24391,N_22975);
nor UO_2494 (O_2494,N_24065,N_24949);
nor UO_2495 (O_2495,N_23554,N_22988);
nor UO_2496 (O_2496,N_24353,N_24692);
nand UO_2497 (O_2497,N_23564,N_23565);
and UO_2498 (O_2498,N_23998,N_23673);
nand UO_2499 (O_2499,N_24521,N_22975);
xor UO_2500 (O_2500,N_23103,N_23173);
or UO_2501 (O_2501,N_24583,N_22929);
nor UO_2502 (O_2502,N_24851,N_24075);
xnor UO_2503 (O_2503,N_23802,N_24656);
or UO_2504 (O_2504,N_23291,N_23031);
nand UO_2505 (O_2505,N_24157,N_24584);
or UO_2506 (O_2506,N_24053,N_24036);
nor UO_2507 (O_2507,N_23093,N_23068);
nor UO_2508 (O_2508,N_22899,N_22991);
xor UO_2509 (O_2509,N_22649,N_24550);
or UO_2510 (O_2510,N_22741,N_24345);
xnor UO_2511 (O_2511,N_24596,N_24723);
xnor UO_2512 (O_2512,N_23647,N_23250);
nor UO_2513 (O_2513,N_24065,N_23587);
or UO_2514 (O_2514,N_23404,N_23686);
nor UO_2515 (O_2515,N_24256,N_24210);
or UO_2516 (O_2516,N_24587,N_22874);
nor UO_2517 (O_2517,N_22839,N_24543);
xnor UO_2518 (O_2518,N_24268,N_24149);
xor UO_2519 (O_2519,N_24879,N_23871);
nor UO_2520 (O_2520,N_23455,N_22608);
or UO_2521 (O_2521,N_23850,N_22631);
nor UO_2522 (O_2522,N_22528,N_23226);
xnor UO_2523 (O_2523,N_24241,N_23555);
nor UO_2524 (O_2524,N_24881,N_23854);
nor UO_2525 (O_2525,N_23845,N_24671);
nor UO_2526 (O_2526,N_23549,N_22992);
and UO_2527 (O_2527,N_23322,N_23807);
nor UO_2528 (O_2528,N_23938,N_23496);
and UO_2529 (O_2529,N_22558,N_22792);
or UO_2530 (O_2530,N_23785,N_24473);
nand UO_2531 (O_2531,N_24700,N_24694);
xor UO_2532 (O_2532,N_24469,N_24483);
nor UO_2533 (O_2533,N_24045,N_22882);
or UO_2534 (O_2534,N_22550,N_24935);
and UO_2535 (O_2535,N_22545,N_22758);
or UO_2536 (O_2536,N_23759,N_23130);
xor UO_2537 (O_2537,N_23291,N_23647);
nor UO_2538 (O_2538,N_24366,N_24710);
and UO_2539 (O_2539,N_22820,N_23232);
nand UO_2540 (O_2540,N_23531,N_22622);
nand UO_2541 (O_2541,N_24465,N_24109);
nand UO_2542 (O_2542,N_24725,N_24381);
xnor UO_2543 (O_2543,N_23829,N_23904);
nand UO_2544 (O_2544,N_24435,N_24144);
nor UO_2545 (O_2545,N_23393,N_24568);
and UO_2546 (O_2546,N_24488,N_23071);
nand UO_2547 (O_2547,N_24371,N_24762);
xnor UO_2548 (O_2548,N_24569,N_23885);
xnor UO_2549 (O_2549,N_24330,N_24509);
nand UO_2550 (O_2550,N_22554,N_23956);
or UO_2551 (O_2551,N_24657,N_24341);
nand UO_2552 (O_2552,N_24447,N_23248);
nand UO_2553 (O_2553,N_23114,N_24618);
or UO_2554 (O_2554,N_23807,N_24509);
xnor UO_2555 (O_2555,N_23106,N_23374);
xnor UO_2556 (O_2556,N_23538,N_22930);
nor UO_2557 (O_2557,N_23870,N_22895);
nand UO_2558 (O_2558,N_23301,N_23926);
nor UO_2559 (O_2559,N_23365,N_23705);
nor UO_2560 (O_2560,N_24612,N_24328);
xor UO_2561 (O_2561,N_22936,N_22783);
nor UO_2562 (O_2562,N_22982,N_24861);
nand UO_2563 (O_2563,N_24341,N_23051);
or UO_2564 (O_2564,N_24526,N_23099);
or UO_2565 (O_2565,N_23085,N_23394);
nor UO_2566 (O_2566,N_22750,N_23255);
xnor UO_2567 (O_2567,N_24052,N_22591);
or UO_2568 (O_2568,N_23976,N_24105);
nand UO_2569 (O_2569,N_22619,N_23653);
nand UO_2570 (O_2570,N_23106,N_24592);
nand UO_2571 (O_2571,N_24727,N_23939);
or UO_2572 (O_2572,N_23672,N_24510);
or UO_2573 (O_2573,N_24505,N_22934);
nor UO_2574 (O_2574,N_23435,N_22978);
or UO_2575 (O_2575,N_23857,N_23577);
and UO_2576 (O_2576,N_24318,N_23801);
nand UO_2577 (O_2577,N_24022,N_24494);
nand UO_2578 (O_2578,N_24081,N_24670);
nor UO_2579 (O_2579,N_23448,N_24952);
and UO_2580 (O_2580,N_22816,N_22697);
xor UO_2581 (O_2581,N_23490,N_23390);
nor UO_2582 (O_2582,N_22606,N_23765);
nor UO_2583 (O_2583,N_23085,N_23827);
or UO_2584 (O_2584,N_24191,N_23364);
xor UO_2585 (O_2585,N_23146,N_23100);
nor UO_2586 (O_2586,N_23337,N_23098);
nand UO_2587 (O_2587,N_23372,N_22823);
xnor UO_2588 (O_2588,N_24017,N_24800);
nand UO_2589 (O_2589,N_24117,N_23940);
xnor UO_2590 (O_2590,N_24632,N_23858);
xnor UO_2591 (O_2591,N_22858,N_23120);
nor UO_2592 (O_2592,N_24407,N_22748);
or UO_2593 (O_2593,N_24793,N_22531);
nand UO_2594 (O_2594,N_23506,N_23004);
or UO_2595 (O_2595,N_22707,N_23229);
and UO_2596 (O_2596,N_24897,N_22583);
and UO_2597 (O_2597,N_23269,N_24677);
nor UO_2598 (O_2598,N_24536,N_24885);
xnor UO_2599 (O_2599,N_23886,N_24252);
or UO_2600 (O_2600,N_24981,N_23781);
and UO_2601 (O_2601,N_23154,N_24741);
xor UO_2602 (O_2602,N_23480,N_24419);
nor UO_2603 (O_2603,N_23513,N_23042);
xor UO_2604 (O_2604,N_24341,N_24876);
xor UO_2605 (O_2605,N_22721,N_24949);
nand UO_2606 (O_2606,N_23901,N_23791);
nor UO_2607 (O_2607,N_23484,N_24604);
nor UO_2608 (O_2608,N_24335,N_24597);
nand UO_2609 (O_2609,N_24518,N_24995);
and UO_2610 (O_2610,N_23542,N_23683);
nor UO_2611 (O_2611,N_24451,N_23579);
or UO_2612 (O_2612,N_24895,N_24364);
nor UO_2613 (O_2613,N_23491,N_24091);
nor UO_2614 (O_2614,N_23172,N_22687);
nor UO_2615 (O_2615,N_23165,N_24152);
nor UO_2616 (O_2616,N_23926,N_24590);
xor UO_2617 (O_2617,N_24210,N_24369);
and UO_2618 (O_2618,N_22937,N_22579);
xor UO_2619 (O_2619,N_24910,N_23371);
and UO_2620 (O_2620,N_24859,N_23070);
and UO_2621 (O_2621,N_23285,N_23921);
nand UO_2622 (O_2622,N_24849,N_23121);
nor UO_2623 (O_2623,N_24896,N_22616);
or UO_2624 (O_2624,N_23417,N_22647);
and UO_2625 (O_2625,N_24310,N_22606);
or UO_2626 (O_2626,N_24849,N_24484);
nor UO_2627 (O_2627,N_22904,N_23460);
or UO_2628 (O_2628,N_23811,N_24586);
nand UO_2629 (O_2629,N_24473,N_23237);
or UO_2630 (O_2630,N_24125,N_24658);
nand UO_2631 (O_2631,N_24313,N_24969);
nand UO_2632 (O_2632,N_24472,N_23212);
and UO_2633 (O_2633,N_24080,N_23924);
nand UO_2634 (O_2634,N_24624,N_23192);
xor UO_2635 (O_2635,N_24853,N_22845);
xor UO_2636 (O_2636,N_24243,N_23417);
and UO_2637 (O_2637,N_22945,N_22746);
nor UO_2638 (O_2638,N_24953,N_23861);
and UO_2639 (O_2639,N_24252,N_22620);
xnor UO_2640 (O_2640,N_22986,N_23016);
nor UO_2641 (O_2641,N_24338,N_23974);
nor UO_2642 (O_2642,N_23364,N_23247);
nand UO_2643 (O_2643,N_24817,N_22647);
nor UO_2644 (O_2644,N_22792,N_24741);
or UO_2645 (O_2645,N_24597,N_24453);
nor UO_2646 (O_2646,N_24971,N_22863);
xor UO_2647 (O_2647,N_23414,N_23516);
or UO_2648 (O_2648,N_24192,N_24353);
nor UO_2649 (O_2649,N_22657,N_22645);
and UO_2650 (O_2650,N_22636,N_24347);
nor UO_2651 (O_2651,N_24759,N_22782);
nand UO_2652 (O_2652,N_24811,N_23346);
and UO_2653 (O_2653,N_22871,N_23048);
nand UO_2654 (O_2654,N_24013,N_22683);
and UO_2655 (O_2655,N_24562,N_24171);
nand UO_2656 (O_2656,N_22967,N_24510);
or UO_2657 (O_2657,N_22848,N_23693);
nor UO_2658 (O_2658,N_24684,N_22572);
nor UO_2659 (O_2659,N_23450,N_24490);
nand UO_2660 (O_2660,N_24000,N_23285);
xnor UO_2661 (O_2661,N_23885,N_24259);
and UO_2662 (O_2662,N_24299,N_22817);
and UO_2663 (O_2663,N_24966,N_24927);
and UO_2664 (O_2664,N_23385,N_23275);
nor UO_2665 (O_2665,N_24419,N_23655);
or UO_2666 (O_2666,N_23441,N_23056);
and UO_2667 (O_2667,N_24747,N_23277);
xor UO_2668 (O_2668,N_24083,N_23660);
or UO_2669 (O_2669,N_24848,N_24795);
or UO_2670 (O_2670,N_24636,N_23311);
nor UO_2671 (O_2671,N_22941,N_24445);
nor UO_2672 (O_2672,N_24760,N_23265);
and UO_2673 (O_2673,N_23878,N_24994);
xnor UO_2674 (O_2674,N_24976,N_24264);
or UO_2675 (O_2675,N_23078,N_22904);
or UO_2676 (O_2676,N_23583,N_23950);
and UO_2677 (O_2677,N_23114,N_24045);
xor UO_2678 (O_2678,N_24214,N_23842);
xnor UO_2679 (O_2679,N_24033,N_24954);
or UO_2680 (O_2680,N_23793,N_24586);
and UO_2681 (O_2681,N_23558,N_23704);
nand UO_2682 (O_2682,N_24727,N_23273);
nor UO_2683 (O_2683,N_24353,N_23808);
xnor UO_2684 (O_2684,N_22732,N_24896);
nand UO_2685 (O_2685,N_24828,N_24544);
nor UO_2686 (O_2686,N_23767,N_24282);
xor UO_2687 (O_2687,N_22974,N_24752);
nor UO_2688 (O_2688,N_24161,N_22980);
or UO_2689 (O_2689,N_22541,N_23298);
nor UO_2690 (O_2690,N_23756,N_22648);
xor UO_2691 (O_2691,N_23586,N_22940);
nand UO_2692 (O_2692,N_23151,N_22600);
and UO_2693 (O_2693,N_23359,N_23805);
and UO_2694 (O_2694,N_24961,N_22811);
nor UO_2695 (O_2695,N_23080,N_23045);
xor UO_2696 (O_2696,N_23396,N_24107);
or UO_2697 (O_2697,N_23529,N_22560);
and UO_2698 (O_2698,N_24162,N_24139);
and UO_2699 (O_2699,N_23247,N_24726);
nor UO_2700 (O_2700,N_23872,N_23107);
nand UO_2701 (O_2701,N_23208,N_24982);
and UO_2702 (O_2702,N_23058,N_24705);
or UO_2703 (O_2703,N_23378,N_23558);
nor UO_2704 (O_2704,N_24598,N_24269);
nand UO_2705 (O_2705,N_24155,N_24904);
or UO_2706 (O_2706,N_23606,N_24810);
xor UO_2707 (O_2707,N_24959,N_23467);
or UO_2708 (O_2708,N_23432,N_23949);
nor UO_2709 (O_2709,N_23588,N_22552);
nor UO_2710 (O_2710,N_24323,N_24964);
xor UO_2711 (O_2711,N_24109,N_24231);
and UO_2712 (O_2712,N_23386,N_22630);
or UO_2713 (O_2713,N_23176,N_23187);
or UO_2714 (O_2714,N_24520,N_24057);
or UO_2715 (O_2715,N_23864,N_22791);
nor UO_2716 (O_2716,N_22722,N_23686);
nand UO_2717 (O_2717,N_23173,N_24533);
nor UO_2718 (O_2718,N_24531,N_23308);
nand UO_2719 (O_2719,N_22845,N_22653);
or UO_2720 (O_2720,N_23855,N_24068);
nor UO_2721 (O_2721,N_24340,N_24498);
xnor UO_2722 (O_2722,N_23250,N_24170);
and UO_2723 (O_2723,N_23252,N_22605);
nor UO_2724 (O_2724,N_24138,N_24047);
or UO_2725 (O_2725,N_23813,N_22773);
nand UO_2726 (O_2726,N_22509,N_24801);
xor UO_2727 (O_2727,N_23298,N_22655);
nand UO_2728 (O_2728,N_24815,N_24171);
nor UO_2729 (O_2729,N_23823,N_24685);
and UO_2730 (O_2730,N_23202,N_24660);
xor UO_2731 (O_2731,N_22762,N_24634);
xor UO_2732 (O_2732,N_22635,N_24965);
and UO_2733 (O_2733,N_22561,N_24939);
nand UO_2734 (O_2734,N_22990,N_22984);
xor UO_2735 (O_2735,N_22748,N_22847);
nand UO_2736 (O_2736,N_23141,N_23867);
or UO_2737 (O_2737,N_23037,N_22918);
xnor UO_2738 (O_2738,N_23101,N_23062);
and UO_2739 (O_2739,N_24589,N_23567);
nor UO_2740 (O_2740,N_24397,N_24271);
xnor UO_2741 (O_2741,N_24785,N_22636);
or UO_2742 (O_2742,N_23915,N_22566);
nor UO_2743 (O_2743,N_23791,N_23441);
nor UO_2744 (O_2744,N_24727,N_24305);
nor UO_2745 (O_2745,N_22521,N_22859);
or UO_2746 (O_2746,N_23305,N_22879);
or UO_2747 (O_2747,N_24468,N_24441);
xor UO_2748 (O_2748,N_23086,N_23560);
xor UO_2749 (O_2749,N_22862,N_23731);
and UO_2750 (O_2750,N_23305,N_23822);
or UO_2751 (O_2751,N_24137,N_22789);
nand UO_2752 (O_2752,N_23391,N_22934);
nand UO_2753 (O_2753,N_23487,N_24978);
nand UO_2754 (O_2754,N_22613,N_23772);
and UO_2755 (O_2755,N_24370,N_23841);
or UO_2756 (O_2756,N_23074,N_23372);
nor UO_2757 (O_2757,N_23762,N_24803);
nand UO_2758 (O_2758,N_23425,N_23929);
or UO_2759 (O_2759,N_23469,N_24385);
or UO_2760 (O_2760,N_24213,N_23839);
nand UO_2761 (O_2761,N_24846,N_24946);
nor UO_2762 (O_2762,N_24977,N_24943);
and UO_2763 (O_2763,N_24403,N_23089);
or UO_2764 (O_2764,N_23630,N_24045);
or UO_2765 (O_2765,N_23625,N_23234);
or UO_2766 (O_2766,N_23111,N_24726);
nor UO_2767 (O_2767,N_23637,N_23786);
nor UO_2768 (O_2768,N_22877,N_24351);
xor UO_2769 (O_2769,N_24953,N_23848);
or UO_2770 (O_2770,N_23221,N_22878);
nor UO_2771 (O_2771,N_24206,N_23951);
xor UO_2772 (O_2772,N_23734,N_23770);
nand UO_2773 (O_2773,N_23870,N_23217);
and UO_2774 (O_2774,N_23166,N_23279);
nand UO_2775 (O_2775,N_23300,N_23512);
nand UO_2776 (O_2776,N_23502,N_22993);
and UO_2777 (O_2777,N_24154,N_24210);
xnor UO_2778 (O_2778,N_24240,N_23567);
or UO_2779 (O_2779,N_23304,N_23739);
xnor UO_2780 (O_2780,N_23179,N_23285);
and UO_2781 (O_2781,N_24308,N_24987);
nor UO_2782 (O_2782,N_22511,N_23902);
nor UO_2783 (O_2783,N_22810,N_24869);
or UO_2784 (O_2784,N_24220,N_23921);
xor UO_2785 (O_2785,N_24925,N_23386);
xor UO_2786 (O_2786,N_23477,N_23867);
or UO_2787 (O_2787,N_23466,N_24276);
nor UO_2788 (O_2788,N_23671,N_24826);
and UO_2789 (O_2789,N_24761,N_23656);
and UO_2790 (O_2790,N_24771,N_24988);
and UO_2791 (O_2791,N_23676,N_24227);
nor UO_2792 (O_2792,N_24880,N_24169);
nor UO_2793 (O_2793,N_23472,N_23823);
or UO_2794 (O_2794,N_23701,N_24768);
nand UO_2795 (O_2795,N_23316,N_22919);
and UO_2796 (O_2796,N_23224,N_24849);
or UO_2797 (O_2797,N_22730,N_22774);
or UO_2798 (O_2798,N_23933,N_24200);
nand UO_2799 (O_2799,N_24188,N_23373);
and UO_2800 (O_2800,N_23521,N_24858);
nor UO_2801 (O_2801,N_23439,N_23009);
xor UO_2802 (O_2802,N_23446,N_24793);
nor UO_2803 (O_2803,N_23751,N_22992);
nor UO_2804 (O_2804,N_23108,N_23291);
nor UO_2805 (O_2805,N_24809,N_23616);
nor UO_2806 (O_2806,N_23612,N_24030);
nand UO_2807 (O_2807,N_24808,N_23516);
nor UO_2808 (O_2808,N_24323,N_24748);
nand UO_2809 (O_2809,N_23401,N_24973);
and UO_2810 (O_2810,N_23086,N_22741);
nand UO_2811 (O_2811,N_24391,N_23163);
or UO_2812 (O_2812,N_23950,N_23511);
or UO_2813 (O_2813,N_24345,N_24007);
xor UO_2814 (O_2814,N_24825,N_23449);
or UO_2815 (O_2815,N_22516,N_22799);
nand UO_2816 (O_2816,N_24141,N_24127);
xnor UO_2817 (O_2817,N_24666,N_22708);
nor UO_2818 (O_2818,N_24039,N_23937);
and UO_2819 (O_2819,N_24489,N_24301);
or UO_2820 (O_2820,N_24388,N_24371);
nand UO_2821 (O_2821,N_24365,N_23395);
and UO_2822 (O_2822,N_23882,N_23150);
nand UO_2823 (O_2823,N_24863,N_23150);
nor UO_2824 (O_2824,N_24889,N_24176);
xnor UO_2825 (O_2825,N_23171,N_23606);
or UO_2826 (O_2826,N_22746,N_24428);
and UO_2827 (O_2827,N_23434,N_23064);
nand UO_2828 (O_2828,N_24353,N_23831);
nand UO_2829 (O_2829,N_23535,N_22690);
or UO_2830 (O_2830,N_22572,N_22509);
or UO_2831 (O_2831,N_22573,N_23133);
and UO_2832 (O_2832,N_24603,N_24028);
nand UO_2833 (O_2833,N_22954,N_23391);
nand UO_2834 (O_2834,N_24052,N_22557);
nand UO_2835 (O_2835,N_22653,N_24494);
and UO_2836 (O_2836,N_22516,N_24141);
or UO_2837 (O_2837,N_22808,N_24100);
nand UO_2838 (O_2838,N_23843,N_23414);
nand UO_2839 (O_2839,N_24724,N_23811);
xor UO_2840 (O_2840,N_22841,N_24973);
and UO_2841 (O_2841,N_23461,N_23152);
nor UO_2842 (O_2842,N_22790,N_23981);
nand UO_2843 (O_2843,N_24198,N_23229);
nand UO_2844 (O_2844,N_24126,N_24677);
xor UO_2845 (O_2845,N_24020,N_24538);
nor UO_2846 (O_2846,N_23646,N_23346);
xnor UO_2847 (O_2847,N_23997,N_24649);
nor UO_2848 (O_2848,N_24335,N_22827);
nor UO_2849 (O_2849,N_23048,N_23784);
nor UO_2850 (O_2850,N_24901,N_23840);
xnor UO_2851 (O_2851,N_22724,N_23339);
and UO_2852 (O_2852,N_22699,N_22588);
nand UO_2853 (O_2853,N_24251,N_23805);
nand UO_2854 (O_2854,N_24825,N_23169);
and UO_2855 (O_2855,N_23305,N_24932);
nor UO_2856 (O_2856,N_23225,N_22805);
and UO_2857 (O_2857,N_22771,N_22911);
xor UO_2858 (O_2858,N_24741,N_22817);
nand UO_2859 (O_2859,N_24040,N_24108);
and UO_2860 (O_2860,N_22932,N_24005);
and UO_2861 (O_2861,N_23464,N_23379);
xor UO_2862 (O_2862,N_24410,N_24316);
and UO_2863 (O_2863,N_22600,N_22504);
or UO_2864 (O_2864,N_24141,N_23987);
or UO_2865 (O_2865,N_23596,N_22888);
nand UO_2866 (O_2866,N_24733,N_22792);
nor UO_2867 (O_2867,N_23294,N_23324);
or UO_2868 (O_2868,N_23913,N_24459);
or UO_2869 (O_2869,N_23702,N_24358);
and UO_2870 (O_2870,N_24415,N_23184);
nand UO_2871 (O_2871,N_23787,N_24687);
and UO_2872 (O_2872,N_23991,N_24533);
nand UO_2873 (O_2873,N_24402,N_23305);
or UO_2874 (O_2874,N_24193,N_24805);
xnor UO_2875 (O_2875,N_22579,N_24106);
nor UO_2876 (O_2876,N_22625,N_23653);
nand UO_2877 (O_2877,N_23507,N_23518);
xor UO_2878 (O_2878,N_23388,N_23024);
nor UO_2879 (O_2879,N_22949,N_22660);
or UO_2880 (O_2880,N_24941,N_23529);
nor UO_2881 (O_2881,N_24997,N_22794);
nand UO_2882 (O_2882,N_24299,N_23347);
nor UO_2883 (O_2883,N_24984,N_24369);
xnor UO_2884 (O_2884,N_22506,N_23825);
or UO_2885 (O_2885,N_23270,N_22715);
and UO_2886 (O_2886,N_23457,N_22515);
and UO_2887 (O_2887,N_24652,N_23016);
nor UO_2888 (O_2888,N_24786,N_23972);
xnor UO_2889 (O_2889,N_22730,N_23406);
or UO_2890 (O_2890,N_24479,N_23303);
nor UO_2891 (O_2891,N_22962,N_22841);
xor UO_2892 (O_2892,N_24972,N_22806);
nor UO_2893 (O_2893,N_23287,N_24247);
nand UO_2894 (O_2894,N_23946,N_23048);
nor UO_2895 (O_2895,N_24342,N_24615);
and UO_2896 (O_2896,N_23144,N_24962);
or UO_2897 (O_2897,N_24386,N_24097);
nor UO_2898 (O_2898,N_24593,N_22538);
nor UO_2899 (O_2899,N_23342,N_23282);
nand UO_2900 (O_2900,N_23691,N_22960);
or UO_2901 (O_2901,N_23462,N_23684);
xor UO_2902 (O_2902,N_24807,N_22612);
or UO_2903 (O_2903,N_23800,N_23236);
or UO_2904 (O_2904,N_24800,N_23358);
nor UO_2905 (O_2905,N_24583,N_22851);
xor UO_2906 (O_2906,N_24441,N_23151);
nor UO_2907 (O_2907,N_23142,N_24681);
nor UO_2908 (O_2908,N_23575,N_24539);
or UO_2909 (O_2909,N_23661,N_23869);
nand UO_2910 (O_2910,N_23835,N_24784);
nor UO_2911 (O_2911,N_22982,N_23829);
nand UO_2912 (O_2912,N_23811,N_24126);
nand UO_2913 (O_2913,N_22505,N_24726);
nor UO_2914 (O_2914,N_24456,N_23857);
and UO_2915 (O_2915,N_22550,N_24244);
and UO_2916 (O_2916,N_23165,N_23515);
or UO_2917 (O_2917,N_23877,N_23911);
or UO_2918 (O_2918,N_24701,N_22819);
nor UO_2919 (O_2919,N_23286,N_24393);
or UO_2920 (O_2920,N_24277,N_23759);
or UO_2921 (O_2921,N_24731,N_23034);
and UO_2922 (O_2922,N_23254,N_23806);
nand UO_2923 (O_2923,N_22655,N_24961);
xnor UO_2924 (O_2924,N_24065,N_23836);
nand UO_2925 (O_2925,N_23404,N_22786);
nand UO_2926 (O_2926,N_22787,N_23176);
nor UO_2927 (O_2927,N_24499,N_24582);
and UO_2928 (O_2928,N_22904,N_24539);
xor UO_2929 (O_2929,N_23746,N_22524);
and UO_2930 (O_2930,N_23884,N_24091);
and UO_2931 (O_2931,N_24048,N_23507);
xnor UO_2932 (O_2932,N_22771,N_24207);
nand UO_2933 (O_2933,N_22861,N_24219);
xor UO_2934 (O_2934,N_24915,N_23373);
or UO_2935 (O_2935,N_22735,N_24928);
nand UO_2936 (O_2936,N_23330,N_22611);
nor UO_2937 (O_2937,N_23186,N_23552);
nor UO_2938 (O_2938,N_23821,N_22984);
and UO_2939 (O_2939,N_22543,N_24506);
nand UO_2940 (O_2940,N_23094,N_22902);
nand UO_2941 (O_2941,N_22824,N_23221);
or UO_2942 (O_2942,N_24848,N_23044);
and UO_2943 (O_2943,N_23852,N_24627);
and UO_2944 (O_2944,N_24200,N_22829);
xnor UO_2945 (O_2945,N_23185,N_23904);
nor UO_2946 (O_2946,N_22519,N_24374);
xor UO_2947 (O_2947,N_24350,N_23596);
xor UO_2948 (O_2948,N_24849,N_23618);
and UO_2949 (O_2949,N_23679,N_22868);
nand UO_2950 (O_2950,N_23705,N_24457);
nand UO_2951 (O_2951,N_22686,N_24034);
nor UO_2952 (O_2952,N_23475,N_24125);
nand UO_2953 (O_2953,N_23041,N_23834);
nor UO_2954 (O_2954,N_24266,N_22993);
and UO_2955 (O_2955,N_23051,N_24624);
xor UO_2956 (O_2956,N_24099,N_23195);
and UO_2957 (O_2957,N_24594,N_23002);
xnor UO_2958 (O_2958,N_24474,N_23186);
xnor UO_2959 (O_2959,N_22501,N_23865);
or UO_2960 (O_2960,N_24053,N_23537);
nor UO_2961 (O_2961,N_24893,N_24066);
xor UO_2962 (O_2962,N_23202,N_24379);
or UO_2963 (O_2963,N_24424,N_24688);
nand UO_2964 (O_2964,N_24797,N_22688);
nand UO_2965 (O_2965,N_23051,N_24710);
nor UO_2966 (O_2966,N_22723,N_23149);
and UO_2967 (O_2967,N_24015,N_24322);
nor UO_2968 (O_2968,N_23056,N_23284);
or UO_2969 (O_2969,N_22627,N_22857);
xnor UO_2970 (O_2970,N_22669,N_22550);
xor UO_2971 (O_2971,N_24035,N_24707);
and UO_2972 (O_2972,N_24653,N_23882);
nand UO_2973 (O_2973,N_24388,N_22681);
nor UO_2974 (O_2974,N_24828,N_24629);
and UO_2975 (O_2975,N_23825,N_24407);
nor UO_2976 (O_2976,N_23673,N_23699);
xor UO_2977 (O_2977,N_24259,N_24913);
and UO_2978 (O_2978,N_24834,N_24244);
xor UO_2979 (O_2979,N_24727,N_23397);
nand UO_2980 (O_2980,N_24460,N_24847);
nand UO_2981 (O_2981,N_23312,N_24679);
nor UO_2982 (O_2982,N_24079,N_24054);
or UO_2983 (O_2983,N_24534,N_23959);
or UO_2984 (O_2984,N_23731,N_24569);
nand UO_2985 (O_2985,N_23569,N_23455);
and UO_2986 (O_2986,N_24941,N_23436);
nand UO_2987 (O_2987,N_24111,N_24544);
nor UO_2988 (O_2988,N_24351,N_24157);
xor UO_2989 (O_2989,N_24762,N_22695);
nor UO_2990 (O_2990,N_22759,N_24111);
nor UO_2991 (O_2991,N_24379,N_22638);
xnor UO_2992 (O_2992,N_24422,N_24864);
and UO_2993 (O_2993,N_24052,N_24242);
and UO_2994 (O_2994,N_23223,N_24750);
nand UO_2995 (O_2995,N_24578,N_24334);
nand UO_2996 (O_2996,N_24147,N_24089);
or UO_2997 (O_2997,N_23292,N_22637);
and UO_2998 (O_2998,N_22539,N_22807);
nor UO_2999 (O_2999,N_22862,N_23324);
endmodule