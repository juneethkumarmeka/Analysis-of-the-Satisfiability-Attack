module basic_1500_15000_2000_100_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
xnor U0 (N_0,In_376,In_957);
or U1 (N_1,In_135,In_219);
nor U2 (N_2,In_1363,In_400);
nand U3 (N_3,In_491,In_122);
nor U4 (N_4,In_928,In_521);
nor U5 (N_5,In_790,In_719);
nand U6 (N_6,In_1186,In_296);
and U7 (N_7,In_967,In_819);
nand U8 (N_8,In_1098,In_1355);
or U9 (N_9,In_1494,In_862);
or U10 (N_10,In_745,In_752);
or U11 (N_11,In_1128,In_1307);
xor U12 (N_12,In_1065,In_482);
nor U13 (N_13,In_299,In_1177);
xor U14 (N_14,In_120,In_365);
xor U15 (N_15,In_1377,In_825);
or U16 (N_16,In_938,In_635);
or U17 (N_17,In_1053,In_751);
nor U18 (N_18,In_1288,In_1178);
nand U19 (N_19,In_177,In_1235);
nor U20 (N_20,In_735,In_650);
and U21 (N_21,In_214,In_382);
and U22 (N_22,In_168,In_1077);
xor U23 (N_23,In_600,In_1035);
nor U24 (N_24,In_785,In_802);
or U25 (N_25,In_555,In_822);
or U26 (N_26,In_658,In_1193);
or U27 (N_27,In_551,In_272);
nand U28 (N_28,In_1020,In_99);
xnor U29 (N_29,In_750,In_370);
and U30 (N_30,In_60,In_150);
xnor U31 (N_31,In_1245,In_1084);
nand U32 (N_32,In_298,In_534);
nor U33 (N_33,In_260,In_746);
xnor U34 (N_34,In_1069,In_1075);
xor U35 (N_35,In_1331,In_1366);
xnor U36 (N_36,In_730,In_309);
nor U37 (N_37,In_328,In_1419);
nor U38 (N_38,In_619,In_721);
or U39 (N_39,In_1091,In_1292);
xor U40 (N_40,In_960,In_1085);
nor U41 (N_41,In_1064,In_1231);
nand U42 (N_42,In_109,In_1176);
xnor U43 (N_43,In_458,In_627);
nor U44 (N_44,In_212,In_171);
xnor U45 (N_45,In_300,In_1353);
nor U46 (N_46,In_1442,In_451);
nand U47 (N_47,In_1259,In_203);
xnor U48 (N_48,In_1341,In_925);
xnor U49 (N_49,In_844,In_1452);
nor U50 (N_50,In_1291,In_565);
nor U51 (N_51,In_991,In_607);
or U52 (N_52,In_1301,In_1309);
xnor U53 (N_53,In_722,In_715);
nor U54 (N_54,In_502,In_392);
xor U55 (N_55,In_30,In_1112);
nand U56 (N_56,In_1016,In_1086);
and U57 (N_57,In_73,In_1451);
nor U58 (N_58,In_791,In_1456);
nor U59 (N_59,In_577,In_383);
or U60 (N_60,In_548,In_562);
xnor U61 (N_61,In_630,In_853);
nand U62 (N_62,In_833,In_852);
or U63 (N_63,In_1125,In_1191);
and U64 (N_64,In_1026,In_229);
or U65 (N_65,In_836,In_44);
nand U66 (N_66,In_995,In_1232);
nor U67 (N_67,In_312,In_1019);
xor U68 (N_68,In_660,In_1047);
and U69 (N_69,In_553,In_238);
xor U70 (N_70,In_1478,In_977);
and U71 (N_71,In_835,In_818);
nor U72 (N_72,In_531,In_1246);
and U73 (N_73,In_1411,In_446);
nor U74 (N_74,In_330,In_37);
and U75 (N_75,In_505,In_2);
xnor U76 (N_76,In_448,In_367);
nand U77 (N_77,In_388,In_485);
nand U78 (N_78,In_1345,In_1261);
nor U79 (N_79,In_682,In_36);
nor U80 (N_80,In_209,In_1145);
nand U81 (N_81,In_659,In_1276);
or U82 (N_82,In_1289,In_1332);
or U83 (N_83,In_1201,In_107);
or U84 (N_84,In_1150,In_806);
and U85 (N_85,In_795,In_249);
and U86 (N_86,In_695,In_5);
xor U87 (N_87,In_63,In_1044);
xnor U88 (N_88,In_1117,In_517);
xnor U89 (N_89,In_205,In_59);
xnor U90 (N_90,In_245,In_1168);
and U91 (N_91,In_713,In_1290);
and U92 (N_92,In_871,In_436);
or U93 (N_93,In_754,In_1444);
or U94 (N_94,In_151,In_158);
and U95 (N_95,In_687,In_1080);
or U96 (N_96,In_596,In_242);
and U97 (N_97,In_613,In_899);
or U98 (N_98,In_574,In_1446);
and U99 (N_99,In_1467,In_804);
nor U100 (N_100,In_435,In_199);
xor U101 (N_101,In_114,In_493);
nand U102 (N_102,In_167,In_759);
and U103 (N_103,In_442,In_616);
nor U104 (N_104,In_605,In_1265);
nor U105 (N_105,In_610,In_936);
nand U106 (N_106,In_592,In_1129);
and U107 (N_107,In_1347,In_344);
nand U108 (N_108,In_1425,In_947);
and U109 (N_109,In_340,In_1094);
nor U110 (N_110,In_47,In_923);
nor U111 (N_111,In_137,In_384);
xnor U112 (N_112,In_52,In_744);
xor U113 (N_113,In_1491,In_90);
and U114 (N_114,In_969,In_1378);
nor U115 (N_115,In_1106,In_82);
nor U116 (N_116,In_1154,In_1316);
and U117 (N_117,In_667,In_1063);
and U118 (N_118,In_766,In_1163);
nand U119 (N_119,In_612,In_1293);
and U120 (N_120,In_526,In_879);
and U121 (N_121,In_1413,In_1438);
or U122 (N_122,In_1382,In_462);
nand U123 (N_123,In_1306,In_1090);
and U124 (N_124,In_1387,In_780);
or U125 (N_125,In_823,In_1267);
nand U126 (N_126,In_520,In_1471);
or U127 (N_127,In_768,In_758);
nor U128 (N_128,In_302,In_1092);
or U129 (N_129,In_1134,In_208);
nand U130 (N_130,In_1473,In_1322);
nand U131 (N_131,In_256,In_511);
nor U132 (N_132,In_1173,In_631);
nor U133 (N_133,In_821,In_1405);
nand U134 (N_134,In_901,In_147);
nand U135 (N_135,In_11,In_83);
xor U136 (N_136,In_50,In_268);
or U137 (N_137,In_1399,In_69);
nor U138 (N_138,In_655,In_569);
nor U139 (N_139,In_697,In_471);
and U140 (N_140,In_1251,In_727);
and U141 (N_141,In_1083,In_181);
or U142 (N_142,In_132,In_352);
nor U143 (N_143,In_1192,In_41);
nand U144 (N_144,In_430,In_914);
or U145 (N_145,In_789,In_628);
xor U146 (N_146,In_717,In_1459);
or U147 (N_147,In_1321,In_98);
xnor U148 (N_148,In_454,In_504);
xor U149 (N_149,In_918,In_1006);
and U150 (N_150,In_684,In_677);
nand U151 (N_151,In_1249,In_239);
xnor U152 (N_152,In_926,In_519);
xnor U153 (N_153,In_664,In_1118);
and U154 (N_154,In_621,In_1130);
nor U155 (N_155,In_1463,In_770);
or U156 (N_156,In_1317,N_13);
xor U157 (N_157,In_525,In_438);
and U158 (N_158,In_142,In_557);
and U159 (N_159,In_467,In_1000);
nand U160 (N_160,N_76,In_1385);
nand U161 (N_161,In_351,N_100);
nor U162 (N_162,In_1258,In_463);
and U163 (N_163,In_705,N_37);
nand U164 (N_164,N_73,In_1350);
and U165 (N_165,N_47,N_21);
or U166 (N_166,In_7,N_72);
or U167 (N_167,In_381,In_247);
and U168 (N_168,In_1038,In_892);
nand U169 (N_169,In_1270,In_1423);
and U170 (N_170,In_950,In_774);
xnor U171 (N_171,In_803,In_93);
xnor U172 (N_172,In_1171,In_1361);
and U173 (N_173,In_134,In_1359);
xnor U174 (N_174,In_127,In_1212);
or U175 (N_175,In_198,In_495);
nor U176 (N_176,In_461,In_1052);
and U177 (N_177,In_210,In_545);
and U178 (N_178,In_255,In_43);
xor U179 (N_179,In_14,In_1062);
nor U180 (N_180,In_753,N_141);
or U181 (N_181,In_1081,In_372);
xnor U182 (N_182,In_742,In_787);
and U183 (N_183,In_1257,In_117);
nand U184 (N_184,In_455,N_25);
nand U185 (N_185,In_536,N_65);
nand U186 (N_186,N_136,In_1137);
and U187 (N_187,N_92,In_395);
nor U188 (N_188,In_952,In_817);
xnor U189 (N_189,In_1389,In_1078);
nor U190 (N_190,In_941,In_139);
nand U191 (N_191,In_942,In_406);
or U192 (N_192,In_543,In_8);
nor U193 (N_193,In_1298,In_761);
nor U194 (N_194,N_42,In_972);
nand U195 (N_195,In_1184,In_642);
nand U196 (N_196,In_1138,In_1430);
xnor U197 (N_197,N_148,In_1082);
nor U198 (N_198,In_149,In_207);
or U199 (N_199,In_637,In_830);
nor U200 (N_200,In_1021,In_1202);
nor U201 (N_201,In_1144,In_813);
xor U202 (N_202,In_691,In_893);
or U203 (N_203,In_1023,In_475);
xor U204 (N_204,In_1189,In_638);
nand U205 (N_205,In_1343,In_1054);
nand U206 (N_206,In_1320,In_19);
and U207 (N_207,In_9,N_52);
and U208 (N_208,In_934,In_1131);
nand U209 (N_209,In_561,In_85);
xnor U210 (N_210,In_832,In_1179);
nor U211 (N_211,In_1216,In_601);
or U212 (N_212,In_1376,In_775);
xor U213 (N_213,In_1205,In_10);
or U214 (N_214,In_550,In_478);
nand U215 (N_215,In_634,In_1498);
or U216 (N_216,In_854,In_1402);
or U217 (N_217,In_827,In_1421);
or U218 (N_218,In_261,N_10);
nor U219 (N_219,In_760,In_796);
xor U220 (N_220,In_1194,In_13);
or U221 (N_221,In_808,In_213);
and U222 (N_222,In_464,N_16);
or U223 (N_223,In_1400,In_427);
xor U224 (N_224,In_1370,N_19);
or U225 (N_225,In_466,In_162);
and U226 (N_226,In_444,In_424);
xnor U227 (N_227,In_843,N_85);
nor U228 (N_228,N_102,In_554);
xor U229 (N_229,In_902,In_1260);
or U230 (N_230,In_360,In_1417);
and U231 (N_231,In_81,In_1066);
nand U232 (N_232,In_129,In_962);
or U233 (N_233,In_1381,In_1076);
nand U234 (N_234,In_76,In_1479);
nand U235 (N_235,In_1356,In_1156);
nor U236 (N_236,In_645,In_1334);
nor U237 (N_237,In_1283,In_200);
xnor U238 (N_238,N_139,In_593);
xor U239 (N_239,In_812,In_397);
and U240 (N_240,In_178,In_323);
nand U241 (N_241,In_1256,In_319);
or U242 (N_242,In_416,In_1455);
and U243 (N_243,In_1217,N_40);
nand U244 (N_244,N_87,In_1308);
xnor U245 (N_245,In_332,In_980);
nand U246 (N_246,In_18,In_1036);
or U247 (N_247,In_377,In_116);
xor U248 (N_248,In_1474,In_762);
or U249 (N_249,In_1379,In_1364);
nand U250 (N_250,N_1,In_288);
xnor U251 (N_251,In_155,In_673);
nor U252 (N_252,In_737,In_1155);
nor U253 (N_253,In_1342,In_1485);
or U254 (N_254,In_1277,In_341);
nor U255 (N_255,In_253,In_1482);
and U256 (N_256,In_1059,In_643);
and U257 (N_257,In_529,N_2);
xor U258 (N_258,In_46,In_724);
nor U259 (N_259,In_1010,In_170);
or U260 (N_260,In_1073,In_1214);
and U261 (N_261,In_878,In_257);
nor U262 (N_262,In_233,In_723);
nor U263 (N_263,In_1149,In_978);
xnor U264 (N_264,In_1029,In_767);
nand U265 (N_265,In_685,In_161);
nor U266 (N_266,In_575,In_647);
xor U267 (N_267,In_1369,In_845);
or U268 (N_268,N_104,In_935);
or U269 (N_269,In_1057,N_66);
xnor U270 (N_270,In_387,In_1027);
nand U271 (N_271,In_437,In_496);
or U272 (N_272,In_183,In_1237);
nand U273 (N_273,In_349,In_994);
nor U274 (N_274,In_407,In_1056);
nor U275 (N_275,In_1286,N_9);
or U276 (N_276,In_1305,In_680);
and U277 (N_277,In_235,In_856);
nand U278 (N_278,In_710,In_598);
nor U279 (N_279,N_23,In_426);
xor U280 (N_280,In_749,In_1042);
nand U281 (N_281,In_1050,In_1101);
xor U282 (N_282,In_809,N_114);
nand U283 (N_283,In_1311,In_670);
nand U284 (N_284,In_265,In_1172);
nor U285 (N_285,In_1412,In_1367);
and U286 (N_286,In_1008,In_528);
xnor U287 (N_287,In_133,In_350);
xnor U288 (N_288,In_867,In_39);
xor U289 (N_289,In_468,In_291);
xnor U290 (N_290,In_986,In_16);
xor U291 (N_291,In_681,In_1335);
nor U292 (N_292,In_62,In_56);
nor U293 (N_293,N_75,N_48);
nand U294 (N_294,N_122,In_949);
and U295 (N_295,In_215,In_346);
nor U296 (N_296,N_27,In_194);
nand U297 (N_297,In_527,In_1159);
xor U298 (N_298,In_379,In_23);
xor U299 (N_299,In_1152,In_731);
or U300 (N_300,In_483,N_280);
and U301 (N_301,In_898,In_917);
and U302 (N_302,In_188,N_112);
nand U303 (N_303,In_646,In_927);
xnor U304 (N_304,In_439,In_1440);
nor U305 (N_305,In_985,N_71);
nor U306 (N_306,In_1093,In_1097);
nor U307 (N_307,In_396,In_1060);
and U308 (N_308,In_320,In_699);
or U309 (N_309,In_304,In_22);
or U310 (N_310,In_378,N_276);
nor U311 (N_311,In_1354,In_1041);
xor U312 (N_312,N_227,In_999);
nor U313 (N_313,In_1282,In_763);
nor U314 (N_314,In_273,In_870);
nand U315 (N_315,In_123,In_595);
xor U316 (N_316,In_267,In_1233);
and U317 (N_317,In_961,N_181);
or U318 (N_318,In_153,In_837);
nor U319 (N_319,In_1380,In_362);
or U320 (N_320,In_1229,In_987);
and U321 (N_321,In_71,In_417);
nand U322 (N_322,N_242,In_1104);
nor U323 (N_323,In_712,In_1344);
nor U324 (N_324,In_625,In_1487);
nor U325 (N_325,N_249,In_269);
nor U326 (N_326,In_259,In_289);
nor U327 (N_327,In_706,In_1161);
xnor U328 (N_328,In_49,N_158);
nor U329 (N_329,In_811,In_1348);
nor U330 (N_330,In_580,In_115);
or U331 (N_331,In_686,In_908);
xor U332 (N_332,In_1011,In_709);
nand U333 (N_333,In_1174,In_944);
or U334 (N_334,In_951,In_87);
or U335 (N_335,In_1074,In_903);
or U336 (N_336,In_1218,N_33);
nand U337 (N_337,In_512,In_939);
and U338 (N_338,In_1222,In_1484);
or U339 (N_339,In_310,In_1210);
and U340 (N_340,N_213,N_30);
or U341 (N_341,N_254,In_230);
nand U342 (N_342,In_1181,In_541);
xnor U343 (N_343,In_1158,In_973);
nor U344 (N_344,In_1271,N_152);
nor U345 (N_345,In_1169,In_875);
or U346 (N_346,In_588,In_1426);
nand U347 (N_347,In_798,In_640);
and U348 (N_348,In_1424,In_481);
or U349 (N_349,In_1116,In_539);
nor U350 (N_350,In_386,In_606);
xnor U351 (N_351,In_1133,In_347);
or U352 (N_352,In_1190,In_412);
xor U353 (N_353,N_177,In_698);
nor U354 (N_354,In_755,In_61);
xnor U355 (N_355,In_477,In_1365);
xnor U356 (N_356,In_1015,In_1230);
nor U357 (N_357,In_916,In_104);
nor U358 (N_358,In_1318,In_954);
nand U359 (N_359,In_278,In_842);
and U360 (N_360,In_1462,In_275);
xnor U361 (N_361,N_176,N_145);
xnor U362 (N_362,N_147,In_1394);
nand U363 (N_363,In_583,N_39);
nand U364 (N_364,N_3,In_78);
or U365 (N_365,In_1032,In_847);
nand U366 (N_366,N_140,In_964);
or U367 (N_367,In_1295,In_348);
nor U368 (N_368,In_1457,In_1466);
xor U369 (N_369,In_1211,In_157);
and U370 (N_370,In_846,In_1071);
and U371 (N_371,In_500,In_223);
xor U372 (N_372,In_848,In_538);
xor U373 (N_373,In_1495,In_1022);
and U374 (N_374,In_469,In_1046);
and U375 (N_375,In_301,N_68);
xnor U376 (N_376,In_1488,In_315);
xor U377 (N_377,In_708,In_51);
or U378 (N_378,In_110,In_476);
xor U379 (N_379,In_373,In_1285);
and U380 (N_380,In_937,In_581);
nor U381 (N_381,N_273,N_224);
xor U382 (N_382,In_1051,In_799);
xor U383 (N_383,N_264,In_415);
or U384 (N_384,In_425,In_326);
xor U385 (N_385,In_264,In_544);
or U386 (N_386,N_172,N_154);
and U387 (N_387,In_945,N_204);
nand U388 (N_388,In_1004,In_884);
or U389 (N_389,In_79,In_841);
nor U390 (N_390,N_219,N_26);
nor U391 (N_391,In_1362,In_1325);
nand U392 (N_392,In_154,In_958);
nand U393 (N_393,In_933,In_277);
and U394 (N_394,N_150,In_112);
xnor U395 (N_395,In_943,N_103);
or U396 (N_396,N_196,In_982);
nand U397 (N_397,In_876,N_216);
and U398 (N_398,N_261,N_164);
xnor U399 (N_399,In_1453,In_21);
or U400 (N_400,In_1127,In_840);
nand U401 (N_401,In_96,In_1242);
and U402 (N_402,N_189,In_932);
nand U403 (N_403,In_979,In_187);
nor U404 (N_404,In_1266,In_1352);
or U405 (N_405,In_897,In_1135);
or U406 (N_406,In_1096,In_159);
and U407 (N_407,In_689,N_81);
or U408 (N_408,In_904,N_101);
or U409 (N_409,N_185,N_61);
and U410 (N_410,N_171,N_250);
and U411 (N_411,In_1340,In_1328);
nand U412 (N_412,In_447,In_887);
nand U413 (N_413,In_290,In_358);
nand U414 (N_414,In_414,In_1486);
xnor U415 (N_415,In_891,In_981);
nor U416 (N_416,In_393,In_308);
nor U417 (N_417,In_1262,In_108);
nor U418 (N_418,In_629,In_1204);
xnor U419 (N_419,In_164,N_86);
xnor U420 (N_420,In_1119,In_357);
or U421 (N_421,In_820,N_146);
xnor U422 (N_422,In_1220,In_1025);
nand U423 (N_423,In_1396,In_111);
or U424 (N_424,In_1414,N_24);
nand U425 (N_425,In_998,N_186);
or U426 (N_426,In_40,In_390);
nand U427 (N_427,In_889,In_1165);
xor U428 (N_428,N_131,N_14);
or U429 (N_429,In_95,N_118);
xnor U430 (N_430,N_230,In_1164);
nor U431 (N_431,In_72,In_498);
nor U432 (N_432,In_678,In_402);
nand U433 (N_433,N_64,In_281);
xor U434 (N_434,In_1199,In_1209);
nor U435 (N_435,N_255,In_1294);
xnor U436 (N_436,In_1147,In_1383);
nor U437 (N_437,In_1250,In_152);
and U438 (N_438,In_55,In_620);
nor U439 (N_439,In_53,In_459);
and U440 (N_440,In_510,In_1252);
nor U441 (N_441,N_58,N_127);
nor U442 (N_442,In_196,In_912);
nor U443 (N_443,In_1033,In_355);
nor U444 (N_444,In_1140,In_1226);
xnor U445 (N_445,In_35,In_524);
nor U446 (N_446,In_585,In_570);
nand U447 (N_447,In_1089,N_289);
nand U448 (N_448,In_1493,N_259);
and U449 (N_449,In_615,In_1225);
and U450 (N_450,N_297,In_1392);
xnor U451 (N_451,In_696,In_515);
or U452 (N_452,N_310,In_1088);
nand U453 (N_453,In_1003,In_850);
nand U454 (N_454,N_41,In_490);
xnor U455 (N_455,In_262,In_280);
or U456 (N_456,In_389,In_156);
and U457 (N_457,N_334,In_486);
nor U458 (N_458,N_142,N_99);
xor U459 (N_459,N_281,In_869);
or U460 (N_460,In_1441,In_503);
nor U461 (N_461,N_208,In_1481);
nand U462 (N_462,N_195,N_178);
nor U463 (N_463,N_315,In_246);
and U464 (N_464,In_67,N_190);
nor U465 (N_465,In_86,In_31);
xnor U466 (N_466,In_586,In_404);
nor U467 (N_467,In_990,In_956);
nor U468 (N_468,N_44,In_1284);
or U469 (N_469,N_174,In_700);
or U470 (N_470,In_1475,In_29);
or U471 (N_471,In_48,In_984);
and U472 (N_472,N_212,In_1420);
and U473 (N_473,In_399,N_420);
nor U474 (N_474,In_174,In_801);
or U475 (N_475,In_353,In_191);
and U476 (N_476,In_189,N_275);
nor U477 (N_477,N_153,In_1200);
or U478 (N_478,In_1448,In_1429);
and U479 (N_479,In_547,In_287);
and U480 (N_480,In_1110,In_465);
and U481 (N_481,In_366,N_49);
and U482 (N_482,In_1304,N_238);
nor U483 (N_483,In_1312,In_1049);
nand U484 (N_484,In_1195,N_434);
nand U485 (N_485,N_271,In_38);
and U486 (N_486,N_312,In_248);
nand U487 (N_487,In_1433,In_329);
nor U488 (N_488,In_757,In_317);
nand U489 (N_489,In_1449,N_165);
or U490 (N_490,In_974,In_136);
nand U491 (N_491,In_421,N_79);
nor U492 (N_492,N_416,In_922);
nor U493 (N_493,In_1275,N_53);
nand U494 (N_494,N_63,N_5);
xor U495 (N_495,In_513,In_861);
nand U496 (N_496,N_294,In_125);
or U497 (N_497,In_651,In_608);
and U498 (N_498,N_395,In_1464);
xor U499 (N_499,N_188,In_829);
xnor U500 (N_500,N_210,In_27);
or U501 (N_501,N_372,In_614);
nor U502 (N_502,In_431,In_364);
or U503 (N_503,In_231,N_262);
xnor U504 (N_504,N_78,N_388);
nand U505 (N_505,N_365,In_649);
nor U506 (N_506,N_411,In_924);
or U507 (N_507,In_285,In_1302);
nand U508 (N_508,In_1197,In_1326);
and U509 (N_509,In_327,In_1017);
and U510 (N_510,N_322,N_265);
xnor U511 (N_511,N_313,In_911);
xnor U512 (N_512,In_669,In_1268);
or U513 (N_513,In_997,In_736);
or U514 (N_514,N_392,In_509);
xnor U515 (N_515,In_1319,N_419);
xor U516 (N_516,In_1329,N_236);
xnor U517 (N_517,N_246,In_690);
nand U518 (N_518,In_487,N_401);
nand U519 (N_519,In_533,N_390);
xor U520 (N_520,N_440,In_506);
or U521 (N_521,In_211,N_340);
and U522 (N_522,In_148,In_814);
nand U523 (N_523,N_400,In_703);
nand U524 (N_524,In_1447,In_1313);
nand U525 (N_525,In_1269,In_335);
or U526 (N_526,N_394,In_250);
or U527 (N_527,In_1492,In_702);
nand U528 (N_528,In_1095,In_1439);
nand U529 (N_529,In_743,N_202);
or U530 (N_530,In_756,N_260);
and U531 (N_531,In_410,In_391);
nand U532 (N_532,In_401,In_1315);
or U533 (N_533,N_137,In_218);
or U534 (N_534,In_1368,In_1079);
and U535 (N_535,In_666,In_734);
and U536 (N_536,In_1386,In_609);
nor U537 (N_537,In_572,In_910);
and U538 (N_538,In_1111,In_241);
nand U539 (N_539,In_1034,N_126);
or U540 (N_540,N_423,In_1287);
nor U541 (N_541,In_786,In_618);
xor U542 (N_542,In_484,In_636);
or U543 (N_543,N_125,In_1167);
nor U544 (N_544,N_336,In_1055);
or U545 (N_545,In_206,In_929);
and U546 (N_546,In_885,In_675);
nand U547 (N_547,N_0,In_1043);
nor U548 (N_548,N_298,In_334);
nand U549 (N_549,In_668,In_1136);
xnor U550 (N_550,In_429,In_890);
nand U551 (N_551,In_792,In_361);
or U552 (N_552,In_450,In_1480);
nor U553 (N_553,N_4,In_418);
nor U554 (N_554,In_815,N_96);
nand U555 (N_555,N_199,In_222);
and U556 (N_556,In_542,N_97);
nor U557 (N_557,In_913,In_976);
nor U558 (N_558,In_474,N_359);
nor U559 (N_559,N_54,In_1415);
or U560 (N_560,N_402,In_858);
nand U561 (N_561,In_769,N_428);
nor U562 (N_562,In_1296,In_748);
and U563 (N_563,N_200,In_508);
nand U564 (N_564,In_324,In_732);
nand U565 (N_565,In_345,N_351);
xor U566 (N_566,N_413,In_432);
or U567 (N_567,In_639,In_94);
and U568 (N_568,In_1224,N_306);
nor U569 (N_569,In_688,In_694);
nand U570 (N_570,In_725,N_51);
and U571 (N_571,N_128,In_1166);
nand U572 (N_572,In_1120,N_414);
and U573 (N_573,In_704,In_1397);
or U574 (N_574,In_1005,In_1244);
xnor U575 (N_575,In_881,N_397);
and U576 (N_576,N_117,In_292);
or U577 (N_577,In_226,In_64);
xnor U578 (N_578,In_656,In_1461);
and U579 (N_579,N_191,In_1146);
or U580 (N_580,N_377,In_1018);
nand U581 (N_581,In_707,In_1039);
or U582 (N_582,N_333,N_354);
xnor U583 (N_583,In_514,N_20);
nand U584 (N_584,In_1472,In_185);
and U585 (N_585,N_295,In_359);
nand U586 (N_586,N_441,In_314);
or U587 (N_587,In_1143,In_657);
or U588 (N_588,In_1,N_132);
or U589 (N_589,In_70,N_316);
nand U590 (N_590,In_948,N_396);
nand U591 (N_591,In_644,In_1351);
or U592 (N_592,In_566,In_1483);
nor U593 (N_593,In_343,In_626);
or U594 (N_594,In_441,N_218);
nor U595 (N_595,In_1437,In_354);
xnor U596 (N_596,In_1072,In_1434);
xor U597 (N_597,In_1395,In_409);
nand U598 (N_598,In_186,In_338);
and U599 (N_599,N_143,N_194);
nand U600 (N_600,In_12,N_393);
xor U601 (N_601,In_1151,In_1279);
nor U602 (N_602,In_28,N_376);
and U603 (N_603,In_624,In_896);
nor U604 (N_604,In_130,In_693);
and U605 (N_605,N_348,N_408);
nor U606 (N_606,In_1103,N_578);
nor U607 (N_607,N_221,In_333);
and U608 (N_608,In_729,In_331);
nand U609 (N_609,N_527,In_68);
or U610 (N_610,N_450,N_231);
nor U611 (N_611,In_1241,N_121);
and U612 (N_612,N_571,In_192);
nand U613 (N_613,In_1123,N_317);
nand U614 (N_614,N_379,In_1374);
or U615 (N_615,In_1323,In_955);
xor U616 (N_616,N_162,In_552);
nor U617 (N_617,N_134,In_92);
xor U618 (N_618,In_282,N_198);
and U619 (N_619,N_356,N_113);
or U620 (N_620,In_403,In_470);
xor U621 (N_621,N_504,In_141);
nor U622 (N_622,N_382,In_782);
or U623 (N_623,In_143,In_1153);
nor U624 (N_624,In_1254,In_276);
or U625 (N_625,N_458,N_311);
or U626 (N_626,N_485,In_591);
nand U627 (N_627,In_1132,N_339);
nand U628 (N_628,In_113,N_508);
and U629 (N_629,In_368,In_1024);
and U630 (N_630,In_779,N_309);
nor U631 (N_631,N_569,N_580);
and U632 (N_632,N_18,In_385);
and U633 (N_633,In_422,N_360);
xnor U634 (N_634,N_577,N_551);
and U635 (N_635,N_451,N_192);
nor U636 (N_636,N_268,In_1338);
nand U637 (N_637,In_499,In_930);
or U638 (N_638,N_179,In_472);
nand U639 (N_639,In_1234,N_587);
nor U640 (N_640,N_28,N_373);
nand U641 (N_641,N_163,In_1198);
xnor U642 (N_642,N_93,In_838);
nor U643 (N_643,In_776,N_549);
nor U644 (N_644,N_288,N_522);
nor U645 (N_645,In_1219,In_1272);
and U646 (N_646,N_464,In_169);
or U647 (N_647,In_866,N_417);
xor U648 (N_648,In_633,In_1333);
nand U649 (N_649,In_1398,In_578);
nor U650 (N_650,N_352,In_91);
or U651 (N_651,In_26,In_394);
nor U652 (N_652,N_248,N_307);
xor U653 (N_653,In_860,N_335);
xor U654 (N_654,In_316,N_77);
and U655 (N_655,N_540,N_243);
nand U656 (N_656,In_456,N_206);
xnor U657 (N_657,In_131,N_449);
and U658 (N_658,N_244,N_521);
nand U659 (N_659,In_537,N_553);
nor U660 (N_660,N_594,In_1109);
or U661 (N_661,In_1496,In_1409);
nor U662 (N_662,In_234,In_532);
xor U663 (N_663,In_325,In_144);
or U664 (N_664,In_805,In_1113);
nand U665 (N_665,In_293,In_1373);
or U666 (N_666,N_545,N_537);
nand U667 (N_667,In_263,In_921);
nand U668 (N_668,In_313,N_523);
and U669 (N_669,In_1099,In_371);
nor U670 (N_670,In_662,In_225);
nand U671 (N_671,In_232,N_237);
xnor U672 (N_672,In_413,In_720);
nand U673 (N_673,N_363,In_568);
xnor U674 (N_674,N_465,In_1454);
nand U675 (N_675,In_182,In_84);
nand U676 (N_676,In_1139,In_679);
and U677 (N_677,In_42,In_184);
nand U678 (N_678,In_1490,In_77);
and U679 (N_679,N_287,In_1460);
and U680 (N_680,N_323,In_88);
and U681 (N_681,In_356,N_557);
nor U682 (N_682,N_576,In_166);
and U683 (N_683,In_118,N_479);
or U684 (N_684,In_160,In_797);
xor U685 (N_685,N_169,In_286);
xor U686 (N_686,N_380,In_434);
xor U687 (N_687,N_229,In_227);
nand U688 (N_688,In_1358,N_496);
xor U689 (N_689,N_431,N_34);
or U690 (N_690,In_4,N_149);
or U691 (N_691,In_179,N_476);
nor U692 (N_692,N_70,N_562);
nand U693 (N_693,N_130,N_473);
nand U694 (N_694,In_74,In_1067);
xnor U695 (N_695,N_326,N_536);
xnor U696 (N_696,In_318,In_54);
xnor U697 (N_697,In_560,In_602);
nor U698 (N_698,N_568,N_168);
and U699 (N_699,In_663,In_1427);
and U700 (N_700,In_1435,N_561);
or U701 (N_701,N_490,In_103);
nor U702 (N_702,N_371,N_207);
nor U703 (N_703,N_156,In_1497);
nor U704 (N_704,In_738,In_599);
and U705 (N_705,N_258,In_764);
or U706 (N_706,N_314,N_456);
nand U707 (N_707,N_489,N_487);
nand U708 (N_708,In_172,In_1105);
nor U709 (N_709,In_20,In_237);
xor U710 (N_710,N_572,In_909);
or U711 (N_711,In_119,N_403);
xor U712 (N_712,In_1228,N_593);
xor U713 (N_713,N_447,N_483);
xor U714 (N_714,In_872,N_386);
xnor U715 (N_715,N_599,In_1121);
nor U716 (N_716,In_522,N_596);
xor U717 (N_717,N_528,In_197);
or U718 (N_718,N_110,In_701);
xnor U719 (N_719,N_43,N_209);
and U720 (N_720,N_484,In_1375);
or U721 (N_721,In_411,In_1239);
and U722 (N_722,N_89,N_296);
and U723 (N_723,In_1458,N_269);
nand U724 (N_724,N_510,In_398);
and U725 (N_725,In_374,N_470);
nor U726 (N_726,In_919,N_247);
or U727 (N_727,N_409,N_437);
or U728 (N_728,N_430,In_1180);
nand U729 (N_729,N_155,In_558);
nand U730 (N_730,N_538,N_303);
xnor U731 (N_731,In_1141,In_1390);
and U732 (N_732,N_277,N_385);
or U733 (N_733,N_107,In_1040);
nand U734 (N_734,In_865,In_741);
xor U735 (N_735,N_45,In_303);
and U736 (N_736,In_907,In_1048);
or U737 (N_737,In_777,N_173);
nand U738 (N_738,In_1223,N_83);
nand U739 (N_739,N_29,In_254);
and U740 (N_740,In_1388,In_1248);
nor U741 (N_741,N_11,In_1371);
and U742 (N_742,In_251,In_1002);
or U743 (N_743,In_623,N_407);
or U744 (N_744,N_525,In_1170);
xor U745 (N_745,In_33,In_1330);
or U746 (N_746,In_1247,N_498);
nor U747 (N_747,N_475,In_17);
xnor U748 (N_748,In_1013,In_988);
nor U749 (N_749,In_863,N_548);
xnor U750 (N_750,N_628,In_216);
or U751 (N_751,N_272,In_874);
xor U752 (N_752,N_556,In_445);
and U753 (N_753,N_418,N_604);
xnor U754 (N_754,N_629,N_445);
or U755 (N_755,N_129,N_645);
nor U756 (N_756,N_364,In_877);
nor U757 (N_757,N_727,N_613);
xnor U758 (N_758,In_1114,In_3);
or U759 (N_759,N_575,N_453);
and U760 (N_760,N_144,In_571);
or U761 (N_761,N_555,N_602);
and U762 (N_762,N_358,In_582);
and U763 (N_763,In_665,In_252);
and U764 (N_764,N_318,In_1031);
and U765 (N_765,N_350,N_435);
nand U766 (N_766,N_399,In_518);
xor U767 (N_767,In_128,N_15);
and U768 (N_768,N_582,In_1281);
nor U769 (N_769,N_506,N_341);
nand U770 (N_770,N_542,In_1100);
nand U771 (N_771,N_387,N_444);
nor U772 (N_772,N_22,In_617);
or U773 (N_773,In_1227,N_480);
and U774 (N_774,In_692,In_683);
or U775 (N_775,In_1274,In_1207);
and U776 (N_776,In_886,In_653);
or U777 (N_777,N_325,N_80);
and U778 (N_778,In_295,In_1443);
xor U779 (N_779,N_598,N_225);
nand U780 (N_780,N_454,In_530);
nor U781 (N_781,N_726,N_452);
and U782 (N_782,In_632,In_479);
nor U783 (N_783,In_1310,N_74);
and U784 (N_784,In_563,In_1470);
and U785 (N_785,N_201,N_516);
and U786 (N_786,In_1160,In_900);
or U787 (N_787,N_671,In_66);
xnor U788 (N_788,N_500,N_560);
xnor U789 (N_789,N_205,N_714);
or U790 (N_790,N_514,N_566);
or U791 (N_791,N_337,In_106);
and U792 (N_792,N_279,N_94);
nor U793 (N_793,In_294,N_366);
or U794 (N_794,In_369,In_1213);
nand U795 (N_795,N_291,N_650);
and U796 (N_796,N_6,N_639);
or U797 (N_797,N_211,N_672);
nand U798 (N_798,In_202,In_140);
or U799 (N_799,In_501,N_503);
xor U800 (N_800,N_461,N_109);
and U801 (N_801,In_940,In_584);
xnor U802 (N_802,N_711,In_375);
nand U803 (N_803,In_1221,N_175);
or U804 (N_804,In_1422,N_180);
or U805 (N_805,In_816,In_857);
or U806 (N_806,N_438,In_258);
or U807 (N_807,N_600,In_771);
nor U808 (N_808,In_652,In_1273);
nor U809 (N_809,N_320,N_730);
nand U810 (N_810,In_1157,N_706);
nand U811 (N_811,In_240,In_1108);
or U812 (N_812,In_718,In_810);
or U813 (N_813,In_45,In_672);
or U814 (N_814,In_983,N_362);
nor U815 (N_815,In_32,In_674);
or U816 (N_816,N_667,In_1431);
and U817 (N_817,N_491,N_235);
xnor U818 (N_818,N_8,N_513);
xor U819 (N_819,In_1476,N_448);
nor U820 (N_820,N_460,In_497);
nor U821 (N_821,N_278,N_135);
xor U822 (N_822,In_97,N_655);
nor U823 (N_823,N_46,N_404);
and U824 (N_824,In_535,N_232);
xor U825 (N_825,N_656,N_632);
or U826 (N_826,N_328,N_304);
nand U827 (N_827,N_668,N_446);
nor U828 (N_828,In_1183,In_460);
and U829 (N_829,N_634,N_738);
and U830 (N_830,N_736,N_731);
or U831 (N_831,N_515,In_888);
nand U832 (N_832,In_305,N_625);
or U833 (N_833,In_180,N_517);
xor U834 (N_834,In_1314,N_241);
or U835 (N_835,N_676,N_374);
nand U836 (N_836,N_694,In_839);
nand U837 (N_837,In_363,In_579);
nor U838 (N_838,In_1499,N_182);
nor U839 (N_839,N_215,In_165);
and U840 (N_840,N_718,N_222);
nand U841 (N_841,N_626,In_1401);
or U842 (N_842,N_108,In_1142);
and U843 (N_843,N_471,N_357);
or U844 (N_844,In_126,In_173);
nand U845 (N_845,N_518,N_405);
and U846 (N_846,In_726,N_35);
nor U847 (N_847,N_308,N_466);
and U848 (N_848,In_221,In_915);
xnor U849 (N_849,N_734,N_633);
or U850 (N_850,N_338,N_84);
and U851 (N_851,N_747,N_737);
nor U852 (N_852,In_297,N_90);
and U853 (N_853,In_1030,N_695);
and U854 (N_854,N_220,In_1243);
or U855 (N_855,N_36,N_123);
nor U856 (N_856,N_647,N_327);
xnor U857 (N_857,N_98,N_744);
and U858 (N_858,In_1406,N_627);
nor U859 (N_859,In_220,In_217);
nand U860 (N_860,N_330,N_443);
or U861 (N_861,In_567,In_772);
or U862 (N_862,N_708,In_1124);
nand U863 (N_863,N_214,N_590);
nor U864 (N_864,N_203,N_618);
nand U865 (N_865,N_601,In_831);
and U866 (N_866,In_824,N_410);
or U867 (N_867,N_111,N_492);
nor U868 (N_868,N_240,N_709);
or U869 (N_869,N_167,N_728);
nand U870 (N_870,N_457,In_953);
or U871 (N_871,N_369,N_505);
or U872 (N_872,In_714,N_432);
xnor U873 (N_873,N_55,In_1408);
nor U874 (N_874,In_546,N_620);
and U875 (N_875,N_116,N_299);
xnor U876 (N_876,N_720,In_963);
xor U877 (N_877,N_597,N_270);
and U878 (N_878,In_965,N_381);
nand U879 (N_879,N_50,In_788);
nor U880 (N_880,N_106,In_270);
nand U881 (N_881,N_653,N_17);
or U882 (N_882,In_778,In_1384);
xnor U883 (N_883,In_283,In_145);
nor U884 (N_884,In_611,N_529);
xor U885 (N_885,N_591,N_406);
xnor U886 (N_886,N_666,N_91);
nor U887 (N_887,In_1012,In_1175);
nor U888 (N_888,In_1477,In_1436);
nand U889 (N_889,N_748,N_285);
or U890 (N_890,N_670,N_697);
nor U891 (N_891,N_550,N_115);
or U892 (N_892,N_319,In_307);
and U893 (N_893,In_1360,In_1346);
nand U894 (N_894,N_654,In_906);
or U895 (N_895,N_644,In_740);
nor U896 (N_896,N_422,In_175);
nand U897 (N_897,In_781,In_492);
xnor U898 (N_898,In_784,N_368);
nand U899 (N_899,In_556,N_60);
and U900 (N_900,N_67,N_674);
nor U901 (N_901,N_534,N_552);
xnor U902 (N_902,N_843,N_161);
and U903 (N_903,N_783,In_433);
nor U904 (N_904,N_785,In_1182);
nor U905 (N_905,N_693,In_266);
and U906 (N_906,N_740,N_349);
nand U907 (N_907,In_124,In_243);
and U908 (N_908,In_1263,N_468);
nand U909 (N_909,N_38,N_520);
or U910 (N_910,In_880,N_784);
nand U911 (N_911,N_868,N_539);
or U912 (N_912,N_831,In_1045);
and U913 (N_913,N_253,N_331);
nand U914 (N_914,N_332,In_773);
and U915 (N_915,N_226,N_426);
or U916 (N_916,N_512,N_690);
nor U917 (N_917,In_24,N_563);
and U918 (N_918,In_337,N_606);
or U919 (N_919,In_661,In_931);
nor U920 (N_920,In_1126,N_689);
nand U921 (N_921,N_7,In_408);
nor U922 (N_922,N_691,N_680);
or U923 (N_923,In_959,N_669);
or U924 (N_924,N_879,In_224);
nor U925 (N_925,In_279,N_355);
nand U926 (N_926,N_558,In_1450);
or U927 (N_927,In_507,N_157);
nor U928 (N_928,N_554,In_89);
xor U929 (N_929,In_1336,In_868);
and U930 (N_930,N_716,In_1107);
and U931 (N_931,In_306,N_802);
or U932 (N_932,N_830,N_751);
nor U933 (N_933,N_502,N_733);
or U934 (N_934,N_849,In_1007);
xnor U935 (N_935,N_488,N_699);
nor U936 (N_936,In_728,N_455);
nor U937 (N_937,N_790,N_859);
nor U938 (N_938,N_251,N_725);
and U939 (N_939,N_702,N_894);
nor U940 (N_940,N_884,In_587);
and U941 (N_941,N_780,N_823);
nor U942 (N_942,In_834,In_1407);
or U943 (N_943,In_1028,N_592);
and U944 (N_944,N_245,N_833);
nand U945 (N_945,N_615,N_547);
xor U946 (N_946,In_603,N_658);
and U947 (N_947,N_133,N_605);
xor U948 (N_948,N_703,In_1148);
xor U949 (N_949,N_217,In_1324);
xnor U950 (N_950,N_759,N_760);
nor U951 (N_951,In_1403,In_711);
nor U952 (N_952,N_721,In_1236);
or U953 (N_953,N_885,N_588);
nor U954 (N_954,In_195,N_384);
nor U955 (N_955,N_467,N_624);
or U956 (N_956,N_752,N_813);
nand U957 (N_957,N_573,N_698);
nor U958 (N_958,N_878,N_797);
xor U959 (N_959,N_638,N_678);
nor U960 (N_960,N_809,N_846);
xnor U961 (N_961,N_607,N_685);
xor U962 (N_962,N_874,N_700);
or U963 (N_963,In_0,N_353);
and U964 (N_964,N_769,N_616);
nand U965 (N_965,N_804,In_873);
and U966 (N_966,N_570,N_757);
nor U967 (N_967,In_274,N_741);
nand U968 (N_968,N_798,N_687);
and U969 (N_969,N_818,N_415);
nor U970 (N_970,N_775,In_65);
and U971 (N_971,N_746,N_442);
xnor U972 (N_972,In_1187,In_1445);
or U973 (N_973,N_729,In_342);
or U974 (N_974,N_819,N_880);
and U975 (N_975,In_419,N_439);
and U976 (N_976,In_1404,In_564);
xor U977 (N_977,N_772,N_779);
nand U978 (N_978,N_835,N_789);
xor U979 (N_979,N_829,In_989);
or U980 (N_980,In_966,N_824);
xor U981 (N_981,N_756,N_660);
and U982 (N_982,In_1255,In_105);
or U983 (N_983,N_595,N_637);
and U984 (N_984,In_146,N_329);
or U985 (N_985,N_887,In_1185);
and U986 (N_986,N_640,In_859);
and U987 (N_987,N_223,In_1297);
nand U988 (N_988,N_799,N_302);
or U989 (N_989,In_573,N_701);
or U990 (N_990,N_425,In_58);
nand U991 (N_991,In_851,N_888);
and U992 (N_992,N_614,N_621);
and U993 (N_993,In_1122,N_864);
xnor U994 (N_994,N_792,N_586);
or U995 (N_995,N_367,In_1393);
nand U996 (N_996,N_742,In_405);
nand U997 (N_997,N_531,In_793);
and U998 (N_998,N_800,In_449);
and U999 (N_999,N_463,In_807);
nor U1000 (N_1000,N_803,N_541);
nand U1001 (N_1001,N_766,N_712);
nand U1002 (N_1002,N_657,N_682);
xor U1003 (N_1003,N_895,N_519);
and U1004 (N_1004,N_543,In_1327);
xnor U1005 (N_1005,N_583,In_604);
nand U1006 (N_1006,N_482,N_750);
xnor U1007 (N_1007,In_176,In_1432);
or U1008 (N_1008,N_836,In_339);
xnor U1009 (N_1009,N_481,In_1215);
and U1010 (N_1010,In_523,N_872);
or U1011 (N_1011,In_1349,N_858);
and U1012 (N_1012,N_429,In_1037);
nand U1013 (N_1013,N_891,In_1416);
or U1014 (N_1014,In_488,In_747);
and U1015 (N_1015,In_102,N_659);
or U1016 (N_1016,N_494,N_795);
xnor U1017 (N_1017,In_57,In_648);
xnor U1018 (N_1018,N_893,In_783);
or U1019 (N_1019,N_56,N_898);
nor U1020 (N_1020,In_163,In_75);
nand U1021 (N_1021,N_524,N_641);
and U1022 (N_1022,N_826,N_873);
and U1023 (N_1023,N_840,In_975);
and U1024 (N_1024,N_762,In_25);
nand U1025 (N_1025,N_346,In_1489);
and U1026 (N_1026,N_233,N_427);
xor U1027 (N_1027,In_864,N_814);
nand U1028 (N_1028,N_239,N_193);
nor U1029 (N_1029,In_882,N_391);
xnor U1030 (N_1030,N_739,N_497);
xor U1031 (N_1031,N_673,In_1240);
xnor U1032 (N_1032,N_724,N_343);
nor U1033 (N_1033,N_683,N_870);
nor U1034 (N_1034,N_839,In_800);
or U1035 (N_1035,In_1391,N_665);
nand U1036 (N_1036,N_652,N_692);
nand U1037 (N_1037,In_271,In_739);
nor U1038 (N_1038,In_968,N_636);
or U1039 (N_1039,In_473,N_877);
or U1040 (N_1040,N_875,N_677);
and U1041 (N_1041,N_663,In_1068);
and U1042 (N_1042,In_920,N_623);
and U1043 (N_1043,In_423,N_170);
nand U1044 (N_1044,N_754,N_662);
xor U1045 (N_1045,N_684,N_882);
and U1046 (N_1046,N_735,N_822);
or U1047 (N_1047,N_794,N_617);
xnor U1048 (N_1048,In_1196,In_321);
nand U1049 (N_1049,N_853,N_765);
or U1050 (N_1050,N_773,N_1017);
xnor U1051 (N_1051,In_34,N_758);
xnor U1052 (N_1052,N_704,N_183);
and U1053 (N_1053,N_948,N_854);
or U1054 (N_1054,N_286,N_764);
nor U1055 (N_1055,In_1337,In_1087);
nor U1056 (N_1056,In_1280,N_723);
or U1057 (N_1057,In_826,N_324);
nor U1058 (N_1058,N_984,N_459);
and U1059 (N_1059,N_812,N_974);
nand U1060 (N_1060,N_389,N_908);
nor U1061 (N_1061,N_782,N_119);
and U1062 (N_1062,N_832,N_941);
nor U1063 (N_1063,N_361,In_1299);
and U1064 (N_1064,N_646,N_184);
nand U1065 (N_1065,N_844,N_862);
or U1066 (N_1066,N_584,N_904);
nor U1067 (N_1067,In_540,N_57);
and U1068 (N_1068,N_533,N_983);
xor U1069 (N_1069,N_424,N_890);
xor U1070 (N_1070,N_856,N_907);
nor U1071 (N_1071,N_970,In_576);
and U1072 (N_1072,N_935,N_1001);
nor U1073 (N_1073,N_883,N_960);
xnor U1074 (N_1074,N_850,N_828);
nand U1075 (N_1075,N_1049,In_1206);
xor U1076 (N_1076,N_1006,N_713);
nor U1077 (N_1077,N_151,N_911);
or U1078 (N_1078,N_1035,N_462);
nand U1079 (N_1079,In_716,In_676);
or U1080 (N_1080,In_443,N_937);
and U1081 (N_1081,In_1357,N_398);
xnor U1082 (N_1082,In_1001,N_501);
nand U1083 (N_1083,N_651,N_661);
nand U1084 (N_1084,N_1026,N_947);
or U1085 (N_1085,In_828,In_1203);
xor U1086 (N_1086,N_923,N_965);
nand U1087 (N_1087,N_915,N_889);
nor U1088 (N_1088,In_228,In_190);
nand U1089 (N_1089,N_421,N_378);
or U1090 (N_1090,In_1208,N_589);
nor U1091 (N_1091,N_997,N_778);
xor U1092 (N_1092,In_80,N_585);
xor U1093 (N_1093,In_452,N_383);
nand U1094 (N_1094,N_929,N_477);
and U1095 (N_1095,N_1042,N_950);
and U1096 (N_1096,N_851,N_901);
xor U1097 (N_1097,N_902,In_1339);
nand U1098 (N_1098,In_970,N_630);
xor U1099 (N_1099,N_912,N_32);
nand U1100 (N_1100,N_228,N_95);
and U1101 (N_1101,N_991,N_707);
nand U1102 (N_1102,N_648,N_881);
xor U1103 (N_1103,In_100,In_1238);
and U1104 (N_1104,N_909,N_567);
or U1105 (N_1105,In_590,N_897);
or U1106 (N_1106,N_1021,N_924);
nor U1107 (N_1107,N_293,N_966);
nor U1108 (N_1108,N_375,N_838);
nor U1109 (N_1109,N_474,In_516);
nor U1110 (N_1110,N_544,N_917);
or U1111 (N_1111,N_949,N_943);
or U1112 (N_1112,N_282,In_101);
or U1113 (N_1113,N_1012,In_284);
nand U1114 (N_1114,N_913,In_336);
or U1115 (N_1115,N_914,N_753);
and U1116 (N_1116,N_69,N_953);
nand U1117 (N_1117,N_942,In_236);
or U1118 (N_1118,In_855,In_849);
nor U1119 (N_1119,N_611,N_886);
and U1120 (N_1120,N_925,N_867);
xnor U1121 (N_1121,In_420,N_982);
or U1122 (N_1122,N_964,N_972);
xnor U1123 (N_1123,In_733,N_1003);
nand U1124 (N_1124,N_786,In_244);
xnor U1125 (N_1125,N_939,N_252);
xor U1126 (N_1126,N_1041,N_848);
nor U1127 (N_1127,N_857,In_765);
nor U1128 (N_1128,In_1009,N_918);
xnor U1129 (N_1129,N_951,In_946);
nor U1130 (N_1130,N_1031,In_654);
nand U1131 (N_1131,N_934,N_808);
and U1132 (N_1132,In_1410,N_952);
nor U1133 (N_1133,N_342,N_810);
or U1134 (N_1134,N_841,N_1016);
or U1135 (N_1135,N_159,N_234);
or U1136 (N_1136,N_852,N_834);
and U1137 (N_1137,N_827,N_688);
nor U1138 (N_1138,N_847,N_933);
nand U1139 (N_1139,N_990,N_936);
nand U1140 (N_1140,N_1044,In_6);
xor U1141 (N_1141,N_986,N_1020);
or U1142 (N_1142,N_82,N_985);
or U1143 (N_1143,N_643,N_681);
nor U1144 (N_1144,N_987,N_1014);
or U1145 (N_1145,N_187,N_928);
and U1146 (N_1146,N_732,N_526);
and U1147 (N_1147,N_821,In_204);
or U1148 (N_1148,N_805,N_820);
nand U1149 (N_1149,N_511,N_749);
and U1150 (N_1150,N_1040,N_994);
and U1151 (N_1151,N_1048,In_996);
and U1152 (N_1152,N_581,N_274);
xor U1153 (N_1153,N_62,N_1024);
and U1154 (N_1154,N_105,N_530);
nor U1155 (N_1155,N_609,N_1009);
xor U1156 (N_1156,In_641,N_412);
xor U1157 (N_1157,N_1027,In_121);
nand U1158 (N_1158,N_921,N_1036);
nor U1159 (N_1159,N_675,In_428);
and U1160 (N_1160,N_866,N_816);
or U1161 (N_1161,N_876,N_993);
nand U1162 (N_1162,In_1303,In_494);
xor U1163 (N_1163,N_971,In_1058);
and U1164 (N_1164,In_440,N_979);
or U1165 (N_1165,N_996,In_457);
xnor U1166 (N_1166,In_597,N_975);
or U1167 (N_1167,N_1022,In_1372);
nor U1168 (N_1168,N_981,N_493);
xnor U1169 (N_1169,N_1038,N_256);
xor U1170 (N_1170,N_787,N_290);
xor U1171 (N_1171,N_469,N_845);
nand U1172 (N_1172,N_1008,In_894);
xnor U1173 (N_1173,N_869,N_301);
or U1174 (N_1174,N_903,N_166);
or U1175 (N_1175,In_559,N_59);
or U1176 (N_1176,N_767,N_370);
or U1177 (N_1177,N_499,In_1061);
or U1178 (N_1178,N_1034,N_686);
nand U1179 (N_1179,In_622,N_961);
xnor U1180 (N_1180,In_1428,N_926);
nor U1181 (N_1181,N_1033,N_777);
nand U1182 (N_1182,N_980,N_956);
xnor U1183 (N_1183,In_15,N_292);
or U1184 (N_1184,N_478,In_193);
xor U1185 (N_1185,N_969,In_138);
nand U1186 (N_1186,N_978,N_719);
xor U1187 (N_1187,In_794,N_321);
xnor U1188 (N_1188,N_998,N_1005);
xnor U1189 (N_1189,N_768,N_1043);
or U1190 (N_1190,N_679,N_930);
nor U1191 (N_1191,N_955,N_559);
nor U1192 (N_1192,N_1000,N_865);
nor U1193 (N_1193,N_305,N_124);
nand U1194 (N_1194,N_761,N_992);
nand U1195 (N_1195,N_257,N_1045);
and U1196 (N_1196,N_959,N_1037);
or U1197 (N_1197,N_664,In_895);
xor U1198 (N_1198,N_284,N_300);
or U1199 (N_1199,N_815,N_954);
nand U1200 (N_1200,N_1134,N_1146);
nor U1201 (N_1201,N_1032,N_1172);
or U1202 (N_1202,In_589,N_871);
xnor U1203 (N_1203,N_1199,In_1070);
xor U1204 (N_1204,N_1129,N_900);
or U1205 (N_1205,N_1158,In_993);
or U1206 (N_1206,N_345,N_1063);
xnor U1207 (N_1207,N_1030,N_1190);
nand U1208 (N_1208,N_1023,In_1278);
or U1209 (N_1209,N_1093,N_811);
nor U1210 (N_1210,N_1067,N_938);
and U1211 (N_1211,N_1094,N_1053);
and U1212 (N_1212,N_433,In_1469);
nor U1213 (N_1213,N_1102,N_1140);
nor U1214 (N_1214,In_905,N_932);
nor U1215 (N_1215,N_906,N_1196);
and U1216 (N_1216,In_1253,N_1002);
nor U1217 (N_1217,N_1188,N_1055);
xor U1218 (N_1218,N_1100,N_892);
nor U1219 (N_1219,N_1056,N_774);
xnor U1220 (N_1220,In_201,N_1082);
and U1221 (N_1221,N_855,N_1039);
nor U1222 (N_1222,N_612,N_631);
xnor U1223 (N_1223,N_1123,N_1113);
nor U1224 (N_1224,N_1091,In_1418);
or U1225 (N_1225,N_1092,N_1083);
xnor U1226 (N_1226,In_311,N_1075);
and U1227 (N_1227,N_1046,N_1077);
nor U1228 (N_1228,N_860,N_1028);
or U1229 (N_1229,N_1098,N_495);
or U1230 (N_1230,N_1121,N_1173);
or U1231 (N_1231,N_931,In_1188);
or U1232 (N_1232,N_1114,N_1163);
xor U1233 (N_1233,N_1195,N_1192);
nand U1234 (N_1234,N_1115,N_842);
and U1235 (N_1235,N_619,N_715);
or U1236 (N_1236,N_1175,N_564);
nor U1237 (N_1237,N_1128,N_1178);
and U1238 (N_1238,N_717,N_31);
or U1239 (N_1239,N_283,N_1078);
or U1240 (N_1240,N_837,N_796);
and U1241 (N_1241,N_968,N_603);
nand U1242 (N_1242,N_574,N_1051);
and U1243 (N_1243,N_1150,N_999);
and U1244 (N_1244,N_896,N_1165);
and U1245 (N_1245,N_1097,N_944);
and U1246 (N_1246,N_771,N_946);
xor U1247 (N_1247,In_971,N_1193);
nand U1248 (N_1248,N_863,N_1066);
nand U1249 (N_1249,N_1015,N_120);
nor U1250 (N_1250,N_1139,N_1060);
or U1251 (N_1251,N_989,N_1111);
nand U1252 (N_1252,N_976,N_1174);
xor U1253 (N_1253,N_910,N_1068);
and U1254 (N_1254,N_807,In_1264);
and U1255 (N_1255,N_266,N_1180);
nor U1256 (N_1256,N_1166,In_489);
or U1257 (N_1257,N_138,N_197);
xnor U1258 (N_1258,In_1300,N_817);
or U1259 (N_1259,N_755,N_899);
nor U1260 (N_1260,N_649,N_1118);
and U1261 (N_1261,N_1061,N_1103);
nor U1262 (N_1262,N_622,N_945);
and U1263 (N_1263,N_344,N_988);
or U1264 (N_1264,N_1176,N_1155);
nor U1265 (N_1265,N_957,N_1096);
or U1266 (N_1266,N_1159,In_992);
or U1267 (N_1267,N_486,N_1029);
and U1268 (N_1268,N_1189,N_1057);
and U1269 (N_1269,N_1137,N_579);
or U1270 (N_1270,N_608,In_1162);
nor U1271 (N_1271,N_642,N_1161);
nor U1272 (N_1272,N_1141,N_1117);
nand U1273 (N_1273,N_1144,N_722);
or U1274 (N_1274,N_1164,N_1122);
nand U1275 (N_1275,N_1064,In_1102);
xor U1276 (N_1276,N_436,N_1127);
and U1277 (N_1277,N_781,In_453);
or U1278 (N_1278,In_1014,In_549);
nand U1279 (N_1279,N_535,In_322);
nor U1280 (N_1280,N_263,N_1151);
xnor U1281 (N_1281,N_1120,N_532);
xnor U1282 (N_1282,N_635,N_1145);
nor U1283 (N_1283,N_793,N_1126);
xnor U1284 (N_1284,N_1149,N_1105);
nand U1285 (N_1285,N_1110,N_1184);
nor U1286 (N_1286,N_776,N_1076);
xnor U1287 (N_1287,N_1177,N_472);
nor U1288 (N_1288,N_1050,N_1011);
or U1289 (N_1289,N_1080,N_745);
and U1290 (N_1290,N_1168,N_1054);
xor U1291 (N_1291,N_791,N_1079);
xor U1292 (N_1292,N_1152,N_919);
nand U1293 (N_1293,N_1047,N_1157);
nor U1294 (N_1294,N_1081,N_1090);
nor U1295 (N_1295,N_1133,N_763);
nand U1296 (N_1296,N_1085,N_1101);
xor U1297 (N_1297,N_967,N_1132);
nand U1298 (N_1298,N_806,N_1135);
xor U1299 (N_1299,N_940,N_1019);
or U1300 (N_1300,N_1147,In_1468);
nor U1301 (N_1301,N_347,N_1194);
xnor U1302 (N_1302,N_1073,N_267);
xnor U1303 (N_1303,N_995,N_1197);
and U1304 (N_1304,N_1071,N_1116);
nand U1305 (N_1305,N_1125,N_1104);
or U1306 (N_1306,N_861,N_610);
nor U1307 (N_1307,N_1167,N_1131);
nand U1308 (N_1308,N_963,N_1058);
nand U1309 (N_1309,N_1108,N_1185);
nor U1310 (N_1310,N_1065,In_380);
and U1311 (N_1311,N_1062,N_12);
or U1312 (N_1312,N_920,N_1013);
nand U1313 (N_1313,N_927,N_1086);
xnor U1314 (N_1314,N_1109,N_1010);
and U1315 (N_1315,In_671,N_1162);
nor U1316 (N_1316,N_509,N_565);
nor U1317 (N_1317,N_770,N_1181);
xnor U1318 (N_1318,N_546,N_1025);
nor U1319 (N_1319,N_1004,In_1115);
nor U1320 (N_1320,N_1112,In_594);
and U1321 (N_1321,N_977,N_1187);
nand U1322 (N_1322,N_1095,N_1148);
and U1323 (N_1323,N_743,N_1087);
or U1324 (N_1324,N_1130,N_973);
nand U1325 (N_1325,N_922,N_705);
nand U1326 (N_1326,N_916,N_1018);
nor U1327 (N_1327,N_1138,N_1136);
nand U1328 (N_1328,N_1052,N_1069);
and U1329 (N_1329,N_1106,N_696);
and U1330 (N_1330,N_905,In_1465);
and U1331 (N_1331,N_1160,N_1124);
nor U1332 (N_1332,N_788,N_1198);
or U1333 (N_1333,N_88,N_1169);
and U1334 (N_1334,N_825,N_801);
xor U1335 (N_1335,N_1007,N_1070);
nor U1336 (N_1336,N_1088,N_1099);
and U1337 (N_1337,N_1143,N_1119);
or U1338 (N_1338,N_1153,N_160);
nor U1339 (N_1339,N_1107,N_1186);
nand U1340 (N_1340,N_1182,N_1183);
nor U1341 (N_1341,N_1156,N_1142);
nand U1342 (N_1342,In_883,N_1089);
xor U1343 (N_1343,N_958,N_1072);
xnor U1344 (N_1344,N_1171,N_1154);
or U1345 (N_1345,N_507,N_1170);
nand U1346 (N_1346,N_1179,In_480);
xor U1347 (N_1347,N_710,N_1084);
xnor U1348 (N_1348,N_962,N_1191);
nor U1349 (N_1349,N_1074,N_1059);
nor U1350 (N_1350,N_1346,N_1287);
or U1351 (N_1351,N_1331,N_1236);
and U1352 (N_1352,N_1204,N_1223);
nor U1353 (N_1353,N_1263,N_1239);
and U1354 (N_1354,N_1318,N_1249);
nand U1355 (N_1355,N_1271,N_1290);
nand U1356 (N_1356,N_1269,N_1265);
nand U1357 (N_1357,N_1264,N_1222);
nand U1358 (N_1358,N_1225,N_1235);
nand U1359 (N_1359,N_1304,N_1319);
xor U1360 (N_1360,N_1343,N_1294);
and U1361 (N_1361,N_1254,N_1330);
or U1362 (N_1362,N_1293,N_1237);
and U1363 (N_1363,N_1207,N_1209);
nand U1364 (N_1364,N_1276,N_1257);
and U1365 (N_1365,N_1344,N_1274);
and U1366 (N_1366,N_1256,N_1255);
nor U1367 (N_1367,N_1252,N_1324);
xnor U1368 (N_1368,N_1266,N_1213);
nand U1369 (N_1369,N_1317,N_1312);
nand U1370 (N_1370,N_1268,N_1218);
nor U1371 (N_1371,N_1258,N_1342);
and U1372 (N_1372,N_1297,N_1285);
or U1373 (N_1373,N_1273,N_1212);
nand U1374 (N_1374,N_1250,N_1329);
or U1375 (N_1375,N_1248,N_1334);
xnor U1376 (N_1376,N_1201,N_1336);
and U1377 (N_1377,N_1205,N_1338);
or U1378 (N_1378,N_1227,N_1216);
nor U1379 (N_1379,N_1251,N_1314);
nand U1380 (N_1380,N_1291,N_1347);
and U1381 (N_1381,N_1206,N_1284);
nand U1382 (N_1382,N_1247,N_1322);
nor U1383 (N_1383,N_1337,N_1242);
nand U1384 (N_1384,N_1303,N_1217);
or U1385 (N_1385,N_1323,N_1226);
and U1386 (N_1386,N_1305,N_1241);
and U1387 (N_1387,N_1240,N_1260);
nand U1388 (N_1388,N_1210,N_1211);
xor U1389 (N_1389,N_1296,N_1325);
and U1390 (N_1390,N_1261,N_1214);
and U1391 (N_1391,N_1288,N_1326);
nand U1392 (N_1392,N_1219,N_1341);
xor U1393 (N_1393,N_1306,N_1327);
nand U1394 (N_1394,N_1308,N_1300);
and U1395 (N_1395,N_1215,N_1243);
nor U1396 (N_1396,N_1286,N_1229);
xor U1397 (N_1397,N_1224,N_1299);
xnor U1398 (N_1398,N_1281,N_1272);
xnor U1399 (N_1399,N_1253,N_1321);
nand U1400 (N_1400,N_1289,N_1280);
nor U1401 (N_1401,N_1233,N_1320);
and U1402 (N_1402,N_1283,N_1234);
nand U1403 (N_1403,N_1310,N_1339);
xnor U1404 (N_1404,N_1220,N_1275);
nand U1405 (N_1405,N_1246,N_1228);
nor U1406 (N_1406,N_1301,N_1333);
nor U1407 (N_1407,N_1262,N_1277);
and U1408 (N_1408,N_1309,N_1328);
nor U1409 (N_1409,N_1270,N_1298);
nand U1410 (N_1410,N_1302,N_1345);
xor U1411 (N_1411,N_1238,N_1282);
xnor U1412 (N_1412,N_1278,N_1292);
xnor U1413 (N_1413,N_1313,N_1340);
xnor U1414 (N_1414,N_1311,N_1200);
xor U1415 (N_1415,N_1208,N_1267);
nor U1416 (N_1416,N_1295,N_1202);
nor U1417 (N_1417,N_1307,N_1203);
or U1418 (N_1418,N_1232,N_1244);
nand U1419 (N_1419,N_1315,N_1348);
or U1420 (N_1420,N_1349,N_1259);
and U1421 (N_1421,N_1230,N_1245);
or U1422 (N_1422,N_1279,N_1335);
xnor U1423 (N_1423,N_1316,N_1221);
xor U1424 (N_1424,N_1231,N_1332);
nand U1425 (N_1425,N_1298,N_1211);
nand U1426 (N_1426,N_1217,N_1333);
xnor U1427 (N_1427,N_1242,N_1267);
nor U1428 (N_1428,N_1233,N_1239);
or U1429 (N_1429,N_1301,N_1257);
xor U1430 (N_1430,N_1290,N_1227);
nor U1431 (N_1431,N_1204,N_1298);
nor U1432 (N_1432,N_1234,N_1282);
nor U1433 (N_1433,N_1213,N_1317);
xnor U1434 (N_1434,N_1326,N_1319);
nor U1435 (N_1435,N_1214,N_1216);
or U1436 (N_1436,N_1291,N_1240);
and U1437 (N_1437,N_1203,N_1334);
or U1438 (N_1438,N_1322,N_1321);
or U1439 (N_1439,N_1292,N_1209);
and U1440 (N_1440,N_1223,N_1333);
and U1441 (N_1441,N_1205,N_1285);
nor U1442 (N_1442,N_1201,N_1253);
and U1443 (N_1443,N_1218,N_1225);
and U1444 (N_1444,N_1262,N_1291);
nand U1445 (N_1445,N_1211,N_1242);
xnor U1446 (N_1446,N_1230,N_1339);
nand U1447 (N_1447,N_1245,N_1278);
nor U1448 (N_1448,N_1278,N_1255);
or U1449 (N_1449,N_1276,N_1227);
or U1450 (N_1450,N_1218,N_1215);
and U1451 (N_1451,N_1251,N_1323);
xor U1452 (N_1452,N_1294,N_1252);
and U1453 (N_1453,N_1223,N_1312);
nand U1454 (N_1454,N_1311,N_1305);
xor U1455 (N_1455,N_1230,N_1272);
nand U1456 (N_1456,N_1309,N_1243);
or U1457 (N_1457,N_1333,N_1228);
or U1458 (N_1458,N_1250,N_1320);
nor U1459 (N_1459,N_1208,N_1326);
xor U1460 (N_1460,N_1241,N_1255);
nor U1461 (N_1461,N_1233,N_1319);
nand U1462 (N_1462,N_1320,N_1314);
and U1463 (N_1463,N_1278,N_1201);
nand U1464 (N_1464,N_1324,N_1346);
xor U1465 (N_1465,N_1284,N_1274);
nor U1466 (N_1466,N_1313,N_1348);
nand U1467 (N_1467,N_1258,N_1273);
nand U1468 (N_1468,N_1325,N_1260);
nor U1469 (N_1469,N_1270,N_1216);
nand U1470 (N_1470,N_1284,N_1283);
or U1471 (N_1471,N_1218,N_1273);
xnor U1472 (N_1472,N_1335,N_1201);
xnor U1473 (N_1473,N_1286,N_1273);
xnor U1474 (N_1474,N_1286,N_1260);
or U1475 (N_1475,N_1200,N_1341);
nand U1476 (N_1476,N_1263,N_1275);
and U1477 (N_1477,N_1261,N_1325);
xor U1478 (N_1478,N_1343,N_1287);
and U1479 (N_1479,N_1330,N_1216);
and U1480 (N_1480,N_1299,N_1216);
or U1481 (N_1481,N_1281,N_1291);
nor U1482 (N_1482,N_1291,N_1300);
xor U1483 (N_1483,N_1345,N_1260);
xnor U1484 (N_1484,N_1283,N_1342);
nor U1485 (N_1485,N_1274,N_1304);
and U1486 (N_1486,N_1283,N_1269);
nand U1487 (N_1487,N_1240,N_1233);
nor U1488 (N_1488,N_1261,N_1284);
nand U1489 (N_1489,N_1261,N_1269);
xor U1490 (N_1490,N_1240,N_1236);
or U1491 (N_1491,N_1236,N_1313);
xnor U1492 (N_1492,N_1268,N_1332);
xnor U1493 (N_1493,N_1282,N_1210);
nor U1494 (N_1494,N_1248,N_1217);
nor U1495 (N_1495,N_1340,N_1247);
or U1496 (N_1496,N_1348,N_1253);
xnor U1497 (N_1497,N_1335,N_1274);
nor U1498 (N_1498,N_1319,N_1318);
or U1499 (N_1499,N_1313,N_1235);
xor U1500 (N_1500,N_1492,N_1400);
xnor U1501 (N_1501,N_1352,N_1394);
and U1502 (N_1502,N_1459,N_1481);
or U1503 (N_1503,N_1429,N_1443);
nand U1504 (N_1504,N_1413,N_1447);
nand U1505 (N_1505,N_1361,N_1393);
nand U1506 (N_1506,N_1441,N_1367);
and U1507 (N_1507,N_1437,N_1427);
nor U1508 (N_1508,N_1353,N_1409);
or U1509 (N_1509,N_1499,N_1480);
nor U1510 (N_1510,N_1460,N_1381);
and U1511 (N_1511,N_1373,N_1478);
nand U1512 (N_1512,N_1363,N_1425);
xnor U1513 (N_1513,N_1479,N_1490);
nor U1514 (N_1514,N_1396,N_1484);
xnor U1515 (N_1515,N_1466,N_1389);
and U1516 (N_1516,N_1464,N_1406);
or U1517 (N_1517,N_1402,N_1370);
nor U1518 (N_1518,N_1401,N_1374);
nand U1519 (N_1519,N_1412,N_1472);
nor U1520 (N_1520,N_1485,N_1498);
nor U1521 (N_1521,N_1390,N_1392);
nand U1522 (N_1522,N_1365,N_1428);
xnor U1523 (N_1523,N_1458,N_1491);
xor U1524 (N_1524,N_1436,N_1358);
or U1525 (N_1525,N_1475,N_1493);
or U1526 (N_1526,N_1430,N_1391);
and U1527 (N_1527,N_1372,N_1462);
or U1528 (N_1528,N_1465,N_1411);
nand U1529 (N_1529,N_1482,N_1467);
xor U1530 (N_1530,N_1356,N_1453);
nand U1531 (N_1531,N_1420,N_1378);
or U1532 (N_1532,N_1380,N_1446);
nand U1533 (N_1533,N_1438,N_1452);
nor U1534 (N_1534,N_1422,N_1359);
nor U1535 (N_1535,N_1410,N_1404);
xor U1536 (N_1536,N_1399,N_1483);
nor U1537 (N_1537,N_1377,N_1355);
xnor U1538 (N_1538,N_1418,N_1494);
nor U1539 (N_1539,N_1432,N_1360);
nor U1540 (N_1540,N_1371,N_1445);
and U1541 (N_1541,N_1468,N_1486);
and U1542 (N_1542,N_1397,N_1385);
and U1543 (N_1543,N_1379,N_1423);
and U1544 (N_1544,N_1461,N_1398);
and U1545 (N_1545,N_1419,N_1449);
nor U1546 (N_1546,N_1471,N_1434);
or U1547 (N_1547,N_1444,N_1414);
or U1548 (N_1548,N_1448,N_1488);
nand U1549 (N_1549,N_1382,N_1439);
xor U1550 (N_1550,N_1388,N_1426);
or U1551 (N_1551,N_1497,N_1416);
or U1552 (N_1552,N_1431,N_1408);
nand U1553 (N_1553,N_1407,N_1433);
nand U1554 (N_1554,N_1487,N_1376);
nor U1555 (N_1555,N_1421,N_1366);
xor U1556 (N_1556,N_1369,N_1384);
xnor U1557 (N_1557,N_1450,N_1354);
nor U1558 (N_1558,N_1417,N_1489);
and U1559 (N_1559,N_1477,N_1424);
xnor U1560 (N_1560,N_1368,N_1387);
nor U1561 (N_1561,N_1403,N_1435);
or U1562 (N_1562,N_1375,N_1362);
or U1563 (N_1563,N_1386,N_1454);
nor U1564 (N_1564,N_1364,N_1442);
or U1565 (N_1565,N_1470,N_1474);
nor U1566 (N_1566,N_1496,N_1469);
nor U1567 (N_1567,N_1351,N_1350);
nor U1568 (N_1568,N_1357,N_1476);
and U1569 (N_1569,N_1440,N_1395);
and U1570 (N_1570,N_1457,N_1415);
nor U1571 (N_1571,N_1463,N_1473);
nand U1572 (N_1572,N_1451,N_1405);
nor U1573 (N_1573,N_1495,N_1383);
xor U1574 (N_1574,N_1455,N_1456);
nor U1575 (N_1575,N_1478,N_1495);
and U1576 (N_1576,N_1444,N_1468);
or U1577 (N_1577,N_1465,N_1419);
and U1578 (N_1578,N_1462,N_1484);
nand U1579 (N_1579,N_1466,N_1395);
nand U1580 (N_1580,N_1369,N_1399);
xor U1581 (N_1581,N_1444,N_1459);
and U1582 (N_1582,N_1451,N_1378);
nor U1583 (N_1583,N_1476,N_1450);
or U1584 (N_1584,N_1489,N_1440);
xor U1585 (N_1585,N_1497,N_1406);
nand U1586 (N_1586,N_1403,N_1436);
and U1587 (N_1587,N_1439,N_1360);
nand U1588 (N_1588,N_1458,N_1497);
xor U1589 (N_1589,N_1368,N_1495);
and U1590 (N_1590,N_1359,N_1473);
nor U1591 (N_1591,N_1448,N_1378);
or U1592 (N_1592,N_1445,N_1456);
nor U1593 (N_1593,N_1368,N_1438);
and U1594 (N_1594,N_1415,N_1485);
and U1595 (N_1595,N_1469,N_1444);
and U1596 (N_1596,N_1354,N_1395);
nor U1597 (N_1597,N_1390,N_1389);
and U1598 (N_1598,N_1426,N_1411);
and U1599 (N_1599,N_1479,N_1394);
and U1600 (N_1600,N_1424,N_1354);
xnor U1601 (N_1601,N_1432,N_1400);
nand U1602 (N_1602,N_1386,N_1451);
xor U1603 (N_1603,N_1359,N_1483);
nor U1604 (N_1604,N_1458,N_1447);
or U1605 (N_1605,N_1374,N_1456);
xnor U1606 (N_1606,N_1444,N_1405);
nand U1607 (N_1607,N_1439,N_1428);
nand U1608 (N_1608,N_1360,N_1352);
nand U1609 (N_1609,N_1384,N_1359);
and U1610 (N_1610,N_1497,N_1367);
nor U1611 (N_1611,N_1363,N_1458);
nand U1612 (N_1612,N_1377,N_1409);
and U1613 (N_1613,N_1406,N_1484);
nor U1614 (N_1614,N_1394,N_1365);
nand U1615 (N_1615,N_1477,N_1487);
xor U1616 (N_1616,N_1491,N_1381);
or U1617 (N_1617,N_1372,N_1416);
and U1618 (N_1618,N_1471,N_1424);
xnor U1619 (N_1619,N_1477,N_1413);
nand U1620 (N_1620,N_1375,N_1499);
or U1621 (N_1621,N_1470,N_1453);
or U1622 (N_1622,N_1495,N_1392);
nor U1623 (N_1623,N_1488,N_1464);
nor U1624 (N_1624,N_1491,N_1468);
or U1625 (N_1625,N_1494,N_1351);
or U1626 (N_1626,N_1372,N_1383);
or U1627 (N_1627,N_1454,N_1481);
xor U1628 (N_1628,N_1366,N_1489);
or U1629 (N_1629,N_1457,N_1401);
or U1630 (N_1630,N_1467,N_1450);
or U1631 (N_1631,N_1355,N_1488);
xor U1632 (N_1632,N_1444,N_1420);
xor U1633 (N_1633,N_1420,N_1493);
xnor U1634 (N_1634,N_1389,N_1427);
nor U1635 (N_1635,N_1455,N_1351);
and U1636 (N_1636,N_1401,N_1447);
nand U1637 (N_1637,N_1468,N_1472);
nor U1638 (N_1638,N_1369,N_1370);
xor U1639 (N_1639,N_1350,N_1452);
nor U1640 (N_1640,N_1425,N_1483);
or U1641 (N_1641,N_1499,N_1492);
or U1642 (N_1642,N_1419,N_1396);
nor U1643 (N_1643,N_1463,N_1355);
nand U1644 (N_1644,N_1423,N_1494);
and U1645 (N_1645,N_1420,N_1492);
or U1646 (N_1646,N_1492,N_1485);
or U1647 (N_1647,N_1353,N_1399);
nand U1648 (N_1648,N_1470,N_1353);
nand U1649 (N_1649,N_1387,N_1494);
and U1650 (N_1650,N_1506,N_1580);
nand U1651 (N_1651,N_1573,N_1579);
or U1652 (N_1652,N_1643,N_1637);
or U1653 (N_1653,N_1563,N_1531);
and U1654 (N_1654,N_1575,N_1620);
or U1655 (N_1655,N_1644,N_1560);
xor U1656 (N_1656,N_1610,N_1537);
or U1657 (N_1657,N_1603,N_1594);
nor U1658 (N_1658,N_1562,N_1585);
nor U1659 (N_1659,N_1642,N_1626);
nor U1660 (N_1660,N_1527,N_1534);
or U1661 (N_1661,N_1606,N_1515);
xor U1662 (N_1662,N_1523,N_1646);
xor U1663 (N_1663,N_1533,N_1535);
or U1664 (N_1664,N_1616,N_1553);
nand U1665 (N_1665,N_1538,N_1524);
nand U1666 (N_1666,N_1526,N_1541);
nand U1667 (N_1667,N_1544,N_1501);
or U1668 (N_1668,N_1631,N_1597);
nor U1669 (N_1669,N_1512,N_1624);
and U1670 (N_1670,N_1511,N_1532);
and U1671 (N_1671,N_1525,N_1557);
xnor U1672 (N_1672,N_1561,N_1551);
xnor U1673 (N_1673,N_1582,N_1618);
nand U1674 (N_1674,N_1507,N_1649);
nand U1675 (N_1675,N_1564,N_1529);
nand U1676 (N_1676,N_1550,N_1530);
xor U1677 (N_1677,N_1503,N_1513);
xor U1678 (N_1678,N_1641,N_1542);
and U1679 (N_1679,N_1548,N_1565);
nor U1680 (N_1680,N_1614,N_1622);
xnor U1681 (N_1681,N_1632,N_1590);
nor U1682 (N_1682,N_1546,N_1543);
xor U1683 (N_1683,N_1566,N_1587);
and U1684 (N_1684,N_1558,N_1568);
and U1685 (N_1685,N_1628,N_1522);
nand U1686 (N_1686,N_1648,N_1520);
or U1687 (N_1687,N_1549,N_1619);
xor U1688 (N_1688,N_1581,N_1601);
or U1689 (N_1689,N_1630,N_1502);
xor U1690 (N_1690,N_1623,N_1504);
or U1691 (N_1691,N_1647,N_1540);
xnor U1692 (N_1692,N_1559,N_1574);
or U1693 (N_1693,N_1547,N_1600);
or U1694 (N_1694,N_1640,N_1612);
xor U1695 (N_1695,N_1584,N_1500);
and U1696 (N_1696,N_1617,N_1621);
xnor U1697 (N_1697,N_1536,N_1636);
or U1698 (N_1698,N_1576,N_1517);
nor U1699 (N_1699,N_1510,N_1608);
and U1700 (N_1700,N_1629,N_1552);
and U1701 (N_1701,N_1516,N_1583);
nand U1702 (N_1702,N_1607,N_1602);
and U1703 (N_1703,N_1609,N_1596);
nor U1704 (N_1704,N_1613,N_1625);
nand U1705 (N_1705,N_1505,N_1635);
xnor U1706 (N_1706,N_1591,N_1539);
and U1707 (N_1707,N_1554,N_1598);
nor U1708 (N_1708,N_1627,N_1599);
and U1709 (N_1709,N_1509,N_1528);
nor U1710 (N_1710,N_1615,N_1508);
or U1711 (N_1711,N_1555,N_1556);
and U1712 (N_1712,N_1589,N_1595);
nor U1713 (N_1713,N_1593,N_1633);
and U1714 (N_1714,N_1514,N_1571);
and U1715 (N_1715,N_1570,N_1572);
or U1716 (N_1716,N_1545,N_1592);
xnor U1717 (N_1717,N_1611,N_1567);
or U1718 (N_1718,N_1588,N_1518);
and U1719 (N_1719,N_1604,N_1521);
and U1720 (N_1720,N_1605,N_1578);
nor U1721 (N_1721,N_1634,N_1639);
or U1722 (N_1722,N_1519,N_1577);
xor U1723 (N_1723,N_1645,N_1638);
nand U1724 (N_1724,N_1586,N_1569);
xor U1725 (N_1725,N_1538,N_1594);
and U1726 (N_1726,N_1639,N_1500);
and U1727 (N_1727,N_1612,N_1581);
xor U1728 (N_1728,N_1632,N_1508);
xnor U1729 (N_1729,N_1558,N_1562);
xor U1730 (N_1730,N_1574,N_1530);
xor U1731 (N_1731,N_1647,N_1500);
or U1732 (N_1732,N_1631,N_1635);
nand U1733 (N_1733,N_1504,N_1634);
nand U1734 (N_1734,N_1623,N_1577);
xor U1735 (N_1735,N_1520,N_1569);
xnor U1736 (N_1736,N_1541,N_1610);
nand U1737 (N_1737,N_1634,N_1573);
and U1738 (N_1738,N_1514,N_1638);
and U1739 (N_1739,N_1552,N_1573);
and U1740 (N_1740,N_1629,N_1509);
nor U1741 (N_1741,N_1587,N_1549);
nand U1742 (N_1742,N_1604,N_1515);
and U1743 (N_1743,N_1532,N_1614);
xor U1744 (N_1744,N_1613,N_1573);
nand U1745 (N_1745,N_1607,N_1644);
nor U1746 (N_1746,N_1596,N_1523);
xor U1747 (N_1747,N_1556,N_1586);
xor U1748 (N_1748,N_1585,N_1638);
and U1749 (N_1749,N_1631,N_1528);
xnor U1750 (N_1750,N_1627,N_1562);
nor U1751 (N_1751,N_1541,N_1558);
or U1752 (N_1752,N_1604,N_1631);
or U1753 (N_1753,N_1606,N_1545);
nor U1754 (N_1754,N_1602,N_1638);
nor U1755 (N_1755,N_1510,N_1648);
and U1756 (N_1756,N_1595,N_1636);
or U1757 (N_1757,N_1635,N_1521);
nand U1758 (N_1758,N_1566,N_1536);
or U1759 (N_1759,N_1597,N_1545);
or U1760 (N_1760,N_1571,N_1616);
nor U1761 (N_1761,N_1618,N_1638);
nand U1762 (N_1762,N_1571,N_1538);
nand U1763 (N_1763,N_1544,N_1602);
or U1764 (N_1764,N_1512,N_1501);
or U1765 (N_1765,N_1578,N_1586);
nand U1766 (N_1766,N_1508,N_1578);
nor U1767 (N_1767,N_1560,N_1592);
nand U1768 (N_1768,N_1632,N_1521);
xor U1769 (N_1769,N_1602,N_1636);
nand U1770 (N_1770,N_1534,N_1615);
nand U1771 (N_1771,N_1631,N_1508);
and U1772 (N_1772,N_1532,N_1580);
or U1773 (N_1773,N_1549,N_1561);
xnor U1774 (N_1774,N_1575,N_1587);
and U1775 (N_1775,N_1503,N_1529);
and U1776 (N_1776,N_1562,N_1534);
xnor U1777 (N_1777,N_1617,N_1563);
nor U1778 (N_1778,N_1625,N_1641);
xnor U1779 (N_1779,N_1627,N_1515);
and U1780 (N_1780,N_1554,N_1587);
nand U1781 (N_1781,N_1607,N_1516);
and U1782 (N_1782,N_1599,N_1558);
xor U1783 (N_1783,N_1502,N_1520);
xor U1784 (N_1784,N_1600,N_1532);
xor U1785 (N_1785,N_1577,N_1544);
xnor U1786 (N_1786,N_1585,N_1625);
or U1787 (N_1787,N_1555,N_1566);
and U1788 (N_1788,N_1559,N_1565);
nor U1789 (N_1789,N_1515,N_1529);
xor U1790 (N_1790,N_1561,N_1613);
nor U1791 (N_1791,N_1605,N_1632);
nand U1792 (N_1792,N_1567,N_1510);
nand U1793 (N_1793,N_1524,N_1601);
or U1794 (N_1794,N_1537,N_1534);
xnor U1795 (N_1795,N_1619,N_1502);
nor U1796 (N_1796,N_1547,N_1593);
or U1797 (N_1797,N_1641,N_1620);
nand U1798 (N_1798,N_1594,N_1576);
or U1799 (N_1799,N_1575,N_1615);
or U1800 (N_1800,N_1685,N_1764);
xor U1801 (N_1801,N_1682,N_1720);
or U1802 (N_1802,N_1748,N_1694);
nor U1803 (N_1803,N_1690,N_1683);
and U1804 (N_1804,N_1740,N_1776);
and U1805 (N_1805,N_1793,N_1708);
nand U1806 (N_1806,N_1657,N_1772);
or U1807 (N_1807,N_1782,N_1735);
nand U1808 (N_1808,N_1754,N_1786);
xor U1809 (N_1809,N_1670,N_1766);
and U1810 (N_1810,N_1680,N_1741);
or U1811 (N_1811,N_1790,N_1781);
or U1812 (N_1812,N_1799,N_1695);
xor U1813 (N_1813,N_1699,N_1662);
nand U1814 (N_1814,N_1664,N_1678);
nand U1815 (N_1815,N_1715,N_1779);
nor U1816 (N_1816,N_1794,N_1763);
or U1817 (N_1817,N_1796,N_1673);
nand U1818 (N_1818,N_1739,N_1744);
and U1819 (N_1819,N_1788,N_1711);
nor U1820 (N_1820,N_1671,N_1791);
nor U1821 (N_1821,N_1755,N_1674);
xor U1822 (N_1822,N_1768,N_1784);
nor U1823 (N_1823,N_1652,N_1752);
and U1824 (N_1824,N_1718,N_1713);
and U1825 (N_1825,N_1717,N_1653);
and U1826 (N_1826,N_1660,N_1730);
or U1827 (N_1827,N_1751,N_1736);
nand U1828 (N_1828,N_1734,N_1709);
xor U1829 (N_1829,N_1780,N_1700);
nand U1830 (N_1830,N_1756,N_1667);
nand U1831 (N_1831,N_1691,N_1759);
nor U1832 (N_1832,N_1797,N_1686);
or U1833 (N_1833,N_1760,N_1672);
xnor U1834 (N_1834,N_1723,N_1714);
xor U1835 (N_1835,N_1746,N_1687);
xnor U1836 (N_1836,N_1765,N_1719);
nor U1837 (N_1837,N_1656,N_1777);
nor U1838 (N_1838,N_1750,N_1679);
or U1839 (N_1839,N_1761,N_1704);
or U1840 (N_1840,N_1659,N_1721);
and U1841 (N_1841,N_1669,N_1731);
xor U1842 (N_1842,N_1698,N_1753);
and U1843 (N_1843,N_1775,N_1676);
nor U1844 (N_1844,N_1798,N_1666);
nor U1845 (N_1845,N_1702,N_1749);
and U1846 (N_1846,N_1738,N_1722);
nand U1847 (N_1847,N_1688,N_1651);
and U1848 (N_1848,N_1758,N_1701);
and U1849 (N_1849,N_1726,N_1650);
and U1850 (N_1850,N_1743,N_1706);
nand U1851 (N_1851,N_1693,N_1703);
xor U1852 (N_1852,N_1684,N_1737);
nand U1853 (N_1853,N_1774,N_1771);
and U1854 (N_1854,N_1729,N_1795);
xor U1855 (N_1855,N_1747,N_1707);
nand U1856 (N_1856,N_1785,N_1725);
and U1857 (N_1857,N_1792,N_1783);
nor U1858 (N_1858,N_1665,N_1769);
and U1859 (N_1859,N_1767,N_1727);
nor U1860 (N_1860,N_1677,N_1675);
nor U1861 (N_1861,N_1668,N_1654);
nand U1862 (N_1862,N_1689,N_1770);
nor U1863 (N_1863,N_1732,N_1663);
and U1864 (N_1864,N_1692,N_1745);
and U1865 (N_1865,N_1697,N_1716);
nand U1866 (N_1866,N_1757,N_1705);
nand U1867 (N_1867,N_1661,N_1787);
nand U1868 (N_1868,N_1724,N_1655);
nor U1869 (N_1869,N_1710,N_1733);
nor U1870 (N_1870,N_1658,N_1696);
and U1871 (N_1871,N_1789,N_1681);
or U1872 (N_1872,N_1773,N_1778);
xnor U1873 (N_1873,N_1762,N_1728);
xnor U1874 (N_1874,N_1712,N_1742);
or U1875 (N_1875,N_1786,N_1672);
or U1876 (N_1876,N_1739,N_1750);
nor U1877 (N_1877,N_1764,N_1669);
xor U1878 (N_1878,N_1731,N_1682);
xnor U1879 (N_1879,N_1695,N_1775);
nor U1880 (N_1880,N_1664,N_1778);
nand U1881 (N_1881,N_1700,N_1687);
or U1882 (N_1882,N_1687,N_1711);
and U1883 (N_1883,N_1792,N_1756);
and U1884 (N_1884,N_1721,N_1779);
nand U1885 (N_1885,N_1661,N_1778);
xor U1886 (N_1886,N_1650,N_1677);
xnor U1887 (N_1887,N_1686,N_1683);
or U1888 (N_1888,N_1674,N_1733);
nor U1889 (N_1889,N_1793,N_1771);
and U1890 (N_1890,N_1662,N_1786);
nand U1891 (N_1891,N_1736,N_1673);
or U1892 (N_1892,N_1672,N_1716);
or U1893 (N_1893,N_1796,N_1765);
nor U1894 (N_1894,N_1735,N_1744);
xor U1895 (N_1895,N_1660,N_1755);
nor U1896 (N_1896,N_1698,N_1694);
or U1897 (N_1897,N_1722,N_1791);
nand U1898 (N_1898,N_1758,N_1680);
nor U1899 (N_1899,N_1784,N_1755);
and U1900 (N_1900,N_1652,N_1688);
nor U1901 (N_1901,N_1683,N_1710);
nor U1902 (N_1902,N_1702,N_1665);
nand U1903 (N_1903,N_1772,N_1693);
and U1904 (N_1904,N_1760,N_1694);
and U1905 (N_1905,N_1685,N_1763);
nand U1906 (N_1906,N_1799,N_1762);
and U1907 (N_1907,N_1782,N_1653);
or U1908 (N_1908,N_1767,N_1794);
or U1909 (N_1909,N_1687,N_1690);
or U1910 (N_1910,N_1673,N_1658);
xor U1911 (N_1911,N_1692,N_1739);
nand U1912 (N_1912,N_1749,N_1676);
and U1913 (N_1913,N_1736,N_1786);
xor U1914 (N_1914,N_1656,N_1715);
and U1915 (N_1915,N_1798,N_1706);
xor U1916 (N_1916,N_1709,N_1794);
xnor U1917 (N_1917,N_1679,N_1747);
nand U1918 (N_1918,N_1683,N_1793);
xnor U1919 (N_1919,N_1672,N_1677);
nor U1920 (N_1920,N_1657,N_1698);
and U1921 (N_1921,N_1671,N_1677);
nand U1922 (N_1922,N_1755,N_1718);
nand U1923 (N_1923,N_1759,N_1689);
nand U1924 (N_1924,N_1673,N_1680);
xor U1925 (N_1925,N_1679,N_1761);
nand U1926 (N_1926,N_1724,N_1728);
and U1927 (N_1927,N_1687,N_1748);
xnor U1928 (N_1928,N_1702,N_1662);
nor U1929 (N_1929,N_1659,N_1652);
and U1930 (N_1930,N_1658,N_1747);
nor U1931 (N_1931,N_1761,N_1720);
nand U1932 (N_1932,N_1721,N_1766);
and U1933 (N_1933,N_1781,N_1658);
nor U1934 (N_1934,N_1742,N_1704);
nand U1935 (N_1935,N_1771,N_1789);
nand U1936 (N_1936,N_1799,N_1664);
or U1937 (N_1937,N_1745,N_1798);
nor U1938 (N_1938,N_1777,N_1760);
xor U1939 (N_1939,N_1677,N_1685);
nor U1940 (N_1940,N_1673,N_1671);
nand U1941 (N_1941,N_1655,N_1652);
nand U1942 (N_1942,N_1799,N_1739);
nor U1943 (N_1943,N_1680,N_1743);
or U1944 (N_1944,N_1656,N_1766);
xor U1945 (N_1945,N_1666,N_1653);
and U1946 (N_1946,N_1666,N_1791);
or U1947 (N_1947,N_1701,N_1770);
nor U1948 (N_1948,N_1657,N_1712);
and U1949 (N_1949,N_1675,N_1663);
and U1950 (N_1950,N_1841,N_1892);
or U1951 (N_1951,N_1847,N_1881);
nand U1952 (N_1952,N_1896,N_1816);
nand U1953 (N_1953,N_1909,N_1932);
or U1954 (N_1954,N_1890,N_1948);
nor U1955 (N_1955,N_1928,N_1913);
nor U1956 (N_1956,N_1897,N_1858);
and U1957 (N_1957,N_1856,N_1840);
xor U1958 (N_1958,N_1862,N_1832);
nor U1959 (N_1959,N_1888,N_1905);
nand U1960 (N_1960,N_1808,N_1926);
nand U1961 (N_1961,N_1949,N_1884);
and U1962 (N_1962,N_1901,N_1865);
nor U1963 (N_1963,N_1921,N_1895);
and U1964 (N_1964,N_1887,N_1923);
nor U1965 (N_1965,N_1920,N_1813);
nand U1966 (N_1966,N_1947,N_1937);
or U1967 (N_1967,N_1803,N_1922);
and U1968 (N_1968,N_1942,N_1906);
xnor U1969 (N_1969,N_1836,N_1869);
nand U1970 (N_1970,N_1938,N_1883);
and U1971 (N_1971,N_1860,N_1844);
nand U1972 (N_1972,N_1886,N_1830);
nand U1973 (N_1973,N_1857,N_1822);
nor U1974 (N_1974,N_1910,N_1839);
and U1975 (N_1975,N_1902,N_1874);
xnor U1976 (N_1976,N_1826,N_1848);
nand U1977 (N_1977,N_1835,N_1815);
and U1978 (N_1978,N_1801,N_1919);
xor U1979 (N_1979,N_1802,N_1871);
and U1980 (N_1980,N_1870,N_1939);
and U1981 (N_1981,N_1931,N_1846);
nand U1982 (N_1982,N_1821,N_1804);
nand U1983 (N_1983,N_1861,N_1929);
nor U1984 (N_1984,N_1899,N_1805);
nand U1985 (N_1985,N_1807,N_1936);
and U1986 (N_1986,N_1907,N_1838);
nor U1987 (N_1987,N_1849,N_1814);
nor U1988 (N_1988,N_1818,N_1908);
xor U1989 (N_1989,N_1806,N_1934);
nand U1990 (N_1990,N_1851,N_1893);
nand U1991 (N_1991,N_1875,N_1876);
and U1992 (N_1992,N_1943,N_1903);
xnor U1993 (N_1993,N_1915,N_1940);
nor U1994 (N_1994,N_1900,N_1850);
nor U1995 (N_1995,N_1837,N_1911);
nor U1996 (N_1996,N_1852,N_1800);
and U1997 (N_1997,N_1864,N_1918);
nand U1998 (N_1998,N_1872,N_1941);
xor U1999 (N_1999,N_1817,N_1853);
nor U2000 (N_2000,N_1944,N_1879);
xnor U2001 (N_2001,N_1946,N_1882);
and U2002 (N_2002,N_1825,N_1820);
nand U2003 (N_2003,N_1885,N_1891);
or U2004 (N_2004,N_1824,N_1819);
and U2005 (N_2005,N_1845,N_1878);
nor U2006 (N_2006,N_1810,N_1866);
and U2007 (N_2007,N_1912,N_1868);
or U2008 (N_2008,N_1809,N_1925);
and U2009 (N_2009,N_1842,N_1855);
nand U2010 (N_2010,N_1914,N_1927);
nand U2011 (N_2011,N_1889,N_1823);
nor U2012 (N_2012,N_1877,N_1843);
nor U2013 (N_2013,N_1828,N_1859);
nor U2014 (N_2014,N_1863,N_1873);
and U2015 (N_2015,N_1827,N_1811);
or U2016 (N_2016,N_1930,N_1917);
and U2017 (N_2017,N_1834,N_1829);
nor U2018 (N_2018,N_1833,N_1894);
nand U2019 (N_2019,N_1924,N_1812);
xor U2020 (N_2020,N_1831,N_1935);
nand U2021 (N_2021,N_1945,N_1933);
xnor U2022 (N_2022,N_1867,N_1904);
xnor U2023 (N_2023,N_1898,N_1880);
or U2024 (N_2024,N_1854,N_1916);
xnor U2025 (N_2025,N_1930,N_1923);
and U2026 (N_2026,N_1869,N_1841);
xor U2027 (N_2027,N_1890,N_1856);
nor U2028 (N_2028,N_1806,N_1895);
or U2029 (N_2029,N_1939,N_1844);
xnor U2030 (N_2030,N_1833,N_1934);
nand U2031 (N_2031,N_1885,N_1876);
and U2032 (N_2032,N_1940,N_1931);
nand U2033 (N_2033,N_1875,N_1898);
and U2034 (N_2034,N_1836,N_1880);
nand U2035 (N_2035,N_1822,N_1890);
or U2036 (N_2036,N_1899,N_1852);
nor U2037 (N_2037,N_1844,N_1857);
nor U2038 (N_2038,N_1814,N_1830);
nand U2039 (N_2039,N_1933,N_1859);
nand U2040 (N_2040,N_1941,N_1806);
xnor U2041 (N_2041,N_1909,N_1895);
nand U2042 (N_2042,N_1873,N_1881);
and U2043 (N_2043,N_1899,N_1825);
xor U2044 (N_2044,N_1946,N_1943);
xnor U2045 (N_2045,N_1929,N_1903);
nand U2046 (N_2046,N_1912,N_1861);
and U2047 (N_2047,N_1816,N_1815);
xnor U2048 (N_2048,N_1878,N_1902);
nor U2049 (N_2049,N_1939,N_1823);
or U2050 (N_2050,N_1946,N_1902);
nand U2051 (N_2051,N_1835,N_1859);
or U2052 (N_2052,N_1916,N_1891);
xor U2053 (N_2053,N_1927,N_1898);
nand U2054 (N_2054,N_1924,N_1860);
nand U2055 (N_2055,N_1938,N_1934);
nor U2056 (N_2056,N_1863,N_1827);
nand U2057 (N_2057,N_1916,N_1931);
xor U2058 (N_2058,N_1867,N_1885);
nor U2059 (N_2059,N_1865,N_1949);
xor U2060 (N_2060,N_1924,N_1929);
and U2061 (N_2061,N_1923,N_1825);
and U2062 (N_2062,N_1923,N_1890);
and U2063 (N_2063,N_1858,N_1861);
or U2064 (N_2064,N_1877,N_1824);
and U2065 (N_2065,N_1915,N_1853);
xnor U2066 (N_2066,N_1895,N_1941);
or U2067 (N_2067,N_1892,N_1925);
and U2068 (N_2068,N_1812,N_1877);
and U2069 (N_2069,N_1854,N_1839);
nand U2070 (N_2070,N_1895,N_1866);
and U2071 (N_2071,N_1863,N_1896);
or U2072 (N_2072,N_1918,N_1884);
xor U2073 (N_2073,N_1858,N_1938);
or U2074 (N_2074,N_1925,N_1939);
nand U2075 (N_2075,N_1813,N_1816);
or U2076 (N_2076,N_1859,N_1838);
or U2077 (N_2077,N_1841,N_1876);
nand U2078 (N_2078,N_1891,N_1871);
nor U2079 (N_2079,N_1922,N_1907);
and U2080 (N_2080,N_1881,N_1836);
or U2081 (N_2081,N_1810,N_1898);
nand U2082 (N_2082,N_1898,N_1832);
or U2083 (N_2083,N_1895,N_1914);
and U2084 (N_2084,N_1924,N_1803);
xor U2085 (N_2085,N_1897,N_1940);
nand U2086 (N_2086,N_1808,N_1866);
or U2087 (N_2087,N_1938,N_1813);
nor U2088 (N_2088,N_1933,N_1848);
or U2089 (N_2089,N_1887,N_1864);
or U2090 (N_2090,N_1897,N_1947);
nor U2091 (N_2091,N_1920,N_1847);
or U2092 (N_2092,N_1880,N_1812);
and U2093 (N_2093,N_1935,N_1934);
nand U2094 (N_2094,N_1814,N_1913);
nand U2095 (N_2095,N_1836,N_1902);
and U2096 (N_2096,N_1890,N_1928);
and U2097 (N_2097,N_1850,N_1918);
xnor U2098 (N_2098,N_1875,N_1851);
and U2099 (N_2099,N_1943,N_1818);
nand U2100 (N_2100,N_2095,N_1951);
and U2101 (N_2101,N_2094,N_2078);
nand U2102 (N_2102,N_2085,N_2071);
xor U2103 (N_2103,N_2021,N_2017);
or U2104 (N_2104,N_1974,N_2042);
and U2105 (N_2105,N_2072,N_2059);
or U2106 (N_2106,N_2055,N_2057);
xnor U2107 (N_2107,N_2052,N_1968);
xnor U2108 (N_2108,N_2050,N_2013);
nand U2109 (N_2109,N_2043,N_2046);
nand U2110 (N_2110,N_2090,N_1966);
nor U2111 (N_2111,N_2022,N_2033);
nor U2112 (N_2112,N_2012,N_2025);
xor U2113 (N_2113,N_2028,N_2038);
xnor U2114 (N_2114,N_1989,N_2091);
xor U2115 (N_2115,N_2014,N_2084);
and U2116 (N_2116,N_1986,N_1998);
and U2117 (N_2117,N_1967,N_2099);
nand U2118 (N_2118,N_2073,N_1961);
and U2119 (N_2119,N_2077,N_2067);
and U2120 (N_2120,N_2079,N_1956);
and U2121 (N_2121,N_2004,N_2096);
nand U2122 (N_2122,N_2026,N_1976);
nor U2123 (N_2123,N_2058,N_1955);
nand U2124 (N_2124,N_1973,N_2069);
or U2125 (N_2125,N_1965,N_1971);
nand U2126 (N_2126,N_1991,N_2063);
nor U2127 (N_2127,N_1979,N_2092);
nor U2128 (N_2128,N_2054,N_2035);
or U2129 (N_2129,N_2068,N_2056);
or U2130 (N_2130,N_2074,N_2034);
nand U2131 (N_2131,N_2001,N_2005);
or U2132 (N_2132,N_1950,N_1984);
or U2133 (N_2133,N_2062,N_1982);
and U2134 (N_2134,N_2082,N_2008);
and U2135 (N_2135,N_1972,N_2076);
nand U2136 (N_2136,N_1977,N_1953);
nand U2137 (N_2137,N_1999,N_2019);
or U2138 (N_2138,N_2051,N_2053);
xor U2139 (N_2139,N_1992,N_2002);
and U2140 (N_2140,N_2087,N_2049);
xnor U2141 (N_2141,N_2009,N_2086);
and U2142 (N_2142,N_2083,N_1958);
and U2143 (N_2143,N_2036,N_1970);
and U2144 (N_2144,N_2020,N_1980);
nand U2145 (N_2145,N_1987,N_2070);
and U2146 (N_2146,N_1985,N_2015);
or U2147 (N_2147,N_2029,N_1990);
xor U2148 (N_2148,N_2064,N_1996);
and U2149 (N_2149,N_2060,N_2024);
xnor U2150 (N_2150,N_2027,N_2081);
nand U2151 (N_2151,N_2047,N_1952);
or U2152 (N_2152,N_2000,N_2093);
or U2153 (N_2153,N_1983,N_1997);
and U2154 (N_2154,N_2044,N_2031);
nor U2155 (N_2155,N_1988,N_2011);
or U2156 (N_2156,N_1981,N_2080);
nor U2157 (N_2157,N_2097,N_1978);
xnor U2158 (N_2158,N_2041,N_2066);
or U2159 (N_2159,N_2065,N_1975);
and U2160 (N_2160,N_1969,N_2010);
and U2161 (N_2161,N_2018,N_1954);
or U2162 (N_2162,N_1960,N_1962);
and U2163 (N_2163,N_2003,N_1993);
xnor U2164 (N_2164,N_2089,N_1994);
and U2165 (N_2165,N_2037,N_2023);
or U2166 (N_2166,N_2039,N_2016);
and U2167 (N_2167,N_2032,N_2040);
nor U2168 (N_2168,N_1995,N_2007);
xnor U2169 (N_2169,N_2098,N_2048);
nand U2170 (N_2170,N_2030,N_2088);
or U2171 (N_2171,N_2045,N_1957);
nor U2172 (N_2172,N_2061,N_1959);
or U2173 (N_2173,N_2075,N_2006);
nor U2174 (N_2174,N_1964,N_1963);
and U2175 (N_2175,N_2005,N_2064);
or U2176 (N_2176,N_2073,N_2061);
or U2177 (N_2177,N_2058,N_2097);
nor U2178 (N_2178,N_2085,N_1987);
xnor U2179 (N_2179,N_2071,N_1995);
and U2180 (N_2180,N_2065,N_2063);
or U2181 (N_2181,N_1950,N_2039);
nor U2182 (N_2182,N_2045,N_1954);
nand U2183 (N_2183,N_2021,N_2048);
and U2184 (N_2184,N_2009,N_1959);
xor U2185 (N_2185,N_2041,N_2083);
nor U2186 (N_2186,N_2089,N_2058);
and U2187 (N_2187,N_2072,N_2056);
nor U2188 (N_2188,N_2036,N_2005);
or U2189 (N_2189,N_2007,N_2068);
or U2190 (N_2190,N_1955,N_1983);
nor U2191 (N_2191,N_2041,N_2072);
and U2192 (N_2192,N_2005,N_1984);
and U2193 (N_2193,N_1950,N_2088);
or U2194 (N_2194,N_2013,N_2034);
nor U2195 (N_2195,N_2042,N_1998);
and U2196 (N_2196,N_2079,N_2025);
and U2197 (N_2197,N_2026,N_2086);
or U2198 (N_2198,N_2079,N_2072);
and U2199 (N_2199,N_2088,N_2081);
nor U2200 (N_2200,N_1981,N_1957);
and U2201 (N_2201,N_1954,N_2047);
nand U2202 (N_2202,N_2096,N_1990);
xor U2203 (N_2203,N_2026,N_2055);
and U2204 (N_2204,N_1996,N_1965);
xor U2205 (N_2205,N_1968,N_2050);
nand U2206 (N_2206,N_2041,N_2010);
nor U2207 (N_2207,N_2049,N_2071);
xor U2208 (N_2208,N_1962,N_2045);
nand U2209 (N_2209,N_2046,N_2007);
xor U2210 (N_2210,N_2046,N_2036);
xor U2211 (N_2211,N_1966,N_2021);
or U2212 (N_2212,N_1982,N_1997);
and U2213 (N_2213,N_2065,N_1960);
nor U2214 (N_2214,N_2022,N_2084);
or U2215 (N_2215,N_2089,N_2095);
or U2216 (N_2216,N_2020,N_2090);
or U2217 (N_2217,N_2036,N_2098);
nand U2218 (N_2218,N_2059,N_1956);
xnor U2219 (N_2219,N_2010,N_2019);
nor U2220 (N_2220,N_2000,N_1989);
xnor U2221 (N_2221,N_2061,N_2097);
nand U2222 (N_2222,N_2034,N_1992);
xor U2223 (N_2223,N_2068,N_2041);
nor U2224 (N_2224,N_2036,N_2050);
nand U2225 (N_2225,N_2054,N_2031);
xnor U2226 (N_2226,N_1970,N_2063);
xnor U2227 (N_2227,N_2014,N_1952);
xor U2228 (N_2228,N_1993,N_2097);
xor U2229 (N_2229,N_1969,N_1983);
nor U2230 (N_2230,N_2087,N_2043);
or U2231 (N_2231,N_1967,N_1960);
or U2232 (N_2232,N_2090,N_2023);
and U2233 (N_2233,N_2047,N_1993);
nor U2234 (N_2234,N_2097,N_1998);
xnor U2235 (N_2235,N_2046,N_2011);
and U2236 (N_2236,N_2013,N_1955);
and U2237 (N_2237,N_2068,N_1960);
and U2238 (N_2238,N_2017,N_2076);
or U2239 (N_2239,N_1978,N_1953);
and U2240 (N_2240,N_2089,N_2068);
nor U2241 (N_2241,N_2073,N_2086);
xnor U2242 (N_2242,N_2070,N_2093);
xnor U2243 (N_2243,N_1976,N_1974);
or U2244 (N_2244,N_2019,N_1970);
nor U2245 (N_2245,N_1988,N_1979);
nand U2246 (N_2246,N_2021,N_1975);
or U2247 (N_2247,N_2005,N_2013);
nand U2248 (N_2248,N_2034,N_2033);
and U2249 (N_2249,N_2077,N_1993);
or U2250 (N_2250,N_2156,N_2177);
xnor U2251 (N_2251,N_2172,N_2248);
or U2252 (N_2252,N_2249,N_2158);
nor U2253 (N_2253,N_2194,N_2100);
or U2254 (N_2254,N_2227,N_2154);
and U2255 (N_2255,N_2126,N_2245);
nand U2256 (N_2256,N_2131,N_2180);
nand U2257 (N_2257,N_2215,N_2109);
nor U2258 (N_2258,N_2107,N_2173);
nand U2259 (N_2259,N_2179,N_2188);
nor U2260 (N_2260,N_2239,N_2151);
nand U2261 (N_2261,N_2136,N_2103);
and U2262 (N_2262,N_2138,N_2175);
nand U2263 (N_2263,N_2114,N_2149);
nor U2264 (N_2264,N_2160,N_2208);
nor U2265 (N_2265,N_2152,N_2241);
or U2266 (N_2266,N_2236,N_2168);
or U2267 (N_2267,N_2247,N_2157);
xnor U2268 (N_2268,N_2231,N_2133);
nor U2269 (N_2269,N_2161,N_2176);
nand U2270 (N_2270,N_2198,N_2190);
or U2271 (N_2271,N_2106,N_2203);
nor U2272 (N_2272,N_2134,N_2132);
xnor U2273 (N_2273,N_2225,N_2178);
nor U2274 (N_2274,N_2145,N_2214);
nor U2275 (N_2275,N_2135,N_2235);
and U2276 (N_2276,N_2234,N_2219);
nand U2277 (N_2277,N_2102,N_2246);
nand U2278 (N_2278,N_2229,N_2116);
xor U2279 (N_2279,N_2101,N_2207);
nand U2280 (N_2280,N_2221,N_2123);
or U2281 (N_2281,N_2184,N_2205);
or U2282 (N_2282,N_2144,N_2113);
nor U2283 (N_2283,N_2223,N_2125);
xor U2284 (N_2284,N_2118,N_2202);
nor U2285 (N_2285,N_2159,N_2108);
and U2286 (N_2286,N_2186,N_2199);
and U2287 (N_2287,N_2197,N_2164);
xor U2288 (N_2288,N_2212,N_2139);
and U2289 (N_2289,N_2233,N_2121);
and U2290 (N_2290,N_2153,N_2204);
and U2291 (N_2291,N_2182,N_2147);
or U2292 (N_2292,N_2104,N_2142);
nor U2293 (N_2293,N_2240,N_2238);
xor U2294 (N_2294,N_2185,N_2243);
xor U2295 (N_2295,N_2146,N_2213);
and U2296 (N_2296,N_2115,N_2226);
nand U2297 (N_2297,N_2209,N_2148);
nor U2298 (N_2298,N_2230,N_2206);
and U2299 (N_2299,N_2187,N_2143);
xor U2300 (N_2300,N_2150,N_2242);
or U2301 (N_2301,N_2192,N_2232);
and U2302 (N_2302,N_2110,N_2211);
nand U2303 (N_2303,N_2218,N_2137);
and U2304 (N_2304,N_2155,N_2162);
and U2305 (N_2305,N_2127,N_2111);
nor U2306 (N_2306,N_2228,N_2112);
and U2307 (N_2307,N_2196,N_2122);
nand U2308 (N_2308,N_2128,N_2124);
nand U2309 (N_2309,N_2189,N_2220);
nand U2310 (N_2310,N_2166,N_2191);
nand U2311 (N_2311,N_2167,N_2237);
nand U2312 (N_2312,N_2244,N_2120);
or U2313 (N_2313,N_2174,N_2117);
nand U2314 (N_2314,N_2171,N_2224);
and U2315 (N_2315,N_2183,N_2181);
nand U2316 (N_2316,N_2195,N_2222);
and U2317 (N_2317,N_2163,N_2210);
xnor U2318 (N_2318,N_2140,N_2201);
nand U2319 (N_2319,N_2129,N_2130);
nor U2320 (N_2320,N_2193,N_2170);
xor U2321 (N_2321,N_2165,N_2216);
xnor U2322 (N_2322,N_2200,N_2217);
or U2323 (N_2323,N_2169,N_2119);
nor U2324 (N_2324,N_2105,N_2141);
nand U2325 (N_2325,N_2234,N_2247);
or U2326 (N_2326,N_2128,N_2142);
xor U2327 (N_2327,N_2212,N_2132);
or U2328 (N_2328,N_2137,N_2109);
and U2329 (N_2329,N_2138,N_2198);
nor U2330 (N_2330,N_2214,N_2248);
xnor U2331 (N_2331,N_2193,N_2160);
xor U2332 (N_2332,N_2106,N_2229);
xnor U2333 (N_2333,N_2127,N_2187);
xnor U2334 (N_2334,N_2153,N_2149);
nor U2335 (N_2335,N_2136,N_2198);
and U2336 (N_2336,N_2173,N_2233);
and U2337 (N_2337,N_2226,N_2119);
and U2338 (N_2338,N_2167,N_2150);
nand U2339 (N_2339,N_2103,N_2145);
nor U2340 (N_2340,N_2119,N_2104);
or U2341 (N_2341,N_2147,N_2112);
or U2342 (N_2342,N_2111,N_2126);
nand U2343 (N_2343,N_2226,N_2178);
and U2344 (N_2344,N_2116,N_2140);
or U2345 (N_2345,N_2146,N_2127);
nand U2346 (N_2346,N_2125,N_2175);
nand U2347 (N_2347,N_2218,N_2105);
xor U2348 (N_2348,N_2114,N_2226);
and U2349 (N_2349,N_2123,N_2237);
nand U2350 (N_2350,N_2220,N_2151);
xor U2351 (N_2351,N_2179,N_2218);
xnor U2352 (N_2352,N_2150,N_2212);
and U2353 (N_2353,N_2118,N_2107);
nor U2354 (N_2354,N_2169,N_2129);
nand U2355 (N_2355,N_2193,N_2214);
or U2356 (N_2356,N_2209,N_2161);
nor U2357 (N_2357,N_2170,N_2165);
and U2358 (N_2358,N_2168,N_2209);
or U2359 (N_2359,N_2198,N_2152);
and U2360 (N_2360,N_2196,N_2182);
nand U2361 (N_2361,N_2206,N_2238);
xor U2362 (N_2362,N_2107,N_2232);
xor U2363 (N_2363,N_2128,N_2159);
nor U2364 (N_2364,N_2230,N_2102);
nand U2365 (N_2365,N_2100,N_2206);
and U2366 (N_2366,N_2146,N_2106);
xor U2367 (N_2367,N_2190,N_2166);
and U2368 (N_2368,N_2112,N_2229);
or U2369 (N_2369,N_2174,N_2233);
xor U2370 (N_2370,N_2240,N_2219);
nand U2371 (N_2371,N_2245,N_2117);
nor U2372 (N_2372,N_2194,N_2187);
and U2373 (N_2373,N_2220,N_2228);
nor U2374 (N_2374,N_2150,N_2103);
nor U2375 (N_2375,N_2175,N_2229);
or U2376 (N_2376,N_2130,N_2213);
nor U2377 (N_2377,N_2131,N_2235);
nand U2378 (N_2378,N_2103,N_2185);
nor U2379 (N_2379,N_2146,N_2165);
nor U2380 (N_2380,N_2202,N_2238);
nor U2381 (N_2381,N_2238,N_2199);
or U2382 (N_2382,N_2183,N_2121);
or U2383 (N_2383,N_2149,N_2223);
or U2384 (N_2384,N_2109,N_2204);
and U2385 (N_2385,N_2191,N_2100);
and U2386 (N_2386,N_2128,N_2106);
and U2387 (N_2387,N_2108,N_2147);
nand U2388 (N_2388,N_2115,N_2179);
xnor U2389 (N_2389,N_2188,N_2123);
and U2390 (N_2390,N_2143,N_2115);
xnor U2391 (N_2391,N_2131,N_2151);
and U2392 (N_2392,N_2130,N_2144);
nand U2393 (N_2393,N_2129,N_2213);
and U2394 (N_2394,N_2224,N_2132);
nor U2395 (N_2395,N_2220,N_2221);
nor U2396 (N_2396,N_2110,N_2130);
and U2397 (N_2397,N_2219,N_2162);
nor U2398 (N_2398,N_2114,N_2157);
nand U2399 (N_2399,N_2123,N_2114);
xor U2400 (N_2400,N_2363,N_2289);
or U2401 (N_2401,N_2354,N_2299);
or U2402 (N_2402,N_2393,N_2310);
nor U2403 (N_2403,N_2397,N_2311);
or U2404 (N_2404,N_2366,N_2318);
and U2405 (N_2405,N_2307,N_2344);
nand U2406 (N_2406,N_2385,N_2290);
xnor U2407 (N_2407,N_2297,N_2362);
nor U2408 (N_2408,N_2263,N_2364);
nand U2409 (N_2409,N_2360,N_2296);
xor U2410 (N_2410,N_2250,N_2379);
nand U2411 (N_2411,N_2356,N_2301);
nand U2412 (N_2412,N_2267,N_2367);
xnor U2413 (N_2413,N_2352,N_2317);
xnor U2414 (N_2414,N_2359,N_2348);
or U2415 (N_2415,N_2328,N_2373);
xnor U2416 (N_2416,N_2315,N_2386);
nor U2417 (N_2417,N_2275,N_2351);
nor U2418 (N_2418,N_2293,N_2375);
and U2419 (N_2419,N_2376,N_2336);
and U2420 (N_2420,N_2399,N_2346);
nand U2421 (N_2421,N_2285,N_2277);
nand U2422 (N_2422,N_2276,N_2253);
nor U2423 (N_2423,N_2282,N_2353);
and U2424 (N_2424,N_2323,N_2347);
nand U2425 (N_2425,N_2326,N_2278);
nor U2426 (N_2426,N_2398,N_2370);
or U2427 (N_2427,N_2388,N_2316);
and U2428 (N_2428,N_2339,N_2264);
xor U2429 (N_2429,N_2258,N_2334);
nand U2430 (N_2430,N_2383,N_2343);
and U2431 (N_2431,N_2325,N_2368);
nand U2432 (N_2432,N_2262,N_2371);
nor U2433 (N_2433,N_2377,N_2329);
and U2434 (N_2434,N_2302,N_2279);
nand U2435 (N_2435,N_2303,N_2252);
nor U2436 (N_2436,N_2345,N_2309);
or U2437 (N_2437,N_2389,N_2271);
nor U2438 (N_2438,N_2322,N_2300);
nor U2439 (N_2439,N_2392,N_2298);
nand U2440 (N_2440,N_2292,N_2324);
nor U2441 (N_2441,N_2284,N_2306);
nor U2442 (N_2442,N_2261,N_2270);
xnor U2443 (N_2443,N_2381,N_2280);
xnor U2444 (N_2444,N_2387,N_2361);
nor U2445 (N_2445,N_2327,N_2272);
nor U2446 (N_2446,N_2396,N_2255);
xor U2447 (N_2447,N_2283,N_2286);
xnor U2448 (N_2448,N_2287,N_2294);
xor U2449 (N_2449,N_2358,N_2305);
xor U2450 (N_2450,N_2395,N_2333);
and U2451 (N_2451,N_2357,N_2365);
nand U2452 (N_2452,N_2332,N_2384);
or U2453 (N_2453,N_2268,N_2372);
xnor U2454 (N_2454,N_2338,N_2391);
nor U2455 (N_2455,N_2340,N_2259);
and U2456 (N_2456,N_2320,N_2319);
nand U2457 (N_2457,N_2256,N_2394);
nand U2458 (N_2458,N_2313,N_2291);
nor U2459 (N_2459,N_2269,N_2349);
and U2460 (N_2460,N_2350,N_2341);
and U2461 (N_2461,N_2342,N_2390);
or U2462 (N_2462,N_2265,N_2260);
or U2463 (N_2463,N_2314,N_2335);
nand U2464 (N_2464,N_2281,N_2254);
and U2465 (N_2465,N_2380,N_2337);
xor U2466 (N_2466,N_2378,N_2295);
and U2467 (N_2467,N_2266,N_2308);
nand U2468 (N_2468,N_2321,N_2257);
or U2469 (N_2469,N_2273,N_2330);
and U2470 (N_2470,N_2382,N_2355);
xnor U2471 (N_2471,N_2304,N_2331);
nand U2472 (N_2472,N_2312,N_2274);
nand U2473 (N_2473,N_2288,N_2374);
xnor U2474 (N_2474,N_2369,N_2251);
and U2475 (N_2475,N_2273,N_2372);
or U2476 (N_2476,N_2380,N_2306);
and U2477 (N_2477,N_2392,N_2317);
or U2478 (N_2478,N_2394,N_2361);
nor U2479 (N_2479,N_2320,N_2289);
and U2480 (N_2480,N_2258,N_2378);
xnor U2481 (N_2481,N_2280,N_2265);
nor U2482 (N_2482,N_2377,N_2303);
nand U2483 (N_2483,N_2277,N_2345);
nor U2484 (N_2484,N_2352,N_2306);
xnor U2485 (N_2485,N_2293,N_2354);
or U2486 (N_2486,N_2390,N_2280);
and U2487 (N_2487,N_2260,N_2339);
and U2488 (N_2488,N_2283,N_2341);
and U2489 (N_2489,N_2353,N_2399);
nand U2490 (N_2490,N_2274,N_2303);
xor U2491 (N_2491,N_2372,N_2354);
xor U2492 (N_2492,N_2359,N_2277);
nor U2493 (N_2493,N_2377,N_2260);
and U2494 (N_2494,N_2271,N_2330);
and U2495 (N_2495,N_2276,N_2267);
or U2496 (N_2496,N_2341,N_2290);
or U2497 (N_2497,N_2375,N_2374);
nor U2498 (N_2498,N_2280,N_2285);
or U2499 (N_2499,N_2290,N_2359);
nand U2500 (N_2500,N_2257,N_2330);
xnor U2501 (N_2501,N_2272,N_2308);
or U2502 (N_2502,N_2297,N_2361);
nand U2503 (N_2503,N_2379,N_2361);
xor U2504 (N_2504,N_2336,N_2398);
or U2505 (N_2505,N_2370,N_2284);
and U2506 (N_2506,N_2365,N_2322);
xor U2507 (N_2507,N_2382,N_2386);
nor U2508 (N_2508,N_2269,N_2348);
nor U2509 (N_2509,N_2393,N_2305);
and U2510 (N_2510,N_2394,N_2385);
or U2511 (N_2511,N_2367,N_2295);
and U2512 (N_2512,N_2384,N_2373);
and U2513 (N_2513,N_2319,N_2355);
or U2514 (N_2514,N_2252,N_2355);
or U2515 (N_2515,N_2331,N_2364);
nand U2516 (N_2516,N_2378,N_2360);
xor U2517 (N_2517,N_2386,N_2304);
nand U2518 (N_2518,N_2366,N_2336);
xor U2519 (N_2519,N_2290,N_2260);
nor U2520 (N_2520,N_2300,N_2364);
xnor U2521 (N_2521,N_2317,N_2393);
and U2522 (N_2522,N_2376,N_2326);
xor U2523 (N_2523,N_2289,N_2360);
nand U2524 (N_2524,N_2281,N_2320);
and U2525 (N_2525,N_2338,N_2385);
nand U2526 (N_2526,N_2283,N_2357);
and U2527 (N_2527,N_2383,N_2263);
and U2528 (N_2528,N_2336,N_2256);
or U2529 (N_2529,N_2304,N_2337);
and U2530 (N_2530,N_2359,N_2302);
nor U2531 (N_2531,N_2270,N_2333);
xnor U2532 (N_2532,N_2319,N_2343);
or U2533 (N_2533,N_2339,N_2332);
nand U2534 (N_2534,N_2332,N_2337);
nand U2535 (N_2535,N_2371,N_2369);
xnor U2536 (N_2536,N_2389,N_2331);
and U2537 (N_2537,N_2346,N_2393);
nor U2538 (N_2538,N_2330,N_2260);
nand U2539 (N_2539,N_2270,N_2276);
nand U2540 (N_2540,N_2262,N_2325);
and U2541 (N_2541,N_2306,N_2267);
or U2542 (N_2542,N_2297,N_2294);
nand U2543 (N_2543,N_2327,N_2281);
xnor U2544 (N_2544,N_2266,N_2336);
nand U2545 (N_2545,N_2296,N_2397);
or U2546 (N_2546,N_2295,N_2269);
or U2547 (N_2547,N_2284,N_2312);
nor U2548 (N_2548,N_2250,N_2261);
xnor U2549 (N_2549,N_2257,N_2342);
nand U2550 (N_2550,N_2473,N_2437);
and U2551 (N_2551,N_2500,N_2429);
and U2552 (N_2552,N_2509,N_2477);
or U2553 (N_2553,N_2415,N_2517);
and U2554 (N_2554,N_2432,N_2430);
xnor U2555 (N_2555,N_2458,N_2427);
or U2556 (N_2556,N_2408,N_2405);
and U2557 (N_2557,N_2443,N_2495);
xnor U2558 (N_2558,N_2478,N_2486);
or U2559 (N_2559,N_2439,N_2460);
nor U2560 (N_2560,N_2491,N_2422);
and U2561 (N_2561,N_2526,N_2503);
nor U2562 (N_2562,N_2488,N_2501);
xor U2563 (N_2563,N_2534,N_2521);
and U2564 (N_2564,N_2523,N_2406);
and U2565 (N_2565,N_2410,N_2411);
nor U2566 (N_2566,N_2531,N_2476);
and U2567 (N_2567,N_2515,N_2423);
and U2568 (N_2568,N_2440,N_2483);
nor U2569 (N_2569,N_2434,N_2524);
nand U2570 (N_2570,N_2419,N_2433);
nor U2571 (N_2571,N_2409,N_2431);
nand U2572 (N_2572,N_2442,N_2487);
and U2573 (N_2573,N_2507,N_2412);
or U2574 (N_2574,N_2413,N_2479);
nand U2575 (N_2575,N_2504,N_2513);
xor U2576 (N_2576,N_2428,N_2470);
xor U2577 (N_2577,N_2529,N_2444);
or U2578 (N_2578,N_2485,N_2497);
nor U2579 (N_2579,N_2545,N_2400);
and U2580 (N_2580,N_2541,N_2401);
and U2581 (N_2581,N_2445,N_2516);
nand U2582 (N_2582,N_2455,N_2425);
nor U2583 (N_2583,N_2481,N_2530);
and U2584 (N_2584,N_2493,N_2424);
nor U2585 (N_2585,N_2449,N_2543);
and U2586 (N_2586,N_2540,N_2511);
nand U2587 (N_2587,N_2480,N_2537);
nor U2588 (N_2588,N_2466,N_2402);
xnor U2589 (N_2589,N_2448,N_2520);
or U2590 (N_2590,N_2453,N_2418);
or U2591 (N_2591,N_2414,N_2452);
xnor U2592 (N_2592,N_2417,N_2519);
and U2593 (N_2593,N_2490,N_2514);
or U2594 (N_2594,N_2535,N_2438);
or U2595 (N_2595,N_2538,N_2505);
and U2596 (N_2596,N_2469,N_2461);
xnor U2597 (N_2597,N_2518,N_2489);
nand U2598 (N_2598,N_2435,N_2484);
or U2599 (N_2599,N_2482,N_2512);
nor U2600 (N_2600,N_2462,N_2421);
nand U2601 (N_2601,N_2522,N_2498);
nand U2602 (N_2602,N_2510,N_2536);
xor U2603 (N_2603,N_2471,N_2467);
xnor U2604 (N_2604,N_2463,N_2451);
nor U2605 (N_2605,N_2508,N_2527);
and U2606 (N_2606,N_2464,N_2416);
or U2607 (N_2607,N_2426,N_2454);
nand U2608 (N_2608,N_2502,N_2499);
or U2609 (N_2609,N_2549,N_2547);
and U2610 (N_2610,N_2468,N_2472);
nor U2611 (N_2611,N_2474,N_2492);
or U2612 (N_2612,N_2407,N_2542);
nand U2613 (N_2613,N_2533,N_2494);
xor U2614 (N_2614,N_2450,N_2457);
or U2615 (N_2615,N_2441,N_2456);
xor U2616 (N_2616,N_2446,N_2496);
xor U2617 (N_2617,N_2548,N_2475);
and U2618 (N_2618,N_2532,N_2447);
nor U2619 (N_2619,N_2420,N_2544);
xor U2620 (N_2620,N_2465,N_2404);
nor U2621 (N_2621,N_2459,N_2546);
xor U2622 (N_2622,N_2525,N_2403);
nand U2623 (N_2623,N_2506,N_2528);
or U2624 (N_2624,N_2539,N_2436);
nor U2625 (N_2625,N_2438,N_2523);
nand U2626 (N_2626,N_2426,N_2409);
or U2627 (N_2627,N_2462,N_2504);
and U2628 (N_2628,N_2468,N_2492);
nand U2629 (N_2629,N_2415,N_2429);
and U2630 (N_2630,N_2440,N_2531);
nand U2631 (N_2631,N_2520,N_2417);
and U2632 (N_2632,N_2462,N_2484);
or U2633 (N_2633,N_2516,N_2510);
nor U2634 (N_2634,N_2469,N_2473);
or U2635 (N_2635,N_2538,N_2456);
or U2636 (N_2636,N_2460,N_2536);
and U2637 (N_2637,N_2468,N_2405);
or U2638 (N_2638,N_2439,N_2427);
nor U2639 (N_2639,N_2517,N_2493);
and U2640 (N_2640,N_2415,N_2483);
xor U2641 (N_2641,N_2539,N_2425);
nor U2642 (N_2642,N_2512,N_2450);
and U2643 (N_2643,N_2534,N_2457);
xnor U2644 (N_2644,N_2463,N_2498);
nand U2645 (N_2645,N_2544,N_2523);
or U2646 (N_2646,N_2415,N_2435);
or U2647 (N_2647,N_2519,N_2407);
or U2648 (N_2648,N_2546,N_2472);
or U2649 (N_2649,N_2487,N_2505);
or U2650 (N_2650,N_2477,N_2501);
or U2651 (N_2651,N_2522,N_2470);
nor U2652 (N_2652,N_2529,N_2482);
nand U2653 (N_2653,N_2494,N_2447);
nand U2654 (N_2654,N_2428,N_2440);
or U2655 (N_2655,N_2511,N_2507);
nand U2656 (N_2656,N_2529,N_2408);
and U2657 (N_2657,N_2545,N_2473);
nand U2658 (N_2658,N_2412,N_2461);
nor U2659 (N_2659,N_2460,N_2438);
or U2660 (N_2660,N_2492,N_2521);
nor U2661 (N_2661,N_2512,N_2459);
xor U2662 (N_2662,N_2543,N_2495);
or U2663 (N_2663,N_2458,N_2483);
nand U2664 (N_2664,N_2538,N_2437);
xnor U2665 (N_2665,N_2475,N_2468);
nor U2666 (N_2666,N_2480,N_2512);
nor U2667 (N_2667,N_2412,N_2411);
nor U2668 (N_2668,N_2463,N_2497);
nor U2669 (N_2669,N_2538,N_2515);
and U2670 (N_2670,N_2466,N_2420);
or U2671 (N_2671,N_2470,N_2471);
or U2672 (N_2672,N_2531,N_2478);
and U2673 (N_2673,N_2510,N_2446);
and U2674 (N_2674,N_2510,N_2475);
xor U2675 (N_2675,N_2457,N_2540);
nor U2676 (N_2676,N_2523,N_2443);
xor U2677 (N_2677,N_2535,N_2452);
or U2678 (N_2678,N_2480,N_2447);
or U2679 (N_2679,N_2467,N_2448);
nor U2680 (N_2680,N_2406,N_2473);
nand U2681 (N_2681,N_2485,N_2434);
or U2682 (N_2682,N_2456,N_2478);
or U2683 (N_2683,N_2523,N_2529);
nor U2684 (N_2684,N_2484,N_2517);
xnor U2685 (N_2685,N_2513,N_2488);
and U2686 (N_2686,N_2545,N_2474);
nand U2687 (N_2687,N_2498,N_2521);
nor U2688 (N_2688,N_2546,N_2436);
xor U2689 (N_2689,N_2505,N_2442);
nor U2690 (N_2690,N_2545,N_2528);
nor U2691 (N_2691,N_2528,N_2470);
xnor U2692 (N_2692,N_2520,N_2447);
or U2693 (N_2693,N_2418,N_2484);
nor U2694 (N_2694,N_2498,N_2429);
nor U2695 (N_2695,N_2539,N_2508);
xnor U2696 (N_2696,N_2421,N_2436);
or U2697 (N_2697,N_2438,N_2542);
or U2698 (N_2698,N_2430,N_2403);
or U2699 (N_2699,N_2481,N_2547);
nand U2700 (N_2700,N_2664,N_2658);
and U2701 (N_2701,N_2688,N_2572);
and U2702 (N_2702,N_2565,N_2552);
nand U2703 (N_2703,N_2586,N_2686);
xnor U2704 (N_2704,N_2645,N_2581);
or U2705 (N_2705,N_2588,N_2638);
and U2706 (N_2706,N_2644,N_2598);
nor U2707 (N_2707,N_2673,N_2680);
xor U2708 (N_2708,N_2619,N_2568);
xor U2709 (N_2709,N_2640,N_2639);
or U2710 (N_2710,N_2560,N_2609);
and U2711 (N_2711,N_2555,N_2596);
nor U2712 (N_2712,N_2667,N_2550);
or U2713 (N_2713,N_2659,N_2695);
nand U2714 (N_2714,N_2582,N_2627);
and U2715 (N_2715,N_2583,N_2577);
nor U2716 (N_2716,N_2625,N_2635);
nand U2717 (N_2717,N_2630,N_2672);
and U2718 (N_2718,N_2674,N_2629);
and U2719 (N_2719,N_2636,N_2571);
or U2720 (N_2720,N_2570,N_2553);
nand U2721 (N_2721,N_2601,N_2624);
xor U2722 (N_2722,N_2612,N_2592);
or U2723 (N_2723,N_2590,N_2575);
and U2724 (N_2724,N_2623,N_2566);
xor U2725 (N_2725,N_2668,N_2670);
and U2726 (N_2726,N_2675,N_2613);
nor U2727 (N_2727,N_2681,N_2618);
nand U2728 (N_2728,N_2676,N_2634);
xor U2729 (N_2729,N_2585,N_2696);
nand U2730 (N_2730,N_2648,N_2600);
or U2731 (N_2731,N_2655,N_2628);
nor U2732 (N_2732,N_2578,N_2605);
nor U2733 (N_2733,N_2606,N_2699);
nor U2734 (N_2734,N_2573,N_2642);
nor U2735 (N_2735,N_2621,N_2599);
nor U2736 (N_2736,N_2663,N_2679);
nor U2737 (N_2737,N_2656,N_2554);
and U2738 (N_2738,N_2692,N_2567);
or U2739 (N_2739,N_2652,N_2631);
xor U2740 (N_2740,N_2689,N_2595);
and U2741 (N_2741,N_2690,N_2579);
nand U2742 (N_2742,N_2671,N_2661);
xor U2743 (N_2743,N_2591,N_2620);
xnor U2744 (N_2744,N_2587,N_2647);
nand U2745 (N_2745,N_2589,N_2693);
nor U2746 (N_2746,N_2564,N_2683);
and U2747 (N_2747,N_2641,N_2684);
nor U2748 (N_2748,N_2657,N_2559);
xor U2749 (N_2749,N_2584,N_2615);
and U2750 (N_2750,N_2593,N_2614);
nor U2751 (N_2751,N_2604,N_2602);
and U2752 (N_2752,N_2563,N_2687);
or U2753 (N_2753,N_2643,N_2646);
and U2754 (N_2754,N_2653,N_2561);
and U2755 (N_2755,N_2685,N_2662);
xnor U2756 (N_2756,N_2569,N_2649);
nand U2757 (N_2757,N_2691,N_2597);
and U2758 (N_2758,N_2651,N_2650);
nand U2759 (N_2759,N_2580,N_2637);
nand U2760 (N_2760,N_2682,N_2576);
nor U2761 (N_2761,N_2660,N_2617);
nand U2762 (N_2762,N_2654,N_2574);
nand U2763 (N_2763,N_2698,N_2666);
and U2764 (N_2764,N_2607,N_2611);
or U2765 (N_2765,N_2603,N_2665);
and U2766 (N_2766,N_2622,N_2626);
nor U2767 (N_2767,N_2558,N_2694);
nand U2768 (N_2768,N_2616,N_2610);
and U2769 (N_2769,N_2669,N_2594);
nand U2770 (N_2770,N_2678,N_2677);
or U2771 (N_2771,N_2551,N_2557);
nand U2772 (N_2772,N_2632,N_2556);
xnor U2773 (N_2773,N_2697,N_2608);
or U2774 (N_2774,N_2633,N_2562);
xnor U2775 (N_2775,N_2576,N_2638);
nor U2776 (N_2776,N_2589,N_2677);
nand U2777 (N_2777,N_2579,N_2551);
xnor U2778 (N_2778,N_2679,N_2692);
nand U2779 (N_2779,N_2655,N_2686);
and U2780 (N_2780,N_2663,N_2602);
xor U2781 (N_2781,N_2551,N_2575);
and U2782 (N_2782,N_2606,N_2557);
nand U2783 (N_2783,N_2620,N_2583);
nand U2784 (N_2784,N_2596,N_2595);
or U2785 (N_2785,N_2596,N_2611);
and U2786 (N_2786,N_2653,N_2652);
or U2787 (N_2787,N_2611,N_2556);
or U2788 (N_2788,N_2607,N_2557);
xor U2789 (N_2789,N_2637,N_2599);
nor U2790 (N_2790,N_2654,N_2583);
xnor U2791 (N_2791,N_2684,N_2588);
nand U2792 (N_2792,N_2560,N_2664);
and U2793 (N_2793,N_2668,N_2629);
and U2794 (N_2794,N_2597,N_2616);
nand U2795 (N_2795,N_2697,N_2605);
nor U2796 (N_2796,N_2658,N_2590);
and U2797 (N_2797,N_2638,N_2652);
nor U2798 (N_2798,N_2597,N_2614);
and U2799 (N_2799,N_2561,N_2628);
or U2800 (N_2800,N_2593,N_2570);
nand U2801 (N_2801,N_2563,N_2694);
and U2802 (N_2802,N_2668,N_2574);
nor U2803 (N_2803,N_2568,N_2641);
nor U2804 (N_2804,N_2663,N_2680);
nor U2805 (N_2805,N_2692,N_2553);
xnor U2806 (N_2806,N_2602,N_2558);
xor U2807 (N_2807,N_2678,N_2635);
nand U2808 (N_2808,N_2599,N_2674);
nor U2809 (N_2809,N_2570,N_2638);
and U2810 (N_2810,N_2555,N_2653);
and U2811 (N_2811,N_2609,N_2581);
nand U2812 (N_2812,N_2653,N_2574);
or U2813 (N_2813,N_2637,N_2671);
or U2814 (N_2814,N_2567,N_2634);
nand U2815 (N_2815,N_2607,N_2696);
and U2816 (N_2816,N_2698,N_2555);
nand U2817 (N_2817,N_2568,N_2690);
and U2818 (N_2818,N_2561,N_2550);
nor U2819 (N_2819,N_2558,N_2693);
or U2820 (N_2820,N_2568,N_2682);
nand U2821 (N_2821,N_2634,N_2655);
or U2822 (N_2822,N_2658,N_2680);
xnor U2823 (N_2823,N_2693,N_2669);
nor U2824 (N_2824,N_2646,N_2620);
nor U2825 (N_2825,N_2656,N_2618);
nor U2826 (N_2826,N_2597,N_2638);
nor U2827 (N_2827,N_2690,N_2552);
nor U2828 (N_2828,N_2610,N_2633);
or U2829 (N_2829,N_2647,N_2658);
and U2830 (N_2830,N_2614,N_2694);
xor U2831 (N_2831,N_2592,N_2694);
nand U2832 (N_2832,N_2667,N_2639);
xnor U2833 (N_2833,N_2618,N_2608);
nor U2834 (N_2834,N_2672,N_2698);
nor U2835 (N_2835,N_2555,N_2680);
nor U2836 (N_2836,N_2697,N_2677);
nand U2837 (N_2837,N_2657,N_2651);
xor U2838 (N_2838,N_2651,N_2587);
nand U2839 (N_2839,N_2606,N_2647);
nand U2840 (N_2840,N_2586,N_2672);
and U2841 (N_2841,N_2674,N_2581);
xor U2842 (N_2842,N_2664,N_2587);
nor U2843 (N_2843,N_2678,N_2686);
nor U2844 (N_2844,N_2672,N_2690);
nand U2845 (N_2845,N_2696,N_2583);
or U2846 (N_2846,N_2562,N_2665);
xor U2847 (N_2847,N_2550,N_2581);
nand U2848 (N_2848,N_2697,N_2669);
or U2849 (N_2849,N_2681,N_2652);
nor U2850 (N_2850,N_2788,N_2836);
and U2851 (N_2851,N_2775,N_2732);
and U2852 (N_2852,N_2751,N_2748);
nand U2853 (N_2853,N_2796,N_2703);
xor U2854 (N_2854,N_2705,N_2780);
xnor U2855 (N_2855,N_2849,N_2835);
xor U2856 (N_2856,N_2818,N_2839);
or U2857 (N_2857,N_2706,N_2712);
nor U2858 (N_2858,N_2816,N_2797);
nand U2859 (N_2859,N_2746,N_2726);
and U2860 (N_2860,N_2792,N_2795);
or U2861 (N_2861,N_2725,N_2729);
or U2862 (N_2862,N_2824,N_2762);
and U2863 (N_2863,N_2700,N_2822);
xnor U2864 (N_2864,N_2769,N_2845);
nor U2865 (N_2865,N_2842,N_2757);
nand U2866 (N_2866,N_2765,N_2728);
or U2867 (N_2867,N_2803,N_2782);
and U2868 (N_2868,N_2791,N_2801);
nor U2869 (N_2869,N_2814,N_2794);
and U2870 (N_2870,N_2826,N_2740);
nor U2871 (N_2871,N_2830,N_2766);
or U2872 (N_2872,N_2808,N_2711);
xor U2873 (N_2873,N_2734,N_2821);
nor U2874 (N_2874,N_2843,N_2846);
nand U2875 (N_2875,N_2815,N_2767);
and U2876 (N_2876,N_2749,N_2825);
nand U2877 (N_2877,N_2848,N_2753);
xnor U2878 (N_2878,N_2736,N_2754);
nor U2879 (N_2879,N_2781,N_2752);
nand U2880 (N_2880,N_2829,N_2770);
nor U2881 (N_2881,N_2776,N_2722);
or U2882 (N_2882,N_2745,N_2798);
nor U2883 (N_2883,N_2727,N_2760);
nor U2884 (N_2884,N_2723,N_2755);
nand U2885 (N_2885,N_2789,N_2840);
nand U2886 (N_2886,N_2820,N_2730);
nor U2887 (N_2887,N_2817,N_2810);
and U2888 (N_2888,N_2714,N_2758);
or U2889 (N_2889,N_2811,N_2793);
and U2890 (N_2890,N_2716,N_2715);
or U2891 (N_2891,N_2779,N_2783);
or U2892 (N_2892,N_2717,N_2771);
nor U2893 (N_2893,N_2731,N_2806);
xnor U2894 (N_2894,N_2805,N_2784);
or U2895 (N_2895,N_2813,N_2764);
nor U2896 (N_2896,N_2790,N_2744);
xnor U2897 (N_2897,N_2763,N_2713);
or U2898 (N_2898,N_2787,N_2809);
xor U2899 (N_2899,N_2719,N_2823);
nand U2900 (N_2900,N_2802,N_2701);
xnor U2901 (N_2901,N_2733,N_2738);
xnor U2902 (N_2902,N_2831,N_2804);
xor U2903 (N_2903,N_2710,N_2743);
and U2904 (N_2904,N_2747,N_2844);
xnor U2905 (N_2905,N_2837,N_2841);
nand U2906 (N_2906,N_2759,N_2709);
or U2907 (N_2907,N_2721,N_2702);
nand U2908 (N_2908,N_2774,N_2739);
xor U2909 (N_2909,N_2756,N_2704);
or U2910 (N_2910,N_2724,N_2827);
and U2911 (N_2911,N_2800,N_2737);
or U2912 (N_2912,N_2799,N_2832);
and U2913 (N_2913,N_2828,N_2807);
xnor U2914 (N_2914,N_2750,N_2707);
xor U2915 (N_2915,N_2777,N_2847);
or U2916 (N_2916,N_2741,N_2708);
xor U2917 (N_2917,N_2838,N_2718);
and U2918 (N_2918,N_2778,N_2785);
nor U2919 (N_2919,N_2773,N_2742);
or U2920 (N_2920,N_2833,N_2720);
xnor U2921 (N_2921,N_2772,N_2812);
nand U2922 (N_2922,N_2761,N_2786);
and U2923 (N_2923,N_2735,N_2819);
xnor U2924 (N_2924,N_2834,N_2768);
xor U2925 (N_2925,N_2792,N_2821);
xor U2926 (N_2926,N_2797,N_2732);
xnor U2927 (N_2927,N_2772,N_2800);
or U2928 (N_2928,N_2711,N_2749);
nor U2929 (N_2929,N_2803,N_2817);
xnor U2930 (N_2930,N_2819,N_2822);
nand U2931 (N_2931,N_2741,N_2812);
and U2932 (N_2932,N_2771,N_2812);
and U2933 (N_2933,N_2778,N_2716);
xnor U2934 (N_2934,N_2808,N_2769);
xor U2935 (N_2935,N_2731,N_2739);
or U2936 (N_2936,N_2795,N_2794);
nand U2937 (N_2937,N_2835,N_2766);
or U2938 (N_2938,N_2705,N_2740);
nor U2939 (N_2939,N_2841,N_2782);
or U2940 (N_2940,N_2812,N_2716);
nor U2941 (N_2941,N_2814,N_2812);
and U2942 (N_2942,N_2768,N_2778);
nor U2943 (N_2943,N_2765,N_2759);
and U2944 (N_2944,N_2718,N_2724);
or U2945 (N_2945,N_2832,N_2778);
nor U2946 (N_2946,N_2788,N_2798);
or U2947 (N_2947,N_2820,N_2700);
or U2948 (N_2948,N_2735,N_2816);
xor U2949 (N_2949,N_2736,N_2741);
and U2950 (N_2950,N_2837,N_2744);
nand U2951 (N_2951,N_2825,N_2707);
nand U2952 (N_2952,N_2705,N_2734);
and U2953 (N_2953,N_2818,N_2737);
nor U2954 (N_2954,N_2789,N_2803);
xor U2955 (N_2955,N_2738,N_2800);
xor U2956 (N_2956,N_2786,N_2711);
nor U2957 (N_2957,N_2703,N_2748);
nor U2958 (N_2958,N_2744,N_2764);
xnor U2959 (N_2959,N_2787,N_2781);
xnor U2960 (N_2960,N_2714,N_2794);
or U2961 (N_2961,N_2826,N_2737);
or U2962 (N_2962,N_2738,N_2812);
and U2963 (N_2963,N_2788,N_2792);
xor U2964 (N_2964,N_2701,N_2703);
xnor U2965 (N_2965,N_2711,N_2725);
nor U2966 (N_2966,N_2804,N_2836);
or U2967 (N_2967,N_2825,N_2782);
and U2968 (N_2968,N_2711,N_2775);
nor U2969 (N_2969,N_2809,N_2756);
or U2970 (N_2970,N_2791,N_2817);
xnor U2971 (N_2971,N_2783,N_2727);
or U2972 (N_2972,N_2710,N_2744);
nand U2973 (N_2973,N_2760,N_2748);
and U2974 (N_2974,N_2817,N_2768);
xnor U2975 (N_2975,N_2713,N_2751);
or U2976 (N_2976,N_2777,N_2831);
or U2977 (N_2977,N_2765,N_2762);
xor U2978 (N_2978,N_2818,N_2831);
and U2979 (N_2979,N_2796,N_2791);
or U2980 (N_2980,N_2803,N_2718);
nor U2981 (N_2981,N_2818,N_2749);
xor U2982 (N_2982,N_2800,N_2742);
xor U2983 (N_2983,N_2806,N_2826);
and U2984 (N_2984,N_2807,N_2745);
or U2985 (N_2985,N_2794,N_2712);
or U2986 (N_2986,N_2718,N_2773);
and U2987 (N_2987,N_2729,N_2773);
xor U2988 (N_2988,N_2746,N_2836);
or U2989 (N_2989,N_2788,N_2775);
xor U2990 (N_2990,N_2732,N_2713);
or U2991 (N_2991,N_2820,N_2829);
nand U2992 (N_2992,N_2783,N_2750);
nand U2993 (N_2993,N_2739,N_2725);
nand U2994 (N_2994,N_2706,N_2730);
or U2995 (N_2995,N_2806,N_2736);
and U2996 (N_2996,N_2753,N_2731);
nand U2997 (N_2997,N_2804,N_2782);
nor U2998 (N_2998,N_2799,N_2844);
and U2999 (N_2999,N_2834,N_2704);
and U3000 (N_3000,N_2880,N_2933);
xnor U3001 (N_3001,N_2958,N_2985);
nand U3002 (N_3002,N_2912,N_2938);
and U3003 (N_3003,N_2910,N_2855);
xnor U3004 (N_3004,N_2991,N_2995);
and U3005 (N_3005,N_2914,N_2884);
xnor U3006 (N_3006,N_2960,N_2881);
nand U3007 (N_3007,N_2871,N_2930);
nand U3008 (N_3008,N_2886,N_2916);
or U3009 (N_3009,N_2962,N_2997);
nand U3010 (N_3010,N_2926,N_2919);
and U3011 (N_3011,N_2992,N_2892);
nor U3012 (N_3012,N_2878,N_2925);
and U3013 (N_3013,N_2928,N_2856);
and U3014 (N_3014,N_2896,N_2969);
nor U3015 (N_3015,N_2959,N_2851);
nor U3016 (N_3016,N_2929,N_2874);
nand U3017 (N_3017,N_2879,N_2857);
xor U3018 (N_3018,N_2966,N_2872);
nor U3019 (N_3019,N_2976,N_2898);
and U3020 (N_3020,N_2924,N_2998);
and U3021 (N_3021,N_2935,N_2980);
nand U3022 (N_3022,N_2890,N_2852);
nor U3023 (N_3023,N_2887,N_2865);
and U3024 (N_3024,N_2949,N_2902);
xor U3025 (N_3025,N_2940,N_2897);
or U3026 (N_3026,N_2868,N_2955);
or U3027 (N_3027,N_2971,N_2920);
or U3028 (N_3028,N_2999,N_2888);
nand U3029 (N_3029,N_2983,N_2921);
or U3030 (N_3030,N_2883,N_2970);
nor U3031 (N_3031,N_2987,N_2864);
nor U3032 (N_3032,N_2946,N_2931);
xnor U3033 (N_3033,N_2917,N_2978);
xnor U3034 (N_3034,N_2950,N_2953);
or U3035 (N_3035,N_2965,N_2901);
nand U3036 (N_3036,N_2984,N_2952);
xor U3037 (N_3037,N_2894,N_2968);
or U3038 (N_3038,N_2945,N_2891);
nor U3039 (N_3039,N_2850,N_2957);
nor U3040 (N_3040,N_2909,N_2990);
nor U3041 (N_3041,N_2853,N_2932);
or U3042 (N_3042,N_2936,N_2911);
nand U3043 (N_3043,N_2963,N_2906);
xor U3044 (N_3044,N_2904,N_2981);
xor U3045 (N_3045,N_2972,N_2895);
and U3046 (N_3046,N_2988,N_2903);
and U3047 (N_3047,N_2875,N_2882);
or U3048 (N_3048,N_2893,N_2908);
nor U3049 (N_3049,N_2885,N_2961);
and U3050 (N_3050,N_2859,N_2867);
or U3051 (N_3051,N_2934,N_2964);
or U3052 (N_3052,N_2861,N_2900);
nor U3053 (N_3053,N_2907,N_2913);
nand U3054 (N_3054,N_2923,N_2956);
and U3055 (N_3055,N_2876,N_2905);
or U3056 (N_3056,N_2877,N_2967);
or U3057 (N_3057,N_2860,N_2873);
or U3058 (N_3058,N_2941,N_2986);
nand U3059 (N_3059,N_2973,N_2870);
or U3060 (N_3060,N_2948,N_2858);
nand U3061 (N_3061,N_2996,N_2977);
or U3062 (N_3062,N_2982,N_2954);
and U3063 (N_3063,N_2918,N_2927);
or U3064 (N_3064,N_2947,N_2989);
xnor U3065 (N_3065,N_2974,N_2994);
and U3066 (N_3066,N_2854,N_2922);
or U3067 (N_3067,N_2863,N_2942);
nor U3068 (N_3068,N_2944,N_2869);
or U3069 (N_3069,N_2975,N_2899);
nor U3070 (N_3070,N_2866,N_2939);
or U3071 (N_3071,N_2943,N_2862);
or U3072 (N_3072,N_2951,N_2889);
or U3073 (N_3073,N_2979,N_2993);
nor U3074 (N_3074,N_2937,N_2915);
and U3075 (N_3075,N_2912,N_2914);
and U3076 (N_3076,N_2997,N_2969);
nor U3077 (N_3077,N_2879,N_2909);
xnor U3078 (N_3078,N_2986,N_2882);
xnor U3079 (N_3079,N_2947,N_2967);
or U3080 (N_3080,N_2856,N_2964);
or U3081 (N_3081,N_2942,N_2980);
or U3082 (N_3082,N_2872,N_2915);
xnor U3083 (N_3083,N_2929,N_2969);
and U3084 (N_3084,N_2894,N_2905);
and U3085 (N_3085,N_2875,N_2879);
and U3086 (N_3086,N_2868,N_2897);
and U3087 (N_3087,N_2856,N_2999);
xor U3088 (N_3088,N_2884,N_2954);
and U3089 (N_3089,N_2942,N_2952);
and U3090 (N_3090,N_2878,N_2922);
or U3091 (N_3091,N_2867,N_2987);
nor U3092 (N_3092,N_2861,N_2992);
and U3093 (N_3093,N_2999,N_2962);
or U3094 (N_3094,N_2874,N_2915);
xnor U3095 (N_3095,N_2960,N_2885);
xor U3096 (N_3096,N_2971,N_2910);
nand U3097 (N_3097,N_2941,N_2938);
nor U3098 (N_3098,N_2991,N_2986);
nand U3099 (N_3099,N_2940,N_2996);
xnor U3100 (N_3100,N_2910,N_2915);
nor U3101 (N_3101,N_2942,N_2886);
and U3102 (N_3102,N_2960,N_2906);
nor U3103 (N_3103,N_2929,N_2863);
or U3104 (N_3104,N_2924,N_2973);
nand U3105 (N_3105,N_2987,N_2944);
and U3106 (N_3106,N_2941,N_2931);
and U3107 (N_3107,N_2972,N_2898);
xnor U3108 (N_3108,N_2915,N_2893);
or U3109 (N_3109,N_2906,N_2902);
nor U3110 (N_3110,N_2918,N_2925);
nand U3111 (N_3111,N_2925,N_2876);
nand U3112 (N_3112,N_2967,N_2869);
nand U3113 (N_3113,N_2944,N_2931);
or U3114 (N_3114,N_2916,N_2969);
xnor U3115 (N_3115,N_2948,N_2887);
or U3116 (N_3116,N_2863,N_2878);
xnor U3117 (N_3117,N_2976,N_2980);
xor U3118 (N_3118,N_2991,N_2865);
xor U3119 (N_3119,N_2942,N_2944);
and U3120 (N_3120,N_2873,N_2952);
nor U3121 (N_3121,N_2885,N_2956);
xor U3122 (N_3122,N_2943,N_2931);
nor U3123 (N_3123,N_2858,N_2994);
nand U3124 (N_3124,N_2905,N_2940);
and U3125 (N_3125,N_2987,N_2930);
nor U3126 (N_3126,N_2908,N_2990);
nor U3127 (N_3127,N_2889,N_2910);
or U3128 (N_3128,N_2872,N_2858);
or U3129 (N_3129,N_2940,N_2945);
nor U3130 (N_3130,N_2986,N_2935);
nand U3131 (N_3131,N_2908,N_2961);
nand U3132 (N_3132,N_2975,N_2940);
xnor U3133 (N_3133,N_2911,N_2988);
nand U3134 (N_3134,N_2902,N_2915);
nand U3135 (N_3135,N_2964,N_2943);
and U3136 (N_3136,N_2920,N_2880);
nand U3137 (N_3137,N_2911,N_2908);
nand U3138 (N_3138,N_2923,N_2913);
nor U3139 (N_3139,N_2956,N_2929);
or U3140 (N_3140,N_2954,N_2987);
nand U3141 (N_3141,N_2973,N_2944);
or U3142 (N_3142,N_2859,N_2915);
or U3143 (N_3143,N_2858,N_2934);
nor U3144 (N_3144,N_2961,N_2910);
and U3145 (N_3145,N_2959,N_2991);
nand U3146 (N_3146,N_2899,N_2992);
xnor U3147 (N_3147,N_2882,N_2852);
or U3148 (N_3148,N_2992,N_2974);
nor U3149 (N_3149,N_2933,N_2862);
nor U3150 (N_3150,N_3036,N_3064);
nor U3151 (N_3151,N_3073,N_3030);
nor U3152 (N_3152,N_3117,N_3074);
and U3153 (N_3153,N_3069,N_3054);
xor U3154 (N_3154,N_3127,N_3094);
or U3155 (N_3155,N_3115,N_3021);
or U3156 (N_3156,N_3012,N_3029);
and U3157 (N_3157,N_3035,N_3131);
or U3158 (N_3158,N_3050,N_3134);
or U3159 (N_3159,N_3038,N_3007);
and U3160 (N_3160,N_3025,N_3044);
xor U3161 (N_3161,N_3121,N_3002);
nor U3162 (N_3162,N_3106,N_3084);
nor U3163 (N_3163,N_3087,N_3057);
xnor U3164 (N_3164,N_3081,N_3129);
and U3165 (N_3165,N_3022,N_3041);
nand U3166 (N_3166,N_3070,N_3143);
nor U3167 (N_3167,N_3120,N_3045);
xnor U3168 (N_3168,N_3093,N_3104);
nor U3169 (N_3169,N_3048,N_3008);
xor U3170 (N_3170,N_3149,N_3001);
xnor U3171 (N_3171,N_3031,N_3138);
and U3172 (N_3172,N_3090,N_3013);
or U3173 (N_3173,N_3046,N_3072);
nand U3174 (N_3174,N_3082,N_3039);
or U3175 (N_3175,N_3078,N_3068);
xor U3176 (N_3176,N_3133,N_3040);
or U3177 (N_3177,N_3124,N_3111);
nor U3178 (N_3178,N_3066,N_3098);
or U3179 (N_3179,N_3023,N_3063);
nand U3180 (N_3180,N_3055,N_3095);
nor U3181 (N_3181,N_3026,N_3005);
or U3182 (N_3182,N_3062,N_3125);
nand U3183 (N_3183,N_3059,N_3071);
xnor U3184 (N_3184,N_3010,N_3102);
nor U3185 (N_3185,N_3088,N_3146);
nand U3186 (N_3186,N_3032,N_3122);
or U3187 (N_3187,N_3105,N_3142);
nand U3188 (N_3188,N_3006,N_3101);
and U3189 (N_3189,N_3085,N_3080);
nor U3190 (N_3190,N_3027,N_3060);
or U3191 (N_3191,N_3089,N_3037);
xnor U3192 (N_3192,N_3003,N_3028);
and U3193 (N_3193,N_3053,N_3096);
nor U3194 (N_3194,N_3083,N_3019);
nand U3195 (N_3195,N_3017,N_3067);
nand U3196 (N_3196,N_3148,N_3015);
and U3197 (N_3197,N_3092,N_3100);
nor U3198 (N_3198,N_3043,N_3014);
nor U3199 (N_3199,N_3033,N_3110);
or U3200 (N_3200,N_3123,N_3077);
nand U3201 (N_3201,N_3056,N_3034);
xnor U3202 (N_3202,N_3061,N_3049);
nor U3203 (N_3203,N_3075,N_3147);
and U3204 (N_3204,N_3145,N_3116);
nand U3205 (N_3205,N_3103,N_3058);
nand U3206 (N_3206,N_3132,N_3108);
or U3207 (N_3207,N_3144,N_3000);
and U3208 (N_3208,N_3139,N_3136);
nor U3209 (N_3209,N_3091,N_3112);
or U3210 (N_3210,N_3042,N_3119);
nand U3211 (N_3211,N_3079,N_3107);
nor U3212 (N_3212,N_3020,N_3140);
and U3213 (N_3213,N_3065,N_3076);
or U3214 (N_3214,N_3024,N_3099);
nor U3215 (N_3215,N_3128,N_3113);
or U3216 (N_3216,N_3047,N_3004);
xor U3217 (N_3217,N_3016,N_3130);
nand U3218 (N_3218,N_3114,N_3137);
or U3219 (N_3219,N_3009,N_3118);
or U3220 (N_3220,N_3141,N_3109);
xor U3221 (N_3221,N_3052,N_3086);
nand U3222 (N_3222,N_3018,N_3011);
nand U3223 (N_3223,N_3051,N_3135);
nand U3224 (N_3224,N_3097,N_3126);
xor U3225 (N_3225,N_3081,N_3092);
nor U3226 (N_3226,N_3101,N_3029);
nor U3227 (N_3227,N_3128,N_3023);
nand U3228 (N_3228,N_3131,N_3115);
and U3229 (N_3229,N_3115,N_3078);
xor U3230 (N_3230,N_3060,N_3066);
nand U3231 (N_3231,N_3096,N_3144);
xnor U3232 (N_3232,N_3020,N_3108);
and U3233 (N_3233,N_3010,N_3092);
or U3234 (N_3234,N_3015,N_3109);
or U3235 (N_3235,N_3089,N_3010);
or U3236 (N_3236,N_3146,N_3094);
nor U3237 (N_3237,N_3130,N_3045);
and U3238 (N_3238,N_3121,N_3149);
xnor U3239 (N_3239,N_3042,N_3031);
and U3240 (N_3240,N_3019,N_3089);
or U3241 (N_3241,N_3041,N_3080);
nor U3242 (N_3242,N_3004,N_3117);
xnor U3243 (N_3243,N_3043,N_3025);
xor U3244 (N_3244,N_3072,N_3132);
xor U3245 (N_3245,N_3133,N_3122);
nand U3246 (N_3246,N_3077,N_3082);
nor U3247 (N_3247,N_3059,N_3082);
nand U3248 (N_3248,N_3141,N_3128);
nand U3249 (N_3249,N_3051,N_3028);
xor U3250 (N_3250,N_3093,N_3120);
nor U3251 (N_3251,N_3012,N_3107);
and U3252 (N_3252,N_3049,N_3073);
nor U3253 (N_3253,N_3086,N_3064);
and U3254 (N_3254,N_3015,N_3099);
or U3255 (N_3255,N_3049,N_3048);
and U3256 (N_3256,N_3091,N_3137);
xor U3257 (N_3257,N_3088,N_3134);
nand U3258 (N_3258,N_3042,N_3100);
nand U3259 (N_3259,N_3040,N_3113);
or U3260 (N_3260,N_3064,N_3045);
and U3261 (N_3261,N_3004,N_3048);
and U3262 (N_3262,N_3118,N_3123);
and U3263 (N_3263,N_3056,N_3067);
or U3264 (N_3264,N_3078,N_3137);
and U3265 (N_3265,N_3017,N_3131);
xnor U3266 (N_3266,N_3049,N_3078);
nor U3267 (N_3267,N_3054,N_3067);
nand U3268 (N_3268,N_3126,N_3110);
nand U3269 (N_3269,N_3118,N_3024);
nor U3270 (N_3270,N_3010,N_3115);
nor U3271 (N_3271,N_3017,N_3071);
nor U3272 (N_3272,N_3036,N_3033);
or U3273 (N_3273,N_3116,N_3047);
nor U3274 (N_3274,N_3111,N_3059);
and U3275 (N_3275,N_3084,N_3105);
or U3276 (N_3276,N_3034,N_3117);
nor U3277 (N_3277,N_3135,N_3033);
and U3278 (N_3278,N_3044,N_3047);
nand U3279 (N_3279,N_3072,N_3042);
nand U3280 (N_3280,N_3112,N_3122);
nand U3281 (N_3281,N_3073,N_3102);
nand U3282 (N_3282,N_3018,N_3141);
or U3283 (N_3283,N_3035,N_3002);
nor U3284 (N_3284,N_3009,N_3096);
nor U3285 (N_3285,N_3029,N_3037);
xor U3286 (N_3286,N_3136,N_3005);
or U3287 (N_3287,N_3129,N_3053);
nand U3288 (N_3288,N_3083,N_3043);
or U3289 (N_3289,N_3115,N_3011);
nand U3290 (N_3290,N_3037,N_3093);
and U3291 (N_3291,N_3133,N_3041);
nand U3292 (N_3292,N_3042,N_3103);
nand U3293 (N_3293,N_3068,N_3149);
xor U3294 (N_3294,N_3072,N_3032);
nand U3295 (N_3295,N_3027,N_3073);
nor U3296 (N_3296,N_3116,N_3149);
nor U3297 (N_3297,N_3091,N_3104);
nand U3298 (N_3298,N_3027,N_3128);
or U3299 (N_3299,N_3005,N_3070);
and U3300 (N_3300,N_3254,N_3171);
nor U3301 (N_3301,N_3165,N_3232);
nor U3302 (N_3302,N_3278,N_3219);
or U3303 (N_3303,N_3183,N_3271);
xnor U3304 (N_3304,N_3213,N_3262);
xnor U3305 (N_3305,N_3204,N_3273);
nand U3306 (N_3306,N_3186,N_3181);
xnor U3307 (N_3307,N_3276,N_3241);
xnor U3308 (N_3308,N_3228,N_3281);
and U3309 (N_3309,N_3184,N_3237);
nor U3310 (N_3310,N_3260,N_3298);
nor U3311 (N_3311,N_3190,N_3217);
xnor U3312 (N_3312,N_3177,N_3221);
or U3313 (N_3313,N_3272,N_3198);
and U3314 (N_3314,N_3176,N_3191);
xor U3315 (N_3315,N_3253,N_3290);
xor U3316 (N_3316,N_3231,N_3170);
xnor U3317 (N_3317,N_3275,N_3280);
nor U3318 (N_3318,N_3156,N_3182);
nand U3319 (N_3319,N_3267,N_3255);
and U3320 (N_3320,N_3207,N_3222);
xor U3321 (N_3321,N_3268,N_3189);
nor U3322 (N_3322,N_3194,N_3175);
xor U3323 (N_3323,N_3265,N_3153);
nor U3324 (N_3324,N_3244,N_3203);
xor U3325 (N_3325,N_3205,N_3295);
nand U3326 (N_3326,N_3292,N_3226);
xnor U3327 (N_3327,N_3266,N_3235);
and U3328 (N_3328,N_3199,N_3179);
xnor U3329 (N_3329,N_3251,N_3291);
or U3330 (N_3330,N_3178,N_3167);
nor U3331 (N_3331,N_3212,N_3279);
xor U3332 (N_3332,N_3258,N_3214);
nand U3333 (N_3333,N_3158,N_3236);
nand U3334 (N_3334,N_3173,N_3211);
xor U3335 (N_3335,N_3159,N_3169);
or U3336 (N_3336,N_3287,N_3192);
and U3337 (N_3337,N_3261,N_3157);
and U3338 (N_3338,N_3188,N_3166);
nand U3339 (N_3339,N_3282,N_3277);
nand U3340 (N_3340,N_3201,N_3187);
nor U3341 (N_3341,N_3168,N_3155);
or U3342 (N_3342,N_3216,N_3234);
and U3343 (N_3343,N_3296,N_3163);
xnor U3344 (N_3344,N_3224,N_3264);
nor U3345 (N_3345,N_3162,N_3161);
xor U3346 (N_3346,N_3257,N_3154);
and U3347 (N_3347,N_3172,N_3248);
nand U3348 (N_3348,N_3200,N_3283);
nand U3349 (N_3349,N_3197,N_3208);
and U3350 (N_3350,N_3150,N_3239);
nor U3351 (N_3351,N_3256,N_3289);
and U3352 (N_3352,N_3263,N_3229);
nor U3353 (N_3353,N_3246,N_3288);
xnor U3354 (N_3354,N_3180,N_3220);
nor U3355 (N_3355,N_3152,N_3270);
nand U3356 (N_3356,N_3223,N_3206);
nor U3357 (N_3357,N_3174,N_3274);
nor U3358 (N_3358,N_3209,N_3240);
xor U3359 (N_3359,N_3294,N_3250);
or U3360 (N_3360,N_3238,N_3210);
nor U3361 (N_3361,N_3193,N_3247);
nor U3362 (N_3362,N_3164,N_3245);
or U3363 (N_3363,N_3160,N_3252);
and U3364 (N_3364,N_3284,N_3233);
nand U3365 (N_3365,N_3243,N_3286);
xnor U3366 (N_3366,N_3151,N_3227);
or U3367 (N_3367,N_3299,N_3215);
or U3368 (N_3368,N_3297,N_3225);
xor U3369 (N_3369,N_3293,N_3259);
nor U3370 (N_3370,N_3242,N_3195);
or U3371 (N_3371,N_3202,N_3218);
nand U3372 (N_3372,N_3230,N_3185);
and U3373 (N_3373,N_3196,N_3249);
xnor U3374 (N_3374,N_3285,N_3269);
and U3375 (N_3375,N_3237,N_3225);
nor U3376 (N_3376,N_3235,N_3176);
xor U3377 (N_3377,N_3243,N_3258);
and U3378 (N_3378,N_3261,N_3187);
xor U3379 (N_3379,N_3261,N_3212);
nand U3380 (N_3380,N_3292,N_3254);
nor U3381 (N_3381,N_3242,N_3232);
nor U3382 (N_3382,N_3175,N_3267);
and U3383 (N_3383,N_3270,N_3255);
xnor U3384 (N_3384,N_3238,N_3285);
nor U3385 (N_3385,N_3152,N_3179);
nand U3386 (N_3386,N_3160,N_3240);
nor U3387 (N_3387,N_3173,N_3263);
xnor U3388 (N_3388,N_3188,N_3261);
and U3389 (N_3389,N_3207,N_3252);
xnor U3390 (N_3390,N_3285,N_3200);
nand U3391 (N_3391,N_3156,N_3259);
nor U3392 (N_3392,N_3285,N_3206);
xnor U3393 (N_3393,N_3232,N_3237);
xor U3394 (N_3394,N_3253,N_3279);
and U3395 (N_3395,N_3242,N_3175);
xor U3396 (N_3396,N_3242,N_3294);
nand U3397 (N_3397,N_3256,N_3169);
xnor U3398 (N_3398,N_3248,N_3152);
or U3399 (N_3399,N_3291,N_3285);
and U3400 (N_3400,N_3258,N_3170);
or U3401 (N_3401,N_3226,N_3242);
and U3402 (N_3402,N_3261,N_3241);
and U3403 (N_3403,N_3284,N_3293);
nand U3404 (N_3404,N_3167,N_3248);
or U3405 (N_3405,N_3245,N_3258);
or U3406 (N_3406,N_3211,N_3154);
or U3407 (N_3407,N_3235,N_3245);
nor U3408 (N_3408,N_3170,N_3265);
xor U3409 (N_3409,N_3246,N_3174);
or U3410 (N_3410,N_3220,N_3176);
or U3411 (N_3411,N_3272,N_3174);
xnor U3412 (N_3412,N_3245,N_3229);
and U3413 (N_3413,N_3229,N_3296);
nand U3414 (N_3414,N_3252,N_3288);
and U3415 (N_3415,N_3157,N_3274);
nand U3416 (N_3416,N_3159,N_3154);
and U3417 (N_3417,N_3173,N_3235);
nand U3418 (N_3418,N_3179,N_3270);
and U3419 (N_3419,N_3212,N_3216);
xor U3420 (N_3420,N_3291,N_3297);
nor U3421 (N_3421,N_3259,N_3199);
xnor U3422 (N_3422,N_3239,N_3195);
and U3423 (N_3423,N_3155,N_3159);
or U3424 (N_3424,N_3271,N_3272);
or U3425 (N_3425,N_3181,N_3224);
nor U3426 (N_3426,N_3214,N_3253);
nand U3427 (N_3427,N_3194,N_3205);
nand U3428 (N_3428,N_3155,N_3186);
nand U3429 (N_3429,N_3257,N_3296);
nor U3430 (N_3430,N_3166,N_3173);
xnor U3431 (N_3431,N_3211,N_3290);
nor U3432 (N_3432,N_3297,N_3250);
xor U3433 (N_3433,N_3291,N_3235);
nand U3434 (N_3434,N_3252,N_3255);
and U3435 (N_3435,N_3296,N_3249);
nand U3436 (N_3436,N_3206,N_3241);
and U3437 (N_3437,N_3247,N_3164);
and U3438 (N_3438,N_3274,N_3195);
and U3439 (N_3439,N_3209,N_3182);
xnor U3440 (N_3440,N_3221,N_3236);
xnor U3441 (N_3441,N_3162,N_3155);
xnor U3442 (N_3442,N_3286,N_3262);
nand U3443 (N_3443,N_3285,N_3198);
nand U3444 (N_3444,N_3280,N_3289);
nand U3445 (N_3445,N_3165,N_3231);
and U3446 (N_3446,N_3284,N_3294);
or U3447 (N_3447,N_3249,N_3188);
xnor U3448 (N_3448,N_3162,N_3240);
and U3449 (N_3449,N_3235,N_3169);
xnor U3450 (N_3450,N_3347,N_3382);
or U3451 (N_3451,N_3374,N_3375);
nor U3452 (N_3452,N_3430,N_3324);
or U3453 (N_3453,N_3318,N_3412);
or U3454 (N_3454,N_3411,N_3360);
xnor U3455 (N_3455,N_3428,N_3400);
nand U3456 (N_3456,N_3404,N_3418);
or U3457 (N_3457,N_3389,N_3367);
or U3458 (N_3458,N_3442,N_3427);
or U3459 (N_3459,N_3397,N_3387);
nor U3460 (N_3460,N_3363,N_3338);
and U3461 (N_3461,N_3345,N_3386);
and U3462 (N_3462,N_3312,N_3405);
nor U3463 (N_3463,N_3408,N_3316);
nand U3464 (N_3464,N_3393,N_3425);
nor U3465 (N_3465,N_3369,N_3368);
nor U3466 (N_3466,N_3351,N_3438);
nand U3467 (N_3467,N_3334,N_3422);
and U3468 (N_3468,N_3417,N_3445);
xor U3469 (N_3469,N_3407,N_3329);
xnor U3470 (N_3470,N_3413,N_3327);
and U3471 (N_3471,N_3331,N_3305);
or U3472 (N_3472,N_3307,N_3356);
or U3473 (N_3473,N_3362,N_3403);
xnor U3474 (N_3474,N_3301,N_3306);
nand U3475 (N_3475,N_3392,N_3402);
nor U3476 (N_3476,N_3309,N_3359);
nand U3477 (N_3477,N_3373,N_3391);
and U3478 (N_3478,N_3320,N_3381);
or U3479 (N_3479,N_3416,N_3390);
and U3480 (N_3480,N_3419,N_3313);
xnor U3481 (N_3481,N_3343,N_3336);
and U3482 (N_3482,N_3434,N_3401);
xnor U3483 (N_3483,N_3321,N_3439);
xnor U3484 (N_3484,N_3447,N_3429);
nand U3485 (N_3485,N_3361,N_3328);
or U3486 (N_3486,N_3372,N_3437);
nor U3487 (N_3487,N_3352,N_3423);
nand U3488 (N_3488,N_3433,N_3409);
nor U3489 (N_3489,N_3371,N_3326);
nand U3490 (N_3490,N_3365,N_3432);
xnor U3491 (N_3491,N_3317,N_3308);
and U3492 (N_3492,N_3376,N_3380);
nor U3493 (N_3493,N_3384,N_3424);
or U3494 (N_3494,N_3431,N_3446);
nor U3495 (N_3495,N_3344,N_3399);
nand U3496 (N_3496,N_3332,N_3339);
and U3497 (N_3497,N_3366,N_3346);
or U3498 (N_3498,N_3337,N_3342);
nor U3499 (N_3499,N_3394,N_3333);
and U3500 (N_3500,N_3449,N_3304);
xor U3501 (N_3501,N_3421,N_3311);
xor U3502 (N_3502,N_3448,N_3314);
nand U3503 (N_3503,N_3410,N_3440);
nand U3504 (N_3504,N_3300,N_3378);
or U3505 (N_3505,N_3420,N_3323);
or U3506 (N_3506,N_3398,N_3443);
nor U3507 (N_3507,N_3357,N_3340);
and U3508 (N_3508,N_3349,N_3444);
and U3509 (N_3509,N_3325,N_3441);
nand U3510 (N_3510,N_3350,N_3303);
nand U3511 (N_3511,N_3396,N_3355);
nor U3512 (N_3512,N_3348,N_3385);
and U3513 (N_3513,N_3414,N_3426);
and U3514 (N_3514,N_3310,N_3315);
nand U3515 (N_3515,N_3383,N_3395);
xor U3516 (N_3516,N_3353,N_3364);
nand U3517 (N_3517,N_3379,N_3335);
or U3518 (N_3518,N_3322,N_3436);
nand U3519 (N_3519,N_3354,N_3377);
or U3520 (N_3520,N_3415,N_3370);
nor U3521 (N_3521,N_3388,N_3358);
and U3522 (N_3522,N_3435,N_3319);
nor U3523 (N_3523,N_3406,N_3330);
or U3524 (N_3524,N_3341,N_3302);
or U3525 (N_3525,N_3319,N_3395);
nor U3526 (N_3526,N_3370,N_3374);
nand U3527 (N_3527,N_3360,N_3394);
nor U3528 (N_3528,N_3328,N_3435);
or U3529 (N_3529,N_3377,N_3402);
and U3530 (N_3530,N_3432,N_3404);
nor U3531 (N_3531,N_3373,N_3393);
nand U3532 (N_3532,N_3375,N_3357);
or U3533 (N_3533,N_3335,N_3384);
xor U3534 (N_3534,N_3421,N_3371);
xor U3535 (N_3535,N_3355,N_3327);
nor U3536 (N_3536,N_3310,N_3449);
nor U3537 (N_3537,N_3419,N_3436);
nor U3538 (N_3538,N_3412,N_3378);
nand U3539 (N_3539,N_3353,N_3319);
or U3540 (N_3540,N_3371,N_3359);
nor U3541 (N_3541,N_3324,N_3303);
or U3542 (N_3542,N_3329,N_3429);
nor U3543 (N_3543,N_3425,N_3365);
nor U3544 (N_3544,N_3307,N_3318);
xnor U3545 (N_3545,N_3316,N_3344);
and U3546 (N_3546,N_3444,N_3425);
nand U3547 (N_3547,N_3440,N_3365);
or U3548 (N_3548,N_3344,N_3382);
and U3549 (N_3549,N_3343,N_3370);
xor U3550 (N_3550,N_3417,N_3305);
nand U3551 (N_3551,N_3340,N_3325);
or U3552 (N_3552,N_3351,N_3403);
and U3553 (N_3553,N_3378,N_3377);
nand U3554 (N_3554,N_3430,N_3383);
xnor U3555 (N_3555,N_3304,N_3300);
or U3556 (N_3556,N_3397,N_3372);
xnor U3557 (N_3557,N_3302,N_3399);
nand U3558 (N_3558,N_3423,N_3323);
and U3559 (N_3559,N_3389,N_3407);
nor U3560 (N_3560,N_3436,N_3391);
nor U3561 (N_3561,N_3418,N_3440);
nor U3562 (N_3562,N_3355,N_3406);
and U3563 (N_3563,N_3445,N_3318);
and U3564 (N_3564,N_3437,N_3385);
nand U3565 (N_3565,N_3449,N_3401);
and U3566 (N_3566,N_3362,N_3427);
nand U3567 (N_3567,N_3370,N_3329);
nor U3568 (N_3568,N_3388,N_3332);
nor U3569 (N_3569,N_3360,N_3344);
nor U3570 (N_3570,N_3306,N_3333);
or U3571 (N_3571,N_3409,N_3392);
nor U3572 (N_3572,N_3431,N_3421);
nor U3573 (N_3573,N_3313,N_3305);
nand U3574 (N_3574,N_3435,N_3361);
nor U3575 (N_3575,N_3366,N_3306);
nor U3576 (N_3576,N_3437,N_3314);
nor U3577 (N_3577,N_3424,N_3359);
nand U3578 (N_3578,N_3358,N_3341);
xor U3579 (N_3579,N_3401,N_3370);
nor U3580 (N_3580,N_3418,N_3416);
nor U3581 (N_3581,N_3353,N_3317);
nor U3582 (N_3582,N_3304,N_3403);
or U3583 (N_3583,N_3411,N_3315);
xor U3584 (N_3584,N_3401,N_3393);
and U3585 (N_3585,N_3339,N_3310);
nor U3586 (N_3586,N_3354,N_3310);
nand U3587 (N_3587,N_3433,N_3416);
nor U3588 (N_3588,N_3396,N_3412);
or U3589 (N_3589,N_3311,N_3304);
xor U3590 (N_3590,N_3439,N_3373);
xor U3591 (N_3591,N_3449,N_3301);
or U3592 (N_3592,N_3444,N_3422);
xor U3593 (N_3593,N_3431,N_3350);
nor U3594 (N_3594,N_3379,N_3333);
nand U3595 (N_3595,N_3308,N_3381);
nor U3596 (N_3596,N_3414,N_3408);
or U3597 (N_3597,N_3319,N_3372);
or U3598 (N_3598,N_3351,N_3344);
nor U3599 (N_3599,N_3411,N_3397);
and U3600 (N_3600,N_3491,N_3587);
nand U3601 (N_3601,N_3540,N_3493);
nor U3602 (N_3602,N_3497,N_3543);
nand U3603 (N_3603,N_3511,N_3490);
nor U3604 (N_3604,N_3456,N_3506);
xnor U3605 (N_3605,N_3520,N_3564);
or U3606 (N_3606,N_3551,N_3522);
nor U3607 (N_3607,N_3568,N_3527);
and U3608 (N_3608,N_3457,N_3577);
and U3609 (N_3609,N_3598,N_3516);
nor U3610 (N_3610,N_3596,N_3574);
nand U3611 (N_3611,N_3452,N_3459);
nor U3612 (N_3612,N_3525,N_3555);
nor U3613 (N_3613,N_3501,N_3484);
or U3614 (N_3614,N_3559,N_3470);
nor U3615 (N_3615,N_3474,N_3450);
or U3616 (N_3616,N_3544,N_3558);
xnor U3617 (N_3617,N_3451,N_3585);
or U3618 (N_3618,N_3479,N_3510);
nand U3619 (N_3619,N_3513,N_3458);
nor U3620 (N_3620,N_3553,N_3469);
xor U3621 (N_3621,N_3579,N_3461);
and U3622 (N_3622,N_3465,N_3578);
xnor U3623 (N_3623,N_3523,N_3582);
xnor U3624 (N_3624,N_3498,N_3466);
xnor U3625 (N_3625,N_3560,N_3580);
or U3626 (N_3626,N_3489,N_3499);
nor U3627 (N_3627,N_3495,N_3554);
and U3628 (N_3628,N_3533,N_3519);
or U3629 (N_3629,N_3473,N_3486);
nor U3630 (N_3630,N_3531,N_3581);
and U3631 (N_3631,N_3464,N_3562);
and U3632 (N_3632,N_3488,N_3462);
xor U3633 (N_3633,N_3595,N_3512);
nor U3634 (N_3634,N_3463,N_3590);
nand U3635 (N_3635,N_3541,N_3475);
xnor U3636 (N_3636,N_3573,N_3583);
nand U3637 (N_3637,N_3536,N_3570);
xor U3638 (N_3638,N_3478,N_3561);
or U3639 (N_3639,N_3552,N_3539);
nor U3640 (N_3640,N_3548,N_3576);
or U3641 (N_3641,N_3530,N_3584);
nand U3642 (N_3642,N_3467,N_3556);
nor U3643 (N_3643,N_3592,N_3494);
nand U3644 (N_3644,N_3481,N_3594);
nand U3645 (N_3645,N_3485,N_3477);
or U3646 (N_3646,N_3472,N_3455);
and U3647 (N_3647,N_3524,N_3597);
nor U3648 (N_3648,N_3507,N_3476);
nor U3649 (N_3649,N_3487,N_3542);
and U3650 (N_3650,N_3593,N_3502);
and U3651 (N_3651,N_3503,N_3566);
nor U3652 (N_3652,N_3454,N_3550);
nand U3653 (N_3653,N_3528,N_3534);
and U3654 (N_3654,N_3508,N_3535);
or U3655 (N_3655,N_3526,N_3599);
nand U3656 (N_3656,N_3569,N_3588);
xnor U3657 (N_3657,N_3586,N_3529);
nor U3658 (N_3658,N_3496,N_3483);
nand U3659 (N_3659,N_3505,N_3571);
xor U3660 (N_3660,N_3538,N_3471);
nand U3661 (N_3661,N_3460,N_3480);
nand U3662 (N_3662,N_3557,N_3504);
or U3663 (N_3663,N_3545,N_3575);
nand U3664 (N_3664,N_3509,N_3572);
nor U3665 (N_3665,N_3500,N_3515);
nor U3666 (N_3666,N_3468,N_3492);
xnor U3667 (N_3667,N_3521,N_3567);
nand U3668 (N_3668,N_3453,N_3546);
and U3669 (N_3669,N_3589,N_3591);
nor U3670 (N_3670,N_3537,N_3565);
nand U3671 (N_3671,N_3532,N_3563);
xnor U3672 (N_3672,N_3514,N_3547);
nand U3673 (N_3673,N_3517,N_3518);
xnor U3674 (N_3674,N_3549,N_3482);
or U3675 (N_3675,N_3518,N_3555);
nor U3676 (N_3676,N_3512,N_3478);
or U3677 (N_3677,N_3594,N_3592);
and U3678 (N_3678,N_3596,N_3594);
or U3679 (N_3679,N_3486,N_3513);
and U3680 (N_3680,N_3587,N_3498);
xnor U3681 (N_3681,N_3549,N_3502);
xor U3682 (N_3682,N_3529,N_3561);
nand U3683 (N_3683,N_3592,N_3458);
xor U3684 (N_3684,N_3557,N_3596);
or U3685 (N_3685,N_3585,N_3493);
xor U3686 (N_3686,N_3504,N_3474);
or U3687 (N_3687,N_3512,N_3532);
or U3688 (N_3688,N_3462,N_3569);
xor U3689 (N_3689,N_3565,N_3499);
and U3690 (N_3690,N_3597,N_3463);
xnor U3691 (N_3691,N_3584,N_3489);
nand U3692 (N_3692,N_3490,N_3586);
nor U3693 (N_3693,N_3519,N_3570);
nor U3694 (N_3694,N_3577,N_3505);
or U3695 (N_3695,N_3544,N_3454);
or U3696 (N_3696,N_3551,N_3487);
and U3697 (N_3697,N_3485,N_3468);
or U3698 (N_3698,N_3578,N_3551);
nand U3699 (N_3699,N_3454,N_3540);
xnor U3700 (N_3700,N_3585,N_3577);
or U3701 (N_3701,N_3576,N_3522);
nand U3702 (N_3702,N_3520,N_3506);
or U3703 (N_3703,N_3540,N_3462);
xor U3704 (N_3704,N_3575,N_3462);
xor U3705 (N_3705,N_3505,N_3451);
and U3706 (N_3706,N_3578,N_3564);
and U3707 (N_3707,N_3514,N_3588);
and U3708 (N_3708,N_3535,N_3538);
xnor U3709 (N_3709,N_3501,N_3539);
nor U3710 (N_3710,N_3547,N_3553);
xor U3711 (N_3711,N_3523,N_3491);
and U3712 (N_3712,N_3530,N_3474);
or U3713 (N_3713,N_3477,N_3560);
nand U3714 (N_3714,N_3546,N_3597);
and U3715 (N_3715,N_3547,N_3598);
nand U3716 (N_3716,N_3554,N_3501);
xor U3717 (N_3717,N_3575,N_3467);
nor U3718 (N_3718,N_3585,N_3500);
and U3719 (N_3719,N_3507,N_3484);
xnor U3720 (N_3720,N_3461,N_3547);
nand U3721 (N_3721,N_3587,N_3531);
or U3722 (N_3722,N_3515,N_3528);
nor U3723 (N_3723,N_3574,N_3561);
or U3724 (N_3724,N_3559,N_3554);
xor U3725 (N_3725,N_3573,N_3525);
and U3726 (N_3726,N_3521,N_3528);
xor U3727 (N_3727,N_3539,N_3496);
and U3728 (N_3728,N_3597,N_3488);
xor U3729 (N_3729,N_3570,N_3549);
and U3730 (N_3730,N_3590,N_3511);
xnor U3731 (N_3731,N_3517,N_3588);
and U3732 (N_3732,N_3562,N_3555);
or U3733 (N_3733,N_3499,N_3494);
xnor U3734 (N_3734,N_3513,N_3484);
and U3735 (N_3735,N_3522,N_3507);
or U3736 (N_3736,N_3506,N_3498);
xnor U3737 (N_3737,N_3584,N_3573);
or U3738 (N_3738,N_3494,N_3495);
nand U3739 (N_3739,N_3503,N_3572);
nand U3740 (N_3740,N_3528,N_3533);
and U3741 (N_3741,N_3487,N_3528);
or U3742 (N_3742,N_3453,N_3593);
xor U3743 (N_3743,N_3557,N_3469);
or U3744 (N_3744,N_3451,N_3532);
nor U3745 (N_3745,N_3566,N_3465);
xor U3746 (N_3746,N_3533,N_3564);
xor U3747 (N_3747,N_3459,N_3478);
or U3748 (N_3748,N_3490,N_3470);
or U3749 (N_3749,N_3472,N_3533);
and U3750 (N_3750,N_3696,N_3671);
nor U3751 (N_3751,N_3604,N_3639);
nor U3752 (N_3752,N_3676,N_3672);
nand U3753 (N_3753,N_3673,N_3711);
xor U3754 (N_3754,N_3707,N_3685);
xor U3755 (N_3755,N_3718,N_3746);
or U3756 (N_3756,N_3723,N_3636);
nor U3757 (N_3757,N_3675,N_3640);
nand U3758 (N_3758,N_3682,N_3619);
nor U3759 (N_3759,N_3691,N_3627);
nor U3760 (N_3760,N_3611,N_3720);
nand U3761 (N_3761,N_3662,N_3621);
nand U3762 (N_3762,N_3688,N_3724);
and U3763 (N_3763,N_3674,N_3609);
xnor U3764 (N_3764,N_3658,N_3721);
nor U3765 (N_3765,N_3747,N_3679);
nand U3766 (N_3766,N_3706,N_3633);
nor U3767 (N_3767,N_3717,N_3697);
nor U3768 (N_3768,N_3749,N_3622);
nand U3769 (N_3769,N_3702,N_3714);
nor U3770 (N_3770,N_3629,N_3712);
nor U3771 (N_3771,N_3728,N_3738);
nand U3772 (N_3772,N_3722,N_3654);
nand U3773 (N_3773,N_3678,N_3740);
or U3774 (N_3774,N_3715,N_3603);
nand U3775 (N_3775,N_3652,N_3613);
xnor U3776 (N_3776,N_3726,N_3680);
nand U3777 (N_3777,N_3624,N_3687);
xnor U3778 (N_3778,N_3625,N_3745);
nand U3779 (N_3779,N_3735,N_3660);
nor U3780 (N_3780,N_3616,N_3701);
and U3781 (N_3781,N_3642,N_3665);
and U3782 (N_3782,N_3704,N_3607);
nand U3783 (N_3783,N_3661,N_3689);
nand U3784 (N_3784,N_3628,N_3709);
and U3785 (N_3785,N_3666,N_3647);
nand U3786 (N_3786,N_3730,N_3681);
or U3787 (N_3787,N_3641,N_3653);
nor U3788 (N_3788,N_3731,N_3668);
nand U3789 (N_3789,N_3732,N_3686);
xnor U3790 (N_3790,N_3631,N_3612);
or U3791 (N_3791,N_3693,N_3727);
xnor U3792 (N_3792,N_3708,N_3614);
or U3793 (N_3793,N_3618,N_3667);
and U3794 (N_3794,N_3610,N_3734);
or U3795 (N_3795,N_3669,N_3656);
and U3796 (N_3796,N_3637,N_3695);
nand U3797 (N_3797,N_3606,N_3705);
and U3798 (N_3798,N_3655,N_3736);
nor U3799 (N_3799,N_3626,N_3617);
xor U3800 (N_3800,N_3700,N_3684);
nand U3801 (N_3801,N_3743,N_3645);
or U3802 (N_3802,N_3634,N_3649);
nand U3803 (N_3803,N_3690,N_3657);
and U3804 (N_3804,N_3632,N_3659);
xor U3805 (N_3805,N_3670,N_3615);
nor U3806 (N_3806,N_3748,N_3744);
xnor U3807 (N_3807,N_3663,N_3698);
or U3808 (N_3808,N_3733,N_3644);
nor U3809 (N_3809,N_3694,N_3648);
xnor U3810 (N_3810,N_3608,N_3623);
nor U3811 (N_3811,N_3713,N_3630);
and U3812 (N_3812,N_3719,N_3703);
or U3813 (N_3813,N_3638,N_3600);
and U3814 (N_3814,N_3741,N_3710);
nand U3815 (N_3815,N_3739,N_3643);
nand U3816 (N_3816,N_3725,N_3646);
nor U3817 (N_3817,N_3716,N_3683);
and U3818 (N_3818,N_3699,N_3602);
and U3819 (N_3819,N_3635,N_3677);
nor U3820 (N_3820,N_3729,N_3651);
nand U3821 (N_3821,N_3650,N_3742);
xor U3822 (N_3822,N_3601,N_3664);
xor U3823 (N_3823,N_3692,N_3737);
and U3824 (N_3824,N_3620,N_3605);
and U3825 (N_3825,N_3600,N_3734);
and U3826 (N_3826,N_3734,N_3743);
or U3827 (N_3827,N_3716,N_3746);
and U3828 (N_3828,N_3720,N_3697);
nor U3829 (N_3829,N_3674,N_3646);
or U3830 (N_3830,N_3633,N_3623);
xor U3831 (N_3831,N_3705,N_3653);
nor U3832 (N_3832,N_3725,N_3727);
nand U3833 (N_3833,N_3722,N_3695);
nor U3834 (N_3834,N_3705,N_3733);
xnor U3835 (N_3835,N_3667,N_3688);
or U3836 (N_3836,N_3606,N_3610);
xor U3837 (N_3837,N_3732,N_3711);
nor U3838 (N_3838,N_3670,N_3741);
and U3839 (N_3839,N_3624,N_3731);
and U3840 (N_3840,N_3647,N_3726);
xor U3841 (N_3841,N_3738,N_3639);
and U3842 (N_3842,N_3749,N_3735);
and U3843 (N_3843,N_3668,N_3721);
or U3844 (N_3844,N_3722,N_3660);
or U3845 (N_3845,N_3681,N_3643);
nor U3846 (N_3846,N_3652,N_3601);
nor U3847 (N_3847,N_3741,N_3714);
and U3848 (N_3848,N_3635,N_3668);
nand U3849 (N_3849,N_3607,N_3635);
or U3850 (N_3850,N_3709,N_3727);
and U3851 (N_3851,N_3704,N_3696);
xor U3852 (N_3852,N_3624,N_3643);
and U3853 (N_3853,N_3601,N_3670);
nor U3854 (N_3854,N_3730,N_3740);
nor U3855 (N_3855,N_3625,N_3700);
nand U3856 (N_3856,N_3737,N_3627);
and U3857 (N_3857,N_3660,N_3620);
nor U3858 (N_3858,N_3722,N_3693);
or U3859 (N_3859,N_3602,N_3705);
or U3860 (N_3860,N_3716,N_3713);
and U3861 (N_3861,N_3715,N_3609);
and U3862 (N_3862,N_3703,N_3660);
and U3863 (N_3863,N_3618,N_3727);
xor U3864 (N_3864,N_3714,N_3707);
nor U3865 (N_3865,N_3676,N_3679);
nand U3866 (N_3866,N_3724,N_3726);
and U3867 (N_3867,N_3721,N_3673);
and U3868 (N_3868,N_3679,N_3675);
or U3869 (N_3869,N_3673,N_3702);
nor U3870 (N_3870,N_3635,N_3672);
or U3871 (N_3871,N_3659,N_3639);
or U3872 (N_3872,N_3635,N_3673);
nor U3873 (N_3873,N_3641,N_3658);
nor U3874 (N_3874,N_3635,N_3718);
and U3875 (N_3875,N_3661,N_3631);
xnor U3876 (N_3876,N_3665,N_3748);
and U3877 (N_3877,N_3640,N_3611);
and U3878 (N_3878,N_3616,N_3633);
nor U3879 (N_3879,N_3641,N_3718);
nand U3880 (N_3880,N_3710,N_3697);
xnor U3881 (N_3881,N_3618,N_3658);
nor U3882 (N_3882,N_3654,N_3733);
or U3883 (N_3883,N_3741,N_3745);
nand U3884 (N_3884,N_3726,N_3634);
or U3885 (N_3885,N_3634,N_3708);
xor U3886 (N_3886,N_3717,N_3715);
xor U3887 (N_3887,N_3642,N_3617);
xnor U3888 (N_3888,N_3666,N_3610);
nor U3889 (N_3889,N_3672,N_3663);
and U3890 (N_3890,N_3630,N_3736);
nor U3891 (N_3891,N_3659,N_3705);
nand U3892 (N_3892,N_3706,N_3650);
xnor U3893 (N_3893,N_3744,N_3667);
nand U3894 (N_3894,N_3610,N_3730);
and U3895 (N_3895,N_3740,N_3622);
or U3896 (N_3896,N_3746,N_3671);
nor U3897 (N_3897,N_3649,N_3718);
and U3898 (N_3898,N_3638,N_3723);
or U3899 (N_3899,N_3614,N_3652);
nor U3900 (N_3900,N_3793,N_3857);
xnor U3901 (N_3901,N_3822,N_3883);
nor U3902 (N_3902,N_3758,N_3898);
and U3903 (N_3903,N_3808,N_3866);
or U3904 (N_3904,N_3761,N_3787);
or U3905 (N_3905,N_3868,N_3786);
nand U3906 (N_3906,N_3755,N_3897);
or U3907 (N_3907,N_3794,N_3893);
and U3908 (N_3908,N_3819,N_3825);
or U3909 (N_3909,N_3899,N_3885);
nand U3910 (N_3910,N_3867,N_3790);
nor U3911 (N_3911,N_3849,N_3775);
nor U3912 (N_3912,N_3799,N_3778);
xnor U3913 (N_3913,N_3768,N_3835);
nand U3914 (N_3914,N_3862,N_3880);
xnor U3915 (N_3915,N_3788,N_3792);
or U3916 (N_3916,N_3896,N_3865);
xor U3917 (N_3917,N_3826,N_3895);
xnor U3918 (N_3918,N_3784,N_3751);
and U3919 (N_3919,N_3800,N_3884);
or U3920 (N_3920,N_3860,N_3797);
xnor U3921 (N_3921,N_3873,N_3767);
nand U3922 (N_3922,N_3765,N_3769);
and U3923 (N_3923,N_3839,N_3887);
nand U3924 (N_3924,N_3891,N_3756);
and U3925 (N_3925,N_3806,N_3757);
nor U3926 (N_3926,N_3877,N_3779);
and U3927 (N_3927,N_3856,N_3759);
and U3928 (N_3928,N_3843,N_3871);
nor U3929 (N_3929,N_3801,N_3760);
xor U3930 (N_3930,N_3804,N_3753);
nand U3931 (N_3931,N_3850,N_3782);
nand U3932 (N_3932,N_3817,N_3879);
and U3933 (N_3933,N_3878,N_3805);
xnor U3934 (N_3934,N_3776,N_3771);
and U3935 (N_3935,N_3859,N_3861);
nand U3936 (N_3936,N_3803,N_3831);
or U3937 (N_3937,N_3837,N_3763);
or U3938 (N_3938,N_3858,N_3762);
and U3939 (N_3939,N_3876,N_3841);
xor U3940 (N_3940,N_3844,N_3874);
nand U3941 (N_3941,N_3802,N_3882);
or U3942 (N_3942,N_3824,N_3845);
nand U3943 (N_3943,N_3796,N_3846);
nand U3944 (N_3944,N_3812,N_3811);
or U3945 (N_3945,N_3870,N_3892);
and U3946 (N_3946,N_3886,N_3823);
and U3947 (N_3947,N_3814,N_3783);
xnor U3948 (N_3948,N_3863,N_3789);
nor U3949 (N_3949,N_3752,N_3832);
nor U3950 (N_3950,N_3872,N_3773);
nand U3951 (N_3951,N_3777,N_3809);
nand U3952 (N_3952,N_3798,N_3816);
nand U3953 (N_3953,N_3869,N_3847);
xor U3954 (N_3954,N_3772,N_3795);
xor U3955 (N_3955,N_3855,N_3854);
or U3956 (N_3956,N_3791,N_3894);
nand U3957 (N_3957,N_3770,N_3766);
nor U3958 (N_3958,N_3780,N_3827);
or U3959 (N_3959,N_3807,N_3853);
and U3960 (N_3960,N_3852,N_3813);
nand U3961 (N_3961,N_3851,N_3820);
nand U3962 (N_3962,N_3810,N_3818);
nand U3963 (N_3963,N_3875,N_3834);
and U3964 (N_3964,N_3815,N_3848);
or U3965 (N_3965,N_3785,N_3830);
nor U3966 (N_3966,N_3829,N_3750);
or U3967 (N_3967,N_3889,N_3842);
or U3968 (N_3968,N_3781,N_3838);
nor U3969 (N_3969,N_3840,N_3833);
nand U3970 (N_3970,N_3774,N_3890);
nand U3971 (N_3971,N_3764,N_3881);
xor U3972 (N_3972,N_3754,N_3864);
xor U3973 (N_3973,N_3888,N_3836);
nor U3974 (N_3974,N_3821,N_3828);
nand U3975 (N_3975,N_3767,N_3882);
xor U3976 (N_3976,N_3789,N_3857);
nand U3977 (N_3977,N_3834,N_3802);
nor U3978 (N_3978,N_3830,N_3804);
or U3979 (N_3979,N_3796,N_3813);
nor U3980 (N_3980,N_3862,N_3829);
nor U3981 (N_3981,N_3752,N_3889);
nand U3982 (N_3982,N_3777,N_3817);
and U3983 (N_3983,N_3898,N_3760);
nor U3984 (N_3984,N_3860,N_3863);
xor U3985 (N_3985,N_3815,N_3762);
nor U3986 (N_3986,N_3890,N_3782);
or U3987 (N_3987,N_3798,N_3776);
xor U3988 (N_3988,N_3787,N_3829);
xnor U3989 (N_3989,N_3788,N_3779);
xor U3990 (N_3990,N_3844,N_3836);
xor U3991 (N_3991,N_3812,N_3830);
nand U3992 (N_3992,N_3758,N_3790);
and U3993 (N_3993,N_3851,N_3761);
and U3994 (N_3994,N_3876,N_3758);
nor U3995 (N_3995,N_3783,N_3823);
xor U3996 (N_3996,N_3795,N_3874);
and U3997 (N_3997,N_3760,N_3851);
nor U3998 (N_3998,N_3832,N_3808);
nor U3999 (N_3999,N_3802,N_3849);
or U4000 (N_4000,N_3815,N_3764);
nor U4001 (N_4001,N_3784,N_3793);
nand U4002 (N_4002,N_3841,N_3862);
nor U4003 (N_4003,N_3867,N_3795);
nand U4004 (N_4004,N_3780,N_3846);
or U4005 (N_4005,N_3759,N_3889);
xor U4006 (N_4006,N_3806,N_3783);
xnor U4007 (N_4007,N_3780,N_3838);
and U4008 (N_4008,N_3763,N_3859);
or U4009 (N_4009,N_3793,N_3800);
and U4010 (N_4010,N_3793,N_3794);
and U4011 (N_4011,N_3834,N_3884);
nor U4012 (N_4012,N_3870,N_3875);
or U4013 (N_4013,N_3842,N_3792);
nor U4014 (N_4014,N_3816,N_3796);
nor U4015 (N_4015,N_3886,N_3845);
or U4016 (N_4016,N_3874,N_3876);
nand U4017 (N_4017,N_3815,N_3867);
nor U4018 (N_4018,N_3899,N_3750);
xor U4019 (N_4019,N_3764,N_3756);
xor U4020 (N_4020,N_3831,N_3897);
or U4021 (N_4021,N_3847,N_3895);
and U4022 (N_4022,N_3844,N_3777);
nor U4023 (N_4023,N_3794,N_3813);
or U4024 (N_4024,N_3847,N_3892);
xnor U4025 (N_4025,N_3760,N_3765);
or U4026 (N_4026,N_3803,N_3752);
and U4027 (N_4027,N_3877,N_3808);
and U4028 (N_4028,N_3814,N_3863);
nor U4029 (N_4029,N_3759,N_3773);
and U4030 (N_4030,N_3885,N_3809);
and U4031 (N_4031,N_3838,N_3811);
nor U4032 (N_4032,N_3859,N_3761);
xor U4033 (N_4033,N_3837,N_3830);
or U4034 (N_4034,N_3759,N_3819);
xor U4035 (N_4035,N_3859,N_3849);
nor U4036 (N_4036,N_3847,N_3891);
or U4037 (N_4037,N_3810,N_3808);
and U4038 (N_4038,N_3831,N_3801);
nand U4039 (N_4039,N_3893,N_3766);
and U4040 (N_4040,N_3859,N_3827);
nand U4041 (N_4041,N_3759,N_3836);
nor U4042 (N_4042,N_3758,N_3777);
nand U4043 (N_4043,N_3776,N_3784);
nand U4044 (N_4044,N_3860,N_3835);
xnor U4045 (N_4045,N_3868,N_3765);
and U4046 (N_4046,N_3883,N_3815);
nor U4047 (N_4047,N_3813,N_3863);
and U4048 (N_4048,N_3784,N_3765);
nor U4049 (N_4049,N_3887,N_3824);
nor U4050 (N_4050,N_3947,N_3909);
and U4051 (N_4051,N_3994,N_3925);
nand U4052 (N_4052,N_3923,N_3977);
or U4053 (N_4053,N_3942,N_3971);
xnor U4054 (N_4054,N_3902,N_4017);
xor U4055 (N_4055,N_3970,N_3935);
nor U4056 (N_4056,N_3991,N_3975);
or U4057 (N_4057,N_4018,N_4022);
and U4058 (N_4058,N_4006,N_4048);
nor U4059 (N_4059,N_3905,N_4001);
and U4060 (N_4060,N_4003,N_3950);
or U4061 (N_4061,N_3912,N_3922);
and U4062 (N_4062,N_4012,N_3965);
nand U4063 (N_4063,N_3963,N_3946);
nand U4064 (N_4064,N_3939,N_4008);
xor U4065 (N_4065,N_4047,N_3998);
or U4066 (N_4066,N_3957,N_4016);
nand U4067 (N_4067,N_4023,N_3927);
xor U4068 (N_4068,N_4034,N_3936);
or U4069 (N_4069,N_4004,N_4030);
xor U4070 (N_4070,N_3982,N_3937);
and U4071 (N_4071,N_4041,N_3916);
nand U4072 (N_4072,N_4042,N_3926);
and U4073 (N_4073,N_4045,N_4040);
xnor U4074 (N_4074,N_3969,N_3979);
nor U4075 (N_4075,N_3958,N_3906);
and U4076 (N_4076,N_3949,N_4020);
xor U4077 (N_4077,N_4002,N_3938);
or U4078 (N_4078,N_4026,N_3934);
and U4079 (N_4079,N_3993,N_3904);
xnor U4080 (N_4080,N_4044,N_3917);
nor U4081 (N_4081,N_3953,N_4021);
nor U4082 (N_4082,N_3992,N_3951);
nor U4083 (N_4083,N_4035,N_4024);
xor U4084 (N_4084,N_3995,N_4027);
nor U4085 (N_4085,N_3972,N_3929);
nand U4086 (N_4086,N_4029,N_3983);
nor U4087 (N_4087,N_3945,N_3908);
xor U4088 (N_4088,N_3997,N_4014);
xnor U4089 (N_4089,N_3985,N_3964);
nand U4090 (N_4090,N_3932,N_3940);
nand U4091 (N_4091,N_3941,N_4005);
or U4092 (N_4092,N_3943,N_3907);
or U4093 (N_4093,N_4038,N_3903);
nor U4094 (N_4094,N_3999,N_4011);
or U4095 (N_4095,N_3980,N_4046);
and U4096 (N_4096,N_4019,N_3901);
or U4097 (N_4097,N_4036,N_4031);
and U4098 (N_4098,N_4028,N_3955);
xnor U4099 (N_4099,N_3910,N_3959);
or U4100 (N_4100,N_3984,N_3933);
or U4101 (N_4101,N_3948,N_3973);
or U4102 (N_4102,N_3962,N_3968);
and U4103 (N_4103,N_3988,N_4000);
nand U4104 (N_4104,N_3990,N_4009);
nor U4105 (N_4105,N_4015,N_3928);
nand U4106 (N_4106,N_4039,N_3961);
and U4107 (N_4107,N_3921,N_3919);
nor U4108 (N_4108,N_3924,N_4043);
nand U4109 (N_4109,N_3976,N_3986);
or U4110 (N_4110,N_4013,N_4007);
or U4111 (N_4111,N_3900,N_3944);
nand U4112 (N_4112,N_3954,N_3974);
nor U4113 (N_4113,N_3967,N_3960);
and U4114 (N_4114,N_4033,N_3978);
or U4115 (N_4115,N_3914,N_3981);
nor U4116 (N_4116,N_3930,N_3996);
and U4117 (N_4117,N_3920,N_3918);
and U4118 (N_4118,N_3913,N_3915);
and U4119 (N_4119,N_3956,N_4010);
nor U4120 (N_4120,N_3989,N_4037);
and U4121 (N_4121,N_4049,N_3911);
nor U4122 (N_4122,N_3987,N_4032);
and U4123 (N_4123,N_3966,N_3931);
and U4124 (N_4124,N_3952,N_4025);
xnor U4125 (N_4125,N_3907,N_4014);
nand U4126 (N_4126,N_3956,N_3955);
and U4127 (N_4127,N_3951,N_4015);
or U4128 (N_4128,N_3928,N_4030);
xor U4129 (N_4129,N_3946,N_3932);
nand U4130 (N_4130,N_4022,N_3968);
nor U4131 (N_4131,N_3981,N_4041);
nand U4132 (N_4132,N_3984,N_4021);
and U4133 (N_4133,N_3994,N_3917);
and U4134 (N_4134,N_3928,N_3988);
nor U4135 (N_4135,N_3928,N_3900);
and U4136 (N_4136,N_3912,N_4022);
nor U4137 (N_4137,N_3962,N_3955);
and U4138 (N_4138,N_3958,N_3983);
xnor U4139 (N_4139,N_4006,N_4029);
or U4140 (N_4140,N_3903,N_3986);
xor U4141 (N_4141,N_3961,N_4025);
xnor U4142 (N_4142,N_3930,N_3954);
nand U4143 (N_4143,N_3938,N_3976);
or U4144 (N_4144,N_4033,N_4049);
nand U4145 (N_4145,N_4040,N_4005);
or U4146 (N_4146,N_4001,N_3901);
nor U4147 (N_4147,N_3928,N_3914);
nor U4148 (N_4148,N_4044,N_3992);
nor U4149 (N_4149,N_3915,N_3907);
xnor U4150 (N_4150,N_3901,N_4004);
and U4151 (N_4151,N_3917,N_4007);
xor U4152 (N_4152,N_4009,N_3984);
or U4153 (N_4153,N_3935,N_3953);
xnor U4154 (N_4154,N_3920,N_4005);
or U4155 (N_4155,N_3997,N_3902);
nand U4156 (N_4156,N_3925,N_3976);
xnor U4157 (N_4157,N_4027,N_4045);
nand U4158 (N_4158,N_3954,N_4025);
nand U4159 (N_4159,N_3965,N_3948);
or U4160 (N_4160,N_4036,N_3972);
nand U4161 (N_4161,N_4014,N_3957);
nand U4162 (N_4162,N_3970,N_4024);
and U4163 (N_4163,N_3940,N_3909);
nand U4164 (N_4164,N_3931,N_3936);
xnor U4165 (N_4165,N_3984,N_4041);
and U4166 (N_4166,N_3971,N_4037);
nor U4167 (N_4167,N_4028,N_4047);
nand U4168 (N_4168,N_3996,N_3978);
or U4169 (N_4169,N_4036,N_3926);
nor U4170 (N_4170,N_3919,N_4043);
xnor U4171 (N_4171,N_4035,N_3950);
nor U4172 (N_4172,N_3935,N_3915);
nor U4173 (N_4173,N_3932,N_4015);
nand U4174 (N_4174,N_3941,N_3913);
and U4175 (N_4175,N_4044,N_4009);
nor U4176 (N_4176,N_3971,N_4045);
or U4177 (N_4177,N_3923,N_3940);
nand U4178 (N_4178,N_4028,N_4042);
nand U4179 (N_4179,N_3989,N_4046);
and U4180 (N_4180,N_3993,N_3980);
or U4181 (N_4181,N_3929,N_3995);
nand U4182 (N_4182,N_3972,N_4045);
or U4183 (N_4183,N_4031,N_3925);
nor U4184 (N_4184,N_3976,N_3942);
and U4185 (N_4185,N_3982,N_4019);
xor U4186 (N_4186,N_3930,N_4034);
and U4187 (N_4187,N_3933,N_3903);
or U4188 (N_4188,N_4048,N_4040);
and U4189 (N_4189,N_3935,N_3902);
nand U4190 (N_4190,N_3942,N_3907);
xor U4191 (N_4191,N_3919,N_3970);
nor U4192 (N_4192,N_3985,N_4024);
and U4193 (N_4193,N_3934,N_3907);
xnor U4194 (N_4194,N_4036,N_4049);
nor U4195 (N_4195,N_3976,N_3933);
or U4196 (N_4196,N_3984,N_4011);
nor U4197 (N_4197,N_3982,N_3985);
xnor U4198 (N_4198,N_3939,N_3947);
nor U4199 (N_4199,N_3918,N_3922);
or U4200 (N_4200,N_4193,N_4093);
or U4201 (N_4201,N_4075,N_4092);
and U4202 (N_4202,N_4157,N_4172);
or U4203 (N_4203,N_4082,N_4171);
nor U4204 (N_4204,N_4123,N_4133);
xnor U4205 (N_4205,N_4154,N_4135);
or U4206 (N_4206,N_4168,N_4127);
nand U4207 (N_4207,N_4177,N_4083);
xnor U4208 (N_4208,N_4118,N_4152);
xnor U4209 (N_4209,N_4132,N_4078);
and U4210 (N_4210,N_4179,N_4189);
nand U4211 (N_4211,N_4130,N_4164);
nor U4212 (N_4212,N_4180,N_4141);
nor U4213 (N_4213,N_4151,N_4125);
nand U4214 (N_4214,N_4073,N_4117);
or U4215 (N_4215,N_4190,N_4086);
nand U4216 (N_4216,N_4158,N_4116);
nand U4217 (N_4217,N_4070,N_4150);
nand U4218 (N_4218,N_4120,N_4091);
xor U4219 (N_4219,N_4145,N_4050);
nand U4220 (N_4220,N_4143,N_4183);
nor U4221 (N_4221,N_4098,N_4079);
or U4222 (N_4222,N_4191,N_4119);
xnor U4223 (N_4223,N_4069,N_4066);
or U4224 (N_4224,N_4174,N_4065);
and U4225 (N_4225,N_4140,N_4194);
nand U4226 (N_4226,N_4192,N_4068);
or U4227 (N_4227,N_4060,N_4095);
or U4228 (N_4228,N_4181,N_4109);
nor U4229 (N_4229,N_4102,N_4188);
nand U4230 (N_4230,N_4111,N_4090);
and U4231 (N_4231,N_4103,N_4175);
or U4232 (N_4232,N_4182,N_4122);
and U4233 (N_4233,N_4121,N_4162);
or U4234 (N_4234,N_4055,N_4147);
nand U4235 (N_4235,N_4063,N_4056);
or U4236 (N_4236,N_4074,N_4161);
and U4237 (N_4237,N_4081,N_4131);
xor U4238 (N_4238,N_4061,N_4053);
nand U4239 (N_4239,N_4088,N_4195);
xor U4240 (N_4240,N_4072,N_4185);
nor U4241 (N_4241,N_4051,N_4169);
nor U4242 (N_4242,N_4197,N_4139);
and U4243 (N_4243,N_4176,N_4144);
or U4244 (N_4244,N_4080,N_4062);
and U4245 (N_4245,N_4128,N_4097);
xnor U4246 (N_4246,N_4084,N_4108);
xnor U4247 (N_4247,N_4054,N_4166);
or U4248 (N_4248,N_4187,N_4129);
nand U4249 (N_4249,N_4134,N_4057);
nor U4250 (N_4250,N_4178,N_4160);
nand U4251 (N_4251,N_4124,N_4085);
xnor U4252 (N_4252,N_4155,N_4126);
nand U4253 (N_4253,N_4142,N_4058);
or U4254 (N_4254,N_4067,N_4099);
nor U4255 (N_4255,N_4184,N_4159);
nor U4256 (N_4256,N_4115,N_4105);
nor U4257 (N_4257,N_4146,N_4167);
nor U4258 (N_4258,N_4163,N_4052);
and U4259 (N_4259,N_4138,N_4064);
and U4260 (N_4260,N_4136,N_4071);
nand U4261 (N_4261,N_4096,N_4100);
xor U4262 (N_4262,N_4107,N_4077);
nor U4263 (N_4263,N_4199,N_4196);
or U4264 (N_4264,N_4089,N_4087);
and U4265 (N_4265,N_4165,N_4112);
xnor U4266 (N_4266,N_4149,N_4076);
nand U4267 (N_4267,N_4101,N_4186);
nor U4268 (N_4268,N_4153,N_4106);
or U4269 (N_4269,N_4173,N_4110);
nand U4270 (N_4270,N_4156,N_4170);
nor U4271 (N_4271,N_4113,N_4104);
or U4272 (N_4272,N_4114,N_4094);
nand U4273 (N_4273,N_4059,N_4137);
xnor U4274 (N_4274,N_4198,N_4148);
xnor U4275 (N_4275,N_4158,N_4162);
and U4276 (N_4276,N_4151,N_4183);
nand U4277 (N_4277,N_4070,N_4132);
or U4278 (N_4278,N_4185,N_4070);
and U4279 (N_4279,N_4195,N_4183);
xnor U4280 (N_4280,N_4175,N_4050);
nand U4281 (N_4281,N_4152,N_4194);
nand U4282 (N_4282,N_4117,N_4174);
and U4283 (N_4283,N_4158,N_4131);
or U4284 (N_4284,N_4058,N_4084);
or U4285 (N_4285,N_4182,N_4147);
xor U4286 (N_4286,N_4106,N_4112);
nand U4287 (N_4287,N_4133,N_4073);
or U4288 (N_4288,N_4063,N_4082);
nor U4289 (N_4289,N_4164,N_4117);
and U4290 (N_4290,N_4064,N_4198);
nor U4291 (N_4291,N_4116,N_4148);
nand U4292 (N_4292,N_4109,N_4175);
or U4293 (N_4293,N_4065,N_4177);
and U4294 (N_4294,N_4069,N_4115);
nor U4295 (N_4295,N_4100,N_4194);
xnor U4296 (N_4296,N_4123,N_4196);
xor U4297 (N_4297,N_4127,N_4155);
nor U4298 (N_4298,N_4148,N_4137);
nand U4299 (N_4299,N_4158,N_4167);
nand U4300 (N_4300,N_4064,N_4162);
xor U4301 (N_4301,N_4159,N_4134);
nand U4302 (N_4302,N_4118,N_4092);
and U4303 (N_4303,N_4123,N_4163);
nand U4304 (N_4304,N_4087,N_4186);
xor U4305 (N_4305,N_4083,N_4180);
xnor U4306 (N_4306,N_4151,N_4051);
or U4307 (N_4307,N_4168,N_4126);
nand U4308 (N_4308,N_4100,N_4189);
and U4309 (N_4309,N_4192,N_4054);
nor U4310 (N_4310,N_4104,N_4128);
and U4311 (N_4311,N_4065,N_4064);
or U4312 (N_4312,N_4147,N_4080);
or U4313 (N_4313,N_4063,N_4171);
nor U4314 (N_4314,N_4073,N_4061);
and U4315 (N_4315,N_4097,N_4197);
xnor U4316 (N_4316,N_4149,N_4111);
or U4317 (N_4317,N_4110,N_4054);
nand U4318 (N_4318,N_4199,N_4178);
nand U4319 (N_4319,N_4149,N_4082);
or U4320 (N_4320,N_4060,N_4068);
or U4321 (N_4321,N_4168,N_4199);
nand U4322 (N_4322,N_4186,N_4137);
nor U4323 (N_4323,N_4179,N_4190);
and U4324 (N_4324,N_4133,N_4137);
and U4325 (N_4325,N_4153,N_4085);
nor U4326 (N_4326,N_4072,N_4093);
nor U4327 (N_4327,N_4097,N_4194);
or U4328 (N_4328,N_4088,N_4186);
or U4329 (N_4329,N_4067,N_4085);
nor U4330 (N_4330,N_4187,N_4143);
nor U4331 (N_4331,N_4118,N_4124);
xnor U4332 (N_4332,N_4120,N_4097);
or U4333 (N_4333,N_4094,N_4184);
nand U4334 (N_4334,N_4176,N_4157);
nand U4335 (N_4335,N_4176,N_4187);
xnor U4336 (N_4336,N_4084,N_4177);
and U4337 (N_4337,N_4165,N_4053);
xnor U4338 (N_4338,N_4058,N_4104);
and U4339 (N_4339,N_4056,N_4115);
and U4340 (N_4340,N_4137,N_4150);
xor U4341 (N_4341,N_4092,N_4158);
xnor U4342 (N_4342,N_4192,N_4076);
nand U4343 (N_4343,N_4197,N_4056);
or U4344 (N_4344,N_4183,N_4164);
xnor U4345 (N_4345,N_4145,N_4068);
nor U4346 (N_4346,N_4083,N_4141);
and U4347 (N_4347,N_4099,N_4103);
or U4348 (N_4348,N_4083,N_4098);
xor U4349 (N_4349,N_4165,N_4070);
and U4350 (N_4350,N_4251,N_4298);
xnor U4351 (N_4351,N_4202,N_4214);
and U4352 (N_4352,N_4256,N_4280);
nor U4353 (N_4353,N_4286,N_4334);
nor U4354 (N_4354,N_4246,N_4331);
and U4355 (N_4355,N_4259,N_4215);
or U4356 (N_4356,N_4294,N_4221);
nand U4357 (N_4357,N_4348,N_4243);
nand U4358 (N_4358,N_4233,N_4349);
nand U4359 (N_4359,N_4289,N_4278);
nor U4360 (N_4360,N_4228,N_4307);
and U4361 (N_4361,N_4328,N_4212);
xor U4362 (N_4362,N_4231,N_4264);
and U4363 (N_4363,N_4238,N_4338);
or U4364 (N_4364,N_4330,N_4325);
nand U4365 (N_4365,N_4222,N_4271);
and U4366 (N_4366,N_4322,N_4345);
nor U4367 (N_4367,N_4227,N_4300);
xor U4368 (N_4368,N_4290,N_4230);
nand U4369 (N_4369,N_4200,N_4323);
nor U4370 (N_4370,N_4210,N_4255);
xnor U4371 (N_4371,N_4253,N_4275);
nor U4372 (N_4372,N_4213,N_4287);
or U4373 (N_4373,N_4269,N_4288);
or U4374 (N_4374,N_4292,N_4297);
or U4375 (N_4375,N_4232,N_4225);
or U4376 (N_4376,N_4262,N_4314);
or U4377 (N_4377,N_4299,N_4240);
nand U4378 (N_4378,N_4235,N_4295);
xor U4379 (N_4379,N_4320,N_4205);
nand U4380 (N_4380,N_4250,N_4335);
and U4381 (N_4381,N_4241,N_4234);
nor U4382 (N_4382,N_4284,N_4267);
or U4383 (N_4383,N_4301,N_4327);
xnor U4384 (N_4384,N_4317,N_4333);
or U4385 (N_4385,N_4293,N_4344);
nor U4386 (N_4386,N_4305,N_4310);
and U4387 (N_4387,N_4265,N_4216);
xor U4388 (N_4388,N_4260,N_4272);
nor U4389 (N_4389,N_4340,N_4203);
xnor U4390 (N_4390,N_4343,N_4220);
xor U4391 (N_4391,N_4311,N_4326);
or U4392 (N_4392,N_4204,N_4341);
nor U4393 (N_4393,N_4291,N_4211);
nand U4394 (N_4394,N_4342,N_4242);
nor U4395 (N_4395,N_4270,N_4226);
xor U4396 (N_4396,N_4223,N_4324);
nand U4397 (N_4397,N_4347,N_4249);
or U4398 (N_4398,N_4277,N_4304);
nand U4399 (N_4399,N_4303,N_4337);
nand U4400 (N_4400,N_4279,N_4257);
or U4401 (N_4401,N_4296,N_4261);
xor U4402 (N_4402,N_4208,N_4254);
and U4403 (N_4403,N_4285,N_4329);
or U4404 (N_4404,N_4302,N_4319);
and U4405 (N_4405,N_4206,N_4339);
and U4406 (N_4406,N_4244,N_4224);
and U4407 (N_4407,N_4252,N_4312);
nand U4408 (N_4408,N_4306,N_4273);
nand U4409 (N_4409,N_4321,N_4318);
nand U4410 (N_4410,N_4217,N_4316);
and U4411 (N_4411,N_4283,N_4309);
or U4412 (N_4412,N_4276,N_4207);
and U4413 (N_4413,N_4245,N_4218);
nand U4414 (N_4414,N_4268,N_4274);
or U4415 (N_4415,N_4308,N_4209);
xor U4416 (N_4416,N_4236,N_4315);
nor U4417 (N_4417,N_4201,N_4266);
xor U4418 (N_4418,N_4282,N_4248);
nand U4419 (N_4419,N_4313,N_4229);
xor U4420 (N_4420,N_4239,N_4237);
nor U4421 (N_4421,N_4263,N_4336);
nor U4422 (N_4422,N_4258,N_4332);
xnor U4423 (N_4423,N_4219,N_4346);
or U4424 (N_4424,N_4247,N_4281);
nand U4425 (N_4425,N_4242,N_4250);
nand U4426 (N_4426,N_4320,N_4300);
xor U4427 (N_4427,N_4278,N_4261);
and U4428 (N_4428,N_4266,N_4295);
or U4429 (N_4429,N_4239,N_4202);
xor U4430 (N_4430,N_4257,N_4347);
nand U4431 (N_4431,N_4222,N_4300);
nor U4432 (N_4432,N_4239,N_4331);
or U4433 (N_4433,N_4304,N_4267);
or U4434 (N_4434,N_4298,N_4308);
or U4435 (N_4435,N_4209,N_4255);
nand U4436 (N_4436,N_4279,N_4329);
nor U4437 (N_4437,N_4273,N_4253);
and U4438 (N_4438,N_4232,N_4308);
nor U4439 (N_4439,N_4231,N_4259);
and U4440 (N_4440,N_4312,N_4310);
or U4441 (N_4441,N_4343,N_4245);
and U4442 (N_4442,N_4209,N_4302);
nor U4443 (N_4443,N_4279,N_4243);
and U4444 (N_4444,N_4295,N_4239);
nor U4445 (N_4445,N_4289,N_4214);
nand U4446 (N_4446,N_4340,N_4347);
or U4447 (N_4447,N_4278,N_4208);
nand U4448 (N_4448,N_4206,N_4201);
and U4449 (N_4449,N_4266,N_4321);
and U4450 (N_4450,N_4293,N_4229);
and U4451 (N_4451,N_4256,N_4303);
nand U4452 (N_4452,N_4319,N_4305);
xnor U4453 (N_4453,N_4209,N_4300);
and U4454 (N_4454,N_4278,N_4336);
nor U4455 (N_4455,N_4327,N_4285);
nor U4456 (N_4456,N_4291,N_4324);
and U4457 (N_4457,N_4348,N_4295);
or U4458 (N_4458,N_4289,N_4293);
xor U4459 (N_4459,N_4252,N_4349);
nor U4460 (N_4460,N_4278,N_4253);
nor U4461 (N_4461,N_4331,N_4247);
and U4462 (N_4462,N_4204,N_4217);
or U4463 (N_4463,N_4213,N_4314);
and U4464 (N_4464,N_4216,N_4248);
and U4465 (N_4465,N_4273,N_4332);
xor U4466 (N_4466,N_4302,N_4247);
nand U4467 (N_4467,N_4297,N_4242);
nand U4468 (N_4468,N_4293,N_4246);
nand U4469 (N_4469,N_4325,N_4293);
nor U4470 (N_4470,N_4283,N_4341);
xnor U4471 (N_4471,N_4279,N_4332);
and U4472 (N_4472,N_4232,N_4327);
xor U4473 (N_4473,N_4303,N_4246);
and U4474 (N_4474,N_4331,N_4343);
and U4475 (N_4475,N_4315,N_4342);
nor U4476 (N_4476,N_4273,N_4291);
and U4477 (N_4477,N_4200,N_4310);
and U4478 (N_4478,N_4216,N_4241);
and U4479 (N_4479,N_4239,N_4245);
and U4480 (N_4480,N_4230,N_4213);
xnor U4481 (N_4481,N_4271,N_4246);
xnor U4482 (N_4482,N_4276,N_4294);
and U4483 (N_4483,N_4213,N_4316);
nor U4484 (N_4484,N_4279,N_4242);
and U4485 (N_4485,N_4324,N_4277);
nand U4486 (N_4486,N_4318,N_4313);
xor U4487 (N_4487,N_4263,N_4272);
nand U4488 (N_4488,N_4317,N_4233);
nor U4489 (N_4489,N_4247,N_4330);
and U4490 (N_4490,N_4279,N_4216);
and U4491 (N_4491,N_4302,N_4282);
nand U4492 (N_4492,N_4226,N_4342);
nand U4493 (N_4493,N_4277,N_4206);
and U4494 (N_4494,N_4286,N_4320);
xnor U4495 (N_4495,N_4304,N_4264);
and U4496 (N_4496,N_4250,N_4229);
nand U4497 (N_4497,N_4302,N_4345);
nand U4498 (N_4498,N_4267,N_4237);
or U4499 (N_4499,N_4242,N_4240);
nor U4500 (N_4500,N_4421,N_4367);
and U4501 (N_4501,N_4375,N_4453);
nor U4502 (N_4502,N_4420,N_4378);
xnor U4503 (N_4503,N_4483,N_4432);
nor U4504 (N_4504,N_4406,N_4393);
nor U4505 (N_4505,N_4369,N_4429);
or U4506 (N_4506,N_4419,N_4492);
nand U4507 (N_4507,N_4400,N_4407);
nor U4508 (N_4508,N_4449,N_4499);
nand U4509 (N_4509,N_4409,N_4403);
nand U4510 (N_4510,N_4477,N_4436);
or U4511 (N_4511,N_4490,N_4451);
nor U4512 (N_4512,N_4374,N_4404);
nand U4513 (N_4513,N_4356,N_4416);
and U4514 (N_4514,N_4484,N_4379);
nand U4515 (N_4515,N_4445,N_4359);
nor U4516 (N_4516,N_4458,N_4351);
or U4517 (N_4517,N_4468,N_4464);
xnor U4518 (N_4518,N_4385,N_4396);
or U4519 (N_4519,N_4399,N_4497);
nor U4520 (N_4520,N_4434,N_4493);
and U4521 (N_4521,N_4370,N_4461);
xor U4522 (N_4522,N_4414,N_4474);
and U4523 (N_4523,N_4422,N_4470);
or U4524 (N_4524,N_4485,N_4450);
xor U4525 (N_4525,N_4427,N_4465);
and U4526 (N_4526,N_4352,N_4439);
nand U4527 (N_4527,N_4447,N_4415);
nor U4528 (N_4528,N_4428,N_4491);
nand U4529 (N_4529,N_4394,N_4452);
nor U4530 (N_4530,N_4486,N_4489);
or U4531 (N_4531,N_4395,N_4357);
nand U4532 (N_4532,N_4408,N_4362);
nand U4533 (N_4533,N_4381,N_4411);
and U4534 (N_4534,N_4469,N_4397);
nor U4535 (N_4535,N_4425,N_4361);
and U4536 (N_4536,N_4457,N_4388);
xor U4537 (N_4537,N_4460,N_4437);
and U4538 (N_4538,N_4401,N_4467);
nand U4539 (N_4539,N_4478,N_4480);
or U4540 (N_4540,N_4417,N_4424);
or U4541 (N_4541,N_4440,N_4372);
or U4542 (N_4542,N_4373,N_4456);
xnor U4543 (N_4543,N_4444,N_4472);
xnor U4544 (N_4544,N_4398,N_4368);
xor U4545 (N_4545,N_4441,N_4380);
nor U4546 (N_4546,N_4471,N_4389);
xor U4547 (N_4547,N_4423,N_4353);
or U4548 (N_4548,N_4387,N_4402);
xnor U4549 (N_4549,N_4496,N_4476);
or U4550 (N_4550,N_4355,N_4482);
and U4551 (N_4551,N_4390,N_4405);
nor U4552 (N_4552,N_4454,N_4443);
or U4553 (N_4553,N_4376,N_4494);
or U4554 (N_4554,N_4358,N_4366);
nand U4555 (N_4555,N_4455,N_4413);
xnor U4556 (N_4556,N_4383,N_4364);
and U4557 (N_4557,N_4495,N_4412);
nand U4558 (N_4558,N_4410,N_4365);
nor U4559 (N_4559,N_4462,N_4426);
nand U4560 (N_4560,N_4430,N_4463);
and U4561 (N_4561,N_4488,N_4446);
and U4562 (N_4562,N_4431,N_4386);
nor U4563 (N_4563,N_4391,N_4487);
nor U4564 (N_4564,N_4479,N_4438);
or U4565 (N_4565,N_4466,N_4354);
or U4566 (N_4566,N_4377,N_4433);
xnor U4567 (N_4567,N_4360,N_4498);
xor U4568 (N_4568,N_4350,N_4442);
and U4569 (N_4569,N_4392,N_4384);
or U4570 (N_4570,N_4475,N_4448);
nand U4571 (N_4571,N_4382,N_4459);
nand U4572 (N_4572,N_4371,N_4473);
nand U4573 (N_4573,N_4363,N_4435);
or U4574 (N_4574,N_4418,N_4481);
xor U4575 (N_4575,N_4393,N_4398);
nor U4576 (N_4576,N_4354,N_4404);
xnor U4577 (N_4577,N_4447,N_4434);
nor U4578 (N_4578,N_4437,N_4388);
xnor U4579 (N_4579,N_4428,N_4373);
nor U4580 (N_4580,N_4416,N_4473);
or U4581 (N_4581,N_4434,N_4454);
nor U4582 (N_4582,N_4364,N_4480);
and U4583 (N_4583,N_4391,N_4447);
nand U4584 (N_4584,N_4421,N_4452);
nand U4585 (N_4585,N_4401,N_4379);
nor U4586 (N_4586,N_4438,N_4397);
and U4587 (N_4587,N_4419,N_4493);
nand U4588 (N_4588,N_4354,N_4385);
or U4589 (N_4589,N_4382,N_4383);
or U4590 (N_4590,N_4412,N_4449);
or U4591 (N_4591,N_4410,N_4490);
and U4592 (N_4592,N_4414,N_4478);
or U4593 (N_4593,N_4453,N_4364);
nor U4594 (N_4594,N_4417,N_4453);
nand U4595 (N_4595,N_4483,N_4379);
xnor U4596 (N_4596,N_4435,N_4356);
nand U4597 (N_4597,N_4483,N_4413);
nand U4598 (N_4598,N_4410,N_4493);
xnor U4599 (N_4599,N_4446,N_4368);
nand U4600 (N_4600,N_4481,N_4442);
or U4601 (N_4601,N_4473,N_4495);
or U4602 (N_4602,N_4463,N_4449);
or U4603 (N_4603,N_4380,N_4474);
or U4604 (N_4604,N_4416,N_4392);
nor U4605 (N_4605,N_4438,N_4492);
and U4606 (N_4606,N_4469,N_4419);
xor U4607 (N_4607,N_4402,N_4428);
xor U4608 (N_4608,N_4390,N_4439);
or U4609 (N_4609,N_4430,N_4363);
and U4610 (N_4610,N_4460,N_4369);
xor U4611 (N_4611,N_4377,N_4470);
nand U4612 (N_4612,N_4393,N_4394);
and U4613 (N_4613,N_4411,N_4417);
nand U4614 (N_4614,N_4492,N_4432);
and U4615 (N_4615,N_4395,N_4458);
and U4616 (N_4616,N_4492,N_4441);
and U4617 (N_4617,N_4439,N_4489);
and U4618 (N_4618,N_4449,N_4382);
and U4619 (N_4619,N_4475,N_4409);
or U4620 (N_4620,N_4429,N_4434);
nand U4621 (N_4621,N_4441,N_4403);
xnor U4622 (N_4622,N_4366,N_4406);
xnor U4623 (N_4623,N_4373,N_4432);
and U4624 (N_4624,N_4376,N_4434);
nor U4625 (N_4625,N_4417,N_4448);
or U4626 (N_4626,N_4390,N_4381);
nor U4627 (N_4627,N_4433,N_4486);
nor U4628 (N_4628,N_4376,N_4370);
and U4629 (N_4629,N_4361,N_4455);
nor U4630 (N_4630,N_4429,N_4401);
xor U4631 (N_4631,N_4494,N_4402);
xnor U4632 (N_4632,N_4352,N_4375);
xor U4633 (N_4633,N_4468,N_4426);
or U4634 (N_4634,N_4482,N_4454);
and U4635 (N_4635,N_4406,N_4405);
xor U4636 (N_4636,N_4493,N_4476);
and U4637 (N_4637,N_4415,N_4369);
or U4638 (N_4638,N_4490,N_4400);
and U4639 (N_4639,N_4405,N_4413);
nand U4640 (N_4640,N_4412,N_4499);
or U4641 (N_4641,N_4421,N_4359);
nand U4642 (N_4642,N_4438,N_4488);
xnor U4643 (N_4643,N_4374,N_4368);
and U4644 (N_4644,N_4433,N_4387);
nor U4645 (N_4645,N_4461,N_4431);
nor U4646 (N_4646,N_4429,N_4441);
nand U4647 (N_4647,N_4428,N_4451);
nor U4648 (N_4648,N_4455,N_4405);
nand U4649 (N_4649,N_4395,N_4495);
or U4650 (N_4650,N_4558,N_4602);
or U4651 (N_4651,N_4632,N_4503);
and U4652 (N_4652,N_4633,N_4603);
nand U4653 (N_4653,N_4639,N_4548);
xnor U4654 (N_4654,N_4635,N_4581);
and U4655 (N_4655,N_4568,N_4502);
xnor U4656 (N_4656,N_4642,N_4580);
nor U4657 (N_4657,N_4544,N_4560);
nor U4658 (N_4658,N_4554,N_4509);
nand U4659 (N_4659,N_4647,N_4569);
nor U4660 (N_4660,N_4645,N_4611);
nor U4661 (N_4661,N_4621,N_4625);
nand U4662 (N_4662,N_4521,N_4643);
nor U4663 (N_4663,N_4616,N_4613);
nor U4664 (N_4664,N_4595,N_4592);
nand U4665 (N_4665,N_4529,N_4511);
nand U4666 (N_4666,N_4619,N_4517);
xnor U4667 (N_4667,N_4577,N_4598);
or U4668 (N_4668,N_4646,N_4505);
or U4669 (N_4669,N_4510,N_4593);
xor U4670 (N_4670,N_4518,N_4527);
and U4671 (N_4671,N_4586,N_4617);
and U4672 (N_4672,N_4584,N_4561);
nor U4673 (N_4673,N_4623,N_4629);
or U4674 (N_4674,N_4588,N_4530);
nand U4675 (N_4675,N_4612,N_4536);
xor U4676 (N_4676,N_4594,N_4501);
xor U4677 (N_4677,N_4547,N_4600);
nand U4678 (N_4678,N_4624,N_4615);
and U4679 (N_4679,N_4582,N_4535);
nand U4680 (N_4680,N_4513,N_4634);
nor U4681 (N_4681,N_4543,N_4608);
nor U4682 (N_4682,N_4553,N_4541);
and U4683 (N_4683,N_4609,N_4542);
nor U4684 (N_4684,N_4525,N_4638);
and U4685 (N_4685,N_4538,N_4567);
nand U4686 (N_4686,N_4531,N_4583);
xnor U4687 (N_4687,N_4636,N_4599);
and U4688 (N_4688,N_4637,N_4585);
or U4689 (N_4689,N_4515,N_4626);
nand U4690 (N_4690,N_4557,N_4622);
or U4691 (N_4691,N_4545,N_4564);
xnor U4692 (N_4692,N_4648,N_4533);
nand U4693 (N_4693,N_4504,N_4562);
nor U4694 (N_4694,N_4596,N_4508);
xnor U4695 (N_4695,N_4630,N_4565);
and U4696 (N_4696,N_4539,N_4575);
or U4697 (N_4697,N_4571,N_4590);
xor U4698 (N_4698,N_4519,N_4512);
or U4699 (N_4699,N_4500,N_4641);
nor U4700 (N_4700,N_4644,N_4627);
and U4701 (N_4701,N_4532,N_4589);
nor U4702 (N_4702,N_4576,N_4540);
nor U4703 (N_4703,N_4526,N_4572);
xor U4704 (N_4704,N_4573,N_4552);
nor U4705 (N_4705,N_4523,N_4507);
nor U4706 (N_4706,N_4506,N_4579);
or U4707 (N_4707,N_4597,N_4606);
xor U4708 (N_4708,N_4537,N_4555);
xnor U4709 (N_4709,N_4520,N_4570);
or U4710 (N_4710,N_4566,N_4556);
nand U4711 (N_4711,N_4534,N_4546);
nand U4712 (N_4712,N_4628,N_4640);
and U4713 (N_4713,N_4604,N_4550);
nand U4714 (N_4714,N_4578,N_4563);
nor U4715 (N_4715,N_4514,N_4559);
or U4716 (N_4716,N_4522,N_4516);
and U4717 (N_4717,N_4620,N_4605);
or U4718 (N_4718,N_4524,N_4587);
nand U4719 (N_4719,N_4618,N_4574);
or U4720 (N_4720,N_4551,N_4649);
or U4721 (N_4721,N_4607,N_4591);
or U4722 (N_4722,N_4614,N_4549);
nand U4723 (N_4723,N_4610,N_4631);
or U4724 (N_4724,N_4601,N_4528);
nand U4725 (N_4725,N_4598,N_4575);
nand U4726 (N_4726,N_4604,N_4555);
nor U4727 (N_4727,N_4642,N_4583);
or U4728 (N_4728,N_4623,N_4511);
xnor U4729 (N_4729,N_4626,N_4600);
and U4730 (N_4730,N_4648,N_4633);
and U4731 (N_4731,N_4548,N_4616);
nor U4732 (N_4732,N_4614,N_4582);
nand U4733 (N_4733,N_4608,N_4520);
and U4734 (N_4734,N_4534,N_4582);
and U4735 (N_4735,N_4555,N_4642);
nand U4736 (N_4736,N_4546,N_4555);
or U4737 (N_4737,N_4636,N_4533);
and U4738 (N_4738,N_4587,N_4546);
nor U4739 (N_4739,N_4508,N_4585);
xnor U4740 (N_4740,N_4637,N_4566);
or U4741 (N_4741,N_4578,N_4527);
nor U4742 (N_4742,N_4571,N_4526);
nand U4743 (N_4743,N_4601,N_4563);
nand U4744 (N_4744,N_4541,N_4620);
nor U4745 (N_4745,N_4556,N_4614);
or U4746 (N_4746,N_4524,N_4648);
xor U4747 (N_4747,N_4512,N_4636);
nor U4748 (N_4748,N_4553,N_4631);
or U4749 (N_4749,N_4546,N_4600);
or U4750 (N_4750,N_4529,N_4553);
and U4751 (N_4751,N_4518,N_4596);
nor U4752 (N_4752,N_4525,N_4609);
nor U4753 (N_4753,N_4605,N_4538);
xor U4754 (N_4754,N_4518,N_4610);
and U4755 (N_4755,N_4588,N_4546);
xnor U4756 (N_4756,N_4603,N_4575);
and U4757 (N_4757,N_4613,N_4503);
or U4758 (N_4758,N_4588,N_4592);
nand U4759 (N_4759,N_4609,N_4552);
nand U4760 (N_4760,N_4625,N_4513);
nor U4761 (N_4761,N_4587,N_4633);
xnor U4762 (N_4762,N_4621,N_4648);
xnor U4763 (N_4763,N_4592,N_4519);
xor U4764 (N_4764,N_4605,N_4536);
nor U4765 (N_4765,N_4582,N_4595);
nor U4766 (N_4766,N_4530,N_4512);
xnor U4767 (N_4767,N_4557,N_4558);
nor U4768 (N_4768,N_4587,N_4542);
and U4769 (N_4769,N_4532,N_4606);
nor U4770 (N_4770,N_4584,N_4573);
xnor U4771 (N_4771,N_4570,N_4574);
nand U4772 (N_4772,N_4629,N_4544);
xnor U4773 (N_4773,N_4622,N_4600);
nor U4774 (N_4774,N_4600,N_4604);
nor U4775 (N_4775,N_4546,N_4519);
and U4776 (N_4776,N_4571,N_4640);
nor U4777 (N_4777,N_4526,N_4597);
and U4778 (N_4778,N_4595,N_4541);
xnor U4779 (N_4779,N_4523,N_4627);
or U4780 (N_4780,N_4646,N_4641);
nor U4781 (N_4781,N_4514,N_4599);
nand U4782 (N_4782,N_4594,N_4593);
and U4783 (N_4783,N_4635,N_4618);
and U4784 (N_4784,N_4537,N_4524);
or U4785 (N_4785,N_4571,N_4586);
nand U4786 (N_4786,N_4644,N_4638);
or U4787 (N_4787,N_4557,N_4576);
xnor U4788 (N_4788,N_4514,N_4547);
nor U4789 (N_4789,N_4507,N_4629);
nor U4790 (N_4790,N_4631,N_4512);
and U4791 (N_4791,N_4537,N_4508);
nand U4792 (N_4792,N_4517,N_4602);
nor U4793 (N_4793,N_4591,N_4571);
nor U4794 (N_4794,N_4556,N_4572);
and U4795 (N_4795,N_4594,N_4560);
xor U4796 (N_4796,N_4613,N_4632);
nor U4797 (N_4797,N_4622,N_4645);
nor U4798 (N_4798,N_4592,N_4598);
xnor U4799 (N_4799,N_4535,N_4575);
and U4800 (N_4800,N_4664,N_4764);
nor U4801 (N_4801,N_4696,N_4728);
nand U4802 (N_4802,N_4798,N_4737);
and U4803 (N_4803,N_4703,N_4661);
and U4804 (N_4804,N_4770,N_4766);
nor U4805 (N_4805,N_4683,N_4685);
or U4806 (N_4806,N_4657,N_4656);
xnor U4807 (N_4807,N_4694,N_4773);
and U4808 (N_4808,N_4788,N_4699);
and U4809 (N_4809,N_4697,N_4675);
or U4810 (N_4810,N_4763,N_4780);
nand U4811 (N_4811,N_4722,N_4721);
and U4812 (N_4812,N_4712,N_4786);
xor U4813 (N_4813,N_4669,N_4708);
nor U4814 (N_4814,N_4672,N_4774);
nor U4815 (N_4815,N_4755,N_4713);
nand U4816 (N_4816,N_4715,N_4779);
and U4817 (N_4817,N_4794,N_4783);
xor U4818 (N_4818,N_4692,N_4736);
xnor U4819 (N_4819,N_4787,N_4727);
or U4820 (N_4820,N_4701,N_4725);
or U4821 (N_4821,N_4778,N_4709);
nor U4822 (N_4822,N_4761,N_4673);
nand U4823 (N_4823,N_4732,N_4670);
xnor U4824 (N_4824,N_4665,N_4777);
nand U4825 (N_4825,N_4793,N_4710);
and U4826 (N_4826,N_4738,N_4759);
or U4827 (N_4827,N_4726,N_4686);
xnor U4828 (N_4828,N_4754,N_4681);
xor U4829 (N_4829,N_4771,N_4693);
xor U4830 (N_4830,N_4730,N_4739);
and U4831 (N_4831,N_4796,N_4716);
nor U4832 (N_4832,N_4799,N_4653);
nor U4833 (N_4833,N_4680,N_4769);
nor U4834 (N_4834,N_4706,N_4668);
nor U4835 (N_4835,N_4695,N_4782);
and U4836 (N_4836,N_4731,N_4658);
and U4837 (N_4837,N_4678,N_4729);
and U4838 (N_4838,N_4688,N_4742);
or U4839 (N_4839,N_4785,N_4790);
xnor U4840 (N_4840,N_4768,N_4765);
and U4841 (N_4841,N_4659,N_4700);
xnor U4842 (N_4842,N_4652,N_4751);
xor U4843 (N_4843,N_4679,N_4714);
or U4844 (N_4844,N_4744,N_4662);
nand U4845 (N_4845,N_4789,N_4667);
and U4846 (N_4846,N_4682,N_4747);
xor U4847 (N_4847,N_4740,N_4752);
nor U4848 (N_4848,N_4767,N_4756);
nor U4849 (N_4849,N_4689,N_4760);
or U4850 (N_4850,N_4775,N_4758);
or U4851 (N_4851,N_4677,N_4797);
nand U4852 (N_4852,N_4684,N_4733);
or U4853 (N_4853,N_4663,N_4750);
nor U4854 (N_4854,N_4746,N_4745);
xor U4855 (N_4855,N_4717,N_4650);
xnor U4856 (N_4856,N_4691,N_4784);
nor U4857 (N_4857,N_4749,N_4723);
nor U4858 (N_4858,N_4705,N_4674);
xor U4859 (N_4859,N_4698,N_4690);
or U4860 (N_4860,N_4743,N_4791);
and U4861 (N_4861,N_4707,N_4734);
and U4862 (N_4862,N_4776,N_4655);
or U4863 (N_4863,N_4781,N_4748);
nand U4864 (N_4864,N_4702,N_4741);
xor U4865 (N_4865,N_4651,N_4757);
or U4866 (N_4866,N_4666,N_4772);
or U4867 (N_4867,N_4654,N_4687);
nor U4868 (N_4868,N_4753,N_4718);
nor U4869 (N_4869,N_4719,N_4795);
nand U4870 (N_4870,N_4660,N_4711);
nand U4871 (N_4871,N_4704,N_4735);
nand U4872 (N_4872,N_4720,N_4724);
nor U4873 (N_4873,N_4762,N_4676);
or U4874 (N_4874,N_4671,N_4792);
and U4875 (N_4875,N_4718,N_4660);
and U4876 (N_4876,N_4669,N_4685);
and U4877 (N_4877,N_4785,N_4748);
nand U4878 (N_4878,N_4747,N_4780);
or U4879 (N_4879,N_4686,N_4680);
and U4880 (N_4880,N_4717,N_4674);
nand U4881 (N_4881,N_4650,N_4796);
nand U4882 (N_4882,N_4751,N_4712);
nor U4883 (N_4883,N_4684,N_4739);
or U4884 (N_4884,N_4756,N_4716);
xnor U4885 (N_4885,N_4685,N_4739);
nor U4886 (N_4886,N_4681,N_4706);
nand U4887 (N_4887,N_4724,N_4723);
or U4888 (N_4888,N_4729,N_4655);
xor U4889 (N_4889,N_4672,N_4730);
or U4890 (N_4890,N_4716,N_4653);
nand U4891 (N_4891,N_4710,N_4704);
and U4892 (N_4892,N_4768,N_4742);
or U4893 (N_4893,N_4797,N_4757);
nor U4894 (N_4894,N_4799,N_4697);
or U4895 (N_4895,N_4684,N_4797);
nand U4896 (N_4896,N_4729,N_4728);
and U4897 (N_4897,N_4757,N_4756);
nor U4898 (N_4898,N_4749,N_4740);
nor U4899 (N_4899,N_4666,N_4695);
nor U4900 (N_4900,N_4774,N_4736);
and U4901 (N_4901,N_4706,N_4765);
nor U4902 (N_4902,N_4751,N_4654);
or U4903 (N_4903,N_4762,N_4662);
nor U4904 (N_4904,N_4678,N_4746);
and U4905 (N_4905,N_4680,N_4787);
and U4906 (N_4906,N_4686,N_4795);
and U4907 (N_4907,N_4661,N_4664);
nand U4908 (N_4908,N_4676,N_4688);
and U4909 (N_4909,N_4695,N_4743);
nor U4910 (N_4910,N_4712,N_4709);
nand U4911 (N_4911,N_4697,N_4701);
nor U4912 (N_4912,N_4753,N_4751);
nand U4913 (N_4913,N_4772,N_4796);
nand U4914 (N_4914,N_4687,N_4679);
nor U4915 (N_4915,N_4753,N_4729);
xor U4916 (N_4916,N_4777,N_4679);
nor U4917 (N_4917,N_4775,N_4672);
xnor U4918 (N_4918,N_4767,N_4722);
and U4919 (N_4919,N_4681,N_4718);
nor U4920 (N_4920,N_4731,N_4743);
nand U4921 (N_4921,N_4773,N_4744);
and U4922 (N_4922,N_4719,N_4754);
nand U4923 (N_4923,N_4659,N_4675);
nor U4924 (N_4924,N_4781,N_4669);
or U4925 (N_4925,N_4722,N_4715);
nor U4926 (N_4926,N_4751,N_4681);
nand U4927 (N_4927,N_4667,N_4754);
and U4928 (N_4928,N_4676,N_4693);
and U4929 (N_4929,N_4671,N_4789);
nor U4930 (N_4930,N_4664,N_4657);
nor U4931 (N_4931,N_4657,N_4737);
xor U4932 (N_4932,N_4678,N_4747);
or U4933 (N_4933,N_4768,N_4696);
and U4934 (N_4934,N_4736,N_4673);
and U4935 (N_4935,N_4782,N_4729);
nor U4936 (N_4936,N_4746,N_4730);
nand U4937 (N_4937,N_4672,N_4717);
or U4938 (N_4938,N_4696,N_4739);
nor U4939 (N_4939,N_4749,N_4721);
nand U4940 (N_4940,N_4791,N_4779);
nor U4941 (N_4941,N_4668,N_4733);
and U4942 (N_4942,N_4782,N_4775);
nand U4943 (N_4943,N_4734,N_4704);
and U4944 (N_4944,N_4671,N_4668);
and U4945 (N_4945,N_4681,N_4767);
or U4946 (N_4946,N_4758,N_4714);
nor U4947 (N_4947,N_4650,N_4765);
nand U4948 (N_4948,N_4748,N_4720);
xnor U4949 (N_4949,N_4777,N_4736);
or U4950 (N_4950,N_4882,N_4826);
nand U4951 (N_4951,N_4816,N_4917);
nor U4952 (N_4952,N_4836,N_4805);
and U4953 (N_4953,N_4810,N_4932);
nand U4954 (N_4954,N_4913,N_4832);
nor U4955 (N_4955,N_4938,N_4900);
xnor U4956 (N_4956,N_4827,N_4860);
or U4957 (N_4957,N_4891,N_4875);
nor U4958 (N_4958,N_4859,N_4817);
nor U4959 (N_4959,N_4918,N_4946);
nor U4960 (N_4960,N_4842,N_4925);
and U4961 (N_4961,N_4916,N_4858);
nand U4962 (N_4962,N_4895,N_4942);
nor U4963 (N_4963,N_4949,N_4829);
and U4964 (N_4964,N_4864,N_4933);
and U4965 (N_4965,N_4929,N_4930);
nor U4966 (N_4966,N_4905,N_4894);
and U4967 (N_4967,N_4849,N_4838);
and U4968 (N_4968,N_4856,N_4893);
and U4969 (N_4969,N_4907,N_4800);
and U4970 (N_4970,N_4825,N_4945);
or U4971 (N_4971,N_4897,N_4921);
and U4972 (N_4972,N_4877,N_4948);
or U4973 (N_4973,N_4820,N_4926);
and U4974 (N_4974,N_4815,N_4874);
nand U4975 (N_4975,N_4837,N_4892);
nor U4976 (N_4976,N_4867,N_4915);
and U4977 (N_4977,N_4927,N_4821);
xnor U4978 (N_4978,N_4863,N_4833);
nor U4979 (N_4979,N_4939,N_4830);
and U4980 (N_4980,N_4852,N_4808);
nand U4981 (N_4981,N_4886,N_4888);
nand U4982 (N_4982,N_4865,N_4919);
or U4983 (N_4983,N_4869,N_4881);
nor U4984 (N_4984,N_4861,N_4901);
and U4985 (N_4985,N_4890,N_4831);
nor U4986 (N_4986,N_4801,N_4844);
and U4987 (N_4987,N_4899,N_4871);
nand U4988 (N_4988,N_4944,N_4850);
or U4989 (N_4989,N_4904,N_4868);
nor U4990 (N_4990,N_4846,N_4922);
nor U4991 (N_4991,N_4873,N_4823);
nand U4992 (N_4992,N_4806,N_4885);
xnor U4993 (N_4993,N_4883,N_4937);
or U4994 (N_4994,N_4924,N_4862);
nand U4995 (N_4995,N_4870,N_4876);
nor U4996 (N_4996,N_4809,N_4824);
and U4997 (N_4997,N_4934,N_4845);
nand U4998 (N_4998,N_4872,N_4866);
nor U4999 (N_4999,N_4828,N_4841);
nand U5000 (N_5000,N_4848,N_4855);
or U5001 (N_5001,N_4943,N_4908);
nand U5002 (N_5002,N_4887,N_4879);
nand U5003 (N_5003,N_4902,N_4803);
nor U5004 (N_5004,N_4931,N_4853);
nand U5005 (N_5005,N_4851,N_4889);
or U5006 (N_5006,N_4822,N_4909);
nand U5007 (N_5007,N_4839,N_4910);
nand U5008 (N_5008,N_4923,N_4804);
nor U5009 (N_5009,N_4912,N_4914);
nand U5010 (N_5010,N_4928,N_4818);
nor U5011 (N_5011,N_4947,N_4807);
and U5012 (N_5012,N_4843,N_4911);
or U5013 (N_5013,N_4878,N_4906);
or U5014 (N_5014,N_4813,N_4811);
or U5015 (N_5015,N_4840,N_4812);
and U5016 (N_5016,N_4935,N_4903);
nand U5017 (N_5017,N_4857,N_4847);
or U5018 (N_5018,N_4884,N_4854);
nor U5019 (N_5019,N_4814,N_4835);
nand U5020 (N_5020,N_4819,N_4880);
nand U5021 (N_5021,N_4940,N_4802);
nand U5022 (N_5022,N_4898,N_4936);
nand U5023 (N_5023,N_4920,N_4896);
or U5024 (N_5024,N_4941,N_4834);
nand U5025 (N_5025,N_4821,N_4924);
xnor U5026 (N_5026,N_4941,N_4892);
and U5027 (N_5027,N_4882,N_4840);
nor U5028 (N_5028,N_4940,N_4895);
and U5029 (N_5029,N_4891,N_4906);
and U5030 (N_5030,N_4923,N_4921);
nor U5031 (N_5031,N_4838,N_4804);
and U5032 (N_5032,N_4917,N_4901);
nor U5033 (N_5033,N_4945,N_4909);
xnor U5034 (N_5034,N_4901,N_4845);
xor U5035 (N_5035,N_4816,N_4916);
xor U5036 (N_5036,N_4890,N_4863);
and U5037 (N_5037,N_4809,N_4940);
xnor U5038 (N_5038,N_4918,N_4906);
nand U5039 (N_5039,N_4924,N_4894);
or U5040 (N_5040,N_4884,N_4858);
and U5041 (N_5041,N_4803,N_4820);
or U5042 (N_5042,N_4835,N_4824);
and U5043 (N_5043,N_4891,N_4936);
and U5044 (N_5044,N_4803,N_4843);
nor U5045 (N_5045,N_4895,N_4918);
and U5046 (N_5046,N_4899,N_4857);
and U5047 (N_5047,N_4841,N_4904);
xor U5048 (N_5048,N_4907,N_4878);
nand U5049 (N_5049,N_4849,N_4805);
or U5050 (N_5050,N_4839,N_4838);
nor U5051 (N_5051,N_4850,N_4821);
nand U5052 (N_5052,N_4893,N_4927);
and U5053 (N_5053,N_4840,N_4910);
xor U5054 (N_5054,N_4830,N_4946);
xnor U5055 (N_5055,N_4826,N_4874);
or U5056 (N_5056,N_4800,N_4913);
and U5057 (N_5057,N_4909,N_4867);
xnor U5058 (N_5058,N_4838,N_4828);
nand U5059 (N_5059,N_4834,N_4851);
nand U5060 (N_5060,N_4820,N_4844);
and U5061 (N_5061,N_4910,N_4883);
and U5062 (N_5062,N_4820,N_4830);
and U5063 (N_5063,N_4911,N_4940);
and U5064 (N_5064,N_4821,N_4879);
nor U5065 (N_5065,N_4913,N_4868);
nand U5066 (N_5066,N_4867,N_4925);
nor U5067 (N_5067,N_4939,N_4878);
nor U5068 (N_5068,N_4917,N_4895);
or U5069 (N_5069,N_4928,N_4923);
nand U5070 (N_5070,N_4947,N_4894);
nor U5071 (N_5071,N_4814,N_4933);
xnor U5072 (N_5072,N_4890,N_4888);
and U5073 (N_5073,N_4895,N_4825);
nor U5074 (N_5074,N_4919,N_4904);
nor U5075 (N_5075,N_4916,N_4899);
nor U5076 (N_5076,N_4893,N_4883);
nor U5077 (N_5077,N_4831,N_4891);
xor U5078 (N_5078,N_4813,N_4836);
nand U5079 (N_5079,N_4901,N_4803);
xnor U5080 (N_5080,N_4803,N_4817);
nor U5081 (N_5081,N_4859,N_4844);
and U5082 (N_5082,N_4899,N_4911);
or U5083 (N_5083,N_4836,N_4894);
or U5084 (N_5084,N_4820,N_4871);
nand U5085 (N_5085,N_4880,N_4806);
nor U5086 (N_5086,N_4854,N_4919);
and U5087 (N_5087,N_4927,N_4863);
or U5088 (N_5088,N_4922,N_4918);
or U5089 (N_5089,N_4875,N_4927);
nor U5090 (N_5090,N_4915,N_4848);
xnor U5091 (N_5091,N_4825,N_4914);
or U5092 (N_5092,N_4920,N_4841);
nand U5093 (N_5093,N_4814,N_4926);
nand U5094 (N_5094,N_4896,N_4808);
nor U5095 (N_5095,N_4806,N_4901);
or U5096 (N_5096,N_4811,N_4845);
nand U5097 (N_5097,N_4907,N_4810);
or U5098 (N_5098,N_4873,N_4813);
xnor U5099 (N_5099,N_4810,N_4918);
nand U5100 (N_5100,N_5099,N_4964);
xor U5101 (N_5101,N_5097,N_5026);
nor U5102 (N_5102,N_5015,N_4978);
or U5103 (N_5103,N_5021,N_5066);
nand U5104 (N_5104,N_5048,N_5014);
and U5105 (N_5105,N_4969,N_4961);
xnor U5106 (N_5106,N_5050,N_5057);
xnor U5107 (N_5107,N_4959,N_5042);
or U5108 (N_5108,N_5046,N_5069);
nor U5109 (N_5109,N_5055,N_4968);
or U5110 (N_5110,N_5071,N_4966);
and U5111 (N_5111,N_5004,N_4956);
nor U5112 (N_5112,N_4998,N_5008);
nand U5113 (N_5113,N_4954,N_5003);
xnor U5114 (N_5114,N_4979,N_5025);
nand U5115 (N_5115,N_4995,N_5088);
and U5116 (N_5116,N_5063,N_5047);
nor U5117 (N_5117,N_5058,N_4971);
nand U5118 (N_5118,N_5023,N_4957);
xnor U5119 (N_5119,N_4996,N_5051);
xnor U5120 (N_5120,N_5022,N_5028);
nand U5121 (N_5121,N_4977,N_5061);
nand U5122 (N_5122,N_5054,N_5020);
or U5123 (N_5123,N_5011,N_5018);
nor U5124 (N_5124,N_5037,N_5078);
or U5125 (N_5125,N_4986,N_4997);
nor U5126 (N_5126,N_4965,N_5034);
or U5127 (N_5127,N_5062,N_4990);
xnor U5128 (N_5128,N_5039,N_5036);
or U5129 (N_5129,N_5079,N_5052);
or U5130 (N_5130,N_4980,N_4970);
and U5131 (N_5131,N_5000,N_4958);
nor U5132 (N_5132,N_5010,N_5087);
xnor U5133 (N_5133,N_5038,N_5049);
xnor U5134 (N_5134,N_5012,N_5029);
xnor U5135 (N_5135,N_4999,N_5043);
and U5136 (N_5136,N_5094,N_5096);
xor U5137 (N_5137,N_5060,N_5009);
xor U5138 (N_5138,N_4955,N_5032);
or U5139 (N_5139,N_5002,N_5027);
or U5140 (N_5140,N_5089,N_5041);
and U5141 (N_5141,N_4950,N_5077);
nand U5142 (N_5142,N_5074,N_5067);
xor U5143 (N_5143,N_5007,N_4952);
nor U5144 (N_5144,N_5065,N_5086);
xnor U5145 (N_5145,N_4973,N_4953);
xnor U5146 (N_5146,N_5068,N_5092);
and U5147 (N_5147,N_5030,N_5059);
nor U5148 (N_5148,N_4981,N_5081);
or U5149 (N_5149,N_4987,N_5016);
and U5150 (N_5150,N_5090,N_5056);
xnor U5151 (N_5151,N_5005,N_4982);
or U5152 (N_5152,N_4984,N_4974);
xnor U5153 (N_5153,N_5093,N_4960);
and U5154 (N_5154,N_5095,N_5006);
and U5155 (N_5155,N_4975,N_4993);
and U5156 (N_5156,N_4967,N_5040);
nor U5157 (N_5157,N_5024,N_4963);
and U5158 (N_5158,N_5031,N_5080);
nor U5159 (N_5159,N_5035,N_5072);
xor U5160 (N_5160,N_4962,N_5064);
nand U5161 (N_5161,N_5075,N_5073);
xor U5162 (N_5162,N_5001,N_4994);
nand U5163 (N_5163,N_5070,N_4985);
nor U5164 (N_5164,N_4972,N_5091);
nand U5165 (N_5165,N_4976,N_5083);
nand U5166 (N_5166,N_5045,N_5084);
nor U5167 (N_5167,N_5076,N_4989);
nand U5168 (N_5168,N_5013,N_4988);
and U5169 (N_5169,N_4983,N_5082);
xor U5170 (N_5170,N_5098,N_4991);
or U5171 (N_5171,N_5053,N_4992);
xnor U5172 (N_5172,N_5044,N_5017);
nand U5173 (N_5173,N_5019,N_5085);
or U5174 (N_5174,N_4951,N_5033);
nor U5175 (N_5175,N_5091,N_4991);
nor U5176 (N_5176,N_5013,N_4976);
and U5177 (N_5177,N_5099,N_4996);
nand U5178 (N_5178,N_4999,N_5017);
and U5179 (N_5179,N_5004,N_4983);
or U5180 (N_5180,N_5018,N_5092);
xor U5181 (N_5181,N_5006,N_4960);
xnor U5182 (N_5182,N_5094,N_4984);
or U5183 (N_5183,N_4960,N_5097);
or U5184 (N_5184,N_5055,N_4971);
or U5185 (N_5185,N_5058,N_5029);
xor U5186 (N_5186,N_4992,N_5095);
nor U5187 (N_5187,N_5026,N_4958);
nor U5188 (N_5188,N_5063,N_5052);
and U5189 (N_5189,N_5054,N_5029);
nor U5190 (N_5190,N_5079,N_4984);
and U5191 (N_5191,N_4984,N_5043);
xor U5192 (N_5192,N_5060,N_4966);
nor U5193 (N_5193,N_5075,N_5098);
xor U5194 (N_5194,N_5019,N_5071);
nor U5195 (N_5195,N_5025,N_4975);
and U5196 (N_5196,N_5012,N_5097);
or U5197 (N_5197,N_4988,N_5003);
xnor U5198 (N_5198,N_4982,N_5028);
nor U5199 (N_5199,N_4973,N_4956);
nand U5200 (N_5200,N_5084,N_4980);
and U5201 (N_5201,N_5057,N_5002);
nand U5202 (N_5202,N_5059,N_4973);
or U5203 (N_5203,N_5080,N_5037);
nor U5204 (N_5204,N_5091,N_5074);
xor U5205 (N_5205,N_5097,N_5011);
xor U5206 (N_5206,N_5053,N_5061);
nor U5207 (N_5207,N_4963,N_5075);
and U5208 (N_5208,N_5002,N_4959);
or U5209 (N_5209,N_5079,N_4981);
nand U5210 (N_5210,N_5094,N_4957);
nand U5211 (N_5211,N_4960,N_5010);
nor U5212 (N_5212,N_5053,N_5062);
and U5213 (N_5213,N_4963,N_5042);
nand U5214 (N_5214,N_5080,N_5064);
and U5215 (N_5215,N_4954,N_5077);
xnor U5216 (N_5216,N_5000,N_5070);
xnor U5217 (N_5217,N_5077,N_5009);
and U5218 (N_5218,N_5093,N_5090);
nor U5219 (N_5219,N_5053,N_5003);
nand U5220 (N_5220,N_5046,N_4989);
nand U5221 (N_5221,N_5048,N_5068);
nand U5222 (N_5222,N_5016,N_5043);
xor U5223 (N_5223,N_4967,N_5078);
xor U5224 (N_5224,N_4983,N_4966);
nor U5225 (N_5225,N_5052,N_5009);
nor U5226 (N_5226,N_5096,N_4971);
nand U5227 (N_5227,N_5076,N_5045);
and U5228 (N_5228,N_5014,N_5080);
xnor U5229 (N_5229,N_5053,N_5040);
nor U5230 (N_5230,N_5031,N_4968);
nor U5231 (N_5231,N_5082,N_5075);
and U5232 (N_5232,N_5093,N_5012);
or U5233 (N_5233,N_5069,N_4963);
nor U5234 (N_5234,N_4985,N_5047);
xor U5235 (N_5235,N_4999,N_5029);
or U5236 (N_5236,N_5001,N_4971);
and U5237 (N_5237,N_4997,N_4973);
or U5238 (N_5238,N_5061,N_4994);
nor U5239 (N_5239,N_5056,N_5016);
xor U5240 (N_5240,N_4971,N_5023);
xor U5241 (N_5241,N_5034,N_5060);
nor U5242 (N_5242,N_5043,N_4969);
xnor U5243 (N_5243,N_4984,N_5056);
and U5244 (N_5244,N_4956,N_5064);
or U5245 (N_5245,N_5027,N_5014);
nand U5246 (N_5246,N_4961,N_5069);
or U5247 (N_5247,N_5063,N_4998);
and U5248 (N_5248,N_5064,N_5012);
nor U5249 (N_5249,N_5057,N_5025);
or U5250 (N_5250,N_5160,N_5135);
or U5251 (N_5251,N_5151,N_5192);
and U5252 (N_5252,N_5134,N_5209);
and U5253 (N_5253,N_5215,N_5133);
nor U5254 (N_5254,N_5204,N_5180);
nand U5255 (N_5255,N_5223,N_5111);
xor U5256 (N_5256,N_5155,N_5173);
nand U5257 (N_5257,N_5200,N_5186);
or U5258 (N_5258,N_5236,N_5211);
or U5259 (N_5259,N_5143,N_5125);
nor U5260 (N_5260,N_5237,N_5231);
or U5261 (N_5261,N_5241,N_5185);
and U5262 (N_5262,N_5116,N_5233);
nand U5263 (N_5263,N_5183,N_5187);
or U5264 (N_5264,N_5194,N_5170);
nand U5265 (N_5265,N_5174,N_5196);
or U5266 (N_5266,N_5219,N_5218);
xor U5267 (N_5267,N_5229,N_5130);
nand U5268 (N_5268,N_5113,N_5195);
xnor U5269 (N_5269,N_5238,N_5172);
nor U5270 (N_5270,N_5189,N_5127);
xor U5271 (N_5271,N_5107,N_5145);
nand U5272 (N_5272,N_5157,N_5190);
nor U5273 (N_5273,N_5106,N_5142);
nor U5274 (N_5274,N_5217,N_5199);
and U5275 (N_5275,N_5166,N_5132);
nor U5276 (N_5276,N_5240,N_5137);
and U5277 (N_5277,N_5176,N_5129);
and U5278 (N_5278,N_5210,N_5126);
or U5279 (N_5279,N_5118,N_5152);
nand U5280 (N_5280,N_5239,N_5184);
nor U5281 (N_5281,N_5246,N_5109);
and U5282 (N_5282,N_5191,N_5161);
or U5283 (N_5283,N_5245,N_5188);
nand U5284 (N_5284,N_5207,N_5220);
or U5285 (N_5285,N_5150,N_5197);
nor U5286 (N_5286,N_5122,N_5104);
or U5287 (N_5287,N_5226,N_5242);
xnor U5288 (N_5288,N_5216,N_5202);
nand U5289 (N_5289,N_5158,N_5178);
nand U5290 (N_5290,N_5201,N_5153);
or U5291 (N_5291,N_5119,N_5131);
or U5292 (N_5292,N_5103,N_5140);
nor U5293 (N_5293,N_5206,N_5227);
nor U5294 (N_5294,N_5165,N_5105);
or U5295 (N_5295,N_5171,N_5232);
nor U5296 (N_5296,N_5225,N_5120);
and U5297 (N_5297,N_5128,N_5168);
or U5298 (N_5298,N_5100,N_5205);
or U5299 (N_5299,N_5146,N_5243);
nand U5300 (N_5300,N_5212,N_5247);
nor U5301 (N_5301,N_5169,N_5121);
nor U5302 (N_5302,N_5235,N_5147);
and U5303 (N_5303,N_5234,N_5222);
nand U5304 (N_5304,N_5136,N_5248);
and U5305 (N_5305,N_5163,N_5148);
and U5306 (N_5306,N_5138,N_5182);
and U5307 (N_5307,N_5249,N_5139);
and U5308 (N_5308,N_5101,N_5164);
nand U5309 (N_5309,N_5177,N_5167);
nand U5310 (N_5310,N_5141,N_5208);
nand U5311 (N_5311,N_5193,N_5203);
nor U5312 (N_5312,N_5175,N_5159);
nor U5313 (N_5313,N_5102,N_5123);
nand U5314 (N_5314,N_5154,N_5115);
nor U5315 (N_5315,N_5108,N_5156);
or U5316 (N_5316,N_5214,N_5213);
xnor U5317 (N_5317,N_5149,N_5181);
or U5318 (N_5318,N_5162,N_5144);
or U5319 (N_5319,N_5110,N_5117);
and U5320 (N_5320,N_5198,N_5244);
or U5321 (N_5321,N_5230,N_5112);
nor U5322 (N_5322,N_5224,N_5228);
and U5323 (N_5323,N_5221,N_5124);
or U5324 (N_5324,N_5179,N_5114);
xor U5325 (N_5325,N_5114,N_5226);
xnor U5326 (N_5326,N_5168,N_5232);
xnor U5327 (N_5327,N_5189,N_5160);
nor U5328 (N_5328,N_5136,N_5112);
nor U5329 (N_5329,N_5162,N_5238);
and U5330 (N_5330,N_5166,N_5196);
nand U5331 (N_5331,N_5114,N_5121);
and U5332 (N_5332,N_5190,N_5184);
nand U5333 (N_5333,N_5134,N_5110);
and U5334 (N_5334,N_5155,N_5195);
xnor U5335 (N_5335,N_5117,N_5129);
or U5336 (N_5336,N_5230,N_5126);
nand U5337 (N_5337,N_5221,N_5248);
or U5338 (N_5338,N_5212,N_5218);
xnor U5339 (N_5339,N_5107,N_5244);
and U5340 (N_5340,N_5228,N_5103);
nor U5341 (N_5341,N_5135,N_5103);
or U5342 (N_5342,N_5208,N_5113);
or U5343 (N_5343,N_5246,N_5145);
xnor U5344 (N_5344,N_5242,N_5198);
and U5345 (N_5345,N_5164,N_5196);
and U5346 (N_5346,N_5231,N_5141);
nor U5347 (N_5347,N_5229,N_5162);
nand U5348 (N_5348,N_5124,N_5233);
nand U5349 (N_5349,N_5190,N_5192);
or U5350 (N_5350,N_5144,N_5125);
nor U5351 (N_5351,N_5151,N_5105);
and U5352 (N_5352,N_5230,N_5213);
nor U5353 (N_5353,N_5100,N_5234);
xor U5354 (N_5354,N_5221,N_5161);
nor U5355 (N_5355,N_5211,N_5248);
and U5356 (N_5356,N_5176,N_5240);
and U5357 (N_5357,N_5191,N_5189);
nand U5358 (N_5358,N_5221,N_5131);
or U5359 (N_5359,N_5118,N_5151);
xor U5360 (N_5360,N_5166,N_5211);
or U5361 (N_5361,N_5126,N_5238);
or U5362 (N_5362,N_5200,N_5163);
nor U5363 (N_5363,N_5175,N_5238);
xor U5364 (N_5364,N_5136,N_5193);
xor U5365 (N_5365,N_5220,N_5233);
nor U5366 (N_5366,N_5207,N_5239);
or U5367 (N_5367,N_5144,N_5189);
and U5368 (N_5368,N_5102,N_5225);
and U5369 (N_5369,N_5150,N_5183);
nand U5370 (N_5370,N_5196,N_5146);
or U5371 (N_5371,N_5227,N_5121);
or U5372 (N_5372,N_5184,N_5202);
and U5373 (N_5373,N_5108,N_5215);
or U5374 (N_5374,N_5157,N_5184);
nand U5375 (N_5375,N_5245,N_5230);
or U5376 (N_5376,N_5163,N_5155);
or U5377 (N_5377,N_5222,N_5239);
nand U5378 (N_5378,N_5232,N_5166);
nand U5379 (N_5379,N_5244,N_5160);
xnor U5380 (N_5380,N_5249,N_5212);
or U5381 (N_5381,N_5200,N_5165);
xnor U5382 (N_5382,N_5242,N_5186);
nor U5383 (N_5383,N_5181,N_5194);
and U5384 (N_5384,N_5186,N_5129);
xor U5385 (N_5385,N_5241,N_5141);
and U5386 (N_5386,N_5212,N_5143);
nor U5387 (N_5387,N_5153,N_5126);
nor U5388 (N_5388,N_5107,N_5215);
nand U5389 (N_5389,N_5206,N_5221);
nand U5390 (N_5390,N_5119,N_5220);
or U5391 (N_5391,N_5110,N_5120);
nand U5392 (N_5392,N_5138,N_5183);
nor U5393 (N_5393,N_5159,N_5240);
nor U5394 (N_5394,N_5200,N_5238);
nand U5395 (N_5395,N_5193,N_5219);
nand U5396 (N_5396,N_5122,N_5136);
nand U5397 (N_5397,N_5165,N_5138);
or U5398 (N_5398,N_5197,N_5218);
xnor U5399 (N_5399,N_5149,N_5228);
or U5400 (N_5400,N_5258,N_5363);
xor U5401 (N_5401,N_5340,N_5341);
nor U5402 (N_5402,N_5299,N_5384);
nor U5403 (N_5403,N_5254,N_5297);
xor U5404 (N_5404,N_5264,N_5255);
xor U5405 (N_5405,N_5323,N_5399);
xnor U5406 (N_5406,N_5262,N_5312);
xnor U5407 (N_5407,N_5390,N_5337);
or U5408 (N_5408,N_5383,N_5291);
xnor U5409 (N_5409,N_5273,N_5349);
xor U5410 (N_5410,N_5376,N_5360);
xnor U5411 (N_5411,N_5282,N_5388);
or U5412 (N_5412,N_5310,N_5303);
nor U5413 (N_5413,N_5329,N_5276);
nand U5414 (N_5414,N_5306,N_5294);
xnor U5415 (N_5415,N_5304,N_5257);
or U5416 (N_5416,N_5356,N_5320);
nand U5417 (N_5417,N_5277,N_5298);
and U5418 (N_5418,N_5319,N_5366);
xnor U5419 (N_5419,N_5346,N_5293);
nand U5420 (N_5420,N_5268,N_5382);
and U5421 (N_5421,N_5370,N_5335);
or U5422 (N_5422,N_5362,N_5342);
nand U5423 (N_5423,N_5317,N_5321);
nand U5424 (N_5424,N_5330,N_5266);
nor U5425 (N_5425,N_5379,N_5386);
nand U5426 (N_5426,N_5283,N_5375);
and U5427 (N_5427,N_5269,N_5345);
nor U5428 (N_5428,N_5353,N_5261);
or U5429 (N_5429,N_5309,N_5389);
or U5430 (N_5430,N_5271,N_5290);
and U5431 (N_5431,N_5252,N_5336);
or U5432 (N_5432,N_5365,N_5259);
nand U5433 (N_5433,N_5387,N_5324);
nand U5434 (N_5434,N_5274,N_5393);
and U5435 (N_5435,N_5352,N_5316);
nor U5436 (N_5436,N_5380,N_5272);
nand U5437 (N_5437,N_5275,N_5250);
or U5438 (N_5438,N_5333,N_5367);
and U5439 (N_5439,N_5301,N_5281);
nor U5440 (N_5440,N_5339,N_5343);
nand U5441 (N_5441,N_5295,N_5394);
or U5442 (N_5442,N_5357,N_5289);
nor U5443 (N_5443,N_5397,N_5334);
nand U5444 (N_5444,N_5260,N_5358);
and U5445 (N_5445,N_5286,N_5308);
and U5446 (N_5446,N_5398,N_5256);
or U5447 (N_5447,N_5338,N_5285);
and U5448 (N_5448,N_5287,N_5265);
nor U5449 (N_5449,N_5392,N_5300);
nand U5450 (N_5450,N_5251,N_5278);
nand U5451 (N_5451,N_5348,N_5396);
nand U5452 (N_5452,N_5270,N_5327);
and U5453 (N_5453,N_5369,N_5263);
and U5454 (N_5454,N_5280,N_5332);
and U5455 (N_5455,N_5381,N_5311);
and U5456 (N_5456,N_5347,N_5322);
or U5457 (N_5457,N_5279,N_5315);
or U5458 (N_5458,N_5373,N_5364);
nor U5459 (N_5459,N_5378,N_5328);
and U5460 (N_5460,N_5359,N_5371);
xor U5461 (N_5461,N_5350,N_5325);
and U5462 (N_5462,N_5288,N_5313);
xnor U5463 (N_5463,N_5296,N_5372);
and U5464 (N_5464,N_5331,N_5318);
nor U5465 (N_5465,N_5267,N_5284);
nand U5466 (N_5466,N_5302,N_5354);
and U5467 (N_5467,N_5314,N_5377);
or U5468 (N_5468,N_5326,N_5292);
nor U5469 (N_5469,N_5344,N_5385);
xnor U5470 (N_5470,N_5368,N_5361);
or U5471 (N_5471,N_5305,N_5355);
or U5472 (N_5472,N_5374,N_5351);
and U5473 (N_5473,N_5307,N_5253);
and U5474 (N_5474,N_5395,N_5391);
xnor U5475 (N_5475,N_5273,N_5357);
xor U5476 (N_5476,N_5324,N_5255);
nor U5477 (N_5477,N_5281,N_5272);
xnor U5478 (N_5478,N_5285,N_5328);
nand U5479 (N_5479,N_5260,N_5326);
nor U5480 (N_5480,N_5359,N_5335);
xor U5481 (N_5481,N_5276,N_5398);
and U5482 (N_5482,N_5350,N_5383);
nor U5483 (N_5483,N_5288,N_5292);
xnor U5484 (N_5484,N_5393,N_5375);
and U5485 (N_5485,N_5283,N_5294);
nand U5486 (N_5486,N_5271,N_5321);
xor U5487 (N_5487,N_5288,N_5269);
nand U5488 (N_5488,N_5263,N_5281);
nand U5489 (N_5489,N_5361,N_5263);
nor U5490 (N_5490,N_5347,N_5339);
or U5491 (N_5491,N_5381,N_5346);
or U5492 (N_5492,N_5274,N_5379);
xor U5493 (N_5493,N_5332,N_5298);
xor U5494 (N_5494,N_5323,N_5392);
xnor U5495 (N_5495,N_5311,N_5304);
xnor U5496 (N_5496,N_5265,N_5333);
nor U5497 (N_5497,N_5308,N_5319);
nand U5498 (N_5498,N_5282,N_5380);
and U5499 (N_5499,N_5311,N_5252);
nand U5500 (N_5500,N_5297,N_5376);
nor U5501 (N_5501,N_5264,N_5308);
nand U5502 (N_5502,N_5284,N_5263);
or U5503 (N_5503,N_5275,N_5255);
or U5504 (N_5504,N_5302,N_5266);
nand U5505 (N_5505,N_5357,N_5353);
or U5506 (N_5506,N_5379,N_5324);
or U5507 (N_5507,N_5375,N_5321);
and U5508 (N_5508,N_5289,N_5376);
nor U5509 (N_5509,N_5330,N_5380);
or U5510 (N_5510,N_5313,N_5341);
nand U5511 (N_5511,N_5362,N_5300);
xor U5512 (N_5512,N_5385,N_5369);
nor U5513 (N_5513,N_5266,N_5327);
or U5514 (N_5514,N_5266,N_5292);
nand U5515 (N_5515,N_5259,N_5285);
and U5516 (N_5516,N_5352,N_5270);
and U5517 (N_5517,N_5264,N_5272);
nor U5518 (N_5518,N_5381,N_5297);
nor U5519 (N_5519,N_5312,N_5379);
xor U5520 (N_5520,N_5300,N_5352);
xnor U5521 (N_5521,N_5267,N_5258);
or U5522 (N_5522,N_5271,N_5377);
or U5523 (N_5523,N_5307,N_5383);
xor U5524 (N_5524,N_5320,N_5339);
nand U5525 (N_5525,N_5271,N_5297);
nor U5526 (N_5526,N_5345,N_5355);
nor U5527 (N_5527,N_5344,N_5255);
nor U5528 (N_5528,N_5273,N_5341);
xor U5529 (N_5529,N_5386,N_5306);
nand U5530 (N_5530,N_5363,N_5374);
nor U5531 (N_5531,N_5357,N_5397);
xnor U5532 (N_5532,N_5264,N_5344);
nand U5533 (N_5533,N_5355,N_5370);
or U5534 (N_5534,N_5389,N_5357);
xnor U5535 (N_5535,N_5316,N_5267);
or U5536 (N_5536,N_5301,N_5320);
or U5537 (N_5537,N_5327,N_5393);
or U5538 (N_5538,N_5328,N_5292);
and U5539 (N_5539,N_5319,N_5281);
nand U5540 (N_5540,N_5299,N_5317);
or U5541 (N_5541,N_5325,N_5339);
or U5542 (N_5542,N_5331,N_5292);
and U5543 (N_5543,N_5257,N_5376);
and U5544 (N_5544,N_5315,N_5357);
xor U5545 (N_5545,N_5282,N_5344);
nand U5546 (N_5546,N_5316,N_5328);
nor U5547 (N_5547,N_5323,N_5361);
xor U5548 (N_5548,N_5308,N_5269);
xor U5549 (N_5549,N_5265,N_5346);
and U5550 (N_5550,N_5444,N_5427);
and U5551 (N_5551,N_5442,N_5413);
xnor U5552 (N_5552,N_5545,N_5517);
xor U5553 (N_5553,N_5541,N_5499);
xnor U5554 (N_5554,N_5529,N_5497);
and U5555 (N_5555,N_5480,N_5428);
nor U5556 (N_5556,N_5492,N_5511);
and U5557 (N_5557,N_5403,N_5530);
and U5558 (N_5558,N_5487,N_5464);
xor U5559 (N_5559,N_5482,N_5440);
nor U5560 (N_5560,N_5512,N_5515);
nor U5561 (N_5561,N_5520,N_5420);
nand U5562 (N_5562,N_5411,N_5435);
or U5563 (N_5563,N_5546,N_5498);
or U5564 (N_5564,N_5489,N_5475);
nor U5565 (N_5565,N_5449,N_5485);
xnor U5566 (N_5566,N_5412,N_5457);
xnor U5567 (N_5567,N_5453,N_5402);
nand U5568 (N_5568,N_5407,N_5510);
or U5569 (N_5569,N_5465,N_5491);
xor U5570 (N_5570,N_5494,N_5523);
nand U5571 (N_5571,N_5547,N_5404);
nor U5572 (N_5572,N_5421,N_5532);
nand U5573 (N_5573,N_5437,N_5509);
or U5574 (N_5574,N_5496,N_5500);
and U5575 (N_5575,N_5549,N_5466);
or U5576 (N_5576,N_5531,N_5528);
nand U5577 (N_5577,N_5486,N_5460);
and U5578 (N_5578,N_5524,N_5448);
nor U5579 (N_5579,N_5534,N_5405);
nor U5580 (N_5580,N_5470,N_5483);
nor U5581 (N_5581,N_5414,N_5468);
or U5582 (N_5582,N_5533,N_5406);
xor U5583 (N_5583,N_5472,N_5518);
and U5584 (N_5584,N_5543,N_5436);
xnor U5585 (N_5585,N_5501,N_5521);
nand U5586 (N_5586,N_5503,N_5538);
nor U5587 (N_5587,N_5454,N_5445);
nor U5588 (N_5588,N_5474,N_5456);
xor U5589 (N_5589,N_5416,N_5459);
nor U5590 (N_5590,N_5537,N_5479);
nand U5591 (N_5591,N_5410,N_5493);
or U5592 (N_5592,N_5471,N_5504);
xnor U5593 (N_5593,N_5495,N_5455);
xnor U5594 (N_5594,N_5525,N_5522);
or U5595 (N_5595,N_5422,N_5544);
xnor U5596 (N_5596,N_5490,N_5450);
xnor U5597 (N_5597,N_5513,N_5452);
or U5598 (N_5598,N_5408,N_5432);
or U5599 (N_5599,N_5514,N_5548);
nor U5600 (N_5600,N_5478,N_5540);
or U5601 (N_5601,N_5400,N_5476);
and U5602 (N_5602,N_5401,N_5481);
or U5603 (N_5603,N_5535,N_5516);
xor U5604 (N_5604,N_5461,N_5429);
nand U5605 (N_5605,N_5419,N_5441);
nand U5606 (N_5606,N_5488,N_5484);
and U5607 (N_5607,N_5446,N_5438);
or U5608 (N_5608,N_5542,N_5502);
xnor U5609 (N_5609,N_5477,N_5431);
xnor U5610 (N_5610,N_5539,N_5505);
nand U5611 (N_5611,N_5467,N_5473);
xnor U5612 (N_5612,N_5433,N_5409);
or U5613 (N_5613,N_5443,N_5424);
nand U5614 (N_5614,N_5526,N_5506);
xor U5615 (N_5615,N_5425,N_5458);
or U5616 (N_5616,N_5519,N_5463);
and U5617 (N_5617,N_5423,N_5462);
nor U5618 (N_5618,N_5536,N_5527);
nand U5619 (N_5619,N_5447,N_5417);
nor U5620 (N_5620,N_5418,N_5508);
nor U5621 (N_5621,N_5415,N_5507);
and U5622 (N_5622,N_5451,N_5469);
nand U5623 (N_5623,N_5434,N_5426);
nor U5624 (N_5624,N_5430,N_5439);
and U5625 (N_5625,N_5531,N_5529);
xnor U5626 (N_5626,N_5435,N_5538);
xnor U5627 (N_5627,N_5499,N_5549);
nand U5628 (N_5628,N_5408,N_5528);
nand U5629 (N_5629,N_5410,N_5440);
nand U5630 (N_5630,N_5419,N_5460);
xor U5631 (N_5631,N_5532,N_5438);
xor U5632 (N_5632,N_5539,N_5511);
nand U5633 (N_5633,N_5548,N_5444);
or U5634 (N_5634,N_5524,N_5461);
or U5635 (N_5635,N_5547,N_5545);
and U5636 (N_5636,N_5543,N_5499);
or U5637 (N_5637,N_5475,N_5432);
and U5638 (N_5638,N_5426,N_5457);
and U5639 (N_5639,N_5420,N_5473);
nor U5640 (N_5640,N_5476,N_5523);
nor U5641 (N_5641,N_5515,N_5426);
nor U5642 (N_5642,N_5411,N_5469);
xnor U5643 (N_5643,N_5501,N_5470);
or U5644 (N_5644,N_5474,N_5524);
or U5645 (N_5645,N_5529,N_5408);
nand U5646 (N_5646,N_5406,N_5461);
nor U5647 (N_5647,N_5449,N_5524);
and U5648 (N_5648,N_5451,N_5521);
nor U5649 (N_5649,N_5466,N_5537);
or U5650 (N_5650,N_5463,N_5439);
nor U5651 (N_5651,N_5537,N_5515);
nand U5652 (N_5652,N_5522,N_5427);
nor U5653 (N_5653,N_5543,N_5510);
nor U5654 (N_5654,N_5430,N_5414);
nor U5655 (N_5655,N_5496,N_5477);
or U5656 (N_5656,N_5441,N_5405);
nand U5657 (N_5657,N_5425,N_5450);
and U5658 (N_5658,N_5465,N_5479);
or U5659 (N_5659,N_5512,N_5421);
and U5660 (N_5660,N_5523,N_5438);
or U5661 (N_5661,N_5452,N_5511);
nor U5662 (N_5662,N_5505,N_5474);
nor U5663 (N_5663,N_5536,N_5487);
or U5664 (N_5664,N_5403,N_5419);
nor U5665 (N_5665,N_5498,N_5463);
xnor U5666 (N_5666,N_5475,N_5434);
nand U5667 (N_5667,N_5518,N_5544);
nand U5668 (N_5668,N_5549,N_5543);
and U5669 (N_5669,N_5536,N_5508);
and U5670 (N_5670,N_5406,N_5439);
nand U5671 (N_5671,N_5466,N_5455);
or U5672 (N_5672,N_5456,N_5423);
xnor U5673 (N_5673,N_5541,N_5486);
nor U5674 (N_5674,N_5540,N_5503);
or U5675 (N_5675,N_5473,N_5437);
or U5676 (N_5676,N_5463,N_5402);
and U5677 (N_5677,N_5518,N_5406);
and U5678 (N_5678,N_5512,N_5431);
nand U5679 (N_5679,N_5422,N_5522);
xor U5680 (N_5680,N_5540,N_5420);
or U5681 (N_5681,N_5533,N_5415);
or U5682 (N_5682,N_5463,N_5452);
or U5683 (N_5683,N_5416,N_5498);
xnor U5684 (N_5684,N_5411,N_5499);
and U5685 (N_5685,N_5427,N_5545);
and U5686 (N_5686,N_5409,N_5478);
xnor U5687 (N_5687,N_5422,N_5512);
nor U5688 (N_5688,N_5517,N_5528);
and U5689 (N_5689,N_5459,N_5466);
xor U5690 (N_5690,N_5524,N_5452);
and U5691 (N_5691,N_5502,N_5472);
nor U5692 (N_5692,N_5488,N_5476);
nor U5693 (N_5693,N_5462,N_5401);
nor U5694 (N_5694,N_5537,N_5477);
nand U5695 (N_5695,N_5494,N_5461);
and U5696 (N_5696,N_5504,N_5534);
nor U5697 (N_5697,N_5452,N_5521);
and U5698 (N_5698,N_5499,N_5510);
nor U5699 (N_5699,N_5413,N_5495);
nor U5700 (N_5700,N_5599,N_5566);
or U5701 (N_5701,N_5697,N_5581);
nand U5702 (N_5702,N_5678,N_5551);
nand U5703 (N_5703,N_5654,N_5683);
and U5704 (N_5704,N_5668,N_5629);
and U5705 (N_5705,N_5635,N_5589);
nor U5706 (N_5706,N_5613,N_5680);
nor U5707 (N_5707,N_5661,N_5602);
nor U5708 (N_5708,N_5575,N_5659);
and U5709 (N_5709,N_5649,N_5699);
nand U5710 (N_5710,N_5582,N_5553);
and U5711 (N_5711,N_5615,N_5552);
and U5712 (N_5712,N_5648,N_5651);
xnor U5713 (N_5713,N_5671,N_5669);
nand U5714 (N_5714,N_5611,N_5591);
and U5715 (N_5715,N_5637,N_5624);
xor U5716 (N_5716,N_5638,N_5647);
xor U5717 (N_5717,N_5567,N_5593);
or U5718 (N_5718,N_5564,N_5627);
and U5719 (N_5719,N_5557,N_5662);
nand U5720 (N_5720,N_5586,N_5633);
nor U5721 (N_5721,N_5685,N_5691);
nand U5722 (N_5722,N_5643,N_5574);
and U5723 (N_5723,N_5622,N_5621);
and U5724 (N_5724,N_5609,N_5561);
and U5725 (N_5725,N_5558,N_5687);
nor U5726 (N_5726,N_5568,N_5618);
nand U5727 (N_5727,N_5597,N_5625);
or U5728 (N_5728,N_5628,N_5692);
xor U5729 (N_5729,N_5681,N_5610);
and U5730 (N_5730,N_5579,N_5570);
nor U5731 (N_5731,N_5601,N_5630);
and U5732 (N_5732,N_5682,N_5690);
xnor U5733 (N_5733,N_5631,N_5612);
and U5734 (N_5734,N_5600,N_5657);
nor U5735 (N_5735,N_5584,N_5693);
nor U5736 (N_5736,N_5587,N_5652);
xnor U5737 (N_5737,N_5595,N_5658);
and U5738 (N_5738,N_5555,N_5644);
and U5739 (N_5739,N_5619,N_5585);
nor U5740 (N_5740,N_5620,N_5688);
or U5741 (N_5741,N_5604,N_5663);
nor U5742 (N_5742,N_5560,N_5623);
or U5743 (N_5743,N_5675,N_5590);
nor U5744 (N_5744,N_5642,N_5580);
or U5745 (N_5745,N_5684,N_5641);
and U5746 (N_5746,N_5640,N_5565);
nand U5747 (N_5747,N_5686,N_5606);
or U5748 (N_5748,N_5650,N_5656);
nor U5749 (N_5749,N_5616,N_5634);
nor U5750 (N_5750,N_5603,N_5592);
nand U5751 (N_5751,N_5576,N_5563);
nand U5752 (N_5752,N_5673,N_5596);
and U5753 (N_5753,N_5588,N_5598);
xnor U5754 (N_5754,N_5639,N_5646);
or U5755 (N_5755,N_5617,N_5569);
xor U5756 (N_5756,N_5556,N_5571);
nand U5757 (N_5757,N_5632,N_5605);
nor U5758 (N_5758,N_5562,N_5664);
nand U5759 (N_5759,N_5666,N_5583);
and U5760 (N_5760,N_5653,N_5572);
and U5761 (N_5761,N_5655,N_5607);
and U5762 (N_5762,N_5698,N_5660);
and U5763 (N_5763,N_5573,N_5689);
or U5764 (N_5764,N_5550,N_5578);
or U5765 (N_5765,N_5594,N_5608);
or U5766 (N_5766,N_5670,N_5667);
nor U5767 (N_5767,N_5554,N_5645);
and U5768 (N_5768,N_5577,N_5665);
nand U5769 (N_5769,N_5677,N_5679);
nand U5770 (N_5770,N_5636,N_5694);
and U5771 (N_5771,N_5674,N_5696);
and U5772 (N_5772,N_5559,N_5614);
or U5773 (N_5773,N_5672,N_5676);
nand U5774 (N_5774,N_5626,N_5695);
xor U5775 (N_5775,N_5666,N_5615);
nor U5776 (N_5776,N_5554,N_5600);
nand U5777 (N_5777,N_5662,N_5555);
nor U5778 (N_5778,N_5617,N_5586);
nand U5779 (N_5779,N_5678,N_5550);
nand U5780 (N_5780,N_5580,N_5698);
nor U5781 (N_5781,N_5563,N_5662);
nand U5782 (N_5782,N_5613,N_5585);
xor U5783 (N_5783,N_5610,N_5618);
nor U5784 (N_5784,N_5579,N_5687);
or U5785 (N_5785,N_5595,N_5607);
xor U5786 (N_5786,N_5629,N_5579);
xnor U5787 (N_5787,N_5633,N_5671);
nor U5788 (N_5788,N_5678,N_5604);
nor U5789 (N_5789,N_5595,N_5602);
xor U5790 (N_5790,N_5681,N_5642);
nor U5791 (N_5791,N_5602,N_5610);
or U5792 (N_5792,N_5552,N_5622);
or U5793 (N_5793,N_5569,N_5591);
nand U5794 (N_5794,N_5630,N_5662);
or U5795 (N_5795,N_5657,N_5595);
or U5796 (N_5796,N_5644,N_5626);
xor U5797 (N_5797,N_5590,N_5575);
nor U5798 (N_5798,N_5608,N_5665);
xor U5799 (N_5799,N_5606,N_5605);
nand U5800 (N_5800,N_5674,N_5636);
xor U5801 (N_5801,N_5638,N_5583);
or U5802 (N_5802,N_5672,N_5571);
xnor U5803 (N_5803,N_5599,N_5607);
and U5804 (N_5804,N_5665,N_5616);
or U5805 (N_5805,N_5667,N_5695);
and U5806 (N_5806,N_5693,N_5684);
or U5807 (N_5807,N_5605,N_5589);
or U5808 (N_5808,N_5583,N_5694);
nor U5809 (N_5809,N_5578,N_5568);
xnor U5810 (N_5810,N_5628,N_5662);
xnor U5811 (N_5811,N_5607,N_5561);
or U5812 (N_5812,N_5601,N_5600);
nand U5813 (N_5813,N_5621,N_5592);
nand U5814 (N_5814,N_5673,N_5672);
or U5815 (N_5815,N_5590,N_5684);
or U5816 (N_5816,N_5668,N_5648);
xnor U5817 (N_5817,N_5646,N_5615);
or U5818 (N_5818,N_5695,N_5591);
or U5819 (N_5819,N_5613,N_5557);
nor U5820 (N_5820,N_5643,N_5572);
and U5821 (N_5821,N_5648,N_5650);
and U5822 (N_5822,N_5631,N_5595);
nand U5823 (N_5823,N_5583,N_5614);
or U5824 (N_5824,N_5559,N_5582);
and U5825 (N_5825,N_5649,N_5673);
nand U5826 (N_5826,N_5659,N_5650);
nor U5827 (N_5827,N_5698,N_5596);
nand U5828 (N_5828,N_5640,N_5669);
and U5829 (N_5829,N_5623,N_5644);
xnor U5830 (N_5830,N_5666,N_5562);
nor U5831 (N_5831,N_5620,N_5696);
nand U5832 (N_5832,N_5589,N_5654);
and U5833 (N_5833,N_5567,N_5615);
nand U5834 (N_5834,N_5689,N_5675);
xnor U5835 (N_5835,N_5583,N_5570);
and U5836 (N_5836,N_5682,N_5593);
nor U5837 (N_5837,N_5679,N_5658);
xor U5838 (N_5838,N_5634,N_5569);
xnor U5839 (N_5839,N_5579,N_5697);
or U5840 (N_5840,N_5578,N_5698);
xnor U5841 (N_5841,N_5578,N_5553);
and U5842 (N_5842,N_5621,N_5579);
or U5843 (N_5843,N_5664,N_5596);
nor U5844 (N_5844,N_5616,N_5632);
nand U5845 (N_5845,N_5626,N_5658);
nand U5846 (N_5846,N_5624,N_5551);
nor U5847 (N_5847,N_5605,N_5671);
or U5848 (N_5848,N_5664,N_5665);
or U5849 (N_5849,N_5671,N_5569);
or U5850 (N_5850,N_5755,N_5711);
nand U5851 (N_5851,N_5704,N_5786);
and U5852 (N_5852,N_5835,N_5821);
or U5853 (N_5853,N_5778,N_5807);
xor U5854 (N_5854,N_5843,N_5759);
and U5855 (N_5855,N_5839,N_5790);
and U5856 (N_5856,N_5777,N_5830);
xor U5857 (N_5857,N_5770,N_5810);
nand U5858 (N_5858,N_5783,N_5825);
nor U5859 (N_5859,N_5812,N_5708);
nand U5860 (N_5860,N_5822,N_5716);
or U5861 (N_5861,N_5781,N_5706);
or U5862 (N_5862,N_5749,N_5734);
and U5863 (N_5863,N_5774,N_5717);
or U5864 (N_5864,N_5731,N_5780);
nand U5865 (N_5865,N_5827,N_5714);
nor U5866 (N_5866,N_5799,N_5802);
nor U5867 (N_5867,N_5769,N_5739);
nor U5868 (N_5868,N_5838,N_5732);
or U5869 (N_5869,N_5760,N_5744);
nand U5870 (N_5870,N_5775,N_5840);
xor U5871 (N_5871,N_5787,N_5723);
xnor U5872 (N_5872,N_5700,N_5756);
nand U5873 (N_5873,N_5779,N_5742);
or U5874 (N_5874,N_5837,N_5801);
xor U5875 (N_5875,N_5751,N_5746);
nand U5876 (N_5876,N_5727,N_5784);
xor U5877 (N_5877,N_5847,N_5710);
or U5878 (N_5878,N_5738,N_5823);
and U5879 (N_5879,N_5725,N_5792);
xnor U5880 (N_5880,N_5718,N_5720);
nor U5881 (N_5881,N_5788,N_5761);
xnor U5882 (N_5882,N_5757,N_5737);
or U5883 (N_5883,N_5809,N_5758);
xor U5884 (N_5884,N_5771,N_5848);
nor U5885 (N_5885,N_5712,N_5747);
nand U5886 (N_5886,N_5707,N_5730);
or U5887 (N_5887,N_5831,N_5733);
nor U5888 (N_5888,N_5740,N_5842);
or U5889 (N_5889,N_5805,N_5828);
nor U5890 (N_5890,N_5762,N_5798);
or U5891 (N_5891,N_5832,N_5833);
nor U5892 (N_5892,N_5763,N_5817);
xor U5893 (N_5893,N_5849,N_5819);
nor U5894 (N_5894,N_5785,N_5829);
and U5895 (N_5895,N_5841,N_5820);
nor U5896 (N_5896,N_5773,N_5818);
or U5897 (N_5897,N_5728,N_5795);
nor U5898 (N_5898,N_5709,N_5803);
and U5899 (N_5899,N_5750,N_5705);
nand U5900 (N_5900,N_5800,N_5826);
nor U5901 (N_5901,N_5844,N_5726);
xor U5902 (N_5902,N_5765,N_5845);
nor U5903 (N_5903,N_5713,N_5721);
and U5904 (N_5904,N_5702,N_5724);
or U5905 (N_5905,N_5804,N_5715);
or U5906 (N_5906,N_5793,N_5776);
nand U5907 (N_5907,N_5811,N_5736);
and U5908 (N_5908,N_5772,N_5741);
and U5909 (N_5909,N_5794,N_5796);
xnor U5910 (N_5910,N_5797,N_5754);
xor U5911 (N_5911,N_5808,N_5806);
and U5912 (N_5912,N_5766,N_5703);
xor U5913 (N_5913,N_5789,N_5722);
nor U5914 (N_5914,N_5701,N_5836);
nor U5915 (N_5915,N_5767,N_5791);
nor U5916 (N_5916,N_5824,N_5752);
xnor U5917 (N_5917,N_5815,N_5748);
xnor U5918 (N_5918,N_5846,N_5814);
nand U5919 (N_5919,N_5813,N_5753);
nand U5920 (N_5920,N_5782,N_5764);
or U5921 (N_5921,N_5719,N_5735);
nor U5922 (N_5922,N_5816,N_5834);
xor U5923 (N_5923,N_5745,N_5768);
or U5924 (N_5924,N_5743,N_5729);
and U5925 (N_5925,N_5708,N_5798);
nand U5926 (N_5926,N_5737,N_5788);
or U5927 (N_5927,N_5822,N_5846);
nor U5928 (N_5928,N_5715,N_5791);
nand U5929 (N_5929,N_5826,N_5725);
nor U5930 (N_5930,N_5746,N_5791);
or U5931 (N_5931,N_5726,N_5756);
nand U5932 (N_5932,N_5803,N_5814);
and U5933 (N_5933,N_5786,N_5785);
xor U5934 (N_5934,N_5832,N_5839);
nor U5935 (N_5935,N_5739,N_5785);
xor U5936 (N_5936,N_5739,N_5708);
or U5937 (N_5937,N_5794,N_5808);
xor U5938 (N_5938,N_5746,N_5724);
xor U5939 (N_5939,N_5723,N_5763);
nand U5940 (N_5940,N_5795,N_5721);
xnor U5941 (N_5941,N_5758,N_5723);
and U5942 (N_5942,N_5712,N_5751);
nand U5943 (N_5943,N_5807,N_5714);
nand U5944 (N_5944,N_5773,N_5739);
xor U5945 (N_5945,N_5822,N_5701);
xnor U5946 (N_5946,N_5814,N_5779);
nand U5947 (N_5947,N_5714,N_5837);
or U5948 (N_5948,N_5715,N_5833);
nand U5949 (N_5949,N_5712,N_5825);
xnor U5950 (N_5950,N_5730,N_5770);
or U5951 (N_5951,N_5750,N_5849);
and U5952 (N_5952,N_5722,N_5802);
nor U5953 (N_5953,N_5774,N_5733);
xor U5954 (N_5954,N_5829,N_5816);
nand U5955 (N_5955,N_5797,N_5778);
nand U5956 (N_5956,N_5742,N_5703);
or U5957 (N_5957,N_5788,N_5825);
and U5958 (N_5958,N_5729,N_5787);
or U5959 (N_5959,N_5735,N_5838);
xnor U5960 (N_5960,N_5784,N_5752);
nor U5961 (N_5961,N_5748,N_5769);
nor U5962 (N_5962,N_5840,N_5796);
nor U5963 (N_5963,N_5781,N_5727);
and U5964 (N_5964,N_5798,N_5838);
xnor U5965 (N_5965,N_5757,N_5835);
nor U5966 (N_5966,N_5797,N_5819);
nor U5967 (N_5967,N_5746,N_5739);
xor U5968 (N_5968,N_5763,N_5703);
and U5969 (N_5969,N_5767,N_5735);
and U5970 (N_5970,N_5740,N_5831);
xnor U5971 (N_5971,N_5740,N_5762);
or U5972 (N_5972,N_5848,N_5739);
nor U5973 (N_5973,N_5737,N_5715);
xor U5974 (N_5974,N_5841,N_5720);
or U5975 (N_5975,N_5724,N_5822);
nand U5976 (N_5976,N_5747,N_5725);
and U5977 (N_5977,N_5793,N_5771);
nand U5978 (N_5978,N_5839,N_5824);
nand U5979 (N_5979,N_5728,N_5734);
nand U5980 (N_5980,N_5736,N_5750);
nor U5981 (N_5981,N_5701,N_5833);
nor U5982 (N_5982,N_5840,N_5713);
or U5983 (N_5983,N_5797,N_5776);
and U5984 (N_5984,N_5820,N_5762);
nor U5985 (N_5985,N_5716,N_5825);
xor U5986 (N_5986,N_5701,N_5831);
or U5987 (N_5987,N_5843,N_5839);
nor U5988 (N_5988,N_5731,N_5773);
and U5989 (N_5989,N_5797,N_5826);
nor U5990 (N_5990,N_5734,N_5808);
and U5991 (N_5991,N_5836,N_5828);
nor U5992 (N_5992,N_5773,N_5830);
nand U5993 (N_5993,N_5794,N_5795);
and U5994 (N_5994,N_5836,N_5783);
nor U5995 (N_5995,N_5804,N_5727);
nor U5996 (N_5996,N_5791,N_5706);
or U5997 (N_5997,N_5841,N_5717);
and U5998 (N_5998,N_5842,N_5737);
or U5999 (N_5999,N_5822,N_5730);
nand U6000 (N_6000,N_5956,N_5987);
nor U6001 (N_6001,N_5876,N_5861);
xor U6002 (N_6002,N_5863,N_5933);
xor U6003 (N_6003,N_5955,N_5961);
nor U6004 (N_6004,N_5874,N_5879);
and U6005 (N_6005,N_5860,N_5964);
or U6006 (N_6006,N_5993,N_5897);
or U6007 (N_6007,N_5908,N_5853);
or U6008 (N_6008,N_5982,N_5969);
nand U6009 (N_6009,N_5980,N_5923);
xnor U6010 (N_6010,N_5957,N_5951);
and U6011 (N_6011,N_5972,N_5864);
xor U6012 (N_6012,N_5910,N_5890);
nor U6013 (N_6013,N_5950,N_5939);
xor U6014 (N_6014,N_5998,N_5871);
nor U6015 (N_6015,N_5936,N_5935);
nand U6016 (N_6016,N_5938,N_5919);
or U6017 (N_6017,N_5883,N_5959);
nor U6018 (N_6018,N_5877,N_5967);
nor U6019 (N_6019,N_5970,N_5926);
xnor U6020 (N_6020,N_5988,N_5995);
or U6021 (N_6021,N_5997,N_5892);
and U6022 (N_6022,N_5905,N_5893);
xor U6023 (N_6023,N_5852,N_5940);
xor U6024 (N_6024,N_5963,N_5889);
nand U6025 (N_6025,N_5986,N_5896);
and U6026 (N_6026,N_5992,N_5953);
nor U6027 (N_6027,N_5882,N_5932);
and U6028 (N_6028,N_5968,N_5880);
and U6029 (N_6029,N_5974,N_5927);
nor U6030 (N_6030,N_5952,N_5913);
or U6031 (N_6031,N_5916,N_5925);
xor U6032 (N_6032,N_5887,N_5920);
nor U6033 (N_6033,N_5917,N_5903);
nor U6034 (N_6034,N_5898,N_5949);
nand U6035 (N_6035,N_5991,N_5958);
or U6036 (N_6036,N_5895,N_5945);
or U6037 (N_6037,N_5884,N_5858);
nor U6038 (N_6038,N_5866,N_5878);
nor U6039 (N_6039,N_5891,N_5946);
xor U6040 (N_6040,N_5869,N_5990);
and U6041 (N_6041,N_5973,N_5904);
or U6042 (N_6042,N_5962,N_5901);
xor U6043 (N_6043,N_5921,N_5981);
or U6044 (N_6044,N_5965,N_5999);
or U6045 (N_6045,N_5977,N_5954);
and U6046 (N_6046,N_5931,N_5859);
nand U6047 (N_6047,N_5865,N_5857);
nand U6048 (N_6048,N_5856,N_5914);
or U6049 (N_6049,N_5907,N_5886);
nor U6050 (N_6050,N_5875,N_5996);
nor U6051 (N_6051,N_5985,N_5984);
xor U6052 (N_6052,N_5888,N_5976);
nand U6053 (N_6053,N_5943,N_5922);
xor U6054 (N_6054,N_5947,N_5934);
xnor U6055 (N_6055,N_5944,N_5937);
and U6056 (N_6056,N_5912,N_5911);
xnor U6057 (N_6057,N_5924,N_5930);
nand U6058 (N_6058,N_5885,N_5900);
or U6059 (N_6059,N_5971,N_5862);
or U6060 (N_6060,N_5918,N_5979);
nor U6061 (N_6061,N_5854,N_5989);
or U6062 (N_6062,N_5941,N_5942);
and U6063 (N_6063,N_5966,N_5899);
or U6064 (N_6064,N_5870,N_5928);
and U6065 (N_6065,N_5872,N_5868);
nand U6066 (N_6066,N_5855,N_5929);
xor U6067 (N_6067,N_5873,N_5975);
nor U6068 (N_6068,N_5948,N_5983);
nor U6069 (N_6069,N_5915,N_5851);
xor U6070 (N_6070,N_5978,N_5894);
nor U6071 (N_6071,N_5909,N_5902);
or U6072 (N_6072,N_5867,N_5994);
xnor U6073 (N_6073,N_5881,N_5960);
and U6074 (N_6074,N_5906,N_5850);
and U6075 (N_6075,N_5978,N_5997);
xnor U6076 (N_6076,N_5927,N_5855);
nor U6077 (N_6077,N_5975,N_5856);
nor U6078 (N_6078,N_5876,N_5901);
and U6079 (N_6079,N_5974,N_5967);
and U6080 (N_6080,N_5867,N_5956);
and U6081 (N_6081,N_5938,N_5892);
or U6082 (N_6082,N_5869,N_5889);
nor U6083 (N_6083,N_5949,N_5897);
or U6084 (N_6084,N_5939,N_5871);
and U6085 (N_6085,N_5881,N_5909);
or U6086 (N_6086,N_5881,N_5930);
and U6087 (N_6087,N_5963,N_5888);
and U6088 (N_6088,N_5903,N_5864);
or U6089 (N_6089,N_5851,N_5964);
nor U6090 (N_6090,N_5944,N_5918);
or U6091 (N_6091,N_5986,N_5939);
and U6092 (N_6092,N_5992,N_5853);
and U6093 (N_6093,N_5976,N_5991);
nor U6094 (N_6094,N_5860,N_5952);
xnor U6095 (N_6095,N_5887,N_5879);
nand U6096 (N_6096,N_5862,N_5852);
nand U6097 (N_6097,N_5917,N_5895);
nand U6098 (N_6098,N_5993,N_5982);
nor U6099 (N_6099,N_5859,N_5908);
and U6100 (N_6100,N_5891,N_5982);
nor U6101 (N_6101,N_5857,N_5980);
or U6102 (N_6102,N_5959,N_5926);
and U6103 (N_6103,N_5880,N_5928);
or U6104 (N_6104,N_5978,N_5930);
and U6105 (N_6105,N_5931,N_5951);
and U6106 (N_6106,N_5924,N_5852);
xnor U6107 (N_6107,N_5873,N_5988);
nand U6108 (N_6108,N_5926,N_5982);
xnor U6109 (N_6109,N_5901,N_5930);
or U6110 (N_6110,N_5945,N_5927);
or U6111 (N_6111,N_5864,N_5865);
nand U6112 (N_6112,N_5898,N_5972);
and U6113 (N_6113,N_5853,N_5902);
and U6114 (N_6114,N_5999,N_5864);
or U6115 (N_6115,N_5926,N_5921);
nand U6116 (N_6116,N_5946,N_5856);
nand U6117 (N_6117,N_5884,N_5971);
and U6118 (N_6118,N_5982,N_5995);
or U6119 (N_6119,N_5979,N_5854);
nand U6120 (N_6120,N_5862,N_5937);
xor U6121 (N_6121,N_5954,N_5945);
or U6122 (N_6122,N_5961,N_5902);
nand U6123 (N_6123,N_5880,N_5865);
or U6124 (N_6124,N_5932,N_5919);
or U6125 (N_6125,N_5982,N_5894);
xor U6126 (N_6126,N_5873,N_5872);
nor U6127 (N_6127,N_5995,N_5884);
and U6128 (N_6128,N_5889,N_5890);
nand U6129 (N_6129,N_5929,N_5859);
and U6130 (N_6130,N_5971,N_5986);
nand U6131 (N_6131,N_5954,N_5872);
or U6132 (N_6132,N_5928,N_5915);
xnor U6133 (N_6133,N_5881,N_5890);
and U6134 (N_6134,N_5899,N_5859);
xor U6135 (N_6135,N_5927,N_5978);
nand U6136 (N_6136,N_5871,N_5968);
nor U6137 (N_6137,N_5853,N_5976);
and U6138 (N_6138,N_5949,N_5880);
or U6139 (N_6139,N_5918,N_5907);
nand U6140 (N_6140,N_5963,N_5972);
and U6141 (N_6141,N_5906,N_5928);
nand U6142 (N_6142,N_5934,N_5925);
nand U6143 (N_6143,N_5852,N_5958);
xnor U6144 (N_6144,N_5864,N_5943);
nor U6145 (N_6145,N_5923,N_5979);
nand U6146 (N_6146,N_5963,N_5857);
xor U6147 (N_6147,N_5936,N_5874);
nand U6148 (N_6148,N_5949,N_5999);
and U6149 (N_6149,N_5854,N_5868);
or U6150 (N_6150,N_6086,N_6141);
nand U6151 (N_6151,N_6139,N_6022);
nand U6152 (N_6152,N_6008,N_6060);
xnor U6153 (N_6153,N_6013,N_6084);
xnor U6154 (N_6154,N_6029,N_6078);
or U6155 (N_6155,N_6127,N_6074);
and U6156 (N_6156,N_6148,N_6128);
and U6157 (N_6157,N_6147,N_6050);
nand U6158 (N_6158,N_6001,N_6063);
nand U6159 (N_6159,N_6077,N_6027);
nor U6160 (N_6160,N_6107,N_6024);
or U6161 (N_6161,N_6087,N_6104);
or U6162 (N_6162,N_6116,N_6061);
nor U6163 (N_6163,N_6134,N_6059);
nand U6164 (N_6164,N_6085,N_6123);
nor U6165 (N_6165,N_6032,N_6064);
nor U6166 (N_6166,N_6144,N_6115);
nand U6167 (N_6167,N_6025,N_6091);
nand U6168 (N_6168,N_6038,N_6011);
nand U6169 (N_6169,N_6018,N_6037);
nor U6170 (N_6170,N_6019,N_6045);
xor U6171 (N_6171,N_6121,N_6145);
xor U6172 (N_6172,N_6017,N_6110);
nor U6173 (N_6173,N_6143,N_6092);
nand U6174 (N_6174,N_6075,N_6146);
xor U6175 (N_6175,N_6015,N_6020);
xnor U6176 (N_6176,N_6080,N_6002);
and U6177 (N_6177,N_6126,N_6014);
nand U6178 (N_6178,N_6136,N_6108);
and U6179 (N_6179,N_6124,N_6065);
or U6180 (N_6180,N_6125,N_6140);
or U6181 (N_6181,N_6119,N_6000);
xor U6182 (N_6182,N_6005,N_6113);
nand U6183 (N_6183,N_6109,N_6047);
nor U6184 (N_6184,N_6102,N_6082);
nor U6185 (N_6185,N_6030,N_6057);
nor U6186 (N_6186,N_6056,N_6135);
xnor U6187 (N_6187,N_6073,N_6111);
xnor U6188 (N_6188,N_6049,N_6081);
nand U6189 (N_6189,N_6048,N_6122);
and U6190 (N_6190,N_6021,N_6043);
nor U6191 (N_6191,N_6079,N_6106);
or U6192 (N_6192,N_6114,N_6099);
xnor U6193 (N_6193,N_6129,N_6023);
and U6194 (N_6194,N_6066,N_6137);
nor U6195 (N_6195,N_6009,N_6036);
and U6196 (N_6196,N_6062,N_6040);
nor U6197 (N_6197,N_6101,N_6097);
nand U6198 (N_6198,N_6031,N_6133);
and U6199 (N_6199,N_6051,N_6131);
nor U6200 (N_6200,N_6090,N_6069);
and U6201 (N_6201,N_6055,N_6012);
nand U6202 (N_6202,N_6072,N_6076);
xor U6203 (N_6203,N_6026,N_6028);
or U6204 (N_6204,N_6041,N_6089);
nor U6205 (N_6205,N_6006,N_6120);
nor U6206 (N_6206,N_6033,N_6004);
xor U6207 (N_6207,N_6067,N_6034);
or U6208 (N_6208,N_6096,N_6118);
or U6209 (N_6209,N_6095,N_6044);
xor U6210 (N_6210,N_6088,N_6100);
xnor U6211 (N_6211,N_6070,N_6035);
xor U6212 (N_6212,N_6039,N_6053);
xor U6213 (N_6213,N_6052,N_6149);
and U6214 (N_6214,N_6003,N_6083);
and U6215 (N_6215,N_6117,N_6103);
or U6216 (N_6216,N_6098,N_6016);
and U6217 (N_6217,N_6058,N_6010);
nand U6218 (N_6218,N_6112,N_6054);
nand U6219 (N_6219,N_6093,N_6105);
or U6220 (N_6220,N_6071,N_6046);
and U6221 (N_6221,N_6068,N_6130);
nand U6222 (N_6222,N_6094,N_6007);
or U6223 (N_6223,N_6042,N_6142);
nor U6224 (N_6224,N_6138,N_6132);
nand U6225 (N_6225,N_6111,N_6084);
and U6226 (N_6226,N_6119,N_6031);
nor U6227 (N_6227,N_6077,N_6000);
or U6228 (N_6228,N_6110,N_6034);
xor U6229 (N_6229,N_6110,N_6096);
nor U6230 (N_6230,N_6136,N_6133);
xor U6231 (N_6231,N_6065,N_6136);
and U6232 (N_6232,N_6024,N_6006);
nor U6233 (N_6233,N_6098,N_6053);
nand U6234 (N_6234,N_6045,N_6076);
xor U6235 (N_6235,N_6012,N_6073);
nand U6236 (N_6236,N_6094,N_6095);
nor U6237 (N_6237,N_6147,N_6142);
or U6238 (N_6238,N_6024,N_6026);
nand U6239 (N_6239,N_6117,N_6115);
nor U6240 (N_6240,N_6035,N_6059);
and U6241 (N_6241,N_6080,N_6069);
xor U6242 (N_6242,N_6054,N_6130);
nand U6243 (N_6243,N_6017,N_6024);
nor U6244 (N_6244,N_6108,N_6011);
and U6245 (N_6245,N_6061,N_6052);
and U6246 (N_6246,N_6016,N_6103);
nor U6247 (N_6247,N_6110,N_6086);
nand U6248 (N_6248,N_6143,N_6072);
nand U6249 (N_6249,N_6017,N_6087);
xor U6250 (N_6250,N_6066,N_6075);
xnor U6251 (N_6251,N_6127,N_6080);
nor U6252 (N_6252,N_6076,N_6111);
or U6253 (N_6253,N_6079,N_6116);
or U6254 (N_6254,N_6010,N_6147);
nand U6255 (N_6255,N_6107,N_6127);
xnor U6256 (N_6256,N_6142,N_6109);
xor U6257 (N_6257,N_6097,N_6048);
nand U6258 (N_6258,N_6107,N_6081);
or U6259 (N_6259,N_6052,N_6146);
nand U6260 (N_6260,N_6137,N_6064);
or U6261 (N_6261,N_6112,N_6001);
nand U6262 (N_6262,N_6077,N_6057);
and U6263 (N_6263,N_6020,N_6011);
and U6264 (N_6264,N_6012,N_6071);
nand U6265 (N_6265,N_6005,N_6079);
nor U6266 (N_6266,N_6066,N_6045);
nor U6267 (N_6267,N_6082,N_6149);
and U6268 (N_6268,N_6022,N_6146);
or U6269 (N_6269,N_6116,N_6005);
or U6270 (N_6270,N_6038,N_6025);
or U6271 (N_6271,N_6087,N_6113);
or U6272 (N_6272,N_6036,N_6078);
nand U6273 (N_6273,N_6102,N_6145);
nor U6274 (N_6274,N_6002,N_6101);
nor U6275 (N_6275,N_6006,N_6095);
xnor U6276 (N_6276,N_6007,N_6067);
nand U6277 (N_6277,N_6036,N_6020);
xnor U6278 (N_6278,N_6144,N_6080);
nor U6279 (N_6279,N_6041,N_6021);
xnor U6280 (N_6280,N_6141,N_6119);
xor U6281 (N_6281,N_6096,N_6089);
and U6282 (N_6282,N_6096,N_6067);
xor U6283 (N_6283,N_6051,N_6070);
nand U6284 (N_6284,N_6081,N_6054);
and U6285 (N_6285,N_6001,N_6088);
and U6286 (N_6286,N_6085,N_6087);
nand U6287 (N_6287,N_6065,N_6106);
nor U6288 (N_6288,N_6043,N_6088);
and U6289 (N_6289,N_6104,N_6139);
and U6290 (N_6290,N_6027,N_6055);
xnor U6291 (N_6291,N_6087,N_6137);
xor U6292 (N_6292,N_6126,N_6145);
xnor U6293 (N_6293,N_6107,N_6079);
xnor U6294 (N_6294,N_6012,N_6095);
and U6295 (N_6295,N_6092,N_6064);
or U6296 (N_6296,N_6097,N_6148);
nor U6297 (N_6297,N_6120,N_6009);
nand U6298 (N_6298,N_6065,N_6024);
xor U6299 (N_6299,N_6095,N_6144);
xnor U6300 (N_6300,N_6196,N_6162);
and U6301 (N_6301,N_6284,N_6237);
or U6302 (N_6302,N_6199,N_6168);
nand U6303 (N_6303,N_6205,N_6202);
xor U6304 (N_6304,N_6281,N_6183);
or U6305 (N_6305,N_6169,N_6298);
or U6306 (N_6306,N_6152,N_6194);
or U6307 (N_6307,N_6246,N_6158);
nor U6308 (N_6308,N_6193,N_6242);
xor U6309 (N_6309,N_6247,N_6201);
xnor U6310 (N_6310,N_6186,N_6155);
xnor U6311 (N_6311,N_6195,N_6189);
or U6312 (N_6312,N_6211,N_6192);
nor U6313 (N_6313,N_6200,N_6204);
nand U6314 (N_6314,N_6157,N_6160);
nor U6315 (N_6315,N_6236,N_6198);
xnor U6316 (N_6316,N_6280,N_6165);
nor U6317 (N_6317,N_6170,N_6271);
nand U6318 (N_6318,N_6154,N_6219);
nor U6319 (N_6319,N_6248,N_6258);
xnor U6320 (N_6320,N_6164,N_6185);
nand U6321 (N_6321,N_6207,N_6151);
and U6322 (N_6322,N_6214,N_6288);
nor U6323 (N_6323,N_6188,N_6282);
or U6324 (N_6324,N_6159,N_6269);
or U6325 (N_6325,N_6230,N_6239);
nor U6326 (N_6326,N_6263,N_6212);
nor U6327 (N_6327,N_6297,N_6249);
nand U6328 (N_6328,N_6245,N_6291);
or U6329 (N_6329,N_6265,N_6178);
or U6330 (N_6330,N_6250,N_6289);
nand U6331 (N_6331,N_6283,N_6233);
nand U6332 (N_6332,N_6187,N_6272);
or U6333 (N_6333,N_6213,N_6163);
nand U6334 (N_6334,N_6238,N_6203);
nand U6335 (N_6335,N_6252,N_6228);
nand U6336 (N_6336,N_6270,N_6267);
xnor U6337 (N_6337,N_6278,N_6275);
or U6338 (N_6338,N_6184,N_6177);
or U6339 (N_6339,N_6197,N_6251);
xor U6340 (N_6340,N_6217,N_6277);
or U6341 (N_6341,N_6156,N_6166);
xnor U6342 (N_6342,N_6231,N_6174);
nand U6343 (N_6343,N_6215,N_6286);
nor U6344 (N_6344,N_6191,N_6181);
nand U6345 (N_6345,N_6257,N_6222);
xnor U6346 (N_6346,N_6167,N_6253);
nand U6347 (N_6347,N_6210,N_6235);
nor U6348 (N_6348,N_6226,N_6216);
and U6349 (N_6349,N_6227,N_6273);
nor U6350 (N_6350,N_6206,N_6264);
nand U6351 (N_6351,N_6223,N_6287);
nand U6352 (N_6352,N_6285,N_6268);
nand U6353 (N_6353,N_6290,N_6292);
and U6354 (N_6354,N_6161,N_6294);
nor U6355 (N_6355,N_6209,N_6240);
nand U6356 (N_6356,N_6175,N_6232);
and U6357 (N_6357,N_6299,N_6182);
nor U6358 (N_6358,N_6179,N_6279);
nand U6359 (N_6359,N_6255,N_6244);
or U6360 (N_6360,N_6234,N_6153);
xor U6361 (N_6361,N_6266,N_6261);
and U6362 (N_6362,N_6262,N_6208);
or U6363 (N_6363,N_6180,N_6173);
nand U6364 (N_6364,N_6224,N_6176);
nor U6365 (N_6365,N_6260,N_6171);
xor U6366 (N_6366,N_6293,N_6229);
or U6367 (N_6367,N_6254,N_6172);
nand U6368 (N_6368,N_6221,N_6256);
or U6369 (N_6369,N_6241,N_6150);
nand U6370 (N_6370,N_6218,N_6295);
xor U6371 (N_6371,N_6259,N_6276);
nand U6372 (N_6372,N_6296,N_6243);
nor U6373 (N_6373,N_6225,N_6220);
and U6374 (N_6374,N_6190,N_6274);
and U6375 (N_6375,N_6152,N_6267);
or U6376 (N_6376,N_6260,N_6170);
nand U6377 (N_6377,N_6237,N_6233);
nor U6378 (N_6378,N_6214,N_6276);
or U6379 (N_6379,N_6242,N_6284);
nand U6380 (N_6380,N_6280,N_6237);
xor U6381 (N_6381,N_6290,N_6163);
or U6382 (N_6382,N_6263,N_6202);
or U6383 (N_6383,N_6216,N_6274);
and U6384 (N_6384,N_6172,N_6228);
or U6385 (N_6385,N_6178,N_6190);
nand U6386 (N_6386,N_6152,N_6243);
nand U6387 (N_6387,N_6159,N_6299);
or U6388 (N_6388,N_6162,N_6269);
and U6389 (N_6389,N_6249,N_6191);
xnor U6390 (N_6390,N_6152,N_6232);
nand U6391 (N_6391,N_6290,N_6239);
xnor U6392 (N_6392,N_6186,N_6152);
and U6393 (N_6393,N_6254,N_6288);
and U6394 (N_6394,N_6224,N_6218);
xor U6395 (N_6395,N_6237,N_6246);
or U6396 (N_6396,N_6183,N_6227);
and U6397 (N_6397,N_6232,N_6297);
xnor U6398 (N_6398,N_6202,N_6172);
and U6399 (N_6399,N_6229,N_6239);
nor U6400 (N_6400,N_6292,N_6203);
nor U6401 (N_6401,N_6293,N_6169);
nand U6402 (N_6402,N_6154,N_6173);
nand U6403 (N_6403,N_6190,N_6219);
nor U6404 (N_6404,N_6256,N_6162);
or U6405 (N_6405,N_6158,N_6195);
nor U6406 (N_6406,N_6154,N_6194);
nand U6407 (N_6407,N_6255,N_6226);
and U6408 (N_6408,N_6297,N_6286);
nand U6409 (N_6409,N_6211,N_6190);
nand U6410 (N_6410,N_6241,N_6193);
nor U6411 (N_6411,N_6245,N_6223);
nor U6412 (N_6412,N_6239,N_6222);
and U6413 (N_6413,N_6213,N_6188);
xor U6414 (N_6414,N_6175,N_6285);
xnor U6415 (N_6415,N_6240,N_6289);
or U6416 (N_6416,N_6268,N_6265);
and U6417 (N_6417,N_6228,N_6285);
nor U6418 (N_6418,N_6156,N_6173);
or U6419 (N_6419,N_6174,N_6186);
xnor U6420 (N_6420,N_6165,N_6268);
xnor U6421 (N_6421,N_6219,N_6188);
and U6422 (N_6422,N_6298,N_6280);
nand U6423 (N_6423,N_6215,N_6172);
and U6424 (N_6424,N_6222,N_6275);
and U6425 (N_6425,N_6157,N_6273);
and U6426 (N_6426,N_6188,N_6226);
or U6427 (N_6427,N_6264,N_6275);
nand U6428 (N_6428,N_6183,N_6240);
and U6429 (N_6429,N_6180,N_6193);
or U6430 (N_6430,N_6271,N_6220);
nand U6431 (N_6431,N_6169,N_6252);
xnor U6432 (N_6432,N_6289,N_6202);
nor U6433 (N_6433,N_6156,N_6263);
xnor U6434 (N_6434,N_6279,N_6224);
nor U6435 (N_6435,N_6247,N_6274);
xnor U6436 (N_6436,N_6188,N_6298);
or U6437 (N_6437,N_6277,N_6264);
xnor U6438 (N_6438,N_6190,N_6285);
xnor U6439 (N_6439,N_6222,N_6195);
and U6440 (N_6440,N_6290,N_6255);
nand U6441 (N_6441,N_6289,N_6230);
nand U6442 (N_6442,N_6285,N_6214);
nor U6443 (N_6443,N_6293,N_6172);
xnor U6444 (N_6444,N_6187,N_6260);
and U6445 (N_6445,N_6282,N_6296);
or U6446 (N_6446,N_6187,N_6170);
and U6447 (N_6447,N_6244,N_6204);
nand U6448 (N_6448,N_6265,N_6215);
and U6449 (N_6449,N_6237,N_6188);
nor U6450 (N_6450,N_6335,N_6300);
nand U6451 (N_6451,N_6395,N_6362);
xor U6452 (N_6452,N_6429,N_6449);
xnor U6453 (N_6453,N_6319,N_6308);
or U6454 (N_6454,N_6415,N_6385);
or U6455 (N_6455,N_6371,N_6320);
nand U6456 (N_6456,N_6398,N_6324);
or U6457 (N_6457,N_6364,N_6427);
xnor U6458 (N_6458,N_6367,N_6348);
or U6459 (N_6459,N_6325,N_6376);
xor U6460 (N_6460,N_6387,N_6379);
or U6461 (N_6461,N_6309,N_6377);
xor U6462 (N_6462,N_6322,N_6421);
nor U6463 (N_6463,N_6444,N_6321);
nand U6464 (N_6464,N_6368,N_6436);
nand U6465 (N_6465,N_6359,N_6346);
and U6466 (N_6466,N_6396,N_6326);
nor U6467 (N_6467,N_6327,N_6307);
or U6468 (N_6468,N_6388,N_6406);
xor U6469 (N_6469,N_6407,N_6412);
xor U6470 (N_6470,N_6373,N_6446);
or U6471 (N_6471,N_6392,N_6363);
and U6472 (N_6472,N_6370,N_6329);
or U6473 (N_6473,N_6411,N_6357);
nand U6474 (N_6474,N_6426,N_6419);
nand U6475 (N_6475,N_6410,N_6440);
nor U6476 (N_6476,N_6380,N_6397);
or U6477 (N_6477,N_6369,N_6312);
nand U6478 (N_6478,N_6349,N_6438);
and U6479 (N_6479,N_6418,N_6340);
nor U6480 (N_6480,N_6422,N_6430);
xnor U6481 (N_6481,N_6304,N_6400);
xor U6482 (N_6482,N_6434,N_6323);
nand U6483 (N_6483,N_6442,N_6414);
xnor U6484 (N_6484,N_6334,N_6336);
and U6485 (N_6485,N_6306,N_6404);
nor U6486 (N_6486,N_6409,N_6361);
and U6487 (N_6487,N_6330,N_6445);
and U6488 (N_6488,N_6352,N_6317);
or U6489 (N_6489,N_6332,N_6435);
or U6490 (N_6490,N_6439,N_6358);
and U6491 (N_6491,N_6420,N_6428);
nand U6492 (N_6492,N_6303,N_6337);
nand U6493 (N_6493,N_6351,N_6313);
or U6494 (N_6494,N_6356,N_6338);
and U6495 (N_6495,N_6375,N_6353);
nand U6496 (N_6496,N_6433,N_6347);
nor U6497 (N_6497,N_6417,N_6350);
nand U6498 (N_6498,N_6399,N_6394);
nor U6499 (N_6499,N_6447,N_6432);
or U6500 (N_6500,N_6372,N_6443);
nand U6501 (N_6501,N_6402,N_6384);
xor U6502 (N_6502,N_6355,N_6448);
or U6503 (N_6503,N_6301,N_6378);
or U6504 (N_6504,N_6314,N_6344);
or U6505 (N_6505,N_6310,N_6343);
or U6506 (N_6506,N_6366,N_6423);
xnor U6507 (N_6507,N_6305,N_6437);
nor U6508 (N_6508,N_6393,N_6431);
nand U6509 (N_6509,N_6381,N_6386);
or U6510 (N_6510,N_6413,N_6341);
nor U6511 (N_6511,N_6382,N_6333);
nor U6512 (N_6512,N_6408,N_6401);
nand U6513 (N_6513,N_6405,N_6315);
and U6514 (N_6514,N_6441,N_6389);
and U6515 (N_6515,N_6374,N_6342);
and U6516 (N_6516,N_6316,N_6360);
or U6517 (N_6517,N_6390,N_6302);
nand U6518 (N_6518,N_6345,N_6339);
or U6519 (N_6519,N_6331,N_6403);
and U6520 (N_6520,N_6318,N_6328);
and U6521 (N_6521,N_6311,N_6383);
xnor U6522 (N_6522,N_6354,N_6424);
nor U6523 (N_6523,N_6416,N_6391);
and U6524 (N_6524,N_6425,N_6365);
and U6525 (N_6525,N_6362,N_6410);
and U6526 (N_6526,N_6345,N_6443);
nor U6527 (N_6527,N_6432,N_6423);
nand U6528 (N_6528,N_6410,N_6431);
nor U6529 (N_6529,N_6300,N_6429);
or U6530 (N_6530,N_6440,N_6347);
nor U6531 (N_6531,N_6307,N_6410);
nand U6532 (N_6532,N_6357,N_6309);
xnor U6533 (N_6533,N_6442,N_6333);
xnor U6534 (N_6534,N_6330,N_6331);
nor U6535 (N_6535,N_6428,N_6427);
xor U6536 (N_6536,N_6375,N_6384);
nor U6537 (N_6537,N_6415,N_6315);
xnor U6538 (N_6538,N_6348,N_6392);
nor U6539 (N_6539,N_6313,N_6408);
xnor U6540 (N_6540,N_6303,N_6328);
xor U6541 (N_6541,N_6349,N_6319);
or U6542 (N_6542,N_6427,N_6329);
xnor U6543 (N_6543,N_6407,N_6437);
and U6544 (N_6544,N_6323,N_6320);
or U6545 (N_6545,N_6365,N_6338);
and U6546 (N_6546,N_6333,N_6322);
nand U6547 (N_6547,N_6329,N_6351);
and U6548 (N_6548,N_6403,N_6394);
and U6549 (N_6549,N_6433,N_6317);
or U6550 (N_6550,N_6330,N_6361);
nand U6551 (N_6551,N_6445,N_6426);
xor U6552 (N_6552,N_6417,N_6418);
or U6553 (N_6553,N_6399,N_6358);
and U6554 (N_6554,N_6364,N_6330);
xor U6555 (N_6555,N_6421,N_6354);
nor U6556 (N_6556,N_6326,N_6338);
or U6557 (N_6557,N_6311,N_6338);
xnor U6558 (N_6558,N_6341,N_6302);
and U6559 (N_6559,N_6355,N_6319);
nand U6560 (N_6560,N_6334,N_6343);
nor U6561 (N_6561,N_6445,N_6344);
nand U6562 (N_6562,N_6381,N_6378);
and U6563 (N_6563,N_6304,N_6377);
nand U6564 (N_6564,N_6421,N_6383);
nor U6565 (N_6565,N_6310,N_6420);
nand U6566 (N_6566,N_6341,N_6433);
or U6567 (N_6567,N_6303,N_6389);
nand U6568 (N_6568,N_6350,N_6442);
nand U6569 (N_6569,N_6323,N_6316);
nand U6570 (N_6570,N_6334,N_6403);
or U6571 (N_6571,N_6428,N_6405);
nand U6572 (N_6572,N_6323,N_6346);
and U6573 (N_6573,N_6347,N_6310);
and U6574 (N_6574,N_6441,N_6438);
nor U6575 (N_6575,N_6371,N_6337);
xor U6576 (N_6576,N_6388,N_6448);
and U6577 (N_6577,N_6423,N_6354);
and U6578 (N_6578,N_6342,N_6419);
or U6579 (N_6579,N_6380,N_6369);
nand U6580 (N_6580,N_6301,N_6334);
nor U6581 (N_6581,N_6409,N_6423);
and U6582 (N_6582,N_6448,N_6441);
nand U6583 (N_6583,N_6444,N_6341);
nor U6584 (N_6584,N_6412,N_6328);
nand U6585 (N_6585,N_6348,N_6382);
and U6586 (N_6586,N_6318,N_6402);
nand U6587 (N_6587,N_6382,N_6376);
nand U6588 (N_6588,N_6447,N_6442);
and U6589 (N_6589,N_6307,N_6360);
and U6590 (N_6590,N_6410,N_6438);
nand U6591 (N_6591,N_6328,N_6447);
nand U6592 (N_6592,N_6389,N_6369);
or U6593 (N_6593,N_6390,N_6377);
or U6594 (N_6594,N_6402,N_6410);
and U6595 (N_6595,N_6373,N_6308);
nand U6596 (N_6596,N_6326,N_6413);
xnor U6597 (N_6597,N_6398,N_6341);
or U6598 (N_6598,N_6301,N_6380);
nor U6599 (N_6599,N_6301,N_6436);
nor U6600 (N_6600,N_6563,N_6452);
nand U6601 (N_6601,N_6463,N_6591);
xnor U6602 (N_6602,N_6468,N_6450);
nand U6603 (N_6603,N_6571,N_6540);
nor U6604 (N_6604,N_6576,N_6597);
or U6605 (N_6605,N_6475,N_6530);
or U6606 (N_6606,N_6471,N_6488);
or U6607 (N_6607,N_6529,N_6541);
nor U6608 (N_6608,N_6506,N_6596);
xnor U6609 (N_6609,N_6500,N_6570);
or U6610 (N_6610,N_6536,N_6589);
and U6611 (N_6611,N_6521,N_6509);
and U6612 (N_6612,N_6501,N_6527);
nor U6613 (N_6613,N_6533,N_6556);
nand U6614 (N_6614,N_6535,N_6551);
nor U6615 (N_6615,N_6542,N_6557);
nor U6616 (N_6616,N_6507,N_6487);
and U6617 (N_6617,N_6510,N_6553);
and U6618 (N_6618,N_6577,N_6537);
nand U6619 (N_6619,N_6550,N_6493);
and U6620 (N_6620,N_6465,N_6512);
nor U6621 (N_6621,N_6593,N_6528);
and U6622 (N_6622,N_6584,N_6534);
and U6623 (N_6623,N_6595,N_6484);
and U6624 (N_6624,N_6573,N_6594);
xnor U6625 (N_6625,N_6492,N_6472);
or U6626 (N_6626,N_6517,N_6579);
nand U6627 (N_6627,N_6564,N_6457);
nand U6628 (N_6628,N_6590,N_6532);
and U6629 (N_6629,N_6522,N_6474);
nor U6630 (N_6630,N_6453,N_6515);
nand U6631 (N_6631,N_6552,N_6505);
xnor U6632 (N_6632,N_6466,N_6524);
and U6633 (N_6633,N_6566,N_6572);
or U6634 (N_6634,N_6498,N_6479);
and U6635 (N_6635,N_6481,N_6544);
xnor U6636 (N_6636,N_6461,N_6587);
or U6637 (N_6637,N_6539,N_6519);
or U6638 (N_6638,N_6495,N_6555);
or U6639 (N_6639,N_6531,N_6546);
or U6640 (N_6640,N_6559,N_6562);
xnor U6641 (N_6641,N_6508,N_6459);
or U6642 (N_6642,N_6489,N_6494);
or U6643 (N_6643,N_6458,N_6480);
nor U6644 (N_6644,N_6514,N_6598);
and U6645 (N_6645,N_6526,N_6538);
nor U6646 (N_6646,N_6574,N_6588);
xor U6647 (N_6647,N_6568,N_6520);
or U6648 (N_6648,N_6513,N_6560);
or U6649 (N_6649,N_6511,N_6516);
nand U6650 (N_6650,N_6580,N_6578);
nand U6651 (N_6651,N_6473,N_6464);
or U6652 (N_6652,N_6518,N_6499);
nand U6653 (N_6653,N_6460,N_6558);
and U6654 (N_6654,N_6502,N_6454);
nor U6655 (N_6655,N_6467,N_6575);
nand U6656 (N_6656,N_6490,N_6485);
or U6657 (N_6657,N_6496,N_6470);
nor U6658 (N_6658,N_6581,N_6585);
nand U6659 (N_6659,N_6525,N_6455);
xnor U6660 (N_6660,N_6547,N_6476);
nand U6661 (N_6661,N_6451,N_6486);
nor U6662 (N_6662,N_6462,N_6478);
nor U6663 (N_6663,N_6523,N_6545);
and U6664 (N_6664,N_6482,N_6565);
nand U6665 (N_6665,N_6456,N_6583);
nand U6666 (N_6666,N_6504,N_6497);
and U6667 (N_6667,N_6548,N_6477);
nor U6668 (N_6668,N_6592,N_6491);
nand U6669 (N_6669,N_6586,N_6567);
nor U6670 (N_6670,N_6599,N_6469);
or U6671 (N_6671,N_6582,N_6503);
nand U6672 (N_6672,N_6549,N_6554);
nand U6673 (N_6673,N_6561,N_6543);
nand U6674 (N_6674,N_6483,N_6569);
nor U6675 (N_6675,N_6461,N_6570);
and U6676 (N_6676,N_6454,N_6567);
nor U6677 (N_6677,N_6524,N_6517);
or U6678 (N_6678,N_6468,N_6573);
xor U6679 (N_6679,N_6505,N_6489);
nand U6680 (N_6680,N_6536,N_6521);
nor U6681 (N_6681,N_6476,N_6457);
or U6682 (N_6682,N_6533,N_6546);
nand U6683 (N_6683,N_6526,N_6505);
and U6684 (N_6684,N_6522,N_6473);
nand U6685 (N_6685,N_6519,N_6499);
nor U6686 (N_6686,N_6596,N_6457);
nand U6687 (N_6687,N_6471,N_6505);
nor U6688 (N_6688,N_6538,N_6536);
nand U6689 (N_6689,N_6463,N_6585);
nor U6690 (N_6690,N_6466,N_6576);
xor U6691 (N_6691,N_6538,N_6458);
nor U6692 (N_6692,N_6509,N_6536);
nand U6693 (N_6693,N_6576,N_6487);
nand U6694 (N_6694,N_6500,N_6580);
nor U6695 (N_6695,N_6465,N_6460);
nor U6696 (N_6696,N_6455,N_6475);
and U6697 (N_6697,N_6546,N_6537);
nor U6698 (N_6698,N_6474,N_6584);
nand U6699 (N_6699,N_6593,N_6520);
nand U6700 (N_6700,N_6490,N_6541);
xnor U6701 (N_6701,N_6550,N_6489);
and U6702 (N_6702,N_6518,N_6557);
and U6703 (N_6703,N_6551,N_6472);
nand U6704 (N_6704,N_6452,N_6538);
nor U6705 (N_6705,N_6455,N_6592);
and U6706 (N_6706,N_6599,N_6541);
nor U6707 (N_6707,N_6474,N_6498);
nor U6708 (N_6708,N_6519,N_6595);
or U6709 (N_6709,N_6556,N_6489);
nor U6710 (N_6710,N_6567,N_6469);
nor U6711 (N_6711,N_6462,N_6555);
or U6712 (N_6712,N_6493,N_6564);
nor U6713 (N_6713,N_6572,N_6494);
xor U6714 (N_6714,N_6461,N_6568);
and U6715 (N_6715,N_6487,N_6466);
xnor U6716 (N_6716,N_6493,N_6509);
and U6717 (N_6717,N_6500,N_6508);
nand U6718 (N_6718,N_6466,N_6481);
or U6719 (N_6719,N_6532,N_6487);
xnor U6720 (N_6720,N_6582,N_6589);
or U6721 (N_6721,N_6543,N_6516);
and U6722 (N_6722,N_6552,N_6576);
xnor U6723 (N_6723,N_6531,N_6551);
nor U6724 (N_6724,N_6552,N_6475);
xor U6725 (N_6725,N_6494,N_6450);
nand U6726 (N_6726,N_6470,N_6585);
xnor U6727 (N_6727,N_6585,N_6525);
xnor U6728 (N_6728,N_6496,N_6568);
xnor U6729 (N_6729,N_6592,N_6530);
or U6730 (N_6730,N_6490,N_6450);
or U6731 (N_6731,N_6541,N_6501);
nor U6732 (N_6732,N_6583,N_6451);
nor U6733 (N_6733,N_6596,N_6533);
xnor U6734 (N_6734,N_6495,N_6522);
nand U6735 (N_6735,N_6563,N_6488);
nor U6736 (N_6736,N_6540,N_6491);
xnor U6737 (N_6737,N_6459,N_6526);
xor U6738 (N_6738,N_6511,N_6550);
nor U6739 (N_6739,N_6507,N_6525);
nor U6740 (N_6740,N_6462,N_6541);
xor U6741 (N_6741,N_6484,N_6535);
or U6742 (N_6742,N_6464,N_6583);
xnor U6743 (N_6743,N_6518,N_6459);
xnor U6744 (N_6744,N_6517,N_6496);
xnor U6745 (N_6745,N_6537,N_6480);
and U6746 (N_6746,N_6565,N_6477);
or U6747 (N_6747,N_6529,N_6504);
nand U6748 (N_6748,N_6522,N_6450);
or U6749 (N_6749,N_6495,N_6497);
and U6750 (N_6750,N_6715,N_6748);
nor U6751 (N_6751,N_6627,N_6702);
nand U6752 (N_6752,N_6744,N_6692);
nor U6753 (N_6753,N_6687,N_6681);
xnor U6754 (N_6754,N_6619,N_6645);
xor U6755 (N_6755,N_6630,N_6727);
xor U6756 (N_6756,N_6609,N_6699);
and U6757 (N_6757,N_6734,N_6678);
nand U6758 (N_6758,N_6608,N_6672);
and U6759 (N_6759,N_6623,N_6683);
and U6760 (N_6760,N_6724,N_6631);
or U6761 (N_6761,N_6693,N_6709);
or U6762 (N_6762,N_6656,N_6676);
nor U6763 (N_6763,N_6725,N_6714);
or U6764 (N_6764,N_6737,N_6602);
xnor U6765 (N_6765,N_6689,N_6612);
nand U6766 (N_6766,N_6650,N_6695);
nand U6767 (N_6767,N_6604,N_6641);
xor U6768 (N_6768,N_6662,N_6703);
nor U6769 (N_6769,N_6654,N_6664);
and U6770 (N_6770,N_6673,N_6633);
and U6771 (N_6771,N_6732,N_6700);
nand U6772 (N_6772,N_6713,N_6652);
or U6773 (N_6773,N_6697,N_6620);
or U6774 (N_6774,N_6651,N_6730);
and U6775 (N_6775,N_6648,N_6688);
nor U6776 (N_6776,N_6605,N_6660);
nand U6777 (N_6777,N_6741,N_6611);
and U6778 (N_6778,N_6712,N_6669);
nor U6779 (N_6779,N_6615,N_6647);
or U6780 (N_6780,N_6726,N_6642);
nand U6781 (N_6781,N_6632,N_6667);
xnor U6782 (N_6782,N_6607,N_6716);
xnor U6783 (N_6783,N_6655,N_6638);
nand U6784 (N_6784,N_6629,N_6640);
xor U6785 (N_6785,N_6685,N_6749);
or U6786 (N_6786,N_6624,N_6665);
and U6787 (N_6787,N_6696,N_6636);
nand U6788 (N_6788,N_6740,N_6690);
or U6789 (N_6789,N_6677,N_6637);
or U6790 (N_6790,N_6738,N_6718);
and U6791 (N_6791,N_6661,N_6711);
and U6792 (N_6792,N_6601,N_6621);
nand U6793 (N_6793,N_6625,N_6649);
nor U6794 (N_6794,N_6698,N_6663);
nand U6795 (N_6795,N_6668,N_6657);
nand U6796 (N_6796,N_6721,N_6675);
nor U6797 (N_6797,N_6635,N_6701);
xor U6798 (N_6798,N_6682,N_6729);
xnor U6799 (N_6799,N_6706,N_6742);
xnor U6800 (N_6800,N_6707,N_6735);
xor U6801 (N_6801,N_6659,N_6614);
xor U6802 (N_6802,N_6723,N_6720);
nor U6803 (N_6803,N_6731,N_6626);
xor U6804 (N_6804,N_6622,N_6686);
or U6805 (N_6805,N_6617,N_6613);
xor U6806 (N_6806,N_6603,N_6680);
xor U6807 (N_6807,N_6653,N_6710);
nor U6808 (N_6808,N_6610,N_6722);
nand U6809 (N_6809,N_6644,N_6606);
xor U6810 (N_6810,N_6628,N_6739);
nor U6811 (N_6811,N_6708,N_6719);
nor U6812 (N_6812,N_6705,N_6658);
nand U6813 (N_6813,N_6616,N_6745);
xor U6814 (N_6814,N_6639,N_6618);
and U6815 (N_6815,N_6717,N_6746);
nand U6816 (N_6816,N_6634,N_6666);
xnor U6817 (N_6817,N_6728,N_6670);
xnor U6818 (N_6818,N_6643,N_6646);
xor U6819 (N_6819,N_6671,N_6691);
and U6820 (N_6820,N_6600,N_6736);
and U6821 (N_6821,N_6733,N_6704);
xor U6822 (N_6822,N_6679,N_6694);
or U6823 (N_6823,N_6684,N_6747);
nor U6824 (N_6824,N_6743,N_6674);
nor U6825 (N_6825,N_6715,N_6697);
or U6826 (N_6826,N_6626,N_6677);
or U6827 (N_6827,N_6681,N_6664);
nand U6828 (N_6828,N_6680,N_6710);
xnor U6829 (N_6829,N_6625,N_6619);
nand U6830 (N_6830,N_6749,N_6726);
or U6831 (N_6831,N_6748,N_6625);
xnor U6832 (N_6832,N_6676,N_6641);
and U6833 (N_6833,N_6732,N_6632);
nand U6834 (N_6834,N_6641,N_6655);
nand U6835 (N_6835,N_6659,N_6737);
and U6836 (N_6836,N_6616,N_6719);
or U6837 (N_6837,N_6630,N_6657);
xnor U6838 (N_6838,N_6691,N_6661);
nor U6839 (N_6839,N_6691,N_6694);
nor U6840 (N_6840,N_6745,N_6659);
and U6841 (N_6841,N_6647,N_6721);
nor U6842 (N_6842,N_6675,N_6701);
and U6843 (N_6843,N_6696,N_6730);
xnor U6844 (N_6844,N_6698,N_6630);
nor U6845 (N_6845,N_6618,N_6744);
nand U6846 (N_6846,N_6744,N_6716);
or U6847 (N_6847,N_6600,N_6621);
and U6848 (N_6848,N_6634,N_6676);
or U6849 (N_6849,N_6629,N_6614);
nand U6850 (N_6850,N_6628,N_6697);
and U6851 (N_6851,N_6695,N_6744);
nand U6852 (N_6852,N_6653,N_6729);
nor U6853 (N_6853,N_6674,N_6666);
nand U6854 (N_6854,N_6694,N_6639);
and U6855 (N_6855,N_6647,N_6636);
or U6856 (N_6856,N_6641,N_6675);
and U6857 (N_6857,N_6624,N_6687);
nand U6858 (N_6858,N_6746,N_6744);
xnor U6859 (N_6859,N_6690,N_6632);
xor U6860 (N_6860,N_6736,N_6662);
or U6861 (N_6861,N_6705,N_6689);
nor U6862 (N_6862,N_6706,N_6680);
nor U6863 (N_6863,N_6605,N_6696);
or U6864 (N_6864,N_6742,N_6635);
xor U6865 (N_6865,N_6694,N_6738);
or U6866 (N_6866,N_6639,N_6678);
and U6867 (N_6867,N_6677,N_6604);
nor U6868 (N_6868,N_6700,N_6600);
nand U6869 (N_6869,N_6616,N_6618);
nor U6870 (N_6870,N_6696,N_6723);
or U6871 (N_6871,N_6725,N_6642);
nor U6872 (N_6872,N_6745,N_6671);
or U6873 (N_6873,N_6720,N_6739);
nor U6874 (N_6874,N_6748,N_6617);
nand U6875 (N_6875,N_6628,N_6705);
xnor U6876 (N_6876,N_6613,N_6640);
and U6877 (N_6877,N_6687,N_6647);
and U6878 (N_6878,N_6672,N_6724);
or U6879 (N_6879,N_6732,N_6631);
xor U6880 (N_6880,N_6729,N_6602);
nor U6881 (N_6881,N_6640,N_6678);
and U6882 (N_6882,N_6687,N_6707);
and U6883 (N_6883,N_6690,N_6614);
or U6884 (N_6884,N_6696,N_6667);
or U6885 (N_6885,N_6660,N_6650);
or U6886 (N_6886,N_6644,N_6600);
nand U6887 (N_6887,N_6617,N_6677);
xor U6888 (N_6888,N_6671,N_6620);
or U6889 (N_6889,N_6745,N_6733);
or U6890 (N_6890,N_6644,N_6617);
or U6891 (N_6891,N_6707,N_6685);
or U6892 (N_6892,N_6647,N_6736);
nand U6893 (N_6893,N_6730,N_6719);
or U6894 (N_6894,N_6716,N_6734);
or U6895 (N_6895,N_6617,N_6621);
and U6896 (N_6896,N_6674,N_6604);
or U6897 (N_6897,N_6675,N_6728);
or U6898 (N_6898,N_6616,N_6675);
or U6899 (N_6899,N_6627,N_6616);
xor U6900 (N_6900,N_6835,N_6853);
and U6901 (N_6901,N_6824,N_6809);
or U6902 (N_6902,N_6793,N_6764);
xnor U6903 (N_6903,N_6870,N_6899);
xnor U6904 (N_6904,N_6849,N_6894);
or U6905 (N_6905,N_6805,N_6872);
nor U6906 (N_6906,N_6772,N_6862);
nand U6907 (N_6907,N_6780,N_6858);
xor U6908 (N_6908,N_6799,N_6761);
and U6909 (N_6909,N_6814,N_6781);
or U6910 (N_6910,N_6827,N_6783);
or U6911 (N_6911,N_6753,N_6869);
nand U6912 (N_6912,N_6852,N_6757);
or U6913 (N_6913,N_6841,N_6790);
xor U6914 (N_6914,N_6765,N_6759);
nor U6915 (N_6915,N_6777,N_6826);
or U6916 (N_6916,N_6769,N_6878);
nand U6917 (N_6917,N_6791,N_6758);
xor U6918 (N_6918,N_6874,N_6861);
nand U6919 (N_6919,N_6831,N_6773);
and U6920 (N_6920,N_6786,N_6778);
or U6921 (N_6921,N_6821,N_6887);
or U6922 (N_6922,N_6860,N_6843);
or U6923 (N_6923,N_6875,N_6756);
nor U6924 (N_6924,N_6819,N_6762);
and U6925 (N_6925,N_6807,N_6890);
xor U6926 (N_6926,N_6796,N_6760);
and U6927 (N_6927,N_6752,N_6825);
nor U6928 (N_6928,N_6886,N_6897);
nor U6929 (N_6929,N_6863,N_6846);
and U6930 (N_6930,N_6816,N_6794);
nand U6931 (N_6931,N_6820,N_6880);
nor U6932 (N_6932,N_6750,N_6812);
and U6933 (N_6933,N_6848,N_6833);
nor U6934 (N_6934,N_6850,N_6779);
nor U6935 (N_6935,N_6792,N_6832);
xor U6936 (N_6936,N_6871,N_6766);
and U6937 (N_6937,N_6775,N_6891);
xnor U6938 (N_6938,N_6828,N_6802);
nand U6939 (N_6939,N_6804,N_6840);
nand U6940 (N_6940,N_6774,N_6842);
nand U6941 (N_6941,N_6844,N_6788);
xor U6942 (N_6942,N_6813,N_6839);
nand U6943 (N_6943,N_6798,N_6892);
and U6944 (N_6944,N_6789,N_6856);
nand U6945 (N_6945,N_6845,N_6855);
nand U6946 (N_6946,N_6782,N_6876);
nor U6947 (N_6947,N_6768,N_6895);
and U6948 (N_6948,N_6776,N_6823);
xnor U6949 (N_6949,N_6800,N_6836);
nor U6950 (N_6950,N_6865,N_6884);
nor U6951 (N_6951,N_6817,N_6881);
nor U6952 (N_6952,N_6857,N_6851);
nor U6953 (N_6953,N_6818,N_6806);
and U6954 (N_6954,N_6785,N_6801);
nor U6955 (N_6955,N_6803,N_6885);
nor U6956 (N_6956,N_6754,N_6898);
or U6957 (N_6957,N_6888,N_6859);
nand U6958 (N_6958,N_6784,N_6854);
nor U6959 (N_6959,N_6867,N_6883);
and U6960 (N_6960,N_6763,N_6893);
and U6961 (N_6961,N_6873,N_6837);
and U6962 (N_6962,N_6830,N_6815);
nand U6963 (N_6963,N_6868,N_6866);
or U6964 (N_6964,N_6877,N_6864);
nand U6965 (N_6965,N_6834,N_6847);
and U6966 (N_6966,N_6822,N_6882);
and U6967 (N_6967,N_6811,N_6838);
or U6968 (N_6968,N_6770,N_6767);
or U6969 (N_6969,N_6879,N_6771);
or U6970 (N_6970,N_6787,N_6797);
xor U6971 (N_6971,N_6889,N_6751);
nor U6972 (N_6972,N_6755,N_6829);
or U6973 (N_6973,N_6795,N_6810);
and U6974 (N_6974,N_6896,N_6808);
nand U6975 (N_6975,N_6803,N_6880);
or U6976 (N_6976,N_6755,N_6847);
or U6977 (N_6977,N_6774,N_6844);
or U6978 (N_6978,N_6894,N_6769);
or U6979 (N_6979,N_6867,N_6865);
nand U6980 (N_6980,N_6771,N_6872);
xor U6981 (N_6981,N_6830,N_6783);
nor U6982 (N_6982,N_6800,N_6849);
or U6983 (N_6983,N_6871,N_6807);
xnor U6984 (N_6984,N_6894,N_6853);
and U6985 (N_6985,N_6781,N_6867);
or U6986 (N_6986,N_6887,N_6761);
or U6987 (N_6987,N_6865,N_6870);
xor U6988 (N_6988,N_6780,N_6784);
nand U6989 (N_6989,N_6899,N_6767);
nor U6990 (N_6990,N_6779,N_6831);
nand U6991 (N_6991,N_6795,N_6754);
xnor U6992 (N_6992,N_6887,N_6881);
or U6993 (N_6993,N_6867,N_6862);
nand U6994 (N_6994,N_6848,N_6896);
nand U6995 (N_6995,N_6801,N_6869);
nand U6996 (N_6996,N_6899,N_6865);
xor U6997 (N_6997,N_6857,N_6892);
or U6998 (N_6998,N_6821,N_6853);
or U6999 (N_6999,N_6790,N_6828);
and U7000 (N_7000,N_6826,N_6776);
nand U7001 (N_7001,N_6862,N_6840);
nor U7002 (N_7002,N_6854,N_6786);
nand U7003 (N_7003,N_6876,N_6824);
nor U7004 (N_7004,N_6757,N_6853);
and U7005 (N_7005,N_6870,N_6764);
nor U7006 (N_7006,N_6855,N_6889);
or U7007 (N_7007,N_6790,N_6782);
nor U7008 (N_7008,N_6820,N_6847);
or U7009 (N_7009,N_6897,N_6827);
nor U7010 (N_7010,N_6788,N_6848);
xnor U7011 (N_7011,N_6859,N_6777);
and U7012 (N_7012,N_6885,N_6899);
nand U7013 (N_7013,N_6816,N_6897);
and U7014 (N_7014,N_6798,N_6890);
nor U7015 (N_7015,N_6815,N_6763);
and U7016 (N_7016,N_6777,N_6822);
xnor U7017 (N_7017,N_6847,N_6783);
or U7018 (N_7018,N_6833,N_6765);
and U7019 (N_7019,N_6870,N_6770);
and U7020 (N_7020,N_6822,N_6829);
nor U7021 (N_7021,N_6878,N_6810);
or U7022 (N_7022,N_6851,N_6780);
xor U7023 (N_7023,N_6889,N_6882);
or U7024 (N_7024,N_6843,N_6780);
nor U7025 (N_7025,N_6756,N_6893);
nand U7026 (N_7026,N_6750,N_6758);
xor U7027 (N_7027,N_6804,N_6838);
or U7028 (N_7028,N_6760,N_6751);
nand U7029 (N_7029,N_6846,N_6843);
or U7030 (N_7030,N_6782,N_6780);
and U7031 (N_7031,N_6884,N_6889);
nand U7032 (N_7032,N_6856,N_6834);
xnor U7033 (N_7033,N_6836,N_6887);
or U7034 (N_7034,N_6795,N_6751);
xnor U7035 (N_7035,N_6851,N_6841);
or U7036 (N_7036,N_6768,N_6798);
xor U7037 (N_7037,N_6870,N_6835);
xor U7038 (N_7038,N_6835,N_6809);
nand U7039 (N_7039,N_6839,N_6859);
or U7040 (N_7040,N_6862,N_6896);
nor U7041 (N_7041,N_6815,N_6827);
nand U7042 (N_7042,N_6852,N_6874);
and U7043 (N_7043,N_6839,N_6845);
xnor U7044 (N_7044,N_6831,N_6759);
xor U7045 (N_7045,N_6778,N_6755);
xor U7046 (N_7046,N_6793,N_6846);
or U7047 (N_7047,N_6820,N_6833);
xor U7048 (N_7048,N_6768,N_6786);
xor U7049 (N_7049,N_6754,N_6769);
or U7050 (N_7050,N_7019,N_6993);
and U7051 (N_7051,N_7024,N_7049);
nor U7052 (N_7052,N_6909,N_7037);
or U7053 (N_7053,N_6935,N_7026);
or U7054 (N_7054,N_6972,N_6960);
or U7055 (N_7055,N_6924,N_6903);
nand U7056 (N_7056,N_6961,N_6911);
xor U7057 (N_7057,N_6951,N_7018);
or U7058 (N_7058,N_6938,N_7040);
and U7059 (N_7059,N_6954,N_6940);
nor U7060 (N_7060,N_7012,N_6906);
nor U7061 (N_7061,N_6999,N_6988);
or U7062 (N_7062,N_6959,N_6900);
xnor U7063 (N_7063,N_6977,N_7036);
and U7064 (N_7064,N_6910,N_7004);
and U7065 (N_7065,N_7027,N_6933);
nor U7066 (N_7066,N_6952,N_7044);
or U7067 (N_7067,N_6986,N_6942);
and U7068 (N_7068,N_7020,N_6930);
or U7069 (N_7069,N_6958,N_7042);
xnor U7070 (N_7070,N_6949,N_6980);
xor U7071 (N_7071,N_7035,N_6996);
and U7072 (N_7072,N_6981,N_6922);
xnor U7073 (N_7073,N_7028,N_6907);
xor U7074 (N_7074,N_6946,N_6997);
or U7075 (N_7075,N_6927,N_6976);
or U7076 (N_7076,N_6947,N_6948);
nor U7077 (N_7077,N_7008,N_7022);
nor U7078 (N_7078,N_7016,N_6929);
and U7079 (N_7079,N_6912,N_6969);
nor U7080 (N_7080,N_6914,N_6932);
or U7081 (N_7081,N_6901,N_6973);
xor U7082 (N_7082,N_6978,N_6928);
nand U7083 (N_7083,N_6915,N_6943);
nor U7084 (N_7084,N_6925,N_6962);
and U7085 (N_7085,N_6991,N_7011);
xor U7086 (N_7086,N_6939,N_6945);
nand U7087 (N_7087,N_6964,N_7033);
and U7088 (N_7088,N_6992,N_6934);
xor U7089 (N_7089,N_7023,N_6944);
and U7090 (N_7090,N_7038,N_7046);
and U7091 (N_7091,N_7010,N_7025);
and U7092 (N_7092,N_6971,N_6918);
or U7093 (N_7093,N_6989,N_6974);
nor U7094 (N_7094,N_6975,N_6920);
nor U7095 (N_7095,N_6983,N_6904);
xnor U7096 (N_7096,N_6905,N_6956);
nand U7097 (N_7097,N_6937,N_6998);
nor U7098 (N_7098,N_6902,N_6979);
nand U7099 (N_7099,N_7047,N_6950);
xnor U7100 (N_7100,N_7030,N_6985);
nor U7101 (N_7101,N_6963,N_6968);
xnor U7102 (N_7102,N_6926,N_7003);
nand U7103 (N_7103,N_7013,N_6990);
nand U7104 (N_7104,N_6982,N_6967);
nor U7105 (N_7105,N_6955,N_7000);
and U7106 (N_7106,N_7006,N_7041);
nand U7107 (N_7107,N_7001,N_7009);
nand U7108 (N_7108,N_6994,N_6953);
xor U7109 (N_7109,N_7031,N_6965);
nor U7110 (N_7110,N_7015,N_7002);
xor U7111 (N_7111,N_6995,N_6970);
nor U7112 (N_7112,N_7021,N_6923);
or U7113 (N_7113,N_7007,N_7032);
and U7114 (N_7114,N_6984,N_6957);
nand U7115 (N_7115,N_6966,N_7029);
nor U7116 (N_7116,N_7034,N_7014);
and U7117 (N_7117,N_6916,N_6941);
nor U7118 (N_7118,N_7045,N_6913);
nand U7119 (N_7119,N_6921,N_7043);
nand U7120 (N_7120,N_6936,N_6917);
nor U7121 (N_7121,N_7005,N_6908);
nor U7122 (N_7122,N_6919,N_7048);
nor U7123 (N_7123,N_7039,N_7017);
nor U7124 (N_7124,N_6931,N_6987);
or U7125 (N_7125,N_7029,N_7048);
nand U7126 (N_7126,N_6909,N_6973);
xor U7127 (N_7127,N_7007,N_6902);
xor U7128 (N_7128,N_6953,N_6993);
or U7129 (N_7129,N_6922,N_6920);
or U7130 (N_7130,N_6932,N_7013);
or U7131 (N_7131,N_7021,N_7036);
nand U7132 (N_7132,N_6973,N_7033);
nor U7133 (N_7133,N_6999,N_7009);
nor U7134 (N_7134,N_6946,N_6917);
nand U7135 (N_7135,N_6953,N_6936);
xor U7136 (N_7136,N_6954,N_6937);
or U7137 (N_7137,N_7040,N_6902);
nor U7138 (N_7138,N_6989,N_6962);
and U7139 (N_7139,N_6985,N_6927);
nor U7140 (N_7140,N_6905,N_6973);
nor U7141 (N_7141,N_6921,N_7006);
xnor U7142 (N_7142,N_6964,N_6922);
nand U7143 (N_7143,N_6975,N_6985);
xor U7144 (N_7144,N_7001,N_6951);
nand U7145 (N_7145,N_6985,N_6979);
nor U7146 (N_7146,N_6964,N_7042);
nand U7147 (N_7147,N_7004,N_6930);
nor U7148 (N_7148,N_7017,N_6944);
or U7149 (N_7149,N_7023,N_7041);
or U7150 (N_7150,N_6946,N_6974);
nor U7151 (N_7151,N_7018,N_6971);
nor U7152 (N_7152,N_6951,N_7007);
nand U7153 (N_7153,N_6936,N_7034);
xnor U7154 (N_7154,N_7001,N_6910);
xnor U7155 (N_7155,N_6986,N_6971);
xnor U7156 (N_7156,N_6926,N_6950);
or U7157 (N_7157,N_7040,N_7021);
xor U7158 (N_7158,N_6958,N_6999);
nor U7159 (N_7159,N_7042,N_6945);
or U7160 (N_7160,N_6961,N_7018);
and U7161 (N_7161,N_7025,N_7030);
xnor U7162 (N_7162,N_6949,N_7007);
and U7163 (N_7163,N_6920,N_6912);
or U7164 (N_7164,N_6998,N_6941);
or U7165 (N_7165,N_7005,N_6956);
and U7166 (N_7166,N_7011,N_6906);
and U7167 (N_7167,N_7044,N_6934);
or U7168 (N_7168,N_6998,N_7024);
nand U7169 (N_7169,N_7000,N_6966);
nor U7170 (N_7170,N_7009,N_6943);
nor U7171 (N_7171,N_6992,N_6961);
xor U7172 (N_7172,N_6973,N_7013);
and U7173 (N_7173,N_7008,N_6981);
or U7174 (N_7174,N_6961,N_7023);
nand U7175 (N_7175,N_7040,N_7029);
and U7176 (N_7176,N_7014,N_6906);
xnor U7177 (N_7177,N_6919,N_7023);
nor U7178 (N_7178,N_6978,N_7003);
xor U7179 (N_7179,N_7049,N_7034);
nor U7180 (N_7180,N_6920,N_6919);
nand U7181 (N_7181,N_6941,N_6955);
and U7182 (N_7182,N_6929,N_6970);
xor U7183 (N_7183,N_6955,N_7027);
and U7184 (N_7184,N_6981,N_7007);
and U7185 (N_7185,N_6950,N_6960);
and U7186 (N_7186,N_6986,N_6925);
and U7187 (N_7187,N_6927,N_7013);
and U7188 (N_7188,N_7043,N_6944);
and U7189 (N_7189,N_7008,N_7039);
nand U7190 (N_7190,N_6905,N_6948);
xnor U7191 (N_7191,N_6978,N_7030);
and U7192 (N_7192,N_6921,N_7045);
nand U7193 (N_7193,N_7037,N_7043);
and U7194 (N_7194,N_7018,N_6922);
and U7195 (N_7195,N_6995,N_6972);
and U7196 (N_7196,N_7048,N_6954);
nand U7197 (N_7197,N_7043,N_7017);
and U7198 (N_7198,N_7043,N_6985);
nand U7199 (N_7199,N_7016,N_7044);
and U7200 (N_7200,N_7138,N_7086);
nand U7201 (N_7201,N_7123,N_7193);
nand U7202 (N_7202,N_7087,N_7192);
or U7203 (N_7203,N_7052,N_7136);
xor U7204 (N_7204,N_7148,N_7073);
nor U7205 (N_7205,N_7083,N_7116);
nand U7206 (N_7206,N_7174,N_7150);
and U7207 (N_7207,N_7161,N_7183);
and U7208 (N_7208,N_7177,N_7072);
xnor U7209 (N_7209,N_7055,N_7074);
nand U7210 (N_7210,N_7173,N_7190);
and U7211 (N_7211,N_7164,N_7078);
nand U7212 (N_7212,N_7105,N_7062);
nor U7213 (N_7213,N_7071,N_7121);
xnor U7214 (N_7214,N_7088,N_7084);
or U7215 (N_7215,N_7166,N_7097);
or U7216 (N_7216,N_7163,N_7104);
and U7217 (N_7217,N_7149,N_7154);
nand U7218 (N_7218,N_7167,N_7111);
or U7219 (N_7219,N_7195,N_7180);
or U7220 (N_7220,N_7054,N_7144);
xnor U7221 (N_7221,N_7134,N_7142);
or U7222 (N_7222,N_7137,N_7120);
and U7223 (N_7223,N_7053,N_7162);
xor U7224 (N_7224,N_7060,N_7135);
nor U7225 (N_7225,N_7091,N_7095);
and U7226 (N_7226,N_7090,N_7125);
and U7227 (N_7227,N_7160,N_7124);
or U7228 (N_7228,N_7102,N_7185);
nor U7229 (N_7229,N_7169,N_7197);
nand U7230 (N_7230,N_7065,N_7186);
nor U7231 (N_7231,N_7194,N_7069);
nor U7232 (N_7232,N_7122,N_7198);
xor U7233 (N_7233,N_7098,N_7159);
xnor U7234 (N_7234,N_7093,N_7127);
and U7235 (N_7235,N_7176,N_7101);
or U7236 (N_7236,N_7118,N_7109);
nor U7237 (N_7237,N_7155,N_7181);
and U7238 (N_7238,N_7141,N_7115);
or U7239 (N_7239,N_7106,N_7158);
nor U7240 (N_7240,N_7066,N_7050);
and U7241 (N_7241,N_7187,N_7057);
nand U7242 (N_7242,N_7094,N_7099);
or U7243 (N_7243,N_7171,N_7179);
nand U7244 (N_7244,N_7059,N_7153);
or U7245 (N_7245,N_7061,N_7114);
nand U7246 (N_7246,N_7140,N_7165);
nand U7247 (N_7247,N_7082,N_7191);
nor U7248 (N_7248,N_7096,N_7196);
and U7249 (N_7249,N_7058,N_7092);
nor U7250 (N_7250,N_7172,N_7152);
xor U7251 (N_7251,N_7103,N_7128);
nand U7252 (N_7252,N_7064,N_7188);
or U7253 (N_7253,N_7199,N_7067);
nand U7254 (N_7254,N_7139,N_7151);
nand U7255 (N_7255,N_7079,N_7108);
xnor U7256 (N_7256,N_7070,N_7189);
xnor U7257 (N_7257,N_7132,N_7170);
or U7258 (N_7258,N_7130,N_7089);
and U7259 (N_7259,N_7112,N_7056);
and U7260 (N_7260,N_7131,N_7145);
nor U7261 (N_7261,N_7126,N_7175);
xnor U7262 (N_7262,N_7156,N_7051);
or U7263 (N_7263,N_7068,N_7075);
nor U7264 (N_7264,N_7107,N_7182);
nand U7265 (N_7265,N_7146,N_7119);
or U7266 (N_7266,N_7085,N_7143);
or U7267 (N_7267,N_7133,N_7077);
and U7268 (N_7268,N_7168,N_7076);
nand U7269 (N_7269,N_7184,N_7063);
nand U7270 (N_7270,N_7081,N_7147);
or U7271 (N_7271,N_7100,N_7113);
nand U7272 (N_7272,N_7117,N_7110);
and U7273 (N_7273,N_7178,N_7080);
or U7274 (N_7274,N_7157,N_7129);
xnor U7275 (N_7275,N_7104,N_7073);
xnor U7276 (N_7276,N_7179,N_7184);
xnor U7277 (N_7277,N_7154,N_7160);
or U7278 (N_7278,N_7174,N_7179);
or U7279 (N_7279,N_7124,N_7119);
nor U7280 (N_7280,N_7121,N_7082);
or U7281 (N_7281,N_7138,N_7069);
xor U7282 (N_7282,N_7183,N_7050);
xor U7283 (N_7283,N_7139,N_7085);
xnor U7284 (N_7284,N_7185,N_7053);
or U7285 (N_7285,N_7198,N_7174);
nor U7286 (N_7286,N_7152,N_7052);
nand U7287 (N_7287,N_7077,N_7074);
nor U7288 (N_7288,N_7169,N_7104);
or U7289 (N_7289,N_7097,N_7085);
xor U7290 (N_7290,N_7082,N_7193);
xnor U7291 (N_7291,N_7154,N_7054);
nand U7292 (N_7292,N_7106,N_7122);
and U7293 (N_7293,N_7177,N_7137);
xor U7294 (N_7294,N_7141,N_7059);
and U7295 (N_7295,N_7120,N_7189);
xnor U7296 (N_7296,N_7148,N_7070);
or U7297 (N_7297,N_7175,N_7180);
xnor U7298 (N_7298,N_7089,N_7136);
xnor U7299 (N_7299,N_7091,N_7138);
xor U7300 (N_7300,N_7159,N_7169);
or U7301 (N_7301,N_7190,N_7118);
xor U7302 (N_7302,N_7099,N_7098);
nor U7303 (N_7303,N_7104,N_7061);
nand U7304 (N_7304,N_7127,N_7159);
nand U7305 (N_7305,N_7135,N_7181);
or U7306 (N_7306,N_7169,N_7119);
xnor U7307 (N_7307,N_7177,N_7188);
nor U7308 (N_7308,N_7130,N_7096);
nor U7309 (N_7309,N_7066,N_7142);
nand U7310 (N_7310,N_7096,N_7152);
nand U7311 (N_7311,N_7112,N_7119);
and U7312 (N_7312,N_7079,N_7183);
or U7313 (N_7313,N_7111,N_7157);
nand U7314 (N_7314,N_7101,N_7104);
xor U7315 (N_7315,N_7163,N_7057);
or U7316 (N_7316,N_7145,N_7132);
or U7317 (N_7317,N_7184,N_7135);
or U7318 (N_7318,N_7184,N_7140);
and U7319 (N_7319,N_7113,N_7125);
and U7320 (N_7320,N_7086,N_7104);
and U7321 (N_7321,N_7148,N_7173);
or U7322 (N_7322,N_7082,N_7088);
xnor U7323 (N_7323,N_7061,N_7190);
nor U7324 (N_7324,N_7061,N_7157);
nor U7325 (N_7325,N_7098,N_7161);
nor U7326 (N_7326,N_7071,N_7141);
nand U7327 (N_7327,N_7160,N_7059);
nand U7328 (N_7328,N_7098,N_7065);
xor U7329 (N_7329,N_7169,N_7175);
or U7330 (N_7330,N_7187,N_7151);
xnor U7331 (N_7331,N_7112,N_7148);
nor U7332 (N_7332,N_7073,N_7164);
xnor U7333 (N_7333,N_7158,N_7159);
xor U7334 (N_7334,N_7195,N_7111);
or U7335 (N_7335,N_7094,N_7156);
or U7336 (N_7336,N_7112,N_7118);
or U7337 (N_7337,N_7152,N_7105);
xnor U7338 (N_7338,N_7148,N_7136);
xor U7339 (N_7339,N_7066,N_7054);
nor U7340 (N_7340,N_7130,N_7135);
and U7341 (N_7341,N_7171,N_7140);
nand U7342 (N_7342,N_7195,N_7143);
xor U7343 (N_7343,N_7142,N_7125);
nor U7344 (N_7344,N_7083,N_7086);
or U7345 (N_7345,N_7088,N_7159);
xor U7346 (N_7346,N_7192,N_7066);
or U7347 (N_7347,N_7051,N_7191);
nor U7348 (N_7348,N_7126,N_7079);
xor U7349 (N_7349,N_7109,N_7066);
xnor U7350 (N_7350,N_7282,N_7219);
or U7351 (N_7351,N_7218,N_7246);
or U7352 (N_7352,N_7332,N_7271);
and U7353 (N_7353,N_7288,N_7345);
nor U7354 (N_7354,N_7295,N_7245);
and U7355 (N_7355,N_7243,N_7254);
and U7356 (N_7356,N_7286,N_7220);
or U7357 (N_7357,N_7341,N_7340);
and U7358 (N_7358,N_7294,N_7285);
and U7359 (N_7359,N_7274,N_7251);
xnor U7360 (N_7360,N_7256,N_7269);
xor U7361 (N_7361,N_7238,N_7277);
or U7362 (N_7362,N_7334,N_7207);
and U7363 (N_7363,N_7335,N_7339);
xnor U7364 (N_7364,N_7203,N_7284);
or U7365 (N_7365,N_7297,N_7264);
or U7366 (N_7366,N_7221,N_7280);
nor U7367 (N_7367,N_7316,N_7349);
and U7368 (N_7368,N_7231,N_7273);
nor U7369 (N_7369,N_7348,N_7292);
xor U7370 (N_7370,N_7242,N_7208);
or U7371 (N_7371,N_7310,N_7291);
nor U7372 (N_7372,N_7342,N_7287);
xor U7373 (N_7373,N_7213,N_7346);
nand U7374 (N_7374,N_7236,N_7293);
nand U7375 (N_7375,N_7257,N_7263);
nand U7376 (N_7376,N_7312,N_7338);
and U7377 (N_7377,N_7301,N_7202);
and U7378 (N_7378,N_7214,N_7237);
and U7379 (N_7379,N_7252,N_7211);
and U7380 (N_7380,N_7240,N_7321);
xor U7381 (N_7381,N_7331,N_7255);
xnor U7382 (N_7382,N_7215,N_7333);
and U7383 (N_7383,N_7268,N_7308);
and U7384 (N_7384,N_7206,N_7217);
nand U7385 (N_7385,N_7307,N_7212);
nand U7386 (N_7386,N_7311,N_7227);
xnor U7387 (N_7387,N_7262,N_7224);
xnor U7388 (N_7388,N_7247,N_7244);
or U7389 (N_7389,N_7261,N_7283);
or U7390 (N_7390,N_7209,N_7258);
and U7391 (N_7391,N_7309,N_7314);
nor U7392 (N_7392,N_7327,N_7343);
xnor U7393 (N_7393,N_7302,N_7303);
and U7394 (N_7394,N_7241,N_7253);
nand U7395 (N_7395,N_7260,N_7229);
and U7396 (N_7396,N_7330,N_7317);
or U7397 (N_7397,N_7222,N_7228);
nor U7398 (N_7398,N_7235,N_7248);
nor U7399 (N_7399,N_7319,N_7289);
xor U7400 (N_7400,N_7200,N_7249);
and U7401 (N_7401,N_7210,N_7234);
or U7402 (N_7402,N_7344,N_7204);
nand U7403 (N_7403,N_7230,N_7322);
nand U7404 (N_7404,N_7313,N_7300);
and U7405 (N_7405,N_7337,N_7223);
or U7406 (N_7406,N_7225,N_7336);
nor U7407 (N_7407,N_7320,N_7278);
and U7408 (N_7408,N_7265,N_7279);
and U7409 (N_7409,N_7275,N_7329);
xnor U7410 (N_7410,N_7323,N_7304);
xor U7411 (N_7411,N_7328,N_7290);
and U7412 (N_7412,N_7315,N_7299);
nor U7413 (N_7413,N_7232,N_7306);
xnor U7414 (N_7414,N_7226,N_7325);
nor U7415 (N_7415,N_7266,N_7250);
or U7416 (N_7416,N_7326,N_7281);
nor U7417 (N_7417,N_7272,N_7318);
nor U7418 (N_7418,N_7259,N_7296);
or U7419 (N_7419,N_7347,N_7270);
or U7420 (N_7420,N_7267,N_7233);
xor U7421 (N_7421,N_7276,N_7298);
or U7422 (N_7422,N_7239,N_7201);
and U7423 (N_7423,N_7205,N_7324);
or U7424 (N_7424,N_7216,N_7305);
or U7425 (N_7425,N_7254,N_7320);
xnor U7426 (N_7426,N_7267,N_7339);
nor U7427 (N_7427,N_7277,N_7227);
or U7428 (N_7428,N_7228,N_7271);
xnor U7429 (N_7429,N_7203,N_7237);
nand U7430 (N_7430,N_7225,N_7328);
nand U7431 (N_7431,N_7282,N_7344);
nor U7432 (N_7432,N_7280,N_7237);
xor U7433 (N_7433,N_7337,N_7233);
or U7434 (N_7434,N_7250,N_7290);
xnor U7435 (N_7435,N_7275,N_7224);
or U7436 (N_7436,N_7339,N_7271);
or U7437 (N_7437,N_7289,N_7275);
or U7438 (N_7438,N_7321,N_7221);
xnor U7439 (N_7439,N_7243,N_7230);
nor U7440 (N_7440,N_7203,N_7322);
or U7441 (N_7441,N_7306,N_7246);
nor U7442 (N_7442,N_7239,N_7237);
nand U7443 (N_7443,N_7269,N_7253);
xnor U7444 (N_7444,N_7305,N_7315);
nor U7445 (N_7445,N_7266,N_7218);
nor U7446 (N_7446,N_7274,N_7207);
nand U7447 (N_7447,N_7314,N_7226);
and U7448 (N_7448,N_7323,N_7306);
xor U7449 (N_7449,N_7215,N_7292);
or U7450 (N_7450,N_7281,N_7312);
or U7451 (N_7451,N_7344,N_7251);
or U7452 (N_7452,N_7239,N_7224);
and U7453 (N_7453,N_7348,N_7257);
or U7454 (N_7454,N_7339,N_7222);
or U7455 (N_7455,N_7252,N_7284);
nand U7456 (N_7456,N_7341,N_7271);
xor U7457 (N_7457,N_7221,N_7324);
and U7458 (N_7458,N_7309,N_7236);
nand U7459 (N_7459,N_7270,N_7278);
xnor U7460 (N_7460,N_7340,N_7307);
nand U7461 (N_7461,N_7270,N_7219);
or U7462 (N_7462,N_7201,N_7267);
nor U7463 (N_7463,N_7244,N_7227);
and U7464 (N_7464,N_7347,N_7213);
and U7465 (N_7465,N_7342,N_7271);
nand U7466 (N_7466,N_7291,N_7257);
nor U7467 (N_7467,N_7310,N_7253);
xor U7468 (N_7468,N_7300,N_7316);
nand U7469 (N_7469,N_7233,N_7348);
and U7470 (N_7470,N_7238,N_7283);
nor U7471 (N_7471,N_7343,N_7207);
nand U7472 (N_7472,N_7312,N_7239);
nor U7473 (N_7473,N_7226,N_7296);
nand U7474 (N_7474,N_7265,N_7281);
or U7475 (N_7475,N_7298,N_7299);
and U7476 (N_7476,N_7294,N_7345);
and U7477 (N_7477,N_7255,N_7320);
or U7478 (N_7478,N_7327,N_7239);
or U7479 (N_7479,N_7284,N_7317);
xnor U7480 (N_7480,N_7206,N_7220);
or U7481 (N_7481,N_7277,N_7303);
or U7482 (N_7482,N_7286,N_7276);
nor U7483 (N_7483,N_7202,N_7326);
xnor U7484 (N_7484,N_7250,N_7273);
nand U7485 (N_7485,N_7258,N_7260);
and U7486 (N_7486,N_7319,N_7310);
nand U7487 (N_7487,N_7341,N_7327);
or U7488 (N_7488,N_7330,N_7346);
nor U7489 (N_7489,N_7271,N_7235);
nand U7490 (N_7490,N_7323,N_7331);
nand U7491 (N_7491,N_7228,N_7297);
and U7492 (N_7492,N_7333,N_7285);
nand U7493 (N_7493,N_7254,N_7281);
xor U7494 (N_7494,N_7307,N_7261);
and U7495 (N_7495,N_7277,N_7209);
or U7496 (N_7496,N_7260,N_7261);
nor U7497 (N_7497,N_7234,N_7202);
nand U7498 (N_7498,N_7338,N_7267);
and U7499 (N_7499,N_7332,N_7346);
or U7500 (N_7500,N_7441,N_7388);
nor U7501 (N_7501,N_7412,N_7486);
or U7502 (N_7502,N_7399,N_7352);
or U7503 (N_7503,N_7360,N_7458);
nand U7504 (N_7504,N_7408,N_7484);
and U7505 (N_7505,N_7442,N_7480);
and U7506 (N_7506,N_7462,N_7454);
nand U7507 (N_7507,N_7404,N_7495);
nand U7508 (N_7508,N_7471,N_7449);
xnor U7509 (N_7509,N_7405,N_7386);
or U7510 (N_7510,N_7440,N_7420);
xnor U7511 (N_7511,N_7393,N_7467);
xor U7512 (N_7512,N_7409,N_7483);
nor U7513 (N_7513,N_7478,N_7384);
xor U7514 (N_7514,N_7437,N_7391);
and U7515 (N_7515,N_7356,N_7417);
and U7516 (N_7516,N_7455,N_7353);
and U7517 (N_7517,N_7448,N_7445);
xnor U7518 (N_7518,N_7398,N_7379);
and U7519 (N_7519,N_7460,N_7406);
and U7520 (N_7520,N_7362,N_7482);
xnor U7521 (N_7521,N_7392,N_7457);
xor U7522 (N_7522,N_7450,N_7375);
or U7523 (N_7523,N_7401,N_7473);
and U7524 (N_7524,N_7470,N_7456);
xnor U7525 (N_7525,N_7354,N_7387);
and U7526 (N_7526,N_7489,N_7461);
xnor U7527 (N_7527,N_7477,N_7383);
or U7528 (N_7528,N_7370,N_7453);
xnor U7529 (N_7529,N_7373,N_7479);
and U7530 (N_7530,N_7490,N_7430);
or U7531 (N_7531,N_7422,N_7364);
or U7532 (N_7532,N_7425,N_7378);
or U7533 (N_7533,N_7390,N_7363);
xor U7534 (N_7534,N_7367,N_7451);
xnor U7535 (N_7535,N_7444,N_7400);
nand U7536 (N_7536,N_7418,N_7494);
or U7537 (N_7537,N_7468,N_7429);
or U7538 (N_7538,N_7443,N_7433);
xnor U7539 (N_7539,N_7371,N_7491);
nand U7540 (N_7540,N_7350,N_7428);
xor U7541 (N_7541,N_7472,N_7481);
nand U7542 (N_7542,N_7426,N_7488);
nor U7543 (N_7543,N_7366,N_7396);
or U7544 (N_7544,N_7474,N_7434);
xnor U7545 (N_7545,N_7464,N_7436);
and U7546 (N_7546,N_7485,N_7499);
and U7547 (N_7547,N_7452,N_7372);
nor U7548 (N_7548,N_7382,N_7402);
nand U7549 (N_7549,N_7427,N_7377);
or U7550 (N_7550,N_7497,N_7432);
or U7551 (N_7551,N_7431,N_7438);
nor U7552 (N_7552,N_7469,N_7487);
xnor U7553 (N_7553,N_7359,N_7380);
or U7554 (N_7554,N_7435,N_7413);
nor U7555 (N_7555,N_7389,N_7496);
and U7556 (N_7556,N_7424,N_7421);
nor U7557 (N_7557,N_7355,N_7475);
or U7558 (N_7558,N_7439,N_7492);
nand U7559 (N_7559,N_7414,N_7403);
xor U7560 (N_7560,N_7410,N_7374);
and U7561 (N_7561,N_7381,N_7385);
nor U7562 (N_7562,N_7369,N_7416);
nand U7563 (N_7563,N_7395,N_7498);
nand U7564 (N_7564,N_7407,N_7476);
or U7565 (N_7565,N_7357,N_7465);
and U7566 (N_7566,N_7411,N_7423);
and U7567 (N_7567,N_7419,N_7376);
nor U7568 (N_7568,N_7361,N_7447);
or U7569 (N_7569,N_7351,N_7493);
nor U7570 (N_7570,N_7415,N_7368);
or U7571 (N_7571,N_7446,N_7358);
nor U7572 (N_7572,N_7459,N_7466);
xnor U7573 (N_7573,N_7397,N_7463);
nor U7574 (N_7574,N_7365,N_7394);
xor U7575 (N_7575,N_7363,N_7374);
nor U7576 (N_7576,N_7489,N_7399);
xor U7577 (N_7577,N_7436,N_7468);
nor U7578 (N_7578,N_7401,N_7440);
nor U7579 (N_7579,N_7367,N_7355);
and U7580 (N_7580,N_7454,N_7369);
nand U7581 (N_7581,N_7494,N_7393);
or U7582 (N_7582,N_7482,N_7377);
nand U7583 (N_7583,N_7392,N_7486);
xnor U7584 (N_7584,N_7484,N_7406);
nor U7585 (N_7585,N_7417,N_7418);
nor U7586 (N_7586,N_7399,N_7357);
nand U7587 (N_7587,N_7424,N_7429);
and U7588 (N_7588,N_7421,N_7380);
nor U7589 (N_7589,N_7488,N_7423);
xnor U7590 (N_7590,N_7412,N_7401);
nor U7591 (N_7591,N_7452,N_7434);
nor U7592 (N_7592,N_7407,N_7494);
xnor U7593 (N_7593,N_7446,N_7373);
nor U7594 (N_7594,N_7492,N_7386);
nor U7595 (N_7595,N_7413,N_7373);
and U7596 (N_7596,N_7359,N_7452);
nor U7597 (N_7597,N_7358,N_7468);
or U7598 (N_7598,N_7477,N_7494);
and U7599 (N_7599,N_7406,N_7473);
xor U7600 (N_7600,N_7490,N_7382);
and U7601 (N_7601,N_7395,N_7400);
xnor U7602 (N_7602,N_7396,N_7397);
nand U7603 (N_7603,N_7473,N_7381);
and U7604 (N_7604,N_7394,N_7453);
nand U7605 (N_7605,N_7491,N_7430);
nor U7606 (N_7606,N_7369,N_7451);
and U7607 (N_7607,N_7414,N_7457);
or U7608 (N_7608,N_7359,N_7354);
nand U7609 (N_7609,N_7367,N_7363);
or U7610 (N_7610,N_7404,N_7465);
xor U7611 (N_7611,N_7473,N_7361);
and U7612 (N_7612,N_7376,N_7407);
nor U7613 (N_7613,N_7408,N_7390);
or U7614 (N_7614,N_7488,N_7439);
xnor U7615 (N_7615,N_7482,N_7471);
xor U7616 (N_7616,N_7461,N_7452);
nand U7617 (N_7617,N_7491,N_7437);
nor U7618 (N_7618,N_7395,N_7350);
nor U7619 (N_7619,N_7377,N_7450);
xor U7620 (N_7620,N_7419,N_7372);
or U7621 (N_7621,N_7455,N_7381);
nand U7622 (N_7622,N_7411,N_7373);
nand U7623 (N_7623,N_7371,N_7424);
nand U7624 (N_7624,N_7440,N_7426);
or U7625 (N_7625,N_7417,N_7384);
xor U7626 (N_7626,N_7353,N_7424);
or U7627 (N_7627,N_7403,N_7491);
nor U7628 (N_7628,N_7405,N_7419);
and U7629 (N_7629,N_7398,N_7356);
and U7630 (N_7630,N_7401,N_7476);
and U7631 (N_7631,N_7479,N_7416);
xor U7632 (N_7632,N_7401,N_7381);
nand U7633 (N_7633,N_7480,N_7409);
and U7634 (N_7634,N_7399,N_7413);
xnor U7635 (N_7635,N_7425,N_7350);
nand U7636 (N_7636,N_7459,N_7428);
nor U7637 (N_7637,N_7475,N_7488);
nand U7638 (N_7638,N_7412,N_7456);
nand U7639 (N_7639,N_7365,N_7411);
nor U7640 (N_7640,N_7367,N_7467);
nor U7641 (N_7641,N_7370,N_7380);
xor U7642 (N_7642,N_7399,N_7499);
or U7643 (N_7643,N_7419,N_7395);
nor U7644 (N_7644,N_7386,N_7471);
nand U7645 (N_7645,N_7365,N_7389);
nor U7646 (N_7646,N_7385,N_7497);
xor U7647 (N_7647,N_7447,N_7360);
nand U7648 (N_7648,N_7400,N_7480);
or U7649 (N_7649,N_7371,N_7366);
and U7650 (N_7650,N_7620,N_7515);
nand U7651 (N_7651,N_7549,N_7565);
and U7652 (N_7652,N_7590,N_7519);
and U7653 (N_7653,N_7624,N_7625);
or U7654 (N_7654,N_7628,N_7636);
and U7655 (N_7655,N_7638,N_7570);
nor U7656 (N_7656,N_7523,N_7533);
xnor U7657 (N_7657,N_7611,N_7527);
nor U7658 (N_7658,N_7560,N_7524);
nand U7659 (N_7659,N_7574,N_7568);
xnor U7660 (N_7660,N_7631,N_7547);
xnor U7661 (N_7661,N_7613,N_7649);
or U7662 (N_7662,N_7556,N_7554);
nor U7663 (N_7663,N_7516,N_7579);
and U7664 (N_7664,N_7550,N_7542);
nand U7665 (N_7665,N_7511,N_7608);
or U7666 (N_7666,N_7587,N_7629);
xnor U7667 (N_7667,N_7507,N_7537);
xnor U7668 (N_7668,N_7510,N_7630);
nor U7669 (N_7669,N_7581,N_7502);
nand U7670 (N_7670,N_7543,N_7646);
xnor U7671 (N_7671,N_7615,N_7577);
and U7672 (N_7672,N_7597,N_7634);
or U7673 (N_7673,N_7513,N_7569);
nor U7674 (N_7674,N_7605,N_7551);
nand U7675 (N_7675,N_7506,N_7558);
nand U7676 (N_7676,N_7557,N_7528);
or U7677 (N_7677,N_7644,N_7648);
nand U7678 (N_7678,N_7534,N_7616);
or U7679 (N_7679,N_7582,N_7521);
or U7680 (N_7680,N_7633,N_7617);
xor U7681 (N_7681,N_7595,N_7614);
nor U7682 (N_7682,N_7546,N_7517);
xnor U7683 (N_7683,N_7545,N_7562);
xnor U7684 (N_7684,N_7529,N_7532);
xnor U7685 (N_7685,N_7618,N_7573);
xnor U7686 (N_7686,N_7575,N_7591);
or U7687 (N_7687,N_7525,N_7526);
or U7688 (N_7688,N_7621,N_7610);
nor U7689 (N_7689,N_7626,N_7512);
nor U7690 (N_7690,N_7596,N_7602);
or U7691 (N_7691,N_7584,N_7604);
and U7692 (N_7692,N_7623,N_7609);
xnor U7693 (N_7693,N_7592,N_7540);
nand U7694 (N_7694,N_7647,N_7552);
and U7695 (N_7695,N_7603,N_7640);
xnor U7696 (N_7696,N_7500,N_7518);
and U7697 (N_7697,N_7593,N_7645);
and U7698 (N_7698,N_7563,N_7588);
nand U7699 (N_7699,N_7566,N_7561);
and U7700 (N_7700,N_7509,N_7612);
or U7701 (N_7701,N_7559,N_7567);
or U7702 (N_7702,N_7539,N_7553);
nand U7703 (N_7703,N_7514,N_7600);
or U7704 (N_7704,N_7594,N_7578);
nand U7705 (N_7705,N_7522,N_7606);
and U7706 (N_7706,N_7531,N_7583);
xor U7707 (N_7707,N_7548,N_7536);
nor U7708 (N_7708,N_7501,N_7641);
and U7709 (N_7709,N_7639,N_7503);
nand U7710 (N_7710,N_7541,N_7627);
and U7711 (N_7711,N_7642,N_7538);
and U7712 (N_7712,N_7505,N_7643);
or U7713 (N_7713,N_7530,N_7622);
and U7714 (N_7714,N_7598,N_7520);
nor U7715 (N_7715,N_7580,N_7504);
and U7716 (N_7716,N_7571,N_7599);
nor U7717 (N_7717,N_7544,N_7508);
and U7718 (N_7718,N_7637,N_7576);
and U7719 (N_7719,N_7619,N_7635);
and U7720 (N_7720,N_7555,N_7601);
xor U7721 (N_7721,N_7572,N_7632);
nor U7722 (N_7722,N_7589,N_7564);
and U7723 (N_7723,N_7535,N_7586);
nor U7724 (N_7724,N_7585,N_7607);
nand U7725 (N_7725,N_7613,N_7596);
and U7726 (N_7726,N_7577,N_7645);
and U7727 (N_7727,N_7571,N_7607);
and U7728 (N_7728,N_7544,N_7505);
or U7729 (N_7729,N_7612,N_7578);
xnor U7730 (N_7730,N_7568,N_7636);
and U7731 (N_7731,N_7518,N_7633);
xor U7732 (N_7732,N_7509,N_7572);
nor U7733 (N_7733,N_7631,N_7580);
xor U7734 (N_7734,N_7560,N_7630);
xor U7735 (N_7735,N_7603,N_7587);
or U7736 (N_7736,N_7607,N_7600);
xor U7737 (N_7737,N_7583,N_7572);
nor U7738 (N_7738,N_7539,N_7537);
or U7739 (N_7739,N_7563,N_7645);
nor U7740 (N_7740,N_7502,N_7533);
and U7741 (N_7741,N_7596,N_7554);
xor U7742 (N_7742,N_7640,N_7569);
nor U7743 (N_7743,N_7648,N_7568);
nand U7744 (N_7744,N_7588,N_7577);
or U7745 (N_7745,N_7614,N_7543);
nor U7746 (N_7746,N_7572,N_7649);
nor U7747 (N_7747,N_7568,N_7621);
and U7748 (N_7748,N_7639,N_7584);
nand U7749 (N_7749,N_7537,N_7640);
and U7750 (N_7750,N_7598,N_7506);
nand U7751 (N_7751,N_7530,N_7612);
xor U7752 (N_7752,N_7581,N_7617);
nor U7753 (N_7753,N_7646,N_7648);
xor U7754 (N_7754,N_7590,N_7562);
nor U7755 (N_7755,N_7554,N_7557);
and U7756 (N_7756,N_7555,N_7618);
nand U7757 (N_7757,N_7635,N_7593);
nand U7758 (N_7758,N_7642,N_7543);
and U7759 (N_7759,N_7580,N_7593);
and U7760 (N_7760,N_7539,N_7546);
nand U7761 (N_7761,N_7620,N_7550);
nand U7762 (N_7762,N_7604,N_7510);
nand U7763 (N_7763,N_7575,N_7521);
and U7764 (N_7764,N_7601,N_7551);
or U7765 (N_7765,N_7579,N_7527);
xor U7766 (N_7766,N_7634,N_7588);
and U7767 (N_7767,N_7509,N_7598);
and U7768 (N_7768,N_7607,N_7559);
nand U7769 (N_7769,N_7615,N_7568);
nor U7770 (N_7770,N_7585,N_7547);
nand U7771 (N_7771,N_7538,N_7521);
and U7772 (N_7772,N_7645,N_7515);
and U7773 (N_7773,N_7519,N_7552);
xor U7774 (N_7774,N_7541,N_7584);
or U7775 (N_7775,N_7576,N_7638);
nand U7776 (N_7776,N_7555,N_7571);
nor U7777 (N_7777,N_7567,N_7504);
and U7778 (N_7778,N_7531,N_7597);
and U7779 (N_7779,N_7565,N_7553);
or U7780 (N_7780,N_7624,N_7502);
nor U7781 (N_7781,N_7527,N_7648);
nor U7782 (N_7782,N_7504,N_7513);
and U7783 (N_7783,N_7527,N_7550);
nand U7784 (N_7784,N_7600,N_7599);
xnor U7785 (N_7785,N_7560,N_7570);
and U7786 (N_7786,N_7555,N_7556);
and U7787 (N_7787,N_7639,N_7624);
and U7788 (N_7788,N_7521,N_7626);
nor U7789 (N_7789,N_7641,N_7536);
and U7790 (N_7790,N_7597,N_7510);
and U7791 (N_7791,N_7576,N_7560);
and U7792 (N_7792,N_7569,N_7561);
xor U7793 (N_7793,N_7564,N_7544);
and U7794 (N_7794,N_7605,N_7612);
or U7795 (N_7795,N_7538,N_7633);
or U7796 (N_7796,N_7555,N_7512);
nor U7797 (N_7797,N_7506,N_7516);
xnor U7798 (N_7798,N_7608,N_7637);
and U7799 (N_7799,N_7643,N_7615);
nand U7800 (N_7800,N_7673,N_7695);
nor U7801 (N_7801,N_7774,N_7767);
nor U7802 (N_7802,N_7758,N_7656);
or U7803 (N_7803,N_7776,N_7731);
xnor U7804 (N_7804,N_7697,N_7766);
nand U7805 (N_7805,N_7797,N_7718);
nor U7806 (N_7806,N_7662,N_7747);
or U7807 (N_7807,N_7721,N_7663);
or U7808 (N_7808,N_7678,N_7763);
nand U7809 (N_7809,N_7730,N_7769);
nor U7810 (N_7810,N_7729,N_7712);
nor U7811 (N_7811,N_7707,N_7764);
nand U7812 (N_7812,N_7714,N_7740);
xnor U7813 (N_7813,N_7736,N_7752);
xor U7814 (N_7814,N_7798,N_7787);
nand U7815 (N_7815,N_7779,N_7675);
nor U7816 (N_7816,N_7761,N_7759);
nand U7817 (N_7817,N_7749,N_7667);
nor U7818 (N_7818,N_7658,N_7681);
xor U7819 (N_7819,N_7699,N_7757);
nand U7820 (N_7820,N_7724,N_7708);
nor U7821 (N_7821,N_7743,N_7711);
xnor U7822 (N_7822,N_7703,N_7795);
or U7823 (N_7823,N_7702,N_7670);
or U7824 (N_7824,N_7683,N_7793);
or U7825 (N_7825,N_7772,N_7783);
nand U7826 (N_7826,N_7799,N_7684);
nor U7827 (N_7827,N_7728,N_7704);
or U7828 (N_7828,N_7720,N_7796);
or U7829 (N_7829,N_7690,N_7732);
nand U7830 (N_7830,N_7741,N_7661);
and U7831 (N_7831,N_7786,N_7660);
and U7832 (N_7832,N_7745,N_7782);
or U7833 (N_7833,N_7692,N_7655);
and U7834 (N_7834,N_7737,N_7685);
or U7835 (N_7835,N_7665,N_7751);
nand U7836 (N_7836,N_7746,N_7686);
and U7837 (N_7837,N_7722,N_7719);
nor U7838 (N_7838,N_7778,N_7755);
nor U7839 (N_7839,N_7725,N_7726);
or U7840 (N_7840,N_7689,N_7753);
nand U7841 (N_7841,N_7671,N_7768);
xor U7842 (N_7842,N_7693,N_7713);
and U7843 (N_7843,N_7657,N_7676);
and U7844 (N_7844,N_7794,N_7742);
nor U7845 (N_7845,N_7669,N_7650);
or U7846 (N_7846,N_7748,N_7727);
nand U7847 (N_7847,N_7674,N_7754);
or U7848 (N_7848,N_7654,N_7760);
or U7849 (N_7849,N_7750,N_7785);
xnor U7850 (N_7850,N_7775,N_7710);
or U7851 (N_7851,N_7700,N_7706);
xnor U7852 (N_7852,N_7739,N_7780);
nor U7853 (N_7853,N_7738,N_7698);
xnor U7854 (N_7854,N_7672,N_7664);
or U7855 (N_7855,N_7659,N_7696);
or U7856 (N_7856,N_7705,N_7691);
xnor U7857 (N_7857,N_7709,N_7687);
and U7858 (N_7858,N_7789,N_7715);
nand U7859 (N_7859,N_7701,N_7668);
nand U7860 (N_7860,N_7762,N_7733);
and U7861 (N_7861,N_7680,N_7717);
or U7862 (N_7862,N_7781,N_7677);
or U7863 (N_7863,N_7679,N_7694);
xor U7864 (N_7864,N_7788,N_7784);
nand U7865 (N_7865,N_7790,N_7682);
or U7866 (N_7866,N_7744,N_7653);
nand U7867 (N_7867,N_7723,N_7792);
nor U7868 (N_7868,N_7756,N_7666);
or U7869 (N_7869,N_7765,N_7716);
or U7870 (N_7870,N_7770,N_7773);
and U7871 (N_7871,N_7652,N_7688);
nand U7872 (N_7872,N_7735,N_7791);
and U7873 (N_7873,N_7777,N_7734);
xor U7874 (N_7874,N_7771,N_7651);
nor U7875 (N_7875,N_7773,N_7789);
nand U7876 (N_7876,N_7675,N_7727);
xor U7877 (N_7877,N_7744,N_7661);
nor U7878 (N_7878,N_7656,N_7746);
and U7879 (N_7879,N_7708,N_7662);
xor U7880 (N_7880,N_7780,N_7725);
nor U7881 (N_7881,N_7693,N_7654);
xnor U7882 (N_7882,N_7691,N_7732);
xnor U7883 (N_7883,N_7664,N_7730);
nand U7884 (N_7884,N_7658,N_7746);
or U7885 (N_7885,N_7659,N_7725);
nor U7886 (N_7886,N_7740,N_7735);
and U7887 (N_7887,N_7763,N_7691);
and U7888 (N_7888,N_7742,N_7778);
or U7889 (N_7889,N_7766,N_7735);
nand U7890 (N_7890,N_7680,N_7670);
nor U7891 (N_7891,N_7678,N_7687);
or U7892 (N_7892,N_7744,N_7707);
xor U7893 (N_7893,N_7707,N_7653);
nor U7894 (N_7894,N_7689,N_7748);
xnor U7895 (N_7895,N_7666,N_7711);
and U7896 (N_7896,N_7703,N_7717);
or U7897 (N_7897,N_7694,N_7768);
nand U7898 (N_7898,N_7675,N_7673);
nand U7899 (N_7899,N_7761,N_7672);
nor U7900 (N_7900,N_7671,N_7664);
nand U7901 (N_7901,N_7785,N_7720);
and U7902 (N_7902,N_7651,N_7695);
xnor U7903 (N_7903,N_7710,N_7664);
xor U7904 (N_7904,N_7762,N_7659);
xor U7905 (N_7905,N_7683,N_7709);
nand U7906 (N_7906,N_7674,N_7718);
nand U7907 (N_7907,N_7782,N_7686);
nand U7908 (N_7908,N_7770,N_7669);
xor U7909 (N_7909,N_7772,N_7782);
or U7910 (N_7910,N_7677,N_7780);
nor U7911 (N_7911,N_7706,N_7684);
xor U7912 (N_7912,N_7677,N_7691);
and U7913 (N_7913,N_7677,N_7770);
nor U7914 (N_7914,N_7670,N_7732);
xor U7915 (N_7915,N_7793,N_7710);
xnor U7916 (N_7916,N_7700,N_7753);
xor U7917 (N_7917,N_7761,N_7786);
xor U7918 (N_7918,N_7779,N_7794);
nor U7919 (N_7919,N_7714,N_7664);
and U7920 (N_7920,N_7660,N_7726);
nand U7921 (N_7921,N_7772,N_7681);
or U7922 (N_7922,N_7728,N_7707);
and U7923 (N_7923,N_7758,N_7760);
or U7924 (N_7924,N_7770,N_7673);
nor U7925 (N_7925,N_7792,N_7702);
and U7926 (N_7926,N_7768,N_7665);
or U7927 (N_7927,N_7682,N_7694);
nor U7928 (N_7928,N_7797,N_7670);
nand U7929 (N_7929,N_7745,N_7796);
xor U7930 (N_7930,N_7767,N_7742);
nor U7931 (N_7931,N_7789,N_7707);
or U7932 (N_7932,N_7784,N_7763);
or U7933 (N_7933,N_7675,N_7746);
and U7934 (N_7934,N_7759,N_7760);
or U7935 (N_7935,N_7697,N_7659);
nand U7936 (N_7936,N_7758,N_7685);
nor U7937 (N_7937,N_7722,N_7769);
or U7938 (N_7938,N_7771,N_7752);
nand U7939 (N_7939,N_7727,N_7766);
or U7940 (N_7940,N_7677,N_7695);
or U7941 (N_7941,N_7716,N_7656);
nor U7942 (N_7942,N_7727,N_7713);
and U7943 (N_7943,N_7796,N_7783);
xor U7944 (N_7944,N_7681,N_7780);
or U7945 (N_7945,N_7750,N_7689);
nand U7946 (N_7946,N_7743,N_7715);
nand U7947 (N_7947,N_7664,N_7720);
nor U7948 (N_7948,N_7771,N_7698);
and U7949 (N_7949,N_7738,N_7741);
and U7950 (N_7950,N_7899,N_7898);
or U7951 (N_7951,N_7934,N_7849);
nor U7952 (N_7952,N_7812,N_7817);
xor U7953 (N_7953,N_7897,N_7831);
or U7954 (N_7954,N_7815,N_7895);
or U7955 (N_7955,N_7819,N_7901);
or U7956 (N_7956,N_7829,N_7884);
and U7957 (N_7957,N_7919,N_7857);
xnor U7958 (N_7958,N_7927,N_7896);
nand U7959 (N_7959,N_7844,N_7835);
and U7960 (N_7960,N_7802,N_7940);
and U7961 (N_7961,N_7949,N_7843);
xor U7962 (N_7962,N_7839,N_7830);
xor U7963 (N_7963,N_7912,N_7865);
or U7964 (N_7964,N_7806,N_7929);
or U7965 (N_7965,N_7862,N_7905);
nor U7966 (N_7966,N_7917,N_7832);
xor U7967 (N_7967,N_7921,N_7931);
and U7968 (N_7968,N_7932,N_7805);
or U7969 (N_7969,N_7800,N_7878);
xor U7970 (N_7970,N_7814,N_7892);
or U7971 (N_7971,N_7811,N_7913);
or U7972 (N_7972,N_7883,N_7856);
or U7973 (N_7973,N_7942,N_7904);
xor U7974 (N_7974,N_7861,N_7869);
or U7975 (N_7975,N_7909,N_7920);
and U7976 (N_7976,N_7941,N_7885);
nand U7977 (N_7977,N_7866,N_7876);
and U7978 (N_7978,N_7828,N_7890);
nor U7979 (N_7979,N_7947,N_7891);
and U7980 (N_7980,N_7807,N_7848);
nor U7981 (N_7981,N_7834,N_7825);
nand U7982 (N_7982,N_7855,N_7821);
xor U7983 (N_7983,N_7922,N_7945);
and U7984 (N_7984,N_7881,N_7889);
nand U7985 (N_7985,N_7930,N_7933);
and U7986 (N_7986,N_7859,N_7810);
or U7987 (N_7987,N_7867,N_7935);
nor U7988 (N_7988,N_7928,N_7874);
or U7989 (N_7989,N_7937,N_7915);
and U7990 (N_7990,N_7804,N_7880);
xnor U7991 (N_7991,N_7864,N_7902);
nor U7992 (N_7992,N_7946,N_7841);
nand U7993 (N_7993,N_7826,N_7916);
xor U7994 (N_7994,N_7836,N_7944);
xnor U7995 (N_7995,N_7854,N_7906);
xor U7996 (N_7996,N_7850,N_7939);
and U7997 (N_7997,N_7833,N_7816);
or U7998 (N_7998,N_7840,N_7853);
or U7999 (N_7999,N_7893,N_7914);
and U8000 (N_8000,N_7910,N_7938);
nand U8001 (N_8001,N_7948,N_7923);
nor U8002 (N_8002,N_7871,N_7801);
nor U8003 (N_8003,N_7863,N_7943);
nor U8004 (N_8004,N_7907,N_7936);
or U8005 (N_8005,N_7809,N_7908);
nor U8006 (N_8006,N_7847,N_7877);
nor U8007 (N_8007,N_7879,N_7822);
nor U8008 (N_8008,N_7924,N_7870);
nand U8009 (N_8009,N_7845,N_7808);
and U8010 (N_8010,N_7813,N_7803);
or U8011 (N_8011,N_7827,N_7887);
xor U8012 (N_8012,N_7868,N_7837);
and U8013 (N_8013,N_7875,N_7925);
nand U8014 (N_8014,N_7888,N_7911);
nor U8015 (N_8015,N_7823,N_7851);
or U8016 (N_8016,N_7838,N_7882);
nor U8017 (N_8017,N_7842,N_7918);
nor U8018 (N_8018,N_7824,N_7860);
nand U8019 (N_8019,N_7900,N_7873);
or U8020 (N_8020,N_7903,N_7894);
xor U8021 (N_8021,N_7852,N_7858);
or U8022 (N_8022,N_7846,N_7818);
or U8023 (N_8023,N_7820,N_7926);
xor U8024 (N_8024,N_7872,N_7886);
or U8025 (N_8025,N_7924,N_7881);
or U8026 (N_8026,N_7909,N_7899);
and U8027 (N_8027,N_7865,N_7934);
nand U8028 (N_8028,N_7861,N_7880);
nand U8029 (N_8029,N_7806,N_7911);
or U8030 (N_8030,N_7838,N_7880);
nand U8031 (N_8031,N_7820,N_7899);
and U8032 (N_8032,N_7883,N_7811);
nor U8033 (N_8033,N_7865,N_7817);
and U8034 (N_8034,N_7801,N_7899);
and U8035 (N_8035,N_7923,N_7872);
nand U8036 (N_8036,N_7908,N_7888);
or U8037 (N_8037,N_7873,N_7806);
nor U8038 (N_8038,N_7922,N_7930);
or U8039 (N_8039,N_7868,N_7853);
xnor U8040 (N_8040,N_7867,N_7837);
and U8041 (N_8041,N_7899,N_7907);
nor U8042 (N_8042,N_7875,N_7935);
xor U8043 (N_8043,N_7903,N_7896);
nor U8044 (N_8044,N_7827,N_7871);
or U8045 (N_8045,N_7831,N_7924);
nor U8046 (N_8046,N_7843,N_7849);
nand U8047 (N_8047,N_7915,N_7807);
or U8048 (N_8048,N_7840,N_7949);
or U8049 (N_8049,N_7830,N_7819);
xor U8050 (N_8050,N_7890,N_7941);
nand U8051 (N_8051,N_7821,N_7891);
nand U8052 (N_8052,N_7895,N_7880);
nand U8053 (N_8053,N_7893,N_7856);
nor U8054 (N_8054,N_7805,N_7935);
xor U8055 (N_8055,N_7871,N_7821);
nand U8056 (N_8056,N_7910,N_7802);
and U8057 (N_8057,N_7883,N_7909);
xnor U8058 (N_8058,N_7911,N_7851);
or U8059 (N_8059,N_7875,N_7910);
or U8060 (N_8060,N_7944,N_7818);
nand U8061 (N_8061,N_7931,N_7846);
xor U8062 (N_8062,N_7903,N_7892);
and U8063 (N_8063,N_7942,N_7918);
and U8064 (N_8064,N_7922,N_7834);
and U8065 (N_8065,N_7892,N_7904);
or U8066 (N_8066,N_7845,N_7903);
and U8067 (N_8067,N_7903,N_7919);
or U8068 (N_8068,N_7924,N_7916);
xor U8069 (N_8069,N_7803,N_7845);
nor U8070 (N_8070,N_7930,N_7934);
nand U8071 (N_8071,N_7937,N_7896);
or U8072 (N_8072,N_7821,N_7885);
nand U8073 (N_8073,N_7881,N_7914);
or U8074 (N_8074,N_7825,N_7876);
nand U8075 (N_8075,N_7817,N_7828);
or U8076 (N_8076,N_7923,N_7939);
or U8077 (N_8077,N_7863,N_7891);
and U8078 (N_8078,N_7940,N_7820);
nor U8079 (N_8079,N_7935,N_7810);
nand U8080 (N_8080,N_7802,N_7886);
nor U8081 (N_8081,N_7855,N_7891);
and U8082 (N_8082,N_7893,N_7895);
xor U8083 (N_8083,N_7810,N_7906);
nand U8084 (N_8084,N_7945,N_7903);
nor U8085 (N_8085,N_7868,N_7830);
xor U8086 (N_8086,N_7826,N_7869);
nor U8087 (N_8087,N_7872,N_7888);
and U8088 (N_8088,N_7898,N_7822);
nor U8089 (N_8089,N_7922,N_7855);
or U8090 (N_8090,N_7871,N_7811);
xnor U8091 (N_8091,N_7916,N_7842);
xor U8092 (N_8092,N_7899,N_7901);
xnor U8093 (N_8093,N_7862,N_7946);
and U8094 (N_8094,N_7940,N_7911);
nand U8095 (N_8095,N_7866,N_7938);
xnor U8096 (N_8096,N_7897,N_7802);
nor U8097 (N_8097,N_7876,N_7821);
nand U8098 (N_8098,N_7802,N_7889);
xnor U8099 (N_8099,N_7803,N_7911);
xor U8100 (N_8100,N_7970,N_7983);
or U8101 (N_8101,N_8001,N_8067);
nor U8102 (N_8102,N_8051,N_7950);
and U8103 (N_8103,N_8084,N_7977);
and U8104 (N_8104,N_7951,N_7986);
nor U8105 (N_8105,N_8025,N_7988);
xnor U8106 (N_8106,N_8070,N_8064);
nor U8107 (N_8107,N_8020,N_7989);
xnor U8108 (N_8108,N_7958,N_7961);
xnor U8109 (N_8109,N_8037,N_7987);
xor U8110 (N_8110,N_8046,N_8006);
or U8111 (N_8111,N_7990,N_8082);
nand U8112 (N_8112,N_8017,N_8056);
xor U8113 (N_8113,N_8000,N_8054);
nand U8114 (N_8114,N_7996,N_7981);
and U8115 (N_8115,N_8031,N_8069);
nor U8116 (N_8116,N_8048,N_8087);
nand U8117 (N_8117,N_8041,N_8049);
and U8118 (N_8118,N_8095,N_7968);
and U8119 (N_8119,N_7992,N_8066);
xor U8120 (N_8120,N_7999,N_8027);
or U8121 (N_8121,N_7971,N_8080);
nand U8122 (N_8122,N_7975,N_8032);
and U8123 (N_8123,N_8086,N_7960);
nor U8124 (N_8124,N_8085,N_7974);
nor U8125 (N_8125,N_7953,N_8058);
nor U8126 (N_8126,N_8077,N_8047);
nand U8127 (N_8127,N_8030,N_8091);
or U8128 (N_8128,N_7997,N_8038);
nand U8129 (N_8129,N_8013,N_8022);
xnor U8130 (N_8130,N_8083,N_8063);
xor U8131 (N_8131,N_8026,N_8097);
nand U8132 (N_8132,N_8061,N_8043);
xor U8133 (N_8133,N_8023,N_7980);
or U8134 (N_8134,N_8015,N_7964);
or U8135 (N_8135,N_8018,N_8014);
xor U8136 (N_8136,N_8042,N_8005);
xor U8137 (N_8137,N_8050,N_8028);
nand U8138 (N_8138,N_8019,N_8002);
nand U8139 (N_8139,N_7985,N_8081);
nand U8140 (N_8140,N_7965,N_8016);
xor U8141 (N_8141,N_8008,N_8099);
xnor U8142 (N_8142,N_8059,N_8040);
nor U8143 (N_8143,N_8076,N_8089);
nand U8144 (N_8144,N_8052,N_8065);
xnor U8145 (N_8145,N_8045,N_7954);
nand U8146 (N_8146,N_8075,N_8039);
nor U8147 (N_8147,N_8012,N_7973);
or U8148 (N_8148,N_8033,N_8034);
nor U8149 (N_8149,N_8062,N_8094);
nor U8150 (N_8150,N_8071,N_8021);
and U8151 (N_8151,N_8088,N_8024);
xnor U8152 (N_8152,N_8072,N_8010);
xor U8153 (N_8153,N_8074,N_7956);
nand U8154 (N_8154,N_8057,N_8090);
and U8155 (N_8155,N_8035,N_8009);
nand U8156 (N_8156,N_8079,N_7972);
xor U8157 (N_8157,N_8053,N_7967);
or U8158 (N_8158,N_7966,N_7994);
and U8159 (N_8159,N_8093,N_8029);
nand U8160 (N_8160,N_7959,N_7969);
and U8161 (N_8161,N_8098,N_8055);
and U8162 (N_8162,N_7955,N_7995);
nor U8163 (N_8163,N_8044,N_7984);
nor U8164 (N_8164,N_8092,N_7982);
and U8165 (N_8165,N_8078,N_8060);
nand U8166 (N_8166,N_8068,N_8003);
nand U8167 (N_8167,N_7991,N_7952);
or U8168 (N_8168,N_8004,N_7962);
and U8169 (N_8169,N_7978,N_8007);
nor U8170 (N_8170,N_7979,N_7976);
xor U8171 (N_8171,N_8036,N_7993);
nand U8172 (N_8172,N_7998,N_7963);
or U8173 (N_8173,N_8011,N_7957);
and U8174 (N_8174,N_8096,N_8073);
nand U8175 (N_8175,N_7977,N_8086);
nand U8176 (N_8176,N_7987,N_7965);
nor U8177 (N_8177,N_8057,N_8096);
or U8178 (N_8178,N_7954,N_7999);
and U8179 (N_8179,N_7959,N_8014);
nor U8180 (N_8180,N_8088,N_7977);
and U8181 (N_8181,N_7966,N_8093);
nor U8182 (N_8182,N_7955,N_8040);
nand U8183 (N_8183,N_8044,N_8053);
or U8184 (N_8184,N_8011,N_8072);
xnor U8185 (N_8185,N_8030,N_7988);
xor U8186 (N_8186,N_7980,N_8080);
and U8187 (N_8187,N_8088,N_8020);
nor U8188 (N_8188,N_8088,N_8097);
nor U8189 (N_8189,N_8051,N_8046);
and U8190 (N_8190,N_8009,N_8028);
nand U8191 (N_8191,N_8086,N_8044);
xor U8192 (N_8192,N_8005,N_7958);
or U8193 (N_8193,N_8017,N_8036);
xor U8194 (N_8194,N_7956,N_8093);
xnor U8195 (N_8195,N_7974,N_8064);
and U8196 (N_8196,N_7977,N_8073);
nand U8197 (N_8197,N_7953,N_7985);
nor U8198 (N_8198,N_8008,N_8040);
or U8199 (N_8199,N_8068,N_7964);
and U8200 (N_8200,N_8059,N_7985);
nor U8201 (N_8201,N_7955,N_8096);
nor U8202 (N_8202,N_8066,N_7966);
and U8203 (N_8203,N_8055,N_7973);
xnor U8204 (N_8204,N_8078,N_8064);
nor U8205 (N_8205,N_8081,N_8094);
nand U8206 (N_8206,N_7956,N_7981);
nor U8207 (N_8207,N_8046,N_7984);
xnor U8208 (N_8208,N_7999,N_8099);
nand U8209 (N_8209,N_8098,N_8028);
nand U8210 (N_8210,N_7996,N_7956);
or U8211 (N_8211,N_7974,N_8099);
nand U8212 (N_8212,N_8042,N_7969);
nor U8213 (N_8213,N_7988,N_8005);
xnor U8214 (N_8214,N_8000,N_7954);
nand U8215 (N_8215,N_8095,N_7967);
nor U8216 (N_8216,N_7961,N_8048);
and U8217 (N_8217,N_8029,N_8088);
or U8218 (N_8218,N_8058,N_7962);
and U8219 (N_8219,N_7975,N_8094);
and U8220 (N_8220,N_8031,N_8010);
nor U8221 (N_8221,N_8025,N_7997);
and U8222 (N_8222,N_8028,N_7974);
or U8223 (N_8223,N_7960,N_7986);
xor U8224 (N_8224,N_8049,N_8099);
or U8225 (N_8225,N_8051,N_7999);
xor U8226 (N_8226,N_8058,N_8078);
nor U8227 (N_8227,N_8012,N_8004);
and U8228 (N_8228,N_7998,N_8022);
nor U8229 (N_8229,N_8049,N_8019);
nand U8230 (N_8230,N_8073,N_7978);
or U8231 (N_8231,N_7986,N_8065);
nand U8232 (N_8232,N_7964,N_8018);
or U8233 (N_8233,N_7992,N_8081);
and U8234 (N_8234,N_8075,N_8019);
nor U8235 (N_8235,N_7961,N_8042);
and U8236 (N_8236,N_8065,N_8002);
or U8237 (N_8237,N_8072,N_8087);
nor U8238 (N_8238,N_8015,N_8027);
nand U8239 (N_8239,N_8050,N_8086);
nand U8240 (N_8240,N_8095,N_7956);
xnor U8241 (N_8241,N_8012,N_8006);
nor U8242 (N_8242,N_7968,N_7960);
and U8243 (N_8243,N_8045,N_7959);
xor U8244 (N_8244,N_8010,N_7965);
nand U8245 (N_8245,N_8026,N_7985);
and U8246 (N_8246,N_8054,N_8045);
nor U8247 (N_8247,N_8002,N_8075);
nand U8248 (N_8248,N_8086,N_8006);
nor U8249 (N_8249,N_8048,N_7958);
or U8250 (N_8250,N_8163,N_8248);
nand U8251 (N_8251,N_8121,N_8180);
and U8252 (N_8252,N_8198,N_8210);
or U8253 (N_8253,N_8150,N_8201);
nand U8254 (N_8254,N_8179,N_8161);
nor U8255 (N_8255,N_8192,N_8159);
xor U8256 (N_8256,N_8177,N_8129);
nand U8257 (N_8257,N_8138,N_8249);
nor U8258 (N_8258,N_8173,N_8125);
and U8259 (N_8259,N_8244,N_8184);
and U8260 (N_8260,N_8145,N_8170);
nand U8261 (N_8261,N_8228,N_8186);
nor U8262 (N_8262,N_8220,N_8223);
and U8263 (N_8263,N_8225,N_8115);
nand U8264 (N_8264,N_8117,N_8128);
or U8265 (N_8265,N_8221,N_8200);
or U8266 (N_8266,N_8230,N_8235);
nor U8267 (N_8267,N_8151,N_8234);
xnor U8268 (N_8268,N_8156,N_8116);
nor U8269 (N_8269,N_8136,N_8175);
or U8270 (N_8270,N_8229,N_8188);
and U8271 (N_8271,N_8133,N_8135);
and U8272 (N_8272,N_8101,N_8106);
and U8273 (N_8273,N_8141,N_8119);
nand U8274 (N_8274,N_8158,N_8222);
nand U8275 (N_8275,N_8213,N_8237);
or U8276 (N_8276,N_8105,N_8144);
nand U8277 (N_8277,N_8155,N_8242);
or U8278 (N_8278,N_8189,N_8187);
xor U8279 (N_8279,N_8236,N_8232);
nor U8280 (N_8280,N_8137,N_8169);
or U8281 (N_8281,N_8181,N_8131);
nor U8282 (N_8282,N_8238,N_8217);
or U8283 (N_8283,N_8182,N_8108);
nor U8284 (N_8284,N_8203,N_8195);
or U8285 (N_8285,N_8174,N_8172);
nor U8286 (N_8286,N_8111,N_8227);
and U8287 (N_8287,N_8212,N_8240);
or U8288 (N_8288,N_8152,N_8123);
and U8289 (N_8289,N_8214,N_8218);
xnor U8290 (N_8290,N_8168,N_8239);
nand U8291 (N_8291,N_8211,N_8196);
or U8292 (N_8292,N_8208,N_8202);
or U8293 (N_8293,N_8103,N_8219);
nor U8294 (N_8294,N_8148,N_8110);
and U8295 (N_8295,N_8139,N_8157);
or U8296 (N_8296,N_8113,N_8215);
nor U8297 (N_8297,N_8231,N_8246);
and U8298 (N_8298,N_8224,N_8216);
and U8299 (N_8299,N_8143,N_8226);
nand U8300 (N_8300,N_8140,N_8132);
and U8301 (N_8301,N_8191,N_8160);
nand U8302 (N_8302,N_8171,N_8164);
or U8303 (N_8303,N_8104,N_8190);
and U8304 (N_8304,N_8134,N_8100);
xnor U8305 (N_8305,N_8162,N_8166);
or U8306 (N_8306,N_8241,N_8178);
or U8307 (N_8307,N_8127,N_8153);
and U8308 (N_8308,N_8146,N_8165);
or U8309 (N_8309,N_8243,N_8114);
and U8310 (N_8310,N_8245,N_8122);
and U8311 (N_8311,N_8124,N_8109);
or U8312 (N_8312,N_8197,N_8183);
or U8313 (N_8313,N_8147,N_8176);
xnor U8314 (N_8314,N_8154,N_8193);
nand U8315 (N_8315,N_8204,N_8107);
or U8316 (N_8316,N_8194,N_8112);
nand U8317 (N_8317,N_8205,N_8207);
and U8318 (N_8318,N_8118,N_8206);
or U8319 (N_8319,N_8247,N_8120);
or U8320 (N_8320,N_8185,N_8233);
nand U8321 (N_8321,N_8142,N_8167);
nand U8322 (N_8322,N_8102,N_8209);
xnor U8323 (N_8323,N_8199,N_8149);
nand U8324 (N_8324,N_8126,N_8130);
or U8325 (N_8325,N_8162,N_8137);
or U8326 (N_8326,N_8150,N_8171);
nor U8327 (N_8327,N_8131,N_8238);
or U8328 (N_8328,N_8144,N_8202);
nand U8329 (N_8329,N_8195,N_8173);
nand U8330 (N_8330,N_8176,N_8222);
and U8331 (N_8331,N_8175,N_8141);
nor U8332 (N_8332,N_8123,N_8244);
nor U8333 (N_8333,N_8103,N_8238);
or U8334 (N_8334,N_8126,N_8129);
and U8335 (N_8335,N_8173,N_8231);
or U8336 (N_8336,N_8177,N_8119);
nand U8337 (N_8337,N_8245,N_8105);
or U8338 (N_8338,N_8223,N_8203);
and U8339 (N_8339,N_8131,N_8228);
xor U8340 (N_8340,N_8144,N_8245);
nand U8341 (N_8341,N_8174,N_8246);
or U8342 (N_8342,N_8171,N_8182);
or U8343 (N_8343,N_8165,N_8241);
nor U8344 (N_8344,N_8225,N_8139);
or U8345 (N_8345,N_8178,N_8174);
and U8346 (N_8346,N_8103,N_8239);
xnor U8347 (N_8347,N_8177,N_8101);
or U8348 (N_8348,N_8179,N_8208);
and U8349 (N_8349,N_8189,N_8169);
or U8350 (N_8350,N_8210,N_8201);
and U8351 (N_8351,N_8179,N_8213);
and U8352 (N_8352,N_8127,N_8243);
or U8353 (N_8353,N_8190,N_8207);
and U8354 (N_8354,N_8165,N_8192);
and U8355 (N_8355,N_8235,N_8171);
and U8356 (N_8356,N_8212,N_8155);
nor U8357 (N_8357,N_8155,N_8188);
and U8358 (N_8358,N_8210,N_8224);
nand U8359 (N_8359,N_8161,N_8180);
nand U8360 (N_8360,N_8144,N_8216);
and U8361 (N_8361,N_8169,N_8153);
or U8362 (N_8362,N_8233,N_8238);
nand U8363 (N_8363,N_8198,N_8160);
nand U8364 (N_8364,N_8139,N_8246);
nand U8365 (N_8365,N_8223,N_8211);
or U8366 (N_8366,N_8174,N_8116);
nor U8367 (N_8367,N_8210,N_8238);
and U8368 (N_8368,N_8214,N_8202);
nand U8369 (N_8369,N_8241,N_8117);
xor U8370 (N_8370,N_8187,N_8156);
xnor U8371 (N_8371,N_8141,N_8110);
nand U8372 (N_8372,N_8132,N_8197);
nor U8373 (N_8373,N_8220,N_8164);
or U8374 (N_8374,N_8179,N_8159);
nor U8375 (N_8375,N_8248,N_8240);
nand U8376 (N_8376,N_8142,N_8135);
or U8377 (N_8377,N_8231,N_8155);
and U8378 (N_8378,N_8172,N_8183);
nor U8379 (N_8379,N_8210,N_8226);
nor U8380 (N_8380,N_8155,N_8147);
nand U8381 (N_8381,N_8110,N_8173);
nand U8382 (N_8382,N_8213,N_8167);
nand U8383 (N_8383,N_8158,N_8119);
nor U8384 (N_8384,N_8239,N_8181);
and U8385 (N_8385,N_8135,N_8190);
and U8386 (N_8386,N_8101,N_8228);
xnor U8387 (N_8387,N_8206,N_8189);
nor U8388 (N_8388,N_8182,N_8214);
xnor U8389 (N_8389,N_8139,N_8153);
nand U8390 (N_8390,N_8214,N_8210);
nor U8391 (N_8391,N_8183,N_8223);
or U8392 (N_8392,N_8227,N_8210);
xor U8393 (N_8393,N_8171,N_8242);
or U8394 (N_8394,N_8161,N_8236);
or U8395 (N_8395,N_8222,N_8140);
nand U8396 (N_8396,N_8195,N_8170);
nand U8397 (N_8397,N_8138,N_8214);
nor U8398 (N_8398,N_8235,N_8155);
nor U8399 (N_8399,N_8152,N_8118);
nand U8400 (N_8400,N_8310,N_8373);
and U8401 (N_8401,N_8263,N_8375);
nand U8402 (N_8402,N_8264,N_8268);
or U8403 (N_8403,N_8385,N_8338);
and U8404 (N_8404,N_8292,N_8395);
or U8405 (N_8405,N_8289,N_8306);
nand U8406 (N_8406,N_8322,N_8293);
nor U8407 (N_8407,N_8365,N_8258);
xor U8408 (N_8408,N_8255,N_8329);
and U8409 (N_8409,N_8383,N_8314);
nand U8410 (N_8410,N_8303,N_8323);
xor U8411 (N_8411,N_8307,N_8270);
nor U8412 (N_8412,N_8282,N_8250);
nor U8413 (N_8413,N_8336,N_8257);
nor U8414 (N_8414,N_8296,N_8398);
and U8415 (N_8415,N_8388,N_8366);
and U8416 (N_8416,N_8325,N_8266);
and U8417 (N_8417,N_8315,N_8313);
or U8418 (N_8418,N_8275,N_8260);
or U8419 (N_8419,N_8335,N_8269);
nand U8420 (N_8420,N_8261,N_8284);
and U8421 (N_8421,N_8341,N_8381);
or U8422 (N_8422,N_8396,N_8386);
or U8423 (N_8423,N_8251,N_8279);
and U8424 (N_8424,N_8328,N_8276);
nand U8425 (N_8425,N_8360,N_8344);
nor U8426 (N_8426,N_8363,N_8274);
nor U8427 (N_8427,N_8354,N_8283);
and U8428 (N_8428,N_8305,N_8317);
or U8429 (N_8429,N_8297,N_8326);
xnor U8430 (N_8430,N_8308,N_8369);
xnor U8431 (N_8431,N_8343,N_8286);
and U8432 (N_8432,N_8318,N_8285);
xnor U8433 (N_8433,N_8392,N_8324);
xor U8434 (N_8434,N_8265,N_8298);
and U8435 (N_8435,N_8331,N_8330);
nand U8436 (N_8436,N_8301,N_8288);
nor U8437 (N_8437,N_8320,N_8374);
nor U8438 (N_8438,N_8281,N_8252);
or U8439 (N_8439,N_8361,N_8358);
nor U8440 (N_8440,N_8273,N_8349);
nand U8441 (N_8441,N_8347,N_8377);
nand U8442 (N_8442,N_8380,N_8372);
nor U8443 (N_8443,N_8291,N_8378);
nor U8444 (N_8444,N_8340,N_8397);
xor U8445 (N_8445,N_8253,N_8300);
or U8446 (N_8446,N_8389,N_8357);
or U8447 (N_8447,N_8394,N_8387);
nor U8448 (N_8448,N_8271,N_8370);
nor U8449 (N_8449,N_8390,N_8367);
or U8450 (N_8450,N_8254,N_8379);
and U8451 (N_8451,N_8332,N_8309);
nand U8452 (N_8452,N_8368,N_8316);
xor U8453 (N_8453,N_8259,N_8267);
nand U8454 (N_8454,N_8272,N_8327);
xnor U8455 (N_8455,N_8393,N_8339);
xor U8456 (N_8456,N_8304,N_8312);
and U8457 (N_8457,N_8311,N_8352);
or U8458 (N_8458,N_8348,N_8346);
and U8459 (N_8459,N_8345,N_8287);
nor U8460 (N_8460,N_8350,N_8319);
and U8461 (N_8461,N_8355,N_8391);
or U8462 (N_8462,N_8356,N_8302);
or U8463 (N_8463,N_8277,N_8353);
and U8464 (N_8464,N_8280,N_8290);
and U8465 (N_8465,N_8334,N_8376);
xnor U8466 (N_8466,N_8371,N_8256);
and U8467 (N_8467,N_8294,N_8362);
or U8468 (N_8468,N_8384,N_8333);
xnor U8469 (N_8469,N_8278,N_8399);
nand U8470 (N_8470,N_8364,N_8382);
nor U8471 (N_8471,N_8299,N_8262);
nor U8472 (N_8472,N_8337,N_8351);
and U8473 (N_8473,N_8295,N_8321);
nand U8474 (N_8474,N_8359,N_8342);
nand U8475 (N_8475,N_8333,N_8284);
nand U8476 (N_8476,N_8344,N_8362);
nor U8477 (N_8477,N_8256,N_8329);
nor U8478 (N_8478,N_8323,N_8370);
nor U8479 (N_8479,N_8345,N_8384);
or U8480 (N_8480,N_8323,N_8369);
nor U8481 (N_8481,N_8328,N_8319);
or U8482 (N_8482,N_8280,N_8347);
nand U8483 (N_8483,N_8305,N_8293);
xor U8484 (N_8484,N_8354,N_8396);
or U8485 (N_8485,N_8324,N_8363);
and U8486 (N_8486,N_8375,N_8347);
nand U8487 (N_8487,N_8361,N_8256);
nor U8488 (N_8488,N_8289,N_8327);
xnor U8489 (N_8489,N_8342,N_8371);
nand U8490 (N_8490,N_8262,N_8349);
xor U8491 (N_8491,N_8362,N_8368);
nor U8492 (N_8492,N_8306,N_8380);
xor U8493 (N_8493,N_8372,N_8378);
and U8494 (N_8494,N_8314,N_8324);
nor U8495 (N_8495,N_8310,N_8336);
and U8496 (N_8496,N_8307,N_8351);
or U8497 (N_8497,N_8265,N_8282);
or U8498 (N_8498,N_8335,N_8250);
nor U8499 (N_8499,N_8386,N_8324);
or U8500 (N_8500,N_8284,N_8299);
nand U8501 (N_8501,N_8320,N_8283);
and U8502 (N_8502,N_8398,N_8304);
xnor U8503 (N_8503,N_8338,N_8308);
and U8504 (N_8504,N_8296,N_8351);
and U8505 (N_8505,N_8281,N_8332);
xnor U8506 (N_8506,N_8356,N_8279);
xnor U8507 (N_8507,N_8340,N_8282);
xnor U8508 (N_8508,N_8321,N_8357);
and U8509 (N_8509,N_8260,N_8287);
or U8510 (N_8510,N_8306,N_8350);
xor U8511 (N_8511,N_8343,N_8261);
or U8512 (N_8512,N_8304,N_8369);
and U8513 (N_8513,N_8387,N_8283);
and U8514 (N_8514,N_8369,N_8305);
or U8515 (N_8515,N_8343,N_8337);
xor U8516 (N_8516,N_8290,N_8342);
xnor U8517 (N_8517,N_8316,N_8255);
and U8518 (N_8518,N_8278,N_8367);
xor U8519 (N_8519,N_8384,N_8316);
or U8520 (N_8520,N_8314,N_8331);
nor U8521 (N_8521,N_8282,N_8338);
nor U8522 (N_8522,N_8387,N_8280);
xnor U8523 (N_8523,N_8356,N_8323);
nand U8524 (N_8524,N_8251,N_8399);
or U8525 (N_8525,N_8272,N_8251);
nand U8526 (N_8526,N_8253,N_8393);
nor U8527 (N_8527,N_8268,N_8358);
xnor U8528 (N_8528,N_8272,N_8341);
nand U8529 (N_8529,N_8342,N_8328);
and U8530 (N_8530,N_8321,N_8263);
xor U8531 (N_8531,N_8399,N_8385);
or U8532 (N_8532,N_8275,N_8388);
or U8533 (N_8533,N_8384,N_8272);
nor U8534 (N_8534,N_8264,N_8259);
or U8535 (N_8535,N_8363,N_8263);
or U8536 (N_8536,N_8353,N_8292);
or U8537 (N_8537,N_8312,N_8356);
and U8538 (N_8538,N_8261,N_8372);
xnor U8539 (N_8539,N_8390,N_8375);
nand U8540 (N_8540,N_8397,N_8296);
nor U8541 (N_8541,N_8355,N_8344);
and U8542 (N_8542,N_8376,N_8377);
nor U8543 (N_8543,N_8302,N_8358);
or U8544 (N_8544,N_8318,N_8312);
xnor U8545 (N_8545,N_8275,N_8258);
nand U8546 (N_8546,N_8343,N_8396);
and U8547 (N_8547,N_8315,N_8397);
nor U8548 (N_8548,N_8372,N_8314);
and U8549 (N_8549,N_8255,N_8318);
nand U8550 (N_8550,N_8420,N_8405);
or U8551 (N_8551,N_8545,N_8506);
nor U8552 (N_8552,N_8446,N_8539);
or U8553 (N_8553,N_8406,N_8505);
nand U8554 (N_8554,N_8428,N_8458);
nand U8555 (N_8555,N_8513,N_8519);
and U8556 (N_8556,N_8426,N_8542);
nand U8557 (N_8557,N_8417,N_8415);
and U8558 (N_8558,N_8437,N_8548);
xor U8559 (N_8559,N_8477,N_8489);
xor U8560 (N_8560,N_8451,N_8461);
or U8561 (N_8561,N_8530,N_8479);
xnor U8562 (N_8562,N_8543,N_8485);
and U8563 (N_8563,N_8500,N_8510);
xnor U8564 (N_8564,N_8435,N_8464);
nor U8565 (N_8565,N_8468,N_8456);
nor U8566 (N_8566,N_8482,N_8471);
xnor U8567 (N_8567,N_8512,N_8524);
xnor U8568 (N_8568,N_8403,N_8546);
and U8569 (N_8569,N_8438,N_8425);
xor U8570 (N_8570,N_8540,N_8517);
nor U8571 (N_8571,N_8460,N_8432);
or U8572 (N_8572,N_8467,N_8503);
nand U8573 (N_8573,N_8448,N_8408);
and U8574 (N_8574,N_8527,N_8504);
xnor U8575 (N_8575,N_8535,N_8547);
nor U8576 (N_8576,N_8492,N_8533);
and U8577 (N_8577,N_8495,N_8441);
or U8578 (N_8578,N_8444,N_8526);
xnor U8579 (N_8579,N_8509,N_8515);
nand U8580 (N_8580,N_8421,N_8528);
nor U8581 (N_8581,N_8430,N_8439);
nand U8582 (N_8582,N_8499,N_8521);
nor U8583 (N_8583,N_8490,N_8433);
and U8584 (N_8584,N_8537,N_8469);
xnor U8585 (N_8585,N_8449,N_8442);
and U8586 (N_8586,N_8532,N_8445);
and U8587 (N_8587,N_8529,N_8463);
and U8588 (N_8588,N_8538,N_8429);
or U8589 (N_8589,N_8447,N_8472);
nand U8590 (N_8590,N_8427,N_8497);
and U8591 (N_8591,N_8423,N_8531);
nand U8592 (N_8592,N_8484,N_8507);
nor U8593 (N_8593,N_8416,N_8549);
nand U8594 (N_8594,N_8431,N_8491);
nor U8595 (N_8595,N_8411,N_8525);
nand U8596 (N_8596,N_8452,N_8443);
and U8597 (N_8597,N_8412,N_8400);
and U8598 (N_8598,N_8544,N_8459);
xnor U8599 (N_8599,N_8457,N_8409);
nand U8600 (N_8600,N_8454,N_8536);
nor U8601 (N_8601,N_8480,N_8440);
and U8602 (N_8602,N_8422,N_8470);
and U8603 (N_8603,N_8476,N_8410);
nor U8604 (N_8604,N_8418,N_8478);
and U8605 (N_8605,N_8462,N_8508);
and U8606 (N_8606,N_8488,N_8413);
or U8607 (N_8607,N_8401,N_8434);
nor U8608 (N_8608,N_8475,N_8518);
xnor U8609 (N_8609,N_8473,N_8502);
or U8610 (N_8610,N_8520,N_8534);
xnor U8611 (N_8611,N_8404,N_8455);
nor U8612 (N_8612,N_8516,N_8436);
xor U8613 (N_8613,N_8496,N_8419);
nor U8614 (N_8614,N_8486,N_8514);
or U8615 (N_8615,N_8498,N_8402);
xnor U8616 (N_8616,N_8465,N_8511);
nand U8617 (N_8617,N_8541,N_8481);
or U8618 (N_8618,N_8424,N_8522);
nand U8619 (N_8619,N_8494,N_8450);
or U8620 (N_8620,N_8483,N_8474);
xor U8621 (N_8621,N_8487,N_8493);
or U8622 (N_8622,N_8407,N_8466);
nand U8623 (N_8623,N_8501,N_8453);
and U8624 (N_8624,N_8414,N_8523);
or U8625 (N_8625,N_8444,N_8537);
or U8626 (N_8626,N_8494,N_8466);
xor U8627 (N_8627,N_8525,N_8457);
or U8628 (N_8628,N_8536,N_8417);
and U8629 (N_8629,N_8461,N_8547);
nand U8630 (N_8630,N_8454,N_8482);
xnor U8631 (N_8631,N_8537,N_8407);
and U8632 (N_8632,N_8541,N_8494);
and U8633 (N_8633,N_8493,N_8407);
nor U8634 (N_8634,N_8526,N_8411);
and U8635 (N_8635,N_8529,N_8457);
nand U8636 (N_8636,N_8402,N_8465);
or U8637 (N_8637,N_8444,N_8408);
or U8638 (N_8638,N_8467,N_8443);
nand U8639 (N_8639,N_8466,N_8422);
nor U8640 (N_8640,N_8505,N_8482);
or U8641 (N_8641,N_8522,N_8434);
and U8642 (N_8642,N_8429,N_8437);
xnor U8643 (N_8643,N_8494,N_8476);
nor U8644 (N_8644,N_8548,N_8505);
nand U8645 (N_8645,N_8545,N_8461);
or U8646 (N_8646,N_8521,N_8400);
nand U8647 (N_8647,N_8514,N_8521);
and U8648 (N_8648,N_8434,N_8539);
and U8649 (N_8649,N_8507,N_8506);
xnor U8650 (N_8650,N_8521,N_8449);
and U8651 (N_8651,N_8503,N_8501);
nor U8652 (N_8652,N_8491,N_8495);
xnor U8653 (N_8653,N_8497,N_8545);
nand U8654 (N_8654,N_8460,N_8478);
and U8655 (N_8655,N_8540,N_8499);
xor U8656 (N_8656,N_8426,N_8527);
nor U8657 (N_8657,N_8405,N_8540);
or U8658 (N_8658,N_8512,N_8545);
and U8659 (N_8659,N_8412,N_8487);
xnor U8660 (N_8660,N_8461,N_8502);
or U8661 (N_8661,N_8412,N_8485);
nor U8662 (N_8662,N_8542,N_8502);
nor U8663 (N_8663,N_8415,N_8410);
or U8664 (N_8664,N_8414,N_8497);
nand U8665 (N_8665,N_8492,N_8487);
or U8666 (N_8666,N_8439,N_8467);
nand U8667 (N_8667,N_8492,N_8479);
and U8668 (N_8668,N_8406,N_8445);
and U8669 (N_8669,N_8455,N_8528);
or U8670 (N_8670,N_8496,N_8512);
nand U8671 (N_8671,N_8480,N_8474);
nand U8672 (N_8672,N_8514,N_8470);
nor U8673 (N_8673,N_8511,N_8439);
xor U8674 (N_8674,N_8501,N_8534);
or U8675 (N_8675,N_8425,N_8516);
and U8676 (N_8676,N_8465,N_8522);
xor U8677 (N_8677,N_8542,N_8456);
or U8678 (N_8678,N_8423,N_8517);
or U8679 (N_8679,N_8436,N_8416);
xnor U8680 (N_8680,N_8483,N_8485);
nand U8681 (N_8681,N_8487,N_8489);
nor U8682 (N_8682,N_8513,N_8538);
xor U8683 (N_8683,N_8406,N_8515);
nor U8684 (N_8684,N_8444,N_8538);
and U8685 (N_8685,N_8464,N_8483);
and U8686 (N_8686,N_8541,N_8415);
and U8687 (N_8687,N_8419,N_8454);
nand U8688 (N_8688,N_8446,N_8518);
nor U8689 (N_8689,N_8521,N_8436);
and U8690 (N_8690,N_8531,N_8478);
and U8691 (N_8691,N_8419,N_8526);
and U8692 (N_8692,N_8515,N_8439);
xnor U8693 (N_8693,N_8510,N_8503);
nand U8694 (N_8694,N_8513,N_8441);
xnor U8695 (N_8695,N_8444,N_8406);
nor U8696 (N_8696,N_8530,N_8483);
nor U8697 (N_8697,N_8425,N_8472);
nor U8698 (N_8698,N_8476,N_8431);
nor U8699 (N_8699,N_8438,N_8405);
nor U8700 (N_8700,N_8564,N_8611);
or U8701 (N_8701,N_8565,N_8640);
or U8702 (N_8702,N_8690,N_8686);
xnor U8703 (N_8703,N_8677,N_8578);
nand U8704 (N_8704,N_8567,N_8576);
and U8705 (N_8705,N_8650,N_8596);
nand U8706 (N_8706,N_8617,N_8682);
nor U8707 (N_8707,N_8587,N_8626);
xor U8708 (N_8708,N_8642,N_8689);
and U8709 (N_8709,N_8612,N_8603);
and U8710 (N_8710,N_8594,N_8658);
or U8711 (N_8711,N_8562,N_8697);
xor U8712 (N_8712,N_8621,N_8619);
and U8713 (N_8713,N_8613,N_8601);
nand U8714 (N_8714,N_8692,N_8577);
or U8715 (N_8715,N_8665,N_8571);
and U8716 (N_8716,N_8585,N_8561);
xor U8717 (N_8717,N_8678,N_8673);
xnor U8718 (N_8718,N_8655,N_8608);
xor U8719 (N_8719,N_8555,N_8660);
or U8720 (N_8720,N_8674,N_8659);
xor U8721 (N_8721,N_8639,N_8551);
nand U8722 (N_8722,N_8602,N_8590);
and U8723 (N_8723,N_8647,N_8656);
nand U8724 (N_8724,N_8579,N_8609);
and U8725 (N_8725,N_8627,N_8648);
and U8726 (N_8726,N_8610,N_8651);
or U8727 (N_8727,N_8634,N_8550);
or U8728 (N_8728,N_8570,N_8654);
xor U8729 (N_8729,N_8695,N_8676);
or U8730 (N_8730,N_8574,N_8606);
and U8731 (N_8731,N_8556,N_8691);
and U8732 (N_8732,N_8615,N_8652);
or U8733 (N_8733,N_8566,N_8680);
nor U8734 (N_8734,N_8553,N_8604);
nand U8735 (N_8735,N_8672,N_8688);
and U8736 (N_8736,N_8653,N_8671);
nand U8737 (N_8737,N_8698,N_8662);
nand U8738 (N_8738,N_8595,N_8646);
xor U8739 (N_8739,N_8696,N_8558);
nor U8740 (N_8740,N_8694,N_8591);
nand U8741 (N_8741,N_8581,N_8607);
or U8742 (N_8742,N_8573,N_8623);
and U8743 (N_8743,N_8622,N_8636);
nor U8744 (N_8744,N_8563,N_8679);
nand U8745 (N_8745,N_8586,N_8600);
and U8746 (N_8746,N_8667,N_8669);
or U8747 (N_8747,N_8628,N_8664);
nor U8748 (N_8748,N_8631,N_8569);
xor U8749 (N_8749,N_8630,N_8645);
xor U8750 (N_8750,N_8620,N_8560);
xor U8751 (N_8751,N_8599,N_8598);
nand U8752 (N_8752,N_8635,N_8637);
nor U8753 (N_8753,N_8593,N_8552);
and U8754 (N_8754,N_8681,N_8605);
nor U8755 (N_8755,N_8575,N_8588);
nand U8756 (N_8756,N_8644,N_8618);
nor U8757 (N_8757,N_8670,N_8568);
or U8758 (N_8758,N_8661,N_8693);
and U8759 (N_8759,N_8699,N_8616);
and U8760 (N_8760,N_8559,N_8683);
or U8761 (N_8761,N_8572,N_8632);
nor U8762 (N_8762,N_8580,N_8597);
or U8763 (N_8763,N_8629,N_8554);
nand U8764 (N_8764,N_8641,N_8687);
or U8765 (N_8765,N_8685,N_8666);
xnor U8766 (N_8766,N_8657,N_8649);
or U8767 (N_8767,N_8582,N_8557);
and U8768 (N_8768,N_8643,N_8614);
nand U8769 (N_8769,N_8684,N_8675);
nor U8770 (N_8770,N_8638,N_8633);
nor U8771 (N_8771,N_8592,N_8668);
and U8772 (N_8772,N_8583,N_8589);
or U8773 (N_8773,N_8624,N_8584);
or U8774 (N_8774,N_8625,N_8663);
nand U8775 (N_8775,N_8553,N_8551);
nor U8776 (N_8776,N_8620,N_8696);
nor U8777 (N_8777,N_8613,N_8588);
nor U8778 (N_8778,N_8568,N_8583);
or U8779 (N_8779,N_8629,N_8677);
nand U8780 (N_8780,N_8591,N_8551);
nand U8781 (N_8781,N_8667,N_8593);
xor U8782 (N_8782,N_8568,N_8681);
and U8783 (N_8783,N_8651,N_8563);
nand U8784 (N_8784,N_8647,N_8698);
and U8785 (N_8785,N_8635,N_8631);
nand U8786 (N_8786,N_8560,N_8575);
or U8787 (N_8787,N_8678,N_8563);
and U8788 (N_8788,N_8661,N_8596);
and U8789 (N_8789,N_8670,N_8564);
and U8790 (N_8790,N_8669,N_8597);
nor U8791 (N_8791,N_8584,N_8640);
nand U8792 (N_8792,N_8635,N_8577);
nor U8793 (N_8793,N_8645,N_8608);
nor U8794 (N_8794,N_8698,N_8636);
and U8795 (N_8795,N_8633,N_8579);
nor U8796 (N_8796,N_8691,N_8642);
and U8797 (N_8797,N_8596,N_8696);
nor U8798 (N_8798,N_8626,N_8666);
or U8799 (N_8799,N_8550,N_8651);
nor U8800 (N_8800,N_8566,N_8671);
xnor U8801 (N_8801,N_8665,N_8639);
nand U8802 (N_8802,N_8660,N_8580);
nor U8803 (N_8803,N_8559,N_8554);
nand U8804 (N_8804,N_8558,N_8613);
xnor U8805 (N_8805,N_8592,N_8669);
nand U8806 (N_8806,N_8605,N_8580);
xnor U8807 (N_8807,N_8601,N_8637);
or U8808 (N_8808,N_8602,N_8611);
or U8809 (N_8809,N_8624,N_8574);
and U8810 (N_8810,N_8612,N_8641);
nand U8811 (N_8811,N_8657,N_8675);
nand U8812 (N_8812,N_8612,N_8592);
xor U8813 (N_8813,N_8642,N_8677);
nand U8814 (N_8814,N_8590,N_8671);
or U8815 (N_8815,N_8630,N_8665);
and U8816 (N_8816,N_8653,N_8611);
or U8817 (N_8817,N_8695,N_8584);
nor U8818 (N_8818,N_8595,N_8590);
nand U8819 (N_8819,N_8599,N_8551);
and U8820 (N_8820,N_8558,N_8662);
nand U8821 (N_8821,N_8569,N_8683);
xnor U8822 (N_8822,N_8649,N_8650);
nand U8823 (N_8823,N_8652,N_8572);
or U8824 (N_8824,N_8637,N_8570);
xor U8825 (N_8825,N_8675,N_8609);
nand U8826 (N_8826,N_8665,N_8697);
nand U8827 (N_8827,N_8572,N_8631);
or U8828 (N_8828,N_8556,N_8649);
nor U8829 (N_8829,N_8613,N_8633);
xnor U8830 (N_8830,N_8632,N_8662);
nor U8831 (N_8831,N_8649,N_8567);
and U8832 (N_8832,N_8642,N_8662);
and U8833 (N_8833,N_8625,N_8581);
nand U8834 (N_8834,N_8671,N_8584);
nand U8835 (N_8835,N_8662,N_8692);
nor U8836 (N_8836,N_8602,N_8637);
xor U8837 (N_8837,N_8624,N_8554);
or U8838 (N_8838,N_8570,N_8691);
nand U8839 (N_8839,N_8619,N_8668);
nor U8840 (N_8840,N_8629,N_8560);
nand U8841 (N_8841,N_8643,N_8677);
nor U8842 (N_8842,N_8667,N_8690);
and U8843 (N_8843,N_8611,N_8660);
nand U8844 (N_8844,N_8688,N_8587);
and U8845 (N_8845,N_8654,N_8555);
nor U8846 (N_8846,N_8595,N_8607);
or U8847 (N_8847,N_8597,N_8625);
nor U8848 (N_8848,N_8684,N_8612);
nor U8849 (N_8849,N_8603,N_8575);
nor U8850 (N_8850,N_8730,N_8838);
nand U8851 (N_8851,N_8810,N_8849);
nor U8852 (N_8852,N_8771,N_8705);
nor U8853 (N_8853,N_8827,N_8812);
xnor U8854 (N_8854,N_8804,N_8756);
or U8855 (N_8855,N_8744,N_8752);
and U8856 (N_8856,N_8702,N_8842);
nor U8857 (N_8857,N_8807,N_8836);
or U8858 (N_8858,N_8764,N_8727);
and U8859 (N_8859,N_8700,N_8802);
nor U8860 (N_8860,N_8814,N_8723);
nor U8861 (N_8861,N_8798,N_8704);
nor U8862 (N_8862,N_8825,N_8845);
nand U8863 (N_8863,N_8790,N_8758);
nand U8864 (N_8864,N_8767,N_8772);
nor U8865 (N_8865,N_8708,N_8844);
or U8866 (N_8866,N_8725,N_8711);
and U8867 (N_8867,N_8749,N_8745);
nor U8868 (N_8868,N_8788,N_8706);
nand U8869 (N_8869,N_8713,N_8765);
nor U8870 (N_8870,N_8816,N_8829);
nor U8871 (N_8871,N_8714,N_8722);
and U8872 (N_8872,N_8748,N_8775);
and U8873 (N_8873,N_8835,N_8831);
and U8874 (N_8874,N_8709,N_8746);
nor U8875 (N_8875,N_8824,N_8737);
or U8876 (N_8876,N_8747,N_8782);
and U8877 (N_8877,N_8833,N_8834);
xnor U8878 (N_8878,N_8822,N_8735);
nor U8879 (N_8879,N_8741,N_8846);
nand U8880 (N_8880,N_8712,N_8818);
and U8881 (N_8881,N_8776,N_8793);
or U8882 (N_8882,N_8740,N_8753);
and U8883 (N_8883,N_8720,N_8837);
and U8884 (N_8884,N_8808,N_8809);
or U8885 (N_8885,N_8751,N_8774);
nor U8886 (N_8886,N_8715,N_8732);
or U8887 (N_8887,N_8803,N_8847);
nand U8888 (N_8888,N_8716,N_8784);
nand U8889 (N_8889,N_8743,N_8801);
and U8890 (N_8890,N_8777,N_8779);
nand U8891 (N_8891,N_8785,N_8766);
or U8892 (N_8892,N_8721,N_8768);
and U8893 (N_8893,N_8819,N_8736);
xnor U8894 (N_8894,N_8828,N_8791);
xnor U8895 (N_8895,N_8823,N_8761);
xor U8896 (N_8896,N_8789,N_8750);
or U8897 (N_8897,N_8770,N_8830);
nor U8898 (N_8898,N_8707,N_8759);
xnor U8899 (N_8899,N_8760,N_8719);
xor U8900 (N_8900,N_8799,N_8811);
nor U8901 (N_8901,N_8821,N_8832);
nand U8902 (N_8902,N_8710,N_8800);
or U8903 (N_8903,N_8762,N_8703);
nor U8904 (N_8904,N_8734,N_8733);
xnor U8905 (N_8905,N_8796,N_8820);
nor U8906 (N_8906,N_8739,N_8742);
nor U8907 (N_8907,N_8806,N_8773);
or U8908 (N_8908,N_8792,N_8787);
nor U8909 (N_8909,N_8815,N_8731);
nand U8910 (N_8910,N_8786,N_8755);
nand U8911 (N_8911,N_8839,N_8757);
nand U8912 (N_8912,N_8754,N_8724);
and U8913 (N_8913,N_8728,N_8729);
xor U8914 (N_8914,N_8738,N_8848);
nor U8915 (N_8915,N_8794,N_8726);
and U8916 (N_8916,N_8769,N_8840);
and U8917 (N_8917,N_8843,N_8780);
or U8918 (N_8918,N_8781,N_8813);
xor U8919 (N_8919,N_8805,N_8797);
nand U8920 (N_8920,N_8783,N_8795);
nor U8921 (N_8921,N_8763,N_8826);
or U8922 (N_8922,N_8717,N_8841);
nor U8923 (N_8923,N_8718,N_8778);
or U8924 (N_8924,N_8701,N_8817);
nand U8925 (N_8925,N_8827,N_8710);
and U8926 (N_8926,N_8776,N_8733);
xor U8927 (N_8927,N_8841,N_8835);
or U8928 (N_8928,N_8813,N_8769);
nor U8929 (N_8929,N_8762,N_8714);
nand U8930 (N_8930,N_8763,N_8818);
and U8931 (N_8931,N_8796,N_8803);
xor U8932 (N_8932,N_8791,N_8843);
and U8933 (N_8933,N_8777,N_8795);
or U8934 (N_8934,N_8725,N_8709);
or U8935 (N_8935,N_8793,N_8727);
nor U8936 (N_8936,N_8772,N_8728);
nor U8937 (N_8937,N_8775,N_8783);
or U8938 (N_8938,N_8700,N_8826);
nor U8939 (N_8939,N_8772,N_8721);
nor U8940 (N_8940,N_8768,N_8765);
nand U8941 (N_8941,N_8717,N_8834);
or U8942 (N_8942,N_8779,N_8811);
and U8943 (N_8943,N_8751,N_8789);
xor U8944 (N_8944,N_8736,N_8700);
xnor U8945 (N_8945,N_8779,N_8738);
nor U8946 (N_8946,N_8749,N_8724);
or U8947 (N_8947,N_8783,N_8782);
or U8948 (N_8948,N_8831,N_8740);
or U8949 (N_8949,N_8725,N_8701);
nand U8950 (N_8950,N_8804,N_8838);
or U8951 (N_8951,N_8845,N_8819);
nor U8952 (N_8952,N_8768,N_8844);
nand U8953 (N_8953,N_8787,N_8725);
nand U8954 (N_8954,N_8840,N_8807);
or U8955 (N_8955,N_8795,N_8792);
nor U8956 (N_8956,N_8771,N_8730);
and U8957 (N_8957,N_8764,N_8714);
nand U8958 (N_8958,N_8830,N_8812);
xor U8959 (N_8959,N_8777,N_8743);
or U8960 (N_8960,N_8836,N_8797);
or U8961 (N_8961,N_8744,N_8732);
nand U8962 (N_8962,N_8788,N_8834);
or U8963 (N_8963,N_8722,N_8825);
nand U8964 (N_8964,N_8788,N_8832);
xor U8965 (N_8965,N_8705,N_8817);
nor U8966 (N_8966,N_8733,N_8712);
nand U8967 (N_8967,N_8815,N_8838);
nand U8968 (N_8968,N_8717,N_8833);
nand U8969 (N_8969,N_8824,N_8732);
or U8970 (N_8970,N_8747,N_8718);
or U8971 (N_8971,N_8703,N_8820);
or U8972 (N_8972,N_8845,N_8735);
xor U8973 (N_8973,N_8719,N_8741);
or U8974 (N_8974,N_8819,N_8844);
nor U8975 (N_8975,N_8810,N_8727);
xor U8976 (N_8976,N_8753,N_8796);
and U8977 (N_8977,N_8783,N_8733);
or U8978 (N_8978,N_8767,N_8837);
or U8979 (N_8979,N_8835,N_8708);
or U8980 (N_8980,N_8844,N_8737);
and U8981 (N_8981,N_8828,N_8801);
xnor U8982 (N_8982,N_8732,N_8820);
nor U8983 (N_8983,N_8845,N_8801);
or U8984 (N_8984,N_8744,N_8828);
nand U8985 (N_8985,N_8714,N_8790);
xnor U8986 (N_8986,N_8770,N_8720);
and U8987 (N_8987,N_8800,N_8832);
nand U8988 (N_8988,N_8755,N_8750);
nor U8989 (N_8989,N_8740,N_8764);
or U8990 (N_8990,N_8775,N_8836);
or U8991 (N_8991,N_8786,N_8825);
nand U8992 (N_8992,N_8755,N_8824);
xor U8993 (N_8993,N_8774,N_8787);
and U8994 (N_8994,N_8733,N_8849);
and U8995 (N_8995,N_8807,N_8768);
nand U8996 (N_8996,N_8832,N_8829);
xor U8997 (N_8997,N_8700,N_8749);
and U8998 (N_8998,N_8725,N_8790);
or U8999 (N_8999,N_8786,N_8821);
xor U9000 (N_9000,N_8943,N_8921);
nor U9001 (N_9001,N_8981,N_8990);
and U9002 (N_9002,N_8935,N_8890);
or U9003 (N_9003,N_8888,N_8948);
or U9004 (N_9004,N_8862,N_8891);
nor U9005 (N_9005,N_8936,N_8866);
nor U9006 (N_9006,N_8874,N_8980);
and U9007 (N_9007,N_8932,N_8964);
or U9008 (N_9008,N_8957,N_8907);
and U9009 (N_9009,N_8999,N_8996);
or U9010 (N_9010,N_8850,N_8869);
nor U9011 (N_9011,N_8898,N_8880);
or U9012 (N_9012,N_8962,N_8991);
or U9013 (N_9013,N_8940,N_8927);
and U9014 (N_9014,N_8867,N_8913);
nand U9015 (N_9015,N_8883,N_8917);
nand U9016 (N_9016,N_8858,N_8855);
nor U9017 (N_9017,N_8916,N_8876);
nor U9018 (N_9018,N_8914,N_8961);
and U9019 (N_9019,N_8954,N_8877);
nand U9020 (N_9020,N_8909,N_8983);
or U9021 (N_9021,N_8931,N_8944);
and U9022 (N_9022,N_8924,N_8988);
xor U9023 (N_9023,N_8995,N_8859);
xnor U9024 (N_9024,N_8860,N_8972);
nand U9025 (N_9025,N_8947,N_8969);
or U9026 (N_9026,N_8887,N_8977);
nor U9027 (N_9027,N_8863,N_8946);
and U9028 (N_9028,N_8911,N_8974);
xnor U9029 (N_9029,N_8950,N_8951);
nor U9030 (N_9030,N_8992,N_8852);
and U9031 (N_9031,N_8904,N_8856);
and U9032 (N_9032,N_8989,N_8903);
nand U9033 (N_9033,N_8966,N_8857);
or U9034 (N_9034,N_8854,N_8873);
or U9035 (N_9035,N_8945,N_8870);
xnor U9036 (N_9036,N_8926,N_8879);
nor U9037 (N_9037,N_8949,N_8968);
and U9038 (N_9038,N_8939,N_8918);
and U9039 (N_9039,N_8967,N_8889);
nor U9040 (N_9040,N_8982,N_8997);
xnor U9041 (N_9041,N_8985,N_8919);
or U9042 (N_9042,N_8987,N_8942);
nor U9043 (N_9043,N_8871,N_8915);
nor U9044 (N_9044,N_8979,N_8975);
xnor U9045 (N_9045,N_8893,N_8912);
xnor U9046 (N_9046,N_8959,N_8881);
nand U9047 (N_9047,N_8882,N_8925);
and U9048 (N_9048,N_8872,N_8910);
and U9049 (N_9049,N_8958,N_8973);
and U9050 (N_9050,N_8930,N_8923);
and U9051 (N_9051,N_8993,N_8865);
nor U9052 (N_9052,N_8894,N_8956);
nand U9053 (N_9053,N_8878,N_8984);
nor U9054 (N_9054,N_8895,N_8938);
and U9055 (N_9055,N_8929,N_8971);
or U9056 (N_9056,N_8892,N_8902);
and U9057 (N_9057,N_8970,N_8853);
or U9058 (N_9058,N_8896,N_8937);
nand U9059 (N_9059,N_8861,N_8851);
and U9060 (N_9060,N_8933,N_8886);
and U9061 (N_9061,N_8976,N_8953);
or U9062 (N_9062,N_8900,N_8960);
nor U9063 (N_9063,N_8885,N_8955);
and U9064 (N_9064,N_8994,N_8986);
xnor U9065 (N_9065,N_8899,N_8906);
nand U9066 (N_9066,N_8920,N_8868);
and U9067 (N_9067,N_8998,N_8864);
nor U9068 (N_9068,N_8897,N_8934);
nor U9069 (N_9069,N_8908,N_8952);
nand U9070 (N_9070,N_8905,N_8875);
and U9071 (N_9071,N_8963,N_8941);
xor U9072 (N_9072,N_8884,N_8978);
nor U9073 (N_9073,N_8901,N_8922);
nand U9074 (N_9074,N_8965,N_8928);
or U9075 (N_9075,N_8990,N_8960);
xnor U9076 (N_9076,N_8943,N_8968);
nor U9077 (N_9077,N_8894,N_8964);
xor U9078 (N_9078,N_8987,N_8966);
or U9079 (N_9079,N_8970,N_8916);
and U9080 (N_9080,N_8903,N_8924);
or U9081 (N_9081,N_8863,N_8913);
or U9082 (N_9082,N_8958,N_8988);
and U9083 (N_9083,N_8926,N_8861);
or U9084 (N_9084,N_8905,N_8885);
nand U9085 (N_9085,N_8879,N_8977);
nand U9086 (N_9086,N_8962,N_8993);
and U9087 (N_9087,N_8864,N_8867);
nor U9088 (N_9088,N_8926,N_8988);
nor U9089 (N_9089,N_8888,N_8923);
nor U9090 (N_9090,N_8861,N_8924);
xor U9091 (N_9091,N_8965,N_8865);
nand U9092 (N_9092,N_8986,N_8944);
nand U9093 (N_9093,N_8871,N_8979);
nand U9094 (N_9094,N_8906,N_8932);
nor U9095 (N_9095,N_8890,N_8960);
and U9096 (N_9096,N_8938,N_8901);
nand U9097 (N_9097,N_8909,N_8919);
or U9098 (N_9098,N_8957,N_8940);
nor U9099 (N_9099,N_8900,N_8962);
or U9100 (N_9100,N_8882,N_8881);
nand U9101 (N_9101,N_8959,N_8935);
nor U9102 (N_9102,N_8977,N_8960);
xnor U9103 (N_9103,N_8917,N_8989);
or U9104 (N_9104,N_8981,N_8988);
or U9105 (N_9105,N_8901,N_8918);
nor U9106 (N_9106,N_8980,N_8909);
nand U9107 (N_9107,N_8898,N_8933);
xnor U9108 (N_9108,N_8864,N_8974);
nor U9109 (N_9109,N_8996,N_8926);
xnor U9110 (N_9110,N_8976,N_8925);
or U9111 (N_9111,N_8863,N_8908);
nand U9112 (N_9112,N_8988,N_8884);
nor U9113 (N_9113,N_8927,N_8925);
nor U9114 (N_9114,N_8892,N_8998);
and U9115 (N_9115,N_8974,N_8975);
and U9116 (N_9116,N_8971,N_8914);
xor U9117 (N_9117,N_8889,N_8916);
nand U9118 (N_9118,N_8950,N_8869);
nor U9119 (N_9119,N_8961,N_8863);
xor U9120 (N_9120,N_8960,N_8908);
nand U9121 (N_9121,N_8866,N_8930);
or U9122 (N_9122,N_8858,N_8856);
or U9123 (N_9123,N_8864,N_8947);
or U9124 (N_9124,N_8954,N_8921);
nor U9125 (N_9125,N_8909,N_8967);
nand U9126 (N_9126,N_8945,N_8959);
xor U9127 (N_9127,N_8910,N_8890);
nor U9128 (N_9128,N_8991,N_8918);
and U9129 (N_9129,N_8995,N_8912);
nor U9130 (N_9130,N_8970,N_8978);
or U9131 (N_9131,N_8955,N_8939);
nand U9132 (N_9132,N_8909,N_8917);
nor U9133 (N_9133,N_8904,N_8899);
or U9134 (N_9134,N_8857,N_8952);
xor U9135 (N_9135,N_8997,N_8960);
nand U9136 (N_9136,N_8911,N_8937);
nor U9137 (N_9137,N_8981,N_8935);
and U9138 (N_9138,N_8958,N_8894);
nand U9139 (N_9139,N_8862,N_8910);
or U9140 (N_9140,N_8894,N_8980);
and U9141 (N_9141,N_8933,N_8895);
and U9142 (N_9142,N_8943,N_8905);
nor U9143 (N_9143,N_8902,N_8951);
nand U9144 (N_9144,N_8958,N_8969);
nor U9145 (N_9145,N_8860,N_8887);
xnor U9146 (N_9146,N_8971,N_8879);
nor U9147 (N_9147,N_8882,N_8874);
and U9148 (N_9148,N_8952,N_8855);
and U9149 (N_9149,N_8870,N_8975);
nand U9150 (N_9150,N_9107,N_9132);
xor U9151 (N_9151,N_9018,N_9064);
and U9152 (N_9152,N_9131,N_9135);
and U9153 (N_9153,N_9040,N_9014);
nor U9154 (N_9154,N_9020,N_9036);
xnor U9155 (N_9155,N_9122,N_9016);
and U9156 (N_9156,N_9110,N_9124);
xnor U9157 (N_9157,N_9035,N_9062);
nor U9158 (N_9158,N_9061,N_9010);
xor U9159 (N_9159,N_9069,N_9128);
xor U9160 (N_9160,N_9096,N_9049);
or U9161 (N_9161,N_9113,N_9088);
and U9162 (N_9162,N_9045,N_9024);
xnor U9163 (N_9163,N_9146,N_9022);
nand U9164 (N_9164,N_9111,N_9144);
xor U9165 (N_9165,N_9005,N_9136);
nor U9166 (N_9166,N_9077,N_9087);
nand U9167 (N_9167,N_9063,N_9125);
and U9168 (N_9168,N_9026,N_9009);
and U9169 (N_9169,N_9090,N_9104);
xor U9170 (N_9170,N_9067,N_9118);
nor U9171 (N_9171,N_9085,N_9052);
nand U9172 (N_9172,N_9006,N_9027);
nor U9173 (N_9173,N_9115,N_9031);
nor U9174 (N_9174,N_9127,N_9112);
nand U9175 (N_9175,N_9089,N_9083);
or U9176 (N_9176,N_9034,N_9054);
nand U9177 (N_9177,N_9101,N_9143);
xor U9178 (N_9178,N_9126,N_9117);
xor U9179 (N_9179,N_9106,N_9032);
nor U9180 (N_9180,N_9003,N_9147);
or U9181 (N_9181,N_9070,N_9114);
nor U9182 (N_9182,N_9123,N_9109);
and U9183 (N_9183,N_9091,N_9042);
and U9184 (N_9184,N_9138,N_9055);
nand U9185 (N_9185,N_9097,N_9116);
and U9186 (N_9186,N_9142,N_9100);
nor U9187 (N_9187,N_9102,N_9149);
and U9188 (N_9188,N_9043,N_9001);
xor U9189 (N_9189,N_9044,N_9050);
nand U9190 (N_9190,N_9098,N_9021);
nand U9191 (N_9191,N_9025,N_9121);
xnor U9192 (N_9192,N_9080,N_9059);
nor U9193 (N_9193,N_9141,N_9086);
nor U9194 (N_9194,N_9140,N_9007);
nand U9195 (N_9195,N_9039,N_9015);
or U9196 (N_9196,N_9074,N_9019);
or U9197 (N_9197,N_9011,N_9071);
or U9198 (N_9198,N_9017,N_9139);
and U9199 (N_9199,N_9023,N_9129);
and U9200 (N_9200,N_9066,N_9073);
or U9201 (N_9201,N_9033,N_9004);
nor U9202 (N_9202,N_9145,N_9012);
nor U9203 (N_9203,N_9057,N_9060);
and U9204 (N_9204,N_9108,N_9130);
xor U9205 (N_9205,N_9002,N_9053);
xor U9206 (N_9206,N_9076,N_9148);
or U9207 (N_9207,N_9041,N_9093);
nor U9208 (N_9208,N_9029,N_9133);
nor U9209 (N_9209,N_9008,N_9056);
nor U9210 (N_9210,N_9030,N_9048);
or U9211 (N_9211,N_9047,N_9038);
and U9212 (N_9212,N_9013,N_9105);
xnor U9213 (N_9213,N_9092,N_9134);
or U9214 (N_9214,N_9068,N_9051);
nor U9215 (N_9215,N_9075,N_9103);
nand U9216 (N_9216,N_9079,N_9084);
xor U9217 (N_9217,N_9058,N_9072);
nor U9218 (N_9218,N_9000,N_9037);
nand U9219 (N_9219,N_9095,N_9094);
and U9220 (N_9220,N_9081,N_9028);
or U9221 (N_9221,N_9065,N_9099);
xor U9222 (N_9222,N_9137,N_9120);
nor U9223 (N_9223,N_9046,N_9082);
and U9224 (N_9224,N_9078,N_9119);
nand U9225 (N_9225,N_9137,N_9083);
nor U9226 (N_9226,N_9118,N_9081);
or U9227 (N_9227,N_9071,N_9142);
nor U9228 (N_9228,N_9116,N_9079);
and U9229 (N_9229,N_9053,N_9014);
xnor U9230 (N_9230,N_9070,N_9058);
and U9231 (N_9231,N_9080,N_9136);
nand U9232 (N_9232,N_9044,N_9115);
or U9233 (N_9233,N_9147,N_9118);
xor U9234 (N_9234,N_9094,N_9126);
xnor U9235 (N_9235,N_9038,N_9035);
xor U9236 (N_9236,N_9071,N_9062);
nor U9237 (N_9237,N_9074,N_9060);
nand U9238 (N_9238,N_9012,N_9019);
nor U9239 (N_9239,N_9109,N_9011);
xnor U9240 (N_9240,N_9146,N_9013);
or U9241 (N_9241,N_9034,N_9132);
xor U9242 (N_9242,N_9048,N_9066);
nand U9243 (N_9243,N_9041,N_9141);
nand U9244 (N_9244,N_9064,N_9131);
xnor U9245 (N_9245,N_9108,N_9053);
or U9246 (N_9246,N_9101,N_9123);
nand U9247 (N_9247,N_9043,N_9074);
xor U9248 (N_9248,N_9102,N_9148);
xor U9249 (N_9249,N_9119,N_9005);
or U9250 (N_9250,N_9027,N_9042);
or U9251 (N_9251,N_9012,N_9007);
or U9252 (N_9252,N_9040,N_9069);
and U9253 (N_9253,N_9146,N_9148);
nand U9254 (N_9254,N_9099,N_9042);
xnor U9255 (N_9255,N_9122,N_9116);
or U9256 (N_9256,N_9127,N_9048);
xnor U9257 (N_9257,N_9125,N_9110);
and U9258 (N_9258,N_9059,N_9106);
xnor U9259 (N_9259,N_9102,N_9086);
or U9260 (N_9260,N_9095,N_9009);
and U9261 (N_9261,N_9024,N_9033);
and U9262 (N_9262,N_9096,N_9030);
xnor U9263 (N_9263,N_9027,N_9093);
and U9264 (N_9264,N_9036,N_9105);
or U9265 (N_9265,N_9067,N_9043);
nor U9266 (N_9266,N_9119,N_9127);
and U9267 (N_9267,N_9043,N_9100);
nor U9268 (N_9268,N_9001,N_9098);
and U9269 (N_9269,N_9075,N_9109);
nand U9270 (N_9270,N_9101,N_9098);
or U9271 (N_9271,N_9013,N_9107);
nor U9272 (N_9272,N_9035,N_9121);
and U9273 (N_9273,N_9000,N_9060);
and U9274 (N_9274,N_9003,N_9015);
or U9275 (N_9275,N_9102,N_9138);
or U9276 (N_9276,N_9011,N_9119);
xnor U9277 (N_9277,N_9140,N_9127);
or U9278 (N_9278,N_9091,N_9031);
xor U9279 (N_9279,N_9046,N_9054);
xor U9280 (N_9280,N_9046,N_9067);
or U9281 (N_9281,N_9065,N_9106);
or U9282 (N_9282,N_9015,N_9100);
nor U9283 (N_9283,N_9068,N_9070);
nor U9284 (N_9284,N_9018,N_9035);
and U9285 (N_9285,N_9057,N_9051);
or U9286 (N_9286,N_9036,N_9116);
xor U9287 (N_9287,N_9075,N_9017);
nand U9288 (N_9288,N_9046,N_9131);
or U9289 (N_9289,N_9131,N_9055);
and U9290 (N_9290,N_9139,N_9050);
and U9291 (N_9291,N_9049,N_9056);
or U9292 (N_9292,N_9000,N_9145);
or U9293 (N_9293,N_9146,N_9140);
nand U9294 (N_9294,N_9053,N_9028);
or U9295 (N_9295,N_9117,N_9123);
nor U9296 (N_9296,N_9144,N_9048);
nor U9297 (N_9297,N_9044,N_9055);
or U9298 (N_9298,N_9043,N_9034);
and U9299 (N_9299,N_9001,N_9140);
or U9300 (N_9300,N_9261,N_9181);
or U9301 (N_9301,N_9214,N_9186);
or U9302 (N_9302,N_9272,N_9287);
and U9303 (N_9303,N_9232,N_9288);
nor U9304 (N_9304,N_9218,N_9296);
nor U9305 (N_9305,N_9297,N_9273);
xor U9306 (N_9306,N_9276,N_9215);
xnor U9307 (N_9307,N_9153,N_9211);
nand U9308 (N_9308,N_9244,N_9194);
and U9309 (N_9309,N_9195,N_9221);
or U9310 (N_9310,N_9227,N_9197);
xnor U9311 (N_9311,N_9251,N_9274);
xnor U9312 (N_9312,N_9246,N_9280);
or U9313 (N_9313,N_9269,N_9225);
xor U9314 (N_9314,N_9286,N_9185);
xnor U9315 (N_9315,N_9187,N_9266);
or U9316 (N_9316,N_9263,N_9166);
and U9317 (N_9317,N_9293,N_9226);
xnor U9318 (N_9318,N_9169,N_9292);
or U9319 (N_9319,N_9250,N_9283);
and U9320 (N_9320,N_9154,N_9158);
nor U9321 (N_9321,N_9233,N_9179);
nor U9322 (N_9322,N_9204,N_9174);
or U9323 (N_9323,N_9258,N_9254);
xnor U9324 (N_9324,N_9243,N_9260);
xor U9325 (N_9325,N_9285,N_9278);
and U9326 (N_9326,N_9182,N_9290);
and U9327 (N_9327,N_9188,N_9216);
nor U9328 (N_9328,N_9159,N_9198);
or U9329 (N_9329,N_9294,N_9230);
xor U9330 (N_9330,N_9176,N_9267);
and U9331 (N_9331,N_9291,N_9253);
xnor U9332 (N_9332,N_9231,N_9177);
and U9333 (N_9333,N_9203,N_9279);
nor U9334 (N_9334,N_9259,N_9235);
xnor U9335 (N_9335,N_9155,N_9205);
nand U9336 (N_9336,N_9156,N_9284);
xor U9337 (N_9337,N_9196,N_9173);
or U9338 (N_9338,N_9220,N_9209);
xnor U9339 (N_9339,N_9262,N_9150);
and U9340 (N_9340,N_9228,N_9257);
nor U9341 (N_9341,N_9180,N_9178);
nor U9342 (N_9342,N_9170,N_9167);
nor U9343 (N_9343,N_9298,N_9242);
nand U9344 (N_9344,N_9172,N_9252);
and U9345 (N_9345,N_9152,N_9151);
and U9346 (N_9346,N_9222,N_9245);
nand U9347 (N_9347,N_9282,N_9192);
nand U9348 (N_9348,N_9299,N_9175);
nand U9349 (N_9349,N_9162,N_9201);
xor U9350 (N_9350,N_9240,N_9193);
nor U9351 (N_9351,N_9200,N_9265);
xor U9352 (N_9352,N_9247,N_9256);
and U9353 (N_9353,N_9275,N_9165);
and U9354 (N_9354,N_9236,N_9289);
xor U9355 (N_9355,N_9224,N_9189);
or U9356 (N_9356,N_9191,N_9238);
nand U9357 (N_9357,N_9217,N_9207);
xor U9358 (N_9358,N_9161,N_9164);
or U9359 (N_9359,N_9281,N_9268);
xnor U9360 (N_9360,N_9241,N_9237);
xnor U9361 (N_9361,N_9255,N_9202);
or U9362 (N_9362,N_9248,N_9206);
nand U9363 (N_9363,N_9171,N_9168);
nor U9364 (N_9364,N_9271,N_9277);
or U9365 (N_9365,N_9295,N_9249);
or U9366 (N_9366,N_9210,N_9264);
and U9367 (N_9367,N_9183,N_9223);
nand U9368 (N_9368,N_9160,N_9163);
or U9369 (N_9369,N_9184,N_9234);
and U9370 (N_9370,N_9213,N_9199);
nor U9371 (N_9371,N_9270,N_9229);
or U9372 (N_9372,N_9219,N_9190);
xor U9373 (N_9373,N_9212,N_9208);
nand U9374 (N_9374,N_9239,N_9157);
nand U9375 (N_9375,N_9212,N_9206);
or U9376 (N_9376,N_9201,N_9156);
and U9377 (N_9377,N_9204,N_9279);
and U9378 (N_9378,N_9239,N_9296);
nor U9379 (N_9379,N_9228,N_9247);
xor U9380 (N_9380,N_9279,N_9173);
or U9381 (N_9381,N_9294,N_9234);
or U9382 (N_9382,N_9203,N_9181);
and U9383 (N_9383,N_9165,N_9280);
xnor U9384 (N_9384,N_9285,N_9197);
nor U9385 (N_9385,N_9220,N_9281);
nor U9386 (N_9386,N_9218,N_9267);
nand U9387 (N_9387,N_9158,N_9159);
nor U9388 (N_9388,N_9213,N_9267);
xor U9389 (N_9389,N_9257,N_9229);
xnor U9390 (N_9390,N_9255,N_9236);
or U9391 (N_9391,N_9269,N_9239);
or U9392 (N_9392,N_9227,N_9159);
nor U9393 (N_9393,N_9195,N_9194);
nor U9394 (N_9394,N_9267,N_9221);
and U9395 (N_9395,N_9208,N_9265);
nand U9396 (N_9396,N_9257,N_9279);
and U9397 (N_9397,N_9244,N_9274);
nor U9398 (N_9398,N_9171,N_9236);
or U9399 (N_9399,N_9249,N_9152);
and U9400 (N_9400,N_9226,N_9203);
nand U9401 (N_9401,N_9173,N_9292);
or U9402 (N_9402,N_9288,N_9260);
nand U9403 (N_9403,N_9214,N_9197);
nand U9404 (N_9404,N_9290,N_9297);
xnor U9405 (N_9405,N_9210,N_9253);
nor U9406 (N_9406,N_9244,N_9286);
nor U9407 (N_9407,N_9188,N_9179);
and U9408 (N_9408,N_9217,N_9218);
nand U9409 (N_9409,N_9268,N_9289);
xor U9410 (N_9410,N_9264,N_9175);
nand U9411 (N_9411,N_9261,N_9215);
nand U9412 (N_9412,N_9251,N_9252);
and U9413 (N_9413,N_9291,N_9188);
nor U9414 (N_9414,N_9170,N_9267);
xnor U9415 (N_9415,N_9156,N_9259);
xnor U9416 (N_9416,N_9256,N_9282);
or U9417 (N_9417,N_9267,N_9153);
nand U9418 (N_9418,N_9234,N_9173);
and U9419 (N_9419,N_9227,N_9175);
or U9420 (N_9420,N_9234,N_9263);
and U9421 (N_9421,N_9243,N_9178);
nor U9422 (N_9422,N_9280,N_9167);
and U9423 (N_9423,N_9253,N_9208);
nand U9424 (N_9424,N_9193,N_9203);
nand U9425 (N_9425,N_9189,N_9197);
nor U9426 (N_9426,N_9180,N_9270);
nor U9427 (N_9427,N_9157,N_9296);
or U9428 (N_9428,N_9180,N_9255);
and U9429 (N_9429,N_9208,N_9168);
nor U9430 (N_9430,N_9181,N_9278);
nand U9431 (N_9431,N_9206,N_9168);
and U9432 (N_9432,N_9245,N_9283);
nand U9433 (N_9433,N_9218,N_9223);
nand U9434 (N_9434,N_9280,N_9278);
and U9435 (N_9435,N_9174,N_9227);
and U9436 (N_9436,N_9257,N_9261);
nor U9437 (N_9437,N_9257,N_9218);
nand U9438 (N_9438,N_9245,N_9205);
nand U9439 (N_9439,N_9240,N_9260);
or U9440 (N_9440,N_9174,N_9237);
xnor U9441 (N_9441,N_9197,N_9277);
nor U9442 (N_9442,N_9161,N_9157);
xor U9443 (N_9443,N_9199,N_9282);
xnor U9444 (N_9444,N_9248,N_9179);
xor U9445 (N_9445,N_9180,N_9232);
or U9446 (N_9446,N_9239,N_9171);
nand U9447 (N_9447,N_9153,N_9243);
or U9448 (N_9448,N_9246,N_9228);
xnor U9449 (N_9449,N_9222,N_9157);
or U9450 (N_9450,N_9335,N_9315);
nand U9451 (N_9451,N_9310,N_9365);
nor U9452 (N_9452,N_9373,N_9432);
or U9453 (N_9453,N_9403,N_9436);
nand U9454 (N_9454,N_9402,N_9444);
xor U9455 (N_9455,N_9382,N_9336);
or U9456 (N_9456,N_9333,N_9411);
nor U9457 (N_9457,N_9412,N_9375);
xor U9458 (N_9458,N_9337,N_9326);
and U9459 (N_9459,N_9360,N_9407);
nand U9460 (N_9460,N_9354,N_9313);
nor U9461 (N_9461,N_9370,N_9431);
nand U9462 (N_9462,N_9421,N_9307);
xor U9463 (N_9463,N_9417,N_9390);
nor U9464 (N_9464,N_9344,N_9399);
and U9465 (N_9465,N_9334,N_9329);
xnor U9466 (N_9466,N_9353,N_9338);
nor U9467 (N_9467,N_9440,N_9369);
nand U9468 (N_9468,N_9428,N_9367);
nand U9469 (N_9469,N_9433,N_9318);
or U9470 (N_9470,N_9413,N_9327);
nand U9471 (N_9471,N_9355,N_9312);
and U9472 (N_9472,N_9392,N_9426);
nor U9473 (N_9473,N_9358,N_9332);
nand U9474 (N_9474,N_9396,N_9384);
nand U9475 (N_9475,N_9359,N_9328);
nand U9476 (N_9476,N_9429,N_9374);
nand U9477 (N_9477,N_9347,N_9416);
and U9478 (N_9478,N_9325,N_9348);
nor U9479 (N_9479,N_9303,N_9366);
or U9480 (N_9480,N_9340,N_9309);
or U9481 (N_9481,N_9388,N_9314);
nand U9482 (N_9482,N_9443,N_9415);
nand U9483 (N_9483,N_9425,N_9405);
or U9484 (N_9484,N_9317,N_9350);
xor U9485 (N_9485,N_9400,N_9371);
nand U9486 (N_9486,N_9401,N_9387);
or U9487 (N_9487,N_9352,N_9331);
nand U9488 (N_9488,N_9380,N_9386);
nor U9489 (N_9489,N_9306,N_9302);
nand U9490 (N_9490,N_9414,N_9418);
and U9491 (N_9491,N_9383,N_9364);
xnor U9492 (N_9492,N_9361,N_9409);
and U9493 (N_9493,N_9305,N_9324);
xor U9494 (N_9494,N_9389,N_9385);
and U9495 (N_9495,N_9339,N_9434);
nand U9496 (N_9496,N_9449,N_9322);
xnor U9497 (N_9497,N_9419,N_9441);
or U9498 (N_9498,N_9300,N_9378);
and U9499 (N_9499,N_9437,N_9357);
nand U9500 (N_9500,N_9408,N_9404);
nand U9501 (N_9501,N_9342,N_9356);
or U9502 (N_9502,N_9430,N_9372);
and U9503 (N_9503,N_9406,N_9424);
nor U9504 (N_9504,N_9330,N_9423);
and U9505 (N_9505,N_9345,N_9393);
and U9506 (N_9506,N_9368,N_9397);
nor U9507 (N_9507,N_9420,N_9398);
and U9508 (N_9508,N_9301,N_9442);
nor U9509 (N_9509,N_9377,N_9323);
nand U9510 (N_9510,N_9422,N_9363);
xor U9511 (N_9511,N_9395,N_9343);
xor U9512 (N_9512,N_9351,N_9311);
or U9513 (N_9513,N_9319,N_9427);
nand U9514 (N_9514,N_9445,N_9410);
xor U9515 (N_9515,N_9346,N_9316);
nor U9516 (N_9516,N_9349,N_9362);
nor U9517 (N_9517,N_9376,N_9447);
or U9518 (N_9518,N_9308,N_9446);
nor U9519 (N_9519,N_9438,N_9394);
xor U9520 (N_9520,N_9448,N_9320);
nor U9521 (N_9521,N_9391,N_9321);
nand U9522 (N_9522,N_9379,N_9381);
and U9523 (N_9523,N_9341,N_9435);
or U9524 (N_9524,N_9439,N_9304);
nor U9525 (N_9525,N_9349,N_9425);
and U9526 (N_9526,N_9305,N_9432);
xor U9527 (N_9527,N_9343,N_9446);
or U9528 (N_9528,N_9386,N_9387);
or U9529 (N_9529,N_9393,N_9372);
xnor U9530 (N_9530,N_9331,N_9427);
or U9531 (N_9531,N_9416,N_9403);
or U9532 (N_9532,N_9414,N_9319);
or U9533 (N_9533,N_9314,N_9441);
nand U9534 (N_9534,N_9441,N_9374);
nand U9535 (N_9535,N_9424,N_9340);
and U9536 (N_9536,N_9393,N_9384);
and U9537 (N_9537,N_9322,N_9304);
or U9538 (N_9538,N_9449,N_9431);
or U9539 (N_9539,N_9425,N_9397);
nor U9540 (N_9540,N_9344,N_9438);
xor U9541 (N_9541,N_9436,N_9323);
nor U9542 (N_9542,N_9364,N_9394);
or U9543 (N_9543,N_9364,N_9352);
or U9544 (N_9544,N_9416,N_9399);
and U9545 (N_9545,N_9327,N_9307);
or U9546 (N_9546,N_9322,N_9361);
and U9547 (N_9547,N_9440,N_9421);
nand U9548 (N_9548,N_9337,N_9429);
or U9549 (N_9549,N_9369,N_9433);
xnor U9550 (N_9550,N_9423,N_9377);
nand U9551 (N_9551,N_9328,N_9332);
xor U9552 (N_9552,N_9432,N_9354);
nor U9553 (N_9553,N_9355,N_9357);
xor U9554 (N_9554,N_9429,N_9376);
and U9555 (N_9555,N_9321,N_9417);
nand U9556 (N_9556,N_9395,N_9444);
xor U9557 (N_9557,N_9387,N_9439);
nor U9558 (N_9558,N_9351,N_9305);
or U9559 (N_9559,N_9369,N_9324);
nand U9560 (N_9560,N_9363,N_9369);
and U9561 (N_9561,N_9330,N_9376);
nand U9562 (N_9562,N_9380,N_9425);
and U9563 (N_9563,N_9350,N_9383);
nand U9564 (N_9564,N_9389,N_9318);
and U9565 (N_9565,N_9363,N_9323);
or U9566 (N_9566,N_9373,N_9418);
or U9567 (N_9567,N_9379,N_9327);
xor U9568 (N_9568,N_9342,N_9401);
xor U9569 (N_9569,N_9388,N_9320);
nor U9570 (N_9570,N_9414,N_9416);
xor U9571 (N_9571,N_9305,N_9419);
and U9572 (N_9572,N_9442,N_9422);
nor U9573 (N_9573,N_9363,N_9339);
and U9574 (N_9574,N_9419,N_9324);
nand U9575 (N_9575,N_9394,N_9429);
or U9576 (N_9576,N_9310,N_9382);
xor U9577 (N_9577,N_9359,N_9310);
and U9578 (N_9578,N_9367,N_9438);
xor U9579 (N_9579,N_9345,N_9376);
nand U9580 (N_9580,N_9400,N_9440);
or U9581 (N_9581,N_9403,N_9392);
nor U9582 (N_9582,N_9325,N_9313);
or U9583 (N_9583,N_9360,N_9383);
nand U9584 (N_9584,N_9304,N_9406);
or U9585 (N_9585,N_9427,N_9342);
nand U9586 (N_9586,N_9349,N_9405);
and U9587 (N_9587,N_9321,N_9344);
nand U9588 (N_9588,N_9441,N_9326);
nand U9589 (N_9589,N_9348,N_9364);
nand U9590 (N_9590,N_9418,N_9445);
and U9591 (N_9591,N_9330,N_9439);
nand U9592 (N_9592,N_9328,N_9418);
nor U9593 (N_9593,N_9349,N_9429);
and U9594 (N_9594,N_9422,N_9370);
or U9595 (N_9595,N_9337,N_9315);
nand U9596 (N_9596,N_9432,N_9365);
xor U9597 (N_9597,N_9386,N_9411);
or U9598 (N_9598,N_9336,N_9403);
nor U9599 (N_9599,N_9326,N_9429);
nor U9600 (N_9600,N_9548,N_9469);
or U9601 (N_9601,N_9599,N_9479);
and U9602 (N_9602,N_9543,N_9570);
nand U9603 (N_9603,N_9539,N_9538);
nor U9604 (N_9604,N_9509,N_9510);
or U9605 (N_9605,N_9544,N_9527);
nand U9606 (N_9606,N_9526,N_9493);
nand U9607 (N_9607,N_9551,N_9511);
nor U9608 (N_9608,N_9549,N_9468);
nor U9609 (N_9609,N_9576,N_9457);
nand U9610 (N_9610,N_9503,N_9553);
xor U9611 (N_9611,N_9564,N_9451);
xor U9612 (N_9612,N_9536,N_9452);
and U9613 (N_9613,N_9470,N_9546);
and U9614 (N_9614,N_9524,N_9465);
or U9615 (N_9615,N_9577,N_9569);
and U9616 (N_9616,N_9586,N_9597);
nor U9617 (N_9617,N_9547,N_9573);
nand U9618 (N_9618,N_9562,N_9462);
nand U9619 (N_9619,N_9473,N_9537);
xnor U9620 (N_9620,N_9492,N_9561);
and U9621 (N_9621,N_9578,N_9515);
and U9622 (N_9622,N_9521,N_9455);
nand U9623 (N_9623,N_9522,N_9514);
nor U9624 (N_9624,N_9591,N_9460);
nand U9625 (N_9625,N_9485,N_9518);
and U9626 (N_9626,N_9488,N_9520);
xnor U9627 (N_9627,N_9534,N_9582);
xor U9628 (N_9628,N_9472,N_9519);
nor U9629 (N_9629,N_9594,N_9512);
or U9630 (N_9630,N_9500,N_9454);
or U9631 (N_9631,N_9528,N_9506);
nor U9632 (N_9632,N_9489,N_9587);
nand U9633 (N_9633,N_9496,N_9495);
xnor U9634 (N_9634,N_9450,N_9571);
nor U9635 (N_9635,N_9456,N_9580);
and U9636 (N_9636,N_9552,N_9490);
or U9637 (N_9637,N_9533,N_9574);
and U9638 (N_9638,N_9566,N_9463);
and U9639 (N_9639,N_9458,N_9491);
xnor U9640 (N_9640,N_9557,N_9502);
xnor U9641 (N_9641,N_9486,N_9590);
or U9642 (N_9642,N_9477,N_9461);
xnor U9643 (N_9643,N_9579,N_9555);
or U9644 (N_9644,N_9516,N_9530);
and U9645 (N_9645,N_9504,N_9476);
nand U9646 (N_9646,N_9471,N_9542);
and U9647 (N_9647,N_9563,N_9481);
or U9648 (N_9648,N_9584,N_9467);
xnor U9649 (N_9649,N_9592,N_9459);
xor U9650 (N_9650,N_9596,N_9585);
nand U9651 (N_9651,N_9517,N_9453);
and U9652 (N_9652,N_9475,N_9484);
xnor U9653 (N_9653,N_9501,N_9523);
xor U9654 (N_9654,N_9545,N_9593);
and U9655 (N_9655,N_9529,N_9466);
nor U9656 (N_9656,N_9474,N_9482);
xor U9657 (N_9657,N_9483,N_9541);
and U9658 (N_9658,N_9572,N_9568);
nor U9659 (N_9659,N_9556,N_9559);
nor U9660 (N_9660,N_9565,N_9595);
nand U9661 (N_9661,N_9480,N_9494);
nor U9662 (N_9662,N_9560,N_9567);
and U9663 (N_9663,N_9507,N_9558);
xnor U9664 (N_9664,N_9535,N_9531);
or U9665 (N_9665,N_9540,N_9525);
nand U9666 (N_9666,N_9598,N_9532);
xnor U9667 (N_9667,N_9508,N_9589);
nand U9668 (N_9668,N_9575,N_9513);
xor U9669 (N_9669,N_9498,N_9581);
nand U9670 (N_9670,N_9550,N_9554);
nand U9671 (N_9671,N_9497,N_9505);
nor U9672 (N_9672,N_9499,N_9487);
or U9673 (N_9673,N_9588,N_9478);
nand U9674 (N_9674,N_9464,N_9583);
or U9675 (N_9675,N_9517,N_9460);
and U9676 (N_9676,N_9484,N_9518);
or U9677 (N_9677,N_9523,N_9477);
and U9678 (N_9678,N_9550,N_9574);
nand U9679 (N_9679,N_9491,N_9528);
nand U9680 (N_9680,N_9563,N_9498);
nor U9681 (N_9681,N_9551,N_9507);
nor U9682 (N_9682,N_9457,N_9482);
nand U9683 (N_9683,N_9459,N_9474);
nand U9684 (N_9684,N_9583,N_9570);
nor U9685 (N_9685,N_9480,N_9532);
xnor U9686 (N_9686,N_9555,N_9492);
nor U9687 (N_9687,N_9453,N_9547);
xor U9688 (N_9688,N_9564,N_9509);
nor U9689 (N_9689,N_9489,N_9524);
nand U9690 (N_9690,N_9457,N_9532);
or U9691 (N_9691,N_9579,N_9589);
or U9692 (N_9692,N_9559,N_9497);
nand U9693 (N_9693,N_9530,N_9512);
xor U9694 (N_9694,N_9488,N_9599);
xnor U9695 (N_9695,N_9545,N_9506);
nor U9696 (N_9696,N_9471,N_9528);
xor U9697 (N_9697,N_9466,N_9483);
and U9698 (N_9698,N_9583,N_9589);
nor U9699 (N_9699,N_9533,N_9529);
or U9700 (N_9700,N_9461,N_9582);
nand U9701 (N_9701,N_9592,N_9492);
and U9702 (N_9702,N_9566,N_9489);
xnor U9703 (N_9703,N_9498,N_9476);
and U9704 (N_9704,N_9455,N_9471);
nand U9705 (N_9705,N_9460,N_9504);
and U9706 (N_9706,N_9475,N_9499);
and U9707 (N_9707,N_9500,N_9480);
and U9708 (N_9708,N_9466,N_9587);
xnor U9709 (N_9709,N_9595,N_9566);
xor U9710 (N_9710,N_9536,N_9561);
xnor U9711 (N_9711,N_9565,N_9534);
nand U9712 (N_9712,N_9588,N_9470);
xnor U9713 (N_9713,N_9578,N_9520);
and U9714 (N_9714,N_9565,N_9450);
or U9715 (N_9715,N_9557,N_9559);
or U9716 (N_9716,N_9509,N_9503);
or U9717 (N_9717,N_9513,N_9496);
nand U9718 (N_9718,N_9473,N_9584);
or U9719 (N_9719,N_9597,N_9497);
or U9720 (N_9720,N_9521,N_9531);
or U9721 (N_9721,N_9519,N_9532);
xor U9722 (N_9722,N_9456,N_9528);
and U9723 (N_9723,N_9545,N_9527);
nand U9724 (N_9724,N_9559,N_9532);
nand U9725 (N_9725,N_9577,N_9594);
or U9726 (N_9726,N_9479,N_9500);
nand U9727 (N_9727,N_9517,N_9507);
nor U9728 (N_9728,N_9566,N_9518);
nand U9729 (N_9729,N_9586,N_9547);
nor U9730 (N_9730,N_9463,N_9537);
and U9731 (N_9731,N_9472,N_9511);
and U9732 (N_9732,N_9494,N_9519);
nand U9733 (N_9733,N_9531,N_9477);
and U9734 (N_9734,N_9450,N_9486);
nor U9735 (N_9735,N_9591,N_9579);
xnor U9736 (N_9736,N_9488,N_9469);
and U9737 (N_9737,N_9528,N_9523);
nand U9738 (N_9738,N_9492,N_9513);
and U9739 (N_9739,N_9450,N_9454);
or U9740 (N_9740,N_9470,N_9487);
nor U9741 (N_9741,N_9481,N_9539);
nand U9742 (N_9742,N_9530,N_9563);
or U9743 (N_9743,N_9520,N_9575);
nor U9744 (N_9744,N_9509,N_9457);
or U9745 (N_9745,N_9489,N_9471);
xnor U9746 (N_9746,N_9529,N_9528);
and U9747 (N_9747,N_9488,N_9596);
and U9748 (N_9748,N_9537,N_9465);
xnor U9749 (N_9749,N_9489,N_9500);
or U9750 (N_9750,N_9672,N_9735);
or U9751 (N_9751,N_9699,N_9742);
and U9752 (N_9752,N_9630,N_9631);
and U9753 (N_9753,N_9730,N_9635);
nand U9754 (N_9754,N_9613,N_9729);
or U9755 (N_9755,N_9638,N_9634);
and U9756 (N_9756,N_9636,N_9726);
nor U9757 (N_9757,N_9632,N_9698);
nor U9758 (N_9758,N_9719,N_9717);
nand U9759 (N_9759,N_9656,N_9648);
or U9760 (N_9760,N_9695,N_9629);
nand U9761 (N_9761,N_9737,N_9691);
and U9762 (N_9762,N_9675,N_9627);
and U9763 (N_9763,N_9610,N_9714);
and U9764 (N_9764,N_9707,N_9706);
or U9765 (N_9765,N_9653,N_9600);
or U9766 (N_9766,N_9696,N_9621);
xor U9767 (N_9767,N_9747,N_9659);
nand U9768 (N_9768,N_9743,N_9683);
xnor U9769 (N_9769,N_9687,N_9710);
nor U9770 (N_9770,N_9718,N_9657);
and U9771 (N_9771,N_9739,N_9715);
nand U9772 (N_9772,N_9749,N_9611);
and U9773 (N_9773,N_9741,N_9615);
or U9774 (N_9774,N_9664,N_9700);
or U9775 (N_9775,N_9686,N_9626);
xnor U9776 (N_9776,N_9628,N_9668);
xor U9777 (N_9777,N_9666,N_9603);
nand U9778 (N_9778,N_9693,N_9694);
or U9779 (N_9779,N_9640,N_9658);
xor U9780 (N_9780,N_9723,N_9705);
nor U9781 (N_9781,N_9722,N_9692);
xor U9782 (N_9782,N_9732,N_9676);
nand U9783 (N_9783,N_9601,N_9602);
xor U9784 (N_9784,N_9679,N_9620);
and U9785 (N_9785,N_9607,N_9701);
or U9786 (N_9786,N_9684,N_9625);
nor U9787 (N_9787,N_9738,N_9608);
nor U9788 (N_9788,N_9641,N_9736);
nand U9789 (N_9789,N_9680,N_9617);
nor U9790 (N_9790,N_9609,N_9712);
or U9791 (N_9791,N_9746,N_9661);
xor U9792 (N_9792,N_9639,N_9655);
xor U9793 (N_9793,N_9673,N_9623);
and U9794 (N_9794,N_9650,N_9614);
and U9795 (N_9795,N_9667,N_9713);
xor U9796 (N_9796,N_9697,N_9685);
or U9797 (N_9797,N_9646,N_9678);
and U9798 (N_9798,N_9704,N_9702);
and U9799 (N_9799,N_9711,N_9734);
or U9800 (N_9800,N_9633,N_9637);
nor U9801 (N_9801,N_9671,N_9748);
or U9802 (N_9802,N_9604,N_9674);
xor U9803 (N_9803,N_9689,N_9647);
nor U9804 (N_9804,N_9619,N_9642);
and U9805 (N_9805,N_9720,N_9708);
xor U9806 (N_9806,N_9670,N_9727);
or U9807 (N_9807,N_9643,N_9612);
xor U9808 (N_9808,N_9622,N_9703);
nand U9809 (N_9809,N_9624,N_9662);
or U9810 (N_9810,N_9652,N_9733);
or U9811 (N_9811,N_9682,N_9660);
nand U9812 (N_9812,N_9649,N_9688);
nand U9813 (N_9813,N_9725,N_9690);
or U9814 (N_9814,N_9721,N_9665);
and U9815 (N_9815,N_9618,N_9644);
or U9816 (N_9816,N_9663,N_9724);
or U9817 (N_9817,N_9709,N_9716);
and U9818 (N_9818,N_9740,N_9744);
or U9819 (N_9819,N_9654,N_9677);
nor U9820 (N_9820,N_9645,N_9745);
xnor U9821 (N_9821,N_9606,N_9681);
nor U9822 (N_9822,N_9605,N_9669);
nand U9823 (N_9823,N_9651,N_9616);
and U9824 (N_9824,N_9728,N_9731);
xor U9825 (N_9825,N_9730,N_9743);
nor U9826 (N_9826,N_9731,N_9710);
nand U9827 (N_9827,N_9731,N_9735);
or U9828 (N_9828,N_9610,N_9629);
nor U9829 (N_9829,N_9741,N_9679);
and U9830 (N_9830,N_9646,N_9636);
nor U9831 (N_9831,N_9704,N_9634);
nor U9832 (N_9832,N_9729,N_9611);
nand U9833 (N_9833,N_9677,N_9628);
xnor U9834 (N_9834,N_9723,N_9740);
nor U9835 (N_9835,N_9613,N_9714);
and U9836 (N_9836,N_9743,N_9660);
and U9837 (N_9837,N_9607,N_9649);
nand U9838 (N_9838,N_9614,N_9646);
or U9839 (N_9839,N_9649,N_9728);
or U9840 (N_9840,N_9644,N_9684);
or U9841 (N_9841,N_9648,N_9740);
nand U9842 (N_9842,N_9625,N_9695);
nand U9843 (N_9843,N_9714,N_9656);
xor U9844 (N_9844,N_9722,N_9645);
and U9845 (N_9845,N_9727,N_9737);
and U9846 (N_9846,N_9726,N_9680);
nor U9847 (N_9847,N_9621,N_9705);
nand U9848 (N_9848,N_9663,N_9605);
nand U9849 (N_9849,N_9727,N_9671);
or U9850 (N_9850,N_9606,N_9676);
xnor U9851 (N_9851,N_9690,N_9648);
and U9852 (N_9852,N_9621,N_9626);
xor U9853 (N_9853,N_9695,N_9605);
xor U9854 (N_9854,N_9613,N_9718);
and U9855 (N_9855,N_9699,N_9642);
nand U9856 (N_9856,N_9692,N_9656);
nand U9857 (N_9857,N_9661,N_9632);
and U9858 (N_9858,N_9655,N_9625);
or U9859 (N_9859,N_9651,N_9614);
or U9860 (N_9860,N_9653,N_9657);
nor U9861 (N_9861,N_9717,N_9630);
nor U9862 (N_9862,N_9703,N_9642);
and U9863 (N_9863,N_9640,N_9673);
nor U9864 (N_9864,N_9629,N_9678);
or U9865 (N_9865,N_9638,N_9626);
nand U9866 (N_9866,N_9658,N_9624);
and U9867 (N_9867,N_9722,N_9744);
and U9868 (N_9868,N_9746,N_9686);
nand U9869 (N_9869,N_9724,N_9739);
xnor U9870 (N_9870,N_9708,N_9683);
nor U9871 (N_9871,N_9603,N_9657);
and U9872 (N_9872,N_9714,N_9743);
and U9873 (N_9873,N_9743,N_9705);
nand U9874 (N_9874,N_9712,N_9732);
or U9875 (N_9875,N_9610,N_9726);
nor U9876 (N_9876,N_9649,N_9748);
nand U9877 (N_9877,N_9729,N_9681);
and U9878 (N_9878,N_9743,N_9665);
xnor U9879 (N_9879,N_9707,N_9671);
nor U9880 (N_9880,N_9635,N_9742);
and U9881 (N_9881,N_9727,N_9693);
or U9882 (N_9882,N_9661,N_9703);
or U9883 (N_9883,N_9607,N_9660);
xor U9884 (N_9884,N_9706,N_9671);
or U9885 (N_9885,N_9611,N_9682);
or U9886 (N_9886,N_9742,N_9604);
nor U9887 (N_9887,N_9731,N_9658);
or U9888 (N_9888,N_9719,N_9689);
nand U9889 (N_9889,N_9676,N_9638);
nor U9890 (N_9890,N_9695,N_9661);
or U9891 (N_9891,N_9637,N_9649);
or U9892 (N_9892,N_9642,N_9738);
and U9893 (N_9893,N_9662,N_9656);
or U9894 (N_9894,N_9615,N_9685);
and U9895 (N_9895,N_9617,N_9701);
and U9896 (N_9896,N_9680,N_9744);
or U9897 (N_9897,N_9708,N_9678);
nor U9898 (N_9898,N_9620,N_9609);
nor U9899 (N_9899,N_9606,N_9729);
xnor U9900 (N_9900,N_9812,N_9845);
nand U9901 (N_9901,N_9833,N_9885);
or U9902 (N_9902,N_9781,N_9879);
and U9903 (N_9903,N_9884,N_9895);
xnor U9904 (N_9904,N_9838,N_9855);
and U9905 (N_9905,N_9867,N_9829);
nand U9906 (N_9906,N_9762,N_9805);
nand U9907 (N_9907,N_9843,N_9856);
xor U9908 (N_9908,N_9819,N_9763);
nor U9909 (N_9909,N_9751,N_9825);
xnor U9910 (N_9910,N_9821,N_9849);
nor U9911 (N_9911,N_9863,N_9887);
nor U9912 (N_9912,N_9792,N_9777);
xor U9913 (N_9913,N_9857,N_9854);
and U9914 (N_9914,N_9892,N_9767);
xor U9915 (N_9915,N_9774,N_9824);
nand U9916 (N_9916,N_9820,N_9802);
and U9917 (N_9917,N_9823,N_9890);
and U9918 (N_9918,N_9801,N_9883);
nor U9919 (N_9919,N_9769,N_9759);
xor U9920 (N_9920,N_9765,N_9786);
or U9921 (N_9921,N_9780,N_9779);
xor U9922 (N_9922,N_9758,N_9841);
and U9923 (N_9923,N_9782,N_9789);
xnor U9924 (N_9924,N_9875,N_9868);
nand U9925 (N_9925,N_9797,N_9828);
xnor U9926 (N_9926,N_9853,N_9862);
and U9927 (N_9927,N_9778,N_9871);
and U9928 (N_9928,N_9830,N_9865);
or U9929 (N_9929,N_9831,N_9864);
and U9930 (N_9930,N_9835,N_9897);
nor U9931 (N_9931,N_9761,N_9788);
nor U9932 (N_9932,N_9803,N_9896);
xnor U9933 (N_9933,N_9795,N_9878);
nand U9934 (N_9934,N_9794,N_9882);
nor U9935 (N_9935,N_9790,N_9827);
or U9936 (N_9936,N_9813,N_9760);
nor U9937 (N_9937,N_9754,N_9775);
xnor U9938 (N_9938,N_9872,N_9886);
nand U9939 (N_9939,N_9752,N_9889);
xnor U9940 (N_9940,N_9860,N_9832);
xor U9941 (N_9941,N_9861,N_9806);
xor U9942 (N_9942,N_9753,N_9876);
or U9943 (N_9943,N_9766,N_9898);
or U9944 (N_9944,N_9866,N_9816);
and U9945 (N_9945,N_9750,N_9770);
xnor U9946 (N_9946,N_9764,N_9783);
xnor U9947 (N_9947,N_9815,N_9850);
and U9948 (N_9948,N_9877,N_9888);
nand U9949 (N_9949,N_9847,N_9757);
or U9950 (N_9950,N_9811,N_9834);
nand U9951 (N_9951,N_9787,N_9893);
or U9952 (N_9952,N_9796,N_9771);
and U9953 (N_9953,N_9818,N_9848);
xor U9954 (N_9954,N_9839,N_9894);
nor U9955 (N_9955,N_9755,N_9814);
and U9956 (N_9956,N_9809,N_9899);
or U9957 (N_9957,N_9784,N_9881);
nor U9958 (N_9958,N_9768,N_9846);
or U9959 (N_9959,N_9869,N_9817);
nand U9960 (N_9960,N_9793,N_9800);
xor U9961 (N_9961,N_9756,N_9858);
xor U9962 (N_9962,N_9891,N_9772);
and U9963 (N_9963,N_9810,N_9844);
or U9964 (N_9964,N_9799,N_9851);
or U9965 (N_9965,N_9837,N_9859);
nor U9966 (N_9966,N_9791,N_9773);
or U9967 (N_9967,N_9798,N_9874);
or U9968 (N_9968,N_9842,N_9836);
nor U9969 (N_9969,N_9870,N_9826);
and U9970 (N_9970,N_9873,N_9808);
nor U9971 (N_9971,N_9776,N_9822);
nor U9972 (N_9972,N_9852,N_9807);
xor U9973 (N_9973,N_9804,N_9840);
or U9974 (N_9974,N_9785,N_9880);
xor U9975 (N_9975,N_9823,N_9792);
nand U9976 (N_9976,N_9812,N_9884);
nand U9977 (N_9977,N_9831,N_9776);
xnor U9978 (N_9978,N_9772,N_9859);
nand U9979 (N_9979,N_9884,N_9869);
nor U9980 (N_9980,N_9854,N_9831);
nor U9981 (N_9981,N_9755,N_9883);
xnor U9982 (N_9982,N_9756,N_9816);
or U9983 (N_9983,N_9829,N_9853);
nand U9984 (N_9984,N_9846,N_9847);
nor U9985 (N_9985,N_9785,N_9754);
and U9986 (N_9986,N_9816,N_9832);
nor U9987 (N_9987,N_9846,N_9834);
and U9988 (N_9988,N_9826,N_9868);
nand U9989 (N_9989,N_9759,N_9840);
and U9990 (N_9990,N_9847,N_9889);
xnor U9991 (N_9991,N_9842,N_9789);
nor U9992 (N_9992,N_9786,N_9791);
or U9993 (N_9993,N_9806,N_9811);
nand U9994 (N_9994,N_9899,N_9850);
or U9995 (N_9995,N_9896,N_9793);
or U9996 (N_9996,N_9772,N_9895);
and U9997 (N_9997,N_9806,N_9761);
and U9998 (N_9998,N_9841,N_9776);
nor U9999 (N_9999,N_9770,N_9857);
nand U10000 (N_10000,N_9800,N_9788);
nand U10001 (N_10001,N_9850,N_9792);
or U10002 (N_10002,N_9884,N_9867);
and U10003 (N_10003,N_9836,N_9862);
xnor U10004 (N_10004,N_9807,N_9775);
nand U10005 (N_10005,N_9798,N_9789);
xor U10006 (N_10006,N_9895,N_9764);
xor U10007 (N_10007,N_9831,N_9791);
nor U10008 (N_10008,N_9790,N_9821);
or U10009 (N_10009,N_9895,N_9785);
xnor U10010 (N_10010,N_9899,N_9812);
or U10011 (N_10011,N_9770,N_9827);
nand U10012 (N_10012,N_9882,N_9849);
or U10013 (N_10013,N_9881,N_9864);
xnor U10014 (N_10014,N_9795,N_9851);
xor U10015 (N_10015,N_9822,N_9759);
xnor U10016 (N_10016,N_9802,N_9835);
or U10017 (N_10017,N_9891,N_9842);
or U10018 (N_10018,N_9863,N_9826);
nor U10019 (N_10019,N_9769,N_9792);
nor U10020 (N_10020,N_9795,N_9875);
xnor U10021 (N_10021,N_9835,N_9786);
and U10022 (N_10022,N_9804,N_9886);
nor U10023 (N_10023,N_9822,N_9857);
and U10024 (N_10024,N_9877,N_9854);
xor U10025 (N_10025,N_9786,N_9872);
and U10026 (N_10026,N_9804,N_9761);
nor U10027 (N_10027,N_9834,N_9810);
or U10028 (N_10028,N_9838,N_9841);
and U10029 (N_10029,N_9864,N_9859);
xor U10030 (N_10030,N_9851,N_9885);
nand U10031 (N_10031,N_9840,N_9833);
or U10032 (N_10032,N_9860,N_9772);
nand U10033 (N_10033,N_9773,N_9774);
xnor U10034 (N_10034,N_9880,N_9767);
or U10035 (N_10035,N_9858,N_9772);
nand U10036 (N_10036,N_9796,N_9875);
xnor U10037 (N_10037,N_9892,N_9782);
xor U10038 (N_10038,N_9758,N_9891);
nor U10039 (N_10039,N_9783,N_9779);
xor U10040 (N_10040,N_9794,N_9849);
and U10041 (N_10041,N_9892,N_9791);
and U10042 (N_10042,N_9819,N_9801);
nand U10043 (N_10043,N_9845,N_9805);
and U10044 (N_10044,N_9818,N_9816);
or U10045 (N_10045,N_9869,N_9812);
and U10046 (N_10046,N_9879,N_9813);
xor U10047 (N_10047,N_9860,N_9843);
and U10048 (N_10048,N_9877,N_9791);
and U10049 (N_10049,N_9896,N_9792);
or U10050 (N_10050,N_10030,N_9935);
nand U10051 (N_10051,N_9990,N_10014);
nor U10052 (N_10052,N_10021,N_10008);
and U10053 (N_10053,N_9903,N_9987);
or U10054 (N_10054,N_9908,N_9924);
or U10055 (N_10055,N_9926,N_9929);
or U10056 (N_10056,N_9953,N_9976);
or U10057 (N_10057,N_9945,N_10039);
xor U10058 (N_10058,N_9961,N_9927);
nor U10059 (N_10059,N_9925,N_9918);
xnor U10060 (N_10060,N_9993,N_9921);
xnor U10061 (N_10061,N_9956,N_9943);
nor U10062 (N_10062,N_9910,N_9932);
xnor U10063 (N_10063,N_9934,N_9930);
xnor U10064 (N_10064,N_9917,N_9947);
xor U10065 (N_10065,N_10006,N_9994);
xor U10066 (N_10066,N_9951,N_10032);
or U10067 (N_10067,N_9902,N_10034);
and U10068 (N_10068,N_9966,N_9946);
nor U10069 (N_10069,N_9957,N_10000);
nor U10070 (N_10070,N_9998,N_10040);
nor U10071 (N_10071,N_10047,N_10049);
or U10072 (N_10072,N_10041,N_9968);
nor U10073 (N_10073,N_10016,N_10042);
nor U10074 (N_10074,N_9933,N_9915);
xor U10075 (N_10075,N_9937,N_9905);
nor U10076 (N_10076,N_9965,N_9954);
nand U10077 (N_10077,N_9995,N_9955);
nor U10078 (N_10078,N_10027,N_10044);
xnor U10079 (N_10079,N_9942,N_10043);
nor U10080 (N_10080,N_9950,N_9969);
and U10081 (N_10081,N_10009,N_10028);
nor U10082 (N_10082,N_9941,N_9988);
nor U10083 (N_10083,N_9971,N_9958);
xor U10084 (N_10084,N_9973,N_9975);
and U10085 (N_10085,N_9967,N_10025);
or U10086 (N_10086,N_10003,N_9984);
xnor U10087 (N_10087,N_10024,N_9919);
nor U10088 (N_10088,N_9949,N_9986);
nand U10089 (N_10089,N_9922,N_10010);
or U10090 (N_10090,N_10022,N_9979);
nand U10091 (N_10091,N_9900,N_9940);
nor U10092 (N_10092,N_9991,N_9997);
nand U10093 (N_10093,N_9904,N_9952);
nand U10094 (N_10094,N_9980,N_10011);
nand U10095 (N_10095,N_10005,N_9906);
nand U10096 (N_10096,N_10012,N_9963);
nor U10097 (N_10097,N_9977,N_9939);
nor U10098 (N_10098,N_10046,N_10007);
and U10099 (N_10099,N_9985,N_9923);
nand U10100 (N_10100,N_10004,N_9992);
or U10101 (N_10101,N_10045,N_10015);
xor U10102 (N_10102,N_10013,N_10037);
or U10103 (N_10103,N_9972,N_10036);
nand U10104 (N_10104,N_9989,N_9901);
nor U10105 (N_10105,N_10026,N_10029);
or U10106 (N_10106,N_10035,N_9983);
and U10107 (N_10107,N_9978,N_9970);
nor U10108 (N_10108,N_10018,N_9909);
nor U10109 (N_10109,N_9907,N_9913);
xnor U10110 (N_10110,N_9938,N_9960);
nand U10111 (N_10111,N_9912,N_9936);
nor U10112 (N_10112,N_9914,N_9999);
xnor U10113 (N_10113,N_9964,N_9916);
nor U10114 (N_10114,N_9931,N_10031);
nand U10115 (N_10115,N_10023,N_9944);
xor U10116 (N_10116,N_10038,N_10001);
xor U10117 (N_10117,N_9920,N_10002);
and U10118 (N_10118,N_10048,N_9959);
nand U10119 (N_10119,N_10019,N_10020);
nand U10120 (N_10120,N_9911,N_10033);
xnor U10121 (N_10121,N_9996,N_10017);
and U10122 (N_10122,N_9981,N_9948);
and U10123 (N_10123,N_9928,N_9974);
nand U10124 (N_10124,N_9962,N_9982);
nor U10125 (N_10125,N_9903,N_10042);
nand U10126 (N_10126,N_10014,N_9985);
or U10127 (N_10127,N_9970,N_10047);
and U10128 (N_10128,N_10025,N_10042);
xor U10129 (N_10129,N_9986,N_9914);
nand U10130 (N_10130,N_9919,N_10000);
or U10131 (N_10131,N_9919,N_10028);
or U10132 (N_10132,N_10048,N_9940);
xor U10133 (N_10133,N_10034,N_9905);
or U10134 (N_10134,N_9910,N_10033);
or U10135 (N_10135,N_9915,N_10032);
and U10136 (N_10136,N_9935,N_10034);
or U10137 (N_10137,N_9923,N_9928);
nor U10138 (N_10138,N_9914,N_10010);
xnor U10139 (N_10139,N_9984,N_9962);
or U10140 (N_10140,N_9967,N_9939);
nand U10141 (N_10141,N_9973,N_10044);
and U10142 (N_10142,N_9941,N_9922);
xor U10143 (N_10143,N_9938,N_10007);
and U10144 (N_10144,N_9955,N_9963);
nor U10145 (N_10145,N_10022,N_10031);
and U10146 (N_10146,N_10033,N_9949);
nand U10147 (N_10147,N_9984,N_9974);
or U10148 (N_10148,N_9946,N_10013);
xor U10149 (N_10149,N_9997,N_10041);
and U10150 (N_10150,N_10010,N_9971);
xor U10151 (N_10151,N_9964,N_9972);
nand U10152 (N_10152,N_9993,N_10006);
or U10153 (N_10153,N_9974,N_9952);
nor U10154 (N_10154,N_9996,N_10033);
xnor U10155 (N_10155,N_9926,N_9990);
xnor U10156 (N_10156,N_9937,N_10009);
nor U10157 (N_10157,N_9935,N_9928);
and U10158 (N_10158,N_9935,N_10011);
and U10159 (N_10159,N_10002,N_9942);
or U10160 (N_10160,N_10018,N_10045);
or U10161 (N_10161,N_10022,N_10024);
nand U10162 (N_10162,N_10016,N_10001);
nand U10163 (N_10163,N_10017,N_9909);
xor U10164 (N_10164,N_9925,N_9938);
nor U10165 (N_10165,N_9918,N_9912);
or U10166 (N_10166,N_10044,N_9919);
or U10167 (N_10167,N_10048,N_9963);
nand U10168 (N_10168,N_10006,N_9990);
xnor U10169 (N_10169,N_9910,N_10039);
xnor U10170 (N_10170,N_9912,N_9957);
nand U10171 (N_10171,N_9998,N_10008);
xor U10172 (N_10172,N_10000,N_9956);
nor U10173 (N_10173,N_9954,N_9976);
and U10174 (N_10174,N_9931,N_9908);
or U10175 (N_10175,N_9949,N_9958);
xnor U10176 (N_10176,N_10019,N_10042);
nor U10177 (N_10177,N_9974,N_10010);
or U10178 (N_10178,N_10026,N_10037);
and U10179 (N_10179,N_9907,N_10019);
or U10180 (N_10180,N_9941,N_9987);
nand U10181 (N_10181,N_9932,N_9961);
and U10182 (N_10182,N_10030,N_9911);
or U10183 (N_10183,N_9903,N_10012);
nor U10184 (N_10184,N_10002,N_9993);
nand U10185 (N_10185,N_9979,N_9996);
and U10186 (N_10186,N_9978,N_9975);
xnor U10187 (N_10187,N_10027,N_9998);
xor U10188 (N_10188,N_10034,N_10025);
nor U10189 (N_10189,N_9901,N_9927);
nand U10190 (N_10190,N_9902,N_10042);
nand U10191 (N_10191,N_9915,N_10046);
xor U10192 (N_10192,N_10044,N_9904);
or U10193 (N_10193,N_9942,N_9902);
xnor U10194 (N_10194,N_9992,N_9956);
xnor U10195 (N_10195,N_9905,N_9936);
or U10196 (N_10196,N_9914,N_9908);
or U10197 (N_10197,N_9917,N_9912);
nor U10198 (N_10198,N_9965,N_10004);
nand U10199 (N_10199,N_10003,N_9978);
nor U10200 (N_10200,N_10096,N_10113);
nor U10201 (N_10201,N_10150,N_10078);
nor U10202 (N_10202,N_10126,N_10071);
or U10203 (N_10203,N_10132,N_10120);
nor U10204 (N_10204,N_10198,N_10061);
or U10205 (N_10205,N_10172,N_10185);
or U10206 (N_10206,N_10176,N_10140);
nor U10207 (N_10207,N_10190,N_10154);
or U10208 (N_10208,N_10161,N_10170);
xor U10209 (N_10209,N_10106,N_10117);
nor U10210 (N_10210,N_10089,N_10092);
or U10211 (N_10211,N_10111,N_10168);
nor U10212 (N_10212,N_10125,N_10058);
and U10213 (N_10213,N_10116,N_10067);
or U10214 (N_10214,N_10173,N_10133);
or U10215 (N_10215,N_10156,N_10073);
or U10216 (N_10216,N_10129,N_10072);
nor U10217 (N_10217,N_10165,N_10135);
and U10218 (N_10218,N_10199,N_10177);
or U10219 (N_10219,N_10068,N_10075);
xnor U10220 (N_10220,N_10142,N_10145);
or U10221 (N_10221,N_10184,N_10090);
or U10222 (N_10222,N_10196,N_10088);
nand U10223 (N_10223,N_10137,N_10167);
nor U10224 (N_10224,N_10059,N_10085);
nand U10225 (N_10225,N_10153,N_10188);
nand U10226 (N_10226,N_10063,N_10086);
or U10227 (N_10227,N_10077,N_10087);
or U10228 (N_10228,N_10183,N_10157);
or U10229 (N_10229,N_10069,N_10093);
xor U10230 (N_10230,N_10119,N_10064);
or U10231 (N_10231,N_10104,N_10094);
or U10232 (N_10232,N_10155,N_10103);
xnor U10233 (N_10233,N_10151,N_10100);
nor U10234 (N_10234,N_10179,N_10128);
or U10235 (N_10235,N_10175,N_10056);
xnor U10236 (N_10236,N_10197,N_10118);
and U10237 (N_10237,N_10107,N_10180);
nor U10238 (N_10238,N_10174,N_10143);
nor U10239 (N_10239,N_10066,N_10162);
xnor U10240 (N_10240,N_10194,N_10102);
xnor U10241 (N_10241,N_10055,N_10191);
nor U10242 (N_10242,N_10159,N_10079);
or U10243 (N_10243,N_10152,N_10122);
or U10244 (N_10244,N_10192,N_10193);
nand U10245 (N_10245,N_10082,N_10108);
nor U10246 (N_10246,N_10105,N_10115);
and U10247 (N_10247,N_10138,N_10169);
xor U10248 (N_10248,N_10181,N_10139);
nor U10249 (N_10249,N_10171,N_10123);
and U10250 (N_10250,N_10127,N_10062);
or U10251 (N_10251,N_10051,N_10149);
xor U10252 (N_10252,N_10148,N_10109);
xnor U10253 (N_10253,N_10164,N_10130);
xnor U10254 (N_10254,N_10160,N_10187);
or U10255 (N_10255,N_10084,N_10101);
and U10256 (N_10256,N_10141,N_10186);
xnor U10257 (N_10257,N_10124,N_10114);
nor U10258 (N_10258,N_10095,N_10134);
xor U10259 (N_10259,N_10091,N_10131);
nand U10260 (N_10260,N_10112,N_10182);
nor U10261 (N_10261,N_10110,N_10121);
nand U10262 (N_10262,N_10050,N_10195);
xnor U10263 (N_10263,N_10060,N_10070);
nand U10264 (N_10264,N_10054,N_10147);
or U10265 (N_10265,N_10144,N_10163);
nand U10266 (N_10266,N_10081,N_10189);
nand U10267 (N_10267,N_10052,N_10097);
or U10268 (N_10268,N_10158,N_10076);
xnor U10269 (N_10269,N_10057,N_10074);
nor U10270 (N_10270,N_10099,N_10098);
nand U10271 (N_10271,N_10136,N_10178);
nand U10272 (N_10272,N_10146,N_10080);
and U10273 (N_10273,N_10083,N_10166);
xor U10274 (N_10274,N_10065,N_10053);
or U10275 (N_10275,N_10116,N_10197);
xor U10276 (N_10276,N_10191,N_10117);
xor U10277 (N_10277,N_10090,N_10067);
or U10278 (N_10278,N_10108,N_10064);
or U10279 (N_10279,N_10129,N_10156);
and U10280 (N_10280,N_10149,N_10110);
or U10281 (N_10281,N_10133,N_10091);
nand U10282 (N_10282,N_10196,N_10062);
or U10283 (N_10283,N_10156,N_10095);
or U10284 (N_10284,N_10183,N_10085);
and U10285 (N_10285,N_10111,N_10079);
nand U10286 (N_10286,N_10095,N_10151);
xnor U10287 (N_10287,N_10196,N_10054);
xor U10288 (N_10288,N_10169,N_10199);
nand U10289 (N_10289,N_10082,N_10116);
nand U10290 (N_10290,N_10153,N_10082);
nor U10291 (N_10291,N_10186,N_10158);
or U10292 (N_10292,N_10082,N_10181);
and U10293 (N_10293,N_10147,N_10191);
and U10294 (N_10294,N_10123,N_10067);
xor U10295 (N_10295,N_10191,N_10150);
or U10296 (N_10296,N_10083,N_10050);
or U10297 (N_10297,N_10139,N_10126);
xor U10298 (N_10298,N_10072,N_10177);
nor U10299 (N_10299,N_10156,N_10163);
nand U10300 (N_10300,N_10179,N_10078);
nand U10301 (N_10301,N_10147,N_10101);
nand U10302 (N_10302,N_10079,N_10156);
nand U10303 (N_10303,N_10142,N_10094);
nand U10304 (N_10304,N_10191,N_10151);
nor U10305 (N_10305,N_10095,N_10198);
and U10306 (N_10306,N_10145,N_10139);
nor U10307 (N_10307,N_10168,N_10153);
or U10308 (N_10308,N_10069,N_10086);
or U10309 (N_10309,N_10125,N_10054);
or U10310 (N_10310,N_10125,N_10145);
or U10311 (N_10311,N_10144,N_10116);
or U10312 (N_10312,N_10057,N_10188);
or U10313 (N_10313,N_10115,N_10085);
nor U10314 (N_10314,N_10124,N_10107);
or U10315 (N_10315,N_10167,N_10055);
or U10316 (N_10316,N_10091,N_10127);
xnor U10317 (N_10317,N_10153,N_10161);
xor U10318 (N_10318,N_10147,N_10128);
nor U10319 (N_10319,N_10191,N_10190);
and U10320 (N_10320,N_10053,N_10134);
xnor U10321 (N_10321,N_10093,N_10164);
nand U10322 (N_10322,N_10122,N_10084);
xor U10323 (N_10323,N_10172,N_10053);
or U10324 (N_10324,N_10108,N_10179);
xnor U10325 (N_10325,N_10063,N_10142);
nand U10326 (N_10326,N_10077,N_10185);
and U10327 (N_10327,N_10087,N_10122);
nor U10328 (N_10328,N_10064,N_10126);
nor U10329 (N_10329,N_10197,N_10195);
nand U10330 (N_10330,N_10113,N_10154);
nor U10331 (N_10331,N_10164,N_10143);
nor U10332 (N_10332,N_10192,N_10075);
nor U10333 (N_10333,N_10087,N_10107);
and U10334 (N_10334,N_10073,N_10149);
or U10335 (N_10335,N_10082,N_10145);
xnor U10336 (N_10336,N_10110,N_10143);
or U10337 (N_10337,N_10131,N_10098);
nand U10338 (N_10338,N_10094,N_10097);
xnor U10339 (N_10339,N_10169,N_10088);
xnor U10340 (N_10340,N_10180,N_10176);
nand U10341 (N_10341,N_10134,N_10083);
nand U10342 (N_10342,N_10068,N_10127);
nor U10343 (N_10343,N_10106,N_10077);
and U10344 (N_10344,N_10091,N_10056);
nand U10345 (N_10345,N_10066,N_10074);
and U10346 (N_10346,N_10144,N_10189);
xor U10347 (N_10347,N_10068,N_10099);
xnor U10348 (N_10348,N_10126,N_10193);
and U10349 (N_10349,N_10142,N_10089);
nand U10350 (N_10350,N_10215,N_10234);
xor U10351 (N_10351,N_10342,N_10317);
and U10352 (N_10352,N_10264,N_10248);
and U10353 (N_10353,N_10328,N_10263);
nor U10354 (N_10354,N_10226,N_10330);
and U10355 (N_10355,N_10296,N_10216);
or U10356 (N_10356,N_10257,N_10243);
nand U10357 (N_10357,N_10282,N_10224);
nand U10358 (N_10358,N_10325,N_10249);
nand U10359 (N_10359,N_10256,N_10314);
xor U10360 (N_10360,N_10343,N_10303);
xnor U10361 (N_10361,N_10219,N_10336);
and U10362 (N_10362,N_10280,N_10308);
and U10363 (N_10363,N_10202,N_10320);
xnor U10364 (N_10364,N_10220,N_10289);
and U10365 (N_10365,N_10299,N_10246);
xnor U10366 (N_10366,N_10260,N_10205);
and U10367 (N_10367,N_10225,N_10337);
nor U10368 (N_10368,N_10209,N_10231);
nand U10369 (N_10369,N_10228,N_10208);
xnor U10370 (N_10370,N_10276,N_10236);
and U10371 (N_10371,N_10214,N_10211);
nor U10372 (N_10372,N_10212,N_10252);
and U10373 (N_10373,N_10262,N_10223);
xnor U10374 (N_10374,N_10344,N_10233);
and U10375 (N_10375,N_10324,N_10327);
nand U10376 (N_10376,N_10261,N_10270);
nand U10377 (N_10377,N_10309,N_10242);
nand U10378 (N_10378,N_10339,N_10316);
or U10379 (N_10379,N_10245,N_10307);
and U10380 (N_10380,N_10298,N_10302);
and U10381 (N_10381,N_10283,N_10297);
nor U10382 (N_10382,N_10281,N_10285);
or U10383 (N_10383,N_10258,N_10341);
nand U10384 (N_10384,N_10275,N_10291);
nand U10385 (N_10385,N_10311,N_10251);
xor U10386 (N_10386,N_10268,N_10213);
and U10387 (N_10387,N_10259,N_10334);
and U10388 (N_10388,N_10250,N_10207);
nand U10389 (N_10389,N_10203,N_10267);
and U10390 (N_10390,N_10321,N_10210);
nor U10391 (N_10391,N_10201,N_10313);
nand U10392 (N_10392,N_10218,N_10227);
xor U10393 (N_10393,N_10333,N_10312);
xor U10394 (N_10394,N_10235,N_10345);
nor U10395 (N_10395,N_10331,N_10255);
or U10396 (N_10396,N_10329,N_10284);
xnor U10397 (N_10397,N_10304,N_10335);
and U10398 (N_10398,N_10274,N_10319);
and U10399 (N_10399,N_10318,N_10244);
nand U10400 (N_10400,N_10293,N_10266);
or U10401 (N_10401,N_10278,N_10230);
or U10402 (N_10402,N_10279,N_10340);
nand U10403 (N_10403,N_10206,N_10254);
xnor U10404 (N_10404,N_10277,N_10315);
nor U10405 (N_10405,N_10238,N_10290);
nor U10406 (N_10406,N_10295,N_10301);
nor U10407 (N_10407,N_10204,N_10326);
nand U10408 (N_10408,N_10232,N_10286);
nand U10409 (N_10409,N_10253,N_10272);
xor U10410 (N_10410,N_10287,N_10222);
xor U10411 (N_10411,N_10221,N_10237);
nor U10412 (N_10412,N_10322,N_10240);
nor U10413 (N_10413,N_10348,N_10239);
or U10414 (N_10414,N_10247,N_10338);
or U10415 (N_10415,N_10305,N_10265);
nand U10416 (N_10416,N_10349,N_10271);
or U10417 (N_10417,N_10200,N_10294);
xor U10418 (N_10418,N_10229,N_10347);
or U10419 (N_10419,N_10306,N_10288);
nand U10420 (N_10420,N_10292,N_10346);
xor U10421 (N_10421,N_10323,N_10217);
xor U10422 (N_10422,N_10332,N_10300);
nand U10423 (N_10423,N_10310,N_10273);
nor U10424 (N_10424,N_10241,N_10269);
nor U10425 (N_10425,N_10273,N_10319);
nor U10426 (N_10426,N_10291,N_10266);
nor U10427 (N_10427,N_10306,N_10326);
nand U10428 (N_10428,N_10261,N_10324);
xor U10429 (N_10429,N_10229,N_10302);
or U10430 (N_10430,N_10293,N_10209);
nor U10431 (N_10431,N_10287,N_10225);
xor U10432 (N_10432,N_10259,N_10247);
nand U10433 (N_10433,N_10203,N_10318);
nand U10434 (N_10434,N_10262,N_10299);
xnor U10435 (N_10435,N_10319,N_10336);
and U10436 (N_10436,N_10336,N_10321);
and U10437 (N_10437,N_10282,N_10327);
xnor U10438 (N_10438,N_10317,N_10280);
and U10439 (N_10439,N_10305,N_10273);
xnor U10440 (N_10440,N_10328,N_10268);
nand U10441 (N_10441,N_10204,N_10265);
and U10442 (N_10442,N_10313,N_10258);
xor U10443 (N_10443,N_10215,N_10245);
nand U10444 (N_10444,N_10253,N_10333);
nand U10445 (N_10445,N_10206,N_10283);
nand U10446 (N_10446,N_10318,N_10268);
nor U10447 (N_10447,N_10220,N_10259);
or U10448 (N_10448,N_10280,N_10336);
xor U10449 (N_10449,N_10280,N_10278);
nand U10450 (N_10450,N_10232,N_10287);
nor U10451 (N_10451,N_10311,N_10309);
nand U10452 (N_10452,N_10339,N_10274);
and U10453 (N_10453,N_10262,N_10276);
and U10454 (N_10454,N_10235,N_10217);
xnor U10455 (N_10455,N_10312,N_10308);
nor U10456 (N_10456,N_10276,N_10250);
nor U10457 (N_10457,N_10315,N_10267);
or U10458 (N_10458,N_10299,N_10220);
nor U10459 (N_10459,N_10215,N_10338);
xor U10460 (N_10460,N_10252,N_10332);
nor U10461 (N_10461,N_10219,N_10244);
nor U10462 (N_10462,N_10277,N_10311);
nor U10463 (N_10463,N_10260,N_10244);
or U10464 (N_10464,N_10330,N_10297);
xnor U10465 (N_10465,N_10229,N_10320);
nand U10466 (N_10466,N_10222,N_10294);
nand U10467 (N_10467,N_10280,N_10226);
or U10468 (N_10468,N_10246,N_10325);
nand U10469 (N_10469,N_10314,N_10240);
and U10470 (N_10470,N_10296,N_10221);
or U10471 (N_10471,N_10314,N_10231);
or U10472 (N_10472,N_10348,N_10238);
nand U10473 (N_10473,N_10215,N_10221);
or U10474 (N_10474,N_10324,N_10232);
nor U10475 (N_10475,N_10303,N_10348);
xor U10476 (N_10476,N_10298,N_10274);
nand U10477 (N_10477,N_10201,N_10293);
nand U10478 (N_10478,N_10226,N_10302);
xnor U10479 (N_10479,N_10218,N_10304);
nand U10480 (N_10480,N_10243,N_10234);
or U10481 (N_10481,N_10248,N_10214);
nand U10482 (N_10482,N_10238,N_10327);
or U10483 (N_10483,N_10211,N_10294);
nor U10484 (N_10484,N_10299,N_10290);
nor U10485 (N_10485,N_10254,N_10334);
or U10486 (N_10486,N_10273,N_10231);
or U10487 (N_10487,N_10280,N_10337);
and U10488 (N_10488,N_10240,N_10207);
nand U10489 (N_10489,N_10228,N_10331);
nand U10490 (N_10490,N_10348,N_10230);
and U10491 (N_10491,N_10255,N_10340);
nand U10492 (N_10492,N_10250,N_10223);
and U10493 (N_10493,N_10227,N_10342);
xnor U10494 (N_10494,N_10238,N_10225);
nand U10495 (N_10495,N_10278,N_10321);
and U10496 (N_10496,N_10229,N_10238);
nand U10497 (N_10497,N_10206,N_10302);
or U10498 (N_10498,N_10295,N_10275);
or U10499 (N_10499,N_10339,N_10275);
and U10500 (N_10500,N_10405,N_10460);
nand U10501 (N_10501,N_10453,N_10440);
nor U10502 (N_10502,N_10470,N_10352);
or U10503 (N_10503,N_10379,N_10488);
or U10504 (N_10504,N_10441,N_10357);
and U10505 (N_10505,N_10475,N_10464);
nand U10506 (N_10506,N_10437,N_10457);
nand U10507 (N_10507,N_10393,N_10490);
nor U10508 (N_10508,N_10493,N_10424);
nor U10509 (N_10509,N_10499,N_10414);
and U10510 (N_10510,N_10413,N_10487);
xor U10511 (N_10511,N_10353,N_10383);
nand U10512 (N_10512,N_10403,N_10402);
xnor U10513 (N_10513,N_10395,N_10445);
or U10514 (N_10514,N_10369,N_10416);
nand U10515 (N_10515,N_10459,N_10367);
nand U10516 (N_10516,N_10438,N_10350);
and U10517 (N_10517,N_10461,N_10400);
nand U10518 (N_10518,N_10439,N_10496);
or U10519 (N_10519,N_10362,N_10430);
nand U10520 (N_10520,N_10390,N_10417);
nand U10521 (N_10521,N_10387,N_10363);
and U10522 (N_10522,N_10495,N_10486);
nor U10523 (N_10523,N_10492,N_10371);
nand U10524 (N_10524,N_10469,N_10355);
nand U10525 (N_10525,N_10386,N_10477);
nor U10526 (N_10526,N_10384,N_10426);
nand U10527 (N_10527,N_10370,N_10381);
nand U10528 (N_10528,N_10358,N_10435);
nor U10529 (N_10529,N_10449,N_10401);
nor U10530 (N_10530,N_10420,N_10415);
nand U10531 (N_10531,N_10497,N_10354);
nand U10532 (N_10532,N_10376,N_10423);
nand U10533 (N_10533,N_10432,N_10455);
and U10534 (N_10534,N_10473,N_10494);
xor U10535 (N_10535,N_10373,N_10452);
nand U10536 (N_10536,N_10408,N_10471);
and U10537 (N_10537,N_10482,N_10485);
nand U10538 (N_10538,N_10451,N_10454);
nand U10539 (N_10539,N_10377,N_10404);
xnor U10540 (N_10540,N_10388,N_10398);
xor U10541 (N_10541,N_10418,N_10365);
nor U10542 (N_10542,N_10442,N_10351);
nand U10543 (N_10543,N_10465,N_10450);
and U10544 (N_10544,N_10429,N_10456);
and U10545 (N_10545,N_10474,N_10422);
or U10546 (N_10546,N_10396,N_10412);
nand U10547 (N_10547,N_10491,N_10481);
nand U10548 (N_10548,N_10458,N_10436);
and U10549 (N_10549,N_10489,N_10479);
nand U10550 (N_10550,N_10483,N_10462);
nand U10551 (N_10551,N_10463,N_10394);
xnor U10552 (N_10552,N_10434,N_10410);
nand U10553 (N_10553,N_10372,N_10361);
xnor U10554 (N_10554,N_10406,N_10368);
nor U10555 (N_10555,N_10431,N_10467);
nor U10556 (N_10556,N_10380,N_10443);
nand U10557 (N_10557,N_10419,N_10411);
xnor U10558 (N_10558,N_10466,N_10399);
nand U10559 (N_10559,N_10364,N_10480);
nand U10560 (N_10560,N_10378,N_10407);
nand U10561 (N_10561,N_10374,N_10382);
xor U10562 (N_10562,N_10385,N_10446);
xnor U10563 (N_10563,N_10444,N_10359);
and U10564 (N_10564,N_10476,N_10391);
xnor U10565 (N_10565,N_10478,N_10356);
and U10566 (N_10566,N_10421,N_10447);
and U10567 (N_10567,N_10360,N_10428);
or U10568 (N_10568,N_10472,N_10366);
nand U10569 (N_10569,N_10392,N_10448);
xnor U10570 (N_10570,N_10498,N_10375);
nand U10571 (N_10571,N_10397,N_10389);
nand U10572 (N_10572,N_10484,N_10425);
nand U10573 (N_10573,N_10409,N_10433);
nand U10574 (N_10574,N_10468,N_10427);
nand U10575 (N_10575,N_10353,N_10491);
nor U10576 (N_10576,N_10389,N_10372);
nand U10577 (N_10577,N_10370,N_10425);
or U10578 (N_10578,N_10483,N_10397);
xor U10579 (N_10579,N_10380,N_10384);
and U10580 (N_10580,N_10395,N_10373);
or U10581 (N_10581,N_10409,N_10392);
and U10582 (N_10582,N_10378,N_10393);
and U10583 (N_10583,N_10356,N_10359);
xor U10584 (N_10584,N_10468,N_10480);
nor U10585 (N_10585,N_10429,N_10384);
xnor U10586 (N_10586,N_10356,N_10475);
nor U10587 (N_10587,N_10393,N_10408);
nand U10588 (N_10588,N_10409,N_10489);
nand U10589 (N_10589,N_10486,N_10369);
nand U10590 (N_10590,N_10385,N_10444);
nand U10591 (N_10591,N_10404,N_10366);
nor U10592 (N_10592,N_10420,N_10412);
nor U10593 (N_10593,N_10375,N_10426);
nor U10594 (N_10594,N_10423,N_10385);
or U10595 (N_10595,N_10429,N_10417);
nor U10596 (N_10596,N_10439,N_10471);
nor U10597 (N_10597,N_10440,N_10406);
and U10598 (N_10598,N_10422,N_10418);
or U10599 (N_10599,N_10443,N_10368);
and U10600 (N_10600,N_10408,N_10396);
nor U10601 (N_10601,N_10450,N_10452);
nand U10602 (N_10602,N_10387,N_10375);
or U10603 (N_10603,N_10468,N_10440);
or U10604 (N_10604,N_10440,N_10357);
nor U10605 (N_10605,N_10411,N_10365);
xor U10606 (N_10606,N_10385,N_10394);
nand U10607 (N_10607,N_10494,N_10356);
and U10608 (N_10608,N_10402,N_10489);
and U10609 (N_10609,N_10442,N_10443);
xnor U10610 (N_10610,N_10360,N_10453);
xor U10611 (N_10611,N_10386,N_10483);
xnor U10612 (N_10612,N_10435,N_10426);
xnor U10613 (N_10613,N_10357,N_10449);
xnor U10614 (N_10614,N_10436,N_10369);
xnor U10615 (N_10615,N_10374,N_10367);
or U10616 (N_10616,N_10460,N_10426);
xor U10617 (N_10617,N_10497,N_10485);
xnor U10618 (N_10618,N_10387,N_10468);
nand U10619 (N_10619,N_10394,N_10361);
or U10620 (N_10620,N_10357,N_10427);
or U10621 (N_10621,N_10394,N_10366);
or U10622 (N_10622,N_10453,N_10416);
or U10623 (N_10623,N_10363,N_10392);
xnor U10624 (N_10624,N_10377,N_10497);
xnor U10625 (N_10625,N_10455,N_10404);
nand U10626 (N_10626,N_10350,N_10481);
or U10627 (N_10627,N_10367,N_10387);
xor U10628 (N_10628,N_10494,N_10460);
nor U10629 (N_10629,N_10487,N_10445);
or U10630 (N_10630,N_10401,N_10382);
xor U10631 (N_10631,N_10352,N_10465);
and U10632 (N_10632,N_10367,N_10392);
nor U10633 (N_10633,N_10372,N_10396);
nand U10634 (N_10634,N_10374,N_10478);
or U10635 (N_10635,N_10443,N_10490);
xnor U10636 (N_10636,N_10452,N_10488);
and U10637 (N_10637,N_10371,N_10406);
nor U10638 (N_10638,N_10457,N_10423);
xnor U10639 (N_10639,N_10427,N_10485);
nor U10640 (N_10640,N_10459,N_10456);
nor U10641 (N_10641,N_10401,N_10394);
xnor U10642 (N_10642,N_10401,N_10377);
and U10643 (N_10643,N_10488,N_10450);
xor U10644 (N_10644,N_10426,N_10417);
and U10645 (N_10645,N_10430,N_10484);
and U10646 (N_10646,N_10436,N_10463);
nor U10647 (N_10647,N_10481,N_10367);
and U10648 (N_10648,N_10362,N_10397);
xnor U10649 (N_10649,N_10355,N_10400);
nand U10650 (N_10650,N_10553,N_10557);
and U10651 (N_10651,N_10566,N_10588);
nand U10652 (N_10652,N_10520,N_10549);
xnor U10653 (N_10653,N_10603,N_10550);
nand U10654 (N_10654,N_10598,N_10634);
nor U10655 (N_10655,N_10518,N_10514);
and U10656 (N_10656,N_10546,N_10500);
xnor U10657 (N_10657,N_10513,N_10551);
nor U10658 (N_10658,N_10646,N_10534);
or U10659 (N_10659,N_10610,N_10558);
xnor U10660 (N_10660,N_10586,N_10570);
nand U10661 (N_10661,N_10502,N_10568);
and U10662 (N_10662,N_10515,N_10621);
nand U10663 (N_10663,N_10629,N_10583);
nand U10664 (N_10664,N_10615,N_10567);
nor U10665 (N_10665,N_10626,N_10531);
xor U10666 (N_10666,N_10597,N_10563);
and U10667 (N_10667,N_10508,N_10640);
nand U10668 (N_10668,N_10530,N_10596);
nor U10669 (N_10669,N_10647,N_10645);
or U10670 (N_10670,N_10503,N_10639);
nand U10671 (N_10671,N_10554,N_10602);
and U10672 (N_10672,N_10613,N_10556);
or U10673 (N_10673,N_10637,N_10512);
nor U10674 (N_10674,N_10614,N_10577);
xor U10675 (N_10675,N_10519,N_10616);
or U10676 (N_10676,N_10540,N_10587);
or U10677 (N_10677,N_10590,N_10611);
or U10678 (N_10678,N_10607,N_10565);
nor U10679 (N_10679,N_10585,N_10618);
nand U10680 (N_10680,N_10505,N_10578);
nor U10681 (N_10681,N_10525,N_10533);
xor U10682 (N_10682,N_10623,N_10604);
and U10683 (N_10683,N_10605,N_10573);
nand U10684 (N_10684,N_10506,N_10561);
xnor U10685 (N_10685,N_10589,N_10544);
nand U10686 (N_10686,N_10593,N_10641);
and U10687 (N_10687,N_10552,N_10507);
xnor U10688 (N_10688,N_10580,N_10523);
and U10689 (N_10689,N_10582,N_10638);
nand U10690 (N_10690,N_10628,N_10541);
nor U10691 (N_10691,N_10545,N_10526);
nor U10692 (N_10692,N_10547,N_10581);
and U10693 (N_10693,N_10542,N_10584);
xor U10694 (N_10694,N_10608,N_10532);
xnor U10695 (N_10695,N_10627,N_10575);
nor U10696 (N_10696,N_10632,N_10521);
or U10697 (N_10697,N_10600,N_10606);
nor U10698 (N_10698,N_10648,N_10599);
and U10699 (N_10699,N_10501,N_10511);
nand U10700 (N_10700,N_10559,N_10594);
nor U10701 (N_10701,N_10631,N_10562);
and U10702 (N_10702,N_10636,N_10516);
nor U10703 (N_10703,N_10509,N_10569);
xor U10704 (N_10704,N_10504,N_10535);
or U10705 (N_10705,N_10617,N_10649);
and U10706 (N_10706,N_10510,N_10644);
nor U10707 (N_10707,N_10527,N_10543);
nor U10708 (N_10708,N_10524,N_10625);
or U10709 (N_10709,N_10522,N_10571);
or U10710 (N_10710,N_10538,N_10564);
nand U10711 (N_10711,N_10517,N_10560);
or U10712 (N_10712,N_10537,N_10574);
nand U10713 (N_10713,N_10635,N_10624);
or U10714 (N_10714,N_10592,N_10619);
xnor U10715 (N_10715,N_10548,N_10601);
nand U10716 (N_10716,N_10579,N_10576);
and U10717 (N_10717,N_10630,N_10643);
xnor U10718 (N_10718,N_10620,N_10622);
and U10719 (N_10719,N_10591,N_10528);
xor U10720 (N_10720,N_10539,N_10572);
nand U10721 (N_10721,N_10529,N_10555);
nor U10722 (N_10722,N_10609,N_10536);
nand U10723 (N_10723,N_10612,N_10595);
nand U10724 (N_10724,N_10633,N_10642);
nor U10725 (N_10725,N_10623,N_10510);
xnor U10726 (N_10726,N_10513,N_10541);
and U10727 (N_10727,N_10510,N_10593);
nor U10728 (N_10728,N_10581,N_10573);
xor U10729 (N_10729,N_10571,N_10628);
and U10730 (N_10730,N_10616,N_10518);
or U10731 (N_10731,N_10561,N_10529);
xor U10732 (N_10732,N_10518,N_10647);
nor U10733 (N_10733,N_10628,N_10519);
or U10734 (N_10734,N_10596,N_10632);
nand U10735 (N_10735,N_10626,N_10563);
and U10736 (N_10736,N_10624,N_10622);
and U10737 (N_10737,N_10636,N_10550);
nor U10738 (N_10738,N_10649,N_10511);
nand U10739 (N_10739,N_10572,N_10529);
nand U10740 (N_10740,N_10542,N_10629);
xor U10741 (N_10741,N_10603,N_10500);
xor U10742 (N_10742,N_10591,N_10545);
or U10743 (N_10743,N_10511,N_10604);
nand U10744 (N_10744,N_10561,N_10542);
nor U10745 (N_10745,N_10513,N_10629);
or U10746 (N_10746,N_10562,N_10610);
nor U10747 (N_10747,N_10511,N_10534);
and U10748 (N_10748,N_10624,N_10535);
and U10749 (N_10749,N_10503,N_10553);
and U10750 (N_10750,N_10555,N_10599);
xnor U10751 (N_10751,N_10593,N_10616);
and U10752 (N_10752,N_10582,N_10513);
and U10753 (N_10753,N_10645,N_10614);
nand U10754 (N_10754,N_10505,N_10588);
nand U10755 (N_10755,N_10535,N_10626);
nor U10756 (N_10756,N_10523,N_10534);
xor U10757 (N_10757,N_10607,N_10554);
nor U10758 (N_10758,N_10571,N_10598);
or U10759 (N_10759,N_10503,N_10557);
xor U10760 (N_10760,N_10523,N_10537);
and U10761 (N_10761,N_10588,N_10561);
xor U10762 (N_10762,N_10615,N_10557);
xnor U10763 (N_10763,N_10558,N_10594);
xor U10764 (N_10764,N_10577,N_10543);
or U10765 (N_10765,N_10553,N_10575);
or U10766 (N_10766,N_10527,N_10591);
and U10767 (N_10767,N_10547,N_10510);
xor U10768 (N_10768,N_10649,N_10529);
nor U10769 (N_10769,N_10613,N_10574);
nor U10770 (N_10770,N_10520,N_10640);
nor U10771 (N_10771,N_10614,N_10597);
or U10772 (N_10772,N_10638,N_10532);
or U10773 (N_10773,N_10524,N_10561);
nor U10774 (N_10774,N_10527,N_10573);
or U10775 (N_10775,N_10623,N_10533);
nand U10776 (N_10776,N_10549,N_10577);
xor U10777 (N_10777,N_10640,N_10555);
xnor U10778 (N_10778,N_10501,N_10533);
and U10779 (N_10779,N_10581,N_10606);
nand U10780 (N_10780,N_10615,N_10600);
and U10781 (N_10781,N_10514,N_10636);
nor U10782 (N_10782,N_10607,N_10590);
nand U10783 (N_10783,N_10586,N_10529);
nor U10784 (N_10784,N_10647,N_10568);
nor U10785 (N_10785,N_10556,N_10559);
or U10786 (N_10786,N_10577,N_10550);
nor U10787 (N_10787,N_10538,N_10588);
nor U10788 (N_10788,N_10612,N_10601);
xnor U10789 (N_10789,N_10616,N_10547);
nand U10790 (N_10790,N_10545,N_10649);
nand U10791 (N_10791,N_10600,N_10555);
nor U10792 (N_10792,N_10537,N_10606);
or U10793 (N_10793,N_10537,N_10506);
xnor U10794 (N_10794,N_10573,N_10592);
nand U10795 (N_10795,N_10510,N_10609);
nand U10796 (N_10796,N_10507,N_10533);
and U10797 (N_10797,N_10514,N_10545);
nand U10798 (N_10798,N_10538,N_10500);
xnor U10799 (N_10799,N_10534,N_10554);
nand U10800 (N_10800,N_10706,N_10667);
nor U10801 (N_10801,N_10660,N_10747);
nor U10802 (N_10802,N_10704,N_10766);
nand U10803 (N_10803,N_10793,N_10777);
xnor U10804 (N_10804,N_10764,N_10701);
and U10805 (N_10805,N_10705,N_10661);
xor U10806 (N_10806,N_10714,N_10776);
nand U10807 (N_10807,N_10691,N_10670);
and U10808 (N_10808,N_10746,N_10737);
and U10809 (N_10809,N_10708,N_10692);
and U10810 (N_10810,N_10707,N_10712);
or U10811 (N_10811,N_10674,N_10785);
nor U10812 (N_10812,N_10659,N_10763);
xnor U10813 (N_10813,N_10767,N_10745);
and U10814 (N_10814,N_10735,N_10789);
or U10815 (N_10815,N_10754,N_10687);
and U10816 (N_10816,N_10666,N_10734);
nand U10817 (N_10817,N_10662,N_10679);
nor U10818 (N_10818,N_10696,N_10681);
nor U10819 (N_10819,N_10749,N_10740);
nand U10820 (N_10820,N_10653,N_10682);
xor U10821 (N_10821,N_10782,N_10757);
nand U10822 (N_10822,N_10695,N_10664);
xnor U10823 (N_10823,N_10726,N_10671);
xor U10824 (N_10824,N_10773,N_10731);
and U10825 (N_10825,N_10711,N_10694);
xnor U10826 (N_10826,N_10724,N_10713);
xnor U10827 (N_10827,N_10718,N_10794);
nor U10828 (N_10828,N_10790,N_10693);
and U10829 (N_10829,N_10676,N_10672);
nand U10830 (N_10830,N_10750,N_10759);
xnor U10831 (N_10831,N_10795,N_10723);
nor U10832 (N_10832,N_10748,N_10698);
nand U10833 (N_10833,N_10744,N_10733);
and U10834 (N_10834,N_10663,N_10760);
or U10835 (N_10835,N_10739,N_10697);
or U10836 (N_10836,N_10656,N_10689);
and U10837 (N_10837,N_10729,N_10783);
or U10838 (N_10838,N_10797,N_10652);
and U10839 (N_10839,N_10673,N_10732);
and U10840 (N_10840,N_10770,N_10703);
nand U10841 (N_10841,N_10774,N_10772);
xnor U10842 (N_10842,N_10799,N_10686);
or U10843 (N_10843,N_10784,N_10680);
xnor U10844 (N_10844,N_10781,N_10752);
and U10845 (N_10845,N_10651,N_10775);
and U10846 (N_10846,N_10650,N_10677);
nor U10847 (N_10847,N_10758,N_10768);
xor U10848 (N_10848,N_10721,N_10669);
nand U10849 (N_10849,N_10738,N_10716);
nand U10850 (N_10850,N_10778,N_10769);
xor U10851 (N_10851,N_10771,N_10655);
and U10852 (N_10852,N_10709,N_10720);
or U10853 (N_10853,N_10717,N_10791);
or U10854 (N_10854,N_10762,N_10780);
nand U10855 (N_10855,N_10657,N_10796);
nand U10856 (N_10856,N_10741,N_10690);
and U10857 (N_10857,N_10787,N_10719);
and U10858 (N_10858,N_10668,N_10710);
or U10859 (N_10859,N_10753,N_10665);
or U10860 (N_10860,N_10699,N_10722);
or U10861 (N_10861,N_10678,N_10779);
xnor U10862 (N_10862,N_10742,N_10756);
and U10863 (N_10863,N_10730,N_10751);
nand U10864 (N_10864,N_10715,N_10702);
or U10865 (N_10865,N_10658,N_10792);
and U10866 (N_10866,N_10725,N_10755);
nand U10867 (N_10867,N_10798,N_10736);
and U10868 (N_10868,N_10765,N_10688);
nand U10869 (N_10869,N_10685,N_10654);
xor U10870 (N_10870,N_10743,N_10683);
and U10871 (N_10871,N_10727,N_10786);
nand U10872 (N_10872,N_10675,N_10728);
xor U10873 (N_10873,N_10684,N_10788);
or U10874 (N_10874,N_10761,N_10700);
nor U10875 (N_10875,N_10763,N_10790);
xnor U10876 (N_10876,N_10684,N_10798);
nor U10877 (N_10877,N_10689,N_10662);
and U10878 (N_10878,N_10729,N_10741);
xor U10879 (N_10879,N_10782,N_10772);
nand U10880 (N_10880,N_10740,N_10773);
and U10881 (N_10881,N_10662,N_10675);
nand U10882 (N_10882,N_10758,N_10676);
or U10883 (N_10883,N_10773,N_10732);
and U10884 (N_10884,N_10779,N_10702);
and U10885 (N_10885,N_10683,N_10668);
or U10886 (N_10886,N_10700,N_10654);
and U10887 (N_10887,N_10678,N_10651);
and U10888 (N_10888,N_10656,N_10799);
xnor U10889 (N_10889,N_10730,N_10693);
or U10890 (N_10890,N_10758,N_10679);
or U10891 (N_10891,N_10751,N_10790);
nand U10892 (N_10892,N_10698,N_10710);
xor U10893 (N_10893,N_10685,N_10693);
nand U10894 (N_10894,N_10681,N_10772);
xor U10895 (N_10895,N_10726,N_10650);
nor U10896 (N_10896,N_10790,N_10705);
xor U10897 (N_10897,N_10735,N_10725);
nand U10898 (N_10898,N_10704,N_10682);
nand U10899 (N_10899,N_10759,N_10711);
nor U10900 (N_10900,N_10759,N_10738);
xnor U10901 (N_10901,N_10703,N_10685);
xor U10902 (N_10902,N_10711,N_10710);
or U10903 (N_10903,N_10654,N_10653);
nand U10904 (N_10904,N_10663,N_10778);
nand U10905 (N_10905,N_10768,N_10723);
and U10906 (N_10906,N_10666,N_10655);
nand U10907 (N_10907,N_10774,N_10754);
and U10908 (N_10908,N_10766,N_10752);
or U10909 (N_10909,N_10740,N_10736);
and U10910 (N_10910,N_10685,N_10795);
and U10911 (N_10911,N_10743,N_10754);
xnor U10912 (N_10912,N_10694,N_10735);
and U10913 (N_10913,N_10663,N_10795);
xnor U10914 (N_10914,N_10781,N_10713);
xnor U10915 (N_10915,N_10670,N_10759);
nand U10916 (N_10916,N_10655,N_10767);
or U10917 (N_10917,N_10687,N_10681);
or U10918 (N_10918,N_10752,N_10696);
nand U10919 (N_10919,N_10701,N_10664);
xnor U10920 (N_10920,N_10693,N_10792);
nand U10921 (N_10921,N_10750,N_10687);
nor U10922 (N_10922,N_10730,N_10794);
nand U10923 (N_10923,N_10770,N_10731);
and U10924 (N_10924,N_10702,N_10760);
xnor U10925 (N_10925,N_10697,N_10650);
and U10926 (N_10926,N_10757,N_10653);
and U10927 (N_10927,N_10691,N_10777);
or U10928 (N_10928,N_10748,N_10783);
or U10929 (N_10929,N_10653,N_10691);
nand U10930 (N_10930,N_10752,N_10674);
or U10931 (N_10931,N_10754,N_10684);
xnor U10932 (N_10932,N_10674,N_10758);
nand U10933 (N_10933,N_10691,N_10696);
nand U10934 (N_10934,N_10729,N_10773);
xor U10935 (N_10935,N_10778,N_10747);
nand U10936 (N_10936,N_10660,N_10665);
and U10937 (N_10937,N_10782,N_10674);
or U10938 (N_10938,N_10798,N_10796);
nand U10939 (N_10939,N_10752,N_10774);
nor U10940 (N_10940,N_10713,N_10674);
nor U10941 (N_10941,N_10711,N_10651);
and U10942 (N_10942,N_10792,N_10651);
xor U10943 (N_10943,N_10701,N_10722);
nor U10944 (N_10944,N_10733,N_10717);
nand U10945 (N_10945,N_10702,N_10706);
nand U10946 (N_10946,N_10712,N_10770);
or U10947 (N_10947,N_10706,N_10756);
nor U10948 (N_10948,N_10679,N_10736);
xor U10949 (N_10949,N_10695,N_10710);
xor U10950 (N_10950,N_10914,N_10821);
and U10951 (N_10951,N_10836,N_10938);
nand U10952 (N_10952,N_10901,N_10861);
nand U10953 (N_10953,N_10831,N_10838);
and U10954 (N_10954,N_10925,N_10824);
xor U10955 (N_10955,N_10812,N_10937);
and U10956 (N_10956,N_10826,N_10935);
nand U10957 (N_10957,N_10845,N_10895);
nand U10958 (N_10958,N_10857,N_10884);
xor U10959 (N_10959,N_10939,N_10830);
and U10960 (N_10960,N_10891,N_10802);
nor U10961 (N_10961,N_10936,N_10899);
nand U10962 (N_10962,N_10806,N_10909);
xor U10963 (N_10963,N_10819,N_10877);
or U10964 (N_10964,N_10881,N_10853);
xnor U10965 (N_10965,N_10894,N_10848);
nand U10966 (N_10966,N_10888,N_10932);
xnor U10967 (N_10967,N_10869,N_10858);
xnor U10968 (N_10968,N_10942,N_10887);
and U10969 (N_10969,N_10940,N_10911);
xnor U10970 (N_10970,N_10863,N_10832);
or U10971 (N_10971,N_10929,N_10828);
nor U10972 (N_10972,N_10902,N_10804);
and U10973 (N_10973,N_10800,N_10920);
and U10974 (N_10974,N_10834,N_10871);
and U10975 (N_10975,N_10846,N_10870);
xor U10976 (N_10976,N_10842,N_10916);
nor U10977 (N_10977,N_10885,N_10878);
nand U10978 (N_10978,N_10900,N_10837);
and U10979 (N_10979,N_10801,N_10825);
nor U10980 (N_10980,N_10873,N_10944);
xnor U10981 (N_10981,N_10903,N_10913);
nand U10982 (N_10982,N_10809,N_10866);
nand U10983 (N_10983,N_10917,N_10924);
xor U10984 (N_10984,N_10930,N_10813);
nor U10985 (N_10985,N_10859,N_10840);
nand U10986 (N_10986,N_10921,N_10855);
nand U10987 (N_10987,N_10815,N_10822);
nor U10988 (N_10988,N_10880,N_10898);
xor U10989 (N_10989,N_10945,N_10949);
nand U10990 (N_10990,N_10931,N_10864);
and U10991 (N_10991,N_10868,N_10896);
xor U10992 (N_10992,N_10919,N_10892);
or U10993 (N_10993,N_10811,N_10943);
and U10994 (N_10994,N_10839,N_10912);
nor U10995 (N_10995,N_10807,N_10829);
and U10996 (N_10996,N_10854,N_10803);
nand U10997 (N_10997,N_10875,N_10862);
or U10998 (N_10998,N_10927,N_10850);
xor U10999 (N_10999,N_10923,N_10820);
nor U11000 (N_11000,N_10876,N_10841);
nand U11001 (N_11001,N_10843,N_10946);
nor U11002 (N_11002,N_10860,N_10814);
xnor U11003 (N_11003,N_10890,N_10910);
nor U11004 (N_11004,N_10897,N_10879);
nand U11005 (N_11005,N_10844,N_10918);
or U11006 (N_11006,N_10847,N_10882);
and U11007 (N_11007,N_10893,N_10904);
xnor U11008 (N_11008,N_10810,N_10905);
nand U11009 (N_11009,N_10856,N_10865);
nor U11010 (N_11010,N_10933,N_10874);
nor U11011 (N_11011,N_10908,N_10805);
nand U11012 (N_11012,N_10827,N_10872);
nor U11013 (N_11013,N_10889,N_10852);
xor U11014 (N_11014,N_10886,N_10947);
nand U11015 (N_11015,N_10851,N_10808);
nand U11016 (N_11016,N_10922,N_10934);
and U11017 (N_11017,N_10915,N_10906);
xnor U11018 (N_11018,N_10817,N_10867);
nand U11019 (N_11019,N_10926,N_10823);
and U11020 (N_11020,N_10833,N_10907);
nor U11021 (N_11021,N_10816,N_10941);
and U11022 (N_11022,N_10928,N_10883);
nand U11023 (N_11023,N_10835,N_10818);
or U11024 (N_11024,N_10948,N_10849);
xnor U11025 (N_11025,N_10904,N_10855);
or U11026 (N_11026,N_10827,N_10805);
xnor U11027 (N_11027,N_10944,N_10879);
or U11028 (N_11028,N_10925,N_10822);
nor U11029 (N_11029,N_10913,N_10879);
xnor U11030 (N_11030,N_10823,N_10915);
and U11031 (N_11031,N_10856,N_10807);
or U11032 (N_11032,N_10839,N_10949);
and U11033 (N_11033,N_10880,N_10919);
nor U11034 (N_11034,N_10941,N_10910);
or U11035 (N_11035,N_10928,N_10875);
and U11036 (N_11036,N_10916,N_10945);
and U11037 (N_11037,N_10908,N_10810);
or U11038 (N_11038,N_10883,N_10820);
or U11039 (N_11039,N_10847,N_10916);
xnor U11040 (N_11040,N_10834,N_10906);
nand U11041 (N_11041,N_10846,N_10944);
or U11042 (N_11042,N_10861,N_10927);
nand U11043 (N_11043,N_10856,N_10851);
nand U11044 (N_11044,N_10914,N_10917);
nor U11045 (N_11045,N_10902,N_10843);
or U11046 (N_11046,N_10915,N_10850);
nand U11047 (N_11047,N_10924,N_10843);
and U11048 (N_11048,N_10833,N_10803);
and U11049 (N_11049,N_10901,N_10850);
xor U11050 (N_11050,N_10829,N_10912);
nor U11051 (N_11051,N_10900,N_10875);
or U11052 (N_11052,N_10837,N_10946);
nor U11053 (N_11053,N_10948,N_10810);
or U11054 (N_11054,N_10885,N_10806);
xor U11055 (N_11055,N_10877,N_10938);
nor U11056 (N_11056,N_10869,N_10935);
and U11057 (N_11057,N_10841,N_10821);
xor U11058 (N_11058,N_10806,N_10819);
nand U11059 (N_11059,N_10836,N_10846);
nand U11060 (N_11060,N_10935,N_10839);
nand U11061 (N_11061,N_10858,N_10828);
xor U11062 (N_11062,N_10880,N_10854);
xor U11063 (N_11063,N_10910,N_10881);
or U11064 (N_11064,N_10810,N_10858);
and U11065 (N_11065,N_10889,N_10801);
or U11066 (N_11066,N_10805,N_10818);
xnor U11067 (N_11067,N_10804,N_10806);
nand U11068 (N_11068,N_10937,N_10804);
xor U11069 (N_11069,N_10916,N_10888);
xor U11070 (N_11070,N_10913,N_10947);
nor U11071 (N_11071,N_10843,N_10853);
or U11072 (N_11072,N_10918,N_10879);
xnor U11073 (N_11073,N_10823,N_10876);
and U11074 (N_11074,N_10836,N_10805);
or U11075 (N_11075,N_10880,N_10835);
or U11076 (N_11076,N_10876,N_10889);
nor U11077 (N_11077,N_10830,N_10918);
nand U11078 (N_11078,N_10860,N_10810);
xnor U11079 (N_11079,N_10825,N_10861);
nor U11080 (N_11080,N_10845,N_10824);
or U11081 (N_11081,N_10870,N_10819);
nand U11082 (N_11082,N_10912,N_10896);
xor U11083 (N_11083,N_10895,N_10827);
nor U11084 (N_11084,N_10885,N_10838);
nor U11085 (N_11085,N_10937,N_10871);
and U11086 (N_11086,N_10844,N_10828);
or U11087 (N_11087,N_10831,N_10885);
xor U11088 (N_11088,N_10810,N_10814);
and U11089 (N_11089,N_10830,N_10857);
nor U11090 (N_11090,N_10864,N_10832);
nand U11091 (N_11091,N_10861,N_10836);
and U11092 (N_11092,N_10822,N_10932);
nand U11093 (N_11093,N_10915,N_10808);
nand U11094 (N_11094,N_10846,N_10850);
nand U11095 (N_11095,N_10841,N_10839);
and U11096 (N_11096,N_10898,N_10895);
xnor U11097 (N_11097,N_10816,N_10844);
xor U11098 (N_11098,N_10830,N_10927);
nand U11099 (N_11099,N_10905,N_10941);
nor U11100 (N_11100,N_10995,N_11041);
xnor U11101 (N_11101,N_11005,N_11004);
nand U11102 (N_11102,N_10956,N_10960);
nand U11103 (N_11103,N_11019,N_10984);
nor U11104 (N_11104,N_11010,N_11097);
and U11105 (N_11105,N_10978,N_11084);
nor U11106 (N_11106,N_11043,N_11001);
nor U11107 (N_11107,N_11095,N_11098);
nor U11108 (N_11108,N_11058,N_11065);
or U11109 (N_11109,N_11034,N_11025);
xnor U11110 (N_11110,N_11020,N_11032);
xnor U11111 (N_11111,N_11042,N_10991);
nand U11112 (N_11112,N_10977,N_10997);
nor U11113 (N_11113,N_10953,N_11055);
or U11114 (N_11114,N_11014,N_11089);
and U11115 (N_11115,N_11096,N_11062);
or U11116 (N_11116,N_11064,N_11052);
nor U11117 (N_11117,N_11056,N_10965);
or U11118 (N_11118,N_11008,N_10976);
or U11119 (N_11119,N_10996,N_11057);
and U11120 (N_11120,N_11093,N_11028);
or U11121 (N_11121,N_11018,N_11031);
and U11122 (N_11122,N_11072,N_11080);
or U11123 (N_11123,N_11037,N_11012);
and U11124 (N_11124,N_11090,N_10955);
and U11125 (N_11125,N_11051,N_11033);
xnor U11126 (N_11126,N_11044,N_11007);
xor U11127 (N_11127,N_11000,N_11036);
nand U11128 (N_11128,N_10985,N_10967);
nand U11129 (N_11129,N_11040,N_11076);
and U11130 (N_11130,N_11047,N_11071);
nor U11131 (N_11131,N_10962,N_11024);
and U11132 (N_11132,N_11049,N_11068);
or U11133 (N_11133,N_10987,N_11092);
xor U11134 (N_11134,N_10968,N_10981);
xnor U11135 (N_11135,N_11039,N_10958);
nor U11136 (N_11136,N_10998,N_10993);
xnor U11137 (N_11137,N_11022,N_10966);
nor U11138 (N_11138,N_11046,N_11099);
and U11139 (N_11139,N_10970,N_11015);
or U11140 (N_11140,N_10974,N_11077);
nand U11141 (N_11141,N_11023,N_11091);
nor U11142 (N_11142,N_11002,N_10988);
nand U11143 (N_11143,N_10975,N_11073);
xor U11144 (N_11144,N_11038,N_11003);
or U11145 (N_11145,N_11035,N_11066);
and U11146 (N_11146,N_11067,N_10999);
or U11147 (N_11147,N_11060,N_11045);
nor U11148 (N_11148,N_11081,N_10986);
xor U11149 (N_11149,N_10964,N_11026);
and U11150 (N_11150,N_11009,N_11021);
xor U11151 (N_11151,N_11054,N_11016);
xor U11152 (N_11152,N_10994,N_10951);
nand U11153 (N_11153,N_10973,N_10982);
xor U11154 (N_11154,N_11070,N_10961);
and U11155 (N_11155,N_10972,N_11050);
nand U11156 (N_11156,N_11063,N_11069);
xor U11157 (N_11157,N_10957,N_11075);
or U11158 (N_11158,N_11013,N_10959);
nor U11159 (N_11159,N_11094,N_11078);
nor U11160 (N_11160,N_10952,N_10980);
and U11161 (N_11161,N_10963,N_11030);
or U11162 (N_11162,N_11086,N_11079);
xnor U11163 (N_11163,N_11059,N_10954);
and U11164 (N_11164,N_10983,N_11029);
nor U11165 (N_11165,N_11017,N_11027);
nor U11166 (N_11166,N_11011,N_11074);
nor U11167 (N_11167,N_10989,N_11083);
nor U11168 (N_11168,N_11006,N_10992);
nand U11169 (N_11169,N_10990,N_10979);
nand U11170 (N_11170,N_10969,N_11082);
xnor U11171 (N_11171,N_11048,N_11088);
nand U11172 (N_11172,N_11061,N_10950);
nand U11173 (N_11173,N_11053,N_11085);
or U11174 (N_11174,N_10971,N_11087);
nor U11175 (N_11175,N_11090,N_11062);
xnor U11176 (N_11176,N_11019,N_11045);
or U11177 (N_11177,N_11076,N_11099);
and U11178 (N_11178,N_11075,N_11004);
nor U11179 (N_11179,N_11067,N_11031);
xor U11180 (N_11180,N_10980,N_11075);
or U11181 (N_11181,N_11025,N_11038);
xor U11182 (N_11182,N_11013,N_10982);
or U11183 (N_11183,N_11080,N_10974);
xnor U11184 (N_11184,N_11042,N_11044);
and U11185 (N_11185,N_11038,N_11054);
nor U11186 (N_11186,N_11045,N_10955);
and U11187 (N_11187,N_11051,N_10978);
nand U11188 (N_11188,N_11035,N_11002);
nor U11189 (N_11189,N_11095,N_11062);
or U11190 (N_11190,N_10993,N_11061);
nand U11191 (N_11191,N_11064,N_11036);
nand U11192 (N_11192,N_11047,N_10965);
xnor U11193 (N_11193,N_11048,N_11060);
nand U11194 (N_11194,N_11011,N_11065);
or U11195 (N_11195,N_11058,N_10952);
xnor U11196 (N_11196,N_10994,N_10960);
nand U11197 (N_11197,N_11029,N_10958);
and U11198 (N_11198,N_10966,N_10956);
nand U11199 (N_11199,N_10985,N_10968);
nand U11200 (N_11200,N_11060,N_11020);
nor U11201 (N_11201,N_11048,N_10973);
nand U11202 (N_11202,N_11094,N_10981);
nor U11203 (N_11203,N_11086,N_11057);
or U11204 (N_11204,N_11095,N_11028);
xnor U11205 (N_11205,N_11003,N_11018);
and U11206 (N_11206,N_11095,N_11012);
nand U11207 (N_11207,N_11031,N_10961);
and U11208 (N_11208,N_10990,N_10950);
nand U11209 (N_11209,N_10953,N_10964);
or U11210 (N_11210,N_11084,N_11057);
nor U11211 (N_11211,N_11033,N_11062);
nor U11212 (N_11212,N_11060,N_11006);
xnor U11213 (N_11213,N_11046,N_11027);
xor U11214 (N_11214,N_11053,N_10958);
nand U11215 (N_11215,N_11056,N_11060);
or U11216 (N_11216,N_11074,N_11037);
or U11217 (N_11217,N_10955,N_11088);
nor U11218 (N_11218,N_10954,N_11013);
and U11219 (N_11219,N_11038,N_11091);
or U11220 (N_11220,N_10957,N_11060);
nand U11221 (N_11221,N_11008,N_11077);
nand U11222 (N_11222,N_11033,N_11037);
nand U11223 (N_11223,N_11004,N_11030);
nor U11224 (N_11224,N_11064,N_11023);
or U11225 (N_11225,N_11083,N_10979);
xor U11226 (N_11226,N_10957,N_11030);
nand U11227 (N_11227,N_11028,N_10954);
and U11228 (N_11228,N_10970,N_11075);
nor U11229 (N_11229,N_11094,N_10982);
nand U11230 (N_11230,N_11048,N_10995);
xnor U11231 (N_11231,N_11051,N_11020);
nor U11232 (N_11232,N_11085,N_11037);
xor U11233 (N_11233,N_11060,N_11063);
xnor U11234 (N_11234,N_11022,N_11029);
xnor U11235 (N_11235,N_11015,N_11045);
and U11236 (N_11236,N_11060,N_11069);
nand U11237 (N_11237,N_11032,N_11078);
or U11238 (N_11238,N_11012,N_10971);
nor U11239 (N_11239,N_11096,N_10961);
xor U11240 (N_11240,N_11051,N_10989);
or U11241 (N_11241,N_11089,N_11091);
nor U11242 (N_11242,N_11097,N_11013);
nor U11243 (N_11243,N_10973,N_10976);
and U11244 (N_11244,N_11065,N_11022);
nand U11245 (N_11245,N_11092,N_11049);
nor U11246 (N_11246,N_11031,N_10965);
xnor U11247 (N_11247,N_11014,N_11003);
and U11248 (N_11248,N_11035,N_10980);
nand U11249 (N_11249,N_11038,N_11057);
or U11250 (N_11250,N_11129,N_11124);
nor U11251 (N_11251,N_11199,N_11155);
nand U11252 (N_11252,N_11176,N_11216);
xnor U11253 (N_11253,N_11131,N_11117);
or U11254 (N_11254,N_11148,N_11239);
or U11255 (N_11255,N_11163,N_11231);
nand U11256 (N_11256,N_11197,N_11198);
or U11257 (N_11257,N_11234,N_11185);
xor U11258 (N_11258,N_11146,N_11166);
or U11259 (N_11259,N_11217,N_11100);
and U11260 (N_11260,N_11107,N_11210);
nand U11261 (N_11261,N_11211,N_11133);
or U11262 (N_11262,N_11174,N_11167);
xor U11263 (N_11263,N_11147,N_11161);
or U11264 (N_11264,N_11201,N_11221);
or U11265 (N_11265,N_11249,N_11108);
and U11266 (N_11266,N_11156,N_11180);
nor U11267 (N_11267,N_11179,N_11128);
xnor U11268 (N_11268,N_11123,N_11119);
nor U11269 (N_11269,N_11175,N_11103);
xnor U11270 (N_11270,N_11144,N_11187);
or U11271 (N_11271,N_11152,N_11140);
and U11272 (N_11272,N_11173,N_11106);
nand U11273 (N_11273,N_11135,N_11208);
nor U11274 (N_11274,N_11127,N_11118);
nor U11275 (N_11275,N_11220,N_11192);
and U11276 (N_11276,N_11157,N_11182);
nor U11277 (N_11277,N_11242,N_11115);
nor U11278 (N_11278,N_11223,N_11111);
nor U11279 (N_11279,N_11139,N_11238);
and U11280 (N_11280,N_11241,N_11142);
xor U11281 (N_11281,N_11102,N_11159);
and U11282 (N_11282,N_11134,N_11164);
and U11283 (N_11283,N_11141,N_11245);
xor U11284 (N_11284,N_11230,N_11171);
and U11285 (N_11285,N_11219,N_11177);
nor U11286 (N_11286,N_11204,N_11137);
or U11287 (N_11287,N_11168,N_11112);
and U11288 (N_11288,N_11113,N_11150);
and U11289 (N_11289,N_11122,N_11172);
or U11290 (N_11290,N_11184,N_11224);
xor U11291 (N_11291,N_11186,N_11105);
and U11292 (N_11292,N_11158,N_11153);
nor U11293 (N_11293,N_11183,N_11110);
or U11294 (N_11294,N_11188,N_11226);
nand U11295 (N_11295,N_11194,N_11240);
xor U11296 (N_11296,N_11160,N_11228);
xnor U11297 (N_11297,N_11178,N_11248);
nand U11298 (N_11298,N_11181,N_11114);
and U11299 (N_11299,N_11229,N_11143);
and U11300 (N_11300,N_11233,N_11214);
nor U11301 (N_11301,N_11209,N_11195);
and U11302 (N_11302,N_11222,N_11244);
nand U11303 (N_11303,N_11232,N_11132);
nand U11304 (N_11304,N_11225,N_11218);
or U11305 (N_11305,N_11190,N_11149);
nor U11306 (N_11306,N_11235,N_11205);
nand U11307 (N_11307,N_11203,N_11121);
or U11308 (N_11308,N_11116,N_11165);
and U11309 (N_11309,N_11136,N_11162);
and U11310 (N_11310,N_11154,N_11247);
xnor U11311 (N_11311,N_11109,N_11236);
and U11312 (N_11312,N_11212,N_11104);
or U11313 (N_11313,N_11125,N_11193);
nand U11314 (N_11314,N_11246,N_11215);
nor U11315 (N_11315,N_11138,N_11191);
nand U11316 (N_11316,N_11243,N_11151);
or U11317 (N_11317,N_11227,N_11130);
or U11318 (N_11318,N_11202,N_11206);
xnor U11319 (N_11319,N_11169,N_11101);
xor U11320 (N_11320,N_11189,N_11120);
and U11321 (N_11321,N_11170,N_11196);
xor U11322 (N_11322,N_11126,N_11145);
nand U11323 (N_11323,N_11237,N_11213);
xor U11324 (N_11324,N_11207,N_11200);
xnor U11325 (N_11325,N_11172,N_11137);
nor U11326 (N_11326,N_11117,N_11174);
or U11327 (N_11327,N_11162,N_11113);
nor U11328 (N_11328,N_11116,N_11226);
or U11329 (N_11329,N_11214,N_11141);
and U11330 (N_11330,N_11121,N_11164);
nand U11331 (N_11331,N_11216,N_11220);
nand U11332 (N_11332,N_11229,N_11220);
nand U11333 (N_11333,N_11120,N_11245);
nand U11334 (N_11334,N_11125,N_11202);
or U11335 (N_11335,N_11203,N_11235);
xor U11336 (N_11336,N_11215,N_11184);
or U11337 (N_11337,N_11244,N_11118);
nor U11338 (N_11338,N_11213,N_11191);
and U11339 (N_11339,N_11119,N_11177);
nand U11340 (N_11340,N_11199,N_11214);
or U11341 (N_11341,N_11149,N_11209);
nand U11342 (N_11342,N_11179,N_11151);
nor U11343 (N_11343,N_11236,N_11225);
nand U11344 (N_11344,N_11169,N_11124);
nand U11345 (N_11345,N_11245,N_11169);
or U11346 (N_11346,N_11204,N_11241);
or U11347 (N_11347,N_11101,N_11153);
xor U11348 (N_11348,N_11246,N_11222);
xnor U11349 (N_11349,N_11188,N_11155);
nor U11350 (N_11350,N_11119,N_11147);
nor U11351 (N_11351,N_11214,N_11170);
and U11352 (N_11352,N_11196,N_11148);
and U11353 (N_11353,N_11152,N_11188);
or U11354 (N_11354,N_11127,N_11165);
and U11355 (N_11355,N_11140,N_11101);
nor U11356 (N_11356,N_11130,N_11189);
nor U11357 (N_11357,N_11139,N_11219);
nor U11358 (N_11358,N_11112,N_11107);
and U11359 (N_11359,N_11164,N_11113);
nor U11360 (N_11360,N_11248,N_11239);
nand U11361 (N_11361,N_11115,N_11236);
nand U11362 (N_11362,N_11137,N_11160);
or U11363 (N_11363,N_11196,N_11110);
or U11364 (N_11364,N_11147,N_11211);
xnor U11365 (N_11365,N_11244,N_11126);
and U11366 (N_11366,N_11146,N_11120);
xor U11367 (N_11367,N_11114,N_11245);
xnor U11368 (N_11368,N_11156,N_11164);
or U11369 (N_11369,N_11201,N_11152);
nand U11370 (N_11370,N_11247,N_11164);
nand U11371 (N_11371,N_11212,N_11211);
nand U11372 (N_11372,N_11189,N_11127);
xor U11373 (N_11373,N_11150,N_11210);
xnor U11374 (N_11374,N_11111,N_11197);
nand U11375 (N_11375,N_11150,N_11129);
or U11376 (N_11376,N_11119,N_11197);
or U11377 (N_11377,N_11169,N_11138);
xor U11378 (N_11378,N_11237,N_11236);
nor U11379 (N_11379,N_11201,N_11165);
and U11380 (N_11380,N_11217,N_11166);
nand U11381 (N_11381,N_11249,N_11117);
xor U11382 (N_11382,N_11238,N_11120);
nand U11383 (N_11383,N_11204,N_11120);
nor U11384 (N_11384,N_11109,N_11184);
or U11385 (N_11385,N_11114,N_11207);
or U11386 (N_11386,N_11182,N_11166);
nor U11387 (N_11387,N_11193,N_11190);
nand U11388 (N_11388,N_11162,N_11238);
xnor U11389 (N_11389,N_11203,N_11239);
nand U11390 (N_11390,N_11187,N_11213);
nand U11391 (N_11391,N_11239,N_11192);
nor U11392 (N_11392,N_11231,N_11219);
nor U11393 (N_11393,N_11208,N_11125);
or U11394 (N_11394,N_11135,N_11153);
or U11395 (N_11395,N_11123,N_11112);
nand U11396 (N_11396,N_11219,N_11213);
and U11397 (N_11397,N_11151,N_11229);
xnor U11398 (N_11398,N_11232,N_11233);
nand U11399 (N_11399,N_11199,N_11145);
nand U11400 (N_11400,N_11342,N_11333);
nand U11401 (N_11401,N_11330,N_11291);
xnor U11402 (N_11402,N_11263,N_11325);
nand U11403 (N_11403,N_11279,N_11345);
nand U11404 (N_11404,N_11281,N_11394);
nand U11405 (N_11405,N_11332,N_11354);
nand U11406 (N_11406,N_11328,N_11377);
nand U11407 (N_11407,N_11310,N_11397);
nand U11408 (N_11408,N_11275,N_11372);
nand U11409 (N_11409,N_11350,N_11259);
nand U11410 (N_11410,N_11351,N_11305);
and U11411 (N_11411,N_11341,N_11296);
nand U11412 (N_11412,N_11361,N_11321);
xor U11413 (N_11413,N_11356,N_11260);
and U11414 (N_11414,N_11368,N_11312);
nand U11415 (N_11415,N_11274,N_11300);
nor U11416 (N_11416,N_11386,N_11339);
xor U11417 (N_11417,N_11393,N_11271);
or U11418 (N_11418,N_11252,N_11384);
nor U11419 (N_11419,N_11284,N_11264);
and U11420 (N_11420,N_11290,N_11313);
nor U11421 (N_11421,N_11383,N_11396);
xor U11422 (N_11422,N_11295,N_11348);
nor U11423 (N_11423,N_11278,N_11374);
and U11424 (N_11424,N_11331,N_11294);
and U11425 (N_11425,N_11380,N_11307);
nor U11426 (N_11426,N_11316,N_11326);
or U11427 (N_11427,N_11327,N_11317);
xnor U11428 (N_11428,N_11304,N_11258);
and U11429 (N_11429,N_11262,N_11349);
xnor U11430 (N_11430,N_11297,N_11253);
xor U11431 (N_11431,N_11254,N_11390);
and U11432 (N_11432,N_11324,N_11309);
xor U11433 (N_11433,N_11335,N_11385);
nand U11434 (N_11434,N_11399,N_11355);
and U11435 (N_11435,N_11255,N_11378);
nor U11436 (N_11436,N_11314,N_11251);
and U11437 (N_11437,N_11299,N_11315);
nor U11438 (N_11438,N_11273,N_11371);
and U11439 (N_11439,N_11343,N_11357);
nor U11440 (N_11440,N_11398,N_11306);
xnor U11441 (N_11441,N_11344,N_11270);
or U11442 (N_11442,N_11347,N_11308);
and U11443 (N_11443,N_11319,N_11340);
nor U11444 (N_11444,N_11375,N_11302);
nor U11445 (N_11445,N_11277,N_11250);
xnor U11446 (N_11446,N_11266,N_11322);
or U11447 (N_11447,N_11318,N_11379);
nor U11448 (N_11448,N_11293,N_11288);
xor U11449 (N_11449,N_11329,N_11320);
or U11450 (N_11450,N_11387,N_11336);
or U11451 (N_11451,N_11257,N_11298);
or U11452 (N_11452,N_11352,N_11280);
nor U11453 (N_11453,N_11272,N_11311);
xor U11454 (N_11454,N_11365,N_11334);
nor U11455 (N_11455,N_11289,N_11287);
nand U11456 (N_11456,N_11268,N_11338);
or U11457 (N_11457,N_11367,N_11276);
nand U11458 (N_11458,N_11285,N_11358);
nand U11459 (N_11459,N_11256,N_11360);
nor U11460 (N_11460,N_11376,N_11267);
nor U11461 (N_11461,N_11301,N_11389);
or U11462 (N_11462,N_11337,N_11292);
nor U11463 (N_11463,N_11282,N_11373);
and U11464 (N_11464,N_11346,N_11370);
xnor U11465 (N_11465,N_11363,N_11391);
or U11466 (N_11466,N_11353,N_11382);
and U11467 (N_11467,N_11392,N_11362);
and U11468 (N_11468,N_11286,N_11283);
xnor U11469 (N_11469,N_11323,N_11269);
or U11470 (N_11470,N_11265,N_11364);
xnor U11471 (N_11471,N_11359,N_11366);
nor U11472 (N_11472,N_11261,N_11395);
nand U11473 (N_11473,N_11369,N_11303);
xnor U11474 (N_11474,N_11381,N_11388);
nor U11475 (N_11475,N_11351,N_11361);
nand U11476 (N_11476,N_11350,N_11363);
or U11477 (N_11477,N_11281,N_11374);
nor U11478 (N_11478,N_11359,N_11340);
nand U11479 (N_11479,N_11293,N_11284);
nor U11480 (N_11480,N_11315,N_11378);
nand U11481 (N_11481,N_11315,N_11258);
xor U11482 (N_11482,N_11397,N_11320);
xnor U11483 (N_11483,N_11375,N_11360);
or U11484 (N_11484,N_11273,N_11390);
xor U11485 (N_11485,N_11327,N_11356);
and U11486 (N_11486,N_11324,N_11280);
xnor U11487 (N_11487,N_11283,N_11293);
nor U11488 (N_11488,N_11277,N_11292);
nand U11489 (N_11489,N_11356,N_11373);
and U11490 (N_11490,N_11305,N_11294);
nand U11491 (N_11491,N_11356,N_11259);
or U11492 (N_11492,N_11334,N_11253);
and U11493 (N_11493,N_11326,N_11263);
xnor U11494 (N_11494,N_11369,N_11351);
nand U11495 (N_11495,N_11273,N_11320);
nor U11496 (N_11496,N_11346,N_11335);
nor U11497 (N_11497,N_11272,N_11396);
or U11498 (N_11498,N_11360,N_11295);
nor U11499 (N_11499,N_11337,N_11333);
xnor U11500 (N_11500,N_11303,N_11257);
xor U11501 (N_11501,N_11310,N_11304);
nor U11502 (N_11502,N_11291,N_11320);
nor U11503 (N_11503,N_11314,N_11299);
xnor U11504 (N_11504,N_11321,N_11318);
nand U11505 (N_11505,N_11289,N_11283);
xnor U11506 (N_11506,N_11275,N_11276);
nor U11507 (N_11507,N_11361,N_11251);
nand U11508 (N_11508,N_11276,N_11385);
nand U11509 (N_11509,N_11340,N_11321);
nor U11510 (N_11510,N_11334,N_11283);
or U11511 (N_11511,N_11293,N_11377);
or U11512 (N_11512,N_11335,N_11294);
and U11513 (N_11513,N_11252,N_11262);
or U11514 (N_11514,N_11274,N_11316);
and U11515 (N_11515,N_11253,N_11393);
nor U11516 (N_11516,N_11303,N_11358);
nand U11517 (N_11517,N_11330,N_11273);
and U11518 (N_11518,N_11276,N_11383);
nor U11519 (N_11519,N_11390,N_11358);
and U11520 (N_11520,N_11307,N_11324);
or U11521 (N_11521,N_11329,N_11312);
xor U11522 (N_11522,N_11279,N_11276);
xor U11523 (N_11523,N_11397,N_11313);
xor U11524 (N_11524,N_11285,N_11324);
nand U11525 (N_11525,N_11268,N_11324);
or U11526 (N_11526,N_11386,N_11253);
nor U11527 (N_11527,N_11286,N_11348);
or U11528 (N_11528,N_11278,N_11372);
nor U11529 (N_11529,N_11315,N_11298);
and U11530 (N_11530,N_11315,N_11273);
or U11531 (N_11531,N_11289,N_11325);
or U11532 (N_11532,N_11389,N_11315);
or U11533 (N_11533,N_11360,N_11259);
nand U11534 (N_11534,N_11258,N_11277);
or U11535 (N_11535,N_11297,N_11384);
or U11536 (N_11536,N_11268,N_11270);
and U11537 (N_11537,N_11258,N_11281);
nand U11538 (N_11538,N_11370,N_11379);
or U11539 (N_11539,N_11283,N_11331);
or U11540 (N_11540,N_11281,N_11260);
and U11541 (N_11541,N_11263,N_11304);
xor U11542 (N_11542,N_11307,N_11362);
and U11543 (N_11543,N_11274,N_11280);
or U11544 (N_11544,N_11391,N_11290);
nand U11545 (N_11545,N_11254,N_11344);
and U11546 (N_11546,N_11377,N_11334);
nand U11547 (N_11547,N_11340,N_11373);
nand U11548 (N_11548,N_11264,N_11259);
nor U11549 (N_11549,N_11324,N_11317);
or U11550 (N_11550,N_11489,N_11537);
xor U11551 (N_11551,N_11479,N_11503);
nand U11552 (N_11552,N_11407,N_11443);
nor U11553 (N_11553,N_11510,N_11437);
nand U11554 (N_11554,N_11487,N_11473);
nand U11555 (N_11555,N_11468,N_11496);
and U11556 (N_11556,N_11416,N_11514);
nor U11557 (N_11557,N_11474,N_11475);
and U11558 (N_11558,N_11452,N_11485);
nand U11559 (N_11559,N_11449,N_11453);
or U11560 (N_11560,N_11448,N_11430);
and U11561 (N_11561,N_11547,N_11492);
xor U11562 (N_11562,N_11436,N_11435);
or U11563 (N_11563,N_11450,N_11490);
xor U11564 (N_11564,N_11405,N_11446);
xor U11565 (N_11565,N_11497,N_11543);
and U11566 (N_11566,N_11458,N_11427);
nor U11567 (N_11567,N_11517,N_11403);
nor U11568 (N_11568,N_11419,N_11418);
nand U11569 (N_11569,N_11525,N_11549);
nor U11570 (N_11570,N_11417,N_11522);
nor U11571 (N_11571,N_11493,N_11513);
and U11572 (N_11572,N_11457,N_11494);
nor U11573 (N_11573,N_11472,N_11504);
and U11574 (N_11574,N_11433,N_11544);
and U11575 (N_11575,N_11536,N_11486);
or U11576 (N_11576,N_11455,N_11546);
xor U11577 (N_11577,N_11477,N_11515);
xor U11578 (N_11578,N_11509,N_11422);
nand U11579 (N_11579,N_11439,N_11408);
xor U11580 (N_11580,N_11415,N_11476);
nor U11581 (N_11581,N_11548,N_11523);
nor U11582 (N_11582,N_11482,N_11481);
xor U11583 (N_11583,N_11429,N_11451);
and U11584 (N_11584,N_11532,N_11438);
and U11585 (N_11585,N_11465,N_11484);
nand U11586 (N_11586,N_11542,N_11411);
nor U11587 (N_11587,N_11441,N_11471);
nand U11588 (N_11588,N_11464,N_11512);
xnor U11589 (N_11589,N_11483,N_11404);
nor U11590 (N_11590,N_11432,N_11533);
nand U11591 (N_11591,N_11425,N_11420);
or U11592 (N_11592,N_11531,N_11511);
or U11593 (N_11593,N_11456,N_11467);
or U11594 (N_11594,N_11460,N_11488);
or U11595 (N_11595,N_11502,N_11545);
xnor U11596 (N_11596,N_11461,N_11501);
and U11597 (N_11597,N_11541,N_11440);
nand U11598 (N_11598,N_11413,N_11534);
xnor U11599 (N_11599,N_11466,N_11530);
nor U11600 (N_11600,N_11538,N_11499);
nor U11601 (N_11601,N_11402,N_11535);
nor U11602 (N_11602,N_11521,N_11507);
xnor U11603 (N_11603,N_11423,N_11414);
nand U11604 (N_11604,N_11498,N_11406);
xor U11605 (N_11605,N_11428,N_11444);
nand U11606 (N_11606,N_11478,N_11463);
or U11607 (N_11607,N_11528,N_11410);
and U11608 (N_11608,N_11500,N_11445);
and U11609 (N_11609,N_11442,N_11400);
nor U11610 (N_11610,N_11401,N_11470);
nor U11611 (N_11611,N_11540,N_11469);
xor U11612 (N_11612,N_11539,N_11516);
and U11613 (N_11613,N_11505,N_11506);
xor U11614 (N_11614,N_11519,N_11412);
nor U11615 (N_11615,N_11480,N_11529);
nor U11616 (N_11616,N_11526,N_11518);
nand U11617 (N_11617,N_11454,N_11434);
xor U11618 (N_11618,N_11520,N_11431);
nor U11619 (N_11619,N_11426,N_11524);
xor U11620 (N_11620,N_11462,N_11447);
nand U11621 (N_11621,N_11459,N_11495);
nand U11622 (N_11622,N_11421,N_11527);
and U11623 (N_11623,N_11424,N_11508);
and U11624 (N_11624,N_11491,N_11409);
or U11625 (N_11625,N_11482,N_11401);
xnor U11626 (N_11626,N_11497,N_11498);
nand U11627 (N_11627,N_11429,N_11530);
nor U11628 (N_11628,N_11456,N_11419);
xnor U11629 (N_11629,N_11471,N_11409);
nand U11630 (N_11630,N_11524,N_11443);
and U11631 (N_11631,N_11448,N_11439);
nor U11632 (N_11632,N_11515,N_11406);
nand U11633 (N_11633,N_11438,N_11499);
and U11634 (N_11634,N_11436,N_11461);
xor U11635 (N_11635,N_11461,N_11487);
nor U11636 (N_11636,N_11544,N_11476);
and U11637 (N_11637,N_11446,N_11425);
and U11638 (N_11638,N_11429,N_11508);
xor U11639 (N_11639,N_11509,N_11508);
xnor U11640 (N_11640,N_11468,N_11490);
nand U11641 (N_11641,N_11464,N_11461);
nand U11642 (N_11642,N_11410,N_11424);
and U11643 (N_11643,N_11412,N_11469);
and U11644 (N_11644,N_11456,N_11504);
nor U11645 (N_11645,N_11440,N_11435);
xor U11646 (N_11646,N_11410,N_11508);
xnor U11647 (N_11647,N_11536,N_11471);
or U11648 (N_11648,N_11400,N_11545);
nand U11649 (N_11649,N_11459,N_11433);
nand U11650 (N_11650,N_11421,N_11533);
xnor U11651 (N_11651,N_11490,N_11482);
nand U11652 (N_11652,N_11540,N_11439);
nand U11653 (N_11653,N_11426,N_11520);
and U11654 (N_11654,N_11470,N_11440);
nand U11655 (N_11655,N_11537,N_11419);
and U11656 (N_11656,N_11463,N_11439);
or U11657 (N_11657,N_11400,N_11542);
xnor U11658 (N_11658,N_11499,N_11470);
and U11659 (N_11659,N_11417,N_11528);
or U11660 (N_11660,N_11523,N_11403);
and U11661 (N_11661,N_11470,N_11439);
xnor U11662 (N_11662,N_11545,N_11512);
or U11663 (N_11663,N_11462,N_11520);
nand U11664 (N_11664,N_11453,N_11504);
nand U11665 (N_11665,N_11492,N_11416);
nand U11666 (N_11666,N_11470,N_11549);
or U11667 (N_11667,N_11443,N_11525);
or U11668 (N_11668,N_11415,N_11543);
and U11669 (N_11669,N_11469,N_11506);
and U11670 (N_11670,N_11481,N_11478);
xor U11671 (N_11671,N_11474,N_11515);
nor U11672 (N_11672,N_11518,N_11469);
and U11673 (N_11673,N_11439,N_11498);
and U11674 (N_11674,N_11485,N_11522);
or U11675 (N_11675,N_11452,N_11507);
nor U11676 (N_11676,N_11488,N_11496);
and U11677 (N_11677,N_11412,N_11492);
xnor U11678 (N_11678,N_11517,N_11414);
nor U11679 (N_11679,N_11529,N_11418);
nand U11680 (N_11680,N_11434,N_11409);
nand U11681 (N_11681,N_11453,N_11434);
nor U11682 (N_11682,N_11525,N_11427);
nor U11683 (N_11683,N_11422,N_11459);
xnor U11684 (N_11684,N_11460,N_11445);
or U11685 (N_11685,N_11517,N_11489);
and U11686 (N_11686,N_11517,N_11484);
nor U11687 (N_11687,N_11411,N_11403);
nand U11688 (N_11688,N_11465,N_11413);
xor U11689 (N_11689,N_11519,N_11541);
nor U11690 (N_11690,N_11441,N_11446);
nand U11691 (N_11691,N_11527,N_11423);
or U11692 (N_11692,N_11549,N_11462);
nand U11693 (N_11693,N_11524,N_11464);
nor U11694 (N_11694,N_11487,N_11442);
or U11695 (N_11695,N_11549,N_11512);
or U11696 (N_11696,N_11508,N_11428);
nor U11697 (N_11697,N_11545,N_11513);
or U11698 (N_11698,N_11471,N_11524);
nand U11699 (N_11699,N_11438,N_11411);
or U11700 (N_11700,N_11550,N_11627);
or U11701 (N_11701,N_11659,N_11689);
nand U11702 (N_11702,N_11555,N_11693);
and U11703 (N_11703,N_11600,N_11612);
nand U11704 (N_11704,N_11674,N_11619);
or U11705 (N_11705,N_11556,N_11561);
and U11706 (N_11706,N_11587,N_11610);
or U11707 (N_11707,N_11684,N_11665);
nand U11708 (N_11708,N_11590,N_11598);
or U11709 (N_11709,N_11569,N_11616);
xnor U11710 (N_11710,N_11611,N_11573);
or U11711 (N_11711,N_11681,N_11558);
xor U11712 (N_11712,N_11680,N_11635);
nor U11713 (N_11713,N_11634,N_11622);
and U11714 (N_11714,N_11579,N_11554);
xnor U11715 (N_11715,N_11588,N_11669);
nor U11716 (N_11716,N_11652,N_11583);
nand U11717 (N_11717,N_11624,N_11581);
xor U11718 (N_11718,N_11575,N_11676);
or U11719 (N_11719,N_11553,N_11636);
and U11720 (N_11720,N_11577,N_11586);
or U11721 (N_11721,N_11580,N_11621);
nor U11722 (N_11722,N_11566,N_11551);
nor U11723 (N_11723,N_11603,N_11685);
nor U11724 (N_11724,N_11618,N_11668);
xor U11725 (N_11725,N_11691,N_11648);
and U11726 (N_11726,N_11653,N_11585);
nor U11727 (N_11727,N_11678,N_11609);
or U11728 (N_11728,N_11562,N_11655);
xor U11729 (N_11729,N_11630,N_11552);
and U11730 (N_11730,N_11682,N_11620);
nand U11731 (N_11731,N_11660,N_11602);
nor U11732 (N_11732,N_11658,N_11628);
nand U11733 (N_11733,N_11576,N_11560);
nor U11734 (N_11734,N_11606,N_11613);
and U11735 (N_11735,N_11657,N_11557);
and U11736 (N_11736,N_11565,N_11645);
nand U11737 (N_11737,N_11688,N_11671);
nor U11738 (N_11738,N_11574,N_11650);
nor U11739 (N_11739,N_11699,N_11683);
nor U11740 (N_11740,N_11605,N_11638);
or U11741 (N_11741,N_11582,N_11559);
nor U11742 (N_11742,N_11568,N_11649);
and U11743 (N_11743,N_11608,N_11564);
or U11744 (N_11744,N_11595,N_11604);
or U11745 (N_11745,N_11643,N_11696);
or U11746 (N_11746,N_11623,N_11642);
xnor U11747 (N_11747,N_11578,N_11673);
xor U11748 (N_11748,N_11695,N_11632);
or U11749 (N_11749,N_11571,N_11690);
nor U11750 (N_11750,N_11687,N_11640);
nand U11751 (N_11751,N_11654,N_11692);
xor U11752 (N_11752,N_11629,N_11679);
xnor U11753 (N_11753,N_11601,N_11641);
nand U11754 (N_11754,N_11675,N_11617);
and U11755 (N_11755,N_11666,N_11597);
or U11756 (N_11756,N_11662,N_11596);
xor U11757 (N_11757,N_11591,N_11639);
xor U11758 (N_11758,N_11651,N_11594);
or U11759 (N_11759,N_11607,N_11589);
nor U11760 (N_11760,N_11572,N_11656);
and U11761 (N_11761,N_11625,N_11599);
or U11762 (N_11762,N_11631,N_11646);
nand U11763 (N_11763,N_11697,N_11570);
nand U11764 (N_11764,N_11664,N_11567);
nor U11765 (N_11765,N_11670,N_11633);
nor U11766 (N_11766,N_11694,N_11677);
nand U11767 (N_11767,N_11584,N_11614);
nor U11768 (N_11768,N_11647,N_11593);
nand U11769 (N_11769,N_11663,N_11672);
and U11770 (N_11770,N_11698,N_11615);
or U11771 (N_11771,N_11661,N_11644);
and U11772 (N_11772,N_11667,N_11592);
nor U11773 (N_11773,N_11686,N_11626);
nor U11774 (N_11774,N_11637,N_11563);
nor U11775 (N_11775,N_11612,N_11687);
nand U11776 (N_11776,N_11656,N_11686);
nand U11777 (N_11777,N_11585,N_11567);
xor U11778 (N_11778,N_11690,N_11696);
nor U11779 (N_11779,N_11620,N_11671);
nand U11780 (N_11780,N_11616,N_11674);
and U11781 (N_11781,N_11688,N_11568);
and U11782 (N_11782,N_11697,N_11619);
or U11783 (N_11783,N_11634,N_11672);
and U11784 (N_11784,N_11668,N_11672);
nor U11785 (N_11785,N_11651,N_11690);
nand U11786 (N_11786,N_11599,N_11593);
and U11787 (N_11787,N_11584,N_11586);
xor U11788 (N_11788,N_11679,N_11672);
nor U11789 (N_11789,N_11608,N_11557);
or U11790 (N_11790,N_11655,N_11681);
nand U11791 (N_11791,N_11578,N_11644);
xor U11792 (N_11792,N_11686,N_11689);
nand U11793 (N_11793,N_11624,N_11674);
xor U11794 (N_11794,N_11566,N_11603);
nand U11795 (N_11795,N_11579,N_11575);
xor U11796 (N_11796,N_11697,N_11661);
or U11797 (N_11797,N_11667,N_11656);
nand U11798 (N_11798,N_11572,N_11653);
nand U11799 (N_11799,N_11687,N_11668);
or U11800 (N_11800,N_11600,N_11665);
nor U11801 (N_11801,N_11683,N_11668);
nand U11802 (N_11802,N_11570,N_11566);
or U11803 (N_11803,N_11665,N_11689);
or U11804 (N_11804,N_11635,N_11586);
nand U11805 (N_11805,N_11570,N_11575);
nand U11806 (N_11806,N_11663,N_11578);
and U11807 (N_11807,N_11672,N_11585);
and U11808 (N_11808,N_11689,N_11658);
and U11809 (N_11809,N_11656,N_11644);
and U11810 (N_11810,N_11641,N_11673);
nor U11811 (N_11811,N_11653,N_11690);
xor U11812 (N_11812,N_11569,N_11641);
xor U11813 (N_11813,N_11643,N_11616);
or U11814 (N_11814,N_11653,N_11697);
nor U11815 (N_11815,N_11674,N_11620);
and U11816 (N_11816,N_11561,N_11647);
xnor U11817 (N_11817,N_11551,N_11560);
or U11818 (N_11818,N_11603,N_11653);
or U11819 (N_11819,N_11550,N_11570);
and U11820 (N_11820,N_11660,N_11694);
nor U11821 (N_11821,N_11573,N_11689);
or U11822 (N_11822,N_11689,N_11671);
nand U11823 (N_11823,N_11672,N_11698);
nor U11824 (N_11824,N_11630,N_11585);
and U11825 (N_11825,N_11665,N_11579);
or U11826 (N_11826,N_11652,N_11685);
or U11827 (N_11827,N_11571,N_11589);
or U11828 (N_11828,N_11600,N_11664);
nor U11829 (N_11829,N_11628,N_11571);
nor U11830 (N_11830,N_11569,N_11581);
nor U11831 (N_11831,N_11673,N_11579);
nor U11832 (N_11832,N_11670,N_11647);
or U11833 (N_11833,N_11698,N_11685);
nor U11834 (N_11834,N_11642,N_11550);
and U11835 (N_11835,N_11590,N_11684);
xnor U11836 (N_11836,N_11683,N_11567);
nor U11837 (N_11837,N_11651,N_11621);
or U11838 (N_11838,N_11644,N_11643);
or U11839 (N_11839,N_11628,N_11559);
nand U11840 (N_11840,N_11689,N_11569);
xor U11841 (N_11841,N_11680,N_11587);
or U11842 (N_11842,N_11695,N_11600);
nand U11843 (N_11843,N_11661,N_11628);
and U11844 (N_11844,N_11601,N_11634);
or U11845 (N_11845,N_11622,N_11567);
and U11846 (N_11846,N_11655,N_11612);
and U11847 (N_11847,N_11684,N_11591);
xnor U11848 (N_11848,N_11639,N_11621);
xor U11849 (N_11849,N_11607,N_11558);
nor U11850 (N_11850,N_11737,N_11824);
nand U11851 (N_11851,N_11842,N_11712);
or U11852 (N_11852,N_11744,N_11801);
nor U11853 (N_11853,N_11769,N_11732);
xor U11854 (N_11854,N_11826,N_11753);
nor U11855 (N_11855,N_11713,N_11798);
xor U11856 (N_11856,N_11763,N_11849);
nand U11857 (N_11857,N_11750,N_11802);
and U11858 (N_11858,N_11707,N_11848);
nor U11859 (N_11859,N_11803,N_11723);
xor U11860 (N_11860,N_11799,N_11715);
xnor U11861 (N_11861,N_11749,N_11765);
and U11862 (N_11862,N_11787,N_11718);
or U11863 (N_11863,N_11760,N_11836);
and U11864 (N_11864,N_11743,N_11831);
nor U11865 (N_11865,N_11810,N_11817);
or U11866 (N_11866,N_11811,N_11736);
or U11867 (N_11867,N_11785,N_11825);
nand U11868 (N_11868,N_11812,N_11757);
nor U11869 (N_11869,N_11726,N_11729);
xnor U11870 (N_11870,N_11703,N_11704);
nor U11871 (N_11871,N_11780,N_11739);
and U11872 (N_11872,N_11708,N_11700);
or U11873 (N_11873,N_11772,N_11705);
nor U11874 (N_11874,N_11746,N_11791);
nand U11875 (N_11875,N_11773,N_11795);
xnor U11876 (N_11876,N_11834,N_11748);
and U11877 (N_11877,N_11827,N_11719);
nor U11878 (N_11878,N_11820,N_11792);
nor U11879 (N_11879,N_11762,N_11741);
and U11880 (N_11880,N_11828,N_11821);
nor U11881 (N_11881,N_11710,N_11829);
xor U11882 (N_11882,N_11788,N_11756);
nand U11883 (N_11883,N_11776,N_11786);
nor U11884 (N_11884,N_11844,N_11815);
nand U11885 (N_11885,N_11764,N_11774);
or U11886 (N_11886,N_11835,N_11754);
xnor U11887 (N_11887,N_11845,N_11752);
nand U11888 (N_11888,N_11793,N_11777);
nor U11889 (N_11889,N_11721,N_11728);
or U11890 (N_11890,N_11809,N_11755);
or U11891 (N_11891,N_11783,N_11782);
and U11892 (N_11892,N_11709,N_11740);
and U11893 (N_11893,N_11758,N_11790);
and U11894 (N_11894,N_11804,N_11843);
nand U11895 (N_11895,N_11738,N_11701);
nand U11896 (N_11896,N_11784,N_11747);
and U11897 (N_11897,N_11781,N_11720);
xnor U11898 (N_11898,N_11822,N_11800);
xnor U11899 (N_11899,N_11823,N_11805);
nor U11900 (N_11900,N_11761,N_11794);
and U11901 (N_11901,N_11816,N_11711);
or U11902 (N_11902,N_11806,N_11813);
xor U11903 (N_11903,N_11819,N_11797);
nor U11904 (N_11904,N_11847,N_11789);
and U11905 (N_11905,N_11775,N_11742);
xnor U11906 (N_11906,N_11837,N_11839);
nor U11907 (N_11907,N_11796,N_11734);
or U11908 (N_11908,N_11818,N_11735);
nor U11909 (N_11909,N_11832,N_11770);
xor U11910 (N_11910,N_11833,N_11838);
and U11911 (N_11911,N_11722,N_11731);
xor U11912 (N_11912,N_11733,N_11751);
and U11913 (N_11913,N_11814,N_11807);
nand U11914 (N_11914,N_11716,N_11768);
nor U11915 (N_11915,N_11702,N_11724);
nand U11916 (N_11916,N_11846,N_11766);
xnor U11917 (N_11917,N_11841,N_11779);
and U11918 (N_11918,N_11745,N_11830);
or U11919 (N_11919,N_11771,N_11778);
nor U11920 (N_11920,N_11706,N_11808);
nand U11921 (N_11921,N_11725,N_11714);
nand U11922 (N_11922,N_11727,N_11730);
or U11923 (N_11923,N_11767,N_11759);
or U11924 (N_11924,N_11840,N_11717);
nand U11925 (N_11925,N_11842,N_11803);
and U11926 (N_11926,N_11749,N_11798);
nand U11927 (N_11927,N_11708,N_11788);
nand U11928 (N_11928,N_11725,N_11719);
nand U11929 (N_11929,N_11746,N_11828);
xor U11930 (N_11930,N_11848,N_11776);
nand U11931 (N_11931,N_11794,N_11740);
nand U11932 (N_11932,N_11729,N_11801);
nand U11933 (N_11933,N_11813,N_11740);
xnor U11934 (N_11934,N_11737,N_11709);
and U11935 (N_11935,N_11834,N_11846);
xor U11936 (N_11936,N_11827,N_11787);
or U11937 (N_11937,N_11739,N_11808);
nand U11938 (N_11938,N_11791,N_11847);
or U11939 (N_11939,N_11781,N_11746);
nand U11940 (N_11940,N_11831,N_11703);
nand U11941 (N_11941,N_11833,N_11751);
or U11942 (N_11942,N_11721,N_11735);
or U11943 (N_11943,N_11830,N_11789);
nor U11944 (N_11944,N_11843,N_11705);
nand U11945 (N_11945,N_11723,N_11755);
xor U11946 (N_11946,N_11800,N_11752);
xor U11947 (N_11947,N_11715,N_11812);
nand U11948 (N_11948,N_11715,N_11772);
xor U11949 (N_11949,N_11831,N_11720);
and U11950 (N_11950,N_11837,N_11848);
xor U11951 (N_11951,N_11738,N_11837);
or U11952 (N_11952,N_11827,N_11756);
xor U11953 (N_11953,N_11736,N_11784);
and U11954 (N_11954,N_11799,N_11843);
or U11955 (N_11955,N_11748,N_11722);
and U11956 (N_11956,N_11708,N_11779);
and U11957 (N_11957,N_11836,N_11827);
nand U11958 (N_11958,N_11815,N_11818);
nor U11959 (N_11959,N_11709,N_11708);
and U11960 (N_11960,N_11760,N_11791);
or U11961 (N_11961,N_11766,N_11842);
and U11962 (N_11962,N_11700,N_11825);
or U11963 (N_11963,N_11712,N_11766);
or U11964 (N_11964,N_11719,N_11759);
nand U11965 (N_11965,N_11766,N_11708);
nand U11966 (N_11966,N_11789,N_11808);
or U11967 (N_11967,N_11715,N_11733);
nor U11968 (N_11968,N_11804,N_11815);
nor U11969 (N_11969,N_11772,N_11753);
or U11970 (N_11970,N_11738,N_11732);
nor U11971 (N_11971,N_11811,N_11818);
and U11972 (N_11972,N_11787,N_11732);
xor U11973 (N_11973,N_11781,N_11814);
nand U11974 (N_11974,N_11735,N_11822);
nor U11975 (N_11975,N_11723,N_11775);
and U11976 (N_11976,N_11754,N_11728);
nand U11977 (N_11977,N_11726,N_11789);
nand U11978 (N_11978,N_11835,N_11766);
or U11979 (N_11979,N_11847,N_11842);
and U11980 (N_11980,N_11822,N_11813);
and U11981 (N_11981,N_11762,N_11797);
and U11982 (N_11982,N_11791,N_11761);
nor U11983 (N_11983,N_11812,N_11808);
or U11984 (N_11984,N_11766,N_11816);
nand U11985 (N_11985,N_11749,N_11774);
nand U11986 (N_11986,N_11720,N_11742);
and U11987 (N_11987,N_11827,N_11819);
and U11988 (N_11988,N_11711,N_11744);
nor U11989 (N_11989,N_11712,N_11762);
xnor U11990 (N_11990,N_11745,N_11825);
or U11991 (N_11991,N_11835,N_11787);
nor U11992 (N_11992,N_11773,N_11763);
nand U11993 (N_11993,N_11722,N_11750);
nand U11994 (N_11994,N_11821,N_11749);
nor U11995 (N_11995,N_11741,N_11752);
xnor U11996 (N_11996,N_11773,N_11771);
nand U11997 (N_11997,N_11751,N_11798);
and U11998 (N_11998,N_11787,N_11778);
or U11999 (N_11999,N_11828,N_11740);
and U12000 (N_12000,N_11898,N_11913);
nand U12001 (N_12001,N_11901,N_11991);
or U12002 (N_12002,N_11880,N_11930);
nor U12003 (N_12003,N_11928,N_11862);
or U12004 (N_12004,N_11997,N_11932);
nand U12005 (N_12005,N_11863,N_11876);
nor U12006 (N_12006,N_11856,N_11915);
or U12007 (N_12007,N_11900,N_11852);
xnor U12008 (N_12008,N_11916,N_11972);
nand U12009 (N_12009,N_11993,N_11895);
nand U12010 (N_12010,N_11906,N_11927);
nor U12011 (N_12011,N_11929,N_11887);
or U12012 (N_12012,N_11870,N_11944);
nor U12013 (N_12013,N_11851,N_11925);
and U12014 (N_12014,N_11919,N_11949);
or U12015 (N_12015,N_11933,N_11998);
nand U12016 (N_12016,N_11952,N_11867);
nor U12017 (N_12017,N_11853,N_11935);
nand U12018 (N_12018,N_11924,N_11905);
or U12019 (N_12019,N_11987,N_11922);
and U12020 (N_12020,N_11908,N_11926);
or U12021 (N_12021,N_11982,N_11878);
xnor U12022 (N_12022,N_11963,N_11873);
nor U12023 (N_12023,N_11902,N_11921);
xnor U12024 (N_12024,N_11959,N_11977);
xnor U12025 (N_12025,N_11874,N_11970);
or U12026 (N_12026,N_11938,N_11960);
xor U12027 (N_12027,N_11868,N_11897);
nor U12028 (N_12028,N_11988,N_11943);
and U12029 (N_12029,N_11858,N_11883);
or U12030 (N_12030,N_11966,N_11865);
or U12031 (N_12031,N_11990,N_11974);
or U12032 (N_12032,N_11983,N_11886);
xor U12033 (N_12033,N_11885,N_11934);
or U12034 (N_12034,N_11909,N_11892);
xor U12035 (N_12035,N_11891,N_11936);
or U12036 (N_12036,N_11882,N_11854);
nand U12037 (N_12037,N_11911,N_11996);
nor U12038 (N_12038,N_11869,N_11871);
or U12039 (N_12039,N_11945,N_11941);
nor U12040 (N_12040,N_11864,N_11971);
xor U12041 (N_12041,N_11950,N_11903);
nor U12042 (N_12042,N_11956,N_11899);
and U12043 (N_12043,N_11912,N_11957);
nand U12044 (N_12044,N_11910,N_11861);
nand U12045 (N_12045,N_11986,N_11875);
or U12046 (N_12046,N_11969,N_11937);
and U12047 (N_12047,N_11973,N_11954);
or U12048 (N_12048,N_11904,N_11979);
and U12049 (N_12049,N_11964,N_11877);
and U12050 (N_12050,N_11978,N_11980);
or U12051 (N_12051,N_11940,N_11946);
xnor U12052 (N_12052,N_11879,N_11955);
and U12053 (N_12053,N_11889,N_11894);
xor U12054 (N_12054,N_11918,N_11958);
nand U12055 (N_12055,N_11866,N_11914);
or U12056 (N_12056,N_11931,N_11881);
and U12057 (N_12057,N_11907,N_11917);
or U12058 (N_12058,N_11992,N_11995);
nand U12059 (N_12059,N_11994,N_11981);
or U12060 (N_12060,N_11884,N_11999);
or U12061 (N_12061,N_11975,N_11857);
nand U12062 (N_12062,N_11965,N_11947);
and U12063 (N_12063,N_11953,N_11896);
nor U12064 (N_12064,N_11961,N_11942);
or U12065 (N_12065,N_11920,N_11989);
and U12066 (N_12066,N_11984,N_11976);
and U12067 (N_12067,N_11939,N_11850);
nor U12068 (N_12068,N_11967,N_11859);
or U12069 (N_12069,N_11888,N_11855);
nor U12070 (N_12070,N_11985,N_11890);
and U12071 (N_12071,N_11860,N_11962);
xnor U12072 (N_12072,N_11923,N_11951);
nand U12073 (N_12073,N_11872,N_11893);
nor U12074 (N_12074,N_11948,N_11968);
nor U12075 (N_12075,N_11938,N_11874);
and U12076 (N_12076,N_11996,N_11928);
or U12077 (N_12077,N_11966,N_11871);
xnor U12078 (N_12078,N_11906,N_11988);
nor U12079 (N_12079,N_11974,N_11933);
xor U12080 (N_12080,N_11925,N_11942);
or U12081 (N_12081,N_11901,N_11943);
or U12082 (N_12082,N_11953,N_11915);
xor U12083 (N_12083,N_11856,N_11862);
xnor U12084 (N_12084,N_11881,N_11951);
nor U12085 (N_12085,N_11982,N_11918);
and U12086 (N_12086,N_11886,N_11988);
nand U12087 (N_12087,N_11933,N_11946);
and U12088 (N_12088,N_11877,N_11953);
nor U12089 (N_12089,N_11932,N_11949);
or U12090 (N_12090,N_11921,N_11999);
nand U12091 (N_12091,N_11867,N_11931);
nor U12092 (N_12092,N_11866,N_11923);
and U12093 (N_12093,N_11934,N_11933);
nor U12094 (N_12094,N_11873,N_11938);
xor U12095 (N_12095,N_11869,N_11977);
and U12096 (N_12096,N_11961,N_11888);
and U12097 (N_12097,N_11991,N_11872);
xor U12098 (N_12098,N_11902,N_11994);
xor U12099 (N_12099,N_11985,N_11996);
xnor U12100 (N_12100,N_11864,N_11979);
nor U12101 (N_12101,N_11938,N_11984);
nand U12102 (N_12102,N_11953,N_11973);
xnor U12103 (N_12103,N_11958,N_11975);
nor U12104 (N_12104,N_11994,N_11952);
or U12105 (N_12105,N_11863,N_11879);
nor U12106 (N_12106,N_11963,N_11876);
xor U12107 (N_12107,N_11887,N_11968);
nand U12108 (N_12108,N_11860,N_11896);
or U12109 (N_12109,N_11941,N_11933);
nor U12110 (N_12110,N_11945,N_11969);
or U12111 (N_12111,N_11957,N_11954);
or U12112 (N_12112,N_11947,N_11917);
nor U12113 (N_12113,N_11888,N_11913);
nand U12114 (N_12114,N_11935,N_11878);
nor U12115 (N_12115,N_11949,N_11874);
nor U12116 (N_12116,N_11939,N_11957);
nand U12117 (N_12117,N_11996,N_11993);
xor U12118 (N_12118,N_11900,N_11939);
or U12119 (N_12119,N_11943,N_11937);
nand U12120 (N_12120,N_11948,N_11965);
nand U12121 (N_12121,N_11890,N_11855);
nand U12122 (N_12122,N_11977,N_11963);
or U12123 (N_12123,N_11890,N_11867);
nand U12124 (N_12124,N_11858,N_11911);
or U12125 (N_12125,N_11971,N_11894);
xor U12126 (N_12126,N_11944,N_11897);
nand U12127 (N_12127,N_11868,N_11986);
xnor U12128 (N_12128,N_11894,N_11860);
xnor U12129 (N_12129,N_11948,N_11879);
xor U12130 (N_12130,N_11917,N_11884);
or U12131 (N_12131,N_11961,N_11957);
or U12132 (N_12132,N_11953,N_11910);
and U12133 (N_12133,N_11919,N_11898);
and U12134 (N_12134,N_11888,N_11927);
nor U12135 (N_12135,N_11905,N_11868);
and U12136 (N_12136,N_11917,N_11991);
xnor U12137 (N_12137,N_11911,N_11891);
xnor U12138 (N_12138,N_11888,N_11956);
nand U12139 (N_12139,N_11933,N_11908);
or U12140 (N_12140,N_11954,N_11942);
nand U12141 (N_12141,N_11948,N_11972);
or U12142 (N_12142,N_11907,N_11941);
and U12143 (N_12143,N_11958,N_11949);
nor U12144 (N_12144,N_11858,N_11937);
nand U12145 (N_12145,N_11903,N_11981);
nand U12146 (N_12146,N_11956,N_11884);
and U12147 (N_12147,N_11901,N_11853);
nand U12148 (N_12148,N_11869,N_11992);
nor U12149 (N_12149,N_11982,N_11864);
nor U12150 (N_12150,N_12112,N_12120);
xor U12151 (N_12151,N_12077,N_12119);
nor U12152 (N_12152,N_12051,N_12116);
and U12153 (N_12153,N_12066,N_12022);
and U12154 (N_12154,N_12011,N_12067);
or U12155 (N_12155,N_12081,N_12005);
xor U12156 (N_12156,N_12145,N_12125);
or U12157 (N_12157,N_12096,N_12088);
nand U12158 (N_12158,N_12135,N_12035);
xor U12159 (N_12159,N_12020,N_12071);
nand U12160 (N_12160,N_12069,N_12085);
or U12161 (N_12161,N_12059,N_12140);
nand U12162 (N_12162,N_12072,N_12045);
nor U12163 (N_12163,N_12091,N_12047);
and U12164 (N_12164,N_12147,N_12082);
xor U12165 (N_12165,N_12057,N_12117);
or U12166 (N_12166,N_12026,N_12103);
xnor U12167 (N_12167,N_12037,N_12021);
xor U12168 (N_12168,N_12121,N_12108);
or U12169 (N_12169,N_12041,N_12030);
and U12170 (N_12170,N_12074,N_12094);
nand U12171 (N_12171,N_12139,N_12095);
nand U12172 (N_12172,N_12039,N_12040);
and U12173 (N_12173,N_12015,N_12068);
nor U12174 (N_12174,N_12086,N_12075);
xnor U12175 (N_12175,N_12017,N_12031);
xor U12176 (N_12176,N_12093,N_12028);
nor U12177 (N_12177,N_12090,N_12136);
or U12178 (N_12178,N_12054,N_12138);
xor U12179 (N_12179,N_12133,N_12064);
or U12180 (N_12180,N_12043,N_12148);
or U12181 (N_12181,N_12123,N_12027);
or U12182 (N_12182,N_12099,N_12029);
nor U12183 (N_12183,N_12137,N_12058);
nor U12184 (N_12184,N_12019,N_12087);
nor U12185 (N_12185,N_12107,N_12110);
nor U12186 (N_12186,N_12048,N_12053);
nand U12187 (N_12187,N_12126,N_12062);
nand U12188 (N_12188,N_12050,N_12129);
nand U12189 (N_12189,N_12118,N_12024);
nor U12190 (N_12190,N_12052,N_12060);
and U12191 (N_12191,N_12100,N_12008);
and U12192 (N_12192,N_12101,N_12134);
or U12193 (N_12193,N_12084,N_12127);
or U12194 (N_12194,N_12056,N_12128);
nand U12195 (N_12195,N_12013,N_12003);
nor U12196 (N_12196,N_12012,N_12115);
nand U12197 (N_12197,N_12034,N_12073);
and U12198 (N_12198,N_12106,N_12042);
nor U12199 (N_12199,N_12046,N_12124);
nor U12200 (N_12200,N_12033,N_12023);
and U12201 (N_12201,N_12009,N_12063);
or U12202 (N_12202,N_12089,N_12092);
or U12203 (N_12203,N_12114,N_12102);
or U12204 (N_12204,N_12098,N_12016);
or U12205 (N_12205,N_12122,N_12010);
xnor U12206 (N_12206,N_12065,N_12032);
and U12207 (N_12207,N_12076,N_12143);
nand U12208 (N_12208,N_12018,N_12079);
or U12209 (N_12209,N_12004,N_12104);
or U12210 (N_12210,N_12149,N_12083);
xnor U12211 (N_12211,N_12025,N_12131);
nand U12212 (N_12212,N_12014,N_12049);
xor U12213 (N_12213,N_12006,N_12000);
and U12214 (N_12214,N_12105,N_12078);
xor U12215 (N_12215,N_12070,N_12113);
nor U12216 (N_12216,N_12141,N_12142);
or U12217 (N_12217,N_12097,N_12002);
xor U12218 (N_12218,N_12044,N_12111);
xor U12219 (N_12219,N_12080,N_12144);
nor U12220 (N_12220,N_12130,N_12061);
nor U12221 (N_12221,N_12132,N_12001);
or U12222 (N_12222,N_12109,N_12146);
or U12223 (N_12223,N_12055,N_12036);
xor U12224 (N_12224,N_12007,N_12038);
nand U12225 (N_12225,N_12017,N_12082);
nor U12226 (N_12226,N_12087,N_12026);
xnor U12227 (N_12227,N_12010,N_12023);
xor U12228 (N_12228,N_12129,N_12044);
nor U12229 (N_12229,N_12085,N_12053);
nand U12230 (N_12230,N_12122,N_12083);
or U12231 (N_12231,N_12128,N_12089);
xnor U12232 (N_12232,N_12136,N_12089);
or U12233 (N_12233,N_12103,N_12068);
xnor U12234 (N_12234,N_12057,N_12041);
and U12235 (N_12235,N_12090,N_12117);
or U12236 (N_12236,N_12074,N_12017);
and U12237 (N_12237,N_12102,N_12021);
nand U12238 (N_12238,N_12127,N_12055);
or U12239 (N_12239,N_12104,N_12006);
xor U12240 (N_12240,N_12021,N_12126);
nand U12241 (N_12241,N_12102,N_12047);
xor U12242 (N_12242,N_12132,N_12044);
xnor U12243 (N_12243,N_12053,N_12149);
nor U12244 (N_12244,N_12114,N_12066);
xnor U12245 (N_12245,N_12031,N_12096);
nor U12246 (N_12246,N_12097,N_12133);
nor U12247 (N_12247,N_12136,N_12149);
nand U12248 (N_12248,N_12043,N_12075);
and U12249 (N_12249,N_12050,N_12046);
and U12250 (N_12250,N_12025,N_12104);
nor U12251 (N_12251,N_12039,N_12087);
xor U12252 (N_12252,N_12099,N_12085);
or U12253 (N_12253,N_12144,N_12134);
xnor U12254 (N_12254,N_12015,N_12074);
nand U12255 (N_12255,N_12125,N_12058);
nor U12256 (N_12256,N_12073,N_12059);
nor U12257 (N_12257,N_12040,N_12021);
and U12258 (N_12258,N_12053,N_12089);
or U12259 (N_12259,N_12085,N_12097);
xor U12260 (N_12260,N_12102,N_12109);
or U12261 (N_12261,N_12050,N_12104);
xor U12262 (N_12262,N_12083,N_12109);
xor U12263 (N_12263,N_12050,N_12052);
nor U12264 (N_12264,N_12097,N_12018);
and U12265 (N_12265,N_12085,N_12101);
xor U12266 (N_12266,N_12142,N_12095);
nand U12267 (N_12267,N_12053,N_12038);
nor U12268 (N_12268,N_12008,N_12049);
nor U12269 (N_12269,N_12067,N_12115);
and U12270 (N_12270,N_12139,N_12142);
or U12271 (N_12271,N_12110,N_12045);
xnor U12272 (N_12272,N_12050,N_12030);
xor U12273 (N_12273,N_12066,N_12011);
or U12274 (N_12274,N_12125,N_12021);
xor U12275 (N_12275,N_12147,N_12041);
and U12276 (N_12276,N_12087,N_12128);
nor U12277 (N_12277,N_12034,N_12123);
nand U12278 (N_12278,N_12046,N_12101);
or U12279 (N_12279,N_12041,N_12085);
and U12280 (N_12280,N_12090,N_12009);
and U12281 (N_12281,N_12091,N_12059);
xor U12282 (N_12282,N_12145,N_12004);
nand U12283 (N_12283,N_12028,N_12113);
xor U12284 (N_12284,N_12028,N_12148);
nand U12285 (N_12285,N_12077,N_12015);
nor U12286 (N_12286,N_12123,N_12036);
nor U12287 (N_12287,N_12004,N_12024);
nor U12288 (N_12288,N_12020,N_12031);
nor U12289 (N_12289,N_12001,N_12063);
nand U12290 (N_12290,N_12078,N_12070);
nor U12291 (N_12291,N_12083,N_12103);
xnor U12292 (N_12292,N_12073,N_12035);
or U12293 (N_12293,N_12148,N_12016);
or U12294 (N_12294,N_12109,N_12121);
xor U12295 (N_12295,N_12055,N_12082);
or U12296 (N_12296,N_12146,N_12147);
nand U12297 (N_12297,N_12062,N_12013);
or U12298 (N_12298,N_12098,N_12028);
nand U12299 (N_12299,N_12020,N_12033);
nor U12300 (N_12300,N_12199,N_12263);
nand U12301 (N_12301,N_12292,N_12179);
and U12302 (N_12302,N_12283,N_12243);
nand U12303 (N_12303,N_12181,N_12200);
xnor U12304 (N_12304,N_12235,N_12209);
xnor U12305 (N_12305,N_12198,N_12151);
or U12306 (N_12306,N_12239,N_12270);
nor U12307 (N_12307,N_12178,N_12204);
xor U12308 (N_12308,N_12280,N_12272);
nand U12309 (N_12309,N_12177,N_12186);
nor U12310 (N_12310,N_12191,N_12152);
nor U12311 (N_12311,N_12251,N_12176);
xnor U12312 (N_12312,N_12213,N_12234);
nand U12313 (N_12313,N_12217,N_12281);
or U12314 (N_12314,N_12242,N_12159);
and U12315 (N_12315,N_12288,N_12214);
and U12316 (N_12316,N_12228,N_12286);
and U12317 (N_12317,N_12282,N_12299);
or U12318 (N_12318,N_12240,N_12261);
nand U12319 (N_12319,N_12154,N_12211);
xnor U12320 (N_12320,N_12277,N_12188);
or U12321 (N_12321,N_12150,N_12262);
and U12322 (N_12322,N_12201,N_12189);
nand U12323 (N_12323,N_12285,N_12157);
nand U12324 (N_12324,N_12156,N_12265);
and U12325 (N_12325,N_12275,N_12291);
nand U12326 (N_12326,N_12215,N_12252);
and U12327 (N_12327,N_12172,N_12206);
nor U12328 (N_12328,N_12208,N_12203);
nand U12329 (N_12329,N_12212,N_12207);
nor U12330 (N_12330,N_12173,N_12226);
xor U12331 (N_12331,N_12182,N_12169);
or U12332 (N_12332,N_12174,N_12258);
or U12333 (N_12333,N_12225,N_12232);
and U12334 (N_12334,N_12247,N_12210);
or U12335 (N_12335,N_12236,N_12222);
and U12336 (N_12336,N_12278,N_12266);
xnor U12337 (N_12337,N_12295,N_12192);
and U12338 (N_12338,N_12248,N_12153);
nand U12339 (N_12339,N_12268,N_12241);
nor U12340 (N_12340,N_12271,N_12166);
nor U12341 (N_12341,N_12260,N_12162);
and U12342 (N_12342,N_12264,N_12224);
xor U12343 (N_12343,N_12194,N_12257);
nand U12344 (N_12344,N_12233,N_12185);
xor U12345 (N_12345,N_12255,N_12158);
nand U12346 (N_12346,N_12196,N_12168);
xnor U12347 (N_12347,N_12274,N_12287);
xnor U12348 (N_12348,N_12167,N_12227);
nand U12349 (N_12349,N_12273,N_12202);
xor U12350 (N_12350,N_12250,N_12163);
or U12351 (N_12351,N_12279,N_12253);
xnor U12352 (N_12352,N_12171,N_12218);
or U12353 (N_12353,N_12216,N_12297);
nand U12354 (N_12354,N_12259,N_12293);
nand U12355 (N_12355,N_12249,N_12231);
and U12356 (N_12356,N_12164,N_12165);
xor U12357 (N_12357,N_12170,N_12161);
and U12358 (N_12358,N_12269,N_12190);
xor U12359 (N_12359,N_12221,N_12289);
nand U12360 (N_12360,N_12238,N_12175);
xnor U12361 (N_12361,N_12195,N_12220);
and U12362 (N_12362,N_12223,N_12267);
or U12363 (N_12363,N_12205,N_12193);
xnor U12364 (N_12364,N_12298,N_12290);
xnor U12365 (N_12365,N_12284,N_12230);
nand U12366 (N_12366,N_12229,N_12246);
nand U12367 (N_12367,N_12160,N_12245);
nor U12368 (N_12368,N_12180,N_12155);
nand U12369 (N_12369,N_12183,N_12294);
nand U12370 (N_12370,N_12244,N_12187);
and U12371 (N_12371,N_12254,N_12197);
nand U12372 (N_12372,N_12256,N_12184);
or U12373 (N_12373,N_12237,N_12276);
or U12374 (N_12374,N_12296,N_12219);
or U12375 (N_12375,N_12252,N_12262);
nor U12376 (N_12376,N_12213,N_12190);
and U12377 (N_12377,N_12205,N_12288);
nor U12378 (N_12378,N_12151,N_12286);
and U12379 (N_12379,N_12158,N_12241);
or U12380 (N_12380,N_12184,N_12207);
xor U12381 (N_12381,N_12294,N_12164);
nand U12382 (N_12382,N_12256,N_12221);
nand U12383 (N_12383,N_12287,N_12215);
nand U12384 (N_12384,N_12163,N_12239);
nand U12385 (N_12385,N_12271,N_12184);
xor U12386 (N_12386,N_12171,N_12155);
and U12387 (N_12387,N_12163,N_12228);
xnor U12388 (N_12388,N_12151,N_12238);
or U12389 (N_12389,N_12296,N_12263);
nor U12390 (N_12390,N_12158,N_12239);
and U12391 (N_12391,N_12271,N_12266);
xnor U12392 (N_12392,N_12282,N_12156);
nand U12393 (N_12393,N_12246,N_12292);
xnor U12394 (N_12394,N_12229,N_12282);
nor U12395 (N_12395,N_12159,N_12214);
nand U12396 (N_12396,N_12229,N_12160);
or U12397 (N_12397,N_12255,N_12289);
or U12398 (N_12398,N_12295,N_12200);
or U12399 (N_12399,N_12231,N_12236);
nand U12400 (N_12400,N_12271,N_12286);
and U12401 (N_12401,N_12226,N_12294);
nand U12402 (N_12402,N_12172,N_12254);
xnor U12403 (N_12403,N_12154,N_12231);
and U12404 (N_12404,N_12291,N_12264);
nor U12405 (N_12405,N_12243,N_12264);
and U12406 (N_12406,N_12283,N_12172);
xnor U12407 (N_12407,N_12262,N_12255);
or U12408 (N_12408,N_12186,N_12284);
nand U12409 (N_12409,N_12249,N_12162);
nor U12410 (N_12410,N_12203,N_12237);
or U12411 (N_12411,N_12228,N_12298);
or U12412 (N_12412,N_12299,N_12157);
nand U12413 (N_12413,N_12286,N_12199);
and U12414 (N_12414,N_12217,N_12189);
nand U12415 (N_12415,N_12150,N_12282);
or U12416 (N_12416,N_12244,N_12221);
or U12417 (N_12417,N_12151,N_12206);
nand U12418 (N_12418,N_12287,N_12224);
nand U12419 (N_12419,N_12237,N_12207);
and U12420 (N_12420,N_12174,N_12244);
or U12421 (N_12421,N_12266,N_12293);
nand U12422 (N_12422,N_12207,N_12291);
nor U12423 (N_12423,N_12159,N_12287);
nor U12424 (N_12424,N_12160,N_12178);
nor U12425 (N_12425,N_12293,N_12216);
nand U12426 (N_12426,N_12250,N_12196);
and U12427 (N_12427,N_12183,N_12243);
nor U12428 (N_12428,N_12155,N_12217);
xnor U12429 (N_12429,N_12245,N_12274);
nor U12430 (N_12430,N_12272,N_12200);
xnor U12431 (N_12431,N_12262,N_12257);
or U12432 (N_12432,N_12247,N_12189);
xnor U12433 (N_12433,N_12207,N_12254);
nand U12434 (N_12434,N_12156,N_12167);
and U12435 (N_12435,N_12280,N_12275);
nor U12436 (N_12436,N_12179,N_12156);
nand U12437 (N_12437,N_12271,N_12224);
or U12438 (N_12438,N_12192,N_12166);
or U12439 (N_12439,N_12298,N_12220);
nor U12440 (N_12440,N_12185,N_12238);
nand U12441 (N_12441,N_12174,N_12208);
or U12442 (N_12442,N_12202,N_12221);
nand U12443 (N_12443,N_12284,N_12169);
nor U12444 (N_12444,N_12267,N_12161);
and U12445 (N_12445,N_12169,N_12180);
nor U12446 (N_12446,N_12212,N_12186);
and U12447 (N_12447,N_12277,N_12172);
xor U12448 (N_12448,N_12233,N_12168);
and U12449 (N_12449,N_12176,N_12249);
and U12450 (N_12450,N_12321,N_12358);
xnor U12451 (N_12451,N_12383,N_12332);
nor U12452 (N_12452,N_12309,N_12394);
or U12453 (N_12453,N_12374,N_12322);
xor U12454 (N_12454,N_12424,N_12341);
nor U12455 (N_12455,N_12378,N_12313);
and U12456 (N_12456,N_12305,N_12392);
or U12457 (N_12457,N_12344,N_12425);
xnor U12458 (N_12458,N_12333,N_12306);
nand U12459 (N_12459,N_12349,N_12408);
nand U12460 (N_12460,N_12391,N_12380);
xnor U12461 (N_12461,N_12324,N_12367);
nor U12462 (N_12462,N_12303,N_12437);
or U12463 (N_12463,N_12411,N_12304);
nand U12464 (N_12464,N_12444,N_12359);
and U12465 (N_12465,N_12357,N_12347);
nor U12466 (N_12466,N_12387,N_12336);
or U12467 (N_12467,N_12433,N_12429);
nor U12468 (N_12468,N_12366,N_12330);
nor U12469 (N_12469,N_12362,N_12431);
and U12470 (N_12470,N_12370,N_12384);
or U12471 (N_12471,N_12377,N_12334);
or U12472 (N_12472,N_12389,N_12312);
and U12473 (N_12473,N_12420,N_12318);
or U12474 (N_12474,N_12390,N_12368);
nor U12475 (N_12475,N_12413,N_12440);
or U12476 (N_12476,N_12327,N_12421);
xnor U12477 (N_12477,N_12436,N_12400);
and U12478 (N_12478,N_12423,N_12414);
xor U12479 (N_12479,N_12430,N_12398);
nor U12480 (N_12480,N_12361,N_12382);
and U12481 (N_12481,N_12355,N_12376);
nand U12482 (N_12482,N_12308,N_12432);
and U12483 (N_12483,N_12434,N_12315);
nand U12484 (N_12484,N_12375,N_12331);
nor U12485 (N_12485,N_12326,N_12345);
nand U12486 (N_12486,N_12381,N_12350);
xor U12487 (N_12487,N_12438,N_12337);
nor U12488 (N_12488,N_12301,N_12426);
or U12489 (N_12489,N_12415,N_12419);
or U12490 (N_12490,N_12428,N_12353);
nor U12491 (N_12491,N_12365,N_12385);
xnor U12492 (N_12492,N_12447,N_12348);
nand U12493 (N_12493,N_12448,N_12446);
xnor U12494 (N_12494,N_12442,N_12416);
nor U12495 (N_12495,N_12449,N_12339);
nand U12496 (N_12496,N_12397,N_12354);
nand U12497 (N_12497,N_12329,N_12343);
nand U12498 (N_12498,N_12443,N_12328);
nor U12499 (N_12499,N_12311,N_12351);
xor U12500 (N_12500,N_12439,N_12352);
xnor U12501 (N_12501,N_12396,N_12369);
or U12502 (N_12502,N_12372,N_12316);
nand U12503 (N_12503,N_12401,N_12363);
and U12504 (N_12504,N_12417,N_12379);
nor U12505 (N_12505,N_12356,N_12307);
nand U12506 (N_12506,N_12418,N_12364);
xor U12507 (N_12507,N_12373,N_12346);
xor U12508 (N_12508,N_12340,N_12360);
nand U12509 (N_12509,N_12320,N_12371);
nand U12510 (N_12510,N_12388,N_12406);
or U12511 (N_12511,N_12335,N_12393);
nor U12512 (N_12512,N_12402,N_12395);
and U12513 (N_12513,N_12409,N_12422);
or U12514 (N_12514,N_12427,N_12300);
and U12515 (N_12515,N_12325,N_12405);
nor U12516 (N_12516,N_12403,N_12342);
and U12517 (N_12517,N_12404,N_12412);
nand U12518 (N_12518,N_12399,N_12314);
nand U12519 (N_12519,N_12407,N_12319);
or U12520 (N_12520,N_12302,N_12386);
xnor U12521 (N_12521,N_12323,N_12317);
xnor U12522 (N_12522,N_12445,N_12441);
nor U12523 (N_12523,N_12410,N_12338);
nand U12524 (N_12524,N_12435,N_12310);
and U12525 (N_12525,N_12366,N_12398);
and U12526 (N_12526,N_12429,N_12375);
nor U12527 (N_12527,N_12358,N_12311);
or U12528 (N_12528,N_12311,N_12420);
and U12529 (N_12529,N_12409,N_12371);
or U12530 (N_12530,N_12332,N_12379);
nand U12531 (N_12531,N_12341,N_12331);
xor U12532 (N_12532,N_12433,N_12322);
nor U12533 (N_12533,N_12433,N_12435);
xor U12534 (N_12534,N_12375,N_12444);
and U12535 (N_12535,N_12312,N_12378);
or U12536 (N_12536,N_12359,N_12415);
nor U12537 (N_12537,N_12304,N_12438);
nor U12538 (N_12538,N_12390,N_12362);
nor U12539 (N_12539,N_12385,N_12310);
or U12540 (N_12540,N_12431,N_12316);
nand U12541 (N_12541,N_12374,N_12363);
and U12542 (N_12542,N_12340,N_12325);
xnor U12543 (N_12543,N_12331,N_12384);
nor U12544 (N_12544,N_12316,N_12369);
nand U12545 (N_12545,N_12394,N_12373);
xnor U12546 (N_12546,N_12382,N_12431);
or U12547 (N_12547,N_12360,N_12371);
and U12548 (N_12548,N_12415,N_12376);
nor U12549 (N_12549,N_12302,N_12367);
xnor U12550 (N_12550,N_12409,N_12360);
and U12551 (N_12551,N_12406,N_12326);
nor U12552 (N_12552,N_12341,N_12431);
nand U12553 (N_12553,N_12393,N_12322);
nand U12554 (N_12554,N_12446,N_12396);
nand U12555 (N_12555,N_12350,N_12446);
or U12556 (N_12556,N_12325,N_12419);
nand U12557 (N_12557,N_12331,N_12395);
nand U12558 (N_12558,N_12360,N_12308);
and U12559 (N_12559,N_12415,N_12393);
xor U12560 (N_12560,N_12358,N_12372);
nand U12561 (N_12561,N_12393,N_12417);
nor U12562 (N_12562,N_12343,N_12390);
xnor U12563 (N_12563,N_12400,N_12312);
xnor U12564 (N_12564,N_12357,N_12401);
xor U12565 (N_12565,N_12328,N_12338);
nand U12566 (N_12566,N_12328,N_12429);
or U12567 (N_12567,N_12374,N_12428);
nor U12568 (N_12568,N_12427,N_12306);
nand U12569 (N_12569,N_12439,N_12424);
xor U12570 (N_12570,N_12420,N_12373);
nor U12571 (N_12571,N_12342,N_12335);
nor U12572 (N_12572,N_12356,N_12334);
xor U12573 (N_12573,N_12424,N_12325);
or U12574 (N_12574,N_12407,N_12341);
or U12575 (N_12575,N_12331,N_12436);
and U12576 (N_12576,N_12371,N_12340);
or U12577 (N_12577,N_12350,N_12389);
and U12578 (N_12578,N_12305,N_12309);
and U12579 (N_12579,N_12316,N_12362);
xor U12580 (N_12580,N_12353,N_12368);
nor U12581 (N_12581,N_12304,N_12334);
or U12582 (N_12582,N_12318,N_12441);
xnor U12583 (N_12583,N_12402,N_12392);
and U12584 (N_12584,N_12449,N_12380);
nor U12585 (N_12585,N_12357,N_12329);
and U12586 (N_12586,N_12303,N_12401);
nor U12587 (N_12587,N_12427,N_12445);
and U12588 (N_12588,N_12340,N_12439);
or U12589 (N_12589,N_12408,N_12429);
and U12590 (N_12590,N_12378,N_12356);
xor U12591 (N_12591,N_12415,N_12411);
xnor U12592 (N_12592,N_12390,N_12358);
nand U12593 (N_12593,N_12301,N_12443);
or U12594 (N_12594,N_12399,N_12375);
or U12595 (N_12595,N_12446,N_12414);
xor U12596 (N_12596,N_12332,N_12336);
nor U12597 (N_12597,N_12351,N_12359);
xor U12598 (N_12598,N_12302,N_12364);
nor U12599 (N_12599,N_12311,N_12338);
nand U12600 (N_12600,N_12574,N_12583);
nand U12601 (N_12601,N_12513,N_12475);
xnor U12602 (N_12602,N_12451,N_12462);
nand U12603 (N_12603,N_12504,N_12598);
nor U12604 (N_12604,N_12516,N_12535);
or U12605 (N_12605,N_12595,N_12577);
nor U12606 (N_12606,N_12571,N_12537);
xor U12607 (N_12607,N_12532,N_12469);
nor U12608 (N_12608,N_12570,N_12518);
xnor U12609 (N_12609,N_12487,N_12497);
nor U12610 (N_12610,N_12527,N_12556);
and U12611 (N_12611,N_12544,N_12564);
nand U12612 (N_12612,N_12481,N_12576);
or U12613 (N_12613,N_12554,N_12596);
or U12614 (N_12614,N_12508,N_12555);
or U12615 (N_12615,N_12498,N_12530);
or U12616 (N_12616,N_12529,N_12536);
or U12617 (N_12617,N_12483,N_12480);
nand U12618 (N_12618,N_12509,N_12499);
xor U12619 (N_12619,N_12524,N_12495);
xnor U12620 (N_12620,N_12477,N_12579);
xor U12621 (N_12621,N_12492,N_12502);
nand U12622 (N_12622,N_12522,N_12533);
or U12623 (N_12623,N_12540,N_12547);
and U12624 (N_12624,N_12546,N_12455);
nor U12625 (N_12625,N_12501,N_12592);
nand U12626 (N_12626,N_12569,N_12515);
nor U12627 (N_12627,N_12553,N_12461);
xor U12628 (N_12628,N_12534,N_12582);
xor U12629 (N_12629,N_12531,N_12493);
nor U12630 (N_12630,N_12588,N_12568);
nand U12631 (N_12631,N_12463,N_12580);
xnor U12632 (N_12632,N_12542,N_12486);
or U12633 (N_12633,N_12500,N_12484);
nor U12634 (N_12634,N_12511,N_12563);
nor U12635 (N_12635,N_12549,N_12591);
nand U12636 (N_12636,N_12473,N_12528);
nor U12637 (N_12637,N_12586,N_12597);
nor U12638 (N_12638,N_12485,N_12465);
nor U12639 (N_12639,N_12548,N_12454);
and U12640 (N_12640,N_12543,N_12472);
nor U12641 (N_12641,N_12521,N_12452);
nand U12642 (N_12642,N_12457,N_12594);
or U12643 (N_12643,N_12559,N_12482);
xor U12644 (N_12644,N_12471,N_12565);
and U12645 (N_12645,N_12491,N_12494);
nor U12646 (N_12646,N_12599,N_12507);
or U12647 (N_12647,N_12489,N_12470);
xor U12648 (N_12648,N_12593,N_12545);
and U12649 (N_12649,N_12560,N_12572);
or U12650 (N_12650,N_12551,N_12550);
nor U12651 (N_12651,N_12561,N_12519);
xor U12652 (N_12652,N_12562,N_12458);
xor U12653 (N_12653,N_12478,N_12552);
and U12654 (N_12654,N_12558,N_12460);
and U12655 (N_12655,N_12584,N_12566);
nor U12656 (N_12656,N_12474,N_12517);
xor U12657 (N_12657,N_12573,N_12512);
nor U12658 (N_12658,N_12479,N_12456);
and U12659 (N_12659,N_12488,N_12557);
nor U12660 (N_12660,N_12587,N_12539);
and U12661 (N_12661,N_12464,N_12476);
nor U12662 (N_12662,N_12496,N_12490);
nand U12663 (N_12663,N_12590,N_12467);
and U12664 (N_12664,N_12503,N_12453);
or U12665 (N_12665,N_12589,N_12578);
and U12666 (N_12666,N_12538,N_12520);
and U12667 (N_12667,N_12575,N_12567);
nand U12668 (N_12668,N_12525,N_12459);
or U12669 (N_12669,N_12468,N_12585);
nand U12670 (N_12670,N_12505,N_12450);
nand U12671 (N_12671,N_12466,N_12526);
and U12672 (N_12672,N_12581,N_12506);
nor U12673 (N_12673,N_12510,N_12541);
and U12674 (N_12674,N_12514,N_12523);
or U12675 (N_12675,N_12541,N_12598);
and U12676 (N_12676,N_12469,N_12555);
nor U12677 (N_12677,N_12588,N_12453);
nor U12678 (N_12678,N_12509,N_12468);
xnor U12679 (N_12679,N_12483,N_12560);
nor U12680 (N_12680,N_12487,N_12474);
nor U12681 (N_12681,N_12464,N_12572);
xor U12682 (N_12682,N_12511,N_12597);
nor U12683 (N_12683,N_12561,N_12513);
xnor U12684 (N_12684,N_12479,N_12497);
and U12685 (N_12685,N_12474,N_12482);
and U12686 (N_12686,N_12469,N_12482);
xor U12687 (N_12687,N_12549,N_12554);
xor U12688 (N_12688,N_12486,N_12518);
nor U12689 (N_12689,N_12491,N_12592);
or U12690 (N_12690,N_12465,N_12476);
and U12691 (N_12691,N_12499,N_12550);
nor U12692 (N_12692,N_12536,N_12538);
xnor U12693 (N_12693,N_12489,N_12540);
nor U12694 (N_12694,N_12536,N_12475);
xor U12695 (N_12695,N_12524,N_12504);
xnor U12696 (N_12696,N_12580,N_12454);
nor U12697 (N_12697,N_12586,N_12568);
and U12698 (N_12698,N_12544,N_12493);
xor U12699 (N_12699,N_12561,N_12558);
nand U12700 (N_12700,N_12483,N_12485);
nor U12701 (N_12701,N_12459,N_12488);
or U12702 (N_12702,N_12553,N_12499);
and U12703 (N_12703,N_12593,N_12480);
and U12704 (N_12704,N_12594,N_12568);
nor U12705 (N_12705,N_12513,N_12492);
and U12706 (N_12706,N_12546,N_12588);
or U12707 (N_12707,N_12573,N_12472);
nand U12708 (N_12708,N_12503,N_12464);
xor U12709 (N_12709,N_12471,N_12534);
and U12710 (N_12710,N_12594,N_12475);
or U12711 (N_12711,N_12489,N_12592);
or U12712 (N_12712,N_12563,N_12579);
xnor U12713 (N_12713,N_12498,N_12582);
nand U12714 (N_12714,N_12504,N_12479);
or U12715 (N_12715,N_12513,N_12516);
xor U12716 (N_12716,N_12561,N_12599);
and U12717 (N_12717,N_12542,N_12482);
or U12718 (N_12718,N_12576,N_12531);
and U12719 (N_12719,N_12478,N_12488);
and U12720 (N_12720,N_12474,N_12534);
and U12721 (N_12721,N_12472,N_12504);
or U12722 (N_12722,N_12547,N_12566);
nand U12723 (N_12723,N_12479,N_12495);
or U12724 (N_12724,N_12530,N_12472);
and U12725 (N_12725,N_12501,N_12576);
nand U12726 (N_12726,N_12539,N_12518);
or U12727 (N_12727,N_12564,N_12538);
xnor U12728 (N_12728,N_12571,N_12564);
nor U12729 (N_12729,N_12466,N_12524);
and U12730 (N_12730,N_12564,N_12589);
nand U12731 (N_12731,N_12472,N_12582);
nand U12732 (N_12732,N_12535,N_12529);
nor U12733 (N_12733,N_12490,N_12562);
nand U12734 (N_12734,N_12599,N_12496);
and U12735 (N_12735,N_12478,N_12484);
xnor U12736 (N_12736,N_12491,N_12536);
and U12737 (N_12737,N_12458,N_12584);
nand U12738 (N_12738,N_12488,N_12520);
or U12739 (N_12739,N_12584,N_12599);
or U12740 (N_12740,N_12557,N_12534);
or U12741 (N_12741,N_12497,N_12573);
and U12742 (N_12742,N_12490,N_12469);
and U12743 (N_12743,N_12499,N_12459);
nand U12744 (N_12744,N_12528,N_12503);
nand U12745 (N_12745,N_12481,N_12456);
nand U12746 (N_12746,N_12490,N_12524);
nor U12747 (N_12747,N_12551,N_12487);
nor U12748 (N_12748,N_12473,N_12529);
xor U12749 (N_12749,N_12549,N_12513);
nor U12750 (N_12750,N_12726,N_12621);
and U12751 (N_12751,N_12710,N_12651);
or U12752 (N_12752,N_12688,N_12630);
and U12753 (N_12753,N_12639,N_12644);
or U12754 (N_12754,N_12645,N_12615);
and U12755 (N_12755,N_12623,N_12735);
nand U12756 (N_12756,N_12653,N_12665);
and U12757 (N_12757,N_12648,N_12703);
nor U12758 (N_12758,N_12734,N_12696);
nand U12759 (N_12759,N_12633,N_12652);
or U12760 (N_12760,N_12607,N_12698);
and U12761 (N_12761,N_12655,N_12672);
and U12762 (N_12762,N_12641,N_12746);
nor U12763 (N_12763,N_12627,N_12705);
xnor U12764 (N_12764,N_12690,N_12745);
xnor U12765 (N_12765,N_12727,N_12673);
nor U12766 (N_12766,N_12612,N_12663);
nand U12767 (N_12767,N_12724,N_12739);
xor U12768 (N_12768,N_12624,N_12647);
nand U12769 (N_12769,N_12731,N_12674);
or U12770 (N_12770,N_12602,N_12716);
xnor U12771 (N_12771,N_12671,N_12702);
or U12772 (N_12772,N_12650,N_12740);
nand U12773 (N_12773,N_12662,N_12642);
or U12774 (N_12774,N_12631,N_12667);
and U12775 (N_12775,N_12635,N_12747);
nand U12776 (N_12776,N_12658,N_12700);
nand U12777 (N_12777,N_12711,N_12722);
or U12778 (N_12778,N_12725,N_12741);
nor U12779 (N_12779,N_12620,N_12640);
xnor U12780 (N_12780,N_12654,N_12636);
or U12781 (N_12781,N_12697,N_12695);
or U12782 (N_12782,N_12675,N_12719);
or U12783 (N_12783,N_12732,N_12670);
or U12784 (N_12784,N_12669,N_12699);
or U12785 (N_12785,N_12701,N_12613);
nand U12786 (N_12786,N_12738,N_12618);
xnor U12787 (N_12787,N_12714,N_12606);
xor U12788 (N_12788,N_12628,N_12728);
nand U12789 (N_12789,N_12689,N_12609);
and U12790 (N_12790,N_12679,N_12611);
nand U12791 (N_12791,N_12704,N_12638);
nor U12792 (N_12792,N_12718,N_12678);
nand U12793 (N_12793,N_12656,N_12637);
nor U12794 (N_12794,N_12715,N_12707);
or U12795 (N_12795,N_12677,N_12687);
xnor U12796 (N_12796,N_12730,N_12708);
nand U12797 (N_12797,N_12733,N_12604);
xor U12798 (N_12798,N_12717,N_12683);
and U12799 (N_12799,N_12723,N_12619);
and U12800 (N_12800,N_12626,N_12720);
nand U12801 (N_12801,N_12629,N_12692);
nand U12802 (N_12802,N_12676,N_12643);
xnor U12803 (N_12803,N_12691,N_12646);
or U12804 (N_12804,N_12634,N_12729);
or U12805 (N_12805,N_12659,N_12614);
and U12806 (N_12806,N_12749,N_12649);
and U12807 (N_12807,N_12694,N_12601);
and U12808 (N_12808,N_12622,N_12684);
xor U12809 (N_12809,N_12686,N_12743);
nand U12810 (N_12810,N_12617,N_12693);
nor U12811 (N_12811,N_12682,N_12668);
and U12812 (N_12812,N_12742,N_12660);
xnor U12813 (N_12813,N_12657,N_12661);
nand U12814 (N_12814,N_12706,N_12709);
or U12815 (N_12815,N_12736,N_12632);
xor U12816 (N_12816,N_12681,N_12744);
and U12817 (N_12817,N_12608,N_12625);
nand U12818 (N_12818,N_12737,N_12721);
and U12819 (N_12819,N_12680,N_12712);
nand U12820 (N_12820,N_12666,N_12748);
or U12821 (N_12821,N_12610,N_12685);
nor U12822 (N_12822,N_12713,N_12600);
nand U12823 (N_12823,N_12664,N_12605);
and U12824 (N_12824,N_12616,N_12603);
and U12825 (N_12825,N_12600,N_12676);
nand U12826 (N_12826,N_12743,N_12672);
or U12827 (N_12827,N_12717,N_12681);
xnor U12828 (N_12828,N_12648,N_12658);
or U12829 (N_12829,N_12718,N_12615);
nor U12830 (N_12830,N_12629,N_12645);
nand U12831 (N_12831,N_12689,N_12713);
nand U12832 (N_12832,N_12737,N_12618);
and U12833 (N_12833,N_12679,N_12620);
nand U12834 (N_12834,N_12737,N_12654);
nand U12835 (N_12835,N_12673,N_12649);
nor U12836 (N_12836,N_12683,N_12643);
nand U12837 (N_12837,N_12632,N_12684);
or U12838 (N_12838,N_12635,N_12627);
xor U12839 (N_12839,N_12619,N_12616);
nor U12840 (N_12840,N_12680,N_12708);
nor U12841 (N_12841,N_12734,N_12678);
nor U12842 (N_12842,N_12731,N_12610);
nand U12843 (N_12843,N_12677,N_12672);
or U12844 (N_12844,N_12731,N_12683);
nor U12845 (N_12845,N_12624,N_12682);
xor U12846 (N_12846,N_12741,N_12652);
nand U12847 (N_12847,N_12627,N_12636);
or U12848 (N_12848,N_12743,N_12669);
and U12849 (N_12849,N_12650,N_12607);
nor U12850 (N_12850,N_12735,N_12711);
or U12851 (N_12851,N_12743,N_12649);
or U12852 (N_12852,N_12674,N_12650);
nand U12853 (N_12853,N_12723,N_12670);
or U12854 (N_12854,N_12716,N_12672);
or U12855 (N_12855,N_12664,N_12652);
or U12856 (N_12856,N_12730,N_12746);
and U12857 (N_12857,N_12613,N_12617);
and U12858 (N_12858,N_12670,N_12612);
nor U12859 (N_12859,N_12633,N_12604);
nor U12860 (N_12860,N_12647,N_12729);
nor U12861 (N_12861,N_12617,N_12610);
nor U12862 (N_12862,N_12618,N_12609);
xnor U12863 (N_12863,N_12747,N_12602);
nand U12864 (N_12864,N_12674,N_12705);
xnor U12865 (N_12865,N_12718,N_12730);
xnor U12866 (N_12866,N_12667,N_12728);
xor U12867 (N_12867,N_12671,N_12655);
or U12868 (N_12868,N_12624,N_12704);
or U12869 (N_12869,N_12601,N_12628);
xnor U12870 (N_12870,N_12693,N_12732);
nor U12871 (N_12871,N_12720,N_12628);
or U12872 (N_12872,N_12702,N_12707);
nand U12873 (N_12873,N_12681,N_12625);
nand U12874 (N_12874,N_12745,N_12705);
and U12875 (N_12875,N_12728,N_12696);
xor U12876 (N_12876,N_12641,N_12724);
nor U12877 (N_12877,N_12628,N_12704);
or U12878 (N_12878,N_12687,N_12673);
and U12879 (N_12879,N_12666,N_12639);
nor U12880 (N_12880,N_12719,N_12703);
xor U12881 (N_12881,N_12685,N_12733);
nand U12882 (N_12882,N_12609,N_12601);
and U12883 (N_12883,N_12653,N_12724);
xnor U12884 (N_12884,N_12625,N_12631);
nand U12885 (N_12885,N_12731,N_12733);
and U12886 (N_12886,N_12725,N_12654);
nor U12887 (N_12887,N_12654,N_12619);
or U12888 (N_12888,N_12743,N_12651);
nand U12889 (N_12889,N_12612,N_12716);
xnor U12890 (N_12890,N_12626,N_12742);
xor U12891 (N_12891,N_12654,N_12748);
nand U12892 (N_12892,N_12734,N_12647);
nand U12893 (N_12893,N_12696,N_12740);
or U12894 (N_12894,N_12661,N_12686);
xor U12895 (N_12895,N_12604,N_12624);
and U12896 (N_12896,N_12629,N_12684);
nor U12897 (N_12897,N_12639,N_12622);
and U12898 (N_12898,N_12623,N_12629);
and U12899 (N_12899,N_12673,N_12733);
xnor U12900 (N_12900,N_12835,N_12838);
xor U12901 (N_12901,N_12780,N_12881);
xnor U12902 (N_12902,N_12853,N_12788);
nor U12903 (N_12903,N_12766,N_12796);
and U12904 (N_12904,N_12759,N_12842);
or U12905 (N_12905,N_12870,N_12761);
nand U12906 (N_12906,N_12863,N_12809);
or U12907 (N_12907,N_12783,N_12807);
xnor U12908 (N_12908,N_12892,N_12804);
or U12909 (N_12909,N_12754,N_12793);
nand U12910 (N_12910,N_12779,N_12884);
nor U12911 (N_12911,N_12752,N_12841);
nand U12912 (N_12912,N_12786,N_12867);
or U12913 (N_12913,N_12785,N_12760);
nand U12914 (N_12914,N_12768,N_12802);
nor U12915 (N_12915,N_12828,N_12767);
nand U12916 (N_12916,N_12773,N_12826);
or U12917 (N_12917,N_12806,N_12897);
and U12918 (N_12918,N_12869,N_12814);
xor U12919 (N_12919,N_12883,N_12850);
nor U12920 (N_12920,N_12790,N_12891);
xor U12921 (N_12921,N_12758,N_12784);
and U12922 (N_12922,N_12778,N_12844);
xnor U12923 (N_12923,N_12827,N_12868);
nor U12924 (N_12924,N_12765,N_12839);
and U12925 (N_12925,N_12833,N_12840);
nor U12926 (N_12926,N_12820,N_12894);
or U12927 (N_12927,N_12857,N_12771);
xor U12928 (N_12928,N_12750,N_12887);
or U12929 (N_12929,N_12772,N_12871);
nand U12930 (N_12930,N_12782,N_12878);
or U12931 (N_12931,N_12817,N_12764);
and U12932 (N_12932,N_12866,N_12872);
nor U12933 (N_12933,N_12791,N_12873);
or U12934 (N_12934,N_12794,N_12856);
xnor U12935 (N_12935,N_12787,N_12812);
xnor U12936 (N_12936,N_12847,N_12803);
and U12937 (N_12937,N_12769,N_12799);
nand U12938 (N_12938,N_12819,N_12864);
and U12939 (N_12939,N_12755,N_12789);
and U12940 (N_12940,N_12829,N_12805);
and U12941 (N_12941,N_12824,N_12797);
nand U12942 (N_12942,N_12895,N_12899);
and U12943 (N_12943,N_12770,N_12822);
and U12944 (N_12944,N_12823,N_12886);
xor U12945 (N_12945,N_12821,N_12774);
and U12946 (N_12946,N_12811,N_12832);
nor U12947 (N_12947,N_12859,N_12825);
nor U12948 (N_12948,N_12815,N_12795);
xnor U12949 (N_12949,N_12831,N_12776);
or U12950 (N_12950,N_12756,N_12860);
or U12951 (N_12951,N_12851,N_12875);
nor U12952 (N_12952,N_12877,N_12816);
and U12953 (N_12953,N_12862,N_12818);
or U12954 (N_12954,N_12880,N_12876);
nand U12955 (N_12955,N_12893,N_12898);
nor U12956 (N_12956,N_12882,N_12849);
xor U12957 (N_12957,N_12848,N_12874);
or U12958 (N_12958,N_12879,N_12834);
or U12959 (N_12959,N_12753,N_12888);
or U12960 (N_12960,N_12830,N_12792);
nand U12961 (N_12961,N_12855,N_12810);
xnor U12962 (N_12962,N_12896,N_12843);
or U12963 (N_12963,N_12757,N_12845);
xor U12964 (N_12964,N_12781,N_12798);
nor U12965 (N_12965,N_12777,N_12858);
xnor U12966 (N_12966,N_12865,N_12890);
nor U12967 (N_12967,N_12800,N_12751);
nor U12968 (N_12968,N_12861,N_12775);
nor U12969 (N_12969,N_12846,N_12836);
and U12970 (N_12970,N_12854,N_12852);
xor U12971 (N_12971,N_12837,N_12885);
and U12972 (N_12972,N_12889,N_12808);
nand U12973 (N_12973,N_12762,N_12763);
and U12974 (N_12974,N_12813,N_12801);
nor U12975 (N_12975,N_12806,N_12811);
and U12976 (N_12976,N_12891,N_12828);
xnor U12977 (N_12977,N_12897,N_12792);
and U12978 (N_12978,N_12840,N_12885);
xnor U12979 (N_12979,N_12853,N_12859);
xnor U12980 (N_12980,N_12894,N_12818);
or U12981 (N_12981,N_12898,N_12813);
xnor U12982 (N_12982,N_12812,N_12840);
nor U12983 (N_12983,N_12816,N_12892);
xnor U12984 (N_12984,N_12839,N_12815);
nand U12985 (N_12985,N_12859,N_12796);
xnor U12986 (N_12986,N_12884,N_12866);
nand U12987 (N_12987,N_12755,N_12865);
and U12988 (N_12988,N_12803,N_12789);
nor U12989 (N_12989,N_12849,N_12780);
or U12990 (N_12990,N_12766,N_12783);
nor U12991 (N_12991,N_12870,N_12848);
nor U12992 (N_12992,N_12893,N_12791);
xor U12993 (N_12993,N_12760,N_12827);
or U12994 (N_12994,N_12795,N_12892);
or U12995 (N_12995,N_12830,N_12751);
xnor U12996 (N_12996,N_12776,N_12773);
or U12997 (N_12997,N_12827,N_12798);
and U12998 (N_12998,N_12773,N_12815);
or U12999 (N_12999,N_12802,N_12811);
or U13000 (N_13000,N_12782,N_12820);
and U13001 (N_13001,N_12772,N_12812);
xnor U13002 (N_13002,N_12865,N_12857);
xor U13003 (N_13003,N_12769,N_12791);
or U13004 (N_13004,N_12826,N_12837);
nand U13005 (N_13005,N_12819,N_12881);
or U13006 (N_13006,N_12875,N_12823);
xnor U13007 (N_13007,N_12863,N_12899);
or U13008 (N_13008,N_12873,N_12878);
xor U13009 (N_13009,N_12792,N_12815);
and U13010 (N_13010,N_12885,N_12850);
xnor U13011 (N_13011,N_12852,N_12895);
nand U13012 (N_13012,N_12815,N_12753);
and U13013 (N_13013,N_12826,N_12759);
nand U13014 (N_13014,N_12818,N_12765);
nor U13015 (N_13015,N_12792,N_12858);
nor U13016 (N_13016,N_12889,N_12768);
or U13017 (N_13017,N_12760,N_12780);
nor U13018 (N_13018,N_12797,N_12796);
xor U13019 (N_13019,N_12753,N_12854);
and U13020 (N_13020,N_12774,N_12894);
nor U13021 (N_13021,N_12764,N_12868);
xnor U13022 (N_13022,N_12849,N_12816);
nand U13023 (N_13023,N_12820,N_12860);
nor U13024 (N_13024,N_12844,N_12850);
nand U13025 (N_13025,N_12823,N_12761);
nor U13026 (N_13026,N_12870,N_12778);
nand U13027 (N_13027,N_12819,N_12860);
or U13028 (N_13028,N_12756,N_12870);
or U13029 (N_13029,N_12783,N_12888);
xnor U13030 (N_13030,N_12865,N_12754);
or U13031 (N_13031,N_12899,N_12826);
nor U13032 (N_13032,N_12780,N_12888);
xor U13033 (N_13033,N_12766,N_12765);
xnor U13034 (N_13034,N_12757,N_12894);
nand U13035 (N_13035,N_12854,N_12826);
xor U13036 (N_13036,N_12793,N_12845);
and U13037 (N_13037,N_12874,N_12860);
or U13038 (N_13038,N_12880,N_12765);
nand U13039 (N_13039,N_12837,N_12833);
or U13040 (N_13040,N_12817,N_12756);
nor U13041 (N_13041,N_12810,N_12877);
nor U13042 (N_13042,N_12783,N_12842);
nand U13043 (N_13043,N_12852,N_12885);
nor U13044 (N_13044,N_12843,N_12878);
and U13045 (N_13045,N_12794,N_12777);
and U13046 (N_13046,N_12824,N_12891);
nor U13047 (N_13047,N_12763,N_12774);
and U13048 (N_13048,N_12844,N_12776);
nor U13049 (N_13049,N_12767,N_12772);
and U13050 (N_13050,N_12935,N_13041);
nor U13051 (N_13051,N_12947,N_12986);
xnor U13052 (N_13052,N_12999,N_12954);
xor U13053 (N_13053,N_13029,N_12901);
and U13054 (N_13054,N_12932,N_13004);
nor U13055 (N_13055,N_12900,N_12943);
and U13056 (N_13056,N_13035,N_13018);
nand U13057 (N_13057,N_13000,N_13047);
and U13058 (N_13058,N_12916,N_12991);
nand U13059 (N_13059,N_13015,N_12993);
and U13060 (N_13060,N_12975,N_12973);
or U13061 (N_13061,N_13014,N_12974);
and U13062 (N_13062,N_12920,N_12960);
xor U13063 (N_13063,N_13009,N_13011);
or U13064 (N_13064,N_13010,N_13031);
and U13065 (N_13065,N_12915,N_12981);
or U13066 (N_13066,N_12917,N_12979);
nor U13067 (N_13067,N_12955,N_12976);
nor U13068 (N_13068,N_12992,N_12957);
nor U13069 (N_13069,N_13007,N_13001);
nor U13070 (N_13070,N_12950,N_13048);
and U13071 (N_13071,N_12940,N_13034);
xnor U13072 (N_13072,N_13006,N_12987);
nor U13073 (N_13073,N_12971,N_12908);
or U13074 (N_13074,N_13012,N_12951);
and U13075 (N_13075,N_12933,N_12968);
or U13076 (N_13076,N_13027,N_12998);
and U13077 (N_13077,N_13023,N_13013);
xnor U13078 (N_13078,N_12928,N_13042);
nor U13079 (N_13079,N_12913,N_12929);
nand U13080 (N_13080,N_13032,N_13016);
and U13081 (N_13081,N_12983,N_12907);
and U13082 (N_13082,N_12948,N_13039);
nand U13083 (N_13083,N_12994,N_12906);
nand U13084 (N_13084,N_12911,N_13002);
nor U13085 (N_13085,N_12966,N_12938);
or U13086 (N_13086,N_13038,N_12942);
or U13087 (N_13087,N_12980,N_12918);
xor U13088 (N_13088,N_12912,N_12910);
nor U13089 (N_13089,N_13017,N_12962);
or U13090 (N_13090,N_12958,N_12922);
nor U13091 (N_13091,N_12914,N_12924);
or U13092 (N_13092,N_12949,N_12967);
xnor U13093 (N_13093,N_12930,N_13024);
nor U13094 (N_13094,N_12970,N_12977);
or U13095 (N_13095,N_13036,N_12905);
or U13096 (N_13096,N_12946,N_13044);
nand U13097 (N_13097,N_12959,N_12969);
and U13098 (N_13098,N_13030,N_12989);
nand U13099 (N_13099,N_12936,N_13043);
xor U13100 (N_13100,N_12961,N_12904);
nor U13101 (N_13101,N_12921,N_13019);
xnor U13102 (N_13102,N_13028,N_13045);
xor U13103 (N_13103,N_12988,N_12984);
nor U13104 (N_13104,N_13021,N_12978);
nor U13105 (N_13105,N_12923,N_12941);
nor U13106 (N_13106,N_12952,N_12995);
and U13107 (N_13107,N_12903,N_12925);
nor U13108 (N_13108,N_12945,N_13046);
nor U13109 (N_13109,N_13022,N_12944);
xnor U13110 (N_13110,N_12937,N_13005);
xor U13111 (N_13111,N_12956,N_12964);
nand U13112 (N_13112,N_13049,N_12963);
or U13113 (N_13113,N_13008,N_12909);
xnor U13114 (N_13114,N_13026,N_13020);
or U13115 (N_13115,N_12982,N_12919);
or U13116 (N_13116,N_12927,N_12931);
nand U13117 (N_13117,N_12997,N_12965);
xnor U13118 (N_13118,N_13040,N_12972);
xnor U13119 (N_13119,N_12990,N_12996);
nor U13120 (N_13120,N_13003,N_13033);
and U13121 (N_13121,N_12985,N_12939);
and U13122 (N_13122,N_12926,N_12934);
xnor U13123 (N_13123,N_13025,N_12902);
nand U13124 (N_13124,N_13037,N_12953);
or U13125 (N_13125,N_12926,N_13036);
nand U13126 (N_13126,N_12922,N_12918);
or U13127 (N_13127,N_12959,N_13043);
nor U13128 (N_13128,N_13027,N_12949);
and U13129 (N_13129,N_12935,N_12958);
nor U13130 (N_13130,N_12900,N_12995);
nand U13131 (N_13131,N_12970,N_13003);
and U13132 (N_13132,N_12933,N_12950);
nand U13133 (N_13133,N_12920,N_12988);
nand U13134 (N_13134,N_13039,N_13037);
xnor U13135 (N_13135,N_13018,N_12951);
xor U13136 (N_13136,N_13047,N_12914);
nor U13137 (N_13137,N_12939,N_12918);
xor U13138 (N_13138,N_12979,N_12981);
or U13139 (N_13139,N_12993,N_12920);
xnor U13140 (N_13140,N_12925,N_12975);
or U13141 (N_13141,N_12957,N_13029);
xor U13142 (N_13142,N_13048,N_12915);
and U13143 (N_13143,N_13000,N_12979);
and U13144 (N_13144,N_12973,N_12911);
nor U13145 (N_13145,N_12956,N_13001);
nand U13146 (N_13146,N_13041,N_13002);
or U13147 (N_13147,N_12901,N_12937);
nand U13148 (N_13148,N_13039,N_12983);
and U13149 (N_13149,N_12936,N_12986);
nand U13150 (N_13150,N_12902,N_13000);
nor U13151 (N_13151,N_13024,N_13006);
nand U13152 (N_13152,N_12957,N_12917);
xnor U13153 (N_13153,N_12918,N_13023);
xnor U13154 (N_13154,N_12915,N_12991);
nand U13155 (N_13155,N_12958,N_12992);
and U13156 (N_13156,N_13042,N_12976);
nand U13157 (N_13157,N_13035,N_12958);
xnor U13158 (N_13158,N_12913,N_12979);
and U13159 (N_13159,N_13045,N_13000);
xor U13160 (N_13160,N_12988,N_13040);
nand U13161 (N_13161,N_12933,N_13035);
nor U13162 (N_13162,N_12981,N_12912);
nand U13163 (N_13163,N_12973,N_12919);
nand U13164 (N_13164,N_12953,N_12960);
xnor U13165 (N_13165,N_13037,N_12976);
nand U13166 (N_13166,N_12961,N_12973);
nor U13167 (N_13167,N_12906,N_13004);
nand U13168 (N_13168,N_12950,N_12943);
xnor U13169 (N_13169,N_12955,N_13029);
xnor U13170 (N_13170,N_13045,N_12991);
nand U13171 (N_13171,N_13023,N_12964);
xor U13172 (N_13172,N_13013,N_12959);
nand U13173 (N_13173,N_13025,N_12964);
xor U13174 (N_13174,N_12998,N_12937);
xnor U13175 (N_13175,N_12953,N_13040);
or U13176 (N_13176,N_12922,N_12959);
and U13177 (N_13177,N_12926,N_13044);
and U13178 (N_13178,N_12918,N_12971);
or U13179 (N_13179,N_12965,N_13013);
xnor U13180 (N_13180,N_13044,N_12985);
nor U13181 (N_13181,N_12981,N_13008);
or U13182 (N_13182,N_12967,N_12972);
nand U13183 (N_13183,N_12951,N_13002);
nand U13184 (N_13184,N_12984,N_12990);
or U13185 (N_13185,N_12950,N_12957);
nor U13186 (N_13186,N_12935,N_13044);
or U13187 (N_13187,N_12947,N_13042);
nor U13188 (N_13188,N_12988,N_12970);
nor U13189 (N_13189,N_13023,N_12963);
and U13190 (N_13190,N_13032,N_12998);
nand U13191 (N_13191,N_13014,N_13023);
xor U13192 (N_13192,N_12932,N_12936);
nand U13193 (N_13193,N_13046,N_13026);
nor U13194 (N_13194,N_13037,N_12921);
or U13195 (N_13195,N_12903,N_13006);
nand U13196 (N_13196,N_13041,N_12959);
and U13197 (N_13197,N_12913,N_12984);
or U13198 (N_13198,N_13018,N_12995);
xor U13199 (N_13199,N_12956,N_13045);
and U13200 (N_13200,N_13066,N_13069);
nor U13201 (N_13201,N_13158,N_13096);
or U13202 (N_13202,N_13073,N_13074);
or U13203 (N_13203,N_13160,N_13067);
xor U13204 (N_13204,N_13108,N_13175);
nand U13205 (N_13205,N_13087,N_13110);
xnor U13206 (N_13206,N_13093,N_13140);
nor U13207 (N_13207,N_13088,N_13195);
and U13208 (N_13208,N_13144,N_13085);
nand U13209 (N_13209,N_13097,N_13075);
nand U13210 (N_13210,N_13168,N_13135);
and U13211 (N_13211,N_13114,N_13132);
and U13212 (N_13212,N_13070,N_13105);
nand U13213 (N_13213,N_13141,N_13123);
or U13214 (N_13214,N_13167,N_13188);
or U13215 (N_13215,N_13174,N_13082);
and U13216 (N_13216,N_13180,N_13165);
or U13217 (N_13217,N_13111,N_13138);
nor U13218 (N_13218,N_13090,N_13112);
nand U13219 (N_13219,N_13189,N_13133);
and U13220 (N_13220,N_13072,N_13101);
or U13221 (N_13221,N_13117,N_13127);
and U13222 (N_13222,N_13078,N_13062);
xor U13223 (N_13223,N_13171,N_13061);
and U13224 (N_13224,N_13086,N_13058);
nand U13225 (N_13225,N_13169,N_13107);
xnor U13226 (N_13226,N_13193,N_13177);
or U13227 (N_13227,N_13084,N_13191);
xnor U13228 (N_13228,N_13130,N_13151);
nor U13229 (N_13229,N_13059,N_13183);
nand U13230 (N_13230,N_13197,N_13145);
or U13231 (N_13231,N_13190,N_13071);
nor U13232 (N_13232,N_13194,N_13053);
nand U13233 (N_13233,N_13116,N_13162);
nand U13234 (N_13234,N_13179,N_13124);
or U13235 (N_13235,N_13182,N_13060);
nand U13236 (N_13236,N_13054,N_13079);
and U13237 (N_13237,N_13121,N_13184);
nand U13238 (N_13238,N_13064,N_13198);
or U13239 (N_13239,N_13063,N_13125);
nand U13240 (N_13240,N_13081,N_13164);
xor U13241 (N_13241,N_13192,N_13159);
and U13242 (N_13242,N_13122,N_13154);
nor U13243 (N_13243,N_13094,N_13077);
nor U13244 (N_13244,N_13181,N_13118);
or U13245 (N_13245,N_13136,N_13152);
xor U13246 (N_13246,N_13068,N_13089);
nor U13247 (N_13247,N_13142,N_13128);
and U13248 (N_13248,N_13148,N_13137);
xnor U13249 (N_13249,N_13149,N_13050);
nor U13250 (N_13250,N_13157,N_13155);
or U13251 (N_13251,N_13143,N_13131);
nor U13252 (N_13252,N_13099,N_13095);
nor U13253 (N_13253,N_13120,N_13126);
or U13254 (N_13254,N_13163,N_13100);
nor U13255 (N_13255,N_13103,N_13109);
nand U13256 (N_13256,N_13166,N_13092);
and U13257 (N_13257,N_13134,N_13113);
or U13258 (N_13258,N_13057,N_13150);
xnor U13259 (N_13259,N_13076,N_13161);
xor U13260 (N_13260,N_13106,N_13178);
or U13261 (N_13261,N_13187,N_13119);
xor U13262 (N_13262,N_13052,N_13091);
and U13263 (N_13263,N_13146,N_13156);
and U13264 (N_13264,N_13098,N_13185);
nor U13265 (N_13265,N_13186,N_13147);
or U13266 (N_13266,N_13129,N_13065);
xnor U13267 (N_13267,N_13139,N_13102);
xnor U13268 (N_13268,N_13173,N_13104);
nor U13269 (N_13269,N_13172,N_13199);
xor U13270 (N_13270,N_13056,N_13115);
and U13271 (N_13271,N_13153,N_13176);
xor U13272 (N_13272,N_13055,N_13170);
or U13273 (N_13273,N_13083,N_13051);
xnor U13274 (N_13274,N_13080,N_13196);
or U13275 (N_13275,N_13069,N_13154);
nand U13276 (N_13276,N_13188,N_13067);
or U13277 (N_13277,N_13150,N_13157);
nand U13278 (N_13278,N_13059,N_13104);
nor U13279 (N_13279,N_13159,N_13103);
and U13280 (N_13280,N_13128,N_13052);
and U13281 (N_13281,N_13155,N_13075);
and U13282 (N_13282,N_13182,N_13061);
and U13283 (N_13283,N_13147,N_13134);
and U13284 (N_13284,N_13057,N_13072);
nand U13285 (N_13285,N_13153,N_13143);
and U13286 (N_13286,N_13054,N_13174);
and U13287 (N_13287,N_13094,N_13173);
nand U13288 (N_13288,N_13073,N_13122);
or U13289 (N_13289,N_13090,N_13103);
and U13290 (N_13290,N_13185,N_13176);
nor U13291 (N_13291,N_13197,N_13077);
nand U13292 (N_13292,N_13176,N_13069);
or U13293 (N_13293,N_13180,N_13157);
xor U13294 (N_13294,N_13133,N_13073);
and U13295 (N_13295,N_13117,N_13193);
xor U13296 (N_13296,N_13070,N_13189);
xor U13297 (N_13297,N_13099,N_13192);
and U13298 (N_13298,N_13158,N_13066);
and U13299 (N_13299,N_13167,N_13111);
and U13300 (N_13300,N_13106,N_13181);
xnor U13301 (N_13301,N_13132,N_13096);
xnor U13302 (N_13302,N_13130,N_13175);
nor U13303 (N_13303,N_13085,N_13112);
xnor U13304 (N_13304,N_13194,N_13162);
xor U13305 (N_13305,N_13161,N_13129);
or U13306 (N_13306,N_13144,N_13147);
xnor U13307 (N_13307,N_13188,N_13107);
xnor U13308 (N_13308,N_13149,N_13154);
nand U13309 (N_13309,N_13196,N_13147);
and U13310 (N_13310,N_13164,N_13181);
and U13311 (N_13311,N_13061,N_13084);
xor U13312 (N_13312,N_13170,N_13149);
xnor U13313 (N_13313,N_13157,N_13130);
or U13314 (N_13314,N_13189,N_13161);
or U13315 (N_13315,N_13122,N_13166);
nor U13316 (N_13316,N_13085,N_13088);
and U13317 (N_13317,N_13053,N_13107);
and U13318 (N_13318,N_13129,N_13146);
nand U13319 (N_13319,N_13092,N_13177);
and U13320 (N_13320,N_13160,N_13138);
and U13321 (N_13321,N_13073,N_13173);
or U13322 (N_13322,N_13172,N_13056);
nor U13323 (N_13323,N_13129,N_13111);
nor U13324 (N_13324,N_13158,N_13154);
or U13325 (N_13325,N_13064,N_13102);
xor U13326 (N_13326,N_13129,N_13198);
nor U13327 (N_13327,N_13146,N_13170);
xnor U13328 (N_13328,N_13198,N_13191);
nor U13329 (N_13329,N_13149,N_13141);
and U13330 (N_13330,N_13171,N_13192);
xor U13331 (N_13331,N_13078,N_13061);
nor U13332 (N_13332,N_13061,N_13196);
nand U13333 (N_13333,N_13080,N_13088);
nor U13334 (N_13334,N_13171,N_13168);
and U13335 (N_13335,N_13137,N_13102);
nor U13336 (N_13336,N_13062,N_13199);
xor U13337 (N_13337,N_13142,N_13067);
xor U13338 (N_13338,N_13195,N_13078);
or U13339 (N_13339,N_13108,N_13072);
xnor U13340 (N_13340,N_13175,N_13165);
or U13341 (N_13341,N_13112,N_13166);
nand U13342 (N_13342,N_13131,N_13070);
and U13343 (N_13343,N_13092,N_13180);
nor U13344 (N_13344,N_13190,N_13050);
nor U13345 (N_13345,N_13182,N_13050);
or U13346 (N_13346,N_13115,N_13186);
xor U13347 (N_13347,N_13076,N_13070);
or U13348 (N_13348,N_13137,N_13167);
nand U13349 (N_13349,N_13128,N_13179);
nand U13350 (N_13350,N_13309,N_13273);
or U13351 (N_13351,N_13227,N_13281);
nand U13352 (N_13352,N_13320,N_13234);
xor U13353 (N_13353,N_13235,N_13226);
and U13354 (N_13354,N_13339,N_13223);
nor U13355 (N_13355,N_13276,N_13271);
nor U13356 (N_13356,N_13253,N_13217);
or U13357 (N_13357,N_13241,N_13238);
and U13358 (N_13358,N_13325,N_13336);
nand U13359 (N_13359,N_13267,N_13247);
nand U13360 (N_13360,N_13305,N_13278);
or U13361 (N_13361,N_13214,N_13212);
and U13362 (N_13362,N_13261,N_13299);
xnor U13363 (N_13363,N_13264,N_13317);
or U13364 (N_13364,N_13222,N_13313);
or U13365 (N_13365,N_13295,N_13246);
or U13366 (N_13366,N_13286,N_13240);
and U13367 (N_13367,N_13330,N_13208);
nor U13368 (N_13368,N_13279,N_13230);
or U13369 (N_13369,N_13300,N_13314);
xnor U13370 (N_13370,N_13269,N_13291);
and U13371 (N_13371,N_13328,N_13204);
nand U13372 (N_13372,N_13304,N_13254);
or U13373 (N_13373,N_13292,N_13275);
xor U13374 (N_13374,N_13252,N_13256);
nand U13375 (N_13375,N_13329,N_13293);
and U13376 (N_13376,N_13285,N_13298);
xnor U13377 (N_13377,N_13262,N_13341);
or U13378 (N_13378,N_13216,N_13219);
and U13379 (N_13379,N_13348,N_13221);
and U13380 (N_13380,N_13337,N_13296);
nor U13381 (N_13381,N_13260,N_13282);
xor U13382 (N_13382,N_13251,N_13349);
xnor U13383 (N_13383,N_13302,N_13310);
xor U13384 (N_13384,N_13207,N_13255);
xor U13385 (N_13385,N_13259,N_13308);
and U13386 (N_13386,N_13268,N_13239);
nor U13387 (N_13387,N_13233,N_13283);
nor U13388 (N_13388,N_13290,N_13335);
nand U13389 (N_13389,N_13311,N_13345);
nor U13390 (N_13390,N_13323,N_13243);
or U13391 (N_13391,N_13306,N_13284);
xor U13392 (N_13392,N_13327,N_13200);
and U13393 (N_13393,N_13236,N_13312);
or U13394 (N_13394,N_13303,N_13245);
nand U13395 (N_13395,N_13242,N_13224);
nand U13396 (N_13396,N_13321,N_13244);
xor U13397 (N_13397,N_13294,N_13210);
and U13398 (N_13398,N_13334,N_13250);
nand U13399 (N_13399,N_13346,N_13316);
and U13400 (N_13400,N_13213,N_13287);
nand U13401 (N_13401,N_13266,N_13201);
or U13402 (N_13402,N_13326,N_13205);
and U13403 (N_13403,N_13249,N_13270);
and U13404 (N_13404,N_13215,N_13202);
nor U13405 (N_13405,N_13301,N_13225);
nand U13406 (N_13406,N_13322,N_13347);
and U13407 (N_13407,N_13277,N_13218);
nand U13408 (N_13408,N_13248,N_13280);
nand U13409 (N_13409,N_13265,N_13206);
nand U13410 (N_13410,N_13203,N_13307);
nor U13411 (N_13411,N_13257,N_13263);
xnor U13412 (N_13412,N_13220,N_13297);
nand U13413 (N_13413,N_13258,N_13289);
nand U13414 (N_13414,N_13318,N_13338);
nor U13415 (N_13415,N_13324,N_13340);
or U13416 (N_13416,N_13228,N_13231);
nor U13417 (N_13417,N_13331,N_13209);
and U13418 (N_13418,N_13274,N_13232);
and U13419 (N_13419,N_13315,N_13237);
or U13420 (N_13420,N_13211,N_13343);
nor U13421 (N_13421,N_13332,N_13272);
xnor U13422 (N_13422,N_13288,N_13319);
xnor U13423 (N_13423,N_13344,N_13229);
and U13424 (N_13424,N_13342,N_13333);
nor U13425 (N_13425,N_13206,N_13318);
and U13426 (N_13426,N_13205,N_13298);
nor U13427 (N_13427,N_13236,N_13296);
nand U13428 (N_13428,N_13243,N_13275);
and U13429 (N_13429,N_13327,N_13305);
and U13430 (N_13430,N_13234,N_13316);
and U13431 (N_13431,N_13230,N_13335);
and U13432 (N_13432,N_13261,N_13204);
or U13433 (N_13433,N_13319,N_13207);
and U13434 (N_13434,N_13273,N_13294);
and U13435 (N_13435,N_13300,N_13209);
nand U13436 (N_13436,N_13312,N_13278);
xor U13437 (N_13437,N_13349,N_13205);
nor U13438 (N_13438,N_13246,N_13276);
xnor U13439 (N_13439,N_13244,N_13308);
nand U13440 (N_13440,N_13254,N_13291);
or U13441 (N_13441,N_13312,N_13269);
or U13442 (N_13442,N_13247,N_13329);
and U13443 (N_13443,N_13283,N_13245);
nor U13444 (N_13444,N_13301,N_13203);
nor U13445 (N_13445,N_13282,N_13227);
nand U13446 (N_13446,N_13327,N_13340);
nand U13447 (N_13447,N_13249,N_13232);
or U13448 (N_13448,N_13234,N_13296);
xor U13449 (N_13449,N_13237,N_13225);
or U13450 (N_13450,N_13249,N_13330);
and U13451 (N_13451,N_13235,N_13295);
and U13452 (N_13452,N_13255,N_13276);
and U13453 (N_13453,N_13346,N_13260);
or U13454 (N_13454,N_13226,N_13263);
nor U13455 (N_13455,N_13250,N_13324);
and U13456 (N_13456,N_13310,N_13342);
xor U13457 (N_13457,N_13336,N_13204);
or U13458 (N_13458,N_13347,N_13331);
or U13459 (N_13459,N_13214,N_13292);
nor U13460 (N_13460,N_13221,N_13293);
xor U13461 (N_13461,N_13300,N_13205);
nand U13462 (N_13462,N_13221,N_13330);
nand U13463 (N_13463,N_13215,N_13259);
and U13464 (N_13464,N_13264,N_13296);
xnor U13465 (N_13465,N_13344,N_13220);
nor U13466 (N_13466,N_13281,N_13271);
xnor U13467 (N_13467,N_13278,N_13281);
xnor U13468 (N_13468,N_13206,N_13271);
xnor U13469 (N_13469,N_13251,N_13324);
and U13470 (N_13470,N_13245,N_13254);
xor U13471 (N_13471,N_13290,N_13339);
nand U13472 (N_13472,N_13316,N_13226);
and U13473 (N_13473,N_13260,N_13242);
xor U13474 (N_13474,N_13333,N_13237);
nand U13475 (N_13475,N_13327,N_13329);
xor U13476 (N_13476,N_13212,N_13270);
and U13477 (N_13477,N_13255,N_13204);
and U13478 (N_13478,N_13297,N_13265);
nand U13479 (N_13479,N_13336,N_13314);
or U13480 (N_13480,N_13326,N_13285);
xor U13481 (N_13481,N_13250,N_13329);
xnor U13482 (N_13482,N_13290,N_13300);
and U13483 (N_13483,N_13309,N_13290);
nor U13484 (N_13484,N_13342,N_13300);
xnor U13485 (N_13485,N_13330,N_13287);
and U13486 (N_13486,N_13338,N_13247);
nand U13487 (N_13487,N_13281,N_13292);
nand U13488 (N_13488,N_13251,N_13285);
xor U13489 (N_13489,N_13276,N_13226);
nor U13490 (N_13490,N_13244,N_13342);
nand U13491 (N_13491,N_13300,N_13267);
or U13492 (N_13492,N_13238,N_13248);
nor U13493 (N_13493,N_13336,N_13297);
xnor U13494 (N_13494,N_13258,N_13250);
xnor U13495 (N_13495,N_13269,N_13258);
xor U13496 (N_13496,N_13327,N_13236);
nand U13497 (N_13497,N_13249,N_13254);
and U13498 (N_13498,N_13201,N_13271);
and U13499 (N_13499,N_13263,N_13270);
nor U13500 (N_13500,N_13388,N_13489);
nor U13501 (N_13501,N_13427,N_13373);
xor U13502 (N_13502,N_13446,N_13462);
nand U13503 (N_13503,N_13366,N_13405);
nor U13504 (N_13504,N_13494,N_13412);
or U13505 (N_13505,N_13479,N_13417);
or U13506 (N_13506,N_13485,N_13374);
xnor U13507 (N_13507,N_13466,N_13456);
xnor U13508 (N_13508,N_13472,N_13480);
xnor U13509 (N_13509,N_13357,N_13378);
xor U13510 (N_13510,N_13381,N_13395);
and U13511 (N_13511,N_13419,N_13368);
or U13512 (N_13512,N_13415,N_13454);
nand U13513 (N_13513,N_13413,N_13450);
nand U13514 (N_13514,N_13400,N_13396);
xnor U13515 (N_13515,N_13430,N_13362);
nand U13516 (N_13516,N_13445,N_13451);
nor U13517 (N_13517,N_13393,N_13380);
and U13518 (N_13518,N_13499,N_13474);
or U13519 (N_13519,N_13401,N_13429);
and U13520 (N_13520,N_13487,N_13354);
nand U13521 (N_13521,N_13421,N_13464);
or U13522 (N_13522,N_13467,N_13409);
or U13523 (N_13523,N_13498,N_13492);
or U13524 (N_13524,N_13438,N_13434);
xnor U13525 (N_13525,N_13377,N_13390);
and U13526 (N_13526,N_13441,N_13496);
and U13527 (N_13527,N_13414,N_13359);
and U13528 (N_13528,N_13455,N_13444);
nor U13529 (N_13529,N_13387,N_13481);
and U13530 (N_13530,N_13458,N_13365);
nand U13531 (N_13531,N_13392,N_13351);
xnor U13532 (N_13532,N_13482,N_13469);
nor U13533 (N_13533,N_13397,N_13404);
and U13534 (N_13534,N_13361,N_13440);
nand U13535 (N_13535,N_13426,N_13453);
nor U13536 (N_13536,N_13411,N_13422);
or U13537 (N_13537,N_13473,N_13352);
and U13538 (N_13538,N_13486,N_13358);
nor U13539 (N_13539,N_13355,N_13431);
nand U13540 (N_13540,N_13384,N_13398);
xor U13541 (N_13541,N_13428,N_13371);
nand U13542 (N_13542,N_13463,N_13363);
and U13543 (N_13543,N_13442,N_13461);
and U13544 (N_13544,N_13457,N_13459);
or U13545 (N_13545,N_13493,N_13350);
xor U13546 (N_13546,N_13386,N_13448);
nor U13547 (N_13547,N_13407,N_13491);
nor U13548 (N_13548,N_13471,N_13484);
or U13549 (N_13549,N_13402,N_13490);
nand U13550 (N_13550,N_13399,N_13364);
nand U13551 (N_13551,N_13383,N_13391);
and U13552 (N_13552,N_13475,N_13423);
nor U13553 (N_13553,N_13425,N_13452);
nand U13554 (N_13554,N_13372,N_13360);
xor U13555 (N_13555,N_13476,N_13443);
xnor U13556 (N_13556,N_13389,N_13436);
and U13557 (N_13557,N_13483,N_13416);
or U13558 (N_13558,N_13447,N_13370);
and U13559 (N_13559,N_13420,N_13356);
xor U13560 (N_13560,N_13424,N_13433);
nand U13561 (N_13561,N_13470,N_13468);
and U13562 (N_13562,N_13488,N_13497);
and U13563 (N_13563,N_13403,N_13495);
and U13564 (N_13564,N_13375,N_13369);
and U13565 (N_13565,N_13410,N_13394);
or U13566 (N_13566,N_13449,N_13408);
or U13567 (N_13567,N_13385,N_13353);
or U13568 (N_13568,N_13406,N_13376);
xnor U13569 (N_13569,N_13367,N_13418);
xnor U13570 (N_13570,N_13379,N_13477);
nand U13571 (N_13571,N_13382,N_13435);
and U13572 (N_13572,N_13460,N_13478);
or U13573 (N_13573,N_13432,N_13437);
and U13574 (N_13574,N_13465,N_13439);
and U13575 (N_13575,N_13353,N_13417);
nand U13576 (N_13576,N_13358,N_13411);
or U13577 (N_13577,N_13408,N_13470);
nand U13578 (N_13578,N_13363,N_13450);
nand U13579 (N_13579,N_13458,N_13371);
or U13580 (N_13580,N_13479,N_13494);
xnor U13581 (N_13581,N_13386,N_13380);
nor U13582 (N_13582,N_13371,N_13474);
or U13583 (N_13583,N_13394,N_13472);
nand U13584 (N_13584,N_13355,N_13481);
or U13585 (N_13585,N_13423,N_13465);
xor U13586 (N_13586,N_13474,N_13437);
nand U13587 (N_13587,N_13463,N_13429);
or U13588 (N_13588,N_13446,N_13359);
xnor U13589 (N_13589,N_13387,N_13439);
or U13590 (N_13590,N_13446,N_13457);
nor U13591 (N_13591,N_13430,N_13467);
xor U13592 (N_13592,N_13440,N_13461);
and U13593 (N_13593,N_13421,N_13489);
nor U13594 (N_13594,N_13407,N_13467);
nand U13595 (N_13595,N_13363,N_13402);
nor U13596 (N_13596,N_13478,N_13441);
nand U13597 (N_13597,N_13370,N_13475);
xnor U13598 (N_13598,N_13433,N_13456);
xnor U13599 (N_13599,N_13480,N_13360);
xnor U13600 (N_13600,N_13364,N_13446);
or U13601 (N_13601,N_13405,N_13401);
and U13602 (N_13602,N_13367,N_13353);
and U13603 (N_13603,N_13431,N_13432);
xnor U13604 (N_13604,N_13396,N_13437);
nor U13605 (N_13605,N_13386,N_13389);
and U13606 (N_13606,N_13431,N_13449);
and U13607 (N_13607,N_13428,N_13441);
or U13608 (N_13608,N_13477,N_13457);
or U13609 (N_13609,N_13375,N_13423);
or U13610 (N_13610,N_13425,N_13431);
and U13611 (N_13611,N_13369,N_13379);
and U13612 (N_13612,N_13479,N_13459);
nor U13613 (N_13613,N_13447,N_13367);
and U13614 (N_13614,N_13496,N_13360);
xor U13615 (N_13615,N_13437,N_13469);
or U13616 (N_13616,N_13374,N_13441);
nor U13617 (N_13617,N_13392,N_13472);
nor U13618 (N_13618,N_13438,N_13468);
and U13619 (N_13619,N_13456,N_13441);
nor U13620 (N_13620,N_13397,N_13388);
or U13621 (N_13621,N_13471,N_13391);
nor U13622 (N_13622,N_13374,N_13464);
nor U13623 (N_13623,N_13464,N_13357);
and U13624 (N_13624,N_13487,N_13414);
or U13625 (N_13625,N_13429,N_13423);
xor U13626 (N_13626,N_13421,N_13468);
and U13627 (N_13627,N_13466,N_13379);
xnor U13628 (N_13628,N_13430,N_13464);
nand U13629 (N_13629,N_13483,N_13434);
or U13630 (N_13630,N_13498,N_13470);
or U13631 (N_13631,N_13355,N_13451);
xor U13632 (N_13632,N_13465,N_13472);
or U13633 (N_13633,N_13360,N_13466);
nand U13634 (N_13634,N_13450,N_13400);
and U13635 (N_13635,N_13423,N_13359);
and U13636 (N_13636,N_13444,N_13488);
xnor U13637 (N_13637,N_13364,N_13370);
nand U13638 (N_13638,N_13406,N_13411);
nand U13639 (N_13639,N_13477,N_13485);
nand U13640 (N_13640,N_13364,N_13418);
xnor U13641 (N_13641,N_13388,N_13429);
nor U13642 (N_13642,N_13475,N_13390);
xnor U13643 (N_13643,N_13474,N_13388);
and U13644 (N_13644,N_13486,N_13384);
nor U13645 (N_13645,N_13408,N_13378);
or U13646 (N_13646,N_13477,N_13476);
nand U13647 (N_13647,N_13482,N_13389);
nand U13648 (N_13648,N_13425,N_13405);
and U13649 (N_13649,N_13356,N_13454);
or U13650 (N_13650,N_13642,N_13511);
nand U13651 (N_13651,N_13503,N_13570);
nand U13652 (N_13652,N_13524,N_13633);
nand U13653 (N_13653,N_13552,N_13521);
and U13654 (N_13654,N_13558,N_13530);
nor U13655 (N_13655,N_13506,N_13621);
nand U13656 (N_13656,N_13584,N_13575);
or U13657 (N_13657,N_13646,N_13630);
or U13658 (N_13658,N_13618,N_13590);
nor U13659 (N_13659,N_13612,N_13588);
nor U13660 (N_13660,N_13611,N_13632);
or U13661 (N_13661,N_13510,N_13565);
or U13662 (N_13662,N_13581,N_13539);
and U13663 (N_13663,N_13540,N_13609);
and U13664 (N_13664,N_13616,N_13631);
and U13665 (N_13665,N_13537,N_13500);
and U13666 (N_13666,N_13545,N_13567);
nor U13667 (N_13667,N_13624,N_13534);
xnor U13668 (N_13668,N_13580,N_13577);
and U13669 (N_13669,N_13514,N_13525);
nand U13670 (N_13670,N_13505,N_13512);
nor U13671 (N_13671,N_13643,N_13628);
nand U13672 (N_13672,N_13576,N_13555);
or U13673 (N_13673,N_13535,N_13625);
nor U13674 (N_13674,N_13594,N_13509);
nand U13675 (N_13675,N_13639,N_13605);
xor U13676 (N_13676,N_13585,N_13599);
nand U13677 (N_13677,N_13572,N_13635);
or U13678 (N_13678,N_13610,N_13620);
or U13679 (N_13679,N_13607,N_13551);
or U13680 (N_13680,N_13517,N_13533);
nand U13681 (N_13681,N_13638,N_13531);
nor U13682 (N_13682,N_13579,N_13546);
or U13683 (N_13683,N_13574,N_13566);
xor U13684 (N_13684,N_13544,N_13507);
nand U13685 (N_13685,N_13637,N_13562);
and U13686 (N_13686,N_13563,N_13549);
xor U13687 (N_13687,N_13522,N_13541);
or U13688 (N_13688,N_13513,N_13629);
nand U13689 (N_13689,N_13649,N_13583);
nor U13690 (N_13690,N_13564,N_13501);
or U13691 (N_13691,N_13619,N_13593);
nor U13692 (N_13692,N_13557,N_13543);
and U13693 (N_13693,N_13613,N_13634);
or U13694 (N_13694,N_13520,N_13606);
or U13695 (N_13695,N_13603,N_13527);
nor U13696 (N_13696,N_13602,N_13538);
xnor U13697 (N_13697,N_13586,N_13515);
or U13698 (N_13698,N_13554,N_13578);
nand U13699 (N_13699,N_13589,N_13571);
xor U13700 (N_13700,N_13548,N_13640);
and U13701 (N_13701,N_13601,N_13647);
xnor U13702 (N_13702,N_13597,N_13626);
and U13703 (N_13703,N_13542,N_13623);
nor U13704 (N_13704,N_13559,N_13556);
or U13705 (N_13705,N_13504,N_13617);
and U13706 (N_13706,N_13519,N_13645);
and U13707 (N_13707,N_13636,N_13615);
nor U13708 (N_13708,N_13532,N_13604);
xnor U13709 (N_13709,N_13596,N_13516);
xnor U13710 (N_13710,N_13560,N_13561);
nand U13711 (N_13711,N_13627,N_13582);
xor U13712 (N_13712,N_13568,N_13518);
nand U13713 (N_13713,N_13553,N_13595);
nand U13714 (N_13714,N_13608,N_13508);
nand U13715 (N_13715,N_13591,N_13523);
or U13716 (N_13716,N_13529,N_13547);
nor U13717 (N_13717,N_13573,N_13648);
nand U13718 (N_13718,N_13550,N_13587);
xnor U13719 (N_13719,N_13526,N_13502);
xnor U13720 (N_13720,N_13536,N_13622);
nand U13721 (N_13721,N_13569,N_13528);
and U13722 (N_13722,N_13600,N_13641);
or U13723 (N_13723,N_13592,N_13598);
nor U13724 (N_13724,N_13644,N_13614);
or U13725 (N_13725,N_13547,N_13598);
or U13726 (N_13726,N_13525,N_13531);
nand U13727 (N_13727,N_13575,N_13601);
or U13728 (N_13728,N_13593,N_13527);
and U13729 (N_13729,N_13548,N_13578);
or U13730 (N_13730,N_13547,N_13637);
xor U13731 (N_13731,N_13508,N_13563);
nor U13732 (N_13732,N_13513,N_13620);
nand U13733 (N_13733,N_13520,N_13523);
nand U13734 (N_13734,N_13521,N_13525);
and U13735 (N_13735,N_13553,N_13542);
and U13736 (N_13736,N_13508,N_13575);
or U13737 (N_13737,N_13606,N_13555);
nand U13738 (N_13738,N_13636,N_13591);
or U13739 (N_13739,N_13617,N_13544);
nor U13740 (N_13740,N_13515,N_13605);
and U13741 (N_13741,N_13521,N_13580);
xnor U13742 (N_13742,N_13599,N_13561);
and U13743 (N_13743,N_13589,N_13615);
nand U13744 (N_13744,N_13532,N_13599);
xnor U13745 (N_13745,N_13629,N_13618);
nor U13746 (N_13746,N_13586,N_13543);
and U13747 (N_13747,N_13626,N_13578);
or U13748 (N_13748,N_13618,N_13565);
nand U13749 (N_13749,N_13506,N_13635);
and U13750 (N_13750,N_13522,N_13613);
nor U13751 (N_13751,N_13638,N_13544);
and U13752 (N_13752,N_13531,N_13502);
or U13753 (N_13753,N_13578,N_13513);
or U13754 (N_13754,N_13541,N_13507);
nor U13755 (N_13755,N_13540,N_13542);
nand U13756 (N_13756,N_13590,N_13548);
nor U13757 (N_13757,N_13577,N_13501);
nor U13758 (N_13758,N_13607,N_13624);
nor U13759 (N_13759,N_13521,N_13534);
and U13760 (N_13760,N_13550,N_13553);
and U13761 (N_13761,N_13510,N_13519);
or U13762 (N_13762,N_13626,N_13573);
and U13763 (N_13763,N_13610,N_13595);
and U13764 (N_13764,N_13598,N_13557);
nand U13765 (N_13765,N_13567,N_13601);
xor U13766 (N_13766,N_13598,N_13531);
or U13767 (N_13767,N_13645,N_13563);
nand U13768 (N_13768,N_13538,N_13513);
or U13769 (N_13769,N_13532,N_13574);
nor U13770 (N_13770,N_13579,N_13594);
nor U13771 (N_13771,N_13524,N_13591);
nand U13772 (N_13772,N_13571,N_13555);
xnor U13773 (N_13773,N_13576,N_13637);
xor U13774 (N_13774,N_13602,N_13535);
or U13775 (N_13775,N_13557,N_13532);
or U13776 (N_13776,N_13542,N_13514);
or U13777 (N_13777,N_13564,N_13517);
nor U13778 (N_13778,N_13516,N_13553);
and U13779 (N_13779,N_13549,N_13538);
nand U13780 (N_13780,N_13538,N_13633);
and U13781 (N_13781,N_13629,N_13614);
nor U13782 (N_13782,N_13579,N_13538);
nor U13783 (N_13783,N_13617,N_13562);
nor U13784 (N_13784,N_13621,N_13602);
xnor U13785 (N_13785,N_13578,N_13596);
and U13786 (N_13786,N_13560,N_13565);
nand U13787 (N_13787,N_13500,N_13521);
nand U13788 (N_13788,N_13533,N_13637);
xor U13789 (N_13789,N_13646,N_13556);
or U13790 (N_13790,N_13552,N_13561);
and U13791 (N_13791,N_13587,N_13564);
nor U13792 (N_13792,N_13500,N_13505);
nand U13793 (N_13793,N_13638,N_13575);
and U13794 (N_13794,N_13623,N_13564);
xnor U13795 (N_13795,N_13602,N_13590);
nand U13796 (N_13796,N_13591,N_13604);
and U13797 (N_13797,N_13638,N_13599);
or U13798 (N_13798,N_13649,N_13556);
and U13799 (N_13799,N_13614,N_13577);
or U13800 (N_13800,N_13691,N_13749);
or U13801 (N_13801,N_13651,N_13757);
nor U13802 (N_13802,N_13735,N_13718);
xor U13803 (N_13803,N_13728,N_13668);
xor U13804 (N_13804,N_13688,N_13736);
or U13805 (N_13805,N_13710,N_13766);
xnor U13806 (N_13806,N_13698,N_13670);
nor U13807 (N_13807,N_13732,N_13741);
or U13808 (N_13808,N_13661,N_13756);
xnor U13809 (N_13809,N_13733,N_13798);
or U13810 (N_13810,N_13679,N_13775);
and U13811 (N_13811,N_13799,N_13752);
xor U13812 (N_13812,N_13794,N_13774);
and U13813 (N_13813,N_13784,N_13764);
or U13814 (N_13814,N_13695,N_13716);
nor U13815 (N_13815,N_13650,N_13797);
nand U13816 (N_13816,N_13707,N_13771);
and U13817 (N_13817,N_13719,N_13754);
nor U13818 (N_13818,N_13653,N_13705);
and U13819 (N_13819,N_13682,N_13782);
nor U13820 (N_13820,N_13656,N_13663);
nand U13821 (N_13821,N_13660,N_13755);
or U13822 (N_13822,N_13753,N_13795);
and U13823 (N_13823,N_13681,N_13672);
nor U13824 (N_13824,N_13720,N_13700);
and U13825 (N_13825,N_13747,N_13742);
nand U13826 (N_13826,N_13690,N_13748);
and U13827 (N_13827,N_13772,N_13675);
nor U13828 (N_13828,N_13669,N_13791);
nand U13829 (N_13829,N_13738,N_13743);
nand U13830 (N_13830,N_13777,N_13779);
nor U13831 (N_13831,N_13652,N_13740);
nor U13832 (N_13832,N_13677,N_13667);
xnor U13833 (N_13833,N_13796,N_13788);
nand U13834 (N_13834,N_13671,N_13760);
or U13835 (N_13835,N_13726,N_13783);
nor U13836 (N_13836,N_13759,N_13664);
nand U13837 (N_13837,N_13765,N_13725);
xor U13838 (N_13838,N_13686,N_13712);
or U13839 (N_13839,N_13739,N_13790);
nor U13840 (N_13840,N_13704,N_13744);
or U13841 (N_13841,N_13693,N_13711);
or U13842 (N_13842,N_13768,N_13709);
or U13843 (N_13843,N_13708,N_13734);
or U13844 (N_13844,N_13657,N_13792);
nor U13845 (N_13845,N_13659,N_13713);
and U13846 (N_13846,N_13751,N_13787);
or U13847 (N_13847,N_13723,N_13699);
xor U13848 (N_13848,N_13745,N_13666);
nand U13849 (N_13849,N_13750,N_13694);
nor U13850 (N_13850,N_13778,N_13654);
and U13851 (N_13851,N_13689,N_13767);
nand U13852 (N_13852,N_13769,N_13702);
or U13853 (N_13853,N_13746,N_13714);
or U13854 (N_13854,N_13665,N_13685);
or U13855 (N_13855,N_13697,N_13762);
nor U13856 (N_13856,N_13658,N_13729);
and U13857 (N_13857,N_13722,N_13684);
or U13858 (N_13858,N_13696,N_13701);
xnor U13859 (N_13859,N_13773,N_13776);
nor U13860 (N_13860,N_13678,N_13731);
or U13861 (N_13861,N_13724,N_13715);
or U13862 (N_13862,N_13662,N_13676);
nand U13863 (N_13863,N_13770,N_13687);
nor U13864 (N_13864,N_13680,N_13692);
nand U13865 (N_13865,N_13673,N_13703);
and U13866 (N_13866,N_13717,N_13758);
nand U13867 (N_13867,N_13789,N_13721);
nor U13868 (N_13868,N_13727,N_13781);
or U13869 (N_13869,N_13730,N_13780);
nand U13870 (N_13870,N_13763,N_13785);
or U13871 (N_13871,N_13737,N_13761);
xnor U13872 (N_13872,N_13655,N_13793);
or U13873 (N_13873,N_13683,N_13786);
nor U13874 (N_13874,N_13706,N_13674);
or U13875 (N_13875,N_13690,N_13695);
or U13876 (N_13876,N_13753,N_13758);
nor U13877 (N_13877,N_13745,N_13698);
nand U13878 (N_13878,N_13769,N_13747);
xor U13879 (N_13879,N_13668,N_13799);
and U13880 (N_13880,N_13761,N_13660);
or U13881 (N_13881,N_13686,N_13796);
or U13882 (N_13882,N_13734,N_13777);
and U13883 (N_13883,N_13677,N_13741);
nor U13884 (N_13884,N_13768,N_13706);
nand U13885 (N_13885,N_13763,N_13667);
nor U13886 (N_13886,N_13786,N_13769);
and U13887 (N_13887,N_13686,N_13776);
nand U13888 (N_13888,N_13743,N_13681);
nand U13889 (N_13889,N_13688,N_13738);
nand U13890 (N_13890,N_13667,N_13742);
or U13891 (N_13891,N_13679,N_13779);
nor U13892 (N_13892,N_13679,N_13652);
xor U13893 (N_13893,N_13768,N_13798);
nand U13894 (N_13894,N_13777,N_13765);
and U13895 (N_13895,N_13715,N_13791);
nor U13896 (N_13896,N_13704,N_13691);
and U13897 (N_13897,N_13772,N_13769);
nor U13898 (N_13898,N_13675,N_13746);
and U13899 (N_13899,N_13733,N_13790);
nor U13900 (N_13900,N_13697,N_13792);
and U13901 (N_13901,N_13659,N_13789);
xor U13902 (N_13902,N_13718,N_13776);
and U13903 (N_13903,N_13703,N_13662);
and U13904 (N_13904,N_13745,N_13711);
nor U13905 (N_13905,N_13786,N_13700);
nand U13906 (N_13906,N_13763,N_13746);
and U13907 (N_13907,N_13669,N_13799);
xor U13908 (N_13908,N_13796,N_13671);
and U13909 (N_13909,N_13653,N_13771);
xor U13910 (N_13910,N_13781,N_13766);
nand U13911 (N_13911,N_13658,N_13670);
or U13912 (N_13912,N_13661,N_13784);
or U13913 (N_13913,N_13695,N_13739);
or U13914 (N_13914,N_13744,N_13796);
nor U13915 (N_13915,N_13779,N_13685);
and U13916 (N_13916,N_13659,N_13703);
xnor U13917 (N_13917,N_13676,N_13733);
nand U13918 (N_13918,N_13692,N_13761);
xor U13919 (N_13919,N_13665,N_13666);
and U13920 (N_13920,N_13721,N_13687);
xor U13921 (N_13921,N_13698,N_13673);
xnor U13922 (N_13922,N_13686,N_13677);
xor U13923 (N_13923,N_13792,N_13673);
and U13924 (N_13924,N_13734,N_13736);
and U13925 (N_13925,N_13732,N_13728);
xor U13926 (N_13926,N_13717,N_13795);
nor U13927 (N_13927,N_13786,N_13776);
xnor U13928 (N_13928,N_13792,N_13767);
nand U13929 (N_13929,N_13785,N_13661);
and U13930 (N_13930,N_13749,N_13791);
nor U13931 (N_13931,N_13702,N_13662);
nand U13932 (N_13932,N_13696,N_13650);
nand U13933 (N_13933,N_13706,N_13694);
xnor U13934 (N_13934,N_13766,N_13733);
and U13935 (N_13935,N_13793,N_13702);
or U13936 (N_13936,N_13757,N_13766);
xnor U13937 (N_13937,N_13650,N_13704);
or U13938 (N_13938,N_13722,N_13740);
and U13939 (N_13939,N_13674,N_13787);
or U13940 (N_13940,N_13673,N_13701);
and U13941 (N_13941,N_13738,N_13770);
xor U13942 (N_13942,N_13795,N_13784);
nor U13943 (N_13943,N_13757,N_13765);
nand U13944 (N_13944,N_13669,N_13690);
and U13945 (N_13945,N_13735,N_13760);
xor U13946 (N_13946,N_13779,N_13713);
or U13947 (N_13947,N_13738,N_13672);
and U13948 (N_13948,N_13679,N_13663);
nor U13949 (N_13949,N_13657,N_13751);
or U13950 (N_13950,N_13883,N_13910);
nand U13951 (N_13951,N_13949,N_13847);
xnor U13952 (N_13952,N_13853,N_13826);
xor U13953 (N_13953,N_13888,N_13899);
nor U13954 (N_13954,N_13934,N_13931);
nor U13955 (N_13955,N_13900,N_13838);
or U13956 (N_13956,N_13917,N_13856);
nand U13957 (N_13957,N_13803,N_13844);
or U13958 (N_13958,N_13862,N_13897);
and U13959 (N_13959,N_13874,N_13894);
nand U13960 (N_13960,N_13850,N_13808);
nor U13961 (N_13961,N_13896,N_13869);
and U13962 (N_13962,N_13928,N_13807);
nand U13963 (N_13963,N_13851,N_13833);
and U13964 (N_13964,N_13867,N_13906);
nand U13965 (N_13965,N_13938,N_13812);
or U13966 (N_13966,N_13865,N_13944);
or U13967 (N_13967,N_13872,N_13884);
nand U13968 (N_13968,N_13891,N_13834);
and U13969 (N_13969,N_13854,N_13889);
nand U13970 (N_13970,N_13945,N_13887);
nor U13971 (N_13971,N_13827,N_13947);
xor U13972 (N_13972,N_13840,N_13846);
nor U13973 (N_13973,N_13886,N_13805);
nand U13974 (N_13974,N_13809,N_13904);
nor U13975 (N_13975,N_13914,N_13881);
nor U13976 (N_13976,N_13801,N_13836);
xnor U13977 (N_13977,N_13948,N_13913);
or U13978 (N_13978,N_13929,N_13818);
nor U13979 (N_13979,N_13813,N_13939);
and U13980 (N_13980,N_13873,N_13823);
nor U13981 (N_13981,N_13911,N_13860);
xor U13982 (N_13982,N_13879,N_13898);
or U13983 (N_13983,N_13920,N_13880);
xor U13984 (N_13984,N_13863,N_13864);
nand U13985 (N_13985,N_13901,N_13909);
nor U13986 (N_13986,N_13936,N_13830);
or U13987 (N_13987,N_13903,N_13877);
nor U13988 (N_13988,N_13811,N_13822);
xor U13989 (N_13989,N_13814,N_13802);
nor U13990 (N_13990,N_13915,N_13905);
or U13991 (N_13991,N_13942,N_13892);
nand U13992 (N_13992,N_13878,N_13876);
and U13993 (N_13993,N_13875,N_13848);
nand U13994 (N_13994,N_13871,N_13849);
nand U13995 (N_13995,N_13837,N_13916);
nor U13996 (N_13996,N_13890,N_13868);
nand U13997 (N_13997,N_13933,N_13800);
or U13998 (N_13998,N_13882,N_13923);
or U13999 (N_13999,N_13921,N_13843);
xor U14000 (N_14000,N_13918,N_13816);
or U14001 (N_14001,N_13922,N_13820);
or U14002 (N_14002,N_13912,N_13857);
nand U14003 (N_14003,N_13815,N_13852);
xor U14004 (N_14004,N_13832,N_13946);
xnor U14005 (N_14005,N_13919,N_13937);
nor U14006 (N_14006,N_13866,N_13902);
xnor U14007 (N_14007,N_13858,N_13855);
or U14008 (N_14008,N_13925,N_13806);
nor U14009 (N_14009,N_13845,N_13829);
xnor U14010 (N_14010,N_13907,N_13841);
nor U14011 (N_14011,N_13824,N_13821);
nor U14012 (N_14012,N_13940,N_13804);
nand U14013 (N_14013,N_13828,N_13825);
nand U14014 (N_14014,N_13893,N_13895);
xor U14015 (N_14015,N_13842,N_13908);
or U14016 (N_14016,N_13810,N_13819);
nand U14017 (N_14017,N_13861,N_13932);
or U14018 (N_14018,N_13835,N_13831);
nor U14019 (N_14019,N_13926,N_13924);
or U14020 (N_14020,N_13941,N_13930);
nor U14021 (N_14021,N_13943,N_13935);
and U14022 (N_14022,N_13859,N_13927);
or U14023 (N_14023,N_13817,N_13870);
nand U14024 (N_14024,N_13885,N_13839);
xor U14025 (N_14025,N_13898,N_13826);
or U14026 (N_14026,N_13907,N_13822);
xor U14027 (N_14027,N_13812,N_13870);
xnor U14028 (N_14028,N_13876,N_13812);
and U14029 (N_14029,N_13863,N_13855);
nor U14030 (N_14030,N_13843,N_13890);
or U14031 (N_14031,N_13803,N_13828);
nor U14032 (N_14032,N_13821,N_13915);
and U14033 (N_14033,N_13905,N_13865);
nor U14034 (N_14034,N_13940,N_13854);
xor U14035 (N_14035,N_13927,N_13821);
nor U14036 (N_14036,N_13871,N_13876);
nand U14037 (N_14037,N_13891,N_13848);
xnor U14038 (N_14038,N_13835,N_13815);
nor U14039 (N_14039,N_13918,N_13937);
nand U14040 (N_14040,N_13904,N_13940);
and U14041 (N_14041,N_13804,N_13875);
xnor U14042 (N_14042,N_13938,N_13829);
nor U14043 (N_14043,N_13822,N_13914);
xnor U14044 (N_14044,N_13812,N_13805);
and U14045 (N_14045,N_13893,N_13922);
nor U14046 (N_14046,N_13875,N_13829);
xnor U14047 (N_14047,N_13800,N_13824);
nand U14048 (N_14048,N_13861,N_13895);
xnor U14049 (N_14049,N_13909,N_13836);
xor U14050 (N_14050,N_13809,N_13935);
nor U14051 (N_14051,N_13862,N_13805);
nor U14052 (N_14052,N_13860,N_13820);
nor U14053 (N_14053,N_13934,N_13896);
nand U14054 (N_14054,N_13844,N_13861);
nor U14055 (N_14055,N_13800,N_13832);
xnor U14056 (N_14056,N_13840,N_13835);
and U14057 (N_14057,N_13841,N_13881);
nor U14058 (N_14058,N_13914,N_13811);
and U14059 (N_14059,N_13862,N_13881);
nand U14060 (N_14060,N_13842,N_13850);
and U14061 (N_14061,N_13844,N_13916);
nor U14062 (N_14062,N_13806,N_13829);
or U14063 (N_14063,N_13846,N_13895);
xnor U14064 (N_14064,N_13814,N_13883);
xnor U14065 (N_14065,N_13935,N_13905);
or U14066 (N_14066,N_13814,N_13878);
xor U14067 (N_14067,N_13803,N_13907);
nand U14068 (N_14068,N_13844,N_13948);
nand U14069 (N_14069,N_13873,N_13900);
xor U14070 (N_14070,N_13840,N_13868);
and U14071 (N_14071,N_13872,N_13843);
xnor U14072 (N_14072,N_13846,N_13822);
nor U14073 (N_14073,N_13813,N_13886);
or U14074 (N_14074,N_13858,N_13921);
nand U14075 (N_14075,N_13902,N_13949);
nor U14076 (N_14076,N_13820,N_13891);
and U14077 (N_14077,N_13863,N_13881);
nand U14078 (N_14078,N_13858,N_13869);
and U14079 (N_14079,N_13903,N_13947);
or U14080 (N_14080,N_13813,N_13854);
nor U14081 (N_14081,N_13885,N_13897);
or U14082 (N_14082,N_13939,N_13866);
nand U14083 (N_14083,N_13851,N_13865);
and U14084 (N_14084,N_13878,N_13857);
and U14085 (N_14085,N_13933,N_13827);
or U14086 (N_14086,N_13941,N_13915);
and U14087 (N_14087,N_13819,N_13889);
xnor U14088 (N_14088,N_13881,N_13805);
or U14089 (N_14089,N_13936,N_13919);
or U14090 (N_14090,N_13886,N_13921);
nor U14091 (N_14091,N_13808,N_13911);
nand U14092 (N_14092,N_13889,N_13841);
nor U14093 (N_14093,N_13915,N_13920);
and U14094 (N_14094,N_13844,N_13805);
xor U14095 (N_14095,N_13875,N_13889);
nand U14096 (N_14096,N_13918,N_13926);
and U14097 (N_14097,N_13926,N_13858);
and U14098 (N_14098,N_13901,N_13907);
or U14099 (N_14099,N_13807,N_13860);
nand U14100 (N_14100,N_13996,N_14008);
nor U14101 (N_14101,N_13989,N_13969);
nand U14102 (N_14102,N_14087,N_14015);
xor U14103 (N_14103,N_14082,N_13990);
xor U14104 (N_14104,N_13953,N_13986);
and U14105 (N_14105,N_14033,N_13963);
xor U14106 (N_14106,N_13978,N_14064);
nor U14107 (N_14107,N_14060,N_13954);
or U14108 (N_14108,N_14084,N_14017);
nor U14109 (N_14109,N_13955,N_14030);
nor U14110 (N_14110,N_14001,N_14031);
xnor U14111 (N_14111,N_14038,N_14075);
xor U14112 (N_14112,N_13961,N_13972);
and U14113 (N_14113,N_13951,N_14007);
nand U14114 (N_14114,N_14083,N_13980);
and U14115 (N_14115,N_14035,N_13962);
or U14116 (N_14116,N_14046,N_14022);
or U14117 (N_14117,N_14023,N_13999);
and U14118 (N_14118,N_13958,N_13992);
nor U14119 (N_14119,N_14039,N_14071);
and U14120 (N_14120,N_13984,N_14045);
xnor U14121 (N_14121,N_13987,N_13993);
and U14122 (N_14122,N_14029,N_14014);
nand U14123 (N_14123,N_14053,N_14074);
and U14124 (N_14124,N_14054,N_14069);
and U14125 (N_14125,N_14055,N_13957);
and U14126 (N_14126,N_14066,N_14009);
nand U14127 (N_14127,N_14044,N_13979);
and U14128 (N_14128,N_14052,N_14000);
nor U14129 (N_14129,N_14036,N_13994);
nand U14130 (N_14130,N_13968,N_14051);
xnor U14131 (N_14131,N_14097,N_13976);
and U14132 (N_14132,N_13995,N_14024);
or U14133 (N_14133,N_14050,N_13985);
nand U14134 (N_14134,N_14080,N_14081);
or U14135 (N_14135,N_14077,N_14013);
nand U14136 (N_14136,N_14093,N_14010);
and U14137 (N_14137,N_14088,N_14095);
nor U14138 (N_14138,N_14025,N_14004);
xor U14139 (N_14139,N_13998,N_14034);
nor U14140 (N_14140,N_14098,N_14057);
or U14141 (N_14141,N_14076,N_14027);
and U14142 (N_14142,N_14012,N_14028);
nand U14143 (N_14143,N_13950,N_13973);
xnor U14144 (N_14144,N_14002,N_14059);
nor U14145 (N_14145,N_14099,N_14070);
nand U14146 (N_14146,N_14041,N_14063);
nor U14147 (N_14147,N_13991,N_14062);
or U14148 (N_14148,N_14092,N_14037);
nor U14149 (N_14149,N_14061,N_13971);
nor U14150 (N_14150,N_14072,N_14090);
xnor U14151 (N_14151,N_14040,N_14067);
xnor U14152 (N_14152,N_14011,N_13974);
nand U14153 (N_14153,N_14006,N_13967);
nand U14154 (N_14154,N_14094,N_14096);
xor U14155 (N_14155,N_13956,N_14068);
or U14156 (N_14156,N_14005,N_13959);
xnor U14157 (N_14157,N_13982,N_14058);
or U14158 (N_14158,N_14020,N_13997);
nand U14159 (N_14159,N_14042,N_14003);
and U14160 (N_14160,N_14091,N_14078);
or U14161 (N_14161,N_14085,N_14079);
nor U14162 (N_14162,N_14089,N_13983);
nand U14163 (N_14163,N_13960,N_14018);
xnor U14164 (N_14164,N_13966,N_14021);
nand U14165 (N_14165,N_14056,N_13975);
nand U14166 (N_14166,N_14049,N_13964);
and U14167 (N_14167,N_13970,N_14048);
xnor U14168 (N_14168,N_14019,N_14047);
nor U14169 (N_14169,N_13981,N_14026);
nor U14170 (N_14170,N_14016,N_14086);
or U14171 (N_14171,N_13952,N_14065);
and U14172 (N_14172,N_13988,N_14043);
nor U14173 (N_14173,N_13965,N_14032);
nor U14174 (N_14174,N_14073,N_13977);
nand U14175 (N_14175,N_14076,N_14004);
nand U14176 (N_14176,N_14033,N_13962);
and U14177 (N_14177,N_14002,N_13956);
xor U14178 (N_14178,N_14099,N_14055);
xor U14179 (N_14179,N_14021,N_14095);
xor U14180 (N_14180,N_14040,N_14021);
nand U14181 (N_14181,N_14025,N_13951);
nor U14182 (N_14182,N_14044,N_14013);
xnor U14183 (N_14183,N_13954,N_14004);
xnor U14184 (N_14184,N_14047,N_13950);
xor U14185 (N_14185,N_14093,N_14015);
or U14186 (N_14186,N_13959,N_14073);
or U14187 (N_14187,N_13976,N_14055);
nand U14188 (N_14188,N_13960,N_14073);
nand U14189 (N_14189,N_14047,N_13998);
or U14190 (N_14190,N_13990,N_13995);
xor U14191 (N_14191,N_13952,N_14020);
nand U14192 (N_14192,N_14065,N_14094);
or U14193 (N_14193,N_14033,N_13960);
and U14194 (N_14194,N_14087,N_14004);
and U14195 (N_14195,N_14031,N_13981);
or U14196 (N_14196,N_14017,N_14029);
and U14197 (N_14197,N_13969,N_14035);
and U14198 (N_14198,N_14016,N_14010);
xor U14199 (N_14199,N_14076,N_13984);
and U14200 (N_14200,N_14091,N_14047);
or U14201 (N_14201,N_14068,N_13957);
xnor U14202 (N_14202,N_14006,N_14062);
xnor U14203 (N_14203,N_14012,N_14039);
nand U14204 (N_14204,N_13966,N_14009);
and U14205 (N_14205,N_14029,N_13979);
nor U14206 (N_14206,N_14036,N_13971);
nand U14207 (N_14207,N_14070,N_14031);
nand U14208 (N_14208,N_14037,N_14013);
xor U14209 (N_14209,N_13960,N_14030);
or U14210 (N_14210,N_14006,N_14067);
and U14211 (N_14211,N_14066,N_13950);
xnor U14212 (N_14212,N_14018,N_14042);
nor U14213 (N_14213,N_13966,N_14072);
or U14214 (N_14214,N_14082,N_13996);
or U14215 (N_14215,N_14013,N_13977);
and U14216 (N_14216,N_14078,N_13952);
nor U14217 (N_14217,N_14017,N_14099);
nand U14218 (N_14218,N_14043,N_14022);
xor U14219 (N_14219,N_14006,N_14055);
or U14220 (N_14220,N_13976,N_14077);
nand U14221 (N_14221,N_14080,N_14094);
nand U14222 (N_14222,N_14033,N_14029);
xor U14223 (N_14223,N_14079,N_14081);
or U14224 (N_14224,N_13986,N_14091);
nor U14225 (N_14225,N_14004,N_14045);
and U14226 (N_14226,N_13959,N_13986);
or U14227 (N_14227,N_14090,N_13958);
or U14228 (N_14228,N_13982,N_14085);
nand U14229 (N_14229,N_14013,N_14008);
nand U14230 (N_14230,N_14034,N_13979);
nor U14231 (N_14231,N_13994,N_14032);
nand U14232 (N_14232,N_13994,N_14044);
nand U14233 (N_14233,N_14022,N_14020);
nand U14234 (N_14234,N_14009,N_14068);
or U14235 (N_14235,N_13955,N_14029);
xor U14236 (N_14236,N_14060,N_13993);
xnor U14237 (N_14237,N_14036,N_13982);
or U14238 (N_14238,N_14016,N_14064);
nand U14239 (N_14239,N_13974,N_14093);
or U14240 (N_14240,N_13975,N_14044);
and U14241 (N_14241,N_13995,N_14076);
or U14242 (N_14242,N_13965,N_14065);
nor U14243 (N_14243,N_13988,N_14034);
or U14244 (N_14244,N_13992,N_14044);
or U14245 (N_14245,N_13993,N_14048);
and U14246 (N_14246,N_13989,N_14029);
or U14247 (N_14247,N_14095,N_13999);
nand U14248 (N_14248,N_14076,N_14099);
and U14249 (N_14249,N_13954,N_14025);
xor U14250 (N_14250,N_14173,N_14131);
xor U14251 (N_14251,N_14214,N_14125);
xor U14252 (N_14252,N_14197,N_14176);
or U14253 (N_14253,N_14102,N_14191);
and U14254 (N_14254,N_14215,N_14226);
nor U14255 (N_14255,N_14117,N_14127);
and U14256 (N_14256,N_14244,N_14223);
or U14257 (N_14257,N_14248,N_14157);
nand U14258 (N_14258,N_14113,N_14154);
or U14259 (N_14259,N_14241,N_14130);
and U14260 (N_14260,N_14200,N_14218);
or U14261 (N_14261,N_14167,N_14229);
and U14262 (N_14262,N_14118,N_14109);
nand U14263 (N_14263,N_14186,N_14216);
and U14264 (N_14264,N_14202,N_14165);
xor U14265 (N_14265,N_14128,N_14141);
xnor U14266 (N_14266,N_14164,N_14124);
nor U14267 (N_14267,N_14210,N_14213);
xor U14268 (N_14268,N_14103,N_14160);
nand U14269 (N_14269,N_14150,N_14230);
nand U14270 (N_14270,N_14143,N_14169);
xor U14271 (N_14271,N_14132,N_14238);
and U14272 (N_14272,N_14152,N_14201);
and U14273 (N_14273,N_14158,N_14148);
or U14274 (N_14274,N_14174,N_14136);
and U14275 (N_14275,N_14145,N_14196);
and U14276 (N_14276,N_14206,N_14178);
nor U14277 (N_14277,N_14114,N_14190);
or U14278 (N_14278,N_14179,N_14239);
and U14279 (N_14279,N_14107,N_14151);
or U14280 (N_14280,N_14208,N_14108);
and U14281 (N_14281,N_14188,N_14175);
xor U14282 (N_14282,N_14121,N_14246);
and U14283 (N_14283,N_14123,N_14115);
and U14284 (N_14284,N_14224,N_14162);
and U14285 (N_14285,N_14122,N_14180);
xor U14286 (N_14286,N_14189,N_14227);
or U14287 (N_14287,N_14234,N_14116);
and U14288 (N_14288,N_14168,N_14100);
and U14289 (N_14289,N_14187,N_14101);
nand U14290 (N_14290,N_14219,N_14155);
nand U14291 (N_14291,N_14156,N_14171);
and U14292 (N_14292,N_14110,N_14153);
xnor U14293 (N_14293,N_14177,N_14137);
and U14294 (N_14294,N_14233,N_14149);
nand U14295 (N_14295,N_14147,N_14209);
and U14296 (N_14296,N_14184,N_14182);
nand U14297 (N_14297,N_14163,N_14138);
xor U14298 (N_14298,N_14139,N_14211);
xnor U14299 (N_14299,N_14221,N_14237);
xnor U14300 (N_14300,N_14106,N_14183);
nand U14301 (N_14301,N_14135,N_14105);
and U14302 (N_14302,N_14161,N_14193);
or U14303 (N_14303,N_14172,N_14192);
and U14304 (N_14304,N_14129,N_14243);
nand U14305 (N_14305,N_14236,N_14111);
nor U14306 (N_14306,N_14235,N_14198);
or U14307 (N_14307,N_14199,N_14170);
nand U14308 (N_14308,N_14205,N_14232);
and U14309 (N_14309,N_14247,N_14207);
and U14310 (N_14310,N_14245,N_14144);
or U14311 (N_14311,N_14134,N_14194);
and U14312 (N_14312,N_14140,N_14146);
nor U14313 (N_14313,N_14126,N_14231);
or U14314 (N_14314,N_14222,N_14212);
and U14315 (N_14315,N_14225,N_14217);
nand U14316 (N_14316,N_14142,N_14185);
nand U14317 (N_14317,N_14240,N_14104);
or U14318 (N_14318,N_14228,N_14204);
nand U14319 (N_14319,N_14195,N_14133);
nor U14320 (N_14320,N_14203,N_14119);
or U14321 (N_14321,N_14181,N_14249);
nor U14322 (N_14322,N_14120,N_14112);
nand U14323 (N_14323,N_14220,N_14159);
or U14324 (N_14324,N_14166,N_14242);
and U14325 (N_14325,N_14127,N_14228);
nand U14326 (N_14326,N_14197,N_14219);
nor U14327 (N_14327,N_14216,N_14115);
xnor U14328 (N_14328,N_14148,N_14216);
nand U14329 (N_14329,N_14127,N_14186);
xor U14330 (N_14330,N_14111,N_14138);
and U14331 (N_14331,N_14148,N_14115);
nor U14332 (N_14332,N_14186,N_14243);
and U14333 (N_14333,N_14154,N_14146);
xor U14334 (N_14334,N_14235,N_14109);
xor U14335 (N_14335,N_14241,N_14182);
and U14336 (N_14336,N_14234,N_14177);
or U14337 (N_14337,N_14118,N_14225);
and U14338 (N_14338,N_14171,N_14135);
and U14339 (N_14339,N_14142,N_14191);
and U14340 (N_14340,N_14117,N_14141);
or U14341 (N_14341,N_14176,N_14149);
nor U14342 (N_14342,N_14201,N_14232);
xnor U14343 (N_14343,N_14239,N_14236);
and U14344 (N_14344,N_14117,N_14147);
and U14345 (N_14345,N_14200,N_14220);
nand U14346 (N_14346,N_14113,N_14244);
xnor U14347 (N_14347,N_14130,N_14140);
nor U14348 (N_14348,N_14230,N_14168);
and U14349 (N_14349,N_14241,N_14229);
nor U14350 (N_14350,N_14208,N_14118);
nor U14351 (N_14351,N_14158,N_14121);
nor U14352 (N_14352,N_14167,N_14183);
xor U14353 (N_14353,N_14144,N_14240);
nor U14354 (N_14354,N_14237,N_14241);
xnor U14355 (N_14355,N_14177,N_14249);
xnor U14356 (N_14356,N_14112,N_14211);
xor U14357 (N_14357,N_14162,N_14115);
and U14358 (N_14358,N_14232,N_14121);
and U14359 (N_14359,N_14136,N_14124);
nand U14360 (N_14360,N_14108,N_14102);
or U14361 (N_14361,N_14162,N_14205);
or U14362 (N_14362,N_14241,N_14216);
nand U14363 (N_14363,N_14177,N_14166);
or U14364 (N_14364,N_14244,N_14146);
xor U14365 (N_14365,N_14159,N_14113);
or U14366 (N_14366,N_14142,N_14184);
xor U14367 (N_14367,N_14115,N_14204);
and U14368 (N_14368,N_14185,N_14206);
nand U14369 (N_14369,N_14164,N_14191);
nand U14370 (N_14370,N_14238,N_14204);
nor U14371 (N_14371,N_14141,N_14144);
xor U14372 (N_14372,N_14180,N_14126);
nor U14373 (N_14373,N_14111,N_14224);
or U14374 (N_14374,N_14247,N_14119);
nand U14375 (N_14375,N_14157,N_14101);
xor U14376 (N_14376,N_14221,N_14231);
xor U14377 (N_14377,N_14182,N_14138);
xor U14378 (N_14378,N_14129,N_14101);
xnor U14379 (N_14379,N_14173,N_14171);
and U14380 (N_14380,N_14141,N_14230);
nand U14381 (N_14381,N_14101,N_14238);
nand U14382 (N_14382,N_14214,N_14167);
and U14383 (N_14383,N_14248,N_14185);
nor U14384 (N_14384,N_14129,N_14233);
xnor U14385 (N_14385,N_14212,N_14129);
nor U14386 (N_14386,N_14100,N_14180);
nand U14387 (N_14387,N_14139,N_14172);
and U14388 (N_14388,N_14140,N_14216);
and U14389 (N_14389,N_14193,N_14237);
nor U14390 (N_14390,N_14213,N_14115);
or U14391 (N_14391,N_14175,N_14185);
xor U14392 (N_14392,N_14245,N_14128);
nand U14393 (N_14393,N_14219,N_14173);
and U14394 (N_14394,N_14123,N_14131);
xnor U14395 (N_14395,N_14149,N_14177);
nor U14396 (N_14396,N_14165,N_14153);
or U14397 (N_14397,N_14218,N_14117);
or U14398 (N_14398,N_14150,N_14124);
nand U14399 (N_14399,N_14227,N_14197);
nor U14400 (N_14400,N_14252,N_14333);
xnor U14401 (N_14401,N_14298,N_14352);
and U14402 (N_14402,N_14341,N_14317);
and U14403 (N_14403,N_14285,N_14251);
xor U14404 (N_14404,N_14379,N_14388);
xor U14405 (N_14405,N_14353,N_14377);
xor U14406 (N_14406,N_14382,N_14258);
xnor U14407 (N_14407,N_14334,N_14306);
nand U14408 (N_14408,N_14271,N_14354);
or U14409 (N_14409,N_14351,N_14350);
or U14410 (N_14410,N_14301,N_14320);
nor U14411 (N_14411,N_14344,N_14338);
xnor U14412 (N_14412,N_14256,N_14308);
xnor U14413 (N_14413,N_14323,N_14290);
xnor U14414 (N_14414,N_14305,N_14291);
xnor U14415 (N_14415,N_14313,N_14391);
xor U14416 (N_14416,N_14259,N_14385);
xnor U14417 (N_14417,N_14349,N_14342);
nand U14418 (N_14418,N_14277,N_14287);
nor U14419 (N_14419,N_14274,N_14363);
or U14420 (N_14420,N_14369,N_14278);
nor U14421 (N_14421,N_14378,N_14288);
xor U14422 (N_14422,N_14335,N_14370);
nor U14423 (N_14423,N_14264,N_14266);
or U14424 (N_14424,N_14304,N_14282);
xor U14425 (N_14425,N_14325,N_14322);
and U14426 (N_14426,N_14381,N_14366);
nand U14427 (N_14427,N_14260,N_14374);
xnor U14428 (N_14428,N_14254,N_14348);
and U14429 (N_14429,N_14280,N_14272);
nor U14430 (N_14430,N_14293,N_14359);
or U14431 (N_14431,N_14292,N_14289);
nand U14432 (N_14432,N_14358,N_14332);
nor U14433 (N_14433,N_14294,N_14387);
nand U14434 (N_14434,N_14315,N_14362);
nor U14435 (N_14435,N_14283,N_14257);
nand U14436 (N_14436,N_14331,N_14371);
and U14437 (N_14437,N_14311,N_14393);
and U14438 (N_14438,N_14376,N_14398);
or U14439 (N_14439,N_14330,N_14345);
and U14440 (N_14440,N_14383,N_14261);
nand U14441 (N_14441,N_14312,N_14270);
nand U14442 (N_14442,N_14268,N_14314);
nor U14443 (N_14443,N_14250,N_14343);
or U14444 (N_14444,N_14284,N_14321);
nand U14445 (N_14445,N_14375,N_14367);
nand U14446 (N_14446,N_14279,N_14364);
and U14447 (N_14447,N_14255,N_14372);
nand U14448 (N_14448,N_14267,N_14384);
nor U14449 (N_14449,N_14273,N_14275);
nand U14450 (N_14450,N_14397,N_14392);
xor U14451 (N_14451,N_14365,N_14319);
nor U14452 (N_14452,N_14355,N_14390);
nand U14453 (N_14453,N_14328,N_14380);
nor U14454 (N_14454,N_14327,N_14269);
and U14455 (N_14455,N_14329,N_14368);
nor U14456 (N_14456,N_14297,N_14340);
nand U14457 (N_14457,N_14395,N_14263);
nor U14458 (N_14458,N_14326,N_14324);
nand U14459 (N_14459,N_14394,N_14346);
and U14460 (N_14460,N_14310,N_14337);
or U14461 (N_14461,N_14361,N_14253);
xor U14462 (N_14462,N_14399,N_14347);
or U14463 (N_14463,N_14396,N_14302);
xor U14464 (N_14464,N_14295,N_14336);
nand U14465 (N_14465,N_14373,N_14360);
nor U14466 (N_14466,N_14309,N_14318);
and U14467 (N_14467,N_14300,N_14316);
nor U14468 (N_14468,N_14296,N_14276);
xor U14469 (N_14469,N_14339,N_14356);
or U14470 (N_14470,N_14357,N_14386);
and U14471 (N_14471,N_14307,N_14265);
xor U14472 (N_14472,N_14286,N_14389);
nand U14473 (N_14473,N_14281,N_14262);
or U14474 (N_14474,N_14299,N_14303);
xnor U14475 (N_14475,N_14265,N_14368);
nor U14476 (N_14476,N_14353,N_14260);
and U14477 (N_14477,N_14316,N_14339);
and U14478 (N_14478,N_14280,N_14390);
or U14479 (N_14479,N_14270,N_14308);
nand U14480 (N_14480,N_14267,N_14273);
nor U14481 (N_14481,N_14299,N_14338);
nor U14482 (N_14482,N_14267,N_14258);
nor U14483 (N_14483,N_14291,N_14370);
xnor U14484 (N_14484,N_14323,N_14381);
xnor U14485 (N_14485,N_14386,N_14355);
and U14486 (N_14486,N_14380,N_14379);
or U14487 (N_14487,N_14363,N_14280);
nor U14488 (N_14488,N_14250,N_14252);
and U14489 (N_14489,N_14275,N_14276);
nor U14490 (N_14490,N_14375,N_14374);
nand U14491 (N_14491,N_14328,N_14383);
nand U14492 (N_14492,N_14393,N_14383);
or U14493 (N_14493,N_14394,N_14362);
nand U14494 (N_14494,N_14375,N_14351);
nand U14495 (N_14495,N_14271,N_14266);
nand U14496 (N_14496,N_14252,N_14323);
or U14497 (N_14497,N_14304,N_14343);
nor U14498 (N_14498,N_14371,N_14308);
and U14499 (N_14499,N_14355,N_14325);
and U14500 (N_14500,N_14327,N_14367);
xor U14501 (N_14501,N_14278,N_14284);
nor U14502 (N_14502,N_14380,N_14359);
and U14503 (N_14503,N_14339,N_14326);
nand U14504 (N_14504,N_14309,N_14276);
nor U14505 (N_14505,N_14381,N_14370);
xnor U14506 (N_14506,N_14269,N_14255);
nor U14507 (N_14507,N_14254,N_14335);
nor U14508 (N_14508,N_14344,N_14346);
xnor U14509 (N_14509,N_14293,N_14372);
nor U14510 (N_14510,N_14322,N_14397);
nor U14511 (N_14511,N_14363,N_14336);
and U14512 (N_14512,N_14255,N_14277);
xnor U14513 (N_14513,N_14258,N_14385);
or U14514 (N_14514,N_14340,N_14319);
nand U14515 (N_14515,N_14374,N_14360);
nor U14516 (N_14516,N_14394,N_14325);
nor U14517 (N_14517,N_14304,N_14367);
nand U14518 (N_14518,N_14376,N_14300);
xor U14519 (N_14519,N_14353,N_14374);
or U14520 (N_14520,N_14370,N_14351);
and U14521 (N_14521,N_14399,N_14285);
or U14522 (N_14522,N_14325,N_14278);
nand U14523 (N_14523,N_14336,N_14344);
nand U14524 (N_14524,N_14339,N_14283);
nor U14525 (N_14525,N_14375,N_14285);
and U14526 (N_14526,N_14341,N_14302);
nor U14527 (N_14527,N_14261,N_14260);
nor U14528 (N_14528,N_14345,N_14323);
nor U14529 (N_14529,N_14343,N_14382);
or U14530 (N_14530,N_14380,N_14257);
nand U14531 (N_14531,N_14276,N_14331);
nand U14532 (N_14532,N_14379,N_14340);
nor U14533 (N_14533,N_14313,N_14374);
or U14534 (N_14534,N_14262,N_14265);
or U14535 (N_14535,N_14285,N_14397);
xor U14536 (N_14536,N_14312,N_14367);
xnor U14537 (N_14537,N_14340,N_14378);
nand U14538 (N_14538,N_14272,N_14343);
nand U14539 (N_14539,N_14347,N_14344);
and U14540 (N_14540,N_14372,N_14354);
nand U14541 (N_14541,N_14310,N_14324);
xnor U14542 (N_14542,N_14273,N_14268);
nand U14543 (N_14543,N_14288,N_14254);
and U14544 (N_14544,N_14393,N_14250);
and U14545 (N_14545,N_14298,N_14345);
or U14546 (N_14546,N_14352,N_14378);
and U14547 (N_14547,N_14353,N_14271);
and U14548 (N_14548,N_14299,N_14385);
or U14549 (N_14549,N_14381,N_14384);
and U14550 (N_14550,N_14440,N_14404);
nand U14551 (N_14551,N_14519,N_14539);
xor U14552 (N_14552,N_14537,N_14460);
or U14553 (N_14553,N_14464,N_14479);
xor U14554 (N_14554,N_14503,N_14472);
or U14555 (N_14555,N_14480,N_14490);
xnor U14556 (N_14556,N_14531,N_14439);
nand U14557 (N_14557,N_14488,N_14409);
and U14558 (N_14558,N_14415,N_14524);
nor U14559 (N_14559,N_14508,N_14514);
xor U14560 (N_14560,N_14493,N_14471);
nand U14561 (N_14561,N_14529,N_14433);
nor U14562 (N_14562,N_14417,N_14408);
and U14563 (N_14563,N_14434,N_14419);
nor U14564 (N_14564,N_14509,N_14455);
and U14565 (N_14565,N_14459,N_14421);
and U14566 (N_14566,N_14427,N_14468);
nand U14567 (N_14567,N_14424,N_14450);
xor U14568 (N_14568,N_14518,N_14446);
xnor U14569 (N_14569,N_14517,N_14527);
and U14570 (N_14570,N_14512,N_14429);
or U14571 (N_14571,N_14501,N_14444);
or U14572 (N_14572,N_14413,N_14476);
nor U14573 (N_14573,N_14478,N_14422);
and U14574 (N_14574,N_14420,N_14474);
and U14575 (N_14575,N_14410,N_14462);
or U14576 (N_14576,N_14411,N_14454);
and U14577 (N_14577,N_14428,N_14482);
xor U14578 (N_14578,N_14521,N_14532);
nor U14579 (N_14579,N_14447,N_14442);
and U14580 (N_14580,N_14516,N_14485);
or U14581 (N_14581,N_14489,N_14401);
and U14582 (N_14582,N_14522,N_14547);
and U14583 (N_14583,N_14545,N_14469);
xor U14584 (N_14584,N_14473,N_14412);
and U14585 (N_14585,N_14430,N_14494);
xor U14586 (N_14586,N_14465,N_14491);
xnor U14587 (N_14587,N_14477,N_14435);
nand U14588 (N_14588,N_14484,N_14492);
nor U14589 (N_14589,N_14483,N_14470);
xnor U14590 (N_14590,N_14498,N_14418);
nor U14591 (N_14591,N_14438,N_14538);
nand U14592 (N_14592,N_14487,N_14443);
nor U14593 (N_14593,N_14497,N_14405);
or U14594 (N_14594,N_14511,N_14437);
nor U14595 (N_14595,N_14549,N_14402);
nand U14596 (N_14596,N_14431,N_14542);
xnor U14597 (N_14597,N_14504,N_14499);
nor U14598 (N_14598,N_14451,N_14535);
nor U14599 (N_14599,N_14526,N_14533);
nor U14600 (N_14600,N_14448,N_14528);
nand U14601 (N_14601,N_14403,N_14505);
xor U14602 (N_14602,N_14452,N_14453);
xnor U14603 (N_14603,N_14449,N_14400);
or U14604 (N_14604,N_14432,N_14543);
and U14605 (N_14605,N_14507,N_14520);
xnor U14606 (N_14606,N_14544,N_14481);
and U14607 (N_14607,N_14496,N_14534);
xor U14608 (N_14608,N_14467,N_14458);
or U14609 (N_14609,N_14416,N_14515);
xor U14610 (N_14610,N_14461,N_14546);
nor U14611 (N_14611,N_14475,N_14414);
xnor U14612 (N_14612,N_14495,N_14513);
or U14613 (N_14613,N_14407,N_14425);
xnor U14614 (N_14614,N_14506,N_14530);
nand U14615 (N_14615,N_14536,N_14445);
or U14616 (N_14616,N_14502,N_14406);
xor U14617 (N_14617,N_14500,N_14457);
or U14618 (N_14618,N_14510,N_14486);
xor U14619 (N_14619,N_14423,N_14466);
nand U14620 (N_14620,N_14441,N_14548);
xnor U14621 (N_14621,N_14426,N_14523);
xnor U14622 (N_14622,N_14540,N_14463);
nand U14623 (N_14623,N_14436,N_14525);
xnor U14624 (N_14624,N_14541,N_14456);
nor U14625 (N_14625,N_14420,N_14400);
xor U14626 (N_14626,N_14425,N_14478);
xor U14627 (N_14627,N_14476,N_14472);
nor U14628 (N_14628,N_14456,N_14411);
nand U14629 (N_14629,N_14438,N_14439);
and U14630 (N_14630,N_14460,N_14511);
and U14631 (N_14631,N_14403,N_14544);
nand U14632 (N_14632,N_14539,N_14544);
nor U14633 (N_14633,N_14479,N_14538);
xor U14634 (N_14634,N_14463,N_14432);
or U14635 (N_14635,N_14401,N_14472);
or U14636 (N_14636,N_14498,N_14507);
nor U14637 (N_14637,N_14530,N_14430);
nor U14638 (N_14638,N_14429,N_14432);
or U14639 (N_14639,N_14413,N_14475);
xnor U14640 (N_14640,N_14506,N_14516);
xnor U14641 (N_14641,N_14497,N_14450);
xor U14642 (N_14642,N_14471,N_14492);
nand U14643 (N_14643,N_14546,N_14400);
nand U14644 (N_14644,N_14443,N_14426);
xor U14645 (N_14645,N_14485,N_14511);
nor U14646 (N_14646,N_14483,N_14486);
xor U14647 (N_14647,N_14428,N_14404);
and U14648 (N_14648,N_14495,N_14407);
and U14649 (N_14649,N_14464,N_14523);
nor U14650 (N_14650,N_14508,N_14421);
nor U14651 (N_14651,N_14510,N_14445);
nand U14652 (N_14652,N_14417,N_14491);
and U14653 (N_14653,N_14515,N_14402);
nor U14654 (N_14654,N_14475,N_14539);
nand U14655 (N_14655,N_14436,N_14457);
nor U14656 (N_14656,N_14416,N_14477);
nand U14657 (N_14657,N_14473,N_14487);
and U14658 (N_14658,N_14462,N_14471);
nand U14659 (N_14659,N_14410,N_14477);
or U14660 (N_14660,N_14420,N_14491);
xnor U14661 (N_14661,N_14523,N_14511);
or U14662 (N_14662,N_14447,N_14444);
nand U14663 (N_14663,N_14407,N_14504);
xnor U14664 (N_14664,N_14444,N_14548);
or U14665 (N_14665,N_14546,N_14425);
nand U14666 (N_14666,N_14503,N_14493);
or U14667 (N_14667,N_14467,N_14514);
or U14668 (N_14668,N_14464,N_14445);
nor U14669 (N_14669,N_14515,N_14437);
and U14670 (N_14670,N_14405,N_14447);
xor U14671 (N_14671,N_14526,N_14534);
xor U14672 (N_14672,N_14538,N_14543);
and U14673 (N_14673,N_14446,N_14459);
or U14674 (N_14674,N_14446,N_14501);
and U14675 (N_14675,N_14479,N_14546);
and U14676 (N_14676,N_14536,N_14502);
and U14677 (N_14677,N_14504,N_14464);
nand U14678 (N_14678,N_14451,N_14508);
or U14679 (N_14679,N_14518,N_14481);
nand U14680 (N_14680,N_14528,N_14510);
xnor U14681 (N_14681,N_14527,N_14528);
nand U14682 (N_14682,N_14474,N_14411);
xor U14683 (N_14683,N_14411,N_14419);
nor U14684 (N_14684,N_14454,N_14407);
nand U14685 (N_14685,N_14537,N_14420);
nor U14686 (N_14686,N_14429,N_14476);
nor U14687 (N_14687,N_14506,N_14532);
or U14688 (N_14688,N_14474,N_14530);
xnor U14689 (N_14689,N_14543,N_14524);
nor U14690 (N_14690,N_14483,N_14475);
nand U14691 (N_14691,N_14438,N_14504);
and U14692 (N_14692,N_14526,N_14407);
and U14693 (N_14693,N_14442,N_14460);
and U14694 (N_14694,N_14522,N_14520);
and U14695 (N_14695,N_14414,N_14490);
xnor U14696 (N_14696,N_14544,N_14534);
nand U14697 (N_14697,N_14423,N_14535);
or U14698 (N_14698,N_14458,N_14446);
nand U14699 (N_14699,N_14484,N_14531);
and U14700 (N_14700,N_14643,N_14654);
and U14701 (N_14701,N_14552,N_14644);
xnor U14702 (N_14702,N_14669,N_14672);
or U14703 (N_14703,N_14610,N_14587);
nand U14704 (N_14704,N_14699,N_14615);
or U14705 (N_14705,N_14650,N_14664);
xnor U14706 (N_14706,N_14601,N_14653);
and U14707 (N_14707,N_14624,N_14687);
nor U14708 (N_14708,N_14586,N_14594);
and U14709 (N_14709,N_14690,N_14611);
xnor U14710 (N_14710,N_14657,N_14591);
or U14711 (N_14711,N_14625,N_14645);
nand U14712 (N_14712,N_14613,N_14651);
xor U14713 (N_14713,N_14692,N_14550);
nand U14714 (N_14714,N_14562,N_14685);
and U14715 (N_14715,N_14696,N_14668);
xnor U14716 (N_14716,N_14596,N_14676);
nor U14717 (N_14717,N_14678,N_14607);
nand U14718 (N_14718,N_14635,N_14585);
or U14719 (N_14719,N_14560,N_14660);
nand U14720 (N_14720,N_14673,N_14695);
or U14721 (N_14721,N_14572,N_14627);
and U14722 (N_14722,N_14683,N_14632);
nand U14723 (N_14723,N_14659,N_14663);
and U14724 (N_14724,N_14666,N_14598);
and U14725 (N_14725,N_14574,N_14599);
nand U14726 (N_14726,N_14697,N_14569);
nand U14727 (N_14727,N_14583,N_14577);
and U14728 (N_14728,N_14636,N_14584);
xor U14729 (N_14729,N_14553,N_14667);
xor U14730 (N_14730,N_14633,N_14620);
and U14731 (N_14731,N_14680,N_14593);
nand U14732 (N_14732,N_14595,N_14618);
nor U14733 (N_14733,N_14580,N_14564);
nor U14734 (N_14734,N_14665,N_14622);
and U14735 (N_14735,N_14681,N_14619);
nand U14736 (N_14736,N_14565,N_14694);
nand U14737 (N_14737,N_14614,N_14642);
or U14738 (N_14738,N_14629,N_14612);
nand U14739 (N_14739,N_14626,N_14630);
xnor U14740 (N_14740,N_14686,N_14570);
xor U14741 (N_14741,N_14648,N_14617);
or U14742 (N_14742,N_14682,N_14639);
and U14743 (N_14743,N_14606,N_14631);
nand U14744 (N_14744,N_14556,N_14671);
nand U14745 (N_14745,N_14634,N_14641);
or U14746 (N_14746,N_14674,N_14578);
nor U14747 (N_14747,N_14559,N_14688);
nand U14748 (N_14748,N_14608,N_14691);
xnor U14749 (N_14749,N_14621,N_14603);
nand U14750 (N_14750,N_14600,N_14605);
or U14751 (N_14751,N_14662,N_14647);
and U14752 (N_14752,N_14604,N_14675);
xor U14753 (N_14753,N_14581,N_14551);
nand U14754 (N_14754,N_14649,N_14575);
xnor U14755 (N_14755,N_14652,N_14558);
nand U14756 (N_14756,N_14563,N_14589);
and U14757 (N_14757,N_14590,N_14661);
and U14758 (N_14758,N_14561,N_14670);
and U14759 (N_14759,N_14623,N_14592);
nor U14760 (N_14760,N_14698,N_14677);
and U14761 (N_14761,N_14588,N_14571);
and U14762 (N_14762,N_14656,N_14679);
nand U14763 (N_14763,N_14597,N_14655);
xor U14764 (N_14764,N_14637,N_14602);
nand U14765 (N_14765,N_14573,N_14567);
nand U14766 (N_14766,N_14566,N_14576);
and U14767 (N_14767,N_14646,N_14554);
xor U14768 (N_14768,N_14557,N_14616);
nor U14769 (N_14769,N_14555,N_14689);
xor U14770 (N_14770,N_14658,N_14628);
nor U14771 (N_14771,N_14582,N_14609);
or U14772 (N_14772,N_14579,N_14693);
and U14773 (N_14773,N_14638,N_14684);
and U14774 (N_14774,N_14640,N_14568);
nor U14775 (N_14775,N_14691,N_14605);
or U14776 (N_14776,N_14588,N_14553);
nand U14777 (N_14777,N_14618,N_14676);
nor U14778 (N_14778,N_14632,N_14658);
xnor U14779 (N_14779,N_14631,N_14600);
xor U14780 (N_14780,N_14628,N_14698);
nand U14781 (N_14781,N_14553,N_14609);
and U14782 (N_14782,N_14656,N_14646);
and U14783 (N_14783,N_14586,N_14592);
nor U14784 (N_14784,N_14644,N_14683);
or U14785 (N_14785,N_14600,N_14560);
nor U14786 (N_14786,N_14571,N_14641);
and U14787 (N_14787,N_14670,N_14690);
nor U14788 (N_14788,N_14681,N_14652);
xnor U14789 (N_14789,N_14606,N_14638);
xor U14790 (N_14790,N_14592,N_14626);
nand U14791 (N_14791,N_14616,N_14597);
nand U14792 (N_14792,N_14558,N_14551);
nor U14793 (N_14793,N_14564,N_14653);
nor U14794 (N_14794,N_14659,N_14679);
nor U14795 (N_14795,N_14554,N_14683);
nor U14796 (N_14796,N_14686,N_14566);
nand U14797 (N_14797,N_14652,N_14661);
and U14798 (N_14798,N_14590,N_14694);
nor U14799 (N_14799,N_14681,N_14561);
nand U14800 (N_14800,N_14584,N_14639);
xnor U14801 (N_14801,N_14672,N_14665);
nor U14802 (N_14802,N_14564,N_14628);
xor U14803 (N_14803,N_14646,N_14658);
or U14804 (N_14804,N_14615,N_14641);
xnor U14805 (N_14805,N_14682,N_14670);
nand U14806 (N_14806,N_14577,N_14638);
nand U14807 (N_14807,N_14693,N_14554);
and U14808 (N_14808,N_14555,N_14639);
nand U14809 (N_14809,N_14666,N_14683);
nand U14810 (N_14810,N_14641,N_14611);
and U14811 (N_14811,N_14607,N_14664);
nand U14812 (N_14812,N_14668,N_14618);
nand U14813 (N_14813,N_14588,N_14611);
xnor U14814 (N_14814,N_14563,N_14609);
nor U14815 (N_14815,N_14614,N_14654);
xnor U14816 (N_14816,N_14656,N_14613);
and U14817 (N_14817,N_14570,N_14690);
nor U14818 (N_14818,N_14636,N_14595);
xor U14819 (N_14819,N_14558,N_14682);
nor U14820 (N_14820,N_14692,N_14589);
or U14821 (N_14821,N_14552,N_14633);
nand U14822 (N_14822,N_14572,N_14662);
nor U14823 (N_14823,N_14677,N_14570);
xor U14824 (N_14824,N_14652,N_14559);
xnor U14825 (N_14825,N_14624,N_14681);
xnor U14826 (N_14826,N_14682,N_14587);
or U14827 (N_14827,N_14593,N_14555);
nand U14828 (N_14828,N_14618,N_14596);
xnor U14829 (N_14829,N_14574,N_14565);
nand U14830 (N_14830,N_14670,N_14562);
xnor U14831 (N_14831,N_14606,N_14636);
xor U14832 (N_14832,N_14689,N_14582);
or U14833 (N_14833,N_14570,N_14661);
nand U14834 (N_14834,N_14692,N_14556);
xnor U14835 (N_14835,N_14561,N_14687);
xor U14836 (N_14836,N_14614,N_14699);
nor U14837 (N_14837,N_14633,N_14611);
and U14838 (N_14838,N_14600,N_14585);
and U14839 (N_14839,N_14612,N_14552);
nand U14840 (N_14840,N_14689,N_14684);
xnor U14841 (N_14841,N_14687,N_14692);
xor U14842 (N_14842,N_14678,N_14605);
nor U14843 (N_14843,N_14566,N_14577);
and U14844 (N_14844,N_14647,N_14588);
or U14845 (N_14845,N_14550,N_14609);
nand U14846 (N_14846,N_14591,N_14666);
xnor U14847 (N_14847,N_14662,N_14597);
nor U14848 (N_14848,N_14653,N_14689);
nor U14849 (N_14849,N_14558,N_14552);
nor U14850 (N_14850,N_14766,N_14770);
xor U14851 (N_14851,N_14754,N_14779);
and U14852 (N_14852,N_14750,N_14821);
nand U14853 (N_14853,N_14709,N_14728);
nor U14854 (N_14854,N_14820,N_14847);
nor U14855 (N_14855,N_14702,N_14727);
nor U14856 (N_14856,N_14741,N_14735);
and U14857 (N_14857,N_14729,N_14825);
and U14858 (N_14858,N_14849,N_14848);
nand U14859 (N_14859,N_14767,N_14737);
and U14860 (N_14860,N_14831,N_14829);
nor U14861 (N_14861,N_14832,N_14715);
nand U14862 (N_14862,N_14809,N_14733);
nand U14863 (N_14863,N_14710,N_14794);
xnor U14864 (N_14864,N_14802,N_14726);
nand U14865 (N_14865,N_14789,N_14792);
or U14866 (N_14866,N_14839,N_14722);
or U14867 (N_14867,N_14705,N_14747);
nand U14868 (N_14868,N_14842,N_14841);
and U14869 (N_14869,N_14769,N_14778);
or U14870 (N_14870,N_14730,N_14757);
and U14871 (N_14871,N_14781,N_14814);
nor U14872 (N_14872,N_14725,N_14751);
xor U14873 (N_14873,N_14758,N_14817);
xnor U14874 (N_14874,N_14800,N_14837);
nand U14875 (N_14875,N_14761,N_14791);
and U14876 (N_14876,N_14771,N_14810);
nand U14877 (N_14877,N_14703,N_14806);
or U14878 (N_14878,N_14707,N_14813);
nand U14879 (N_14879,N_14811,N_14720);
xor U14880 (N_14880,N_14783,N_14777);
nor U14881 (N_14881,N_14721,N_14723);
and U14882 (N_14882,N_14700,N_14840);
or U14883 (N_14883,N_14819,N_14785);
nand U14884 (N_14884,N_14714,N_14807);
nand U14885 (N_14885,N_14768,N_14774);
and U14886 (N_14886,N_14843,N_14803);
xnor U14887 (N_14887,N_14764,N_14738);
xor U14888 (N_14888,N_14815,N_14846);
or U14889 (N_14889,N_14739,N_14748);
xor U14890 (N_14890,N_14816,N_14743);
and U14891 (N_14891,N_14716,N_14724);
or U14892 (N_14892,N_14706,N_14717);
nor U14893 (N_14893,N_14746,N_14701);
and U14894 (N_14894,N_14736,N_14719);
and U14895 (N_14895,N_14773,N_14732);
xor U14896 (N_14896,N_14772,N_14760);
xnor U14897 (N_14897,N_14765,N_14822);
and U14898 (N_14898,N_14718,N_14740);
and U14899 (N_14899,N_14755,N_14834);
xor U14900 (N_14900,N_14805,N_14708);
nand U14901 (N_14901,N_14845,N_14790);
nor U14902 (N_14902,N_14827,N_14833);
nor U14903 (N_14903,N_14780,N_14711);
nand U14904 (N_14904,N_14745,N_14753);
nor U14905 (N_14905,N_14749,N_14787);
nand U14906 (N_14906,N_14734,N_14712);
xor U14907 (N_14907,N_14844,N_14756);
or U14908 (N_14908,N_14788,N_14826);
and U14909 (N_14909,N_14784,N_14776);
nor U14910 (N_14910,N_14744,N_14828);
xnor U14911 (N_14911,N_14795,N_14824);
nor U14912 (N_14912,N_14797,N_14759);
or U14913 (N_14913,N_14838,N_14731);
xnor U14914 (N_14914,N_14823,N_14796);
and U14915 (N_14915,N_14786,N_14782);
xnor U14916 (N_14916,N_14830,N_14713);
or U14917 (N_14917,N_14799,N_14742);
or U14918 (N_14918,N_14835,N_14804);
or U14919 (N_14919,N_14836,N_14763);
and U14920 (N_14920,N_14752,N_14812);
nand U14921 (N_14921,N_14798,N_14704);
or U14922 (N_14922,N_14818,N_14801);
or U14923 (N_14923,N_14762,N_14793);
xnor U14924 (N_14924,N_14808,N_14775);
and U14925 (N_14925,N_14732,N_14799);
and U14926 (N_14926,N_14841,N_14770);
nor U14927 (N_14927,N_14803,N_14796);
nand U14928 (N_14928,N_14721,N_14739);
and U14929 (N_14929,N_14705,N_14722);
xnor U14930 (N_14930,N_14845,N_14779);
nand U14931 (N_14931,N_14729,N_14768);
nor U14932 (N_14932,N_14713,N_14764);
nand U14933 (N_14933,N_14804,N_14703);
nand U14934 (N_14934,N_14721,N_14843);
xor U14935 (N_14935,N_14823,N_14757);
or U14936 (N_14936,N_14755,N_14786);
nand U14937 (N_14937,N_14702,N_14712);
xor U14938 (N_14938,N_14702,N_14816);
nor U14939 (N_14939,N_14809,N_14760);
and U14940 (N_14940,N_14710,N_14813);
or U14941 (N_14941,N_14793,N_14764);
xnor U14942 (N_14942,N_14714,N_14709);
or U14943 (N_14943,N_14758,N_14712);
xnor U14944 (N_14944,N_14708,N_14806);
nor U14945 (N_14945,N_14736,N_14740);
xor U14946 (N_14946,N_14783,N_14818);
and U14947 (N_14947,N_14849,N_14708);
xor U14948 (N_14948,N_14805,N_14750);
nand U14949 (N_14949,N_14837,N_14839);
nor U14950 (N_14950,N_14839,N_14849);
and U14951 (N_14951,N_14770,N_14849);
and U14952 (N_14952,N_14804,N_14705);
nand U14953 (N_14953,N_14821,N_14797);
or U14954 (N_14954,N_14711,N_14837);
and U14955 (N_14955,N_14805,N_14827);
nand U14956 (N_14956,N_14783,N_14738);
or U14957 (N_14957,N_14798,N_14703);
and U14958 (N_14958,N_14727,N_14707);
nand U14959 (N_14959,N_14765,N_14725);
nor U14960 (N_14960,N_14708,N_14839);
and U14961 (N_14961,N_14776,N_14764);
nor U14962 (N_14962,N_14812,N_14789);
xnor U14963 (N_14963,N_14837,N_14784);
or U14964 (N_14964,N_14818,N_14750);
nor U14965 (N_14965,N_14742,N_14730);
and U14966 (N_14966,N_14763,N_14733);
xor U14967 (N_14967,N_14821,N_14743);
xnor U14968 (N_14968,N_14768,N_14818);
nand U14969 (N_14969,N_14820,N_14752);
or U14970 (N_14970,N_14729,N_14701);
nor U14971 (N_14971,N_14772,N_14832);
xnor U14972 (N_14972,N_14835,N_14796);
xor U14973 (N_14973,N_14838,N_14726);
or U14974 (N_14974,N_14821,N_14734);
nor U14975 (N_14975,N_14710,N_14802);
nand U14976 (N_14976,N_14791,N_14842);
nand U14977 (N_14977,N_14715,N_14820);
and U14978 (N_14978,N_14761,N_14781);
or U14979 (N_14979,N_14777,N_14767);
and U14980 (N_14980,N_14804,N_14842);
nor U14981 (N_14981,N_14758,N_14742);
xnor U14982 (N_14982,N_14743,N_14759);
nor U14983 (N_14983,N_14769,N_14754);
or U14984 (N_14984,N_14735,N_14803);
nand U14985 (N_14985,N_14810,N_14813);
xor U14986 (N_14986,N_14774,N_14820);
xnor U14987 (N_14987,N_14770,N_14848);
nor U14988 (N_14988,N_14832,N_14750);
or U14989 (N_14989,N_14734,N_14792);
nand U14990 (N_14990,N_14795,N_14747);
nand U14991 (N_14991,N_14745,N_14704);
xnor U14992 (N_14992,N_14812,N_14719);
and U14993 (N_14993,N_14839,N_14750);
nor U14994 (N_14994,N_14828,N_14734);
or U14995 (N_14995,N_14799,N_14842);
xor U14996 (N_14996,N_14767,N_14724);
and U14997 (N_14997,N_14838,N_14817);
nor U14998 (N_14998,N_14834,N_14839);
and U14999 (N_14999,N_14820,N_14829);
xor UO_0 (O_0,N_14893,N_14915);
nor UO_1 (O_1,N_14985,N_14866);
or UO_2 (O_2,N_14862,N_14956);
xnor UO_3 (O_3,N_14886,N_14954);
or UO_4 (O_4,N_14879,N_14968);
or UO_5 (O_5,N_14897,N_14878);
or UO_6 (O_6,N_14980,N_14967);
or UO_7 (O_7,N_14913,N_14908);
or UO_8 (O_8,N_14939,N_14871);
and UO_9 (O_9,N_14923,N_14944);
and UO_10 (O_10,N_14912,N_14995);
xor UO_11 (O_11,N_14941,N_14896);
and UO_12 (O_12,N_14924,N_14952);
and UO_13 (O_13,N_14957,N_14929);
nor UO_14 (O_14,N_14977,N_14988);
nand UO_15 (O_15,N_14970,N_14986);
or UO_16 (O_16,N_14940,N_14934);
and UO_17 (O_17,N_14855,N_14919);
and UO_18 (O_18,N_14895,N_14892);
and UO_19 (O_19,N_14991,N_14917);
or UO_20 (O_20,N_14960,N_14853);
nor UO_21 (O_21,N_14906,N_14933);
xnor UO_22 (O_22,N_14935,N_14876);
nor UO_23 (O_23,N_14958,N_14950);
nor UO_24 (O_24,N_14880,N_14877);
and UO_25 (O_25,N_14922,N_14998);
or UO_26 (O_26,N_14850,N_14945);
or UO_27 (O_27,N_14851,N_14969);
or UO_28 (O_28,N_14987,N_14872);
nor UO_29 (O_29,N_14860,N_14927);
or UO_30 (O_30,N_14955,N_14888);
and UO_31 (O_31,N_14914,N_14999);
and UO_32 (O_32,N_14993,N_14964);
and UO_33 (O_33,N_14965,N_14947);
xnor UO_34 (O_34,N_14931,N_14982);
or UO_35 (O_35,N_14979,N_14894);
xnor UO_36 (O_36,N_14902,N_14859);
nand UO_37 (O_37,N_14884,N_14920);
nor UO_38 (O_38,N_14854,N_14910);
nor UO_39 (O_39,N_14904,N_14861);
xnor UO_40 (O_40,N_14921,N_14891);
nand UO_41 (O_41,N_14949,N_14996);
nor UO_42 (O_42,N_14881,N_14946);
xor UO_43 (O_43,N_14926,N_14887);
nand UO_44 (O_44,N_14953,N_14948);
and UO_45 (O_45,N_14959,N_14885);
and UO_46 (O_46,N_14905,N_14990);
xnor UO_47 (O_47,N_14882,N_14962);
nor UO_48 (O_48,N_14869,N_14873);
and UO_49 (O_49,N_14973,N_14972);
nand UO_50 (O_50,N_14981,N_14870);
xor UO_51 (O_51,N_14978,N_14932);
nor UO_52 (O_52,N_14864,N_14966);
nand UO_53 (O_53,N_14916,N_14961);
or UO_54 (O_54,N_14907,N_14858);
nand UO_55 (O_55,N_14868,N_14865);
and UO_56 (O_56,N_14976,N_14903);
or UO_57 (O_57,N_14983,N_14989);
xnor UO_58 (O_58,N_14936,N_14928);
nor UO_59 (O_59,N_14984,N_14937);
nand UO_60 (O_60,N_14857,N_14856);
nor UO_61 (O_61,N_14899,N_14943);
or UO_62 (O_62,N_14994,N_14900);
and UO_63 (O_63,N_14867,N_14925);
nand UO_64 (O_64,N_14883,N_14890);
nor UO_65 (O_65,N_14963,N_14951);
xor UO_66 (O_66,N_14975,N_14863);
nand UO_67 (O_67,N_14898,N_14889);
or UO_68 (O_68,N_14911,N_14901);
and UO_69 (O_69,N_14938,N_14918);
xor UO_70 (O_70,N_14875,N_14930);
or UO_71 (O_71,N_14874,N_14997);
xnor UO_72 (O_72,N_14992,N_14909);
nand UO_73 (O_73,N_14974,N_14971);
xor UO_74 (O_74,N_14942,N_14852);
nand UO_75 (O_75,N_14913,N_14967);
or UO_76 (O_76,N_14874,N_14962);
nand UO_77 (O_77,N_14872,N_14972);
xnor UO_78 (O_78,N_14907,N_14900);
and UO_79 (O_79,N_14998,N_14871);
nand UO_80 (O_80,N_14953,N_14975);
and UO_81 (O_81,N_14930,N_14867);
nor UO_82 (O_82,N_14872,N_14916);
nor UO_83 (O_83,N_14982,N_14954);
or UO_84 (O_84,N_14964,N_14851);
nand UO_85 (O_85,N_14872,N_14931);
nand UO_86 (O_86,N_14864,N_14979);
nor UO_87 (O_87,N_14897,N_14885);
xor UO_88 (O_88,N_14948,N_14961);
or UO_89 (O_89,N_14922,N_14899);
nand UO_90 (O_90,N_14941,N_14992);
nor UO_91 (O_91,N_14899,N_14961);
xnor UO_92 (O_92,N_14922,N_14912);
nand UO_93 (O_93,N_14853,N_14979);
and UO_94 (O_94,N_14904,N_14867);
nand UO_95 (O_95,N_14976,N_14918);
nand UO_96 (O_96,N_14887,N_14985);
nor UO_97 (O_97,N_14856,N_14862);
xor UO_98 (O_98,N_14955,N_14914);
nand UO_99 (O_99,N_14939,N_14988);
nand UO_100 (O_100,N_14862,N_14937);
nor UO_101 (O_101,N_14951,N_14970);
nand UO_102 (O_102,N_14932,N_14917);
or UO_103 (O_103,N_14949,N_14863);
or UO_104 (O_104,N_14947,N_14956);
or UO_105 (O_105,N_14926,N_14989);
nor UO_106 (O_106,N_14944,N_14958);
and UO_107 (O_107,N_14938,N_14852);
or UO_108 (O_108,N_14941,N_14907);
nor UO_109 (O_109,N_14992,N_14907);
and UO_110 (O_110,N_14882,N_14938);
nor UO_111 (O_111,N_14936,N_14960);
nand UO_112 (O_112,N_14955,N_14895);
xnor UO_113 (O_113,N_14867,N_14854);
and UO_114 (O_114,N_14981,N_14877);
and UO_115 (O_115,N_14860,N_14912);
or UO_116 (O_116,N_14983,N_14932);
xnor UO_117 (O_117,N_14938,N_14946);
nor UO_118 (O_118,N_14910,N_14972);
nand UO_119 (O_119,N_14879,N_14997);
nor UO_120 (O_120,N_14853,N_14918);
or UO_121 (O_121,N_14868,N_14904);
or UO_122 (O_122,N_14967,N_14867);
or UO_123 (O_123,N_14871,N_14866);
xnor UO_124 (O_124,N_14966,N_14883);
xor UO_125 (O_125,N_14977,N_14984);
xnor UO_126 (O_126,N_14946,N_14890);
nor UO_127 (O_127,N_14947,N_14940);
nor UO_128 (O_128,N_14977,N_14914);
xor UO_129 (O_129,N_14976,N_14948);
or UO_130 (O_130,N_14940,N_14860);
nand UO_131 (O_131,N_14946,N_14875);
xnor UO_132 (O_132,N_14918,N_14902);
nor UO_133 (O_133,N_14865,N_14863);
nand UO_134 (O_134,N_14901,N_14970);
xnor UO_135 (O_135,N_14854,N_14869);
nor UO_136 (O_136,N_14865,N_14953);
or UO_137 (O_137,N_14918,N_14921);
nor UO_138 (O_138,N_14896,N_14903);
or UO_139 (O_139,N_14922,N_14913);
xor UO_140 (O_140,N_14914,N_14850);
or UO_141 (O_141,N_14954,N_14883);
nand UO_142 (O_142,N_14850,N_14890);
and UO_143 (O_143,N_14861,N_14920);
nand UO_144 (O_144,N_14952,N_14939);
or UO_145 (O_145,N_14895,N_14925);
nand UO_146 (O_146,N_14921,N_14902);
or UO_147 (O_147,N_14970,N_14875);
and UO_148 (O_148,N_14961,N_14921);
or UO_149 (O_149,N_14931,N_14976);
nor UO_150 (O_150,N_14970,N_14859);
xnor UO_151 (O_151,N_14891,N_14945);
nand UO_152 (O_152,N_14883,N_14913);
nand UO_153 (O_153,N_14866,N_14914);
nor UO_154 (O_154,N_14857,N_14884);
xnor UO_155 (O_155,N_14997,N_14971);
and UO_156 (O_156,N_14879,N_14861);
nand UO_157 (O_157,N_14899,N_14927);
or UO_158 (O_158,N_14869,N_14907);
or UO_159 (O_159,N_14880,N_14896);
or UO_160 (O_160,N_14893,N_14867);
and UO_161 (O_161,N_14946,N_14913);
nor UO_162 (O_162,N_14876,N_14955);
xnor UO_163 (O_163,N_14927,N_14997);
nand UO_164 (O_164,N_14929,N_14926);
nor UO_165 (O_165,N_14981,N_14904);
or UO_166 (O_166,N_14894,N_14916);
nand UO_167 (O_167,N_14952,N_14856);
xor UO_168 (O_168,N_14897,N_14892);
xnor UO_169 (O_169,N_14901,N_14881);
nand UO_170 (O_170,N_14913,N_14919);
and UO_171 (O_171,N_14997,N_14982);
nor UO_172 (O_172,N_14916,N_14863);
nand UO_173 (O_173,N_14910,N_14924);
or UO_174 (O_174,N_14922,N_14856);
nand UO_175 (O_175,N_14954,N_14919);
nor UO_176 (O_176,N_14859,N_14869);
and UO_177 (O_177,N_14865,N_14896);
nor UO_178 (O_178,N_14902,N_14900);
xnor UO_179 (O_179,N_14878,N_14916);
or UO_180 (O_180,N_14936,N_14943);
nand UO_181 (O_181,N_14962,N_14897);
nor UO_182 (O_182,N_14939,N_14869);
and UO_183 (O_183,N_14992,N_14863);
nand UO_184 (O_184,N_14920,N_14958);
and UO_185 (O_185,N_14957,N_14900);
nand UO_186 (O_186,N_14977,N_14994);
nand UO_187 (O_187,N_14911,N_14986);
nor UO_188 (O_188,N_14987,N_14855);
xnor UO_189 (O_189,N_14862,N_14977);
or UO_190 (O_190,N_14941,N_14933);
nor UO_191 (O_191,N_14945,N_14957);
and UO_192 (O_192,N_14978,N_14955);
or UO_193 (O_193,N_14920,N_14875);
nor UO_194 (O_194,N_14873,N_14990);
or UO_195 (O_195,N_14928,N_14856);
xor UO_196 (O_196,N_14965,N_14983);
xnor UO_197 (O_197,N_14857,N_14961);
or UO_198 (O_198,N_14944,N_14955);
nand UO_199 (O_199,N_14906,N_14981);
or UO_200 (O_200,N_14912,N_14921);
and UO_201 (O_201,N_14906,N_14970);
and UO_202 (O_202,N_14940,N_14856);
xnor UO_203 (O_203,N_14948,N_14943);
nor UO_204 (O_204,N_14891,N_14906);
or UO_205 (O_205,N_14953,N_14850);
nor UO_206 (O_206,N_14992,N_14948);
xnor UO_207 (O_207,N_14901,N_14961);
nor UO_208 (O_208,N_14949,N_14966);
and UO_209 (O_209,N_14867,N_14929);
or UO_210 (O_210,N_14953,N_14983);
and UO_211 (O_211,N_14961,N_14897);
and UO_212 (O_212,N_14944,N_14896);
or UO_213 (O_213,N_14947,N_14911);
nor UO_214 (O_214,N_14883,N_14855);
or UO_215 (O_215,N_14904,N_14866);
nor UO_216 (O_216,N_14980,N_14944);
and UO_217 (O_217,N_14904,N_14978);
and UO_218 (O_218,N_14987,N_14969);
nand UO_219 (O_219,N_14938,N_14968);
or UO_220 (O_220,N_14922,N_14916);
or UO_221 (O_221,N_14891,N_14857);
or UO_222 (O_222,N_14975,N_14880);
nor UO_223 (O_223,N_14927,N_14974);
and UO_224 (O_224,N_14905,N_14918);
nand UO_225 (O_225,N_14901,N_14891);
or UO_226 (O_226,N_14919,N_14861);
and UO_227 (O_227,N_14945,N_14916);
or UO_228 (O_228,N_14869,N_14892);
xnor UO_229 (O_229,N_14989,N_14909);
and UO_230 (O_230,N_14922,N_14923);
and UO_231 (O_231,N_14893,N_14883);
nand UO_232 (O_232,N_14949,N_14895);
or UO_233 (O_233,N_14881,N_14976);
or UO_234 (O_234,N_14957,N_14914);
nor UO_235 (O_235,N_14891,N_14974);
nand UO_236 (O_236,N_14970,N_14896);
nor UO_237 (O_237,N_14954,N_14851);
nor UO_238 (O_238,N_14895,N_14916);
and UO_239 (O_239,N_14898,N_14924);
or UO_240 (O_240,N_14900,N_14979);
nand UO_241 (O_241,N_14905,N_14989);
or UO_242 (O_242,N_14921,N_14936);
xor UO_243 (O_243,N_14862,N_14869);
nand UO_244 (O_244,N_14996,N_14925);
and UO_245 (O_245,N_14964,N_14933);
nand UO_246 (O_246,N_14994,N_14941);
nand UO_247 (O_247,N_14997,N_14975);
nand UO_248 (O_248,N_14904,N_14999);
nand UO_249 (O_249,N_14992,N_14935);
and UO_250 (O_250,N_14905,N_14909);
or UO_251 (O_251,N_14887,N_14990);
xnor UO_252 (O_252,N_14963,N_14925);
xor UO_253 (O_253,N_14876,N_14856);
nor UO_254 (O_254,N_14926,N_14962);
or UO_255 (O_255,N_14958,N_14886);
or UO_256 (O_256,N_14964,N_14984);
or UO_257 (O_257,N_14962,N_14898);
xor UO_258 (O_258,N_14887,N_14936);
or UO_259 (O_259,N_14933,N_14869);
and UO_260 (O_260,N_14926,N_14964);
xnor UO_261 (O_261,N_14924,N_14945);
nand UO_262 (O_262,N_14979,N_14940);
or UO_263 (O_263,N_14982,N_14951);
nand UO_264 (O_264,N_14903,N_14973);
xnor UO_265 (O_265,N_14855,N_14973);
nand UO_266 (O_266,N_14985,N_14933);
nand UO_267 (O_267,N_14894,N_14901);
or UO_268 (O_268,N_14903,N_14907);
nor UO_269 (O_269,N_14925,N_14898);
nand UO_270 (O_270,N_14916,N_14860);
or UO_271 (O_271,N_14954,N_14946);
or UO_272 (O_272,N_14974,N_14903);
and UO_273 (O_273,N_14920,N_14893);
nand UO_274 (O_274,N_14917,N_14938);
nor UO_275 (O_275,N_14993,N_14903);
nor UO_276 (O_276,N_14882,N_14863);
or UO_277 (O_277,N_14917,N_14883);
and UO_278 (O_278,N_14986,N_14889);
nand UO_279 (O_279,N_14865,N_14966);
xor UO_280 (O_280,N_14920,N_14934);
nor UO_281 (O_281,N_14974,N_14869);
nor UO_282 (O_282,N_14960,N_14856);
or UO_283 (O_283,N_14898,N_14934);
and UO_284 (O_284,N_14922,N_14853);
or UO_285 (O_285,N_14975,N_14983);
xnor UO_286 (O_286,N_14965,N_14996);
nand UO_287 (O_287,N_14966,N_14925);
xnor UO_288 (O_288,N_14863,N_14892);
nor UO_289 (O_289,N_14931,N_14951);
nand UO_290 (O_290,N_14941,N_14900);
nand UO_291 (O_291,N_14910,N_14870);
or UO_292 (O_292,N_14903,N_14970);
or UO_293 (O_293,N_14903,N_14877);
or UO_294 (O_294,N_14852,N_14850);
nand UO_295 (O_295,N_14988,N_14873);
nand UO_296 (O_296,N_14965,N_14978);
nand UO_297 (O_297,N_14969,N_14912);
nand UO_298 (O_298,N_14973,N_14928);
nand UO_299 (O_299,N_14965,N_14970);
nor UO_300 (O_300,N_14956,N_14857);
nand UO_301 (O_301,N_14985,N_14879);
xnor UO_302 (O_302,N_14971,N_14891);
xnor UO_303 (O_303,N_14998,N_14882);
and UO_304 (O_304,N_14994,N_14929);
nor UO_305 (O_305,N_14907,N_14996);
xor UO_306 (O_306,N_14945,N_14952);
nand UO_307 (O_307,N_14963,N_14913);
xnor UO_308 (O_308,N_14966,N_14901);
xnor UO_309 (O_309,N_14924,N_14872);
nor UO_310 (O_310,N_14871,N_14888);
xor UO_311 (O_311,N_14985,N_14964);
xor UO_312 (O_312,N_14866,N_14957);
nor UO_313 (O_313,N_14908,N_14906);
and UO_314 (O_314,N_14944,N_14960);
and UO_315 (O_315,N_14991,N_14877);
and UO_316 (O_316,N_14901,N_14932);
nand UO_317 (O_317,N_14905,N_14946);
and UO_318 (O_318,N_14911,N_14895);
nor UO_319 (O_319,N_14852,N_14944);
xor UO_320 (O_320,N_14953,N_14967);
nand UO_321 (O_321,N_14915,N_14875);
or UO_322 (O_322,N_14908,N_14950);
and UO_323 (O_323,N_14883,N_14981);
and UO_324 (O_324,N_14979,N_14912);
nand UO_325 (O_325,N_14916,N_14854);
nand UO_326 (O_326,N_14876,N_14966);
xor UO_327 (O_327,N_14935,N_14895);
and UO_328 (O_328,N_14851,N_14929);
nor UO_329 (O_329,N_14982,N_14857);
nor UO_330 (O_330,N_14925,N_14938);
or UO_331 (O_331,N_14927,N_14888);
nand UO_332 (O_332,N_14981,N_14990);
or UO_333 (O_333,N_14902,N_14956);
xnor UO_334 (O_334,N_14954,N_14976);
and UO_335 (O_335,N_14996,N_14913);
nand UO_336 (O_336,N_14984,N_14860);
xor UO_337 (O_337,N_14859,N_14901);
xor UO_338 (O_338,N_14997,N_14906);
or UO_339 (O_339,N_14936,N_14922);
nand UO_340 (O_340,N_14947,N_14945);
nor UO_341 (O_341,N_14934,N_14883);
and UO_342 (O_342,N_14893,N_14986);
or UO_343 (O_343,N_14976,N_14962);
and UO_344 (O_344,N_14953,N_14876);
nor UO_345 (O_345,N_14875,N_14975);
xnor UO_346 (O_346,N_14971,N_14939);
nand UO_347 (O_347,N_14994,N_14979);
or UO_348 (O_348,N_14921,N_14991);
nor UO_349 (O_349,N_14907,N_14934);
or UO_350 (O_350,N_14883,N_14896);
nand UO_351 (O_351,N_14896,N_14940);
xnor UO_352 (O_352,N_14911,N_14981);
nand UO_353 (O_353,N_14885,N_14865);
and UO_354 (O_354,N_14962,N_14935);
and UO_355 (O_355,N_14928,N_14908);
nand UO_356 (O_356,N_14935,N_14936);
or UO_357 (O_357,N_14857,N_14920);
or UO_358 (O_358,N_14973,N_14958);
or UO_359 (O_359,N_14905,N_14949);
and UO_360 (O_360,N_14903,N_14893);
or UO_361 (O_361,N_14890,N_14991);
nor UO_362 (O_362,N_14960,N_14894);
and UO_363 (O_363,N_14931,N_14855);
or UO_364 (O_364,N_14927,N_14850);
and UO_365 (O_365,N_14856,N_14934);
nor UO_366 (O_366,N_14854,N_14967);
nand UO_367 (O_367,N_14865,N_14939);
xnor UO_368 (O_368,N_14875,N_14879);
nand UO_369 (O_369,N_14910,N_14943);
nand UO_370 (O_370,N_14999,N_14877);
nor UO_371 (O_371,N_14873,N_14985);
or UO_372 (O_372,N_14967,N_14973);
and UO_373 (O_373,N_14968,N_14975);
xnor UO_374 (O_374,N_14976,N_14939);
nor UO_375 (O_375,N_14872,N_14995);
or UO_376 (O_376,N_14957,N_14861);
and UO_377 (O_377,N_14985,N_14894);
nor UO_378 (O_378,N_14991,N_14927);
and UO_379 (O_379,N_14989,N_14979);
nor UO_380 (O_380,N_14993,N_14969);
or UO_381 (O_381,N_14977,N_14899);
or UO_382 (O_382,N_14950,N_14941);
or UO_383 (O_383,N_14972,N_14999);
and UO_384 (O_384,N_14867,N_14974);
and UO_385 (O_385,N_14944,N_14890);
xnor UO_386 (O_386,N_14933,N_14927);
nand UO_387 (O_387,N_14850,N_14908);
or UO_388 (O_388,N_14987,N_14866);
xor UO_389 (O_389,N_14899,N_14945);
xor UO_390 (O_390,N_14877,N_14987);
xnor UO_391 (O_391,N_14982,N_14921);
nor UO_392 (O_392,N_14899,N_14964);
or UO_393 (O_393,N_14927,N_14887);
nand UO_394 (O_394,N_14872,N_14998);
or UO_395 (O_395,N_14988,N_14926);
xor UO_396 (O_396,N_14965,N_14875);
or UO_397 (O_397,N_14881,N_14855);
nor UO_398 (O_398,N_14850,N_14977);
xor UO_399 (O_399,N_14985,N_14988);
nand UO_400 (O_400,N_14917,N_14967);
nor UO_401 (O_401,N_14969,N_14926);
nor UO_402 (O_402,N_14876,N_14992);
or UO_403 (O_403,N_14896,N_14943);
and UO_404 (O_404,N_14992,N_14951);
or UO_405 (O_405,N_14867,N_14977);
xor UO_406 (O_406,N_14863,N_14936);
and UO_407 (O_407,N_14925,N_14914);
nor UO_408 (O_408,N_14913,N_14860);
or UO_409 (O_409,N_14969,N_14966);
nor UO_410 (O_410,N_14953,N_14916);
xor UO_411 (O_411,N_14940,N_14889);
nand UO_412 (O_412,N_14884,N_14982);
nand UO_413 (O_413,N_14981,N_14872);
or UO_414 (O_414,N_14905,N_14883);
nor UO_415 (O_415,N_14903,N_14908);
or UO_416 (O_416,N_14933,N_14942);
nand UO_417 (O_417,N_14907,N_14914);
and UO_418 (O_418,N_14902,N_14898);
or UO_419 (O_419,N_14964,N_14909);
nor UO_420 (O_420,N_14943,N_14937);
nand UO_421 (O_421,N_14961,N_14895);
or UO_422 (O_422,N_14992,N_14969);
and UO_423 (O_423,N_14986,N_14937);
nor UO_424 (O_424,N_14878,N_14937);
or UO_425 (O_425,N_14946,N_14936);
xor UO_426 (O_426,N_14918,N_14895);
and UO_427 (O_427,N_14865,N_14999);
nor UO_428 (O_428,N_14994,N_14870);
or UO_429 (O_429,N_14947,N_14981);
and UO_430 (O_430,N_14996,N_14862);
or UO_431 (O_431,N_14976,N_14973);
or UO_432 (O_432,N_14946,N_14934);
xor UO_433 (O_433,N_14891,N_14911);
nor UO_434 (O_434,N_14884,N_14888);
and UO_435 (O_435,N_14913,N_14962);
or UO_436 (O_436,N_14898,N_14964);
and UO_437 (O_437,N_14989,N_14904);
xnor UO_438 (O_438,N_14958,N_14933);
nand UO_439 (O_439,N_14995,N_14868);
or UO_440 (O_440,N_14930,N_14876);
xor UO_441 (O_441,N_14953,N_14886);
xnor UO_442 (O_442,N_14909,N_14874);
nand UO_443 (O_443,N_14947,N_14884);
and UO_444 (O_444,N_14946,N_14959);
nor UO_445 (O_445,N_14908,N_14988);
or UO_446 (O_446,N_14991,N_14964);
or UO_447 (O_447,N_14950,N_14990);
xor UO_448 (O_448,N_14931,N_14913);
or UO_449 (O_449,N_14902,N_14932);
or UO_450 (O_450,N_14998,N_14890);
and UO_451 (O_451,N_14931,N_14857);
xor UO_452 (O_452,N_14916,N_14870);
or UO_453 (O_453,N_14951,N_14915);
xor UO_454 (O_454,N_14991,N_14853);
or UO_455 (O_455,N_14933,N_14955);
xor UO_456 (O_456,N_14974,N_14973);
nand UO_457 (O_457,N_14901,N_14903);
and UO_458 (O_458,N_14947,N_14942);
nor UO_459 (O_459,N_14990,N_14901);
or UO_460 (O_460,N_14879,N_14863);
and UO_461 (O_461,N_14891,N_14879);
and UO_462 (O_462,N_14928,N_14870);
nand UO_463 (O_463,N_14910,N_14932);
and UO_464 (O_464,N_14992,N_14981);
or UO_465 (O_465,N_14961,N_14954);
xor UO_466 (O_466,N_14969,N_14910);
nand UO_467 (O_467,N_14852,N_14990);
and UO_468 (O_468,N_14929,N_14976);
nand UO_469 (O_469,N_14869,N_14998);
nand UO_470 (O_470,N_14921,N_14875);
and UO_471 (O_471,N_14898,N_14955);
nor UO_472 (O_472,N_14871,N_14970);
xnor UO_473 (O_473,N_14872,N_14876);
or UO_474 (O_474,N_14850,N_14899);
xor UO_475 (O_475,N_14886,N_14923);
nor UO_476 (O_476,N_14883,N_14887);
xnor UO_477 (O_477,N_14859,N_14985);
xor UO_478 (O_478,N_14919,N_14868);
and UO_479 (O_479,N_14919,N_14850);
or UO_480 (O_480,N_14854,N_14984);
and UO_481 (O_481,N_14872,N_14943);
xor UO_482 (O_482,N_14994,N_14955);
nand UO_483 (O_483,N_14933,N_14934);
nor UO_484 (O_484,N_14942,N_14950);
nor UO_485 (O_485,N_14968,N_14861);
and UO_486 (O_486,N_14997,N_14891);
xor UO_487 (O_487,N_14951,N_14984);
or UO_488 (O_488,N_14876,N_14901);
nor UO_489 (O_489,N_14935,N_14954);
and UO_490 (O_490,N_14999,N_14891);
nor UO_491 (O_491,N_14946,N_14891);
xnor UO_492 (O_492,N_14947,N_14870);
nor UO_493 (O_493,N_14924,N_14965);
nand UO_494 (O_494,N_14899,N_14983);
and UO_495 (O_495,N_14914,N_14919);
xnor UO_496 (O_496,N_14883,N_14923);
nor UO_497 (O_497,N_14957,N_14963);
nor UO_498 (O_498,N_14918,N_14975);
nand UO_499 (O_499,N_14937,N_14996);
nand UO_500 (O_500,N_14926,N_14851);
and UO_501 (O_501,N_14992,N_14875);
nor UO_502 (O_502,N_14981,N_14958);
or UO_503 (O_503,N_14892,N_14914);
xor UO_504 (O_504,N_14895,N_14857);
xor UO_505 (O_505,N_14959,N_14956);
xor UO_506 (O_506,N_14999,N_14893);
xnor UO_507 (O_507,N_14972,N_14996);
nor UO_508 (O_508,N_14924,N_14950);
xor UO_509 (O_509,N_14895,N_14878);
nor UO_510 (O_510,N_14851,N_14864);
nand UO_511 (O_511,N_14961,N_14929);
nand UO_512 (O_512,N_14894,N_14942);
and UO_513 (O_513,N_14875,N_14996);
xor UO_514 (O_514,N_14872,N_14884);
nand UO_515 (O_515,N_14891,N_14919);
xor UO_516 (O_516,N_14978,N_14894);
nor UO_517 (O_517,N_14917,N_14924);
nor UO_518 (O_518,N_14924,N_14862);
nand UO_519 (O_519,N_14911,N_14950);
nand UO_520 (O_520,N_14992,N_14917);
or UO_521 (O_521,N_14854,N_14949);
and UO_522 (O_522,N_14869,N_14992);
nor UO_523 (O_523,N_14888,N_14901);
nand UO_524 (O_524,N_14904,N_14851);
nand UO_525 (O_525,N_14904,N_14901);
and UO_526 (O_526,N_14893,N_14950);
nand UO_527 (O_527,N_14930,N_14872);
or UO_528 (O_528,N_14912,N_14861);
nor UO_529 (O_529,N_14855,N_14864);
nor UO_530 (O_530,N_14988,N_14854);
nand UO_531 (O_531,N_14879,N_14938);
and UO_532 (O_532,N_14938,N_14993);
or UO_533 (O_533,N_14934,N_14905);
nor UO_534 (O_534,N_14962,N_14977);
xnor UO_535 (O_535,N_14982,N_14883);
xnor UO_536 (O_536,N_14963,N_14966);
nand UO_537 (O_537,N_14853,N_14872);
and UO_538 (O_538,N_14934,N_14893);
nor UO_539 (O_539,N_14914,N_14983);
xor UO_540 (O_540,N_14997,N_14921);
xnor UO_541 (O_541,N_14974,N_14944);
xor UO_542 (O_542,N_14949,N_14993);
xor UO_543 (O_543,N_14883,N_14986);
and UO_544 (O_544,N_14976,N_14862);
and UO_545 (O_545,N_14988,N_14944);
nand UO_546 (O_546,N_14945,N_14864);
or UO_547 (O_547,N_14987,N_14880);
nor UO_548 (O_548,N_14890,N_14977);
or UO_549 (O_549,N_14918,N_14954);
xnor UO_550 (O_550,N_14989,N_14924);
nand UO_551 (O_551,N_14928,N_14948);
xor UO_552 (O_552,N_14851,N_14908);
or UO_553 (O_553,N_14856,N_14865);
xnor UO_554 (O_554,N_14896,N_14911);
nor UO_555 (O_555,N_14992,N_14868);
xor UO_556 (O_556,N_14868,N_14857);
and UO_557 (O_557,N_14957,N_14960);
xnor UO_558 (O_558,N_14861,N_14860);
or UO_559 (O_559,N_14917,N_14931);
nor UO_560 (O_560,N_14939,N_14984);
and UO_561 (O_561,N_14877,N_14957);
xor UO_562 (O_562,N_14867,N_14926);
nand UO_563 (O_563,N_14910,N_14906);
nor UO_564 (O_564,N_14953,N_14909);
or UO_565 (O_565,N_14891,N_14865);
and UO_566 (O_566,N_14893,N_14960);
nor UO_567 (O_567,N_14860,N_14985);
xnor UO_568 (O_568,N_14877,N_14955);
nor UO_569 (O_569,N_14951,N_14978);
xnor UO_570 (O_570,N_14946,N_14861);
xnor UO_571 (O_571,N_14996,N_14885);
nand UO_572 (O_572,N_14947,N_14933);
nor UO_573 (O_573,N_14908,N_14991);
xnor UO_574 (O_574,N_14932,N_14897);
nand UO_575 (O_575,N_14901,N_14853);
or UO_576 (O_576,N_14955,N_14935);
nor UO_577 (O_577,N_14854,N_14865);
or UO_578 (O_578,N_14918,N_14970);
nor UO_579 (O_579,N_14982,N_14871);
nor UO_580 (O_580,N_14995,N_14975);
and UO_581 (O_581,N_14869,N_14900);
nor UO_582 (O_582,N_14943,N_14922);
nor UO_583 (O_583,N_14862,N_14904);
or UO_584 (O_584,N_14856,N_14992);
nor UO_585 (O_585,N_14971,N_14935);
xor UO_586 (O_586,N_14957,N_14860);
nor UO_587 (O_587,N_14889,N_14904);
nor UO_588 (O_588,N_14914,N_14929);
nand UO_589 (O_589,N_14998,N_14893);
and UO_590 (O_590,N_14973,N_14963);
or UO_591 (O_591,N_14967,N_14930);
nand UO_592 (O_592,N_14996,N_14864);
nand UO_593 (O_593,N_14913,N_14899);
nand UO_594 (O_594,N_14868,N_14887);
or UO_595 (O_595,N_14941,N_14987);
xor UO_596 (O_596,N_14948,N_14996);
nand UO_597 (O_597,N_14977,N_14971);
and UO_598 (O_598,N_14980,N_14919);
nand UO_599 (O_599,N_14937,N_14989);
nand UO_600 (O_600,N_14925,N_14936);
or UO_601 (O_601,N_14891,N_14867);
or UO_602 (O_602,N_14995,N_14947);
xor UO_603 (O_603,N_14920,N_14969);
nor UO_604 (O_604,N_14916,N_14947);
xnor UO_605 (O_605,N_14891,N_14980);
nand UO_606 (O_606,N_14922,N_14930);
xor UO_607 (O_607,N_14896,N_14964);
or UO_608 (O_608,N_14865,N_14883);
or UO_609 (O_609,N_14897,N_14880);
or UO_610 (O_610,N_14994,N_14931);
and UO_611 (O_611,N_14915,N_14924);
nor UO_612 (O_612,N_14896,N_14933);
nor UO_613 (O_613,N_14936,N_14944);
xnor UO_614 (O_614,N_14937,N_14902);
or UO_615 (O_615,N_14896,N_14957);
or UO_616 (O_616,N_14969,N_14951);
nor UO_617 (O_617,N_14883,N_14900);
xor UO_618 (O_618,N_14877,N_14978);
nand UO_619 (O_619,N_14952,N_14921);
nand UO_620 (O_620,N_14900,N_14913);
and UO_621 (O_621,N_14952,N_14979);
nor UO_622 (O_622,N_14969,N_14872);
nand UO_623 (O_623,N_14899,N_14937);
or UO_624 (O_624,N_14996,N_14935);
or UO_625 (O_625,N_14866,N_14925);
nand UO_626 (O_626,N_14861,N_14871);
nor UO_627 (O_627,N_14850,N_14888);
xor UO_628 (O_628,N_14913,N_14951);
and UO_629 (O_629,N_14901,N_14871);
xnor UO_630 (O_630,N_14963,N_14921);
nand UO_631 (O_631,N_14897,N_14890);
nor UO_632 (O_632,N_14862,N_14886);
nor UO_633 (O_633,N_14978,N_14969);
or UO_634 (O_634,N_14856,N_14902);
nand UO_635 (O_635,N_14999,N_14940);
nor UO_636 (O_636,N_14988,N_14995);
nand UO_637 (O_637,N_14919,N_14870);
or UO_638 (O_638,N_14953,N_14962);
nor UO_639 (O_639,N_14990,N_14955);
xor UO_640 (O_640,N_14873,N_14976);
xnor UO_641 (O_641,N_14904,N_14855);
nor UO_642 (O_642,N_14911,N_14985);
nor UO_643 (O_643,N_14850,N_14990);
and UO_644 (O_644,N_14991,N_14909);
xor UO_645 (O_645,N_14886,N_14968);
xor UO_646 (O_646,N_14985,N_14861);
xor UO_647 (O_647,N_14860,N_14934);
or UO_648 (O_648,N_14922,N_14891);
or UO_649 (O_649,N_14992,N_14945);
and UO_650 (O_650,N_14960,N_14948);
or UO_651 (O_651,N_14912,N_14886);
xnor UO_652 (O_652,N_14921,N_14929);
and UO_653 (O_653,N_14866,N_14867);
nor UO_654 (O_654,N_14904,N_14863);
xor UO_655 (O_655,N_14955,N_14951);
nor UO_656 (O_656,N_14981,N_14936);
nor UO_657 (O_657,N_14902,N_14862);
and UO_658 (O_658,N_14917,N_14970);
nand UO_659 (O_659,N_14888,N_14981);
and UO_660 (O_660,N_14994,N_14858);
nand UO_661 (O_661,N_14993,N_14999);
or UO_662 (O_662,N_14997,N_14883);
nand UO_663 (O_663,N_14973,N_14870);
xor UO_664 (O_664,N_14871,N_14995);
xnor UO_665 (O_665,N_14962,N_14990);
xnor UO_666 (O_666,N_14987,N_14909);
and UO_667 (O_667,N_14888,N_14868);
or UO_668 (O_668,N_14964,N_14871);
or UO_669 (O_669,N_14920,N_14930);
and UO_670 (O_670,N_14916,N_14969);
or UO_671 (O_671,N_14871,N_14851);
and UO_672 (O_672,N_14980,N_14966);
or UO_673 (O_673,N_14871,N_14854);
nor UO_674 (O_674,N_14873,N_14858);
xnor UO_675 (O_675,N_14928,N_14930);
or UO_676 (O_676,N_14870,N_14902);
or UO_677 (O_677,N_14884,N_14954);
and UO_678 (O_678,N_14986,N_14868);
or UO_679 (O_679,N_14950,N_14932);
or UO_680 (O_680,N_14994,N_14876);
nor UO_681 (O_681,N_14901,N_14865);
and UO_682 (O_682,N_14942,N_14962);
xnor UO_683 (O_683,N_14930,N_14866);
or UO_684 (O_684,N_14939,N_14960);
xnor UO_685 (O_685,N_14989,N_14966);
or UO_686 (O_686,N_14861,N_14974);
nor UO_687 (O_687,N_14935,N_14984);
nor UO_688 (O_688,N_14974,N_14871);
xor UO_689 (O_689,N_14982,N_14971);
xnor UO_690 (O_690,N_14988,N_14980);
xor UO_691 (O_691,N_14898,N_14993);
nor UO_692 (O_692,N_14941,N_14923);
nor UO_693 (O_693,N_14878,N_14902);
or UO_694 (O_694,N_14858,N_14909);
xnor UO_695 (O_695,N_14864,N_14927);
or UO_696 (O_696,N_14880,N_14891);
nor UO_697 (O_697,N_14931,N_14956);
and UO_698 (O_698,N_14892,N_14962);
and UO_699 (O_699,N_14873,N_14957);
or UO_700 (O_700,N_14943,N_14851);
or UO_701 (O_701,N_14899,N_14882);
nand UO_702 (O_702,N_14986,N_14961);
and UO_703 (O_703,N_14878,N_14985);
or UO_704 (O_704,N_14938,N_14873);
nand UO_705 (O_705,N_14941,N_14960);
nor UO_706 (O_706,N_14920,N_14879);
nor UO_707 (O_707,N_14940,N_14914);
or UO_708 (O_708,N_14857,N_14870);
nand UO_709 (O_709,N_14890,N_14964);
or UO_710 (O_710,N_14851,N_14869);
nand UO_711 (O_711,N_14912,N_14887);
xor UO_712 (O_712,N_14999,N_14925);
nand UO_713 (O_713,N_14919,N_14948);
xnor UO_714 (O_714,N_14968,N_14898);
and UO_715 (O_715,N_14967,N_14997);
or UO_716 (O_716,N_14975,N_14864);
nor UO_717 (O_717,N_14997,N_14936);
nand UO_718 (O_718,N_14924,N_14998);
nand UO_719 (O_719,N_14952,N_14907);
xor UO_720 (O_720,N_14902,N_14941);
nor UO_721 (O_721,N_14910,N_14963);
nand UO_722 (O_722,N_14936,N_14986);
and UO_723 (O_723,N_14922,N_14992);
nor UO_724 (O_724,N_14988,N_14955);
and UO_725 (O_725,N_14866,N_14859);
xnor UO_726 (O_726,N_14913,N_14999);
nor UO_727 (O_727,N_14984,N_14973);
xnor UO_728 (O_728,N_14859,N_14922);
nor UO_729 (O_729,N_14966,N_14908);
nor UO_730 (O_730,N_14997,N_14898);
nor UO_731 (O_731,N_14920,N_14916);
or UO_732 (O_732,N_14886,N_14910);
nor UO_733 (O_733,N_14881,N_14941);
nand UO_734 (O_734,N_14905,N_14954);
or UO_735 (O_735,N_14907,N_14997);
and UO_736 (O_736,N_14983,N_14907);
nand UO_737 (O_737,N_14978,N_14961);
or UO_738 (O_738,N_14907,N_14945);
nor UO_739 (O_739,N_14853,N_14913);
and UO_740 (O_740,N_14892,N_14918);
nor UO_741 (O_741,N_14947,N_14975);
xnor UO_742 (O_742,N_14927,N_14983);
xnor UO_743 (O_743,N_14948,N_14994);
xor UO_744 (O_744,N_14996,N_14979);
and UO_745 (O_745,N_14964,N_14893);
nor UO_746 (O_746,N_14969,N_14927);
xnor UO_747 (O_747,N_14990,N_14952);
and UO_748 (O_748,N_14855,N_14936);
and UO_749 (O_749,N_14871,N_14885);
or UO_750 (O_750,N_14974,N_14983);
nor UO_751 (O_751,N_14902,N_14971);
or UO_752 (O_752,N_14952,N_14978);
or UO_753 (O_753,N_14857,N_14947);
and UO_754 (O_754,N_14857,N_14963);
nor UO_755 (O_755,N_14934,N_14965);
and UO_756 (O_756,N_14861,N_14939);
or UO_757 (O_757,N_14928,N_14922);
and UO_758 (O_758,N_14852,N_14882);
nand UO_759 (O_759,N_14905,N_14950);
nor UO_760 (O_760,N_14854,N_14902);
xor UO_761 (O_761,N_14919,N_14858);
or UO_762 (O_762,N_14948,N_14969);
xor UO_763 (O_763,N_14975,N_14858);
xor UO_764 (O_764,N_14945,N_14932);
or UO_765 (O_765,N_14949,N_14873);
nor UO_766 (O_766,N_14921,N_14932);
nor UO_767 (O_767,N_14902,N_14899);
nor UO_768 (O_768,N_14966,N_14861);
nand UO_769 (O_769,N_14994,N_14940);
xnor UO_770 (O_770,N_14998,N_14953);
nand UO_771 (O_771,N_14930,N_14956);
or UO_772 (O_772,N_14870,N_14899);
and UO_773 (O_773,N_14858,N_14952);
nor UO_774 (O_774,N_14874,N_14897);
nor UO_775 (O_775,N_14887,N_14991);
nand UO_776 (O_776,N_14984,N_14884);
nand UO_777 (O_777,N_14946,N_14972);
nand UO_778 (O_778,N_14850,N_14893);
nor UO_779 (O_779,N_14914,N_14927);
and UO_780 (O_780,N_14908,N_14972);
nor UO_781 (O_781,N_14861,N_14915);
and UO_782 (O_782,N_14972,N_14896);
xnor UO_783 (O_783,N_14964,N_14916);
xor UO_784 (O_784,N_14933,N_14905);
or UO_785 (O_785,N_14938,N_14865);
nand UO_786 (O_786,N_14879,N_14967);
nand UO_787 (O_787,N_14943,N_14912);
or UO_788 (O_788,N_14919,N_14942);
nor UO_789 (O_789,N_14936,N_14913);
xnor UO_790 (O_790,N_14942,N_14926);
and UO_791 (O_791,N_14971,N_14989);
or UO_792 (O_792,N_14944,N_14919);
xnor UO_793 (O_793,N_14935,N_14958);
xor UO_794 (O_794,N_14935,N_14923);
and UO_795 (O_795,N_14885,N_14957);
and UO_796 (O_796,N_14991,N_14978);
nor UO_797 (O_797,N_14879,N_14986);
and UO_798 (O_798,N_14947,N_14957);
or UO_799 (O_799,N_14896,N_14974);
xnor UO_800 (O_800,N_14969,N_14980);
nand UO_801 (O_801,N_14942,N_14925);
xor UO_802 (O_802,N_14891,N_14937);
nor UO_803 (O_803,N_14968,N_14990);
and UO_804 (O_804,N_14867,N_14918);
nand UO_805 (O_805,N_14875,N_14874);
xnor UO_806 (O_806,N_14894,N_14948);
and UO_807 (O_807,N_14865,N_14852);
or UO_808 (O_808,N_14934,N_14855);
xnor UO_809 (O_809,N_14952,N_14859);
xor UO_810 (O_810,N_14875,N_14895);
and UO_811 (O_811,N_14944,N_14928);
xnor UO_812 (O_812,N_14966,N_14999);
and UO_813 (O_813,N_14978,N_14917);
or UO_814 (O_814,N_14900,N_14858);
and UO_815 (O_815,N_14987,N_14958);
nor UO_816 (O_816,N_14965,N_14891);
nor UO_817 (O_817,N_14889,N_14881);
nor UO_818 (O_818,N_14965,N_14881);
xnor UO_819 (O_819,N_14897,N_14956);
xor UO_820 (O_820,N_14976,N_14940);
xor UO_821 (O_821,N_14918,N_14972);
nor UO_822 (O_822,N_14889,N_14875);
and UO_823 (O_823,N_14906,N_14862);
nor UO_824 (O_824,N_14855,N_14893);
and UO_825 (O_825,N_14955,N_14931);
xor UO_826 (O_826,N_14874,N_14990);
xor UO_827 (O_827,N_14907,N_14995);
xnor UO_828 (O_828,N_14984,N_14946);
nor UO_829 (O_829,N_14985,N_14998);
or UO_830 (O_830,N_14870,N_14940);
nor UO_831 (O_831,N_14904,N_14873);
xnor UO_832 (O_832,N_14883,N_14977);
xnor UO_833 (O_833,N_14874,N_14988);
or UO_834 (O_834,N_14887,N_14908);
or UO_835 (O_835,N_14862,N_14880);
and UO_836 (O_836,N_14906,N_14996);
xor UO_837 (O_837,N_14948,N_14949);
and UO_838 (O_838,N_14967,N_14990);
or UO_839 (O_839,N_14955,N_14952);
or UO_840 (O_840,N_14907,N_14991);
or UO_841 (O_841,N_14863,N_14978);
nand UO_842 (O_842,N_14866,N_14901);
nor UO_843 (O_843,N_14875,N_14880);
nand UO_844 (O_844,N_14881,N_14988);
nor UO_845 (O_845,N_14979,N_14867);
or UO_846 (O_846,N_14958,N_14954);
nor UO_847 (O_847,N_14859,N_14987);
and UO_848 (O_848,N_14973,N_14953);
or UO_849 (O_849,N_14868,N_14907);
xnor UO_850 (O_850,N_14965,N_14957);
or UO_851 (O_851,N_14887,N_14878);
and UO_852 (O_852,N_14892,N_14969);
or UO_853 (O_853,N_14905,N_14962);
nor UO_854 (O_854,N_14976,N_14941);
nor UO_855 (O_855,N_14898,N_14922);
nor UO_856 (O_856,N_14980,N_14904);
xnor UO_857 (O_857,N_14949,N_14906);
and UO_858 (O_858,N_14863,N_14875);
or UO_859 (O_859,N_14974,N_14884);
or UO_860 (O_860,N_14900,N_14939);
xor UO_861 (O_861,N_14942,N_14995);
and UO_862 (O_862,N_14924,N_14963);
nor UO_863 (O_863,N_14984,N_14875);
or UO_864 (O_864,N_14895,N_14964);
nor UO_865 (O_865,N_14935,N_14993);
nand UO_866 (O_866,N_14915,N_14955);
xnor UO_867 (O_867,N_14934,N_14918);
nand UO_868 (O_868,N_14886,N_14872);
xnor UO_869 (O_869,N_14980,N_14868);
and UO_870 (O_870,N_14937,N_14910);
or UO_871 (O_871,N_14975,N_14943);
and UO_872 (O_872,N_14865,N_14918);
or UO_873 (O_873,N_14911,N_14922);
xnor UO_874 (O_874,N_14974,N_14928);
nand UO_875 (O_875,N_14891,N_14855);
nand UO_876 (O_876,N_14879,N_14960);
or UO_877 (O_877,N_14898,N_14929);
xor UO_878 (O_878,N_14940,N_14941);
and UO_879 (O_879,N_14911,N_14944);
and UO_880 (O_880,N_14977,N_14957);
nor UO_881 (O_881,N_14948,N_14959);
and UO_882 (O_882,N_14933,N_14851);
nand UO_883 (O_883,N_14894,N_14904);
nor UO_884 (O_884,N_14906,N_14988);
and UO_885 (O_885,N_14850,N_14915);
or UO_886 (O_886,N_14886,N_14966);
nand UO_887 (O_887,N_14914,N_14879);
and UO_888 (O_888,N_14994,N_14888);
nor UO_889 (O_889,N_14924,N_14973);
nand UO_890 (O_890,N_14981,N_14946);
or UO_891 (O_891,N_14950,N_14895);
xnor UO_892 (O_892,N_14858,N_14996);
and UO_893 (O_893,N_14892,N_14977);
and UO_894 (O_894,N_14916,N_14970);
xor UO_895 (O_895,N_14983,N_14923);
nor UO_896 (O_896,N_14964,N_14956);
xnor UO_897 (O_897,N_14921,N_14907);
nand UO_898 (O_898,N_14983,N_14898);
or UO_899 (O_899,N_14876,N_14939);
nor UO_900 (O_900,N_14924,N_14889);
and UO_901 (O_901,N_14989,N_14930);
and UO_902 (O_902,N_14865,N_14920);
and UO_903 (O_903,N_14882,N_14985);
nand UO_904 (O_904,N_14879,N_14924);
nand UO_905 (O_905,N_14920,N_14983);
nor UO_906 (O_906,N_14977,N_14989);
and UO_907 (O_907,N_14882,N_14862);
xnor UO_908 (O_908,N_14876,N_14866);
xnor UO_909 (O_909,N_14968,N_14997);
xnor UO_910 (O_910,N_14975,N_14859);
nand UO_911 (O_911,N_14994,N_14919);
or UO_912 (O_912,N_14945,N_14946);
or UO_913 (O_913,N_14857,N_14957);
nand UO_914 (O_914,N_14922,N_14909);
nand UO_915 (O_915,N_14941,N_14852);
nor UO_916 (O_916,N_14981,N_14869);
nand UO_917 (O_917,N_14989,N_14986);
or UO_918 (O_918,N_14850,N_14903);
or UO_919 (O_919,N_14866,N_14907);
nor UO_920 (O_920,N_14995,N_14922);
nor UO_921 (O_921,N_14896,N_14986);
xnor UO_922 (O_922,N_14850,N_14873);
nand UO_923 (O_923,N_14973,N_14964);
or UO_924 (O_924,N_14947,N_14974);
and UO_925 (O_925,N_14865,N_14955);
and UO_926 (O_926,N_14887,N_14915);
nand UO_927 (O_927,N_14991,N_14898);
nor UO_928 (O_928,N_14986,N_14912);
and UO_929 (O_929,N_14909,N_14984);
nand UO_930 (O_930,N_14964,N_14912);
or UO_931 (O_931,N_14984,N_14938);
nand UO_932 (O_932,N_14982,N_14936);
and UO_933 (O_933,N_14985,N_14967);
nand UO_934 (O_934,N_14873,N_14887);
xor UO_935 (O_935,N_14932,N_14988);
or UO_936 (O_936,N_14880,N_14950);
or UO_937 (O_937,N_14936,N_14891);
nand UO_938 (O_938,N_14927,N_14879);
nand UO_939 (O_939,N_14924,N_14904);
nor UO_940 (O_940,N_14915,N_14863);
or UO_941 (O_941,N_14987,N_14925);
or UO_942 (O_942,N_14936,N_14961);
nand UO_943 (O_943,N_14871,N_14997);
xnor UO_944 (O_944,N_14858,N_14915);
nor UO_945 (O_945,N_14960,N_14890);
and UO_946 (O_946,N_14915,N_14929);
xnor UO_947 (O_947,N_14974,N_14960);
or UO_948 (O_948,N_14981,N_14862);
nand UO_949 (O_949,N_14907,N_14930);
nand UO_950 (O_950,N_14975,N_14922);
xor UO_951 (O_951,N_14901,N_14882);
nand UO_952 (O_952,N_14851,N_14924);
and UO_953 (O_953,N_14927,N_14912);
xnor UO_954 (O_954,N_14855,N_14991);
or UO_955 (O_955,N_14980,N_14893);
xnor UO_956 (O_956,N_14988,N_14942);
nand UO_957 (O_957,N_14879,N_14934);
and UO_958 (O_958,N_14951,N_14925);
nand UO_959 (O_959,N_14888,N_14957);
nor UO_960 (O_960,N_14854,N_14939);
nor UO_961 (O_961,N_14907,N_14933);
nand UO_962 (O_962,N_14999,N_14866);
nand UO_963 (O_963,N_14888,N_14940);
or UO_964 (O_964,N_14950,N_14885);
xor UO_965 (O_965,N_14893,N_14924);
or UO_966 (O_966,N_14861,N_14956);
xnor UO_967 (O_967,N_14855,N_14879);
and UO_968 (O_968,N_14881,N_14864);
nor UO_969 (O_969,N_14909,N_14911);
and UO_970 (O_970,N_14919,N_14983);
and UO_971 (O_971,N_14866,N_14869);
xor UO_972 (O_972,N_14954,N_14875);
and UO_973 (O_973,N_14922,N_14895);
and UO_974 (O_974,N_14985,N_14970);
or UO_975 (O_975,N_14982,N_14900);
xor UO_976 (O_976,N_14888,N_14895);
nand UO_977 (O_977,N_14965,N_14960);
nand UO_978 (O_978,N_14853,N_14912);
xor UO_979 (O_979,N_14893,N_14982);
and UO_980 (O_980,N_14961,N_14940);
nand UO_981 (O_981,N_14879,N_14964);
and UO_982 (O_982,N_14864,N_14917);
xnor UO_983 (O_983,N_14980,N_14863);
and UO_984 (O_984,N_14852,N_14883);
or UO_985 (O_985,N_14858,N_14918);
and UO_986 (O_986,N_14951,N_14908);
and UO_987 (O_987,N_14887,N_14989);
and UO_988 (O_988,N_14939,N_14974);
nor UO_989 (O_989,N_14978,N_14851);
or UO_990 (O_990,N_14906,N_14878);
xnor UO_991 (O_991,N_14914,N_14985);
nand UO_992 (O_992,N_14965,N_14926);
xnor UO_993 (O_993,N_14936,N_14938);
or UO_994 (O_994,N_14889,N_14887);
nor UO_995 (O_995,N_14927,N_14902);
or UO_996 (O_996,N_14969,N_14930);
xor UO_997 (O_997,N_14895,N_14980);
nand UO_998 (O_998,N_14964,N_14920);
nand UO_999 (O_999,N_14910,N_14948);
or UO_1000 (O_1000,N_14928,N_14888);
or UO_1001 (O_1001,N_14856,N_14901);
or UO_1002 (O_1002,N_14925,N_14879);
nand UO_1003 (O_1003,N_14995,N_14905);
nor UO_1004 (O_1004,N_14988,N_14966);
xor UO_1005 (O_1005,N_14960,N_14857);
nand UO_1006 (O_1006,N_14963,N_14881);
nor UO_1007 (O_1007,N_14940,N_14875);
xor UO_1008 (O_1008,N_14993,N_14926);
nand UO_1009 (O_1009,N_14920,N_14944);
or UO_1010 (O_1010,N_14999,N_14983);
and UO_1011 (O_1011,N_14862,N_14878);
or UO_1012 (O_1012,N_14899,N_14919);
xor UO_1013 (O_1013,N_14914,N_14984);
xor UO_1014 (O_1014,N_14966,N_14874);
xor UO_1015 (O_1015,N_14991,N_14944);
or UO_1016 (O_1016,N_14894,N_14919);
and UO_1017 (O_1017,N_14972,N_14945);
nand UO_1018 (O_1018,N_14971,N_14962);
and UO_1019 (O_1019,N_14984,N_14956);
nand UO_1020 (O_1020,N_14860,N_14881);
and UO_1021 (O_1021,N_14999,N_14857);
and UO_1022 (O_1022,N_14930,N_14941);
nand UO_1023 (O_1023,N_14978,N_14939);
nor UO_1024 (O_1024,N_14926,N_14894);
and UO_1025 (O_1025,N_14856,N_14957);
xor UO_1026 (O_1026,N_14966,N_14879);
xor UO_1027 (O_1027,N_14851,N_14963);
nand UO_1028 (O_1028,N_14853,N_14983);
xnor UO_1029 (O_1029,N_14878,N_14876);
and UO_1030 (O_1030,N_14925,N_14892);
and UO_1031 (O_1031,N_14890,N_14990);
nor UO_1032 (O_1032,N_14936,N_14881);
and UO_1033 (O_1033,N_14904,N_14977);
nand UO_1034 (O_1034,N_14925,N_14947);
or UO_1035 (O_1035,N_14958,N_14966);
nor UO_1036 (O_1036,N_14884,N_14921);
xnor UO_1037 (O_1037,N_14981,N_14975);
nand UO_1038 (O_1038,N_14944,N_14956);
or UO_1039 (O_1039,N_14882,N_14916);
xnor UO_1040 (O_1040,N_14970,N_14889);
or UO_1041 (O_1041,N_14900,N_14867);
nor UO_1042 (O_1042,N_14873,N_14909);
nand UO_1043 (O_1043,N_14934,N_14925);
nor UO_1044 (O_1044,N_14912,N_14881);
nand UO_1045 (O_1045,N_14866,N_14889);
and UO_1046 (O_1046,N_14926,N_14990);
or UO_1047 (O_1047,N_14933,N_14936);
nor UO_1048 (O_1048,N_14956,N_14880);
nor UO_1049 (O_1049,N_14952,N_14912);
nor UO_1050 (O_1050,N_14867,N_14998);
or UO_1051 (O_1051,N_14862,N_14850);
or UO_1052 (O_1052,N_14914,N_14996);
or UO_1053 (O_1053,N_14887,N_14892);
nor UO_1054 (O_1054,N_14990,N_14857);
nor UO_1055 (O_1055,N_14943,N_14892);
nand UO_1056 (O_1056,N_14990,N_14951);
nand UO_1057 (O_1057,N_14941,N_14858);
or UO_1058 (O_1058,N_14958,N_14869);
nor UO_1059 (O_1059,N_14999,N_14854);
nor UO_1060 (O_1060,N_14884,N_14985);
and UO_1061 (O_1061,N_14872,N_14898);
and UO_1062 (O_1062,N_14928,N_14885);
and UO_1063 (O_1063,N_14963,N_14944);
and UO_1064 (O_1064,N_14995,N_14866);
nor UO_1065 (O_1065,N_14900,N_14856);
xnor UO_1066 (O_1066,N_14955,N_14916);
nand UO_1067 (O_1067,N_14979,N_14902);
and UO_1068 (O_1068,N_14990,N_14975);
and UO_1069 (O_1069,N_14902,N_14962);
and UO_1070 (O_1070,N_14927,N_14916);
nand UO_1071 (O_1071,N_14855,N_14902);
and UO_1072 (O_1072,N_14912,N_14945);
or UO_1073 (O_1073,N_14889,N_14996);
and UO_1074 (O_1074,N_14986,N_14885);
xnor UO_1075 (O_1075,N_14924,N_14921);
nand UO_1076 (O_1076,N_14945,N_14950);
or UO_1077 (O_1077,N_14958,N_14899);
nand UO_1078 (O_1078,N_14937,N_14979);
or UO_1079 (O_1079,N_14916,N_14886);
nand UO_1080 (O_1080,N_14876,N_14945);
or UO_1081 (O_1081,N_14902,N_14992);
or UO_1082 (O_1082,N_14986,N_14858);
or UO_1083 (O_1083,N_14895,N_14903);
nor UO_1084 (O_1084,N_14954,N_14908);
nor UO_1085 (O_1085,N_14918,N_14875);
nand UO_1086 (O_1086,N_14854,N_14872);
and UO_1087 (O_1087,N_14860,N_14959);
xnor UO_1088 (O_1088,N_14891,N_14967);
nor UO_1089 (O_1089,N_14943,N_14984);
or UO_1090 (O_1090,N_14917,N_14899);
xnor UO_1091 (O_1091,N_14934,N_14921);
nor UO_1092 (O_1092,N_14921,N_14977);
nor UO_1093 (O_1093,N_14969,N_14925);
and UO_1094 (O_1094,N_14886,N_14944);
or UO_1095 (O_1095,N_14915,N_14971);
nand UO_1096 (O_1096,N_14890,N_14951);
nor UO_1097 (O_1097,N_14942,N_14952);
and UO_1098 (O_1098,N_14911,N_14942);
or UO_1099 (O_1099,N_14907,N_14888);
and UO_1100 (O_1100,N_14891,N_14850);
nand UO_1101 (O_1101,N_14898,N_14915);
nor UO_1102 (O_1102,N_14930,N_14903);
and UO_1103 (O_1103,N_14852,N_14980);
nand UO_1104 (O_1104,N_14961,N_14903);
xor UO_1105 (O_1105,N_14913,N_14937);
and UO_1106 (O_1106,N_14900,N_14945);
xor UO_1107 (O_1107,N_14917,N_14881);
nor UO_1108 (O_1108,N_14992,N_14895);
or UO_1109 (O_1109,N_14883,N_14984);
and UO_1110 (O_1110,N_14972,N_14995);
nor UO_1111 (O_1111,N_14976,N_14850);
nor UO_1112 (O_1112,N_14933,N_14944);
or UO_1113 (O_1113,N_14991,N_14941);
xnor UO_1114 (O_1114,N_14945,N_14858);
xnor UO_1115 (O_1115,N_14962,N_14862);
nor UO_1116 (O_1116,N_14867,N_14860);
and UO_1117 (O_1117,N_14855,N_14986);
nor UO_1118 (O_1118,N_14898,N_14858);
and UO_1119 (O_1119,N_14924,N_14966);
nor UO_1120 (O_1120,N_14996,N_14967);
or UO_1121 (O_1121,N_14963,N_14912);
xnor UO_1122 (O_1122,N_14963,N_14915);
xor UO_1123 (O_1123,N_14866,N_14893);
and UO_1124 (O_1124,N_14982,N_14926);
and UO_1125 (O_1125,N_14886,N_14873);
nand UO_1126 (O_1126,N_14981,N_14942);
nor UO_1127 (O_1127,N_14973,N_14887);
xor UO_1128 (O_1128,N_14859,N_14860);
and UO_1129 (O_1129,N_14863,N_14989);
nand UO_1130 (O_1130,N_14961,N_14910);
nor UO_1131 (O_1131,N_14935,N_14874);
and UO_1132 (O_1132,N_14978,N_14910);
and UO_1133 (O_1133,N_14897,N_14953);
nor UO_1134 (O_1134,N_14885,N_14989);
nor UO_1135 (O_1135,N_14851,N_14940);
xor UO_1136 (O_1136,N_14926,N_14961);
and UO_1137 (O_1137,N_14949,N_14980);
nand UO_1138 (O_1138,N_14982,N_14909);
or UO_1139 (O_1139,N_14903,N_14935);
xor UO_1140 (O_1140,N_14944,N_14925);
xnor UO_1141 (O_1141,N_14976,N_14945);
or UO_1142 (O_1142,N_14956,N_14925);
or UO_1143 (O_1143,N_14945,N_14898);
nor UO_1144 (O_1144,N_14994,N_14992);
nand UO_1145 (O_1145,N_14927,N_14876);
or UO_1146 (O_1146,N_14917,N_14962);
nand UO_1147 (O_1147,N_14850,N_14901);
nor UO_1148 (O_1148,N_14958,N_14866);
nand UO_1149 (O_1149,N_14966,N_14944);
or UO_1150 (O_1150,N_14924,N_14946);
nand UO_1151 (O_1151,N_14863,N_14891);
and UO_1152 (O_1152,N_14987,N_14918);
and UO_1153 (O_1153,N_14948,N_14967);
nand UO_1154 (O_1154,N_14942,N_14903);
nand UO_1155 (O_1155,N_14973,N_14875);
and UO_1156 (O_1156,N_14976,N_14921);
and UO_1157 (O_1157,N_14957,N_14946);
xor UO_1158 (O_1158,N_14977,N_14901);
or UO_1159 (O_1159,N_14897,N_14906);
or UO_1160 (O_1160,N_14985,N_14955);
xnor UO_1161 (O_1161,N_14869,N_14989);
nand UO_1162 (O_1162,N_14983,N_14941);
xor UO_1163 (O_1163,N_14999,N_14922);
or UO_1164 (O_1164,N_14956,N_14903);
or UO_1165 (O_1165,N_14953,N_14990);
xor UO_1166 (O_1166,N_14870,N_14882);
and UO_1167 (O_1167,N_14964,N_14885);
or UO_1168 (O_1168,N_14916,N_14885);
nand UO_1169 (O_1169,N_14989,N_14911);
and UO_1170 (O_1170,N_14947,N_14982);
nor UO_1171 (O_1171,N_14924,N_14858);
or UO_1172 (O_1172,N_14903,N_14860);
or UO_1173 (O_1173,N_14955,N_14857);
or UO_1174 (O_1174,N_14906,N_14873);
xor UO_1175 (O_1175,N_14918,N_14965);
and UO_1176 (O_1176,N_14948,N_14988);
and UO_1177 (O_1177,N_14857,N_14877);
nor UO_1178 (O_1178,N_14996,N_14876);
nand UO_1179 (O_1179,N_14866,N_14936);
or UO_1180 (O_1180,N_14912,N_14928);
or UO_1181 (O_1181,N_14890,N_14904);
and UO_1182 (O_1182,N_14989,N_14938);
nor UO_1183 (O_1183,N_14979,N_14929);
nor UO_1184 (O_1184,N_14951,N_14987);
nand UO_1185 (O_1185,N_14919,N_14889);
and UO_1186 (O_1186,N_14930,N_14880);
and UO_1187 (O_1187,N_14874,N_14888);
or UO_1188 (O_1188,N_14878,N_14894);
nor UO_1189 (O_1189,N_14917,N_14910);
and UO_1190 (O_1190,N_14886,N_14881);
or UO_1191 (O_1191,N_14944,N_14968);
and UO_1192 (O_1192,N_14995,N_14946);
or UO_1193 (O_1193,N_14982,N_14867);
and UO_1194 (O_1194,N_14989,N_14947);
xnor UO_1195 (O_1195,N_14956,N_14954);
xnor UO_1196 (O_1196,N_14892,N_14950);
nor UO_1197 (O_1197,N_14933,N_14948);
nor UO_1198 (O_1198,N_14913,N_14930);
nand UO_1199 (O_1199,N_14985,N_14917);
nor UO_1200 (O_1200,N_14852,N_14950);
and UO_1201 (O_1201,N_14945,N_14869);
or UO_1202 (O_1202,N_14962,N_14867);
nand UO_1203 (O_1203,N_14964,N_14853);
nor UO_1204 (O_1204,N_14891,N_14887);
nor UO_1205 (O_1205,N_14860,N_14942);
nand UO_1206 (O_1206,N_14909,N_14950);
or UO_1207 (O_1207,N_14961,N_14970);
nor UO_1208 (O_1208,N_14971,N_14897);
nand UO_1209 (O_1209,N_14976,N_14978);
nand UO_1210 (O_1210,N_14954,N_14945);
and UO_1211 (O_1211,N_14891,N_14878);
or UO_1212 (O_1212,N_14904,N_14917);
xor UO_1213 (O_1213,N_14877,N_14960);
nor UO_1214 (O_1214,N_14867,N_14949);
or UO_1215 (O_1215,N_14949,N_14992);
nand UO_1216 (O_1216,N_14920,N_14999);
nor UO_1217 (O_1217,N_14915,N_14901);
nand UO_1218 (O_1218,N_14857,N_14976);
xnor UO_1219 (O_1219,N_14940,N_14984);
or UO_1220 (O_1220,N_14971,N_14870);
and UO_1221 (O_1221,N_14941,N_14958);
nand UO_1222 (O_1222,N_14874,N_14936);
xnor UO_1223 (O_1223,N_14990,N_14974);
or UO_1224 (O_1224,N_14984,N_14868);
nand UO_1225 (O_1225,N_14977,N_14920);
and UO_1226 (O_1226,N_14851,N_14905);
or UO_1227 (O_1227,N_14913,N_14968);
and UO_1228 (O_1228,N_14965,N_14878);
and UO_1229 (O_1229,N_14854,N_14954);
and UO_1230 (O_1230,N_14914,N_14890);
nand UO_1231 (O_1231,N_14927,N_14922);
nand UO_1232 (O_1232,N_14930,N_14898);
nor UO_1233 (O_1233,N_14968,N_14974);
nor UO_1234 (O_1234,N_14979,N_14934);
nand UO_1235 (O_1235,N_14871,N_14860);
nor UO_1236 (O_1236,N_14944,N_14967);
and UO_1237 (O_1237,N_14869,N_14909);
nor UO_1238 (O_1238,N_14882,N_14868);
and UO_1239 (O_1239,N_14967,N_14999);
nor UO_1240 (O_1240,N_14905,N_14971);
nor UO_1241 (O_1241,N_14907,N_14859);
nand UO_1242 (O_1242,N_14929,N_14932);
or UO_1243 (O_1243,N_14873,N_14861);
nor UO_1244 (O_1244,N_14927,N_14911);
and UO_1245 (O_1245,N_14983,N_14895);
or UO_1246 (O_1246,N_14928,N_14881);
nor UO_1247 (O_1247,N_14965,N_14861);
nor UO_1248 (O_1248,N_14905,N_14940);
or UO_1249 (O_1249,N_14876,N_14851);
xnor UO_1250 (O_1250,N_14999,N_14901);
and UO_1251 (O_1251,N_14873,N_14961);
or UO_1252 (O_1252,N_14964,N_14927);
and UO_1253 (O_1253,N_14942,N_14886);
nor UO_1254 (O_1254,N_14998,N_14988);
nor UO_1255 (O_1255,N_14969,N_14999);
nand UO_1256 (O_1256,N_14890,N_14898);
nor UO_1257 (O_1257,N_14972,N_14903);
nand UO_1258 (O_1258,N_14850,N_14943);
and UO_1259 (O_1259,N_14971,N_14926);
nor UO_1260 (O_1260,N_14910,N_14980);
xor UO_1261 (O_1261,N_14900,N_14937);
nor UO_1262 (O_1262,N_14898,N_14873);
nor UO_1263 (O_1263,N_14921,N_14958);
xnor UO_1264 (O_1264,N_14946,N_14868);
nor UO_1265 (O_1265,N_14895,N_14933);
or UO_1266 (O_1266,N_14896,N_14884);
nand UO_1267 (O_1267,N_14881,N_14959);
xnor UO_1268 (O_1268,N_14906,N_14992);
or UO_1269 (O_1269,N_14938,N_14900);
and UO_1270 (O_1270,N_14970,N_14934);
nand UO_1271 (O_1271,N_14964,N_14935);
xnor UO_1272 (O_1272,N_14909,N_14887);
or UO_1273 (O_1273,N_14907,N_14959);
and UO_1274 (O_1274,N_14884,N_14998);
or UO_1275 (O_1275,N_14863,N_14964);
and UO_1276 (O_1276,N_14883,N_14963);
nor UO_1277 (O_1277,N_14950,N_14959);
xnor UO_1278 (O_1278,N_14974,N_14914);
nand UO_1279 (O_1279,N_14880,N_14869);
or UO_1280 (O_1280,N_14954,N_14962);
nand UO_1281 (O_1281,N_14952,N_14937);
nor UO_1282 (O_1282,N_14896,N_14915);
nand UO_1283 (O_1283,N_14991,N_14888);
or UO_1284 (O_1284,N_14899,N_14992);
nor UO_1285 (O_1285,N_14887,N_14937);
or UO_1286 (O_1286,N_14927,N_14999);
nor UO_1287 (O_1287,N_14994,N_14946);
or UO_1288 (O_1288,N_14910,N_14982);
or UO_1289 (O_1289,N_14949,N_14857);
nor UO_1290 (O_1290,N_14878,N_14948);
and UO_1291 (O_1291,N_14914,N_14933);
or UO_1292 (O_1292,N_14882,N_14856);
or UO_1293 (O_1293,N_14873,N_14951);
xor UO_1294 (O_1294,N_14940,N_14943);
or UO_1295 (O_1295,N_14913,N_14986);
and UO_1296 (O_1296,N_14917,N_14861);
nor UO_1297 (O_1297,N_14871,N_14904);
xnor UO_1298 (O_1298,N_14894,N_14860);
nand UO_1299 (O_1299,N_14888,N_14947);
nand UO_1300 (O_1300,N_14927,N_14923);
xnor UO_1301 (O_1301,N_14941,N_14868);
nand UO_1302 (O_1302,N_14874,N_14866);
and UO_1303 (O_1303,N_14900,N_14966);
nand UO_1304 (O_1304,N_14861,N_14994);
or UO_1305 (O_1305,N_14890,N_14877);
xor UO_1306 (O_1306,N_14881,N_14967);
nor UO_1307 (O_1307,N_14912,N_14999);
or UO_1308 (O_1308,N_14955,N_14991);
or UO_1309 (O_1309,N_14875,N_14959);
or UO_1310 (O_1310,N_14913,N_14918);
and UO_1311 (O_1311,N_14934,N_14876);
nor UO_1312 (O_1312,N_14939,N_14895);
xor UO_1313 (O_1313,N_14874,N_14984);
or UO_1314 (O_1314,N_14917,N_14905);
or UO_1315 (O_1315,N_14863,N_14969);
and UO_1316 (O_1316,N_14932,N_14937);
nor UO_1317 (O_1317,N_14868,N_14908);
and UO_1318 (O_1318,N_14870,N_14930);
xor UO_1319 (O_1319,N_14900,N_14926);
and UO_1320 (O_1320,N_14890,N_14992);
nor UO_1321 (O_1321,N_14903,N_14985);
nor UO_1322 (O_1322,N_14922,N_14963);
nor UO_1323 (O_1323,N_14897,N_14859);
nand UO_1324 (O_1324,N_14860,N_14998);
nor UO_1325 (O_1325,N_14873,N_14923);
nand UO_1326 (O_1326,N_14874,N_14902);
and UO_1327 (O_1327,N_14958,N_14971);
xor UO_1328 (O_1328,N_14863,N_14905);
and UO_1329 (O_1329,N_14914,N_14969);
nor UO_1330 (O_1330,N_14920,N_14927);
or UO_1331 (O_1331,N_14909,N_14914);
xor UO_1332 (O_1332,N_14923,N_14893);
xnor UO_1333 (O_1333,N_14954,N_14926);
nor UO_1334 (O_1334,N_14866,N_14945);
or UO_1335 (O_1335,N_14890,N_14901);
xnor UO_1336 (O_1336,N_14864,N_14911);
nor UO_1337 (O_1337,N_14974,N_14888);
or UO_1338 (O_1338,N_14856,N_14913);
nand UO_1339 (O_1339,N_14926,N_14959);
xor UO_1340 (O_1340,N_14874,N_14937);
nor UO_1341 (O_1341,N_14918,N_14857);
xor UO_1342 (O_1342,N_14858,N_14932);
and UO_1343 (O_1343,N_14916,N_14949);
xnor UO_1344 (O_1344,N_14888,N_14929);
nor UO_1345 (O_1345,N_14973,N_14891);
nand UO_1346 (O_1346,N_14906,N_14971);
nand UO_1347 (O_1347,N_14954,N_14989);
and UO_1348 (O_1348,N_14973,N_14996);
xor UO_1349 (O_1349,N_14872,N_14852);
or UO_1350 (O_1350,N_14914,N_14982);
nand UO_1351 (O_1351,N_14956,N_14932);
and UO_1352 (O_1352,N_14913,N_14994);
nand UO_1353 (O_1353,N_14858,N_14888);
nor UO_1354 (O_1354,N_14914,N_14908);
xor UO_1355 (O_1355,N_14878,N_14917);
and UO_1356 (O_1356,N_14973,N_14857);
or UO_1357 (O_1357,N_14982,N_14860);
xnor UO_1358 (O_1358,N_14978,N_14869);
nor UO_1359 (O_1359,N_14981,N_14941);
nor UO_1360 (O_1360,N_14925,N_14857);
nor UO_1361 (O_1361,N_14865,N_14873);
xnor UO_1362 (O_1362,N_14912,N_14917);
nor UO_1363 (O_1363,N_14950,N_14863);
nand UO_1364 (O_1364,N_14910,N_14875);
xnor UO_1365 (O_1365,N_14930,N_14993);
nand UO_1366 (O_1366,N_14886,N_14949);
nor UO_1367 (O_1367,N_14999,N_14946);
xor UO_1368 (O_1368,N_14964,N_14883);
nor UO_1369 (O_1369,N_14851,N_14874);
and UO_1370 (O_1370,N_14969,N_14891);
nor UO_1371 (O_1371,N_14980,N_14871);
nor UO_1372 (O_1372,N_14894,N_14900);
or UO_1373 (O_1373,N_14914,N_14880);
nand UO_1374 (O_1374,N_14958,N_14851);
xnor UO_1375 (O_1375,N_14910,N_14964);
and UO_1376 (O_1376,N_14967,N_14979);
and UO_1377 (O_1377,N_14877,N_14868);
nand UO_1378 (O_1378,N_14903,N_14931);
nor UO_1379 (O_1379,N_14889,N_14864);
and UO_1380 (O_1380,N_14901,N_14923);
or UO_1381 (O_1381,N_14862,N_14990);
nand UO_1382 (O_1382,N_14901,N_14954);
nor UO_1383 (O_1383,N_14972,N_14963);
nand UO_1384 (O_1384,N_14851,N_14918);
nand UO_1385 (O_1385,N_14948,N_14873);
nand UO_1386 (O_1386,N_14872,N_14991);
xor UO_1387 (O_1387,N_14934,N_14867);
nand UO_1388 (O_1388,N_14997,N_14942);
nand UO_1389 (O_1389,N_14863,N_14922);
nor UO_1390 (O_1390,N_14871,N_14922);
xor UO_1391 (O_1391,N_14955,N_14863);
or UO_1392 (O_1392,N_14916,N_14858);
or UO_1393 (O_1393,N_14927,N_14894);
or UO_1394 (O_1394,N_14969,N_14933);
nor UO_1395 (O_1395,N_14961,N_14914);
xor UO_1396 (O_1396,N_14921,N_14890);
nor UO_1397 (O_1397,N_14877,N_14958);
and UO_1398 (O_1398,N_14855,N_14970);
xor UO_1399 (O_1399,N_14942,N_14986);
or UO_1400 (O_1400,N_14996,N_14983);
nand UO_1401 (O_1401,N_14899,N_14986);
nand UO_1402 (O_1402,N_14991,N_14985);
and UO_1403 (O_1403,N_14882,N_14876);
nand UO_1404 (O_1404,N_14932,N_14861);
nor UO_1405 (O_1405,N_14967,N_14883);
xor UO_1406 (O_1406,N_14947,N_14969);
xor UO_1407 (O_1407,N_14886,N_14950);
nand UO_1408 (O_1408,N_14862,N_14874);
xor UO_1409 (O_1409,N_14861,N_14925);
nand UO_1410 (O_1410,N_14895,N_14863);
nand UO_1411 (O_1411,N_14926,N_14884);
xnor UO_1412 (O_1412,N_14889,N_14890);
xor UO_1413 (O_1413,N_14963,N_14886);
and UO_1414 (O_1414,N_14921,N_14906);
and UO_1415 (O_1415,N_14961,N_14881);
and UO_1416 (O_1416,N_14981,N_14915);
nand UO_1417 (O_1417,N_14955,N_14970);
and UO_1418 (O_1418,N_14880,N_14892);
nor UO_1419 (O_1419,N_14996,N_14878);
nand UO_1420 (O_1420,N_14938,N_14884);
xnor UO_1421 (O_1421,N_14908,N_14900);
nand UO_1422 (O_1422,N_14886,N_14938);
nand UO_1423 (O_1423,N_14875,N_14917);
xnor UO_1424 (O_1424,N_14994,N_14962);
xor UO_1425 (O_1425,N_14996,N_14985);
and UO_1426 (O_1426,N_14972,N_14893);
xor UO_1427 (O_1427,N_14986,N_14895);
xnor UO_1428 (O_1428,N_14888,N_14983);
nand UO_1429 (O_1429,N_14957,N_14948);
and UO_1430 (O_1430,N_14876,N_14871);
nor UO_1431 (O_1431,N_14910,N_14893);
or UO_1432 (O_1432,N_14969,N_14882);
nor UO_1433 (O_1433,N_14949,N_14990);
nand UO_1434 (O_1434,N_14985,N_14958);
nor UO_1435 (O_1435,N_14987,N_14975);
nor UO_1436 (O_1436,N_14996,N_14861);
or UO_1437 (O_1437,N_14978,N_14934);
xnor UO_1438 (O_1438,N_14909,N_14986);
and UO_1439 (O_1439,N_14963,N_14985);
and UO_1440 (O_1440,N_14910,N_14918);
nor UO_1441 (O_1441,N_14966,N_14930);
and UO_1442 (O_1442,N_14872,N_14874);
nand UO_1443 (O_1443,N_14882,N_14922);
or UO_1444 (O_1444,N_14853,N_14858);
and UO_1445 (O_1445,N_14960,N_14927);
nand UO_1446 (O_1446,N_14944,N_14885);
or UO_1447 (O_1447,N_14974,N_14874);
nor UO_1448 (O_1448,N_14889,N_14869);
and UO_1449 (O_1449,N_14888,N_14982);
xnor UO_1450 (O_1450,N_14913,N_14872);
xnor UO_1451 (O_1451,N_14974,N_14957);
nand UO_1452 (O_1452,N_14875,N_14859);
xnor UO_1453 (O_1453,N_14967,N_14912);
and UO_1454 (O_1454,N_14911,N_14984);
nand UO_1455 (O_1455,N_14854,N_14914);
nor UO_1456 (O_1456,N_14977,N_14978);
nand UO_1457 (O_1457,N_14933,N_14875);
xor UO_1458 (O_1458,N_14937,N_14994);
and UO_1459 (O_1459,N_14941,N_14865);
xor UO_1460 (O_1460,N_14950,N_14961);
and UO_1461 (O_1461,N_14924,N_14884);
and UO_1462 (O_1462,N_14926,N_14881);
nand UO_1463 (O_1463,N_14962,N_14876);
or UO_1464 (O_1464,N_14884,N_14880);
xor UO_1465 (O_1465,N_14877,N_14939);
or UO_1466 (O_1466,N_14857,N_14872);
and UO_1467 (O_1467,N_14923,N_14856);
or UO_1468 (O_1468,N_14938,N_14876);
xor UO_1469 (O_1469,N_14990,N_14963);
nor UO_1470 (O_1470,N_14865,N_14945);
xor UO_1471 (O_1471,N_14887,N_14888);
nand UO_1472 (O_1472,N_14895,N_14890);
or UO_1473 (O_1473,N_14974,N_14910);
nand UO_1474 (O_1474,N_14946,N_14850);
and UO_1475 (O_1475,N_14929,N_14858);
xnor UO_1476 (O_1476,N_14857,N_14882);
and UO_1477 (O_1477,N_14911,N_14965);
nand UO_1478 (O_1478,N_14857,N_14864);
xor UO_1479 (O_1479,N_14955,N_14887);
xor UO_1480 (O_1480,N_14911,N_14875);
nand UO_1481 (O_1481,N_14879,N_14889);
nor UO_1482 (O_1482,N_14930,N_14978);
and UO_1483 (O_1483,N_14937,N_14931);
nor UO_1484 (O_1484,N_14872,N_14976);
or UO_1485 (O_1485,N_14936,N_14897);
nor UO_1486 (O_1486,N_14870,N_14900);
or UO_1487 (O_1487,N_14861,N_14895);
and UO_1488 (O_1488,N_14885,N_14896);
nor UO_1489 (O_1489,N_14902,N_14984);
or UO_1490 (O_1490,N_14853,N_14999);
or UO_1491 (O_1491,N_14905,N_14998);
and UO_1492 (O_1492,N_14913,N_14906);
nor UO_1493 (O_1493,N_14940,N_14938);
xnor UO_1494 (O_1494,N_14885,N_14889);
or UO_1495 (O_1495,N_14898,N_14851);
or UO_1496 (O_1496,N_14883,N_14990);
xnor UO_1497 (O_1497,N_14866,N_14940);
xnor UO_1498 (O_1498,N_14969,N_14986);
and UO_1499 (O_1499,N_14933,N_14879);
nand UO_1500 (O_1500,N_14886,N_14879);
xnor UO_1501 (O_1501,N_14966,N_14903);
xor UO_1502 (O_1502,N_14868,N_14876);
xnor UO_1503 (O_1503,N_14994,N_14906);
nor UO_1504 (O_1504,N_14895,N_14946);
nand UO_1505 (O_1505,N_14983,N_14986);
nor UO_1506 (O_1506,N_14902,N_14945);
or UO_1507 (O_1507,N_14965,N_14892);
nor UO_1508 (O_1508,N_14886,N_14936);
or UO_1509 (O_1509,N_14982,N_14917);
xnor UO_1510 (O_1510,N_14962,N_14985);
xor UO_1511 (O_1511,N_14878,N_14997);
or UO_1512 (O_1512,N_14906,N_14869);
nor UO_1513 (O_1513,N_14896,N_14979);
xor UO_1514 (O_1514,N_14885,N_14983);
and UO_1515 (O_1515,N_14971,N_14996);
nand UO_1516 (O_1516,N_14950,N_14923);
or UO_1517 (O_1517,N_14988,N_14952);
nor UO_1518 (O_1518,N_14908,N_14959);
nor UO_1519 (O_1519,N_14879,N_14957);
nand UO_1520 (O_1520,N_14975,N_14893);
and UO_1521 (O_1521,N_14873,N_14960);
nand UO_1522 (O_1522,N_14944,N_14957);
nand UO_1523 (O_1523,N_14972,N_14902);
nand UO_1524 (O_1524,N_14953,N_14961);
or UO_1525 (O_1525,N_14863,N_14924);
nand UO_1526 (O_1526,N_14890,N_14893);
and UO_1527 (O_1527,N_14947,N_14866);
xor UO_1528 (O_1528,N_14857,N_14924);
nor UO_1529 (O_1529,N_14861,N_14878);
nand UO_1530 (O_1530,N_14920,N_14900);
nor UO_1531 (O_1531,N_14937,N_14981);
and UO_1532 (O_1532,N_14850,N_14887);
or UO_1533 (O_1533,N_14864,N_14926);
and UO_1534 (O_1534,N_14940,N_14985);
nor UO_1535 (O_1535,N_14926,N_14939);
xor UO_1536 (O_1536,N_14889,N_14972);
or UO_1537 (O_1537,N_14863,N_14979);
nand UO_1538 (O_1538,N_14984,N_14983);
or UO_1539 (O_1539,N_14968,N_14991);
or UO_1540 (O_1540,N_14866,N_14905);
xor UO_1541 (O_1541,N_14935,N_14932);
or UO_1542 (O_1542,N_14890,N_14993);
and UO_1543 (O_1543,N_14912,N_14908);
and UO_1544 (O_1544,N_14950,N_14983);
or UO_1545 (O_1545,N_14913,N_14882);
xnor UO_1546 (O_1546,N_14996,N_14998);
nand UO_1547 (O_1547,N_14917,N_14943);
xnor UO_1548 (O_1548,N_14971,N_14904);
nand UO_1549 (O_1549,N_14879,N_14921);
xnor UO_1550 (O_1550,N_14869,N_14874);
nand UO_1551 (O_1551,N_14993,N_14865);
nand UO_1552 (O_1552,N_14991,N_14912);
nand UO_1553 (O_1553,N_14869,N_14985);
and UO_1554 (O_1554,N_14871,N_14886);
or UO_1555 (O_1555,N_14906,N_14959);
and UO_1556 (O_1556,N_14942,N_14853);
or UO_1557 (O_1557,N_14962,N_14893);
xor UO_1558 (O_1558,N_14895,N_14959);
or UO_1559 (O_1559,N_14889,N_14908);
nand UO_1560 (O_1560,N_14925,N_14889);
nor UO_1561 (O_1561,N_14983,N_14960);
or UO_1562 (O_1562,N_14896,N_14856);
nand UO_1563 (O_1563,N_14879,N_14961);
nor UO_1564 (O_1564,N_14973,N_14969);
xor UO_1565 (O_1565,N_14943,N_14968);
nand UO_1566 (O_1566,N_14943,N_14983);
and UO_1567 (O_1567,N_14928,N_14851);
nand UO_1568 (O_1568,N_14866,N_14956);
and UO_1569 (O_1569,N_14970,N_14938);
nand UO_1570 (O_1570,N_14855,N_14989);
nand UO_1571 (O_1571,N_14942,N_14980);
or UO_1572 (O_1572,N_14969,N_14982);
xnor UO_1573 (O_1573,N_14888,N_14963);
or UO_1574 (O_1574,N_14989,N_14965);
and UO_1575 (O_1575,N_14859,N_14933);
nor UO_1576 (O_1576,N_14969,N_14924);
and UO_1577 (O_1577,N_14927,N_14957);
or UO_1578 (O_1578,N_14901,N_14885);
xnor UO_1579 (O_1579,N_14983,N_14992);
nand UO_1580 (O_1580,N_14981,N_14978);
and UO_1581 (O_1581,N_14857,N_14896);
or UO_1582 (O_1582,N_14974,N_14857);
nor UO_1583 (O_1583,N_14866,N_14933);
and UO_1584 (O_1584,N_14960,N_14895);
nor UO_1585 (O_1585,N_14898,N_14862);
or UO_1586 (O_1586,N_14989,N_14948);
or UO_1587 (O_1587,N_14904,N_14969);
and UO_1588 (O_1588,N_14939,N_14911);
nand UO_1589 (O_1589,N_14851,N_14872);
xnor UO_1590 (O_1590,N_14993,N_14876);
nor UO_1591 (O_1591,N_14884,N_14956);
and UO_1592 (O_1592,N_14925,N_14943);
xor UO_1593 (O_1593,N_14951,N_14852);
or UO_1594 (O_1594,N_14971,N_14912);
xnor UO_1595 (O_1595,N_14910,N_14965);
nor UO_1596 (O_1596,N_14924,N_14996);
nor UO_1597 (O_1597,N_14890,N_14938);
or UO_1598 (O_1598,N_14868,N_14977);
and UO_1599 (O_1599,N_14980,N_14937);
nand UO_1600 (O_1600,N_14893,N_14896);
nand UO_1601 (O_1601,N_14918,N_14901);
nor UO_1602 (O_1602,N_14908,N_14960);
xor UO_1603 (O_1603,N_14944,N_14910);
or UO_1604 (O_1604,N_14933,N_14967);
nand UO_1605 (O_1605,N_14878,N_14877);
nor UO_1606 (O_1606,N_14993,N_14968);
nor UO_1607 (O_1607,N_14976,N_14876);
or UO_1608 (O_1608,N_14925,N_14948);
nand UO_1609 (O_1609,N_14953,N_14899);
or UO_1610 (O_1610,N_14885,N_14882);
nand UO_1611 (O_1611,N_14883,N_14935);
or UO_1612 (O_1612,N_14927,N_14985);
and UO_1613 (O_1613,N_14921,N_14962);
xor UO_1614 (O_1614,N_14860,N_14941);
and UO_1615 (O_1615,N_14956,N_14987);
nand UO_1616 (O_1616,N_14894,N_14922);
and UO_1617 (O_1617,N_14967,N_14969);
xnor UO_1618 (O_1618,N_14908,N_14980);
nand UO_1619 (O_1619,N_14937,N_14885);
and UO_1620 (O_1620,N_14957,N_14889);
nand UO_1621 (O_1621,N_14906,N_14978);
or UO_1622 (O_1622,N_14986,N_14890);
or UO_1623 (O_1623,N_14857,N_14983);
nor UO_1624 (O_1624,N_14900,N_14887);
nand UO_1625 (O_1625,N_14896,N_14926);
and UO_1626 (O_1626,N_14917,N_14997);
xnor UO_1627 (O_1627,N_14999,N_14897);
xnor UO_1628 (O_1628,N_14954,N_14853);
xnor UO_1629 (O_1629,N_14960,N_14920);
nor UO_1630 (O_1630,N_14872,N_14986);
xnor UO_1631 (O_1631,N_14866,N_14959);
xor UO_1632 (O_1632,N_14880,N_14999);
or UO_1633 (O_1633,N_14871,N_14902);
nor UO_1634 (O_1634,N_14880,N_14863);
and UO_1635 (O_1635,N_14960,N_14987);
xor UO_1636 (O_1636,N_14934,N_14992);
nor UO_1637 (O_1637,N_14850,N_14962);
xnor UO_1638 (O_1638,N_14933,N_14951);
or UO_1639 (O_1639,N_14899,N_14877);
nor UO_1640 (O_1640,N_14902,N_14890);
xor UO_1641 (O_1641,N_14963,N_14876);
xor UO_1642 (O_1642,N_14911,N_14885);
and UO_1643 (O_1643,N_14988,N_14878);
and UO_1644 (O_1644,N_14999,N_14923);
and UO_1645 (O_1645,N_14995,N_14977);
or UO_1646 (O_1646,N_14885,N_14914);
nor UO_1647 (O_1647,N_14991,N_14972);
nand UO_1648 (O_1648,N_14896,N_14919);
nand UO_1649 (O_1649,N_14977,N_14961);
nand UO_1650 (O_1650,N_14940,N_14871);
xor UO_1651 (O_1651,N_14992,N_14956);
nor UO_1652 (O_1652,N_14867,N_14903);
and UO_1653 (O_1653,N_14916,N_14996);
xnor UO_1654 (O_1654,N_14891,N_14993);
xor UO_1655 (O_1655,N_14991,N_14919);
and UO_1656 (O_1656,N_14936,N_14990);
xor UO_1657 (O_1657,N_14915,N_14904);
xnor UO_1658 (O_1658,N_14986,N_14958);
nand UO_1659 (O_1659,N_14890,N_14988);
xnor UO_1660 (O_1660,N_14969,N_14958);
nand UO_1661 (O_1661,N_14896,N_14905);
and UO_1662 (O_1662,N_14873,N_14930);
and UO_1663 (O_1663,N_14931,N_14904);
nor UO_1664 (O_1664,N_14953,N_14878);
nand UO_1665 (O_1665,N_14865,N_14911);
nand UO_1666 (O_1666,N_14901,N_14920);
or UO_1667 (O_1667,N_14996,N_14865);
xor UO_1668 (O_1668,N_14956,N_14913);
nor UO_1669 (O_1669,N_14939,N_14855);
nand UO_1670 (O_1670,N_14983,N_14962);
nand UO_1671 (O_1671,N_14985,N_14890);
nand UO_1672 (O_1672,N_14989,N_14984);
nor UO_1673 (O_1673,N_14902,N_14994);
xnor UO_1674 (O_1674,N_14957,N_14955);
or UO_1675 (O_1675,N_14970,N_14978);
or UO_1676 (O_1676,N_14998,N_14856);
nand UO_1677 (O_1677,N_14944,N_14954);
nand UO_1678 (O_1678,N_14916,N_14934);
or UO_1679 (O_1679,N_14930,N_14868);
nor UO_1680 (O_1680,N_14955,N_14922);
xnor UO_1681 (O_1681,N_14964,N_14923);
xor UO_1682 (O_1682,N_14928,N_14857);
xor UO_1683 (O_1683,N_14873,N_14868);
and UO_1684 (O_1684,N_14988,N_14986);
and UO_1685 (O_1685,N_14862,N_14883);
nor UO_1686 (O_1686,N_14935,N_14897);
and UO_1687 (O_1687,N_14971,N_14851);
nand UO_1688 (O_1688,N_14992,N_14881);
nor UO_1689 (O_1689,N_14905,N_14915);
or UO_1690 (O_1690,N_14905,N_14994);
and UO_1691 (O_1691,N_14973,N_14877);
and UO_1692 (O_1692,N_14904,N_14954);
or UO_1693 (O_1693,N_14940,N_14945);
nor UO_1694 (O_1694,N_14944,N_14856);
nor UO_1695 (O_1695,N_14972,N_14906);
nand UO_1696 (O_1696,N_14968,N_14897);
nor UO_1697 (O_1697,N_14906,N_14998);
nor UO_1698 (O_1698,N_14928,N_14989);
nor UO_1699 (O_1699,N_14878,N_14855);
and UO_1700 (O_1700,N_14865,N_14904);
xor UO_1701 (O_1701,N_14932,N_14907);
nand UO_1702 (O_1702,N_14867,N_14988);
xnor UO_1703 (O_1703,N_14906,N_14924);
xnor UO_1704 (O_1704,N_14946,N_14872);
or UO_1705 (O_1705,N_14871,N_14934);
nor UO_1706 (O_1706,N_14962,N_14955);
xor UO_1707 (O_1707,N_14867,N_14978);
nor UO_1708 (O_1708,N_14907,N_14852);
xor UO_1709 (O_1709,N_14979,N_14855);
nand UO_1710 (O_1710,N_14920,N_14868);
or UO_1711 (O_1711,N_14975,N_14856);
xor UO_1712 (O_1712,N_14855,N_14951);
or UO_1713 (O_1713,N_14917,N_14850);
or UO_1714 (O_1714,N_14949,N_14869);
nand UO_1715 (O_1715,N_14960,N_14993);
xnor UO_1716 (O_1716,N_14853,N_14963);
nand UO_1717 (O_1717,N_14862,N_14863);
and UO_1718 (O_1718,N_14946,N_14865);
and UO_1719 (O_1719,N_14998,N_14913);
nor UO_1720 (O_1720,N_14871,N_14850);
or UO_1721 (O_1721,N_14904,N_14930);
or UO_1722 (O_1722,N_14988,N_14858);
xor UO_1723 (O_1723,N_14890,N_14936);
or UO_1724 (O_1724,N_14946,N_14965);
nor UO_1725 (O_1725,N_14859,N_14938);
nand UO_1726 (O_1726,N_14919,N_14952);
nor UO_1727 (O_1727,N_14932,N_14960);
or UO_1728 (O_1728,N_14859,N_14884);
xnor UO_1729 (O_1729,N_14921,N_14870);
and UO_1730 (O_1730,N_14936,N_14911);
nand UO_1731 (O_1731,N_14978,N_14879);
nor UO_1732 (O_1732,N_14894,N_14871);
nor UO_1733 (O_1733,N_14912,N_14988);
or UO_1734 (O_1734,N_14993,N_14953);
xnor UO_1735 (O_1735,N_14921,N_14913);
xor UO_1736 (O_1736,N_14935,N_14968);
xor UO_1737 (O_1737,N_14984,N_14965);
nand UO_1738 (O_1738,N_14871,N_14907);
or UO_1739 (O_1739,N_14986,N_14931);
nand UO_1740 (O_1740,N_14980,N_14912);
and UO_1741 (O_1741,N_14879,N_14980);
or UO_1742 (O_1742,N_14970,N_14941);
or UO_1743 (O_1743,N_14874,N_14878);
nand UO_1744 (O_1744,N_14932,N_14909);
or UO_1745 (O_1745,N_14962,N_14922);
or UO_1746 (O_1746,N_14876,N_14923);
and UO_1747 (O_1747,N_14933,N_14873);
xnor UO_1748 (O_1748,N_14902,N_14954);
xnor UO_1749 (O_1749,N_14999,N_14871);
or UO_1750 (O_1750,N_14987,N_14899);
and UO_1751 (O_1751,N_14947,N_14949);
nor UO_1752 (O_1752,N_14921,N_14969);
nand UO_1753 (O_1753,N_14910,N_14850);
nor UO_1754 (O_1754,N_14888,N_14972);
xnor UO_1755 (O_1755,N_14972,N_14981);
nor UO_1756 (O_1756,N_14984,N_14879);
or UO_1757 (O_1757,N_14922,N_14985);
and UO_1758 (O_1758,N_14954,N_14900);
xor UO_1759 (O_1759,N_14945,N_14857);
and UO_1760 (O_1760,N_14970,N_14869);
or UO_1761 (O_1761,N_14992,N_14955);
xnor UO_1762 (O_1762,N_14921,N_14871);
and UO_1763 (O_1763,N_14958,N_14990);
nor UO_1764 (O_1764,N_14890,N_14948);
nand UO_1765 (O_1765,N_14987,N_14942);
or UO_1766 (O_1766,N_14903,N_14865);
and UO_1767 (O_1767,N_14993,N_14937);
nand UO_1768 (O_1768,N_14961,N_14968);
xnor UO_1769 (O_1769,N_14887,N_14965);
or UO_1770 (O_1770,N_14902,N_14952);
xnor UO_1771 (O_1771,N_14922,N_14941);
nand UO_1772 (O_1772,N_14865,N_14989);
nor UO_1773 (O_1773,N_14937,N_14909);
or UO_1774 (O_1774,N_14920,N_14914);
or UO_1775 (O_1775,N_14970,N_14911);
or UO_1776 (O_1776,N_14998,N_14863);
or UO_1777 (O_1777,N_14861,N_14876);
nor UO_1778 (O_1778,N_14974,N_14877);
nand UO_1779 (O_1779,N_14884,N_14866);
nor UO_1780 (O_1780,N_14866,N_14971);
nand UO_1781 (O_1781,N_14907,N_14885);
nand UO_1782 (O_1782,N_14920,N_14906);
and UO_1783 (O_1783,N_14854,N_14915);
xor UO_1784 (O_1784,N_14992,N_14920);
and UO_1785 (O_1785,N_14979,N_14960);
and UO_1786 (O_1786,N_14916,N_14954);
nor UO_1787 (O_1787,N_14925,N_14918);
nor UO_1788 (O_1788,N_14959,N_14937);
or UO_1789 (O_1789,N_14928,N_14993);
nor UO_1790 (O_1790,N_14944,N_14870);
and UO_1791 (O_1791,N_14894,N_14921);
and UO_1792 (O_1792,N_14968,N_14989);
or UO_1793 (O_1793,N_14861,N_14881);
xor UO_1794 (O_1794,N_14884,N_14940);
nand UO_1795 (O_1795,N_14865,N_14982);
nand UO_1796 (O_1796,N_14996,N_14936);
and UO_1797 (O_1797,N_14870,N_14962);
nor UO_1798 (O_1798,N_14963,N_14890);
nor UO_1799 (O_1799,N_14969,N_14883);
xnor UO_1800 (O_1800,N_14996,N_14873);
xnor UO_1801 (O_1801,N_14959,N_14852);
xnor UO_1802 (O_1802,N_14887,N_14922);
and UO_1803 (O_1803,N_14992,N_14916);
and UO_1804 (O_1804,N_14973,N_14947);
or UO_1805 (O_1805,N_14855,N_14905);
nor UO_1806 (O_1806,N_14851,N_14861);
and UO_1807 (O_1807,N_14952,N_14891);
xnor UO_1808 (O_1808,N_14920,N_14976);
nor UO_1809 (O_1809,N_14964,N_14987);
nand UO_1810 (O_1810,N_14883,N_14869);
and UO_1811 (O_1811,N_14997,N_14955);
nor UO_1812 (O_1812,N_14871,N_14865);
nand UO_1813 (O_1813,N_14938,N_14909);
xnor UO_1814 (O_1814,N_14877,N_14965);
nor UO_1815 (O_1815,N_14980,N_14953);
nand UO_1816 (O_1816,N_14960,N_14931);
xnor UO_1817 (O_1817,N_14903,N_14873);
nand UO_1818 (O_1818,N_14877,N_14850);
and UO_1819 (O_1819,N_14929,N_14973);
and UO_1820 (O_1820,N_14919,N_14929);
and UO_1821 (O_1821,N_14858,N_14997);
nor UO_1822 (O_1822,N_14963,N_14919);
and UO_1823 (O_1823,N_14963,N_14953);
nand UO_1824 (O_1824,N_14911,N_14887);
xor UO_1825 (O_1825,N_14924,N_14959);
nor UO_1826 (O_1826,N_14907,N_14870);
and UO_1827 (O_1827,N_14931,N_14884);
or UO_1828 (O_1828,N_14958,N_14905);
nor UO_1829 (O_1829,N_14869,N_14975);
or UO_1830 (O_1830,N_14983,N_14862);
xor UO_1831 (O_1831,N_14891,N_14981);
nor UO_1832 (O_1832,N_14854,N_14952);
nand UO_1833 (O_1833,N_14952,N_14977);
and UO_1834 (O_1834,N_14973,N_14873);
nor UO_1835 (O_1835,N_14998,N_14940);
and UO_1836 (O_1836,N_14980,N_14977);
xnor UO_1837 (O_1837,N_14940,N_14975);
nand UO_1838 (O_1838,N_14948,N_14898);
nor UO_1839 (O_1839,N_14908,N_14969);
or UO_1840 (O_1840,N_14990,N_14940);
or UO_1841 (O_1841,N_14965,N_14990);
nor UO_1842 (O_1842,N_14914,N_14946);
or UO_1843 (O_1843,N_14943,N_14958);
and UO_1844 (O_1844,N_14949,N_14865);
nor UO_1845 (O_1845,N_14854,N_14930);
xnor UO_1846 (O_1846,N_14897,N_14938);
xnor UO_1847 (O_1847,N_14882,N_14960);
nand UO_1848 (O_1848,N_14919,N_14947);
or UO_1849 (O_1849,N_14975,N_14966);
or UO_1850 (O_1850,N_14903,N_14959);
nor UO_1851 (O_1851,N_14961,N_14934);
and UO_1852 (O_1852,N_14987,N_14947);
and UO_1853 (O_1853,N_14944,N_14977);
nor UO_1854 (O_1854,N_14992,N_14965);
or UO_1855 (O_1855,N_14873,N_14944);
nand UO_1856 (O_1856,N_14881,N_14938);
nand UO_1857 (O_1857,N_14918,N_14957);
or UO_1858 (O_1858,N_14915,N_14936);
nor UO_1859 (O_1859,N_14934,N_14899);
and UO_1860 (O_1860,N_14906,N_14885);
xor UO_1861 (O_1861,N_14918,N_14914);
and UO_1862 (O_1862,N_14927,N_14892);
or UO_1863 (O_1863,N_14900,N_14940);
nor UO_1864 (O_1864,N_14920,N_14881);
xnor UO_1865 (O_1865,N_14970,N_14879);
xor UO_1866 (O_1866,N_14931,N_14965);
nand UO_1867 (O_1867,N_14975,N_14927);
nor UO_1868 (O_1868,N_14929,N_14908);
xor UO_1869 (O_1869,N_14999,N_14919);
and UO_1870 (O_1870,N_14949,N_14936);
nand UO_1871 (O_1871,N_14924,N_14974);
nand UO_1872 (O_1872,N_14865,N_14957);
and UO_1873 (O_1873,N_14924,N_14985);
and UO_1874 (O_1874,N_14997,N_14949);
nor UO_1875 (O_1875,N_14987,N_14926);
xor UO_1876 (O_1876,N_14856,N_14889);
or UO_1877 (O_1877,N_14892,N_14967);
and UO_1878 (O_1878,N_14897,N_14867);
or UO_1879 (O_1879,N_14857,N_14871);
nor UO_1880 (O_1880,N_14959,N_14997);
nor UO_1881 (O_1881,N_14998,N_14954);
nor UO_1882 (O_1882,N_14916,N_14932);
nand UO_1883 (O_1883,N_14995,N_14913);
nand UO_1884 (O_1884,N_14978,N_14887);
nor UO_1885 (O_1885,N_14972,N_14907);
or UO_1886 (O_1886,N_14925,N_14873);
nand UO_1887 (O_1887,N_14977,N_14884);
or UO_1888 (O_1888,N_14927,N_14996);
xnor UO_1889 (O_1889,N_14928,N_14855);
xor UO_1890 (O_1890,N_14892,N_14926);
or UO_1891 (O_1891,N_14852,N_14969);
nor UO_1892 (O_1892,N_14868,N_14867);
xnor UO_1893 (O_1893,N_14867,N_14872);
or UO_1894 (O_1894,N_14915,N_14860);
nand UO_1895 (O_1895,N_14877,N_14858);
xor UO_1896 (O_1896,N_14918,N_14961);
nand UO_1897 (O_1897,N_14873,N_14970);
or UO_1898 (O_1898,N_14864,N_14912);
nor UO_1899 (O_1899,N_14858,N_14950);
nand UO_1900 (O_1900,N_14905,N_14966);
and UO_1901 (O_1901,N_14972,N_14951);
nand UO_1902 (O_1902,N_14894,N_14880);
or UO_1903 (O_1903,N_14901,N_14987);
xor UO_1904 (O_1904,N_14946,N_14993);
nor UO_1905 (O_1905,N_14921,N_14919);
nor UO_1906 (O_1906,N_14895,N_14966);
and UO_1907 (O_1907,N_14961,N_14975);
nand UO_1908 (O_1908,N_14992,N_14921);
or UO_1909 (O_1909,N_14871,N_14992);
or UO_1910 (O_1910,N_14875,N_14894);
nor UO_1911 (O_1911,N_14974,N_14894);
xor UO_1912 (O_1912,N_14905,N_14884);
nand UO_1913 (O_1913,N_14879,N_14965);
xor UO_1914 (O_1914,N_14975,N_14958);
nand UO_1915 (O_1915,N_14965,N_14952);
xor UO_1916 (O_1916,N_14938,N_14960);
nand UO_1917 (O_1917,N_14861,N_14967);
or UO_1918 (O_1918,N_14867,N_14944);
nor UO_1919 (O_1919,N_14915,N_14948);
xor UO_1920 (O_1920,N_14858,N_14958);
nand UO_1921 (O_1921,N_14993,N_14954);
nand UO_1922 (O_1922,N_14991,N_14987);
or UO_1923 (O_1923,N_14886,N_14946);
nand UO_1924 (O_1924,N_14912,N_14916);
xor UO_1925 (O_1925,N_14984,N_14862);
or UO_1926 (O_1926,N_14882,N_14881);
nor UO_1927 (O_1927,N_14960,N_14899);
nand UO_1928 (O_1928,N_14852,N_14985);
nor UO_1929 (O_1929,N_14913,N_14894);
xnor UO_1930 (O_1930,N_14939,N_14912);
nor UO_1931 (O_1931,N_14909,N_14962);
nand UO_1932 (O_1932,N_14903,N_14872);
nand UO_1933 (O_1933,N_14943,N_14980);
xnor UO_1934 (O_1934,N_14951,N_14958);
or UO_1935 (O_1935,N_14938,N_14863);
xnor UO_1936 (O_1936,N_14966,N_14915);
and UO_1937 (O_1937,N_14851,N_14948);
nand UO_1938 (O_1938,N_14991,N_14862);
or UO_1939 (O_1939,N_14949,N_14952);
nor UO_1940 (O_1940,N_14899,N_14868);
nor UO_1941 (O_1941,N_14923,N_14940);
or UO_1942 (O_1942,N_14930,N_14869);
nand UO_1943 (O_1943,N_14916,N_14904);
or UO_1944 (O_1944,N_14937,N_14930);
nor UO_1945 (O_1945,N_14940,N_14969);
nand UO_1946 (O_1946,N_14970,N_14956);
nor UO_1947 (O_1947,N_14913,N_14854);
xor UO_1948 (O_1948,N_14876,N_14862);
and UO_1949 (O_1949,N_14966,N_14936);
xor UO_1950 (O_1950,N_14866,N_14909);
and UO_1951 (O_1951,N_14931,N_14972);
xor UO_1952 (O_1952,N_14945,N_14921);
and UO_1953 (O_1953,N_14854,N_14901);
or UO_1954 (O_1954,N_14982,N_14942);
or UO_1955 (O_1955,N_14941,N_14890);
nand UO_1956 (O_1956,N_14921,N_14940);
xnor UO_1957 (O_1957,N_14943,N_14997);
and UO_1958 (O_1958,N_14888,N_14934);
and UO_1959 (O_1959,N_14954,N_14864);
or UO_1960 (O_1960,N_14935,N_14926);
and UO_1961 (O_1961,N_14940,N_14869);
nor UO_1962 (O_1962,N_14939,N_14958);
and UO_1963 (O_1963,N_14879,N_14871);
and UO_1964 (O_1964,N_14927,N_14955);
nand UO_1965 (O_1965,N_14991,N_14950);
nand UO_1966 (O_1966,N_14923,N_14981);
nor UO_1967 (O_1967,N_14944,N_14953);
or UO_1968 (O_1968,N_14924,N_14987);
and UO_1969 (O_1969,N_14956,N_14986);
nor UO_1970 (O_1970,N_14886,N_14976);
xor UO_1971 (O_1971,N_14968,N_14941);
or UO_1972 (O_1972,N_14860,N_14954);
and UO_1973 (O_1973,N_14948,N_14941);
nand UO_1974 (O_1974,N_14889,N_14971);
or UO_1975 (O_1975,N_14951,N_14962);
or UO_1976 (O_1976,N_14993,N_14986);
and UO_1977 (O_1977,N_14859,N_14896);
nand UO_1978 (O_1978,N_14872,N_14993);
xnor UO_1979 (O_1979,N_14904,N_14963);
xor UO_1980 (O_1980,N_14907,N_14851);
or UO_1981 (O_1981,N_14871,N_14895);
and UO_1982 (O_1982,N_14952,N_14951);
xor UO_1983 (O_1983,N_14926,N_14857);
nand UO_1984 (O_1984,N_14971,N_14948);
nor UO_1985 (O_1985,N_14888,N_14980);
xor UO_1986 (O_1986,N_14863,N_14853);
xnor UO_1987 (O_1987,N_14892,N_14853);
nor UO_1988 (O_1988,N_14850,N_14963);
nor UO_1989 (O_1989,N_14951,N_14997);
xor UO_1990 (O_1990,N_14899,N_14990);
and UO_1991 (O_1991,N_14856,N_14983);
nand UO_1992 (O_1992,N_14984,N_14974);
and UO_1993 (O_1993,N_14876,N_14915);
nor UO_1994 (O_1994,N_14952,N_14964);
or UO_1995 (O_1995,N_14925,N_14997);
or UO_1996 (O_1996,N_14863,N_14982);
nand UO_1997 (O_1997,N_14955,N_14986);
or UO_1998 (O_1998,N_14960,N_14887);
and UO_1999 (O_1999,N_14948,N_14877);
endmodule