module basic_500_3000_500_4_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_341,In_487);
nor U1 (N_1,In_85,In_127);
nand U2 (N_2,In_27,In_351);
xor U3 (N_3,In_405,In_419);
nand U4 (N_4,In_11,In_315);
and U5 (N_5,In_91,In_339);
nor U6 (N_6,In_79,In_34);
or U7 (N_7,In_276,In_16);
nand U8 (N_8,In_454,In_61);
nand U9 (N_9,In_427,In_362);
and U10 (N_10,In_322,In_397);
or U11 (N_11,In_131,In_86);
xor U12 (N_12,In_496,In_159);
and U13 (N_13,In_44,In_388);
nor U14 (N_14,In_208,In_437);
nand U15 (N_15,In_122,In_120);
xnor U16 (N_16,In_169,In_289);
nand U17 (N_17,In_170,In_286);
and U18 (N_18,In_469,In_287);
and U19 (N_19,In_9,In_353);
nor U20 (N_20,In_373,In_497);
nor U21 (N_21,In_365,In_30);
nand U22 (N_22,In_165,In_369);
and U23 (N_23,In_87,In_47);
or U24 (N_24,In_393,In_150);
and U25 (N_25,In_266,In_359);
and U26 (N_26,In_107,In_100);
and U27 (N_27,In_300,In_338);
or U28 (N_28,In_46,In_104);
nor U29 (N_29,In_391,In_110);
nor U30 (N_30,In_492,In_458);
and U31 (N_31,In_31,In_255);
nor U32 (N_32,In_400,In_188);
nand U33 (N_33,In_187,In_68);
and U34 (N_34,In_383,In_275);
or U35 (N_35,In_453,In_385);
nand U36 (N_36,In_380,In_396);
or U37 (N_37,In_55,In_433);
and U38 (N_38,In_387,In_270);
nor U39 (N_39,In_456,In_228);
xnor U40 (N_40,In_0,In_316);
nand U41 (N_41,In_312,In_439);
nand U42 (N_42,In_407,In_220);
and U43 (N_43,In_319,In_221);
and U44 (N_44,In_342,In_448);
or U45 (N_45,In_303,In_25);
and U46 (N_46,In_211,In_232);
or U47 (N_47,In_471,In_384);
nor U48 (N_48,In_477,In_89);
and U49 (N_49,In_49,In_82);
nand U50 (N_50,In_146,In_263);
nand U51 (N_51,In_259,In_140);
and U52 (N_52,In_54,In_467);
nor U53 (N_53,In_329,In_426);
xnor U54 (N_54,In_214,In_474);
nand U55 (N_55,In_75,In_52);
or U56 (N_56,In_318,In_445);
or U57 (N_57,In_483,In_175);
and U58 (N_58,In_430,In_145);
nand U59 (N_59,In_475,In_375);
nor U60 (N_60,In_119,In_80);
nor U61 (N_61,In_489,In_148);
nand U62 (N_62,In_77,In_462);
nand U63 (N_63,In_386,In_422);
xor U64 (N_64,In_432,In_434);
or U65 (N_65,In_409,In_283);
and U66 (N_66,In_355,In_334);
or U67 (N_67,In_123,In_56);
and U68 (N_68,In_236,In_247);
nor U69 (N_69,In_317,In_361);
or U70 (N_70,In_128,In_413);
xor U71 (N_71,In_177,In_90);
nand U72 (N_72,In_304,In_443);
and U73 (N_73,In_62,In_313);
xnor U74 (N_74,In_72,In_158);
or U75 (N_75,In_164,In_325);
nand U76 (N_76,In_83,In_218);
or U77 (N_77,In_301,In_449);
nor U78 (N_78,In_229,In_478);
or U79 (N_79,In_424,In_447);
and U80 (N_80,In_94,In_225);
and U81 (N_81,In_84,In_14);
nor U82 (N_82,In_3,In_457);
nor U83 (N_83,In_291,In_411);
or U84 (N_84,In_273,In_436);
nand U85 (N_85,In_118,In_348);
nor U86 (N_86,In_43,In_147);
nand U87 (N_87,In_246,In_404);
nor U88 (N_88,In_162,In_200);
and U89 (N_89,In_192,In_108);
nand U90 (N_90,In_141,In_479);
or U91 (N_91,In_163,In_274);
nand U92 (N_92,In_327,In_293);
nor U93 (N_93,In_425,In_415);
and U94 (N_94,In_258,In_227);
or U95 (N_95,In_60,In_71);
nand U96 (N_96,In_115,In_129);
nand U97 (N_97,In_65,In_395);
and U98 (N_98,In_253,In_367);
or U99 (N_99,In_309,In_18);
xor U100 (N_100,In_113,In_144);
or U101 (N_101,In_473,In_484);
xnor U102 (N_102,In_414,In_331);
or U103 (N_103,In_157,In_189);
or U104 (N_104,In_167,In_238);
nand U105 (N_105,In_444,In_461);
and U106 (N_106,In_185,In_418);
or U107 (N_107,In_372,In_69);
and U108 (N_108,In_138,In_33);
or U109 (N_109,In_38,In_176);
or U110 (N_110,In_32,In_12);
and U111 (N_111,In_335,In_36);
or U112 (N_112,In_398,In_267);
xnor U113 (N_113,In_40,In_51);
or U114 (N_114,In_7,In_336);
nor U115 (N_115,In_321,In_264);
nor U116 (N_116,In_285,In_102);
nor U117 (N_117,In_288,In_96);
nor U118 (N_118,In_241,In_364);
and U119 (N_119,In_310,In_455);
or U120 (N_120,In_168,In_403);
and U121 (N_121,In_178,In_15);
or U122 (N_122,In_166,In_272);
or U123 (N_123,In_254,In_160);
or U124 (N_124,In_21,In_491);
and U125 (N_125,In_222,In_295);
nor U126 (N_126,In_39,In_470);
nor U127 (N_127,In_332,In_5);
or U128 (N_128,In_257,In_13);
or U129 (N_129,In_125,In_121);
nand U130 (N_130,In_132,In_412);
nand U131 (N_131,In_356,In_392);
xor U132 (N_132,In_155,In_233);
nor U133 (N_133,In_344,In_204);
nand U134 (N_134,In_376,In_377);
nor U135 (N_135,In_26,In_378);
and U136 (N_136,In_20,In_248);
and U137 (N_137,In_59,In_459);
nand U138 (N_138,In_139,In_399);
or U139 (N_139,In_88,In_311);
and U140 (N_140,In_114,In_235);
or U141 (N_141,In_302,In_262);
and U142 (N_142,In_494,In_268);
nand U143 (N_143,In_172,In_106);
nand U144 (N_144,In_354,In_63);
xor U145 (N_145,In_223,In_130);
nand U146 (N_146,In_98,In_440);
or U147 (N_147,In_416,In_137);
and U148 (N_148,In_111,In_450);
and U149 (N_149,In_6,In_352);
or U150 (N_150,In_231,In_190);
nor U151 (N_151,In_76,In_50);
and U152 (N_152,In_198,In_429);
xnor U153 (N_153,In_250,In_460);
and U154 (N_154,In_99,In_53);
nand U155 (N_155,In_481,In_486);
and U156 (N_156,In_41,In_294);
nand U157 (N_157,In_368,In_485);
nand U158 (N_158,In_410,In_210);
and U159 (N_159,In_67,In_207);
nand U160 (N_160,In_97,In_382);
and U161 (N_161,In_381,In_463);
or U162 (N_162,In_452,In_371);
or U163 (N_163,In_58,In_366);
and U164 (N_164,In_35,In_126);
xor U165 (N_165,In_451,In_324);
nor U166 (N_166,In_251,In_465);
nand U167 (N_167,In_48,In_151);
and U168 (N_168,In_66,In_464);
xnor U169 (N_169,In_95,In_402);
or U170 (N_170,In_217,In_340);
nor U171 (N_171,In_19,In_156);
nand U172 (N_172,In_64,In_281);
nand U173 (N_173,In_193,In_370);
and U174 (N_174,In_152,In_284);
and U175 (N_175,In_173,In_394);
nor U176 (N_176,In_389,In_244);
nand U177 (N_177,In_8,In_103);
and U178 (N_178,In_112,In_480);
nor U179 (N_179,In_499,In_346);
or U180 (N_180,In_201,In_401);
or U181 (N_181,In_495,In_101);
nor U182 (N_182,In_476,In_57);
and U183 (N_183,In_183,In_423);
or U184 (N_184,In_117,In_149);
and U185 (N_185,In_345,In_493);
and U186 (N_186,In_37,In_135);
nor U187 (N_187,In_358,In_74);
nor U188 (N_188,In_333,In_205);
and U189 (N_189,In_347,In_390);
xor U190 (N_190,In_226,In_282);
xor U191 (N_191,In_468,In_299);
and U192 (N_192,In_191,In_124);
nand U193 (N_193,In_70,In_143);
nand U194 (N_194,In_420,In_184);
and U195 (N_195,In_271,In_28);
nand U196 (N_196,In_245,In_488);
or U197 (N_197,In_197,In_136);
nand U198 (N_198,In_216,In_498);
and U199 (N_199,In_323,In_4);
or U200 (N_200,In_133,In_446);
xor U201 (N_201,In_490,In_357);
nor U202 (N_202,In_242,In_249);
and U203 (N_203,In_442,In_261);
or U204 (N_204,In_213,In_308);
and U205 (N_205,In_202,In_306);
and U206 (N_206,In_17,In_349);
nor U207 (N_207,In_196,In_280);
or U208 (N_208,In_174,In_180);
nand U209 (N_209,In_153,In_278);
nand U210 (N_210,In_93,In_417);
nor U211 (N_211,In_290,In_252);
and U212 (N_212,In_441,In_92);
nand U213 (N_213,In_73,In_142);
nand U214 (N_214,In_305,In_279);
xnor U215 (N_215,In_350,In_134);
and U216 (N_216,In_237,In_116);
nand U217 (N_217,In_209,In_105);
and U218 (N_218,In_292,In_360);
and U219 (N_219,In_78,In_243);
and U220 (N_220,In_269,In_23);
nor U221 (N_221,In_298,In_239);
and U222 (N_222,In_179,In_431);
nand U223 (N_223,In_161,In_374);
nand U224 (N_224,In_379,In_296);
xnor U225 (N_225,In_181,In_277);
xor U226 (N_226,In_199,In_230);
nand U227 (N_227,In_10,In_314);
or U228 (N_228,In_219,In_337);
or U229 (N_229,In_421,In_215);
and U230 (N_230,In_466,In_186);
xor U231 (N_231,In_482,In_1);
and U232 (N_232,In_320,In_438);
xor U233 (N_233,In_435,In_42);
and U234 (N_234,In_326,In_330);
and U235 (N_235,In_29,In_195);
nand U236 (N_236,In_203,In_363);
or U237 (N_237,In_297,In_408);
or U238 (N_238,In_2,In_81);
or U239 (N_239,In_212,In_224);
or U240 (N_240,In_194,In_109);
or U241 (N_241,In_24,In_256);
xor U242 (N_242,In_171,In_328);
xor U243 (N_243,In_206,In_22);
nor U244 (N_244,In_154,In_234);
nor U245 (N_245,In_307,In_45);
or U246 (N_246,In_260,In_265);
or U247 (N_247,In_472,In_343);
and U248 (N_248,In_406,In_182);
and U249 (N_249,In_240,In_428);
or U250 (N_250,In_130,In_252);
or U251 (N_251,In_487,In_207);
xor U252 (N_252,In_355,In_135);
and U253 (N_253,In_457,In_106);
or U254 (N_254,In_396,In_264);
and U255 (N_255,In_304,In_393);
xnor U256 (N_256,In_160,In_26);
or U257 (N_257,In_118,In_209);
or U258 (N_258,In_439,In_314);
nand U259 (N_259,In_84,In_383);
nand U260 (N_260,In_64,In_469);
and U261 (N_261,In_104,In_115);
and U262 (N_262,In_143,In_441);
nor U263 (N_263,In_123,In_194);
nand U264 (N_264,In_79,In_215);
or U265 (N_265,In_444,In_269);
and U266 (N_266,In_423,In_171);
nor U267 (N_267,In_480,In_260);
nand U268 (N_268,In_38,In_215);
nand U269 (N_269,In_265,In_174);
or U270 (N_270,In_288,In_376);
and U271 (N_271,In_210,In_423);
or U272 (N_272,In_371,In_117);
and U273 (N_273,In_369,In_493);
and U274 (N_274,In_458,In_367);
nor U275 (N_275,In_272,In_23);
xor U276 (N_276,In_285,In_176);
and U277 (N_277,In_156,In_432);
or U278 (N_278,In_13,In_72);
xnor U279 (N_279,In_0,In_490);
xor U280 (N_280,In_494,In_433);
nor U281 (N_281,In_391,In_454);
nand U282 (N_282,In_42,In_44);
or U283 (N_283,In_119,In_285);
xnor U284 (N_284,In_141,In_68);
or U285 (N_285,In_107,In_198);
nor U286 (N_286,In_67,In_483);
or U287 (N_287,In_44,In_56);
and U288 (N_288,In_289,In_358);
nor U289 (N_289,In_348,In_315);
and U290 (N_290,In_91,In_119);
or U291 (N_291,In_273,In_429);
nand U292 (N_292,In_237,In_292);
xnor U293 (N_293,In_82,In_154);
nor U294 (N_294,In_495,In_137);
and U295 (N_295,In_258,In_339);
nand U296 (N_296,In_222,In_349);
or U297 (N_297,In_268,In_297);
nor U298 (N_298,In_486,In_14);
nor U299 (N_299,In_95,In_224);
nand U300 (N_300,In_208,In_130);
xnor U301 (N_301,In_463,In_197);
xnor U302 (N_302,In_205,In_458);
nand U303 (N_303,In_377,In_181);
nor U304 (N_304,In_311,In_156);
and U305 (N_305,In_373,In_129);
nand U306 (N_306,In_1,In_173);
and U307 (N_307,In_252,In_307);
nor U308 (N_308,In_224,In_152);
and U309 (N_309,In_102,In_403);
nor U310 (N_310,In_432,In_42);
xor U311 (N_311,In_177,In_36);
and U312 (N_312,In_278,In_102);
and U313 (N_313,In_300,In_293);
nor U314 (N_314,In_124,In_14);
and U315 (N_315,In_347,In_308);
or U316 (N_316,In_105,In_279);
xnor U317 (N_317,In_267,In_233);
nor U318 (N_318,In_277,In_141);
or U319 (N_319,In_46,In_72);
nor U320 (N_320,In_241,In_22);
nor U321 (N_321,In_33,In_245);
xnor U322 (N_322,In_231,In_426);
nand U323 (N_323,In_167,In_357);
or U324 (N_324,In_9,In_3);
and U325 (N_325,In_265,In_430);
or U326 (N_326,In_168,In_155);
and U327 (N_327,In_409,In_340);
or U328 (N_328,In_325,In_158);
nand U329 (N_329,In_246,In_472);
xnor U330 (N_330,In_435,In_433);
nand U331 (N_331,In_205,In_443);
and U332 (N_332,In_182,In_387);
nor U333 (N_333,In_268,In_182);
or U334 (N_334,In_409,In_401);
nor U335 (N_335,In_256,In_482);
nor U336 (N_336,In_63,In_473);
or U337 (N_337,In_426,In_116);
nor U338 (N_338,In_429,In_30);
or U339 (N_339,In_233,In_0);
nand U340 (N_340,In_53,In_170);
or U341 (N_341,In_265,In_299);
and U342 (N_342,In_315,In_333);
or U343 (N_343,In_348,In_225);
nand U344 (N_344,In_382,In_390);
nor U345 (N_345,In_191,In_151);
nor U346 (N_346,In_256,In_364);
nor U347 (N_347,In_68,In_25);
nand U348 (N_348,In_487,In_432);
nand U349 (N_349,In_458,In_396);
and U350 (N_350,In_260,In_479);
and U351 (N_351,In_389,In_276);
or U352 (N_352,In_60,In_486);
nor U353 (N_353,In_44,In_50);
or U354 (N_354,In_15,In_363);
or U355 (N_355,In_483,In_240);
nor U356 (N_356,In_141,In_110);
nand U357 (N_357,In_164,In_400);
xor U358 (N_358,In_103,In_117);
or U359 (N_359,In_131,In_164);
nand U360 (N_360,In_484,In_200);
or U361 (N_361,In_480,In_159);
nor U362 (N_362,In_150,In_107);
nor U363 (N_363,In_390,In_260);
and U364 (N_364,In_79,In_91);
or U365 (N_365,In_143,In_21);
or U366 (N_366,In_440,In_150);
or U367 (N_367,In_341,In_139);
nor U368 (N_368,In_406,In_454);
nor U369 (N_369,In_51,In_70);
or U370 (N_370,In_430,In_292);
and U371 (N_371,In_476,In_31);
and U372 (N_372,In_105,In_124);
nor U373 (N_373,In_457,In_464);
and U374 (N_374,In_173,In_45);
nor U375 (N_375,In_68,In_224);
and U376 (N_376,In_258,In_453);
xor U377 (N_377,In_455,In_71);
or U378 (N_378,In_164,In_192);
or U379 (N_379,In_72,In_485);
nand U380 (N_380,In_486,In_62);
nand U381 (N_381,In_124,In_140);
nand U382 (N_382,In_47,In_14);
nor U383 (N_383,In_474,In_431);
nand U384 (N_384,In_254,In_457);
or U385 (N_385,In_111,In_178);
or U386 (N_386,In_104,In_496);
and U387 (N_387,In_105,In_317);
nor U388 (N_388,In_1,In_223);
xnor U389 (N_389,In_147,In_339);
nand U390 (N_390,In_387,In_16);
or U391 (N_391,In_385,In_399);
and U392 (N_392,In_169,In_329);
nand U393 (N_393,In_379,In_83);
nand U394 (N_394,In_20,In_367);
nor U395 (N_395,In_152,In_193);
nor U396 (N_396,In_156,In_131);
and U397 (N_397,In_216,In_319);
or U398 (N_398,In_1,In_273);
xnor U399 (N_399,In_401,In_96);
nor U400 (N_400,In_468,In_356);
or U401 (N_401,In_175,In_469);
nand U402 (N_402,In_354,In_421);
and U403 (N_403,In_301,In_185);
nor U404 (N_404,In_325,In_296);
nand U405 (N_405,In_368,In_41);
nor U406 (N_406,In_47,In_228);
nand U407 (N_407,In_13,In_79);
nand U408 (N_408,In_327,In_11);
or U409 (N_409,In_430,In_342);
or U410 (N_410,In_404,In_260);
or U411 (N_411,In_20,In_182);
nand U412 (N_412,In_287,In_173);
or U413 (N_413,In_134,In_93);
nand U414 (N_414,In_169,In_356);
nand U415 (N_415,In_276,In_79);
or U416 (N_416,In_415,In_454);
nand U417 (N_417,In_195,In_11);
xnor U418 (N_418,In_39,In_45);
or U419 (N_419,In_101,In_120);
xor U420 (N_420,In_214,In_256);
nor U421 (N_421,In_236,In_436);
xor U422 (N_422,In_116,In_425);
nand U423 (N_423,In_286,In_416);
xor U424 (N_424,In_291,In_103);
nor U425 (N_425,In_216,In_7);
nor U426 (N_426,In_210,In_176);
nand U427 (N_427,In_52,In_267);
or U428 (N_428,In_93,In_389);
nand U429 (N_429,In_329,In_174);
nand U430 (N_430,In_300,In_364);
and U431 (N_431,In_216,In_409);
xnor U432 (N_432,In_416,In_433);
and U433 (N_433,In_265,In_406);
nor U434 (N_434,In_2,In_428);
and U435 (N_435,In_136,In_266);
or U436 (N_436,In_425,In_8);
and U437 (N_437,In_8,In_428);
and U438 (N_438,In_141,In_458);
or U439 (N_439,In_205,In_326);
xnor U440 (N_440,In_21,In_63);
nand U441 (N_441,In_218,In_374);
nand U442 (N_442,In_335,In_87);
and U443 (N_443,In_271,In_415);
and U444 (N_444,In_193,In_153);
nor U445 (N_445,In_136,In_439);
nand U446 (N_446,In_15,In_353);
or U447 (N_447,In_61,In_152);
nand U448 (N_448,In_421,In_442);
nand U449 (N_449,In_5,In_280);
and U450 (N_450,In_344,In_70);
xor U451 (N_451,In_280,In_15);
and U452 (N_452,In_263,In_496);
or U453 (N_453,In_171,In_432);
or U454 (N_454,In_434,In_425);
and U455 (N_455,In_50,In_323);
xor U456 (N_456,In_301,In_441);
and U457 (N_457,In_453,In_128);
xnor U458 (N_458,In_60,In_180);
nor U459 (N_459,In_143,In_251);
or U460 (N_460,In_226,In_197);
nand U461 (N_461,In_193,In_452);
and U462 (N_462,In_247,In_8);
and U463 (N_463,In_471,In_432);
and U464 (N_464,In_274,In_3);
and U465 (N_465,In_144,In_129);
or U466 (N_466,In_490,In_447);
and U467 (N_467,In_282,In_247);
xor U468 (N_468,In_221,In_463);
and U469 (N_469,In_316,In_11);
or U470 (N_470,In_406,In_95);
or U471 (N_471,In_478,In_244);
nor U472 (N_472,In_65,In_392);
nand U473 (N_473,In_190,In_378);
nor U474 (N_474,In_240,In_128);
or U475 (N_475,In_143,In_442);
and U476 (N_476,In_164,In_139);
nand U477 (N_477,In_236,In_54);
nand U478 (N_478,In_290,In_470);
xor U479 (N_479,In_338,In_247);
nor U480 (N_480,In_204,In_71);
nand U481 (N_481,In_4,In_315);
or U482 (N_482,In_415,In_205);
or U483 (N_483,In_312,In_417);
nand U484 (N_484,In_263,In_134);
nand U485 (N_485,In_284,In_91);
nor U486 (N_486,In_22,In_420);
nor U487 (N_487,In_266,In_137);
nor U488 (N_488,In_37,In_464);
xor U489 (N_489,In_197,In_48);
nor U490 (N_490,In_493,In_395);
nand U491 (N_491,In_409,In_272);
nor U492 (N_492,In_23,In_261);
nand U493 (N_493,In_399,In_110);
nand U494 (N_494,In_365,In_437);
xnor U495 (N_495,In_464,In_260);
nor U496 (N_496,In_415,In_329);
nor U497 (N_497,In_24,In_161);
nand U498 (N_498,In_118,In_373);
nand U499 (N_499,In_302,In_465);
or U500 (N_500,In_45,In_129);
and U501 (N_501,In_267,In_190);
nor U502 (N_502,In_384,In_259);
xnor U503 (N_503,In_231,In_309);
or U504 (N_504,In_383,In_227);
and U505 (N_505,In_59,In_131);
and U506 (N_506,In_351,In_228);
nand U507 (N_507,In_482,In_425);
nand U508 (N_508,In_309,In_42);
or U509 (N_509,In_342,In_188);
nand U510 (N_510,In_463,In_468);
nand U511 (N_511,In_405,In_322);
or U512 (N_512,In_312,In_264);
nor U513 (N_513,In_270,In_195);
or U514 (N_514,In_100,In_168);
and U515 (N_515,In_299,In_428);
and U516 (N_516,In_461,In_378);
or U517 (N_517,In_88,In_153);
and U518 (N_518,In_89,In_459);
and U519 (N_519,In_84,In_252);
or U520 (N_520,In_345,In_219);
and U521 (N_521,In_110,In_396);
nand U522 (N_522,In_457,In_316);
nor U523 (N_523,In_426,In_168);
or U524 (N_524,In_379,In_331);
or U525 (N_525,In_138,In_190);
and U526 (N_526,In_85,In_466);
or U527 (N_527,In_185,In_52);
nor U528 (N_528,In_11,In_418);
or U529 (N_529,In_395,In_78);
or U530 (N_530,In_152,In_155);
and U531 (N_531,In_363,In_153);
nand U532 (N_532,In_457,In_95);
nor U533 (N_533,In_286,In_172);
and U534 (N_534,In_321,In_5);
xor U535 (N_535,In_45,In_275);
nor U536 (N_536,In_32,In_375);
or U537 (N_537,In_90,In_372);
and U538 (N_538,In_45,In_110);
nor U539 (N_539,In_414,In_333);
xnor U540 (N_540,In_46,In_154);
and U541 (N_541,In_330,In_33);
or U542 (N_542,In_69,In_479);
or U543 (N_543,In_312,In_304);
and U544 (N_544,In_140,In_112);
and U545 (N_545,In_486,In_334);
nand U546 (N_546,In_412,In_296);
nand U547 (N_547,In_272,In_195);
nand U548 (N_548,In_358,In_477);
and U549 (N_549,In_300,In_280);
or U550 (N_550,In_130,In_182);
or U551 (N_551,In_201,In_205);
or U552 (N_552,In_230,In_112);
or U553 (N_553,In_407,In_346);
nor U554 (N_554,In_374,In_455);
nand U555 (N_555,In_305,In_306);
and U556 (N_556,In_326,In_173);
nand U557 (N_557,In_8,In_85);
or U558 (N_558,In_252,In_207);
and U559 (N_559,In_408,In_34);
or U560 (N_560,In_490,In_302);
or U561 (N_561,In_341,In_289);
or U562 (N_562,In_97,In_232);
nor U563 (N_563,In_353,In_51);
nand U564 (N_564,In_206,In_13);
nand U565 (N_565,In_417,In_157);
xor U566 (N_566,In_434,In_474);
and U567 (N_567,In_283,In_242);
nor U568 (N_568,In_487,In_266);
and U569 (N_569,In_175,In_307);
or U570 (N_570,In_496,In_53);
and U571 (N_571,In_215,In_198);
nand U572 (N_572,In_406,In_369);
xor U573 (N_573,In_406,In_297);
and U574 (N_574,In_111,In_466);
nor U575 (N_575,In_494,In_75);
or U576 (N_576,In_216,In_387);
or U577 (N_577,In_74,In_201);
nor U578 (N_578,In_195,In_122);
or U579 (N_579,In_13,In_171);
xnor U580 (N_580,In_471,In_320);
xor U581 (N_581,In_79,In_136);
or U582 (N_582,In_443,In_94);
nor U583 (N_583,In_373,In_402);
nor U584 (N_584,In_391,In_226);
and U585 (N_585,In_270,In_243);
xnor U586 (N_586,In_9,In_331);
xnor U587 (N_587,In_216,In_217);
and U588 (N_588,In_41,In_272);
nor U589 (N_589,In_283,In_83);
or U590 (N_590,In_128,In_64);
and U591 (N_591,In_160,In_228);
xnor U592 (N_592,In_289,In_494);
and U593 (N_593,In_58,In_411);
or U594 (N_594,In_458,In_79);
nor U595 (N_595,In_117,In_298);
nand U596 (N_596,In_46,In_232);
and U597 (N_597,In_85,In_410);
and U598 (N_598,In_490,In_408);
nand U599 (N_599,In_263,In_35);
xnor U600 (N_600,In_195,In_385);
or U601 (N_601,In_381,In_306);
or U602 (N_602,In_176,In_338);
nand U603 (N_603,In_60,In_178);
nand U604 (N_604,In_299,In_210);
xor U605 (N_605,In_479,In_380);
or U606 (N_606,In_271,In_76);
and U607 (N_607,In_425,In_454);
nor U608 (N_608,In_42,In_298);
xor U609 (N_609,In_129,In_255);
or U610 (N_610,In_105,In_336);
or U611 (N_611,In_450,In_488);
and U612 (N_612,In_403,In_253);
nor U613 (N_613,In_426,In_266);
nand U614 (N_614,In_325,In_456);
nor U615 (N_615,In_112,In_106);
nand U616 (N_616,In_124,In_110);
or U617 (N_617,In_273,In_299);
or U618 (N_618,In_354,In_366);
or U619 (N_619,In_81,In_33);
or U620 (N_620,In_458,In_123);
and U621 (N_621,In_426,In_153);
or U622 (N_622,In_98,In_390);
nor U623 (N_623,In_46,In_197);
nor U624 (N_624,In_327,In_406);
and U625 (N_625,In_360,In_372);
nand U626 (N_626,In_442,In_61);
and U627 (N_627,In_81,In_456);
nor U628 (N_628,In_371,In_473);
and U629 (N_629,In_61,In_156);
nor U630 (N_630,In_327,In_218);
nor U631 (N_631,In_133,In_422);
or U632 (N_632,In_198,In_239);
or U633 (N_633,In_35,In_462);
or U634 (N_634,In_62,In_355);
nor U635 (N_635,In_275,In_89);
and U636 (N_636,In_434,In_214);
or U637 (N_637,In_380,In_323);
nor U638 (N_638,In_448,In_251);
xor U639 (N_639,In_433,In_377);
nand U640 (N_640,In_480,In_267);
nor U641 (N_641,In_493,In_161);
nand U642 (N_642,In_481,In_343);
nor U643 (N_643,In_158,In_239);
xnor U644 (N_644,In_199,In_197);
and U645 (N_645,In_368,In_437);
nand U646 (N_646,In_297,In_251);
nand U647 (N_647,In_38,In_444);
and U648 (N_648,In_341,In_402);
xnor U649 (N_649,In_0,In_439);
nor U650 (N_650,In_380,In_307);
or U651 (N_651,In_479,In_246);
nor U652 (N_652,In_61,In_376);
or U653 (N_653,In_70,In_380);
or U654 (N_654,In_106,In_456);
nand U655 (N_655,In_55,In_158);
nor U656 (N_656,In_454,In_280);
nor U657 (N_657,In_267,In_421);
nand U658 (N_658,In_156,In_442);
or U659 (N_659,In_325,In_202);
or U660 (N_660,In_477,In_432);
xor U661 (N_661,In_378,In_49);
and U662 (N_662,In_403,In_110);
or U663 (N_663,In_55,In_66);
and U664 (N_664,In_352,In_397);
or U665 (N_665,In_21,In_324);
and U666 (N_666,In_383,In_295);
nand U667 (N_667,In_154,In_75);
nor U668 (N_668,In_358,In_373);
nand U669 (N_669,In_499,In_264);
nor U670 (N_670,In_449,In_374);
and U671 (N_671,In_474,In_2);
and U672 (N_672,In_356,In_442);
and U673 (N_673,In_252,In_114);
and U674 (N_674,In_381,In_466);
or U675 (N_675,In_342,In_275);
and U676 (N_676,In_121,In_419);
xnor U677 (N_677,In_362,In_379);
and U678 (N_678,In_463,In_17);
nand U679 (N_679,In_296,In_478);
and U680 (N_680,In_380,In_321);
and U681 (N_681,In_268,In_100);
nor U682 (N_682,In_392,In_228);
nand U683 (N_683,In_98,In_296);
nor U684 (N_684,In_329,In_263);
or U685 (N_685,In_93,In_379);
nor U686 (N_686,In_291,In_499);
nand U687 (N_687,In_283,In_457);
and U688 (N_688,In_444,In_278);
or U689 (N_689,In_492,In_312);
nor U690 (N_690,In_269,In_212);
nand U691 (N_691,In_192,In_472);
and U692 (N_692,In_325,In_37);
or U693 (N_693,In_224,In_148);
xnor U694 (N_694,In_487,In_440);
and U695 (N_695,In_148,In_439);
nand U696 (N_696,In_472,In_426);
and U697 (N_697,In_82,In_10);
and U698 (N_698,In_114,In_272);
and U699 (N_699,In_178,In_41);
and U700 (N_700,In_393,In_282);
or U701 (N_701,In_96,In_340);
and U702 (N_702,In_279,In_202);
nand U703 (N_703,In_461,In_170);
nand U704 (N_704,In_309,In_280);
or U705 (N_705,In_466,In_3);
nor U706 (N_706,In_15,In_490);
nand U707 (N_707,In_185,In_362);
and U708 (N_708,In_145,In_312);
nand U709 (N_709,In_188,In_91);
nand U710 (N_710,In_6,In_65);
nor U711 (N_711,In_42,In_175);
and U712 (N_712,In_109,In_403);
nand U713 (N_713,In_288,In_346);
nor U714 (N_714,In_190,In_445);
and U715 (N_715,In_66,In_251);
and U716 (N_716,In_333,In_428);
or U717 (N_717,In_57,In_89);
nor U718 (N_718,In_36,In_240);
nor U719 (N_719,In_264,In_344);
and U720 (N_720,In_246,In_392);
nor U721 (N_721,In_221,In_17);
nand U722 (N_722,In_17,In_454);
nor U723 (N_723,In_157,In_392);
and U724 (N_724,In_317,In_187);
nand U725 (N_725,In_229,In_46);
nand U726 (N_726,In_484,In_205);
or U727 (N_727,In_290,In_370);
nor U728 (N_728,In_271,In_134);
or U729 (N_729,In_143,In_27);
nor U730 (N_730,In_337,In_33);
and U731 (N_731,In_474,In_496);
nand U732 (N_732,In_238,In_59);
and U733 (N_733,In_445,In_442);
nor U734 (N_734,In_260,In_73);
and U735 (N_735,In_100,In_397);
nand U736 (N_736,In_19,In_394);
nand U737 (N_737,In_24,In_354);
nand U738 (N_738,In_0,In_214);
nand U739 (N_739,In_375,In_285);
nor U740 (N_740,In_422,In_354);
and U741 (N_741,In_10,In_14);
nor U742 (N_742,In_134,In_237);
nand U743 (N_743,In_73,In_415);
nor U744 (N_744,In_6,In_315);
or U745 (N_745,In_321,In_83);
nor U746 (N_746,In_36,In_431);
or U747 (N_747,In_398,In_15);
and U748 (N_748,In_251,In_199);
and U749 (N_749,In_256,In_19);
or U750 (N_750,N_227,N_425);
nor U751 (N_751,N_86,N_666);
and U752 (N_752,N_557,N_741);
or U753 (N_753,N_360,N_132);
nand U754 (N_754,N_598,N_239);
or U755 (N_755,N_603,N_555);
or U756 (N_756,N_322,N_229);
nand U757 (N_757,N_709,N_325);
and U758 (N_758,N_188,N_34);
or U759 (N_759,N_250,N_393);
nand U760 (N_760,N_430,N_120);
nor U761 (N_761,N_33,N_328);
xor U762 (N_762,N_205,N_156);
or U763 (N_763,N_451,N_219);
nor U764 (N_764,N_150,N_542);
nand U765 (N_765,N_53,N_572);
and U766 (N_766,N_701,N_100);
nor U767 (N_767,N_584,N_345);
nor U768 (N_768,N_392,N_333);
or U769 (N_769,N_658,N_577);
or U770 (N_770,N_251,N_326);
nor U771 (N_771,N_614,N_266);
nand U772 (N_772,N_298,N_35);
and U773 (N_773,N_65,N_565);
nor U774 (N_774,N_29,N_58);
nor U775 (N_775,N_471,N_122);
and U776 (N_776,N_302,N_276);
nor U777 (N_777,N_330,N_573);
and U778 (N_778,N_605,N_165);
xor U779 (N_779,N_726,N_138);
nand U780 (N_780,N_194,N_151);
and U781 (N_781,N_59,N_129);
nor U782 (N_782,N_559,N_369);
nand U783 (N_783,N_140,N_288);
xor U784 (N_784,N_331,N_745);
and U785 (N_785,N_632,N_351);
and U786 (N_786,N_622,N_353);
nor U787 (N_787,N_747,N_109);
or U788 (N_788,N_422,N_95);
xnor U789 (N_789,N_241,N_108);
nor U790 (N_790,N_667,N_599);
nor U791 (N_791,N_261,N_399);
and U792 (N_792,N_190,N_230);
nand U793 (N_793,N_708,N_715);
nor U794 (N_794,N_636,N_509);
nand U795 (N_795,N_597,N_304);
and U796 (N_796,N_182,N_590);
nor U797 (N_797,N_394,N_737);
or U798 (N_798,N_349,N_284);
nand U799 (N_799,N_44,N_653);
nor U800 (N_800,N_245,N_20);
xor U801 (N_801,N_327,N_635);
xor U802 (N_802,N_593,N_591);
nand U803 (N_803,N_541,N_644);
nor U804 (N_804,N_534,N_270);
xnor U805 (N_805,N_493,N_407);
or U806 (N_806,N_515,N_136);
and U807 (N_807,N_134,N_640);
or U808 (N_808,N_633,N_544);
nor U809 (N_809,N_69,N_704);
nand U810 (N_810,N_160,N_476);
nor U811 (N_811,N_528,N_348);
nand U812 (N_812,N_153,N_660);
xnor U813 (N_813,N_228,N_490);
xnor U814 (N_814,N_66,N_200);
nand U815 (N_815,N_434,N_426);
and U816 (N_816,N_17,N_255);
nand U817 (N_817,N_749,N_184);
nor U818 (N_818,N_249,N_37);
and U819 (N_819,N_503,N_31);
nand U820 (N_820,N_329,N_281);
and U821 (N_821,N_525,N_400);
or U822 (N_822,N_0,N_639);
or U823 (N_823,N_512,N_114);
nor U824 (N_824,N_39,N_127);
xnor U825 (N_825,N_583,N_566);
and U826 (N_826,N_80,N_403);
or U827 (N_827,N_14,N_432);
or U828 (N_828,N_563,N_536);
nor U829 (N_829,N_11,N_556);
nand U830 (N_830,N_27,N_218);
or U831 (N_831,N_621,N_712);
or U832 (N_832,N_15,N_113);
nor U833 (N_833,N_102,N_22);
nor U834 (N_834,N_208,N_562);
nor U835 (N_835,N_665,N_152);
nand U836 (N_836,N_375,N_339);
and U837 (N_837,N_76,N_111);
and U838 (N_838,N_193,N_404);
nor U839 (N_839,N_693,N_88);
nand U840 (N_840,N_454,N_549);
and U841 (N_841,N_92,N_3);
nand U842 (N_842,N_306,N_180);
xor U843 (N_843,N_386,N_604);
nor U844 (N_844,N_607,N_179);
or U845 (N_845,N_651,N_519);
and U846 (N_846,N_161,N_697);
or U847 (N_847,N_668,N_531);
nand U848 (N_848,N_125,N_104);
and U849 (N_849,N_652,N_547);
and U850 (N_850,N_481,N_681);
nand U851 (N_851,N_199,N_497);
and U852 (N_852,N_10,N_722);
nor U853 (N_853,N_352,N_689);
nand U854 (N_854,N_535,N_647);
nand U855 (N_855,N_378,N_702);
nor U856 (N_856,N_207,N_543);
xor U857 (N_857,N_615,N_720);
or U858 (N_858,N_195,N_540);
nand U859 (N_859,N_506,N_474);
xor U860 (N_860,N_222,N_455);
nand U861 (N_861,N_81,N_415);
nor U862 (N_862,N_587,N_265);
nand U863 (N_863,N_738,N_456);
or U864 (N_864,N_740,N_370);
nor U865 (N_865,N_106,N_387);
or U866 (N_866,N_686,N_186);
or U867 (N_867,N_619,N_52);
xnor U868 (N_868,N_552,N_260);
and U869 (N_869,N_68,N_417);
nand U870 (N_870,N_642,N_680);
nand U871 (N_871,N_428,N_629);
or U872 (N_872,N_297,N_406);
nand U873 (N_873,N_649,N_271);
nor U874 (N_874,N_739,N_731);
and U875 (N_875,N_287,N_162);
nor U876 (N_876,N_61,N_742);
nand U877 (N_877,N_453,N_418);
nor U878 (N_878,N_468,N_643);
and U879 (N_879,N_719,N_168);
xor U880 (N_880,N_486,N_582);
nor U881 (N_881,N_83,N_508);
or U882 (N_882,N_706,N_63);
or U883 (N_883,N_487,N_424);
nor U884 (N_884,N_588,N_146);
nand U885 (N_885,N_214,N_172);
xor U886 (N_886,N_334,N_70);
or U887 (N_887,N_128,N_744);
nor U888 (N_888,N_459,N_93);
and U889 (N_889,N_254,N_209);
and U890 (N_890,N_256,N_291);
nand U891 (N_891,N_317,N_376);
nand U892 (N_892,N_638,N_142);
nand U893 (N_893,N_673,N_514);
and U894 (N_894,N_324,N_383);
nor U895 (N_895,N_247,N_183);
or U896 (N_896,N_283,N_380);
nand U897 (N_897,N_494,N_585);
and U898 (N_898,N_602,N_191);
nor U899 (N_899,N_498,N_171);
nor U900 (N_900,N_561,N_714);
nor U901 (N_901,N_727,N_437);
nand U902 (N_902,N_101,N_467);
or U903 (N_903,N_401,N_650);
nor U904 (N_904,N_610,N_117);
nor U905 (N_905,N_252,N_275);
nor U906 (N_906,N_442,N_212);
xor U907 (N_907,N_396,N_47);
or U908 (N_908,N_410,N_6);
xnor U909 (N_909,N_594,N_734);
nand U910 (N_910,N_21,N_55);
nor U911 (N_911,N_682,N_38);
nor U912 (N_912,N_592,N_743);
nand U913 (N_913,N_159,N_688);
nand U914 (N_914,N_505,N_564);
nor U915 (N_915,N_144,N_164);
nand U916 (N_916,N_596,N_595);
nand U917 (N_917,N_475,N_289);
xnor U918 (N_918,N_700,N_262);
or U919 (N_919,N_463,N_41);
and U920 (N_920,N_457,N_350);
nor U921 (N_921,N_612,N_377);
and U922 (N_922,N_174,N_309);
xnor U923 (N_923,N_630,N_238);
or U924 (N_924,N_570,N_539);
nor U925 (N_925,N_634,N_517);
and U926 (N_926,N_576,N_176);
nand U927 (N_927,N_620,N_705);
xnor U928 (N_928,N_367,N_385);
and U929 (N_929,N_196,N_50);
nor U930 (N_930,N_628,N_692);
and U931 (N_931,N_464,N_248);
nor U932 (N_932,N_641,N_90);
and U933 (N_933,N_272,N_13);
nand U934 (N_934,N_413,N_358);
nor U935 (N_935,N_197,N_145);
or U936 (N_936,N_560,N_683);
nor U937 (N_937,N_480,N_264);
nand U938 (N_938,N_389,N_43);
and U939 (N_939,N_450,N_374);
xnor U940 (N_940,N_510,N_518);
nor U941 (N_941,N_24,N_85);
nand U942 (N_942,N_443,N_500);
or U943 (N_943,N_321,N_589);
and U944 (N_944,N_362,N_571);
or U945 (N_945,N_648,N_491);
nor U946 (N_946,N_492,N_391);
nand U947 (N_947,N_381,N_316);
and U948 (N_948,N_724,N_645);
nand U949 (N_949,N_82,N_233);
xor U950 (N_950,N_520,N_126);
and U951 (N_951,N_263,N_390);
and U952 (N_952,N_716,N_246);
nor U953 (N_953,N_123,N_397);
nand U954 (N_954,N_567,N_273);
nand U955 (N_955,N_730,N_449);
xor U956 (N_956,N_569,N_355);
nand U957 (N_957,N_347,N_242);
nor U958 (N_958,N_96,N_223);
or U959 (N_959,N_746,N_421);
nand U960 (N_960,N_54,N_60);
nand U961 (N_961,N_365,N_478);
nand U962 (N_962,N_473,N_189);
and U963 (N_963,N_729,N_439);
and U964 (N_964,N_48,N_732);
or U965 (N_965,N_616,N_431);
nand U966 (N_966,N_67,N_553);
nor U967 (N_967,N_409,N_600);
or U968 (N_968,N_574,N_575);
and U969 (N_969,N_513,N_684);
and U970 (N_970,N_177,N_346);
xnor U971 (N_971,N_698,N_670);
or U972 (N_972,N_606,N_8);
nand U973 (N_973,N_279,N_213);
nor U974 (N_974,N_16,N_78);
and U975 (N_975,N_303,N_496);
or U976 (N_976,N_408,N_372);
and U977 (N_977,N_466,N_416);
and U978 (N_978,N_135,N_235);
and U979 (N_979,N_234,N_669);
xnor U980 (N_980,N_226,N_268);
nor U981 (N_981,N_656,N_343);
and U982 (N_982,N_672,N_112);
or U983 (N_983,N_484,N_354);
and U984 (N_984,N_141,N_45);
nor U985 (N_985,N_94,N_659);
nor U986 (N_986,N_320,N_98);
and U987 (N_987,N_568,N_299);
or U988 (N_988,N_119,N_655);
xnor U989 (N_989,N_472,N_691);
and U990 (N_990,N_411,N_315);
or U991 (N_991,N_269,N_359);
nand U992 (N_992,N_626,N_545);
nand U993 (N_993,N_26,N_436);
or U994 (N_994,N_723,N_32);
nor U995 (N_995,N_206,N_103);
or U996 (N_996,N_72,N_115);
and U997 (N_997,N_625,N_580);
or U998 (N_998,N_290,N_538);
xor U999 (N_999,N_601,N_91);
xor U1000 (N_1000,N_465,N_460);
and U1001 (N_1001,N_725,N_277);
nand U1002 (N_1002,N_373,N_296);
and U1003 (N_1003,N_139,N_295);
xor U1004 (N_1004,N_257,N_361);
and U1005 (N_1005,N_25,N_446);
nand U1006 (N_1006,N_637,N_447);
nor U1007 (N_1007,N_19,N_504);
and U1008 (N_1008,N_458,N_7);
and U1009 (N_1009,N_395,N_198);
or U1010 (N_1010,N_579,N_558);
nor U1011 (N_1011,N_618,N_533);
and U1012 (N_1012,N_149,N_608);
nand U1013 (N_1013,N_546,N_728);
nor U1014 (N_1014,N_121,N_57);
and U1015 (N_1015,N_323,N_51);
and U1016 (N_1016,N_501,N_676);
and U1017 (N_1017,N_2,N_312);
nor U1018 (N_1018,N_657,N_671);
xor U1019 (N_1019,N_527,N_499);
or U1020 (N_1020,N_4,N_157);
nor U1021 (N_1021,N_523,N_366);
nand U1022 (N_1022,N_1,N_548);
xnor U1023 (N_1023,N_217,N_445);
nor U1024 (N_1024,N_718,N_294);
xnor U1025 (N_1025,N_166,N_364);
or U1026 (N_1026,N_319,N_201);
or U1027 (N_1027,N_9,N_532);
and U1028 (N_1028,N_232,N_178);
or U1029 (N_1029,N_663,N_71);
or U1030 (N_1030,N_748,N_419);
and U1031 (N_1031,N_694,N_721);
nor U1032 (N_1032,N_357,N_259);
xor U1033 (N_1033,N_733,N_89);
or U1034 (N_1034,N_522,N_516);
or U1035 (N_1035,N_384,N_130);
nor U1036 (N_1036,N_46,N_307);
nor U1037 (N_1037,N_97,N_736);
xor U1038 (N_1038,N_342,N_131);
nand U1039 (N_1039,N_405,N_511);
nor U1040 (N_1040,N_285,N_267);
or U1041 (N_1041,N_479,N_550);
xor U1042 (N_1042,N_489,N_105);
nand U1043 (N_1043,N_335,N_203);
nor U1044 (N_1044,N_448,N_382);
nor U1045 (N_1045,N_163,N_631);
or U1046 (N_1046,N_236,N_202);
or U1047 (N_1047,N_707,N_664);
nand U1048 (N_1048,N_332,N_675);
and U1049 (N_1049,N_154,N_99);
nand U1050 (N_1050,N_687,N_107);
or U1051 (N_1051,N_23,N_578);
nand U1052 (N_1052,N_735,N_73);
or U1053 (N_1053,N_215,N_427);
and U1054 (N_1054,N_305,N_158);
and U1055 (N_1055,N_170,N_711);
or U1056 (N_1056,N_87,N_133);
and U1057 (N_1057,N_495,N_175);
nor U1058 (N_1058,N_192,N_338);
nand U1059 (N_1059,N_274,N_482);
and U1060 (N_1060,N_696,N_661);
xnor U1061 (N_1061,N_581,N_18);
nand U1062 (N_1062,N_340,N_356);
nand U1063 (N_1063,N_116,N_155);
nor U1064 (N_1064,N_703,N_662);
nand U1065 (N_1065,N_64,N_678);
and U1066 (N_1066,N_363,N_586);
and U1067 (N_1067,N_440,N_677);
nand U1068 (N_1068,N_685,N_237);
nor U1069 (N_1069,N_485,N_314);
and U1070 (N_1070,N_414,N_646);
nor U1071 (N_1071,N_204,N_221);
or U1072 (N_1072,N_185,N_402);
nor U1073 (N_1073,N_613,N_293);
nor U1074 (N_1074,N_167,N_529);
xnor U1075 (N_1075,N_12,N_477);
nor U1076 (N_1076,N_282,N_674);
and U1077 (N_1077,N_62,N_624);
and U1078 (N_1078,N_713,N_617);
xnor U1079 (N_1079,N_341,N_169);
and U1080 (N_1080,N_181,N_379);
or U1081 (N_1081,N_137,N_224);
nand U1082 (N_1082,N_280,N_258);
and U1083 (N_1083,N_173,N_286);
and U1084 (N_1084,N_79,N_253);
and U1085 (N_1085,N_398,N_110);
nand U1086 (N_1086,N_147,N_452);
or U1087 (N_1087,N_231,N_240);
or U1088 (N_1088,N_461,N_56);
and U1089 (N_1089,N_695,N_717);
nor U1090 (N_1090,N_530,N_143);
or U1091 (N_1091,N_301,N_524);
nor U1092 (N_1092,N_502,N_220);
xnor U1093 (N_1093,N_371,N_84);
and U1094 (N_1094,N_300,N_654);
nor U1095 (N_1095,N_278,N_318);
and U1096 (N_1096,N_225,N_310);
xnor U1097 (N_1097,N_187,N_42);
nand U1098 (N_1098,N_124,N_690);
or U1099 (N_1099,N_292,N_551);
nand U1100 (N_1100,N_313,N_368);
and U1101 (N_1101,N_311,N_210);
or U1102 (N_1102,N_679,N_211);
xor U1103 (N_1103,N_462,N_420);
nand U1104 (N_1104,N_337,N_336);
nor U1105 (N_1105,N_423,N_521);
xor U1106 (N_1106,N_28,N_243);
and U1107 (N_1107,N_5,N_118);
nor U1108 (N_1108,N_344,N_49);
nand U1109 (N_1109,N_77,N_611);
nor U1110 (N_1110,N_429,N_388);
nor U1111 (N_1111,N_74,N_438);
nand U1112 (N_1112,N_470,N_30);
and U1113 (N_1113,N_433,N_627);
or U1114 (N_1114,N_699,N_623);
and U1115 (N_1115,N_609,N_308);
and U1116 (N_1116,N_554,N_40);
nand U1117 (N_1117,N_483,N_244);
nand U1118 (N_1118,N_75,N_488);
nand U1119 (N_1119,N_507,N_435);
nand U1120 (N_1120,N_444,N_441);
and U1121 (N_1121,N_148,N_412);
nand U1122 (N_1122,N_36,N_710);
and U1123 (N_1123,N_469,N_216);
or U1124 (N_1124,N_526,N_537);
nor U1125 (N_1125,N_281,N_60);
or U1126 (N_1126,N_104,N_655);
nor U1127 (N_1127,N_14,N_113);
or U1128 (N_1128,N_27,N_278);
or U1129 (N_1129,N_136,N_224);
xor U1130 (N_1130,N_223,N_108);
nand U1131 (N_1131,N_178,N_349);
nor U1132 (N_1132,N_616,N_713);
nor U1133 (N_1133,N_526,N_647);
or U1134 (N_1134,N_182,N_533);
xnor U1135 (N_1135,N_644,N_9);
nor U1136 (N_1136,N_397,N_173);
and U1137 (N_1137,N_290,N_21);
and U1138 (N_1138,N_259,N_344);
and U1139 (N_1139,N_39,N_277);
nand U1140 (N_1140,N_733,N_10);
xor U1141 (N_1141,N_487,N_584);
and U1142 (N_1142,N_730,N_661);
or U1143 (N_1143,N_726,N_425);
or U1144 (N_1144,N_447,N_66);
xor U1145 (N_1145,N_91,N_613);
nand U1146 (N_1146,N_189,N_345);
or U1147 (N_1147,N_542,N_34);
or U1148 (N_1148,N_657,N_260);
nor U1149 (N_1149,N_514,N_442);
nor U1150 (N_1150,N_67,N_482);
and U1151 (N_1151,N_74,N_320);
or U1152 (N_1152,N_658,N_458);
nand U1153 (N_1153,N_369,N_539);
and U1154 (N_1154,N_308,N_433);
or U1155 (N_1155,N_727,N_567);
nand U1156 (N_1156,N_114,N_25);
or U1157 (N_1157,N_134,N_284);
nand U1158 (N_1158,N_12,N_299);
and U1159 (N_1159,N_65,N_716);
or U1160 (N_1160,N_119,N_426);
nor U1161 (N_1161,N_250,N_730);
xor U1162 (N_1162,N_626,N_89);
nor U1163 (N_1163,N_650,N_309);
nor U1164 (N_1164,N_202,N_652);
and U1165 (N_1165,N_527,N_365);
and U1166 (N_1166,N_741,N_547);
and U1167 (N_1167,N_64,N_165);
xnor U1168 (N_1168,N_290,N_599);
and U1169 (N_1169,N_595,N_269);
and U1170 (N_1170,N_96,N_30);
nor U1171 (N_1171,N_13,N_501);
nor U1172 (N_1172,N_21,N_681);
xor U1173 (N_1173,N_662,N_361);
nand U1174 (N_1174,N_226,N_706);
nor U1175 (N_1175,N_90,N_362);
and U1176 (N_1176,N_390,N_100);
and U1177 (N_1177,N_137,N_232);
nand U1178 (N_1178,N_30,N_24);
nor U1179 (N_1179,N_629,N_268);
nand U1180 (N_1180,N_179,N_302);
or U1181 (N_1181,N_392,N_453);
xor U1182 (N_1182,N_184,N_236);
or U1183 (N_1183,N_510,N_532);
or U1184 (N_1184,N_675,N_304);
nand U1185 (N_1185,N_15,N_695);
nor U1186 (N_1186,N_83,N_451);
nand U1187 (N_1187,N_206,N_220);
nand U1188 (N_1188,N_123,N_30);
nor U1189 (N_1189,N_677,N_178);
nand U1190 (N_1190,N_207,N_723);
nor U1191 (N_1191,N_483,N_131);
xor U1192 (N_1192,N_221,N_115);
nand U1193 (N_1193,N_323,N_271);
xnor U1194 (N_1194,N_231,N_427);
xnor U1195 (N_1195,N_430,N_137);
nor U1196 (N_1196,N_633,N_219);
nor U1197 (N_1197,N_321,N_77);
or U1198 (N_1198,N_483,N_381);
and U1199 (N_1199,N_561,N_607);
nand U1200 (N_1200,N_501,N_336);
and U1201 (N_1201,N_649,N_1);
or U1202 (N_1202,N_108,N_450);
or U1203 (N_1203,N_104,N_720);
and U1204 (N_1204,N_547,N_344);
and U1205 (N_1205,N_412,N_461);
and U1206 (N_1206,N_478,N_259);
and U1207 (N_1207,N_4,N_672);
and U1208 (N_1208,N_90,N_216);
nor U1209 (N_1209,N_677,N_450);
nor U1210 (N_1210,N_83,N_425);
or U1211 (N_1211,N_616,N_436);
and U1212 (N_1212,N_262,N_327);
nand U1213 (N_1213,N_193,N_71);
and U1214 (N_1214,N_592,N_68);
or U1215 (N_1215,N_238,N_229);
or U1216 (N_1216,N_417,N_432);
nand U1217 (N_1217,N_543,N_607);
nor U1218 (N_1218,N_255,N_263);
xnor U1219 (N_1219,N_21,N_220);
nand U1220 (N_1220,N_83,N_220);
and U1221 (N_1221,N_134,N_25);
nand U1222 (N_1222,N_365,N_452);
and U1223 (N_1223,N_728,N_520);
nand U1224 (N_1224,N_312,N_153);
or U1225 (N_1225,N_336,N_485);
nor U1226 (N_1226,N_492,N_723);
or U1227 (N_1227,N_350,N_371);
and U1228 (N_1228,N_416,N_423);
nor U1229 (N_1229,N_520,N_640);
xnor U1230 (N_1230,N_670,N_253);
nor U1231 (N_1231,N_325,N_14);
or U1232 (N_1232,N_693,N_617);
and U1233 (N_1233,N_325,N_561);
nand U1234 (N_1234,N_625,N_190);
nand U1235 (N_1235,N_137,N_311);
nand U1236 (N_1236,N_141,N_654);
or U1237 (N_1237,N_505,N_604);
xor U1238 (N_1238,N_444,N_298);
and U1239 (N_1239,N_250,N_646);
and U1240 (N_1240,N_729,N_525);
nand U1241 (N_1241,N_565,N_10);
xnor U1242 (N_1242,N_432,N_164);
nor U1243 (N_1243,N_179,N_419);
and U1244 (N_1244,N_623,N_358);
and U1245 (N_1245,N_4,N_140);
xor U1246 (N_1246,N_415,N_47);
and U1247 (N_1247,N_364,N_67);
nand U1248 (N_1248,N_713,N_700);
xor U1249 (N_1249,N_122,N_735);
and U1250 (N_1250,N_338,N_264);
nand U1251 (N_1251,N_253,N_320);
and U1252 (N_1252,N_155,N_630);
nand U1253 (N_1253,N_296,N_93);
or U1254 (N_1254,N_337,N_462);
or U1255 (N_1255,N_42,N_538);
and U1256 (N_1256,N_634,N_190);
nand U1257 (N_1257,N_131,N_229);
nand U1258 (N_1258,N_407,N_744);
and U1259 (N_1259,N_337,N_368);
nor U1260 (N_1260,N_262,N_402);
nor U1261 (N_1261,N_579,N_696);
nor U1262 (N_1262,N_577,N_85);
nand U1263 (N_1263,N_289,N_693);
or U1264 (N_1264,N_611,N_583);
or U1265 (N_1265,N_408,N_108);
and U1266 (N_1266,N_116,N_437);
nor U1267 (N_1267,N_598,N_433);
and U1268 (N_1268,N_548,N_665);
nand U1269 (N_1269,N_536,N_468);
nor U1270 (N_1270,N_341,N_390);
nor U1271 (N_1271,N_37,N_431);
nand U1272 (N_1272,N_670,N_226);
or U1273 (N_1273,N_683,N_131);
or U1274 (N_1274,N_709,N_172);
nor U1275 (N_1275,N_379,N_367);
nand U1276 (N_1276,N_325,N_602);
or U1277 (N_1277,N_387,N_473);
nor U1278 (N_1278,N_418,N_396);
or U1279 (N_1279,N_413,N_461);
nand U1280 (N_1280,N_222,N_49);
nor U1281 (N_1281,N_207,N_14);
nor U1282 (N_1282,N_60,N_329);
nor U1283 (N_1283,N_534,N_269);
xor U1284 (N_1284,N_256,N_325);
nor U1285 (N_1285,N_665,N_283);
and U1286 (N_1286,N_210,N_745);
nor U1287 (N_1287,N_571,N_655);
or U1288 (N_1288,N_492,N_525);
nor U1289 (N_1289,N_457,N_312);
nand U1290 (N_1290,N_253,N_220);
and U1291 (N_1291,N_502,N_180);
nor U1292 (N_1292,N_139,N_146);
nand U1293 (N_1293,N_327,N_613);
or U1294 (N_1294,N_356,N_92);
or U1295 (N_1295,N_550,N_241);
or U1296 (N_1296,N_474,N_642);
xnor U1297 (N_1297,N_407,N_146);
or U1298 (N_1298,N_348,N_59);
and U1299 (N_1299,N_484,N_653);
and U1300 (N_1300,N_112,N_593);
nor U1301 (N_1301,N_478,N_538);
xor U1302 (N_1302,N_377,N_56);
nor U1303 (N_1303,N_57,N_637);
nand U1304 (N_1304,N_322,N_22);
nor U1305 (N_1305,N_742,N_115);
and U1306 (N_1306,N_594,N_562);
or U1307 (N_1307,N_383,N_667);
nand U1308 (N_1308,N_620,N_487);
and U1309 (N_1309,N_691,N_28);
nor U1310 (N_1310,N_257,N_267);
or U1311 (N_1311,N_236,N_515);
and U1312 (N_1312,N_365,N_508);
xnor U1313 (N_1313,N_511,N_225);
nand U1314 (N_1314,N_577,N_189);
nor U1315 (N_1315,N_16,N_335);
and U1316 (N_1316,N_420,N_436);
and U1317 (N_1317,N_694,N_660);
or U1318 (N_1318,N_348,N_649);
xnor U1319 (N_1319,N_117,N_422);
nor U1320 (N_1320,N_37,N_159);
xor U1321 (N_1321,N_474,N_650);
nand U1322 (N_1322,N_101,N_246);
and U1323 (N_1323,N_167,N_276);
or U1324 (N_1324,N_227,N_404);
nor U1325 (N_1325,N_504,N_148);
nor U1326 (N_1326,N_704,N_623);
or U1327 (N_1327,N_649,N_549);
xnor U1328 (N_1328,N_63,N_647);
nand U1329 (N_1329,N_551,N_204);
and U1330 (N_1330,N_0,N_669);
xnor U1331 (N_1331,N_598,N_332);
or U1332 (N_1332,N_102,N_236);
and U1333 (N_1333,N_135,N_719);
nand U1334 (N_1334,N_246,N_650);
nor U1335 (N_1335,N_322,N_669);
and U1336 (N_1336,N_344,N_218);
and U1337 (N_1337,N_222,N_406);
nand U1338 (N_1338,N_383,N_548);
and U1339 (N_1339,N_320,N_403);
nand U1340 (N_1340,N_236,N_397);
xor U1341 (N_1341,N_97,N_430);
or U1342 (N_1342,N_341,N_36);
nor U1343 (N_1343,N_569,N_232);
and U1344 (N_1344,N_300,N_502);
xnor U1345 (N_1345,N_566,N_388);
or U1346 (N_1346,N_365,N_369);
nor U1347 (N_1347,N_443,N_491);
or U1348 (N_1348,N_426,N_164);
nand U1349 (N_1349,N_178,N_358);
and U1350 (N_1350,N_465,N_707);
xnor U1351 (N_1351,N_169,N_508);
and U1352 (N_1352,N_140,N_455);
nand U1353 (N_1353,N_435,N_56);
and U1354 (N_1354,N_280,N_68);
nor U1355 (N_1355,N_64,N_420);
xor U1356 (N_1356,N_693,N_69);
nor U1357 (N_1357,N_395,N_562);
or U1358 (N_1358,N_264,N_579);
nor U1359 (N_1359,N_617,N_15);
xnor U1360 (N_1360,N_604,N_510);
and U1361 (N_1361,N_409,N_702);
nand U1362 (N_1362,N_171,N_445);
nor U1363 (N_1363,N_516,N_351);
and U1364 (N_1364,N_402,N_144);
or U1365 (N_1365,N_437,N_502);
and U1366 (N_1366,N_62,N_736);
nor U1367 (N_1367,N_158,N_333);
or U1368 (N_1368,N_23,N_95);
xor U1369 (N_1369,N_569,N_334);
or U1370 (N_1370,N_224,N_322);
nor U1371 (N_1371,N_125,N_298);
or U1372 (N_1372,N_55,N_88);
or U1373 (N_1373,N_347,N_475);
and U1374 (N_1374,N_261,N_635);
and U1375 (N_1375,N_104,N_530);
nor U1376 (N_1376,N_144,N_423);
or U1377 (N_1377,N_30,N_502);
and U1378 (N_1378,N_402,N_455);
nand U1379 (N_1379,N_137,N_86);
nor U1380 (N_1380,N_260,N_197);
nand U1381 (N_1381,N_87,N_419);
or U1382 (N_1382,N_345,N_60);
and U1383 (N_1383,N_628,N_286);
or U1384 (N_1384,N_319,N_483);
nand U1385 (N_1385,N_12,N_40);
or U1386 (N_1386,N_296,N_439);
and U1387 (N_1387,N_380,N_654);
and U1388 (N_1388,N_508,N_92);
nor U1389 (N_1389,N_639,N_50);
nor U1390 (N_1390,N_489,N_503);
nor U1391 (N_1391,N_369,N_291);
nor U1392 (N_1392,N_620,N_114);
nor U1393 (N_1393,N_636,N_658);
nand U1394 (N_1394,N_682,N_530);
and U1395 (N_1395,N_558,N_196);
xnor U1396 (N_1396,N_491,N_387);
and U1397 (N_1397,N_706,N_580);
and U1398 (N_1398,N_460,N_408);
or U1399 (N_1399,N_456,N_596);
or U1400 (N_1400,N_264,N_35);
xnor U1401 (N_1401,N_357,N_575);
or U1402 (N_1402,N_734,N_14);
nor U1403 (N_1403,N_530,N_399);
and U1404 (N_1404,N_367,N_16);
or U1405 (N_1405,N_46,N_386);
nor U1406 (N_1406,N_184,N_197);
nand U1407 (N_1407,N_183,N_107);
nand U1408 (N_1408,N_607,N_388);
and U1409 (N_1409,N_83,N_73);
nor U1410 (N_1410,N_204,N_530);
xor U1411 (N_1411,N_574,N_240);
xor U1412 (N_1412,N_296,N_370);
nand U1413 (N_1413,N_628,N_682);
and U1414 (N_1414,N_428,N_567);
nor U1415 (N_1415,N_518,N_92);
nor U1416 (N_1416,N_51,N_641);
nand U1417 (N_1417,N_746,N_568);
and U1418 (N_1418,N_362,N_625);
or U1419 (N_1419,N_254,N_276);
or U1420 (N_1420,N_461,N_675);
xor U1421 (N_1421,N_650,N_180);
nor U1422 (N_1422,N_33,N_6);
or U1423 (N_1423,N_49,N_680);
or U1424 (N_1424,N_359,N_624);
and U1425 (N_1425,N_190,N_185);
nor U1426 (N_1426,N_223,N_167);
xnor U1427 (N_1427,N_245,N_557);
xnor U1428 (N_1428,N_587,N_651);
nand U1429 (N_1429,N_722,N_345);
or U1430 (N_1430,N_747,N_457);
nor U1431 (N_1431,N_169,N_183);
nand U1432 (N_1432,N_578,N_743);
or U1433 (N_1433,N_36,N_435);
or U1434 (N_1434,N_107,N_560);
nor U1435 (N_1435,N_472,N_159);
and U1436 (N_1436,N_741,N_75);
and U1437 (N_1437,N_179,N_590);
or U1438 (N_1438,N_237,N_244);
nor U1439 (N_1439,N_589,N_201);
xnor U1440 (N_1440,N_438,N_657);
nand U1441 (N_1441,N_432,N_703);
and U1442 (N_1442,N_512,N_431);
nand U1443 (N_1443,N_556,N_188);
and U1444 (N_1444,N_632,N_494);
or U1445 (N_1445,N_623,N_348);
and U1446 (N_1446,N_692,N_474);
nand U1447 (N_1447,N_334,N_371);
or U1448 (N_1448,N_44,N_334);
or U1449 (N_1449,N_682,N_98);
nor U1450 (N_1450,N_99,N_62);
nor U1451 (N_1451,N_271,N_343);
nand U1452 (N_1452,N_489,N_116);
and U1453 (N_1453,N_662,N_711);
nand U1454 (N_1454,N_39,N_154);
or U1455 (N_1455,N_411,N_395);
nand U1456 (N_1456,N_705,N_254);
nand U1457 (N_1457,N_197,N_27);
nand U1458 (N_1458,N_460,N_334);
or U1459 (N_1459,N_480,N_601);
or U1460 (N_1460,N_143,N_624);
or U1461 (N_1461,N_581,N_412);
nor U1462 (N_1462,N_570,N_42);
or U1463 (N_1463,N_696,N_168);
nand U1464 (N_1464,N_119,N_178);
nor U1465 (N_1465,N_732,N_83);
nand U1466 (N_1466,N_19,N_494);
and U1467 (N_1467,N_238,N_487);
nor U1468 (N_1468,N_637,N_301);
or U1469 (N_1469,N_442,N_692);
nand U1470 (N_1470,N_262,N_547);
nor U1471 (N_1471,N_458,N_384);
nand U1472 (N_1472,N_262,N_302);
nor U1473 (N_1473,N_484,N_734);
nor U1474 (N_1474,N_500,N_156);
nor U1475 (N_1475,N_314,N_103);
or U1476 (N_1476,N_506,N_660);
and U1477 (N_1477,N_573,N_690);
nand U1478 (N_1478,N_608,N_605);
and U1479 (N_1479,N_114,N_553);
nand U1480 (N_1480,N_637,N_201);
nand U1481 (N_1481,N_554,N_238);
and U1482 (N_1482,N_84,N_732);
nand U1483 (N_1483,N_334,N_205);
nand U1484 (N_1484,N_28,N_167);
or U1485 (N_1485,N_152,N_540);
nand U1486 (N_1486,N_400,N_499);
and U1487 (N_1487,N_601,N_46);
or U1488 (N_1488,N_52,N_611);
nor U1489 (N_1489,N_445,N_599);
xnor U1490 (N_1490,N_58,N_480);
nand U1491 (N_1491,N_89,N_614);
or U1492 (N_1492,N_565,N_545);
nand U1493 (N_1493,N_345,N_741);
or U1494 (N_1494,N_333,N_544);
nor U1495 (N_1495,N_408,N_3);
and U1496 (N_1496,N_94,N_397);
or U1497 (N_1497,N_17,N_322);
and U1498 (N_1498,N_44,N_697);
and U1499 (N_1499,N_569,N_23);
nor U1500 (N_1500,N_1108,N_1359);
xor U1501 (N_1501,N_1229,N_1417);
nand U1502 (N_1502,N_1284,N_1195);
nand U1503 (N_1503,N_1147,N_1049);
nand U1504 (N_1504,N_1498,N_1414);
and U1505 (N_1505,N_1447,N_1007);
or U1506 (N_1506,N_971,N_1222);
nor U1507 (N_1507,N_1300,N_1278);
xnor U1508 (N_1508,N_829,N_757);
xnor U1509 (N_1509,N_1127,N_1403);
nand U1510 (N_1510,N_1443,N_1390);
or U1511 (N_1511,N_873,N_893);
nand U1512 (N_1512,N_1408,N_1382);
nor U1513 (N_1513,N_854,N_855);
and U1514 (N_1514,N_917,N_1436);
nor U1515 (N_1515,N_1177,N_789);
nand U1516 (N_1516,N_1232,N_859);
nor U1517 (N_1517,N_1435,N_751);
nor U1518 (N_1518,N_1226,N_1404);
and U1519 (N_1519,N_1144,N_1225);
and U1520 (N_1520,N_1441,N_1055);
and U1521 (N_1521,N_1066,N_883);
xor U1522 (N_1522,N_1203,N_1387);
and U1523 (N_1523,N_1161,N_1175);
and U1524 (N_1524,N_1332,N_1352);
or U1525 (N_1525,N_1351,N_1117);
nor U1526 (N_1526,N_1155,N_1385);
and U1527 (N_1527,N_812,N_1025);
nand U1528 (N_1528,N_979,N_759);
and U1529 (N_1529,N_1228,N_1191);
nand U1530 (N_1530,N_1247,N_841);
xnor U1531 (N_1531,N_913,N_922);
nand U1532 (N_1532,N_967,N_1032);
or U1533 (N_1533,N_1085,N_1327);
or U1534 (N_1534,N_1143,N_761);
nand U1535 (N_1535,N_1268,N_1423);
xor U1536 (N_1536,N_1180,N_828);
and U1537 (N_1537,N_765,N_930);
and U1538 (N_1538,N_823,N_1343);
xnor U1539 (N_1539,N_1245,N_991);
nand U1540 (N_1540,N_1335,N_1131);
xnor U1541 (N_1541,N_881,N_1084);
or U1542 (N_1542,N_1054,N_1021);
and U1543 (N_1543,N_908,N_1286);
or U1544 (N_1544,N_997,N_1040);
or U1545 (N_1545,N_1019,N_1028);
or U1546 (N_1546,N_1453,N_1038);
nand U1547 (N_1547,N_1484,N_1016);
nor U1548 (N_1548,N_1336,N_1035);
or U1549 (N_1549,N_996,N_752);
and U1550 (N_1550,N_1018,N_1223);
or U1551 (N_1551,N_1187,N_766);
or U1552 (N_1552,N_1160,N_1276);
or U1553 (N_1553,N_886,N_969);
or U1554 (N_1554,N_1383,N_1046);
or U1555 (N_1555,N_974,N_1063);
nor U1556 (N_1556,N_904,N_846);
xnor U1557 (N_1557,N_1444,N_1000);
nor U1558 (N_1558,N_1365,N_853);
xnor U1559 (N_1559,N_1120,N_1059);
xnor U1560 (N_1560,N_1213,N_1128);
and U1561 (N_1561,N_1297,N_775);
or U1562 (N_1562,N_965,N_921);
nand U1563 (N_1563,N_1197,N_1350);
nor U1564 (N_1564,N_1463,N_1289);
nor U1565 (N_1565,N_815,N_756);
nor U1566 (N_1566,N_1004,N_870);
or U1567 (N_1567,N_1330,N_760);
nor U1568 (N_1568,N_1397,N_882);
or U1569 (N_1569,N_803,N_796);
nor U1570 (N_1570,N_1246,N_1061);
and U1571 (N_1571,N_1031,N_1266);
nand U1572 (N_1572,N_1317,N_1409);
nand U1573 (N_1573,N_1281,N_903);
nand U1574 (N_1574,N_1265,N_1009);
nand U1575 (N_1575,N_1053,N_1258);
and U1576 (N_1576,N_1416,N_982);
nand U1577 (N_1577,N_1043,N_1202);
and U1578 (N_1578,N_1458,N_1377);
nor U1579 (N_1579,N_1366,N_1426);
and U1580 (N_1580,N_1182,N_1311);
and U1581 (N_1581,N_1275,N_1439);
or U1582 (N_1582,N_1233,N_1176);
nor U1583 (N_1583,N_1087,N_1342);
nor U1584 (N_1584,N_915,N_1036);
or U1585 (N_1585,N_1451,N_1494);
nand U1586 (N_1586,N_1427,N_1491);
nor U1587 (N_1587,N_990,N_767);
nand U1588 (N_1588,N_980,N_1483);
nand U1589 (N_1589,N_1138,N_1062);
and U1590 (N_1590,N_1271,N_1430);
and U1591 (N_1591,N_811,N_1140);
and U1592 (N_1592,N_940,N_1077);
nor U1593 (N_1593,N_912,N_1486);
nor U1594 (N_1594,N_1130,N_1279);
or U1595 (N_1595,N_1367,N_1369);
or U1596 (N_1596,N_1238,N_959);
and U1597 (N_1597,N_1466,N_1081);
or U1598 (N_1598,N_1292,N_1163);
xor U1599 (N_1599,N_1401,N_880);
nand U1600 (N_1600,N_852,N_1209);
xnor U1601 (N_1601,N_1211,N_1384);
nand U1602 (N_1602,N_1290,N_1132);
nor U1603 (N_1603,N_1448,N_957);
and U1604 (N_1604,N_929,N_833);
nand U1605 (N_1605,N_1296,N_1406);
and U1606 (N_1606,N_1212,N_1329);
xnor U1607 (N_1607,N_953,N_1378);
or U1608 (N_1608,N_934,N_1099);
nor U1609 (N_1609,N_1188,N_1314);
and U1610 (N_1610,N_1250,N_1456);
nand U1611 (N_1611,N_1142,N_985);
nand U1612 (N_1612,N_1261,N_1418);
or U1613 (N_1613,N_1370,N_1159);
and U1614 (N_1614,N_1057,N_1496);
and U1615 (N_1615,N_1026,N_1361);
nand U1616 (N_1616,N_1264,N_814);
and U1617 (N_1617,N_866,N_1255);
or U1618 (N_1618,N_1432,N_801);
nand U1619 (N_1619,N_1005,N_1259);
nand U1620 (N_1620,N_1368,N_1217);
nor U1621 (N_1621,N_1395,N_1050);
or U1622 (N_1622,N_1339,N_1052);
xor U1623 (N_1623,N_869,N_1241);
and U1624 (N_1624,N_1092,N_879);
nor U1625 (N_1625,N_827,N_781);
or U1626 (N_1626,N_1413,N_1400);
and U1627 (N_1627,N_951,N_1179);
nand U1628 (N_1628,N_1012,N_835);
xor U1629 (N_1629,N_863,N_1164);
or U1630 (N_1630,N_821,N_1149);
nand U1631 (N_1631,N_993,N_1193);
nand U1632 (N_1632,N_1208,N_1481);
nor U1633 (N_1633,N_810,N_1355);
nand U1634 (N_1634,N_837,N_946);
or U1635 (N_1635,N_1080,N_864);
xnor U1636 (N_1636,N_887,N_1362);
or U1637 (N_1637,N_1454,N_1473);
or U1638 (N_1638,N_1151,N_1316);
nand U1639 (N_1639,N_1433,N_795);
nand U1640 (N_1640,N_1106,N_1381);
or U1641 (N_1641,N_1048,N_822);
or U1642 (N_1642,N_1148,N_1083);
nand U1643 (N_1643,N_1319,N_1374);
nor U1644 (N_1644,N_755,N_1020);
xor U1645 (N_1645,N_1499,N_895);
and U1646 (N_1646,N_1474,N_1033);
or U1647 (N_1647,N_889,N_1415);
and U1648 (N_1648,N_876,N_857);
or U1649 (N_1649,N_1285,N_794);
xnor U1650 (N_1650,N_1396,N_1137);
nand U1651 (N_1651,N_1462,N_1065);
nand U1652 (N_1652,N_1119,N_830);
nand U1653 (N_1653,N_955,N_1218);
nor U1654 (N_1654,N_1023,N_954);
nand U1655 (N_1655,N_1328,N_1125);
or U1656 (N_1656,N_1464,N_1412);
xor U1657 (N_1657,N_1006,N_952);
or U1658 (N_1658,N_1470,N_1227);
nand U1659 (N_1659,N_1162,N_1267);
nor U1660 (N_1660,N_1360,N_1001);
nor U1661 (N_1661,N_1394,N_1123);
and U1662 (N_1662,N_806,N_831);
nand U1663 (N_1663,N_1158,N_950);
nand U1664 (N_1664,N_1206,N_838);
and U1665 (N_1665,N_1477,N_798);
and U1666 (N_1666,N_1114,N_1402);
or U1667 (N_1667,N_804,N_832);
or U1668 (N_1668,N_941,N_1022);
nand U1669 (N_1669,N_914,N_1098);
nand U1670 (N_1670,N_1465,N_1221);
or U1671 (N_1671,N_1141,N_768);
or U1672 (N_1672,N_793,N_839);
nand U1673 (N_1673,N_981,N_897);
nor U1674 (N_1674,N_964,N_1455);
nor U1675 (N_1675,N_1488,N_1434);
nor U1676 (N_1676,N_843,N_858);
or U1677 (N_1677,N_1134,N_860);
nand U1678 (N_1678,N_1420,N_1215);
and U1679 (N_1679,N_824,N_1105);
or U1680 (N_1680,N_1078,N_1089);
xor U1681 (N_1681,N_1112,N_896);
and U1682 (N_1682,N_1306,N_1253);
and U1683 (N_1683,N_1174,N_1060);
nand U1684 (N_1684,N_1216,N_1460);
nor U1685 (N_1685,N_1251,N_972);
xnor U1686 (N_1686,N_1459,N_1356);
nor U1687 (N_1687,N_999,N_1047);
or U1688 (N_1688,N_1450,N_773);
nor U1689 (N_1689,N_1091,N_1344);
nand U1690 (N_1690,N_1170,N_1318);
nand U1691 (N_1691,N_845,N_1152);
or U1692 (N_1692,N_984,N_1126);
and U1693 (N_1693,N_1347,N_790);
nor U1694 (N_1694,N_1452,N_762);
nor U1695 (N_1695,N_1257,N_1354);
xnor U1696 (N_1696,N_1348,N_1039);
xnor U1697 (N_1697,N_1479,N_935);
nand U1698 (N_1698,N_1239,N_1219);
and U1699 (N_1699,N_1011,N_1097);
or U1700 (N_1700,N_1118,N_1301);
or U1701 (N_1701,N_1373,N_944);
or U1702 (N_1702,N_792,N_1349);
nor U1703 (N_1703,N_1094,N_840);
xnor U1704 (N_1704,N_1024,N_1399);
and U1705 (N_1705,N_1234,N_899);
nand U1706 (N_1706,N_764,N_937);
or U1707 (N_1707,N_894,N_888);
and U1708 (N_1708,N_868,N_1272);
nand U1709 (N_1709,N_1186,N_1185);
and U1710 (N_1710,N_947,N_1034);
nor U1711 (N_1711,N_1480,N_1371);
or U1712 (N_1712,N_783,N_1201);
nor U1713 (N_1713,N_1475,N_1076);
nand U1714 (N_1714,N_1469,N_1243);
nor U1715 (N_1715,N_1015,N_1291);
or U1716 (N_1716,N_797,N_1424);
nor U1717 (N_1717,N_891,N_1437);
and U1718 (N_1718,N_1472,N_1493);
nor U1719 (N_1719,N_1421,N_1178);
nand U1720 (N_1720,N_1240,N_817);
or U1721 (N_1721,N_834,N_774);
nand U1722 (N_1722,N_1485,N_776);
nor U1723 (N_1723,N_1096,N_1150);
or U1724 (N_1724,N_849,N_1189);
or U1725 (N_1725,N_1045,N_1056);
xnor U1726 (N_1726,N_1183,N_1461);
nor U1727 (N_1727,N_1334,N_1072);
or U1728 (N_1728,N_1487,N_780);
nor U1729 (N_1729,N_928,N_1192);
and U1730 (N_1730,N_1064,N_1313);
nand U1731 (N_1731,N_966,N_963);
or U1732 (N_1732,N_1282,N_987);
and U1733 (N_1733,N_1337,N_1376);
or U1734 (N_1734,N_753,N_1357);
xnor U1735 (N_1735,N_1041,N_1224);
and U1736 (N_1736,N_1405,N_1398);
and U1737 (N_1737,N_1101,N_1363);
and U1738 (N_1738,N_784,N_1214);
nand U1739 (N_1739,N_1322,N_973);
and U1740 (N_1740,N_958,N_1104);
or U1741 (N_1741,N_1478,N_1393);
and U1742 (N_1742,N_1492,N_871);
nor U1743 (N_1743,N_1299,N_754);
and U1744 (N_1744,N_1260,N_885);
or U1745 (N_1745,N_1333,N_1116);
nand U1746 (N_1746,N_1111,N_992);
nor U1747 (N_1747,N_1070,N_918);
nor U1748 (N_1748,N_1310,N_1037);
nand U1749 (N_1749,N_909,N_1497);
and U1750 (N_1750,N_1093,N_1490);
xnor U1751 (N_1751,N_1236,N_1321);
nand U1752 (N_1752,N_779,N_1230);
or U1753 (N_1753,N_924,N_1489);
or U1754 (N_1754,N_902,N_1113);
nand U1755 (N_1755,N_1331,N_936);
and U1756 (N_1756,N_1220,N_1102);
or U1757 (N_1757,N_1156,N_1139);
nor U1758 (N_1758,N_923,N_968);
xor U1759 (N_1759,N_1014,N_1068);
and U1760 (N_1760,N_1157,N_836);
nand U1761 (N_1761,N_1017,N_1090);
or U1762 (N_1762,N_799,N_1495);
or U1763 (N_1763,N_1476,N_1121);
nand U1764 (N_1764,N_1305,N_945);
nand U1765 (N_1765,N_1172,N_983);
or U1766 (N_1766,N_1030,N_1440);
or U1767 (N_1767,N_1198,N_1309);
or U1768 (N_1768,N_842,N_1165);
and U1769 (N_1769,N_809,N_916);
nand U1770 (N_1770,N_1422,N_1302);
and U1771 (N_1771,N_1235,N_942);
nor U1772 (N_1772,N_1287,N_1312);
or U1773 (N_1773,N_1027,N_1295);
nor U1774 (N_1774,N_986,N_1388);
or U1775 (N_1775,N_1358,N_816);
xor U1776 (N_1776,N_1341,N_1181);
nor U1777 (N_1777,N_1073,N_1204);
and U1778 (N_1778,N_1058,N_1129);
or U1779 (N_1779,N_1184,N_800);
or U1780 (N_1780,N_847,N_1283);
nand U1781 (N_1781,N_975,N_1325);
and U1782 (N_1782,N_884,N_905);
nor U1783 (N_1783,N_1392,N_1075);
and U1784 (N_1784,N_802,N_785);
nor U1785 (N_1785,N_1100,N_813);
xnor U1786 (N_1786,N_1168,N_1069);
nor U1787 (N_1787,N_805,N_808);
nor U1788 (N_1788,N_1280,N_970);
xnor U1789 (N_1789,N_1109,N_1298);
nand U1790 (N_1790,N_920,N_875);
xnor U1791 (N_1791,N_851,N_1110);
nor U1792 (N_1792,N_807,N_1242);
nor U1793 (N_1793,N_1379,N_786);
nor U1794 (N_1794,N_1210,N_943);
nand U1795 (N_1795,N_925,N_1438);
or U1796 (N_1796,N_791,N_1372);
and U1797 (N_1797,N_1274,N_932);
nand U1798 (N_1798,N_1107,N_898);
or U1799 (N_1799,N_1375,N_1256);
nor U1800 (N_1800,N_1169,N_1231);
nand U1801 (N_1801,N_1194,N_1145);
nor U1802 (N_1802,N_877,N_938);
nor U1803 (N_1803,N_1449,N_919);
xnor U1804 (N_1804,N_1304,N_892);
and U1805 (N_1805,N_1294,N_1082);
and U1806 (N_1806,N_770,N_862);
nor U1807 (N_1807,N_911,N_856);
xor U1808 (N_1808,N_1095,N_1308);
or U1809 (N_1809,N_1442,N_989);
and U1810 (N_1810,N_1467,N_1252);
and U1811 (N_1811,N_1003,N_926);
nor U1812 (N_1812,N_1153,N_1079);
or U1813 (N_1813,N_1445,N_1270);
nor U1814 (N_1814,N_874,N_1205);
nand U1815 (N_1815,N_865,N_1407);
nor U1816 (N_1816,N_1067,N_1244);
and U1817 (N_1817,N_976,N_988);
nand U1818 (N_1818,N_1171,N_998);
nor U1819 (N_1819,N_994,N_1471);
and U1820 (N_1820,N_1386,N_1273);
or U1821 (N_1821,N_1200,N_948);
and U1822 (N_1822,N_1338,N_1346);
and U1823 (N_1823,N_1410,N_1136);
nor U1824 (N_1824,N_1074,N_900);
nand U1825 (N_1825,N_1269,N_788);
nand U1826 (N_1826,N_750,N_1008);
or U1827 (N_1827,N_758,N_933);
nand U1828 (N_1828,N_818,N_1326);
and U1829 (N_1829,N_1103,N_1446);
nor U1830 (N_1830,N_778,N_956);
xnor U1831 (N_1831,N_1196,N_850);
and U1832 (N_1832,N_1389,N_771);
xnor U1833 (N_1833,N_1166,N_1315);
nand U1834 (N_1834,N_1277,N_819);
and U1835 (N_1835,N_962,N_861);
nor U1836 (N_1836,N_1002,N_977);
or U1837 (N_1837,N_1323,N_1425);
nand U1838 (N_1838,N_960,N_1115);
and U1839 (N_1839,N_1320,N_1124);
or U1840 (N_1840,N_1345,N_1364);
or U1841 (N_1841,N_1482,N_1431);
and U1842 (N_1842,N_1262,N_787);
or U1843 (N_1843,N_1340,N_769);
or U1844 (N_1844,N_878,N_1307);
and U1845 (N_1845,N_1029,N_907);
nand U1846 (N_1846,N_867,N_777);
and U1847 (N_1847,N_1263,N_1088);
nand U1848 (N_1848,N_1122,N_1051);
nand U1849 (N_1849,N_1468,N_772);
and U1850 (N_1850,N_1428,N_1248);
nor U1851 (N_1851,N_1190,N_1199);
and U1852 (N_1852,N_949,N_1324);
nand U1853 (N_1853,N_1411,N_1154);
and U1854 (N_1854,N_931,N_820);
and U1855 (N_1855,N_848,N_782);
nor U1856 (N_1856,N_939,N_890);
and U1857 (N_1857,N_1380,N_1167);
nand U1858 (N_1858,N_1457,N_910);
nor U1859 (N_1859,N_825,N_1207);
nor U1860 (N_1860,N_1419,N_927);
and U1861 (N_1861,N_1086,N_1042);
xnor U1862 (N_1862,N_1173,N_1293);
xnor U1863 (N_1863,N_1146,N_906);
xor U1864 (N_1864,N_844,N_763);
xor U1865 (N_1865,N_1044,N_1353);
nand U1866 (N_1866,N_1249,N_1288);
nand U1867 (N_1867,N_1254,N_1133);
nor U1868 (N_1868,N_1013,N_961);
nand U1869 (N_1869,N_1135,N_1429);
nand U1870 (N_1870,N_1010,N_1237);
and U1871 (N_1871,N_872,N_901);
and U1872 (N_1872,N_826,N_1391);
nand U1873 (N_1873,N_978,N_995);
xnor U1874 (N_1874,N_1071,N_1303);
nor U1875 (N_1875,N_1338,N_754);
or U1876 (N_1876,N_983,N_1335);
and U1877 (N_1877,N_1449,N_900);
xor U1878 (N_1878,N_1313,N_1299);
nor U1879 (N_1879,N_896,N_1053);
and U1880 (N_1880,N_935,N_1208);
nor U1881 (N_1881,N_771,N_1131);
nand U1882 (N_1882,N_1146,N_1338);
xor U1883 (N_1883,N_902,N_1148);
nor U1884 (N_1884,N_1341,N_1120);
nor U1885 (N_1885,N_1494,N_1267);
nor U1886 (N_1886,N_1323,N_764);
nor U1887 (N_1887,N_1292,N_920);
nor U1888 (N_1888,N_1092,N_992);
or U1889 (N_1889,N_1288,N_901);
nand U1890 (N_1890,N_988,N_1231);
nor U1891 (N_1891,N_952,N_1388);
nand U1892 (N_1892,N_1273,N_1293);
xnor U1893 (N_1893,N_1093,N_1310);
nor U1894 (N_1894,N_960,N_1272);
xnor U1895 (N_1895,N_837,N_1358);
and U1896 (N_1896,N_1199,N_1214);
and U1897 (N_1897,N_984,N_1369);
nor U1898 (N_1898,N_1413,N_846);
nand U1899 (N_1899,N_1107,N_962);
nor U1900 (N_1900,N_1157,N_1335);
and U1901 (N_1901,N_1125,N_1322);
or U1902 (N_1902,N_1494,N_1125);
and U1903 (N_1903,N_936,N_1290);
or U1904 (N_1904,N_757,N_1043);
or U1905 (N_1905,N_856,N_819);
and U1906 (N_1906,N_785,N_1451);
or U1907 (N_1907,N_1213,N_1129);
or U1908 (N_1908,N_890,N_1148);
nor U1909 (N_1909,N_1388,N_1112);
nor U1910 (N_1910,N_1110,N_1238);
and U1911 (N_1911,N_967,N_1232);
xor U1912 (N_1912,N_1471,N_1161);
nand U1913 (N_1913,N_1303,N_851);
nor U1914 (N_1914,N_919,N_932);
xor U1915 (N_1915,N_1132,N_1243);
nor U1916 (N_1916,N_949,N_871);
or U1917 (N_1917,N_949,N_783);
xnor U1918 (N_1918,N_1468,N_773);
and U1919 (N_1919,N_1347,N_1481);
nor U1920 (N_1920,N_756,N_1357);
xnor U1921 (N_1921,N_763,N_981);
nor U1922 (N_1922,N_1400,N_1060);
nor U1923 (N_1923,N_753,N_1058);
and U1924 (N_1924,N_1139,N_1367);
or U1925 (N_1925,N_1160,N_1142);
and U1926 (N_1926,N_1323,N_758);
xnor U1927 (N_1927,N_1128,N_902);
xnor U1928 (N_1928,N_1280,N_968);
and U1929 (N_1929,N_1439,N_1250);
nand U1930 (N_1930,N_1455,N_1431);
nor U1931 (N_1931,N_1152,N_1230);
nor U1932 (N_1932,N_1113,N_1066);
nor U1933 (N_1933,N_1005,N_878);
nor U1934 (N_1934,N_964,N_930);
or U1935 (N_1935,N_1161,N_1247);
or U1936 (N_1936,N_1049,N_1166);
or U1937 (N_1937,N_1100,N_1287);
nor U1938 (N_1938,N_1263,N_1141);
nor U1939 (N_1939,N_1181,N_1423);
nor U1940 (N_1940,N_991,N_1162);
or U1941 (N_1941,N_1131,N_1433);
and U1942 (N_1942,N_923,N_1006);
or U1943 (N_1943,N_1101,N_1400);
nand U1944 (N_1944,N_1339,N_1279);
and U1945 (N_1945,N_986,N_1098);
or U1946 (N_1946,N_1280,N_1249);
or U1947 (N_1947,N_1284,N_1084);
and U1948 (N_1948,N_777,N_1408);
nand U1949 (N_1949,N_1183,N_1381);
and U1950 (N_1950,N_1199,N_867);
or U1951 (N_1951,N_1492,N_1108);
and U1952 (N_1952,N_1240,N_1376);
nor U1953 (N_1953,N_1459,N_1074);
nor U1954 (N_1954,N_875,N_1154);
nor U1955 (N_1955,N_1409,N_853);
nand U1956 (N_1956,N_1194,N_843);
and U1957 (N_1957,N_1406,N_997);
and U1958 (N_1958,N_1175,N_1418);
nor U1959 (N_1959,N_1112,N_880);
nor U1960 (N_1960,N_1096,N_1170);
nor U1961 (N_1961,N_879,N_804);
nor U1962 (N_1962,N_1233,N_1448);
and U1963 (N_1963,N_770,N_1366);
nand U1964 (N_1964,N_1275,N_1229);
or U1965 (N_1965,N_1153,N_989);
nand U1966 (N_1966,N_1256,N_1233);
or U1967 (N_1967,N_1344,N_817);
or U1968 (N_1968,N_1202,N_1438);
nor U1969 (N_1969,N_822,N_864);
nor U1970 (N_1970,N_900,N_1067);
nand U1971 (N_1971,N_1033,N_1405);
nor U1972 (N_1972,N_1158,N_1038);
nand U1973 (N_1973,N_1326,N_1052);
or U1974 (N_1974,N_868,N_1106);
and U1975 (N_1975,N_1498,N_815);
nor U1976 (N_1976,N_1457,N_1033);
and U1977 (N_1977,N_1315,N_1171);
or U1978 (N_1978,N_1310,N_1209);
nand U1979 (N_1979,N_911,N_1028);
nand U1980 (N_1980,N_797,N_1113);
nor U1981 (N_1981,N_1166,N_1088);
xnor U1982 (N_1982,N_1344,N_1079);
nand U1983 (N_1983,N_1299,N_1328);
nand U1984 (N_1984,N_1180,N_1449);
xor U1985 (N_1985,N_1259,N_879);
and U1986 (N_1986,N_1441,N_1398);
or U1987 (N_1987,N_1323,N_1184);
nor U1988 (N_1988,N_1010,N_1306);
nand U1989 (N_1989,N_996,N_1110);
nor U1990 (N_1990,N_1330,N_849);
nand U1991 (N_1991,N_878,N_1317);
and U1992 (N_1992,N_850,N_1235);
nand U1993 (N_1993,N_1448,N_761);
nor U1994 (N_1994,N_1423,N_1397);
or U1995 (N_1995,N_783,N_1306);
or U1996 (N_1996,N_1486,N_975);
nand U1997 (N_1997,N_1138,N_1212);
or U1998 (N_1998,N_826,N_1043);
and U1999 (N_1999,N_1404,N_1339);
nor U2000 (N_2000,N_873,N_1407);
nor U2001 (N_2001,N_1083,N_1210);
xor U2002 (N_2002,N_1325,N_1459);
xnor U2003 (N_2003,N_1477,N_1070);
nor U2004 (N_2004,N_1193,N_962);
nor U2005 (N_2005,N_1071,N_1259);
or U2006 (N_2006,N_1270,N_1033);
nand U2007 (N_2007,N_1239,N_990);
or U2008 (N_2008,N_769,N_920);
nand U2009 (N_2009,N_822,N_944);
nand U2010 (N_2010,N_1142,N_1272);
and U2011 (N_2011,N_928,N_1337);
nand U2012 (N_2012,N_822,N_1383);
and U2013 (N_2013,N_813,N_978);
nand U2014 (N_2014,N_802,N_1074);
nand U2015 (N_2015,N_1304,N_1225);
or U2016 (N_2016,N_795,N_1161);
nor U2017 (N_2017,N_938,N_1404);
nand U2018 (N_2018,N_1088,N_1331);
nor U2019 (N_2019,N_1130,N_800);
xor U2020 (N_2020,N_881,N_1125);
nor U2021 (N_2021,N_1000,N_1309);
and U2022 (N_2022,N_1023,N_1478);
nor U2023 (N_2023,N_1377,N_1376);
nor U2024 (N_2024,N_1265,N_911);
nand U2025 (N_2025,N_1400,N_1387);
nand U2026 (N_2026,N_1079,N_801);
and U2027 (N_2027,N_1181,N_1120);
nor U2028 (N_2028,N_978,N_878);
and U2029 (N_2029,N_1113,N_897);
or U2030 (N_2030,N_910,N_915);
xnor U2031 (N_2031,N_981,N_1233);
nor U2032 (N_2032,N_1365,N_972);
nand U2033 (N_2033,N_887,N_849);
xnor U2034 (N_2034,N_1328,N_1492);
and U2035 (N_2035,N_1483,N_828);
or U2036 (N_2036,N_1058,N_990);
nor U2037 (N_2037,N_1359,N_1033);
nand U2038 (N_2038,N_801,N_885);
or U2039 (N_2039,N_1301,N_1308);
nand U2040 (N_2040,N_974,N_1135);
nand U2041 (N_2041,N_1444,N_754);
nor U2042 (N_2042,N_1284,N_1200);
xor U2043 (N_2043,N_1172,N_787);
and U2044 (N_2044,N_1139,N_1345);
nand U2045 (N_2045,N_909,N_962);
nand U2046 (N_2046,N_1114,N_979);
nor U2047 (N_2047,N_1323,N_1182);
nor U2048 (N_2048,N_1362,N_786);
or U2049 (N_2049,N_1442,N_1078);
and U2050 (N_2050,N_783,N_1065);
and U2051 (N_2051,N_1174,N_822);
nor U2052 (N_2052,N_1342,N_1128);
or U2053 (N_2053,N_1012,N_1215);
nand U2054 (N_2054,N_973,N_919);
nor U2055 (N_2055,N_1485,N_891);
and U2056 (N_2056,N_1042,N_1292);
xnor U2057 (N_2057,N_1411,N_1133);
nand U2058 (N_2058,N_1007,N_1066);
and U2059 (N_2059,N_1187,N_1483);
and U2060 (N_2060,N_1279,N_1223);
nand U2061 (N_2061,N_963,N_852);
or U2062 (N_2062,N_913,N_757);
and U2063 (N_2063,N_1475,N_1491);
nor U2064 (N_2064,N_1443,N_1111);
nor U2065 (N_2065,N_1154,N_847);
nor U2066 (N_2066,N_1081,N_1467);
nor U2067 (N_2067,N_886,N_1101);
and U2068 (N_2068,N_1179,N_757);
and U2069 (N_2069,N_1000,N_1138);
nand U2070 (N_2070,N_1301,N_1029);
and U2071 (N_2071,N_1249,N_788);
or U2072 (N_2072,N_837,N_768);
or U2073 (N_2073,N_990,N_1171);
or U2074 (N_2074,N_889,N_882);
nor U2075 (N_2075,N_1295,N_1111);
nand U2076 (N_2076,N_1232,N_937);
and U2077 (N_2077,N_1364,N_1373);
or U2078 (N_2078,N_1127,N_1341);
and U2079 (N_2079,N_896,N_963);
and U2080 (N_2080,N_985,N_1106);
nand U2081 (N_2081,N_1233,N_816);
xor U2082 (N_2082,N_1018,N_796);
or U2083 (N_2083,N_1189,N_954);
or U2084 (N_2084,N_768,N_1281);
and U2085 (N_2085,N_1280,N_1166);
or U2086 (N_2086,N_904,N_1247);
or U2087 (N_2087,N_1401,N_1228);
xor U2088 (N_2088,N_869,N_1082);
nor U2089 (N_2089,N_1349,N_1332);
nand U2090 (N_2090,N_1466,N_1456);
nor U2091 (N_2091,N_1497,N_1195);
and U2092 (N_2092,N_921,N_1083);
nor U2093 (N_2093,N_1248,N_1085);
or U2094 (N_2094,N_1088,N_818);
nor U2095 (N_2095,N_1491,N_1183);
nand U2096 (N_2096,N_881,N_836);
nand U2097 (N_2097,N_1196,N_813);
and U2098 (N_2098,N_1017,N_1439);
and U2099 (N_2099,N_1418,N_1479);
nand U2100 (N_2100,N_989,N_824);
nand U2101 (N_2101,N_1329,N_1422);
nor U2102 (N_2102,N_1316,N_1317);
nand U2103 (N_2103,N_1126,N_800);
or U2104 (N_2104,N_1161,N_1296);
xnor U2105 (N_2105,N_928,N_1467);
nand U2106 (N_2106,N_1176,N_1083);
xnor U2107 (N_2107,N_1142,N_811);
nor U2108 (N_2108,N_775,N_1133);
nor U2109 (N_2109,N_981,N_1078);
nor U2110 (N_2110,N_1010,N_1158);
xor U2111 (N_2111,N_781,N_1233);
nor U2112 (N_2112,N_953,N_969);
nand U2113 (N_2113,N_1133,N_874);
or U2114 (N_2114,N_1015,N_1221);
xor U2115 (N_2115,N_1368,N_952);
and U2116 (N_2116,N_1128,N_1122);
nand U2117 (N_2117,N_1053,N_769);
nor U2118 (N_2118,N_1329,N_914);
or U2119 (N_2119,N_1411,N_1183);
nand U2120 (N_2120,N_819,N_964);
xnor U2121 (N_2121,N_943,N_914);
xor U2122 (N_2122,N_1235,N_1160);
nand U2123 (N_2123,N_1397,N_955);
or U2124 (N_2124,N_1179,N_1263);
and U2125 (N_2125,N_1183,N_918);
nand U2126 (N_2126,N_881,N_1440);
and U2127 (N_2127,N_882,N_833);
nor U2128 (N_2128,N_1374,N_1144);
or U2129 (N_2129,N_893,N_768);
nand U2130 (N_2130,N_869,N_1088);
nand U2131 (N_2131,N_1330,N_1217);
nor U2132 (N_2132,N_870,N_957);
or U2133 (N_2133,N_884,N_1015);
or U2134 (N_2134,N_1129,N_1248);
xor U2135 (N_2135,N_1047,N_1098);
and U2136 (N_2136,N_964,N_1375);
or U2137 (N_2137,N_1422,N_1177);
nand U2138 (N_2138,N_1466,N_854);
and U2139 (N_2139,N_1133,N_928);
nand U2140 (N_2140,N_1497,N_1379);
and U2141 (N_2141,N_978,N_1347);
nand U2142 (N_2142,N_1425,N_1348);
nor U2143 (N_2143,N_1077,N_1330);
nand U2144 (N_2144,N_893,N_818);
nand U2145 (N_2145,N_1277,N_1229);
and U2146 (N_2146,N_1131,N_1458);
nor U2147 (N_2147,N_859,N_1089);
or U2148 (N_2148,N_1131,N_1403);
nor U2149 (N_2149,N_1466,N_797);
or U2150 (N_2150,N_757,N_779);
xnor U2151 (N_2151,N_919,N_1377);
nand U2152 (N_2152,N_1122,N_1315);
nand U2153 (N_2153,N_771,N_1083);
or U2154 (N_2154,N_753,N_1308);
nand U2155 (N_2155,N_1078,N_1476);
and U2156 (N_2156,N_919,N_945);
xor U2157 (N_2157,N_917,N_1169);
nand U2158 (N_2158,N_753,N_1338);
nor U2159 (N_2159,N_840,N_1006);
or U2160 (N_2160,N_1031,N_1476);
or U2161 (N_2161,N_865,N_1106);
or U2162 (N_2162,N_1323,N_1007);
and U2163 (N_2163,N_827,N_1197);
and U2164 (N_2164,N_1045,N_1119);
or U2165 (N_2165,N_1228,N_941);
nor U2166 (N_2166,N_1487,N_1138);
nand U2167 (N_2167,N_827,N_964);
or U2168 (N_2168,N_1402,N_889);
and U2169 (N_2169,N_944,N_761);
nor U2170 (N_2170,N_892,N_1093);
nand U2171 (N_2171,N_987,N_1279);
or U2172 (N_2172,N_1330,N_952);
nor U2173 (N_2173,N_1349,N_1265);
nor U2174 (N_2174,N_939,N_1110);
nor U2175 (N_2175,N_1062,N_1254);
or U2176 (N_2176,N_991,N_959);
nor U2177 (N_2177,N_1349,N_1248);
nand U2178 (N_2178,N_1453,N_1239);
nand U2179 (N_2179,N_1452,N_926);
or U2180 (N_2180,N_1049,N_1246);
and U2181 (N_2181,N_1210,N_889);
and U2182 (N_2182,N_833,N_823);
or U2183 (N_2183,N_1040,N_1006);
or U2184 (N_2184,N_1271,N_760);
and U2185 (N_2185,N_1360,N_1209);
and U2186 (N_2186,N_968,N_802);
or U2187 (N_2187,N_986,N_1118);
xnor U2188 (N_2188,N_1482,N_947);
nand U2189 (N_2189,N_1344,N_1167);
and U2190 (N_2190,N_944,N_1346);
nand U2191 (N_2191,N_1115,N_1474);
or U2192 (N_2192,N_1411,N_755);
nand U2193 (N_2193,N_1020,N_786);
nand U2194 (N_2194,N_844,N_1109);
nor U2195 (N_2195,N_1311,N_1233);
nand U2196 (N_2196,N_990,N_1281);
nand U2197 (N_2197,N_859,N_757);
and U2198 (N_2198,N_770,N_1110);
or U2199 (N_2199,N_1017,N_1318);
xor U2200 (N_2200,N_802,N_845);
and U2201 (N_2201,N_1431,N_1163);
and U2202 (N_2202,N_1273,N_1442);
or U2203 (N_2203,N_1291,N_954);
nor U2204 (N_2204,N_890,N_1410);
and U2205 (N_2205,N_794,N_1151);
xnor U2206 (N_2206,N_1167,N_1234);
and U2207 (N_2207,N_771,N_1070);
nor U2208 (N_2208,N_1420,N_1307);
or U2209 (N_2209,N_881,N_1137);
nor U2210 (N_2210,N_1405,N_1480);
nand U2211 (N_2211,N_883,N_775);
nor U2212 (N_2212,N_1218,N_1151);
nand U2213 (N_2213,N_1198,N_1145);
and U2214 (N_2214,N_1392,N_1011);
nor U2215 (N_2215,N_1141,N_1472);
xor U2216 (N_2216,N_1021,N_1181);
or U2217 (N_2217,N_894,N_1472);
or U2218 (N_2218,N_1059,N_1162);
or U2219 (N_2219,N_1020,N_988);
and U2220 (N_2220,N_1480,N_1462);
nor U2221 (N_2221,N_814,N_1370);
xnor U2222 (N_2222,N_1497,N_1348);
nor U2223 (N_2223,N_1140,N_871);
xor U2224 (N_2224,N_1251,N_1324);
nand U2225 (N_2225,N_1319,N_959);
and U2226 (N_2226,N_1298,N_869);
nand U2227 (N_2227,N_1249,N_905);
nand U2228 (N_2228,N_990,N_1167);
or U2229 (N_2229,N_1477,N_1347);
or U2230 (N_2230,N_1147,N_788);
nor U2231 (N_2231,N_1108,N_768);
xor U2232 (N_2232,N_1261,N_1036);
nor U2233 (N_2233,N_1374,N_1256);
nand U2234 (N_2234,N_1003,N_858);
or U2235 (N_2235,N_1322,N_1397);
xor U2236 (N_2236,N_1073,N_1322);
and U2237 (N_2237,N_855,N_1307);
or U2238 (N_2238,N_928,N_863);
nor U2239 (N_2239,N_1441,N_1493);
xor U2240 (N_2240,N_1446,N_1251);
nor U2241 (N_2241,N_1325,N_1494);
or U2242 (N_2242,N_823,N_1144);
nand U2243 (N_2243,N_1028,N_1276);
nor U2244 (N_2244,N_1353,N_1172);
nand U2245 (N_2245,N_1040,N_1377);
nand U2246 (N_2246,N_1033,N_1060);
nand U2247 (N_2247,N_1427,N_1364);
nand U2248 (N_2248,N_958,N_1219);
or U2249 (N_2249,N_1410,N_1420);
nor U2250 (N_2250,N_2154,N_2182);
and U2251 (N_2251,N_1690,N_2017);
and U2252 (N_2252,N_2167,N_1609);
nand U2253 (N_2253,N_1644,N_2223);
and U2254 (N_2254,N_2115,N_1840);
nand U2255 (N_2255,N_2099,N_2245);
or U2256 (N_2256,N_1809,N_1572);
or U2257 (N_2257,N_1676,N_1632);
xnor U2258 (N_2258,N_1942,N_1618);
and U2259 (N_2259,N_1940,N_1501);
nand U2260 (N_2260,N_1815,N_1622);
nand U2261 (N_2261,N_1711,N_1626);
nand U2262 (N_2262,N_1786,N_2180);
nand U2263 (N_2263,N_1691,N_1750);
and U2264 (N_2264,N_2045,N_1989);
and U2265 (N_2265,N_1623,N_1597);
and U2266 (N_2266,N_1850,N_1699);
nand U2267 (N_2267,N_2240,N_2107);
nand U2268 (N_2268,N_1610,N_2094);
nand U2269 (N_2269,N_1566,N_1900);
nand U2270 (N_2270,N_1865,N_1544);
and U2271 (N_2271,N_1895,N_1546);
nand U2272 (N_2272,N_2236,N_2218);
nand U2273 (N_2273,N_2214,N_1617);
or U2274 (N_2274,N_2241,N_1724);
nor U2275 (N_2275,N_1859,N_1558);
or U2276 (N_2276,N_1993,N_2060);
or U2277 (N_2277,N_2119,N_1928);
and U2278 (N_2278,N_2075,N_2000);
and U2279 (N_2279,N_1514,N_1614);
nor U2280 (N_2280,N_1595,N_1528);
nor U2281 (N_2281,N_1885,N_1944);
nor U2282 (N_2282,N_2133,N_1712);
xnor U2283 (N_2283,N_1822,N_2082);
xor U2284 (N_2284,N_1530,N_1896);
and U2285 (N_2285,N_2196,N_1985);
or U2286 (N_2286,N_2063,N_1592);
nor U2287 (N_2287,N_2046,N_1910);
nand U2288 (N_2288,N_1655,N_1639);
nor U2289 (N_2289,N_1607,N_1999);
nand U2290 (N_2290,N_1882,N_2098);
nor U2291 (N_2291,N_1628,N_1955);
nor U2292 (N_2292,N_1567,N_1722);
nor U2293 (N_2293,N_1769,N_1913);
nand U2294 (N_2294,N_1713,N_2132);
and U2295 (N_2295,N_2148,N_2036);
nor U2296 (N_2296,N_1752,N_1917);
and U2297 (N_2297,N_1813,N_1960);
or U2298 (N_2298,N_1744,N_2034);
nand U2299 (N_2299,N_2248,N_2190);
nor U2300 (N_2300,N_1811,N_1666);
nor U2301 (N_2301,N_2104,N_1714);
and U2302 (N_2302,N_1763,N_1727);
and U2303 (N_2303,N_2142,N_1590);
nand U2304 (N_2304,N_1672,N_1562);
nand U2305 (N_2305,N_1877,N_1717);
and U2306 (N_2306,N_1755,N_2249);
nand U2307 (N_2307,N_1604,N_2210);
or U2308 (N_2308,N_2089,N_2065);
nor U2309 (N_2309,N_2175,N_1762);
nor U2310 (N_2310,N_2111,N_1686);
and U2311 (N_2311,N_1677,N_1543);
nand U2312 (N_2312,N_1720,N_1835);
nor U2313 (N_2313,N_2040,N_1511);
and U2314 (N_2314,N_2007,N_2114);
and U2315 (N_2315,N_2155,N_1751);
and U2316 (N_2316,N_1857,N_1862);
or U2317 (N_2317,N_2209,N_1967);
nor U2318 (N_2318,N_2042,N_2021);
or U2319 (N_2319,N_1941,N_2156);
nor U2320 (N_2320,N_1849,N_1779);
or U2321 (N_2321,N_1746,N_1839);
nand U2322 (N_2322,N_1605,N_1943);
nor U2323 (N_2323,N_1971,N_1659);
or U2324 (N_2324,N_2172,N_1848);
nand U2325 (N_2325,N_2074,N_1945);
or U2326 (N_2326,N_1968,N_1707);
nand U2327 (N_2327,N_1826,N_1902);
and U2328 (N_2328,N_2219,N_1654);
or U2329 (N_2329,N_1990,N_2247);
and U2330 (N_2330,N_1545,N_1536);
and U2331 (N_2331,N_2205,N_1551);
nor U2332 (N_2332,N_2211,N_1819);
or U2333 (N_2333,N_2228,N_1656);
nand U2334 (N_2334,N_1787,N_2083);
nand U2335 (N_2335,N_1650,N_1756);
nand U2336 (N_2336,N_1680,N_2105);
and U2337 (N_2337,N_2173,N_2013);
and U2338 (N_2338,N_1963,N_1782);
or U2339 (N_2339,N_2141,N_2121);
xor U2340 (N_2340,N_2020,N_2224);
xnor U2341 (N_2341,N_1828,N_1802);
xnor U2342 (N_2342,N_1919,N_1522);
or U2343 (N_2343,N_1851,N_1532);
nor U2344 (N_2344,N_2055,N_1638);
nand U2345 (N_2345,N_1582,N_1591);
nand U2346 (N_2346,N_2053,N_1585);
nor U2347 (N_2347,N_2203,N_2122);
xor U2348 (N_2348,N_2022,N_1721);
nor U2349 (N_2349,N_2018,N_1773);
nor U2350 (N_2350,N_1784,N_2170);
or U2351 (N_2351,N_1905,N_1998);
nor U2352 (N_2352,N_1705,N_1619);
nand U2353 (N_2353,N_1737,N_1734);
nand U2354 (N_2354,N_1754,N_1994);
xnor U2355 (N_2355,N_1991,N_1886);
or U2356 (N_2356,N_1890,N_1863);
and U2357 (N_2357,N_2226,N_2169);
nor U2358 (N_2358,N_2126,N_2103);
and U2359 (N_2359,N_2143,N_1620);
or U2360 (N_2360,N_2242,N_1892);
xnor U2361 (N_2361,N_1866,N_1858);
and U2362 (N_2362,N_1510,N_2041);
or U2363 (N_2363,N_2109,N_1838);
nor U2364 (N_2364,N_1818,N_1984);
or U2365 (N_2365,N_1631,N_1834);
nor U2366 (N_2366,N_2061,N_1516);
or U2367 (N_2367,N_2072,N_1759);
or U2368 (N_2368,N_1855,N_1580);
or U2369 (N_2369,N_1698,N_1771);
nor U2370 (N_2370,N_2037,N_2177);
nand U2371 (N_2371,N_2120,N_1788);
xnor U2372 (N_2372,N_2071,N_1780);
nor U2373 (N_2373,N_1660,N_1860);
xor U2374 (N_2374,N_2232,N_2052);
and U2375 (N_2375,N_2005,N_1694);
nor U2376 (N_2376,N_2159,N_2207);
nand U2377 (N_2377,N_2220,N_1870);
or U2378 (N_2378,N_1925,N_2163);
or U2379 (N_2379,N_2181,N_1505);
nor U2380 (N_2380,N_1983,N_1869);
nand U2381 (N_2381,N_2160,N_2183);
nand U2382 (N_2382,N_1824,N_2084);
nand U2383 (N_2383,N_1789,N_2047);
or U2384 (N_2384,N_2006,N_1775);
nand U2385 (N_2385,N_1757,N_2176);
or U2386 (N_2386,N_1842,N_2188);
nor U2387 (N_2387,N_1921,N_2168);
or U2388 (N_2388,N_1864,N_1669);
or U2389 (N_2389,N_2185,N_2035);
or U2390 (N_2390,N_1879,N_1898);
xor U2391 (N_2391,N_2118,N_1966);
nand U2392 (N_2392,N_1957,N_1704);
or U2393 (N_2393,N_2039,N_2234);
nor U2394 (N_2394,N_1633,N_1710);
nand U2395 (N_2395,N_1661,N_1687);
nor U2396 (N_2396,N_1959,N_2191);
nand U2397 (N_2397,N_1569,N_1615);
and U2398 (N_2398,N_2139,N_1949);
or U2399 (N_2399,N_1531,N_1969);
and U2400 (N_2400,N_1647,N_2197);
or U2401 (N_2401,N_2145,N_1608);
and U2402 (N_2402,N_1662,N_1588);
nand U2403 (N_2403,N_1996,N_1743);
nand U2404 (N_2404,N_1652,N_1803);
nand U2405 (N_2405,N_1846,N_2008);
xor U2406 (N_2406,N_2002,N_1593);
and U2407 (N_2407,N_1979,N_1696);
nand U2408 (N_2408,N_1568,N_1715);
or U2409 (N_2409,N_1947,N_1915);
nor U2410 (N_2410,N_1719,N_1520);
nor U2411 (N_2411,N_1795,N_1843);
nand U2412 (N_2412,N_1563,N_1897);
nor U2413 (N_2413,N_1939,N_1946);
nand U2414 (N_2414,N_2201,N_1649);
nand U2415 (N_2415,N_1948,N_2199);
xnor U2416 (N_2416,N_2112,N_2076);
xnor U2417 (N_2417,N_1961,N_1735);
nor U2418 (N_2418,N_2038,N_1922);
and U2419 (N_2419,N_1785,N_1579);
or U2420 (N_2420,N_2009,N_1682);
nand U2421 (N_2421,N_2165,N_1738);
nor U2422 (N_2422,N_2161,N_1517);
or U2423 (N_2423,N_1508,N_1932);
or U2424 (N_2424,N_1548,N_2131);
and U2425 (N_2425,N_1821,N_1596);
nor U2426 (N_2426,N_1874,N_2095);
nor U2427 (N_2427,N_2023,N_1527);
or U2428 (N_2428,N_1761,N_2062);
or U2429 (N_2429,N_2110,N_1663);
and U2430 (N_2430,N_1926,N_2049);
nor U2431 (N_2431,N_2081,N_2054);
or U2432 (N_2432,N_1500,N_1901);
nand U2433 (N_2433,N_1571,N_2166);
nand U2434 (N_2434,N_1800,N_1958);
nand U2435 (N_2435,N_1747,N_2032);
or U2436 (N_2436,N_2238,N_2230);
or U2437 (N_2437,N_2140,N_1702);
or U2438 (N_2438,N_1854,N_2195);
and U2439 (N_2439,N_1630,N_1636);
nor U2440 (N_2440,N_1576,N_2092);
nand U2441 (N_2441,N_1524,N_1564);
nand U2442 (N_2442,N_2019,N_2026);
nand U2443 (N_2443,N_1794,N_2194);
and U2444 (N_2444,N_1978,N_1988);
nand U2445 (N_2445,N_2237,N_1683);
and U2446 (N_2446,N_1982,N_1565);
or U2447 (N_2447,N_2246,N_1541);
nor U2448 (N_2448,N_2048,N_1540);
nor U2449 (N_2449,N_1970,N_2147);
nand U2450 (N_2450,N_2010,N_1889);
or U2451 (N_2451,N_1573,N_1600);
or U2452 (N_2452,N_2030,N_1938);
or U2453 (N_2453,N_2059,N_2158);
nor U2454 (N_2454,N_1550,N_1611);
nor U2455 (N_2455,N_1519,N_1575);
nor U2456 (N_2456,N_1685,N_1515);
nor U2457 (N_2457,N_1513,N_2193);
nor U2458 (N_2458,N_2091,N_1927);
nor U2459 (N_2459,N_1561,N_1742);
nor U2460 (N_2460,N_1692,N_1868);
and U2461 (N_2461,N_1778,N_1693);
xor U2462 (N_2462,N_1976,N_1777);
xnor U2463 (N_2463,N_2198,N_2187);
nand U2464 (N_2464,N_2028,N_1916);
xor U2465 (N_2465,N_2116,N_1668);
and U2466 (N_2466,N_1553,N_2162);
xnor U2467 (N_2467,N_1918,N_1616);
xor U2468 (N_2468,N_1549,N_2130);
and U2469 (N_2469,N_1832,N_1581);
nand U2470 (N_2470,N_1808,N_1766);
nand U2471 (N_2471,N_1881,N_1645);
nand U2472 (N_2472,N_1641,N_1792);
or U2473 (N_2473,N_1760,N_2202);
or U2474 (N_2474,N_1643,N_1560);
and U2475 (N_2475,N_1883,N_1739);
nor U2476 (N_2476,N_2128,N_1844);
nand U2477 (N_2477,N_1853,N_1506);
nor U2478 (N_2478,N_2097,N_1612);
and U2479 (N_2479,N_2152,N_1833);
nor U2480 (N_2480,N_2015,N_1586);
or U2481 (N_2481,N_1523,N_1512);
nor U2482 (N_2482,N_1867,N_2215);
nor U2483 (N_2483,N_2222,N_2085);
nor U2484 (N_2484,N_1981,N_2064);
nand U2485 (N_2485,N_1816,N_1504);
xor U2486 (N_2486,N_2227,N_1629);
nor U2487 (N_2487,N_1951,N_1823);
xnor U2488 (N_2488,N_1906,N_1791);
xnor U2489 (N_2489,N_1741,N_2090);
or U2490 (N_2490,N_1783,N_1749);
and U2491 (N_2491,N_1681,N_2096);
nor U2492 (N_2492,N_1831,N_1873);
nor U2493 (N_2493,N_1665,N_1736);
and U2494 (N_2494,N_1974,N_1776);
nor U2495 (N_2495,N_1678,N_1937);
and U2496 (N_2496,N_1954,N_1716);
or U2497 (N_2497,N_1871,N_1914);
xnor U2498 (N_2498,N_1836,N_1603);
nor U2499 (N_2499,N_2138,N_1542);
xor U2500 (N_2500,N_2216,N_2069);
nor U2501 (N_2501,N_2077,N_1758);
nor U2502 (N_2502,N_2239,N_1554);
or U2503 (N_2503,N_1852,N_1526);
nand U2504 (N_2504,N_1806,N_1675);
or U2505 (N_2505,N_1829,N_1903);
nand U2506 (N_2506,N_1911,N_1804);
nand U2507 (N_2507,N_2129,N_2179);
or U2508 (N_2508,N_2134,N_1725);
or U2509 (N_2509,N_2016,N_1977);
and U2510 (N_2510,N_1509,N_1557);
nor U2511 (N_2511,N_1980,N_1556);
nor U2512 (N_2512,N_2011,N_1875);
nor U2513 (N_2513,N_1887,N_1637);
nor U2514 (N_2514,N_1908,N_1972);
nor U2515 (N_2515,N_1894,N_1807);
or U2516 (N_2516,N_1847,N_2014);
nor U2517 (N_2517,N_2217,N_1667);
nor U2518 (N_2518,N_1805,N_2146);
and U2519 (N_2519,N_1606,N_1728);
and U2520 (N_2520,N_2225,N_1533);
nor U2521 (N_2521,N_1709,N_1930);
or U2522 (N_2522,N_1953,N_1534);
or U2523 (N_2523,N_2079,N_1689);
and U2524 (N_2524,N_1748,N_2192);
nand U2525 (N_2525,N_1539,N_2056);
nor U2526 (N_2526,N_1507,N_2033);
and U2527 (N_2527,N_1934,N_2137);
or U2528 (N_2528,N_1920,N_1729);
and U2529 (N_2529,N_1793,N_1674);
xnor U2530 (N_2530,N_1814,N_1820);
nor U2531 (N_2531,N_2204,N_1731);
xor U2532 (N_2532,N_2024,N_1521);
nor U2533 (N_2533,N_2213,N_2221);
and U2534 (N_2534,N_2057,N_1952);
or U2535 (N_2535,N_1992,N_1975);
and U2536 (N_2536,N_1841,N_2135);
xor U2537 (N_2537,N_2080,N_2149);
nor U2538 (N_2538,N_1798,N_2117);
nor U2539 (N_2539,N_1767,N_1525);
and U2540 (N_2540,N_1825,N_2184);
nand U2541 (N_2541,N_2025,N_1635);
xnor U2542 (N_2542,N_1753,N_1684);
xor U2543 (N_2543,N_1884,N_1923);
nand U2544 (N_2544,N_2100,N_1601);
nand U2545 (N_2545,N_2235,N_1518);
xor U2546 (N_2546,N_1701,N_1673);
nand U2547 (N_2547,N_1730,N_1658);
nor U2548 (N_2548,N_1878,N_1931);
nand U2549 (N_2549,N_1899,N_1765);
and U2550 (N_2550,N_2171,N_1583);
nand U2551 (N_2551,N_2233,N_1613);
or U2552 (N_2552,N_1621,N_2243);
xor U2553 (N_2553,N_1733,N_1912);
and U2554 (N_2554,N_1640,N_1547);
and U2555 (N_2555,N_1997,N_2101);
and U2556 (N_2556,N_2093,N_1837);
xnor U2557 (N_2557,N_1502,N_1781);
nor U2558 (N_2558,N_2051,N_1642);
xor U2559 (N_2559,N_1745,N_1577);
nor U2560 (N_2560,N_1570,N_1797);
nand U2561 (N_2561,N_1587,N_1936);
nor U2562 (N_2562,N_1888,N_1830);
nor U2563 (N_2563,N_1671,N_1964);
nand U2564 (N_2564,N_1774,N_1909);
or U2565 (N_2565,N_1891,N_1657);
or U2566 (N_2566,N_2164,N_1812);
and U2567 (N_2567,N_2044,N_1706);
or U2568 (N_2568,N_2127,N_1634);
and U2569 (N_2569,N_1907,N_1602);
nor U2570 (N_2570,N_2067,N_1856);
or U2571 (N_2571,N_1986,N_1708);
or U2572 (N_2572,N_2066,N_1880);
or U2573 (N_2573,N_1695,N_2186);
xnor U2574 (N_2574,N_1589,N_1726);
xor U2575 (N_2575,N_2108,N_2212);
nor U2576 (N_2576,N_2231,N_1924);
nor U2577 (N_2577,N_2244,N_2144);
xnor U2578 (N_2578,N_1799,N_1653);
nand U2579 (N_2579,N_2078,N_1599);
or U2580 (N_2580,N_2189,N_1772);
nor U2581 (N_2581,N_2208,N_1537);
and U2582 (N_2582,N_1535,N_1700);
or U2583 (N_2583,N_2058,N_1861);
and U2584 (N_2584,N_2073,N_1790);
nor U2585 (N_2585,N_2068,N_1529);
and U2586 (N_2586,N_2001,N_2153);
or U2587 (N_2587,N_1670,N_1555);
nor U2588 (N_2588,N_2050,N_1594);
and U2589 (N_2589,N_2086,N_1552);
nor U2590 (N_2590,N_2113,N_1648);
nor U2591 (N_2591,N_1627,N_2087);
or U2592 (N_2592,N_1965,N_1732);
nand U2593 (N_2593,N_1876,N_1817);
or U2594 (N_2594,N_1904,N_1995);
nand U2595 (N_2595,N_1703,N_2102);
or U2596 (N_2596,N_1827,N_2004);
and U2597 (N_2597,N_2151,N_1625);
nor U2598 (N_2598,N_2125,N_1956);
nand U2599 (N_2599,N_1770,N_2124);
nand U2600 (N_2600,N_1810,N_2150);
or U2601 (N_2601,N_1801,N_1697);
xor U2602 (N_2602,N_1718,N_2070);
or U2603 (N_2603,N_2136,N_2229);
nor U2604 (N_2604,N_2157,N_2088);
and U2605 (N_2605,N_1796,N_1929);
and U2606 (N_2606,N_1872,N_1664);
nand U2607 (N_2607,N_2012,N_2178);
and U2608 (N_2608,N_1768,N_1538);
and U2609 (N_2609,N_1723,N_2206);
or U2610 (N_2610,N_1845,N_1987);
nor U2611 (N_2611,N_1962,N_1559);
and U2612 (N_2612,N_1578,N_1688);
nor U2613 (N_2613,N_1598,N_1740);
or U2614 (N_2614,N_1950,N_1933);
and U2615 (N_2615,N_1624,N_1973);
or U2616 (N_2616,N_1503,N_2003);
nand U2617 (N_2617,N_2027,N_2123);
and U2618 (N_2618,N_2200,N_1651);
and U2619 (N_2619,N_2106,N_1764);
nor U2620 (N_2620,N_2043,N_1574);
nor U2621 (N_2621,N_1893,N_1646);
nor U2622 (N_2622,N_2174,N_2031);
nand U2623 (N_2623,N_2029,N_1679);
nor U2624 (N_2624,N_1584,N_1935);
and U2625 (N_2625,N_1713,N_2072);
nor U2626 (N_2626,N_1519,N_1670);
nor U2627 (N_2627,N_1674,N_1709);
or U2628 (N_2628,N_2098,N_2034);
xor U2629 (N_2629,N_1986,N_1899);
nor U2630 (N_2630,N_1596,N_2240);
or U2631 (N_2631,N_2190,N_2235);
or U2632 (N_2632,N_2230,N_1694);
nor U2633 (N_2633,N_2168,N_1757);
nand U2634 (N_2634,N_2211,N_2051);
nor U2635 (N_2635,N_1968,N_1817);
xor U2636 (N_2636,N_2219,N_1715);
nor U2637 (N_2637,N_1630,N_1956);
or U2638 (N_2638,N_1990,N_1728);
nand U2639 (N_2639,N_2229,N_1516);
and U2640 (N_2640,N_1824,N_1740);
or U2641 (N_2641,N_1804,N_1694);
nand U2642 (N_2642,N_1625,N_2007);
or U2643 (N_2643,N_2071,N_2183);
nor U2644 (N_2644,N_2185,N_1504);
or U2645 (N_2645,N_2031,N_1711);
and U2646 (N_2646,N_1640,N_2114);
or U2647 (N_2647,N_1817,N_1664);
nand U2648 (N_2648,N_1565,N_1860);
or U2649 (N_2649,N_1715,N_1533);
or U2650 (N_2650,N_1635,N_1866);
nand U2651 (N_2651,N_1696,N_1995);
or U2652 (N_2652,N_1981,N_1718);
nand U2653 (N_2653,N_1762,N_1836);
xor U2654 (N_2654,N_1559,N_1927);
nor U2655 (N_2655,N_1968,N_1955);
xnor U2656 (N_2656,N_1616,N_1641);
nor U2657 (N_2657,N_1657,N_1642);
nor U2658 (N_2658,N_2083,N_1625);
nand U2659 (N_2659,N_1729,N_1681);
nor U2660 (N_2660,N_2094,N_1614);
nor U2661 (N_2661,N_2161,N_1929);
or U2662 (N_2662,N_1996,N_1801);
xor U2663 (N_2663,N_2063,N_1901);
and U2664 (N_2664,N_1773,N_2212);
and U2665 (N_2665,N_1902,N_2018);
xor U2666 (N_2666,N_2175,N_2158);
xor U2667 (N_2667,N_1903,N_1660);
and U2668 (N_2668,N_1701,N_1794);
nand U2669 (N_2669,N_1709,N_1963);
and U2670 (N_2670,N_1857,N_2226);
nand U2671 (N_2671,N_2122,N_1579);
and U2672 (N_2672,N_1988,N_1834);
nand U2673 (N_2673,N_1724,N_2111);
and U2674 (N_2674,N_1707,N_2185);
xnor U2675 (N_2675,N_1789,N_2090);
nor U2676 (N_2676,N_1729,N_1984);
and U2677 (N_2677,N_2105,N_1849);
and U2678 (N_2678,N_2028,N_1672);
and U2679 (N_2679,N_1962,N_2248);
nand U2680 (N_2680,N_2069,N_1815);
nand U2681 (N_2681,N_2014,N_1952);
nor U2682 (N_2682,N_1841,N_1559);
and U2683 (N_2683,N_2178,N_1765);
xnor U2684 (N_2684,N_1614,N_1711);
and U2685 (N_2685,N_1557,N_1933);
and U2686 (N_2686,N_1749,N_1522);
or U2687 (N_2687,N_1550,N_2009);
nor U2688 (N_2688,N_1704,N_2221);
and U2689 (N_2689,N_1845,N_1669);
xor U2690 (N_2690,N_1755,N_1929);
xor U2691 (N_2691,N_1956,N_1992);
nor U2692 (N_2692,N_1508,N_1956);
xor U2693 (N_2693,N_1784,N_1863);
and U2694 (N_2694,N_1897,N_2172);
nor U2695 (N_2695,N_2196,N_2023);
and U2696 (N_2696,N_1642,N_1745);
nand U2697 (N_2697,N_2069,N_1572);
and U2698 (N_2698,N_1815,N_1665);
or U2699 (N_2699,N_2218,N_2152);
nand U2700 (N_2700,N_2023,N_1923);
or U2701 (N_2701,N_2146,N_1888);
xor U2702 (N_2702,N_1640,N_1916);
xnor U2703 (N_2703,N_2198,N_1966);
nand U2704 (N_2704,N_1922,N_2129);
nor U2705 (N_2705,N_2157,N_1779);
or U2706 (N_2706,N_2058,N_1729);
nand U2707 (N_2707,N_2190,N_1898);
nor U2708 (N_2708,N_1605,N_1977);
nor U2709 (N_2709,N_2063,N_2085);
xor U2710 (N_2710,N_1724,N_1880);
and U2711 (N_2711,N_1506,N_1731);
or U2712 (N_2712,N_1921,N_1696);
nand U2713 (N_2713,N_1580,N_1799);
nand U2714 (N_2714,N_2035,N_1905);
and U2715 (N_2715,N_1865,N_2112);
and U2716 (N_2716,N_1529,N_1831);
nor U2717 (N_2717,N_1856,N_2223);
nor U2718 (N_2718,N_1945,N_1659);
or U2719 (N_2719,N_1512,N_1601);
nand U2720 (N_2720,N_1612,N_1606);
nor U2721 (N_2721,N_2053,N_2112);
and U2722 (N_2722,N_2186,N_2170);
or U2723 (N_2723,N_1704,N_2072);
or U2724 (N_2724,N_1972,N_1523);
nand U2725 (N_2725,N_2245,N_1917);
nand U2726 (N_2726,N_1954,N_1890);
nor U2727 (N_2727,N_2141,N_1703);
nor U2728 (N_2728,N_1724,N_1841);
nand U2729 (N_2729,N_2082,N_2053);
nor U2730 (N_2730,N_2091,N_2206);
or U2731 (N_2731,N_1965,N_1914);
xnor U2732 (N_2732,N_2205,N_2014);
nand U2733 (N_2733,N_2021,N_1661);
nor U2734 (N_2734,N_2162,N_1636);
and U2735 (N_2735,N_1898,N_1930);
or U2736 (N_2736,N_1805,N_2024);
xor U2737 (N_2737,N_1772,N_1998);
nor U2738 (N_2738,N_1802,N_1600);
or U2739 (N_2739,N_1997,N_1556);
xor U2740 (N_2740,N_1872,N_1918);
nand U2741 (N_2741,N_1536,N_1566);
and U2742 (N_2742,N_2058,N_1761);
nor U2743 (N_2743,N_1824,N_2007);
nor U2744 (N_2744,N_1621,N_2121);
nor U2745 (N_2745,N_2109,N_1958);
nand U2746 (N_2746,N_1655,N_1747);
nand U2747 (N_2747,N_1976,N_1632);
nand U2748 (N_2748,N_1866,N_1821);
xnor U2749 (N_2749,N_1932,N_1928);
nand U2750 (N_2750,N_1671,N_1558);
nor U2751 (N_2751,N_1766,N_1758);
nand U2752 (N_2752,N_1993,N_1797);
nor U2753 (N_2753,N_2137,N_2237);
nor U2754 (N_2754,N_1967,N_1945);
nor U2755 (N_2755,N_1748,N_1865);
nand U2756 (N_2756,N_1838,N_2038);
or U2757 (N_2757,N_2106,N_1896);
nand U2758 (N_2758,N_2232,N_2174);
nand U2759 (N_2759,N_2055,N_1682);
and U2760 (N_2760,N_1749,N_1931);
or U2761 (N_2761,N_1758,N_1980);
or U2762 (N_2762,N_2086,N_2019);
nand U2763 (N_2763,N_2130,N_2141);
nor U2764 (N_2764,N_2015,N_1726);
xnor U2765 (N_2765,N_1902,N_1906);
and U2766 (N_2766,N_1858,N_2118);
and U2767 (N_2767,N_2112,N_1974);
or U2768 (N_2768,N_2046,N_2146);
or U2769 (N_2769,N_1526,N_1900);
nor U2770 (N_2770,N_1887,N_1584);
and U2771 (N_2771,N_1602,N_2040);
and U2772 (N_2772,N_2007,N_1983);
nand U2773 (N_2773,N_1509,N_1614);
and U2774 (N_2774,N_1676,N_1894);
nand U2775 (N_2775,N_2197,N_2024);
and U2776 (N_2776,N_1826,N_1890);
nor U2777 (N_2777,N_1678,N_2015);
nand U2778 (N_2778,N_1765,N_1993);
or U2779 (N_2779,N_2128,N_1835);
or U2780 (N_2780,N_1720,N_1640);
and U2781 (N_2781,N_1603,N_1982);
nand U2782 (N_2782,N_2013,N_1916);
and U2783 (N_2783,N_1987,N_1848);
and U2784 (N_2784,N_2203,N_2054);
xnor U2785 (N_2785,N_2187,N_2235);
nor U2786 (N_2786,N_1524,N_1768);
nand U2787 (N_2787,N_1702,N_1682);
nor U2788 (N_2788,N_1854,N_2127);
nor U2789 (N_2789,N_2017,N_2081);
nor U2790 (N_2790,N_2044,N_2124);
nand U2791 (N_2791,N_1704,N_2154);
or U2792 (N_2792,N_2122,N_1966);
and U2793 (N_2793,N_2000,N_2231);
and U2794 (N_2794,N_2188,N_2041);
xor U2795 (N_2795,N_1820,N_1543);
nor U2796 (N_2796,N_2243,N_1638);
and U2797 (N_2797,N_1509,N_2033);
nor U2798 (N_2798,N_1709,N_1999);
nand U2799 (N_2799,N_1771,N_1821);
or U2800 (N_2800,N_1728,N_2120);
xnor U2801 (N_2801,N_1746,N_1589);
and U2802 (N_2802,N_1856,N_1756);
nand U2803 (N_2803,N_1730,N_1763);
or U2804 (N_2804,N_1954,N_2219);
nand U2805 (N_2805,N_2156,N_1794);
or U2806 (N_2806,N_1916,N_1893);
nand U2807 (N_2807,N_1569,N_2233);
nor U2808 (N_2808,N_1787,N_1588);
and U2809 (N_2809,N_1577,N_2228);
nand U2810 (N_2810,N_1825,N_1549);
and U2811 (N_2811,N_1536,N_2168);
or U2812 (N_2812,N_2209,N_1923);
nand U2813 (N_2813,N_1787,N_1619);
and U2814 (N_2814,N_2248,N_2104);
and U2815 (N_2815,N_1689,N_2091);
nand U2816 (N_2816,N_1848,N_1973);
or U2817 (N_2817,N_1907,N_2108);
nand U2818 (N_2818,N_2163,N_2205);
xnor U2819 (N_2819,N_1512,N_1779);
xor U2820 (N_2820,N_1638,N_1786);
nand U2821 (N_2821,N_1962,N_1527);
and U2822 (N_2822,N_1504,N_1523);
xnor U2823 (N_2823,N_2177,N_1544);
or U2824 (N_2824,N_1543,N_2034);
or U2825 (N_2825,N_1626,N_1531);
or U2826 (N_2826,N_1884,N_1543);
nand U2827 (N_2827,N_1659,N_1632);
or U2828 (N_2828,N_1696,N_1966);
nand U2829 (N_2829,N_2241,N_1716);
nand U2830 (N_2830,N_1820,N_2085);
nor U2831 (N_2831,N_1866,N_2058);
xnor U2832 (N_2832,N_1549,N_2198);
nor U2833 (N_2833,N_2015,N_1986);
nand U2834 (N_2834,N_1835,N_2085);
nor U2835 (N_2835,N_2199,N_1883);
or U2836 (N_2836,N_1630,N_1882);
or U2837 (N_2837,N_2137,N_2218);
and U2838 (N_2838,N_1975,N_1645);
nor U2839 (N_2839,N_2127,N_2141);
or U2840 (N_2840,N_1771,N_1827);
nor U2841 (N_2841,N_1730,N_1511);
or U2842 (N_2842,N_1702,N_2231);
nor U2843 (N_2843,N_1944,N_1997);
nor U2844 (N_2844,N_2148,N_2155);
nand U2845 (N_2845,N_1658,N_1974);
xor U2846 (N_2846,N_2003,N_2150);
or U2847 (N_2847,N_1749,N_1795);
nand U2848 (N_2848,N_1578,N_1966);
or U2849 (N_2849,N_1848,N_1862);
and U2850 (N_2850,N_1506,N_1823);
nand U2851 (N_2851,N_2234,N_2034);
xor U2852 (N_2852,N_2129,N_2116);
or U2853 (N_2853,N_2079,N_1678);
nor U2854 (N_2854,N_1786,N_1941);
and U2855 (N_2855,N_1576,N_1871);
nand U2856 (N_2856,N_1739,N_1898);
nor U2857 (N_2857,N_1932,N_2006);
nor U2858 (N_2858,N_2028,N_1620);
or U2859 (N_2859,N_1767,N_1971);
or U2860 (N_2860,N_2168,N_1737);
nand U2861 (N_2861,N_1510,N_1896);
nand U2862 (N_2862,N_2087,N_1953);
and U2863 (N_2863,N_2233,N_1923);
or U2864 (N_2864,N_2074,N_1613);
and U2865 (N_2865,N_2002,N_2153);
nand U2866 (N_2866,N_2109,N_1601);
and U2867 (N_2867,N_1646,N_1612);
nand U2868 (N_2868,N_1725,N_1851);
nor U2869 (N_2869,N_1998,N_2055);
nand U2870 (N_2870,N_2142,N_1879);
nand U2871 (N_2871,N_1752,N_1858);
or U2872 (N_2872,N_1929,N_2076);
nor U2873 (N_2873,N_2117,N_1664);
nor U2874 (N_2874,N_1727,N_1569);
nor U2875 (N_2875,N_2162,N_1644);
nor U2876 (N_2876,N_1908,N_1619);
nor U2877 (N_2877,N_1862,N_1926);
and U2878 (N_2878,N_1929,N_1841);
xor U2879 (N_2879,N_1889,N_2222);
nor U2880 (N_2880,N_1673,N_1906);
xor U2881 (N_2881,N_1763,N_1540);
and U2882 (N_2882,N_2107,N_1757);
nand U2883 (N_2883,N_1521,N_1516);
or U2884 (N_2884,N_2162,N_2131);
nor U2885 (N_2885,N_1738,N_1793);
nand U2886 (N_2886,N_2047,N_1871);
or U2887 (N_2887,N_2137,N_2117);
nand U2888 (N_2888,N_1633,N_1806);
nor U2889 (N_2889,N_2127,N_2051);
nand U2890 (N_2890,N_2118,N_1520);
nand U2891 (N_2891,N_2101,N_2234);
nor U2892 (N_2892,N_1977,N_1549);
nor U2893 (N_2893,N_1614,N_1530);
xnor U2894 (N_2894,N_2098,N_1980);
or U2895 (N_2895,N_1526,N_1785);
nor U2896 (N_2896,N_2227,N_1805);
nor U2897 (N_2897,N_1815,N_1765);
nand U2898 (N_2898,N_1540,N_2049);
and U2899 (N_2899,N_1878,N_1715);
nor U2900 (N_2900,N_1679,N_1606);
nor U2901 (N_2901,N_2173,N_1658);
or U2902 (N_2902,N_1627,N_1979);
or U2903 (N_2903,N_1906,N_2114);
nand U2904 (N_2904,N_1765,N_1679);
xor U2905 (N_2905,N_2088,N_1977);
xor U2906 (N_2906,N_2114,N_1770);
nor U2907 (N_2907,N_2006,N_1560);
xnor U2908 (N_2908,N_2223,N_1630);
xnor U2909 (N_2909,N_1731,N_1593);
nor U2910 (N_2910,N_2035,N_2125);
and U2911 (N_2911,N_1751,N_1618);
xnor U2912 (N_2912,N_2128,N_1973);
and U2913 (N_2913,N_2144,N_2089);
nor U2914 (N_2914,N_1836,N_1755);
or U2915 (N_2915,N_2244,N_1593);
nand U2916 (N_2916,N_1772,N_1522);
nor U2917 (N_2917,N_1901,N_2097);
and U2918 (N_2918,N_1963,N_1536);
nor U2919 (N_2919,N_2032,N_1558);
nor U2920 (N_2920,N_2226,N_2089);
or U2921 (N_2921,N_1805,N_1855);
or U2922 (N_2922,N_2159,N_1506);
nand U2923 (N_2923,N_1864,N_2155);
or U2924 (N_2924,N_2031,N_1872);
nor U2925 (N_2925,N_1612,N_2048);
nand U2926 (N_2926,N_2101,N_1947);
nor U2927 (N_2927,N_2064,N_1918);
nor U2928 (N_2928,N_2051,N_1626);
xnor U2929 (N_2929,N_2216,N_2242);
or U2930 (N_2930,N_1705,N_2120);
or U2931 (N_2931,N_1813,N_1838);
or U2932 (N_2932,N_2057,N_1923);
or U2933 (N_2933,N_1962,N_2147);
nand U2934 (N_2934,N_2130,N_1664);
nand U2935 (N_2935,N_1574,N_1543);
xnor U2936 (N_2936,N_1945,N_1866);
and U2937 (N_2937,N_2032,N_2005);
or U2938 (N_2938,N_1617,N_2006);
nand U2939 (N_2939,N_1600,N_2237);
or U2940 (N_2940,N_2040,N_2201);
nand U2941 (N_2941,N_1891,N_1597);
and U2942 (N_2942,N_1586,N_1817);
nor U2943 (N_2943,N_2112,N_1954);
nor U2944 (N_2944,N_2169,N_1958);
xnor U2945 (N_2945,N_1612,N_2015);
nand U2946 (N_2946,N_2229,N_2199);
nand U2947 (N_2947,N_1763,N_1859);
nand U2948 (N_2948,N_2083,N_2133);
or U2949 (N_2949,N_1543,N_1985);
and U2950 (N_2950,N_2068,N_2185);
nor U2951 (N_2951,N_2081,N_1675);
nor U2952 (N_2952,N_1851,N_1680);
nor U2953 (N_2953,N_2229,N_2204);
nor U2954 (N_2954,N_1793,N_1538);
and U2955 (N_2955,N_1691,N_1919);
or U2956 (N_2956,N_2075,N_2149);
xnor U2957 (N_2957,N_2005,N_1975);
nand U2958 (N_2958,N_2010,N_1515);
nor U2959 (N_2959,N_2126,N_1610);
and U2960 (N_2960,N_1603,N_1765);
or U2961 (N_2961,N_2158,N_1746);
nand U2962 (N_2962,N_1918,N_1726);
and U2963 (N_2963,N_2111,N_1704);
nand U2964 (N_2964,N_1916,N_2091);
nor U2965 (N_2965,N_1594,N_2151);
or U2966 (N_2966,N_2013,N_1620);
nand U2967 (N_2967,N_2242,N_2048);
nand U2968 (N_2968,N_2032,N_2063);
nor U2969 (N_2969,N_1635,N_1683);
or U2970 (N_2970,N_1978,N_1785);
nor U2971 (N_2971,N_2209,N_2158);
nand U2972 (N_2972,N_2081,N_1520);
or U2973 (N_2973,N_2080,N_1954);
nand U2974 (N_2974,N_1581,N_1789);
or U2975 (N_2975,N_1857,N_2188);
nand U2976 (N_2976,N_2092,N_2155);
xor U2977 (N_2977,N_1635,N_1927);
xor U2978 (N_2978,N_2024,N_1830);
nor U2979 (N_2979,N_2152,N_2225);
or U2980 (N_2980,N_1797,N_2076);
and U2981 (N_2981,N_2110,N_1758);
nand U2982 (N_2982,N_2074,N_1602);
nand U2983 (N_2983,N_2233,N_1824);
nand U2984 (N_2984,N_2084,N_1953);
xnor U2985 (N_2985,N_1573,N_1939);
and U2986 (N_2986,N_2240,N_2143);
nor U2987 (N_2987,N_1932,N_2103);
nand U2988 (N_2988,N_2182,N_1817);
or U2989 (N_2989,N_1830,N_2100);
nor U2990 (N_2990,N_1861,N_1798);
and U2991 (N_2991,N_1524,N_1971);
and U2992 (N_2992,N_2192,N_2009);
nand U2993 (N_2993,N_1623,N_1677);
and U2994 (N_2994,N_1632,N_2151);
nand U2995 (N_2995,N_2063,N_1742);
and U2996 (N_2996,N_1548,N_2115);
nor U2997 (N_2997,N_1517,N_1918);
nor U2998 (N_2998,N_1584,N_2198);
or U2999 (N_2999,N_1621,N_1566);
xor UO_0 (O_0,N_2793,N_2451);
or UO_1 (O_1,N_2782,N_2719);
xor UO_2 (O_2,N_2851,N_2869);
nor UO_3 (O_3,N_2340,N_2597);
xnor UO_4 (O_4,N_2570,N_2263);
nand UO_5 (O_5,N_2726,N_2936);
or UO_6 (O_6,N_2560,N_2567);
or UO_7 (O_7,N_2556,N_2583);
nor UO_8 (O_8,N_2364,N_2693);
nand UO_9 (O_9,N_2659,N_2552);
and UO_10 (O_10,N_2706,N_2434);
nor UO_11 (O_11,N_2800,N_2331);
xor UO_12 (O_12,N_2920,N_2426);
or UO_13 (O_13,N_2632,N_2691);
or UO_14 (O_14,N_2471,N_2943);
or UO_15 (O_15,N_2277,N_2544);
and UO_16 (O_16,N_2348,N_2279);
xnor UO_17 (O_17,N_2836,N_2715);
and UO_18 (O_18,N_2507,N_2728);
and UO_19 (O_19,N_2355,N_2815);
or UO_20 (O_20,N_2984,N_2395);
or UO_21 (O_21,N_2535,N_2673);
or UO_22 (O_22,N_2911,N_2973);
and UO_23 (O_23,N_2498,N_2321);
nor UO_24 (O_24,N_2538,N_2950);
or UO_25 (O_25,N_2690,N_2785);
nor UO_26 (O_26,N_2268,N_2937);
xnor UO_27 (O_27,N_2999,N_2695);
nor UO_28 (O_28,N_2668,N_2998);
and UO_29 (O_29,N_2712,N_2577);
nand UO_30 (O_30,N_2294,N_2772);
nand UO_31 (O_31,N_2788,N_2494);
and UO_32 (O_32,N_2826,N_2926);
nand UO_33 (O_33,N_2502,N_2796);
and UO_34 (O_34,N_2616,N_2529);
xnor UO_35 (O_35,N_2452,N_2311);
and UO_36 (O_36,N_2765,N_2462);
and UO_37 (O_37,N_2805,N_2550);
nand UO_38 (O_38,N_2270,N_2734);
and UO_39 (O_39,N_2993,N_2424);
or UO_40 (O_40,N_2411,N_2795);
and UO_41 (O_41,N_2931,N_2422);
nand UO_42 (O_42,N_2913,N_2915);
nor UO_43 (O_43,N_2446,N_2770);
nand UO_44 (O_44,N_2829,N_2403);
nand UO_45 (O_45,N_2887,N_2359);
and UO_46 (O_46,N_2262,N_2644);
or UO_47 (O_47,N_2580,N_2794);
xnor UO_48 (O_48,N_2724,N_2528);
nor UO_49 (O_49,N_2319,N_2656);
xnor UO_50 (O_50,N_2478,N_2473);
or UO_51 (O_51,N_2375,N_2718);
nor UO_52 (O_52,N_2990,N_2288);
nor UO_53 (O_53,N_2613,N_2429);
or UO_54 (O_54,N_2389,N_2681);
nor UO_55 (O_55,N_2991,N_2628);
or UO_56 (O_56,N_2350,N_2774);
xor UO_57 (O_57,N_2679,N_2463);
nand UO_58 (O_58,N_2781,N_2641);
or UO_59 (O_59,N_2326,N_2773);
or UO_60 (O_60,N_2833,N_2914);
and UO_61 (O_61,N_2401,N_2479);
xnor UO_62 (O_62,N_2338,N_2332);
nand UO_63 (O_63,N_2889,N_2566);
nor UO_64 (O_64,N_2366,N_2299);
nor UO_65 (O_65,N_2652,N_2421);
xnor UO_66 (O_66,N_2777,N_2907);
or UO_67 (O_67,N_2470,N_2514);
or UO_68 (O_68,N_2458,N_2307);
and UO_69 (O_69,N_2428,N_2354);
nand UO_70 (O_70,N_2612,N_2393);
and UO_71 (O_71,N_2454,N_2399);
or UO_72 (O_72,N_2757,N_2947);
nand UO_73 (O_73,N_2368,N_2864);
nor UO_74 (O_74,N_2335,N_2663);
or UO_75 (O_75,N_2832,N_2453);
and UO_76 (O_76,N_2606,N_2658);
nand UO_77 (O_77,N_2349,N_2868);
nor UO_78 (O_78,N_2954,N_2316);
nand UO_79 (O_79,N_2358,N_2992);
and UO_80 (O_80,N_2572,N_2962);
nand UO_81 (O_81,N_2532,N_2251);
nand UO_82 (O_82,N_2447,N_2922);
or UO_83 (O_83,N_2575,N_2825);
nor UO_84 (O_84,N_2394,N_2259);
nand UO_85 (O_85,N_2844,N_2687);
or UO_86 (O_86,N_2599,N_2390);
nor UO_87 (O_87,N_2490,N_2565);
and UO_88 (O_88,N_2571,N_2667);
or UO_89 (O_89,N_2505,N_2787);
nor UO_90 (O_90,N_2645,N_2347);
nor UO_91 (O_91,N_2665,N_2702);
nor UO_92 (O_92,N_2808,N_2305);
nand UO_93 (O_93,N_2703,N_2760);
nand UO_94 (O_94,N_2953,N_2555);
nand UO_95 (O_95,N_2496,N_2798);
nand UO_96 (O_96,N_2847,N_2670);
nor UO_97 (O_97,N_2877,N_2987);
nor UO_98 (O_98,N_2831,N_2743);
nor UO_99 (O_99,N_2725,N_2607);
nor UO_100 (O_100,N_2980,N_2880);
and UO_101 (O_101,N_2482,N_2472);
nand UO_102 (O_102,N_2650,N_2853);
nand UO_103 (O_103,N_2404,N_2465);
or UO_104 (O_104,N_2630,N_2314);
nand UO_105 (O_105,N_2910,N_2308);
xnor UO_106 (O_106,N_2891,N_2686);
and UO_107 (O_107,N_2365,N_2378);
or UO_108 (O_108,N_2736,N_2557);
nand UO_109 (O_109,N_2893,N_2382);
and UO_110 (O_110,N_2791,N_2902);
nand UO_111 (O_111,N_2406,N_2568);
nor UO_112 (O_112,N_2467,N_2336);
and UO_113 (O_113,N_2739,N_2640);
nor UO_114 (O_114,N_2697,N_2339);
and UO_115 (O_115,N_2655,N_2633);
or UO_116 (O_116,N_2723,N_2542);
nor UO_117 (O_117,N_2933,N_2961);
nor UO_118 (O_118,N_2683,N_2301);
or UO_119 (O_119,N_2445,N_2427);
and UO_120 (O_120,N_2412,N_2276);
or UO_121 (O_121,N_2940,N_2518);
and UO_122 (O_122,N_2682,N_2960);
nand UO_123 (O_123,N_2758,N_2879);
and UO_124 (O_124,N_2733,N_2469);
nand UO_125 (O_125,N_2814,N_2964);
or UO_126 (O_126,N_2584,N_2513);
and UO_127 (O_127,N_2374,N_2886);
nand UO_128 (O_128,N_2546,N_2439);
nand UO_129 (O_129,N_2856,N_2563);
nand UO_130 (O_130,N_2692,N_2437);
and UO_131 (O_131,N_2585,N_2545);
or UO_132 (O_132,N_2387,N_2601);
and UO_133 (O_133,N_2315,N_2620);
xor UO_134 (O_134,N_2925,N_2965);
nor UO_135 (O_135,N_2631,N_2731);
or UO_136 (O_136,N_2591,N_2860);
and UO_137 (O_137,N_2430,N_2372);
or UO_138 (O_138,N_2846,N_2417);
or UO_139 (O_139,N_2671,N_2587);
or UO_140 (O_140,N_2713,N_2952);
xnor UO_141 (O_141,N_2290,N_2588);
xnor UO_142 (O_142,N_2254,N_2919);
or UO_143 (O_143,N_2784,N_2958);
and UO_144 (O_144,N_2646,N_2480);
nor UO_145 (O_145,N_2876,N_2678);
nor UO_146 (O_146,N_2603,N_2803);
nor UO_147 (O_147,N_2255,N_2963);
and UO_148 (O_148,N_2975,N_2362);
nor UO_149 (O_149,N_2801,N_2257);
or UO_150 (O_150,N_2780,N_2519);
nand UO_151 (O_151,N_2654,N_2647);
xor UO_152 (O_152,N_2901,N_2256);
and UO_153 (O_153,N_2809,N_2376);
nor UO_154 (O_154,N_2266,N_2865);
and UO_155 (O_155,N_2280,N_2938);
or UO_156 (O_156,N_2615,N_2852);
nor UO_157 (O_157,N_2527,N_2763);
xor UO_158 (O_158,N_2858,N_2870);
nor UO_159 (O_159,N_2735,N_2409);
nor UO_160 (O_160,N_2818,N_2533);
nand UO_161 (O_161,N_2543,N_2344);
nor UO_162 (O_162,N_2432,N_2753);
or UO_163 (O_163,N_2371,N_2540);
and UO_164 (O_164,N_2291,N_2461);
nand UO_165 (O_165,N_2267,N_2275);
nor UO_166 (O_166,N_2709,N_2281);
nand UO_167 (O_167,N_2896,N_2464);
nand UO_168 (O_168,N_2330,N_2804);
and UO_169 (O_169,N_2978,N_2343);
nor UO_170 (O_170,N_2997,N_2730);
or UO_171 (O_171,N_2622,N_2749);
nand UO_172 (O_172,N_2705,N_2329);
and UO_173 (O_173,N_2274,N_2738);
and UO_174 (O_174,N_2611,N_2436);
or UO_175 (O_175,N_2941,N_2841);
or UO_176 (O_176,N_2264,N_2327);
nand UO_177 (O_177,N_2651,N_2413);
xnor UO_178 (O_178,N_2431,N_2768);
nand UO_179 (O_179,N_2306,N_2386);
and UO_180 (O_180,N_2845,N_2410);
and UO_181 (O_181,N_2551,N_2286);
nor UO_182 (O_182,N_2995,N_2842);
xnor UO_183 (O_183,N_2862,N_2523);
nand UO_184 (O_184,N_2521,N_2657);
or UO_185 (O_185,N_2602,N_2750);
nor UO_186 (O_186,N_2293,N_2807);
nand UO_187 (O_187,N_2854,N_2408);
or UO_188 (O_188,N_2271,N_2373);
and UO_189 (O_189,N_2972,N_2252);
xor UO_190 (O_190,N_2967,N_2287);
xor UO_191 (O_191,N_2639,N_2986);
and UO_192 (O_192,N_2666,N_2261);
nor UO_193 (O_193,N_2531,N_2383);
or UO_194 (O_194,N_2617,N_2493);
or UO_195 (O_195,N_2945,N_2677);
and UO_196 (O_196,N_2440,N_2722);
and UO_197 (O_197,N_2970,N_2660);
nand UO_198 (O_198,N_2635,N_2547);
and UO_199 (O_199,N_2448,N_2714);
nand UO_200 (O_200,N_2923,N_2830);
or UO_201 (O_201,N_2912,N_2589);
and UO_202 (O_202,N_2345,N_2495);
nand UO_203 (O_203,N_2694,N_2983);
and UO_204 (O_204,N_2752,N_2619);
or UO_205 (O_205,N_2696,N_2459);
or UO_206 (O_206,N_2699,N_2379);
nand UO_207 (O_207,N_2643,N_2520);
nor UO_208 (O_208,N_2680,N_2392);
or UO_209 (O_209,N_2756,N_2285);
and UO_210 (O_210,N_2346,N_2398);
xor UO_211 (O_211,N_2857,N_2594);
and UO_212 (O_212,N_2561,N_2477);
or UO_213 (O_213,N_2979,N_2466);
or UO_214 (O_214,N_2501,N_2367);
or UO_215 (O_215,N_2593,N_2623);
and UO_216 (O_216,N_2562,N_2894);
and UO_217 (O_217,N_2898,N_2700);
nand UO_218 (O_218,N_2674,N_2312);
nor UO_219 (O_219,N_2884,N_2590);
nor UO_220 (O_220,N_2740,N_2351);
or UO_221 (O_221,N_2637,N_2727);
or UO_222 (O_222,N_2537,N_2377);
nand UO_223 (O_223,N_2303,N_2297);
and UO_224 (O_224,N_2444,N_2614);
nand UO_225 (O_225,N_2746,N_2721);
or UO_226 (O_226,N_2642,N_2875);
nand UO_227 (O_227,N_2323,N_2810);
xnor UO_228 (O_228,N_2258,N_2253);
xnor UO_229 (O_229,N_2318,N_2569);
nand UO_230 (O_230,N_2888,N_2302);
and UO_231 (O_231,N_2957,N_2710);
xnor UO_232 (O_232,N_2755,N_2484);
nor UO_233 (O_233,N_2843,N_2487);
or UO_234 (O_234,N_2554,N_2397);
nand UO_235 (O_235,N_2415,N_2381);
nor UO_236 (O_236,N_2762,N_2491);
nand UO_237 (O_237,N_2488,N_2322);
nor UO_238 (O_238,N_2337,N_2946);
and UO_239 (O_239,N_2859,N_2786);
xnor UO_240 (O_240,N_2300,N_2834);
nor UO_241 (O_241,N_2817,N_2821);
or UO_242 (O_242,N_2419,N_2921);
nand UO_243 (O_243,N_2878,N_2621);
and UO_244 (O_244,N_2511,N_2504);
or UO_245 (O_245,N_2636,N_2476);
and UO_246 (O_246,N_2510,N_2370);
xor UO_247 (O_247,N_2863,N_2483);
and UO_248 (O_248,N_2764,N_2904);
or UO_249 (O_249,N_2400,N_2799);
nor UO_250 (O_250,N_2684,N_2959);
or UO_251 (O_251,N_2396,N_2900);
and UO_252 (O_252,N_2416,N_2595);
nor UO_253 (O_253,N_2775,N_2905);
or UO_254 (O_254,N_2414,N_2872);
and UO_255 (O_255,N_2661,N_2906);
nor UO_256 (O_256,N_2512,N_2530);
nor UO_257 (O_257,N_2363,N_2296);
nand UO_258 (O_258,N_2284,N_2438);
or UO_259 (O_259,N_2481,N_2317);
and UO_260 (O_260,N_2260,N_2295);
and UO_261 (O_261,N_2892,N_2974);
or UO_262 (O_262,N_2790,N_2729);
nand UO_263 (O_263,N_2908,N_2827);
and UO_264 (O_264,N_2352,N_2855);
and UO_265 (O_265,N_2598,N_2435);
nand UO_266 (O_266,N_2420,N_2579);
nand UO_267 (O_267,N_2320,N_2951);
nor UO_268 (O_268,N_2822,N_2341);
xnor UO_269 (O_269,N_2625,N_2298);
or UO_270 (O_270,N_2653,N_2812);
and UO_271 (O_271,N_2485,N_2582);
nor UO_272 (O_272,N_2754,N_2669);
or UO_273 (O_273,N_2909,N_2333);
and UO_274 (O_274,N_2742,N_2450);
and UO_275 (O_275,N_2541,N_2380);
nor UO_276 (O_276,N_2676,N_2313);
nand UO_277 (O_277,N_2353,N_2874);
or UO_278 (O_278,N_2638,N_2456);
and UO_279 (O_279,N_2838,N_2282);
and UO_280 (O_280,N_2948,N_2744);
and UO_281 (O_281,N_2539,N_2745);
nor UO_282 (O_282,N_2581,N_2486);
or UO_283 (O_283,N_2848,N_2985);
nand UO_284 (O_284,N_2866,N_2328);
or UO_285 (O_285,N_2939,N_2342);
nand UO_286 (O_286,N_2806,N_2604);
nand UO_287 (O_287,N_2402,N_2618);
nor UO_288 (O_288,N_2433,N_2309);
nor UO_289 (O_289,N_2867,N_2823);
nor UO_290 (O_290,N_2883,N_2813);
and UO_291 (O_291,N_2917,N_2574);
xor UO_292 (O_292,N_2388,N_2292);
nor UO_293 (O_293,N_2304,N_2732);
or UO_294 (O_294,N_2981,N_2759);
xnor UO_295 (O_295,N_2662,N_2608);
and UO_296 (O_296,N_2776,N_2767);
xor UO_297 (O_297,N_2497,N_2576);
or UO_298 (O_298,N_2384,N_2792);
or UO_299 (O_299,N_2526,N_2811);
nand UO_300 (O_300,N_2553,N_2766);
xor UO_301 (O_301,N_2751,N_2994);
nand UO_302 (O_302,N_2449,N_2391);
nand UO_303 (O_303,N_2927,N_2769);
nand UO_304 (O_304,N_2360,N_2955);
and UO_305 (O_305,N_2839,N_2573);
nor UO_306 (O_306,N_2278,N_2357);
nor UO_307 (O_307,N_2600,N_2559);
nor UO_308 (O_308,N_2506,N_2369);
or UO_309 (O_309,N_2977,N_2624);
nand UO_310 (O_310,N_2897,N_2283);
and UO_311 (O_311,N_2716,N_2492);
nand UO_312 (O_312,N_2949,N_2701);
nand UO_313 (O_313,N_2273,N_2500);
or UO_314 (O_314,N_2688,N_2672);
or UO_315 (O_315,N_2265,N_2996);
or UO_316 (O_316,N_2508,N_2849);
xnor UO_317 (O_317,N_2425,N_2885);
and UO_318 (O_318,N_2976,N_2648);
and UO_319 (O_319,N_2928,N_2988);
nor UO_320 (O_320,N_2711,N_2443);
nor UO_321 (O_321,N_2605,N_2737);
nor UO_322 (O_322,N_2708,N_2356);
xnor UO_323 (O_323,N_2664,N_2861);
nor UO_324 (O_324,N_2442,N_2748);
or UO_325 (O_325,N_2361,N_2525);
and UO_326 (O_326,N_2549,N_2649);
nor UO_327 (O_327,N_2629,N_2460);
xnor UO_328 (O_328,N_2835,N_2837);
nand UO_329 (O_329,N_2468,N_2944);
and UO_330 (O_330,N_2250,N_2578);
xnor UO_331 (O_331,N_2820,N_2689);
or UO_332 (O_332,N_2509,N_2405);
nand UO_333 (O_333,N_2418,N_2685);
and UO_334 (O_334,N_2269,N_2982);
nor UO_335 (O_335,N_2942,N_2890);
and UO_336 (O_336,N_2675,N_2989);
nor UO_337 (O_337,N_2802,N_2441);
nor UO_338 (O_338,N_2517,N_2423);
nand UO_339 (O_339,N_2747,N_2871);
and UO_340 (O_340,N_2407,N_2873);
nand UO_341 (O_341,N_2895,N_2840);
or UO_342 (O_342,N_2828,N_2797);
xor UO_343 (O_343,N_2966,N_2586);
nand UO_344 (O_344,N_2704,N_2819);
xnor UO_345 (O_345,N_2534,N_2881);
and UO_346 (O_346,N_2698,N_2627);
and UO_347 (O_347,N_2761,N_2824);
nor UO_348 (O_348,N_2596,N_2592);
and UO_349 (O_349,N_2524,N_2717);
or UO_350 (O_350,N_2707,N_2385);
and UO_351 (O_351,N_2929,N_2924);
nor UO_352 (O_352,N_2475,N_2903);
nor UO_353 (O_353,N_2522,N_2499);
nor UO_354 (O_354,N_2272,N_2916);
or UO_355 (O_355,N_2325,N_2741);
and UO_356 (O_356,N_2503,N_2455);
or UO_357 (O_357,N_2515,N_2548);
nand UO_358 (O_358,N_2564,N_2610);
nand UO_359 (O_359,N_2626,N_2935);
nor UO_360 (O_360,N_2609,N_2816);
or UO_361 (O_361,N_2930,N_2783);
or UO_362 (O_362,N_2789,N_2969);
or UO_363 (O_363,N_2971,N_2489);
or UO_364 (O_364,N_2850,N_2956);
or UO_365 (O_365,N_2334,N_2968);
or UO_366 (O_366,N_2634,N_2720);
nand UO_367 (O_367,N_2779,N_2932);
nor UO_368 (O_368,N_2516,N_2324);
or UO_369 (O_369,N_2536,N_2918);
and UO_370 (O_370,N_2771,N_2934);
nand UO_371 (O_371,N_2289,N_2310);
or UO_372 (O_372,N_2558,N_2882);
and UO_373 (O_373,N_2778,N_2474);
nand UO_374 (O_374,N_2457,N_2899);
and UO_375 (O_375,N_2722,N_2449);
and UO_376 (O_376,N_2711,N_2320);
nor UO_377 (O_377,N_2414,N_2260);
xor UO_378 (O_378,N_2314,N_2935);
nor UO_379 (O_379,N_2581,N_2467);
and UO_380 (O_380,N_2299,N_2480);
and UO_381 (O_381,N_2874,N_2341);
nor UO_382 (O_382,N_2679,N_2614);
nor UO_383 (O_383,N_2522,N_2420);
and UO_384 (O_384,N_2447,N_2683);
nand UO_385 (O_385,N_2732,N_2445);
nand UO_386 (O_386,N_2443,N_2624);
nand UO_387 (O_387,N_2913,N_2316);
or UO_388 (O_388,N_2685,N_2701);
and UO_389 (O_389,N_2855,N_2431);
nor UO_390 (O_390,N_2889,N_2986);
nand UO_391 (O_391,N_2914,N_2334);
nor UO_392 (O_392,N_2760,N_2339);
or UO_393 (O_393,N_2646,N_2803);
and UO_394 (O_394,N_2848,N_2722);
and UO_395 (O_395,N_2953,N_2747);
and UO_396 (O_396,N_2426,N_2538);
and UO_397 (O_397,N_2620,N_2601);
or UO_398 (O_398,N_2956,N_2360);
xnor UO_399 (O_399,N_2741,N_2299);
nand UO_400 (O_400,N_2307,N_2594);
and UO_401 (O_401,N_2470,N_2328);
and UO_402 (O_402,N_2428,N_2791);
and UO_403 (O_403,N_2803,N_2835);
or UO_404 (O_404,N_2515,N_2918);
or UO_405 (O_405,N_2782,N_2809);
nand UO_406 (O_406,N_2662,N_2330);
and UO_407 (O_407,N_2706,N_2482);
nand UO_408 (O_408,N_2504,N_2722);
or UO_409 (O_409,N_2779,N_2372);
or UO_410 (O_410,N_2513,N_2465);
or UO_411 (O_411,N_2430,N_2481);
or UO_412 (O_412,N_2399,N_2426);
nand UO_413 (O_413,N_2713,N_2873);
nor UO_414 (O_414,N_2658,N_2738);
and UO_415 (O_415,N_2308,N_2926);
and UO_416 (O_416,N_2451,N_2615);
nor UO_417 (O_417,N_2650,N_2942);
nand UO_418 (O_418,N_2704,N_2562);
or UO_419 (O_419,N_2577,N_2937);
nor UO_420 (O_420,N_2485,N_2348);
nand UO_421 (O_421,N_2781,N_2976);
nand UO_422 (O_422,N_2260,N_2931);
xor UO_423 (O_423,N_2801,N_2696);
xor UO_424 (O_424,N_2698,N_2908);
or UO_425 (O_425,N_2307,N_2363);
or UO_426 (O_426,N_2342,N_2947);
nand UO_427 (O_427,N_2305,N_2693);
or UO_428 (O_428,N_2849,N_2429);
nand UO_429 (O_429,N_2456,N_2704);
or UO_430 (O_430,N_2969,N_2540);
xnor UO_431 (O_431,N_2573,N_2253);
nor UO_432 (O_432,N_2513,N_2880);
and UO_433 (O_433,N_2719,N_2784);
xnor UO_434 (O_434,N_2707,N_2355);
nor UO_435 (O_435,N_2549,N_2879);
nand UO_436 (O_436,N_2599,N_2864);
nor UO_437 (O_437,N_2466,N_2397);
nor UO_438 (O_438,N_2868,N_2428);
and UO_439 (O_439,N_2515,N_2695);
and UO_440 (O_440,N_2507,N_2368);
nand UO_441 (O_441,N_2405,N_2649);
or UO_442 (O_442,N_2482,N_2885);
and UO_443 (O_443,N_2625,N_2912);
or UO_444 (O_444,N_2787,N_2695);
or UO_445 (O_445,N_2668,N_2294);
nor UO_446 (O_446,N_2488,N_2415);
or UO_447 (O_447,N_2684,N_2604);
or UO_448 (O_448,N_2969,N_2336);
or UO_449 (O_449,N_2368,N_2993);
nor UO_450 (O_450,N_2609,N_2668);
and UO_451 (O_451,N_2859,N_2997);
and UO_452 (O_452,N_2931,N_2424);
and UO_453 (O_453,N_2340,N_2721);
nor UO_454 (O_454,N_2251,N_2802);
and UO_455 (O_455,N_2654,N_2560);
nand UO_456 (O_456,N_2827,N_2959);
nand UO_457 (O_457,N_2456,N_2420);
and UO_458 (O_458,N_2470,N_2894);
nor UO_459 (O_459,N_2338,N_2493);
and UO_460 (O_460,N_2379,N_2583);
nor UO_461 (O_461,N_2419,N_2699);
or UO_462 (O_462,N_2759,N_2660);
nand UO_463 (O_463,N_2888,N_2890);
xor UO_464 (O_464,N_2862,N_2744);
or UO_465 (O_465,N_2261,N_2826);
nand UO_466 (O_466,N_2723,N_2782);
nand UO_467 (O_467,N_2558,N_2495);
nor UO_468 (O_468,N_2747,N_2318);
or UO_469 (O_469,N_2870,N_2297);
or UO_470 (O_470,N_2313,N_2299);
nand UO_471 (O_471,N_2587,N_2552);
nand UO_472 (O_472,N_2867,N_2662);
nor UO_473 (O_473,N_2379,N_2834);
nand UO_474 (O_474,N_2806,N_2311);
nor UO_475 (O_475,N_2470,N_2346);
and UO_476 (O_476,N_2719,N_2299);
nand UO_477 (O_477,N_2375,N_2839);
or UO_478 (O_478,N_2434,N_2833);
xnor UO_479 (O_479,N_2367,N_2274);
nand UO_480 (O_480,N_2771,N_2329);
nor UO_481 (O_481,N_2547,N_2882);
nand UO_482 (O_482,N_2955,N_2812);
nand UO_483 (O_483,N_2864,N_2282);
nor UO_484 (O_484,N_2618,N_2397);
nor UO_485 (O_485,N_2282,N_2287);
nand UO_486 (O_486,N_2427,N_2361);
nand UO_487 (O_487,N_2447,N_2949);
xor UO_488 (O_488,N_2533,N_2936);
and UO_489 (O_489,N_2857,N_2548);
xor UO_490 (O_490,N_2378,N_2525);
nor UO_491 (O_491,N_2663,N_2832);
and UO_492 (O_492,N_2755,N_2775);
nand UO_493 (O_493,N_2943,N_2826);
and UO_494 (O_494,N_2674,N_2704);
xor UO_495 (O_495,N_2982,N_2556);
nand UO_496 (O_496,N_2333,N_2997);
or UO_497 (O_497,N_2334,N_2896);
nor UO_498 (O_498,N_2814,N_2995);
nand UO_499 (O_499,N_2681,N_2328);
endmodule