module basic_3000_30000_3500_6_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
and U0 (N_0,In_1702,In_625);
xnor U1 (N_1,In_2236,In_1695);
nor U2 (N_2,In_708,In_346);
xnor U3 (N_3,In_2631,In_1763);
or U4 (N_4,In_55,In_282);
or U5 (N_5,In_1304,In_1102);
xor U6 (N_6,In_677,In_1607);
nand U7 (N_7,In_2324,In_1436);
and U8 (N_8,In_1205,In_2347);
nor U9 (N_9,In_1968,In_256);
nand U10 (N_10,In_1747,In_2366);
xnor U11 (N_11,In_1913,In_787);
xor U12 (N_12,In_74,In_2990);
nor U13 (N_13,In_1474,In_1228);
xnor U14 (N_14,In_1641,In_2859);
or U15 (N_15,In_725,In_398);
or U16 (N_16,In_60,In_2800);
or U17 (N_17,In_2734,In_2160);
nand U18 (N_18,In_443,In_185);
nor U19 (N_19,In_1438,In_2280);
or U20 (N_20,In_1579,In_1025);
and U21 (N_21,In_1046,In_1110);
nor U22 (N_22,In_318,In_199);
nand U23 (N_23,In_2822,In_320);
and U24 (N_24,In_959,In_837);
nor U25 (N_25,In_1745,In_2071);
and U26 (N_26,In_2902,In_241);
nor U27 (N_27,In_2300,In_2455);
xnor U28 (N_28,In_802,In_1178);
nor U29 (N_29,In_2422,In_757);
nand U30 (N_30,In_2174,In_2931);
or U31 (N_31,In_1485,In_565);
xnor U32 (N_32,In_2718,In_425);
or U33 (N_33,In_1168,In_2289);
nor U34 (N_34,In_1152,In_184);
xor U35 (N_35,In_975,In_2016);
nand U36 (N_36,In_2814,In_632);
nand U37 (N_37,In_659,In_2510);
and U38 (N_38,In_434,In_807);
nor U39 (N_39,In_2475,In_561);
nor U40 (N_40,In_1639,In_2843);
or U41 (N_41,In_806,In_2942);
and U42 (N_42,In_2924,In_2437);
nor U43 (N_43,In_556,In_675);
xnor U44 (N_44,In_2484,In_712);
nor U45 (N_45,In_2098,In_2737);
xnor U46 (N_46,In_624,In_2257);
or U47 (N_47,In_1016,In_2765);
xnor U48 (N_48,In_224,In_2348);
nor U49 (N_49,In_347,In_2464);
and U50 (N_50,In_1634,In_810);
nor U51 (N_51,In_2959,In_2657);
nor U52 (N_52,In_2430,In_2781);
or U53 (N_53,In_707,In_1728);
and U54 (N_54,In_2395,In_1848);
and U55 (N_55,In_731,In_451);
or U56 (N_56,In_2057,In_843);
and U57 (N_57,In_619,In_2291);
xor U58 (N_58,In_778,In_844);
xnor U59 (N_59,In_2982,In_1940);
and U60 (N_60,In_824,In_2415);
nor U61 (N_61,In_924,In_1213);
nor U62 (N_62,In_2136,In_1788);
and U63 (N_63,In_2222,In_2590);
xor U64 (N_64,In_700,In_1708);
xnor U65 (N_65,In_296,In_1461);
xor U66 (N_66,In_1609,In_1533);
nor U67 (N_67,In_2679,In_1699);
or U68 (N_68,In_96,In_1189);
or U69 (N_69,In_1212,In_1166);
or U70 (N_70,In_121,In_688);
nand U71 (N_71,In_2031,In_1403);
nand U72 (N_72,In_156,In_227);
nor U73 (N_73,In_2082,In_541);
and U74 (N_74,In_2846,In_2500);
and U75 (N_75,In_1693,In_936);
and U76 (N_76,In_1735,In_2709);
nor U77 (N_77,In_2583,In_1587);
and U78 (N_78,In_2239,In_3);
nand U79 (N_79,In_1247,In_2404);
and U80 (N_80,In_498,In_2889);
or U81 (N_81,In_1667,In_995);
or U82 (N_82,In_1821,In_1307);
and U83 (N_83,In_1039,In_20);
xor U84 (N_84,In_140,In_696);
and U85 (N_85,In_1059,In_1749);
nor U86 (N_86,In_506,In_2360);
xor U87 (N_87,In_2490,In_1859);
nand U88 (N_88,In_171,In_883);
and U89 (N_89,In_2162,In_820);
nand U90 (N_90,In_940,In_1395);
and U91 (N_91,In_2084,In_1423);
and U92 (N_92,In_1376,In_59);
or U93 (N_93,In_2904,In_671);
or U94 (N_94,In_2002,In_2301);
xnor U95 (N_95,In_413,In_2813);
and U96 (N_96,In_2454,In_1548);
nor U97 (N_97,In_934,In_2027);
xnor U98 (N_98,In_373,In_190);
or U99 (N_99,In_996,In_2052);
and U100 (N_100,In_1377,In_2024);
xor U101 (N_101,In_962,In_1737);
and U102 (N_102,In_1754,In_1818);
xnor U103 (N_103,In_2154,In_2155);
and U104 (N_104,In_2453,In_1099);
or U105 (N_105,In_1345,In_1159);
or U106 (N_106,In_2327,In_1200);
nor U107 (N_107,In_1922,In_1233);
or U108 (N_108,In_312,In_1620);
or U109 (N_109,In_1909,In_658);
nor U110 (N_110,In_1774,In_31);
and U111 (N_111,In_2400,In_1907);
nand U112 (N_112,In_1912,In_1799);
nor U113 (N_113,In_339,In_1540);
xor U114 (N_114,In_2693,In_2858);
nand U115 (N_115,In_1464,In_875);
and U116 (N_116,In_1545,In_1396);
and U117 (N_117,In_454,In_931);
xnor U118 (N_118,In_1606,In_873);
nand U119 (N_119,In_1574,In_393);
or U120 (N_120,In_238,In_108);
and U121 (N_121,In_1089,In_862);
xnor U122 (N_122,In_1694,In_1479);
and U123 (N_123,In_1552,In_1096);
nand U124 (N_124,In_2887,In_2440);
nand U125 (N_125,In_179,In_402);
xnor U126 (N_126,In_956,In_362);
nand U127 (N_127,In_463,In_419);
or U128 (N_128,In_1585,In_584);
xnor U129 (N_129,In_750,In_775);
nor U130 (N_130,In_2492,In_276);
and U131 (N_131,In_642,In_2479);
nand U132 (N_132,In_1051,In_1174);
and U133 (N_133,In_2288,In_1342);
nand U134 (N_134,In_877,In_1635);
or U135 (N_135,In_1351,In_2383);
or U136 (N_136,In_1203,In_2608);
nand U137 (N_137,In_2518,In_304);
nand U138 (N_138,In_82,In_2939);
xnor U139 (N_139,In_2661,In_2854);
nand U140 (N_140,In_1910,In_702);
or U141 (N_141,In_2164,In_1865);
nand U142 (N_142,In_2549,In_2135);
nand U143 (N_143,In_287,In_508);
xnor U144 (N_144,In_1581,In_247);
or U145 (N_145,In_1452,In_1306);
and U146 (N_146,In_2771,In_1951);
xnor U147 (N_147,In_2306,In_2261);
or U148 (N_148,In_1067,In_1108);
xor U149 (N_149,In_1300,In_2864);
or U150 (N_150,In_472,In_2234);
or U151 (N_151,In_1375,In_131);
nand U152 (N_152,In_485,In_1923);
nor U153 (N_153,In_2824,In_360);
xnor U154 (N_154,In_1294,In_804);
nor U155 (N_155,In_2915,In_1141);
or U156 (N_156,In_1497,In_1723);
or U157 (N_157,In_966,In_583);
nand U158 (N_158,In_1807,In_92);
xnor U159 (N_159,In_1330,In_717);
xor U160 (N_160,In_32,In_1952);
nor U161 (N_161,In_601,In_795);
and U162 (N_162,In_2838,In_706);
nor U163 (N_163,In_1070,In_1144);
and U164 (N_164,In_912,In_1467);
nor U165 (N_165,In_1341,In_1142);
nand U166 (N_166,In_1899,In_621);
nor U167 (N_167,In_1235,In_228);
or U168 (N_168,In_1457,In_2506);
or U169 (N_169,In_2782,In_1008);
and U170 (N_170,In_456,In_16);
nand U171 (N_171,In_311,In_1499);
xnor U172 (N_172,In_2451,In_4);
or U173 (N_173,In_315,In_1369);
or U174 (N_174,In_1543,In_1275);
nand U175 (N_175,In_2157,In_2964);
xor U176 (N_176,In_774,In_1249);
or U177 (N_177,In_1622,In_656);
nand U178 (N_178,In_723,In_2273);
and U179 (N_179,In_1888,In_2783);
and U180 (N_180,In_1947,In_166);
or U181 (N_181,In_1426,In_721);
nand U182 (N_182,In_2739,In_1179);
xnor U183 (N_183,In_78,In_2857);
nor U184 (N_184,In_1934,In_471);
xnor U185 (N_185,In_604,In_2978);
nor U186 (N_186,In_1626,In_466);
xor U187 (N_187,In_2028,In_2791);
nor U188 (N_188,In_520,In_79);
and U189 (N_189,In_2353,In_1315);
and U190 (N_190,In_2703,In_2805);
or U191 (N_191,In_2574,In_2248);
nor U192 (N_192,In_646,In_193);
and U193 (N_193,In_2065,In_816);
nor U194 (N_194,In_2853,In_2364);
xnor U195 (N_195,In_1712,In_1297);
or U196 (N_196,In_1273,In_1534);
and U197 (N_197,In_453,In_490);
and U198 (N_198,In_1822,In_273);
and U199 (N_199,In_474,In_1125);
and U200 (N_200,In_2134,In_662);
nor U201 (N_201,In_2312,In_2972);
and U202 (N_202,In_751,In_1324);
nand U203 (N_203,In_309,In_1811);
or U204 (N_204,In_1107,In_1999);
nor U205 (N_205,In_1379,In_1362);
and U206 (N_206,In_122,In_1953);
nand U207 (N_207,In_730,In_2777);
and U208 (N_208,In_2138,In_2578);
xnor U209 (N_209,In_2756,In_1729);
nor U210 (N_210,In_1224,In_1253);
xnor U211 (N_211,In_1709,In_57);
nand U212 (N_212,In_2705,In_35);
nor U213 (N_213,In_1684,In_2473);
or U214 (N_214,In_316,In_1941);
and U215 (N_215,In_2252,In_1796);
or U216 (N_216,In_1834,In_441);
xnor U217 (N_217,In_2808,In_1828);
nand U218 (N_218,In_831,In_1276);
and U219 (N_219,In_1777,In_1883);
and U220 (N_220,In_1789,In_1531);
and U221 (N_221,In_371,In_1785);
nand U222 (N_222,In_947,In_2670);
nand U223 (N_223,In_667,In_2930);
or U224 (N_224,In_1238,In_2770);
xor U225 (N_225,In_1155,In_803);
nand U226 (N_226,In_2113,In_344);
and U227 (N_227,In_701,In_209);
or U228 (N_228,In_1549,In_827);
xnor U229 (N_229,In_2104,In_2573);
and U230 (N_230,In_1138,In_2097);
nor U231 (N_231,In_1630,In_1407);
nor U232 (N_232,In_1500,In_1658);
or U233 (N_233,In_1528,In_2358);
nand U234 (N_234,In_1193,In_1047);
and U235 (N_235,In_435,In_1196);
or U236 (N_236,In_835,In_697);
nand U237 (N_237,In_181,In_2220);
and U238 (N_238,In_2584,In_777);
nand U239 (N_239,In_1041,In_2493);
or U240 (N_240,In_1456,In_80);
nor U241 (N_241,In_633,In_856);
and U242 (N_242,In_1298,In_1894);
nor U243 (N_243,In_2890,In_2543);
nand U244 (N_244,In_1845,In_1498);
nand U245 (N_245,In_403,In_1425);
nand U246 (N_246,In_997,In_1588);
and U247 (N_247,In_892,In_2431);
nand U248 (N_248,In_1455,In_1829);
nand U249 (N_249,In_1757,In_2319);
and U250 (N_250,In_383,In_1433);
xnor U251 (N_251,In_994,In_400);
nand U252 (N_252,In_2448,In_1553);
nor U253 (N_253,In_1245,In_978);
and U254 (N_254,In_1009,In_1254);
or U255 (N_255,In_1242,In_981);
nand U256 (N_256,In_1378,In_879);
nand U257 (N_257,In_2512,In_1804);
nand U258 (N_258,In_1327,In_1954);
or U259 (N_259,In_2019,In_1871);
nor U260 (N_260,In_889,In_2845);
or U261 (N_261,In_14,In_173);
nor U262 (N_262,In_705,In_1043);
xor U263 (N_263,In_2042,In_977);
or U264 (N_264,In_547,In_1223);
or U265 (N_265,In_1098,In_2260);
nor U266 (N_266,In_1252,In_1201);
nand U267 (N_267,In_202,In_2375);
xor U268 (N_268,In_781,In_2747);
xor U269 (N_269,In_1157,In_72);
and U270 (N_270,In_1838,In_176);
nand U271 (N_271,In_390,In_1270);
nor U272 (N_272,In_1511,In_755);
nand U273 (N_273,In_305,In_524);
nor U274 (N_274,In_1858,In_922);
nand U275 (N_275,In_1786,In_1578);
or U276 (N_276,In_2172,In_2507);
and U277 (N_277,In_175,In_2152);
nor U278 (N_278,In_2898,In_192);
nand U279 (N_279,In_372,In_457);
nor U280 (N_280,In_2109,In_2403);
xor U281 (N_281,In_1901,In_1109);
and U282 (N_282,In_2497,In_615);
xor U283 (N_283,In_481,In_2515);
xor U284 (N_284,In_1759,In_1240);
or U285 (N_285,In_2610,In_1668);
xor U286 (N_286,In_690,In_1033);
or U287 (N_287,In_370,In_1628);
nor U288 (N_288,In_2489,In_2798);
xnor U289 (N_289,In_2390,In_2212);
or U290 (N_290,In_1819,In_380);
or U291 (N_291,In_1536,In_265);
and U292 (N_292,In_2242,In_2246);
xor U293 (N_293,In_1349,In_617);
nor U294 (N_294,In_1840,In_1082);
nand U295 (N_295,In_2,In_507);
or U296 (N_296,In_142,In_1257);
or U297 (N_297,In_2556,In_2208);
and U298 (N_298,In_470,In_1556);
nand U299 (N_299,In_2401,In_1022);
xor U300 (N_300,In_1602,In_2710);
nor U301 (N_301,In_1134,In_871);
nor U302 (N_302,In_2381,In_1830);
or U303 (N_303,In_1244,In_2377);
nor U304 (N_304,In_2344,In_1382);
xor U305 (N_305,In_1,In_2803);
nor U306 (N_306,In_2250,In_447);
nand U307 (N_307,In_118,In_789);
nor U308 (N_308,In_2903,In_2046);
nor U309 (N_309,In_882,In_1598);
and U310 (N_310,In_1736,In_1398);
xnor U311 (N_311,In_292,In_2056);
and U312 (N_312,In_2667,In_973);
nand U313 (N_313,In_2474,In_1592);
or U314 (N_314,In_2732,In_965);
xor U315 (N_315,In_814,In_1064);
nand U316 (N_316,In_2165,In_66);
or U317 (N_317,In_613,In_2588);
nor U318 (N_318,In_575,In_2775);
or U319 (N_319,In_594,In_381);
and U320 (N_320,In_1217,In_2259);
nor U321 (N_321,In_2876,In_2255);
xnor U322 (N_322,In_1226,In_2175);
xnor U323 (N_323,In_2374,In_1204);
xnor U324 (N_324,In_2335,In_1373);
or U325 (N_325,In_1880,In_221);
and U326 (N_326,In_2759,In_1676);
nor U327 (N_327,In_939,In_2856);
nand U328 (N_328,In_2491,In_772);
xor U329 (N_329,In_10,In_2700);
nand U330 (N_330,In_1651,In_351);
nor U331 (N_331,In_2677,In_1250);
nand U332 (N_332,In_1558,In_1363);
nor U333 (N_333,In_2883,In_2309);
or U334 (N_334,In_1529,In_2354);
and U335 (N_335,In_489,In_710);
and U336 (N_336,In_825,In_1271);
and U337 (N_337,In_401,In_155);
xnor U338 (N_338,In_2087,In_2593);
nand U339 (N_339,In_1490,In_2606);
and U340 (N_340,In_1768,In_350);
nand U341 (N_341,In_773,In_2695);
nor U342 (N_342,In_1615,In_25);
and U343 (N_343,In_2287,In_1798);
and U344 (N_344,In_2659,In_429);
or U345 (N_345,In_1586,In_2402);
nor U346 (N_346,In_845,In_426);
or U347 (N_347,In_357,In_955);
and U348 (N_348,In_1756,In_2414);
xnor U349 (N_349,In_1026,In_2412);
or U350 (N_350,In_68,In_2743);
nor U351 (N_351,In_1508,In_1680);
xnor U352 (N_352,In_452,In_1654);
nand U353 (N_353,In_890,In_382);
and U354 (N_354,In_1766,In_2086);
and U355 (N_355,In_124,In_1573);
and U356 (N_356,In_1290,In_93);
nand U357 (N_357,In_1751,In_146);
and U358 (N_358,In_1931,In_993);
nand U359 (N_359,In_805,In_2308);
nand U360 (N_360,In_1862,In_2825);
or U361 (N_361,In_2819,In_98);
nand U362 (N_362,In_2616,In_110);
or U363 (N_363,In_1955,In_321);
xnor U364 (N_364,In_1713,In_48);
xnor U365 (N_365,In_740,In_1846);
nand U366 (N_366,In_2298,In_71);
nor U367 (N_367,In_726,In_1429);
and U368 (N_368,In_150,In_2622);
or U369 (N_369,In_953,In_2350);
xor U370 (N_370,In_1019,In_41);
nor U371 (N_371,In_254,In_249);
or U372 (N_372,In_281,In_2070);
or U373 (N_373,In_958,In_2944);
nand U374 (N_374,In_987,In_512);
nand U375 (N_375,In_2329,In_162);
and U376 (N_376,In_1617,In_1328);
or U377 (N_377,In_2881,In_2371);
or U378 (N_378,In_1946,In_1949);
and U379 (N_379,In_898,In_609);
and U380 (N_380,In_125,In_2839);
nor U381 (N_381,In_216,In_1738);
xnor U382 (N_382,In_1510,In_572);
nor U383 (N_383,In_2158,In_1463);
nor U384 (N_384,In_2468,In_2014);
xnor U385 (N_385,In_670,In_2177);
or U386 (N_386,In_148,In_1715);
nand U387 (N_387,In_2315,In_1052);
nor U388 (N_388,In_1104,In_1430);
or U389 (N_389,In_1685,In_486);
or U390 (N_390,In_1401,In_2276);
xor U391 (N_391,In_2282,In_2950);
or U392 (N_392,In_1895,In_1222);
and U393 (N_393,In_1655,In_2176);
or U394 (N_394,In_2173,In_274);
nand U395 (N_395,In_2551,In_2483);
and U396 (N_396,In_1594,In_1225);
or U397 (N_397,In_1515,In_1760);
nand U398 (N_398,In_830,In_544);
xnor U399 (N_399,In_290,In_1000);
or U400 (N_400,In_523,In_909);
nor U401 (N_401,In_2202,In_2139);
nand U402 (N_402,In_1562,In_1197);
nand U403 (N_403,In_396,In_2534);
and U404 (N_404,In_1465,In_2907);
nand U405 (N_405,In_2116,In_151);
nor U406 (N_406,In_2830,In_170);
and U407 (N_407,In_200,In_1950);
or U408 (N_408,In_2411,In_289);
and U409 (N_409,In_349,In_2762);
or U410 (N_410,In_676,In_1388);
nand U411 (N_411,In_678,In_186);
or U412 (N_412,In_986,In_2832);
xor U413 (N_413,In_138,In_1727);
or U414 (N_414,In_735,In_285);
xor U415 (N_415,In_1336,In_1652);
and U416 (N_416,In_1001,In_2586);
nor U417 (N_417,In_135,In_1487);
nand U418 (N_418,In_460,In_30);
nor U419 (N_419,In_2251,In_1721);
and U420 (N_420,In_2126,In_2117);
nand U421 (N_421,In_2124,In_891);
or U422 (N_422,In_2630,In_720);
nand U423 (N_423,In_2674,In_468);
and U424 (N_424,In_727,In_1672);
or U425 (N_425,In_1967,In_1793);
or U426 (N_426,In_188,In_2744);
and U427 (N_427,In_1177,In_433);
or U428 (N_428,In_2766,In_2788);
and U429 (N_429,In_2977,In_2339);
nand U430 (N_430,In_355,In_2912);
nand U431 (N_431,In_1210,In_2773);
nor U432 (N_432,In_1394,In_1677);
nand U433 (N_433,In_102,In_2432);
nand U434 (N_434,In_644,In_2081);
nand U435 (N_435,In_2682,In_1218);
xnor U436 (N_436,In_2628,In_2882);
xnor U437 (N_437,In_203,In_1664);
nor U438 (N_438,In_1391,In_2449);
and U439 (N_439,In_944,In_872);
and U440 (N_440,In_858,In_1701);
nor U441 (N_441,In_2062,In_598);
nor U442 (N_442,In_1291,In_2672);
nor U443 (N_443,In_1525,In_1933);
xnor U444 (N_444,In_2753,In_1824);
or U445 (N_445,In_1970,In_2342);
and U446 (N_446,In_2382,In_1380);
xor U447 (N_447,In_24,In_1539);
or U448 (N_448,In_2796,In_2642);
nor U449 (N_449,In_2877,In_386);
xnor U450 (N_450,In_376,In_263);
nand U451 (N_451,In_1086,In_709);
nor U452 (N_452,In_1502,In_1886);
xnor U453 (N_453,In_1310,In_999);
nand U454 (N_454,In_2852,In_913);
nand U455 (N_455,In_2511,In_1741);
or U456 (N_456,In_1140,In_923);
or U457 (N_457,In_2643,In_2544);
and U458 (N_458,In_963,In_1803);
or U459 (N_459,In_846,In_2372);
nand U460 (N_460,In_519,In_2336);
or U461 (N_461,In_1454,In_2570);
nor U462 (N_462,In_914,In_2571);
nor U463 (N_463,In_1151,In_2201);
or U464 (N_464,In_1717,In_2069);
xor U465 (N_465,In_219,In_1640);
nand U466 (N_466,In_2923,In_1986);
and U467 (N_467,In_217,In_636);
or U468 (N_468,In_2899,In_2206);
or U469 (N_469,In_2909,In_492);
nor U470 (N_470,In_1800,In_817);
nand U471 (N_471,In_933,In_136);
nor U472 (N_472,In_1903,In_1389);
and U473 (N_473,In_503,In_516);
nand U474 (N_474,In_2987,In_2613);
and U475 (N_475,In_2045,In_374);
or U476 (N_476,In_2524,In_1018);
or U477 (N_477,In_1669,In_552);
nor U478 (N_478,In_2970,In_1877);
nor U479 (N_479,In_724,In_2817);
nor U480 (N_480,In_743,In_2801);
xnor U481 (N_481,In_2235,In_2247);
xnor U482 (N_482,In_2150,In_666);
or U483 (N_483,In_1572,In_2438);
nor U484 (N_484,In_2740,In_611);
nor U485 (N_485,In_2776,In_1136);
or U486 (N_486,In_2078,In_1814);
nor U487 (N_487,In_527,In_39);
nor U488 (N_488,In_300,In_1942);
nor U489 (N_489,In_534,In_13);
or U490 (N_490,In_1753,In_1314);
nor U491 (N_491,In_1731,In_1266);
xnor U492 (N_492,In_1995,In_1841);
nand U493 (N_493,In_2513,In_45);
and U494 (N_494,In_1770,In_2209);
and U495 (N_495,In_405,In_1567);
nand U496 (N_496,In_2553,In_1397);
or U497 (N_497,In_1893,In_2600);
and U498 (N_498,In_2331,In_1471);
xnor U499 (N_499,In_1591,In_1478);
nor U500 (N_500,In_1921,In_1435);
or U501 (N_501,In_64,In_2271);
xor U502 (N_502,In_2216,In_655);
and U503 (N_503,In_1347,In_2582);
nand U504 (N_504,In_38,In_368);
nand U505 (N_505,In_264,In_540);
or U506 (N_506,In_478,In_1065);
nand U507 (N_507,In_1809,In_284);
xnor U508 (N_508,In_1817,In_2170);
and U509 (N_509,In_1897,In_1643);
nor U510 (N_510,In_2860,In_1147);
nand U511 (N_511,In_1126,In_1413);
nand U512 (N_512,In_907,In_900);
nor U513 (N_513,In_1083,In_2316);
nand U514 (N_514,In_2343,In_1480);
nand U515 (N_515,In_2519,In_2279);
xnor U516 (N_516,In_797,In_1679);
or U517 (N_517,In_1343,In_2863);
nor U518 (N_518,In_2146,In_44);
xor U519 (N_519,In_1990,In_2598);
or U520 (N_520,In_1192,In_246);
nand U521 (N_521,In_2665,In_853);
and U522 (N_522,In_1408,In_799);
nand U523 (N_523,In_2419,In_744);
nand U524 (N_524,In_50,In_1501);
nor U525 (N_525,In_448,In_849);
nand U526 (N_526,In_2692,In_1524);
or U527 (N_527,In_2955,In_1227);
or U528 (N_528,In_1614,In_1150);
xor U529 (N_529,In_1782,In_715);
xnor U530 (N_530,In_571,In_1980);
or U531 (N_531,In_1441,In_1936);
xor U532 (N_532,In_607,In_2960);
nand U533 (N_533,In_1207,In_2802);
or U534 (N_534,In_2595,In_437);
nand U535 (N_535,In_2458,In_1028);
or U536 (N_536,In_813,In_301);
nor U537 (N_537,In_2376,In_1687);
nor U538 (N_538,In_1881,In_255);
and U539 (N_539,In_2967,In_1085);
xor U540 (N_540,In_1139,In_1992);
xnor U541 (N_541,In_2660,In_1905);
xor U542 (N_542,In_2694,In_1123);
or U543 (N_543,In_1625,In_1554);
nor U544 (N_544,In_2199,In_1837);
nand U545 (N_545,In_2894,In_1994);
nor U546 (N_546,In_364,In_293);
xnor U547 (N_547,In_243,In_1440);
and U548 (N_548,In_1367,In_1755);
nand U549 (N_549,In_848,In_412);
nand U550 (N_550,In_1977,In_2203);
or U551 (N_551,In_2467,In_828);
and U552 (N_552,In_46,In_1393);
nand U553 (N_553,In_766,In_2159);
or U554 (N_554,In_167,In_197);
xnor U555 (N_555,In_1311,In_1122);
xnor U556 (N_556,In_342,In_1948);
xor U557 (N_557,In_2685,In_183);
nor U558 (N_558,In_2048,In_1808);
xor U559 (N_559,In_432,In_573);
nor U560 (N_560,In_796,In_1078);
nand U561 (N_561,In_2968,In_2131);
nor U562 (N_562,In_563,In_988);
xor U563 (N_563,In_214,In_7);
nand U564 (N_564,In_2962,In_729);
or U565 (N_565,In_1521,In_2644);
nor U566 (N_566,In_1779,In_286);
nor U567 (N_567,In_1621,In_857);
nand U568 (N_568,In_2362,In_2445);
or U569 (N_569,In_1509,In_992);
or U570 (N_570,In_798,In_818);
xor U571 (N_571,In_558,In_2980);
and U572 (N_572,In_1801,In_1131);
and U573 (N_573,In_595,In_1044);
or U574 (N_574,In_2546,In_1726);
or U575 (N_575,In_2984,In_2188);
and U576 (N_576,In_2779,In_2664);
or U577 (N_577,In_272,In_932);
or U578 (N_578,In_925,In_2874);
or U579 (N_579,In_1823,In_770);
and U580 (N_580,In_2318,In_2186);
or U581 (N_581,In_1767,In_1775);
nand U582 (N_582,In_1697,In_1984);
or U583 (N_583,In_1762,In_1188);
and U584 (N_584,In_946,In_1325);
xor U585 (N_585,In_980,In_543);
nand U586 (N_586,In_1989,In_2389);
nand U587 (N_587,In_1666,In_233);
or U588 (N_588,In_1532,In_1095);
nand U589 (N_589,In_267,In_2993);
xor U590 (N_590,In_2089,In_1023);
nand U591 (N_591,In_1156,In_459);
xor U592 (N_592,In_504,In_2397);
xor U593 (N_593,In_1624,In_1983);
xor U594 (N_594,In_2745,In_1100);
xor U595 (N_595,In_733,In_2652);
nor U596 (N_596,In_2722,In_2476);
or U597 (N_597,In_1190,In_1231);
xor U598 (N_598,In_1006,In_1902);
or U599 (N_599,In_546,In_2521);
xnor U600 (N_600,In_592,In_2701);
xor U601 (N_601,In_1170,In_1161);
and U602 (N_602,In_680,In_87);
nand U603 (N_603,In_1494,In_1720);
or U604 (N_604,In_2351,In_1337);
or U605 (N_605,In_1112,In_58);
or U606 (N_606,In_555,In_1725);
or U607 (N_607,In_679,In_2596);
nor U608 (N_608,In_1073,In_1129);
and U609 (N_609,In_377,In_2646);
nor U610 (N_610,In_2442,In_2541);
xnor U611 (N_611,In_1854,In_768);
and U612 (N_612,In_242,In_2168);
xnor U613 (N_613,In_2266,In_876);
or U614 (N_614,In_359,In_1322);
nor U615 (N_615,In_164,In_406);
nor U616 (N_616,In_2020,In_1357);
nor U617 (N_617,In_261,In_2118);
and U618 (N_618,In_325,In_928);
nand U619 (N_619,In_2444,In_1704);
nand U620 (N_620,In_2240,In_1605);
xor U621 (N_621,In_1661,In_1776);
or U622 (N_622,In_208,In_2872);
and U623 (N_623,In_1372,In_2229);
xor U624 (N_624,In_421,In_1505);
nand U625 (N_625,In_2337,In_2058);
nand U626 (N_626,In_551,In_533);
and U627 (N_627,In_2099,In_929);
nand U628 (N_628,In_2880,In_1348);
and U629 (N_629,In_2015,In_2673);
nand U630 (N_630,In_2688,In_1604);
xnor U631 (N_631,In_2244,In_28);
xor U632 (N_632,In_1703,In_2480);
or U633 (N_633,In_1631,In_307);
xnor U634 (N_634,In_673,In_2426);
nor U635 (N_635,In_1450,In_550);
nand U636 (N_636,In_1334,In_972);
and U637 (N_637,In_494,In_2799);
nand U638 (N_638,In_2612,In_340);
nor U639 (N_639,In_2502,In_2999);
and U640 (N_640,In_2560,In_2302);
or U641 (N_641,In_554,In_1647);
nor U642 (N_642,In_2111,In_2778);
and U643 (N_643,In_75,In_605);
and U644 (N_644,In_2568,In_2795);
and U645 (N_645,In_2311,In_2143);
xnor U646 (N_646,In_2698,In_982);
or U647 (N_647,In_1460,In_1048);
or U648 (N_648,In_278,In_1926);
and U649 (N_649,In_37,In_1256);
and U650 (N_650,In_991,In_2580);
xnor U651 (N_651,In_1428,In_2699);
xor U652 (N_652,In_53,In_674);
xnor U653 (N_653,In_1864,In_2072);
xor U654 (N_654,In_424,In_1475);
nand U655 (N_655,In_542,In_1062);
or U656 (N_656,In_1932,In_522);
nand U657 (N_657,In_1234,In_294);
xnor U658 (N_658,In_2809,In_1371);
and U659 (N_659,In_2789,In_366);
nor U660 (N_660,In_2641,In_1042);
xor U661 (N_661,In_1158,In_1982);
or U662 (N_662,In_1623,In_1359);
or U663 (N_663,In_2227,In_1263);
nor U664 (N_664,In_2985,In_589);
nor U665 (N_665,In_2645,In_1660);
or U666 (N_666,In_2041,In_2021);
nand U667 (N_667,In_2446,In_1087);
nand U668 (N_668,In_2530,In_1219);
nor U669 (N_669,In_528,In_505);
xnor U670 (N_670,In_343,In_809);
and U671 (N_671,In_855,In_2563);
nor U672 (N_672,In_230,In_2602);
and U673 (N_673,In_926,In_681);
nor U674 (N_674,In_1557,In_29);
nor U675 (N_675,In_616,In_428);
or U676 (N_676,In_2083,In_2635);
nand U677 (N_677,In_2550,In_2477);
or U678 (N_678,In_2359,In_1507);
xnor U679 (N_679,In_244,In_418);
nand U680 (N_680,In_2953,In_2929);
and U681 (N_681,In_682,In_2460);
xnor U682 (N_682,In_2304,In_2332);
or U683 (N_683,In_1472,In_2334);
xor U684 (N_684,In_888,In_2421);
nor U685 (N_685,In_2529,In_1691);
nor U686 (N_686,In_178,In_1802);
xnor U687 (N_687,In_985,In_392);
and U688 (N_688,In_2161,In_147);
nor U689 (N_689,In_603,In_866);
nand U690 (N_690,In_954,In_2936);
xor U691 (N_691,In_990,In_1560);
xnor U692 (N_692,In_930,In_1146);
nand U693 (N_693,In_1537,In_1262);
nor U694 (N_694,In_117,In_722);
or U695 (N_695,In_1116,In_1050);
and U696 (N_696,In_1503,In_1722);
xnor U697 (N_697,In_2137,In_109);
or U698 (N_698,In_345,In_5);
or U699 (N_699,In_204,In_2913);
nand U700 (N_700,In_518,In_2840);
or U701 (N_701,In_1523,In_1836);
nand U702 (N_702,In_2540,In_308);
and U703 (N_703,In_2253,In_998);
or U704 (N_704,In_1675,In_1128);
or U705 (N_705,In_115,In_1957);
nor U706 (N_706,In_826,In_1851);
or U707 (N_707,In_2156,In_1458);
and U708 (N_708,In_689,In_1874);
nor U709 (N_709,In_562,In_1739);
and U710 (N_710,In_2079,In_2114);
nor U711 (N_711,In_1867,In_2714);
nand U712 (N_712,In_2094,In_1566);
nor U713 (N_713,In_2060,In_538);
nand U714 (N_714,In_660,In_2112);
nor U715 (N_715,In_2533,In_2264);
or U716 (N_716,In_1406,In_1844);
xor U717 (N_717,In_1657,In_1906);
xor U718 (N_718,In_2684,In_1916);
nand U719 (N_719,In_2973,In_1215);
nor U720 (N_720,In_2629,In_2210);
and U721 (N_721,In_2270,In_902);
nand U722 (N_722,In_1520,In_1580);
or U723 (N_723,In_207,In_785);
and U724 (N_724,In_280,In_1415);
nand U725 (N_725,In_2794,In_1610);
or U726 (N_726,In_1462,In_854);
nor U727 (N_727,In_2780,In_8);
nor U728 (N_728,In_252,In_1561);
and U729 (N_729,In_834,In_739);
xnor U730 (N_730,In_250,In_1368);
or U731 (N_731,In_1221,In_2017);
nor U732 (N_732,In_130,In_69);
nand U733 (N_733,In_2163,In_324);
and U734 (N_734,In_158,In_1734);
and U735 (N_735,In_749,In_1716);
nand U736 (N_736,In_476,In_1629);
or U737 (N_737,In_971,In_397);
nor U738 (N_738,In_2368,In_1991);
xor U739 (N_739,In_911,In_654);
nand U740 (N_740,In_411,In_2954);
nand U741 (N_741,In_906,In_2228);
nand U742 (N_742,In_1518,In_2307);
xnor U743 (N_743,In_1259,In_1919);
nor U744 (N_744,In_2249,In_2601);
and U745 (N_745,In_2090,In_1118);
nor U746 (N_746,In_2997,In_2868);
nand U747 (N_747,In_201,In_2604);
and U748 (N_748,In_1364,In_2516);
xor U749 (N_749,In_2408,In_218);
and U750 (N_750,In_1504,In_1381);
xnor U751 (N_751,In_2828,In_1791);
nand U752 (N_752,In_893,In_153);
nor U753 (N_753,In_2963,In_1644);
nor U754 (N_754,In_2012,In_1961);
nand U755 (N_755,In_652,In_1530);
xnor U756 (N_756,In_650,In_2922);
nand U757 (N_757,In_440,In_126);
nor U758 (N_758,In_1339,In_417);
nand U759 (N_759,In_553,In_2865);
xnor U760 (N_760,In_2567,In_322);
xor U761 (N_761,In_1220,In_2810);
nand U762 (N_762,In_537,In_2198);
xor U763 (N_763,In_483,In_2462);
xor U764 (N_764,In_2147,In_194);
or U765 (N_765,In_2891,In_610);
or U766 (N_766,In_2388,In_2503);
nor U767 (N_767,In_2983,In_790);
nand U768 (N_768,In_1084,In_1565);
nor U769 (N_769,In_2182,In_1103);
nor U770 (N_770,In_2407,In_2758);
xor U771 (N_771,In_2785,In_2995);
xor U772 (N_772,In_129,In_976);
nor U773 (N_773,In_375,In_1920);
or U774 (N_774,In_2727,In_2010);
nand U775 (N_775,In_1081,In_436);
and U776 (N_776,In_2958,In_215);
xor U777 (N_777,In_664,In_299);
xnor U778 (N_778,In_532,In_1283);
and U779 (N_779,In_2102,In_886);
or U780 (N_780,In_2768,In_1319);
xor U781 (N_781,In_1175,In_668);
nor U782 (N_782,In_1491,In_657);
nor U783 (N_783,In_1493,In_2585);
nor U784 (N_784,In_67,In_18);
xnor U785 (N_785,In_85,In_2380);
and U786 (N_786,In_1827,In_984);
nand U787 (N_787,In_2893,In_152);
or U788 (N_788,In_2752,In_1974);
xnor U789 (N_789,In_473,In_2634);
nor U790 (N_790,In_33,In_767);
and U791 (N_791,In_143,In_54);
nor U792 (N_792,In_2258,In_2619);
xor U793 (N_793,In_1020,In_608);
and U794 (N_794,In_1277,In_2232);
nor U795 (N_795,In_139,In_2719);
nor U796 (N_796,In_1453,In_623);
xor U797 (N_797,In_253,In_2151);
xor U798 (N_798,In_786,In_630);
or U799 (N_799,In_128,In_2034);
or U800 (N_800,In_765,In_313);
nor U801 (N_801,In_332,In_1133);
xnor U802 (N_802,In_2029,In_2325);
and U803 (N_803,In_1710,In_62);
and U804 (N_804,In_1872,In_1068);
and U805 (N_805,In_1670,In_2620);
or U806 (N_806,In_1535,In_2683);
and U807 (N_807,In_2537,In_387);
nor U808 (N_808,In_865,In_2499);
xor U809 (N_809,In_961,In_1544);
xnor U810 (N_810,In_515,In_2196);
nor U811 (N_811,In_1597,In_1404);
or U812 (N_812,In_2835,In_1815);
xnor U813 (N_813,In_1673,In_1678);
or U814 (N_814,In_1512,In_2394);
nor U815 (N_815,In_491,In_1211);
and U816 (N_816,In_1132,In_1885);
or U817 (N_817,In_859,In_2545);
xor U818 (N_818,In_1130,In_145);
xor U819 (N_819,In_578,In_442);
or U820 (N_820,In_969,In_2225);
xnor U821 (N_821,In_103,In_169);
and U822 (N_822,In_2435,In_2888);
xnor U823 (N_823,In_747,In_1400);
nand U824 (N_824,In_1613,In_2191);
nand U825 (N_825,In_2459,In_2680);
nor U826 (N_826,In_2565,In_2230);
nor U827 (N_827,In_1832,In_2369);
or U828 (N_828,In_1230,In_631);
xor U829 (N_829,In_606,In_1251);
nor U830 (N_830,In_112,In_2416);
nand U831 (N_831,In_2254,In_2772);
or U832 (N_832,In_2532,In_496);
nor U833 (N_833,In_1781,In_277);
or U834 (N_834,In_113,In_842);
xnor U835 (N_835,In_2221,In_1876);
or U836 (N_836,In_1589,In_703);
nand U837 (N_837,In_1825,In_2991);
or U838 (N_838,In_2290,In_1366);
and U839 (N_839,In_2096,In_2330);
nor U840 (N_840,In_275,In_1835);
xor U841 (N_841,In_2187,In_2605);
xnor U842 (N_842,In_568,In_2295);
nor U843 (N_843,In_2572,In_591);
nand U844 (N_844,In_2925,In_2466);
nand U845 (N_845,In_2338,In_365);
xor U846 (N_846,In_1035,In_894);
xnor U847 (N_847,In_2323,In_2640);
nand U848 (N_848,In_1405,In_297);
or U849 (N_849,In_1852,In_1889);
nor U850 (N_850,In_2193,In_2892);
nand U851 (N_851,In_1935,In_51);
and U852 (N_852,In_694,In_475);
and U853 (N_853,In_1261,In_2988);
nand U854 (N_854,In_880,In_1541);
nand U855 (N_855,In_569,In_1317);
or U856 (N_856,In_618,In_2528);
nand U857 (N_857,In_2552,In_2523);
xor U858 (N_858,In_455,In_1833);
xnor U859 (N_859,In_2405,In_2299);
nor U860 (N_860,In_2934,In_2133);
nor U861 (N_861,In_1267,In_1034);
and U862 (N_862,In_960,In_1309);
xor U863 (N_863,In_1484,In_761);
and U864 (N_864,In_1820,In_2636);
nor U865 (N_865,In_2488,In_2428);
or U866 (N_866,In_168,In_2033);
and U867 (N_867,In_1891,In_1476);
or U868 (N_868,In_760,In_764);
nor U869 (N_869,In_577,In_86);
nor U870 (N_870,In_643,In_852);
xor U871 (N_871,In_2310,In_2841);
or U872 (N_872,In_2879,In_1111);
or U873 (N_873,In_141,In_921);
or U874 (N_874,In_754,In_88);
and U875 (N_875,In_1416,In_2757);
nand U876 (N_876,In_323,In_2536);
and U877 (N_877,In_2989,In_306);
or U878 (N_878,In_2294,In_341);
nand U879 (N_879,In_2940,In_1350);
xor U880 (N_880,In_2340,In_1172);
or U881 (N_881,In_1611,In_1017);
xor U882 (N_882,In_235,In_2091);
nand U883 (N_883,In_116,In_2356);
nand U884 (N_884,In_1214,In_649);
or U885 (N_885,In_2439,In_2003);
nor U886 (N_886,In_628,In_2119);
nor U887 (N_887,In_746,In_2836);
xnor U888 (N_888,In_389,In_187);
or U889 (N_889,In_2650,In_1790);
and U890 (N_890,In_915,In_2961);
and U891 (N_891,In_2767,In_1162);
xnor U892 (N_892,In_1706,In_1690);
xnor U893 (N_893,In_2496,In_2243);
xor U894 (N_894,In_2760,In_2952);
nor U895 (N_895,In_1943,In_367);
nor U896 (N_896,In_2615,In_2205);
nand U897 (N_897,In_1121,In_734);
xnor U898 (N_898,In_2938,In_1411);
or U899 (N_899,In_2926,In_2707);
nand U900 (N_900,In_23,In_748);
nand U901 (N_901,In_388,In_535);
nand U902 (N_902,In_714,In_2517);
or U903 (N_903,In_1303,In_378);
nand U904 (N_904,In_2040,In_1882);
and U905 (N_905,In_445,In_2409);
nand U906 (N_906,In_2103,In_2720);
xnor U907 (N_907,In_1320,In_2741);
or U908 (N_908,In_2948,In_1185);
nor U909 (N_909,In_2526,In_1896);
or U910 (N_910,In_469,In_2190);
and U911 (N_911,In_1061,In_531);
nand U912 (N_912,In_1571,In_1482);
xnor U913 (N_913,In_2053,In_614);
and U914 (N_914,In_1032,In_2207);
nor U915 (N_915,In_1232,In_2561);
or U916 (N_916,In_2697,In_1962);
and U917 (N_917,In_196,In_1842);
nor U918 (N_918,In_851,In_2429);
or U919 (N_919,In_2866,In_2215);
xnor U920 (N_920,In_1816,In_2539);
nor U921 (N_921,In_1681,In_2061);
nor U922 (N_922,In_1031,In_2125);
nor U923 (N_923,In_943,In_2321);
and U924 (N_924,In_1074,In_2917);
nor U925 (N_925,In_1884,In_927);
and U926 (N_926,In_391,In_2986);
or U927 (N_927,In_2365,In_15);
or U928 (N_928,In_1618,In_2626);
and U929 (N_929,In_1409,In_2609);
nand U930 (N_930,In_127,In_2844);
xor U931 (N_931,In_314,In_2592);
nand U932 (N_932,In_964,In_2128);
or U933 (N_933,In_1810,In_864);
nor U934 (N_934,In_1608,In_2180);
nand U935 (N_935,In_769,In_1239);
xnor U936 (N_936,In_384,In_2075);
nor U937 (N_937,In_107,In_539);
xnor U938 (N_938,In_2878,In_1517);
nand U939 (N_939,In_97,In_2277);
and U940 (N_940,In_1355,In_2363);
xnor U941 (N_941,In_920,In_1972);
and U942 (N_942,In_27,In_1449);
nand U943 (N_943,In_2218,In_2686);
or U944 (N_944,In_2392,In_1326);
and U945 (N_945,In_2263,In_1787);
nand U946 (N_946,In_728,In_2728);
nor U947 (N_947,In_1612,In_1648);
xor U948 (N_948,In_1633,In_291);
xor U949 (N_949,In_1445,In_1354);
nor U950 (N_950,In_1649,In_637);
or U951 (N_951,In_2815,In_2886);
or U952 (N_952,In_1514,In_1437);
or U953 (N_953,In_1761,In_2461);
or U954 (N_954,In_1293,In_229);
or U955 (N_955,In_1866,In_651);
or U956 (N_956,In_1080,In_1037);
nand U957 (N_957,In_336,In_1489);
or U958 (N_958,In_1595,In_1386);
nand U959 (N_959,In_2875,In_2786);
xor U960 (N_960,In_2478,In_974);
and U961 (N_961,In_240,In_195);
or U962 (N_962,In_841,In_2632);
and U963 (N_963,In_2179,In_869);
and U964 (N_964,In_1194,In_2274);
or U965 (N_965,In_63,In_1575);
xor U966 (N_966,In_2569,In_2554);
and U967 (N_967,In_1850,In_1847);
xnor U968 (N_968,In_2834,In_1091);
nor U969 (N_969,In_951,In_262);
or U970 (N_970,In_1269,In_2725);
nor U971 (N_971,In_1402,In_1124);
nor U972 (N_972,In_1637,In_2373);
and U973 (N_973,In_903,In_821);
nand U974 (N_974,In_719,In_567);
nor U975 (N_975,In_2564,In_2370);
xor U976 (N_976,In_2527,In_2649);
nand U977 (N_977,In_2181,In_114);
and U978 (N_978,In_897,In_1601);
xor U979 (N_979,In_2023,In_99);
nand U980 (N_980,In_2557,In_2357);
xor U981 (N_981,In_1559,In_2945);
or U982 (N_982,In_502,In_2275);
or U983 (N_983,In_811,In_2663);
and U984 (N_984,In_2671,In_1772);
and U985 (N_985,In_1642,In_1358);
nand U986 (N_986,In_331,In_653);
nor U987 (N_987,In_198,In_683);
and U988 (N_988,In_42,In_2847);
xor U989 (N_989,In_641,In_579);
nor U990 (N_990,In_111,In_2666);
xor U991 (N_991,In_1988,In_379);
nor U992 (N_992,In_1279,In_1004);
nand U993 (N_993,In_829,In_957);
nand U994 (N_994,In_1301,In_968);
nor U995 (N_995,In_2214,In_839);
nor U996 (N_996,In_1969,In_1582);
nor U997 (N_997,In_1964,In_1148);
and U998 (N_998,In_1483,In_430);
and U999 (N_999,In_2715,In_2566);
or U1000 (N_1000,In_580,In_752);
or U1001 (N_1001,In_2293,In_2848);
xor U1002 (N_1002,In_65,In_574);
or U1003 (N_1003,In_1094,In_1636);
or U1004 (N_1004,In_509,In_2587);
nor U1005 (N_1005,In_303,In_2811);
or U1006 (N_1006,In_223,In_1295);
and U1007 (N_1007,In_1127,In_501);
and U1008 (N_1008,In_586,In_2004);
xor U1009 (N_1009,In_467,In_385);
nand U1010 (N_1010,In_493,In_1976);
nand U1011 (N_1011,In_1058,In_1996);
or U1012 (N_1012,In_2849,In_950);
and U1013 (N_1013,In_1918,In_222);
nor U1014 (N_1014,In_1195,In_220);
and U1015 (N_1015,In_2504,In_1045);
nand U1016 (N_1016,In_416,In_2842);
xnor U1017 (N_1017,In_2920,In_2080);
xnor U1018 (N_1018,In_2044,In_1076);
and U1019 (N_1019,In_1164,In_2410);
xor U1020 (N_1020,In_395,In_1459);
or U1021 (N_1021,In_2297,In_2471);
or U1022 (N_1022,In_120,In_1105);
and U1023 (N_1023,In_762,In_1333);
xor U1024 (N_1024,In_210,In_2141);
xnor U1025 (N_1025,In_2884,In_1527);
xnor U1026 (N_1026,In_1390,In_536);
and U1027 (N_1027,In_2624,In_500);
xnor U1028 (N_1028,In_2716,In_881);
or U1029 (N_1029,In_1914,In_1998);
nand U1030 (N_1030,In_2738,In_895);
and U1031 (N_1031,In_1199,In_2386);
and U1032 (N_1032,In_1299,In_2054);
and U1033 (N_1033,In_2013,In_1003);
nand U1034 (N_1034,In_0,In_1021);
xnor U1035 (N_1035,In_1958,In_2919);
nand U1036 (N_1036,In_1135,In_1743);
or U1037 (N_1037,In_2036,In_2367);
nor U1038 (N_1038,In_1024,In_919);
and U1039 (N_1039,In_1447,In_2932);
or U1040 (N_1040,In_2267,In_2749);
xor U1041 (N_1041,In_487,In_564);
nand U1042 (N_1042,In_1576,In_2562);
nand U1043 (N_1043,In_1593,In_2030);
xnor U1044 (N_1044,In_1030,In_1446);
and U1045 (N_1045,In_2001,In_1344);
nand U1046 (N_1046,In_1915,In_1711);
nand U1047 (N_1047,In_1027,In_793);
and U1048 (N_1048,In_1714,In_1538);
and U1049 (N_1049,In_288,In_938);
xnor U1050 (N_1050,In_2067,In_159);
xor U1051 (N_1051,In_260,In_1289);
nor U1052 (N_1052,In_1683,In_1857);
and U1053 (N_1053,In_495,In_1900);
xnor U1054 (N_1054,In_1570,In_1010);
nor U1055 (N_1055,In_1181,In_1979);
or U1056 (N_1056,In_1488,In_833);
nor U1057 (N_1057,In_2009,In_2726);
and U1058 (N_1058,In_1577,In_1638);
or U1059 (N_1059,In_2007,In_2706);
xor U1060 (N_1060,In_348,In_2750);
or U1061 (N_1061,In_530,In_2105);
nor U1062 (N_1062,In_1868,In_1937);
nor U1063 (N_1063,In_2482,In_356);
nor U1064 (N_1064,In_2443,In_526);
and U1065 (N_1065,In_908,In_905);
nand U1066 (N_1066,In_1698,In_2943);
nand U1067 (N_1067,In_2059,In_2272);
and U1068 (N_1068,In_2861,In_123);
or U1069 (N_1069,In_2345,In_2827);
or U1070 (N_1070,In_684,In_1981);
or U1071 (N_1071,In_461,In_2463);
xor U1072 (N_1072,In_941,In_2905);
and U1073 (N_1073,In_1853,In_2076);
and U1074 (N_1074,In_1424,In_2217);
nor U1075 (N_1075,In_1163,In_2992);
nor U1076 (N_1076,In_878,In_698);
xor U1077 (N_1077,In_1963,In_352);
and U1078 (N_1078,In_1323,In_1563);
and U1079 (N_1079,In_2712,In_1176);
xnor U1080 (N_1080,In_70,In_1890);
and U1081 (N_1081,In_559,In_2457);
or U1082 (N_1082,In_1443,In_713);
and U1083 (N_1083,In_1384,In_2379);
or U1084 (N_1084,In_2911,In_2807);
or U1085 (N_1085,In_2655,In_446);
nor U1086 (N_1086,In_1928,In_2723);
and U1087 (N_1087,In_134,In_2183);
or U1088 (N_1088,In_1993,In_438);
and U1089 (N_1089,In_259,In_1938);
and U1090 (N_1090,In_1029,In_2495);
nand U1091 (N_1091,In_2730,In_2647);
nor U1092 (N_1092,In_1187,In_225);
or U1093 (N_1093,In_106,In_154);
and U1094 (N_1094,In_1546,In_1778);
nor U1095 (N_1095,In_1662,In_1526);
nand U1096 (N_1096,In_1486,In_557);
or U1097 (N_1097,In_2281,In_2241);
nand U1098 (N_1098,In_1286,In_1113);
or U1099 (N_1099,In_899,In_2656);
nand U1100 (N_1100,In_444,In_1812);
xnor U1101 (N_1101,In_2648,In_2399);
xor U1102 (N_1102,In_144,In_2385);
xor U1103 (N_1103,In_1875,In_1551);
nor U1104 (N_1104,In_1432,In_1764);
xor U1105 (N_1105,In_2178,In_1700);
xor U1106 (N_1106,In_77,In_160);
or U1107 (N_1107,In_672,In_2851);
and U1108 (N_1108,In_2637,In_1473);
xnor U1109 (N_1109,In_1924,In_2333);
or U1110 (N_1110,In_1360,In_1466);
or U1111 (N_1111,In_2897,In_916);
and U1112 (N_1112,In_1412,In_952);
xor U1113 (N_1113,In_791,In_2581);
and U1114 (N_1114,In_669,In_732);
and U1115 (N_1115,In_2855,In_213);
xnor U1116 (N_1116,In_1154,In_2485);
xor U1117 (N_1117,In_2481,In_81);
nand U1118 (N_1118,In_945,In_105);
xnor U1119 (N_1119,In_1939,In_1308);
or U1120 (N_1120,In_2603,In_1237);
xor U1121 (N_1121,In_2623,In_1186);
nand U1122 (N_1122,In_2391,In_1583);
nor U1123 (N_1123,In_1646,In_2812);
nor U1124 (N_1124,In_1481,In_237);
nor U1125 (N_1125,In_1861,In_2039);
nor U1126 (N_1126,In_1236,In_1547);
xnor U1127 (N_1127,In_337,In_465);
nand U1128 (N_1128,In_1863,In_521);
nor U1129 (N_1129,In_2005,In_756);
or U1130 (N_1130,In_1419,In_1014);
nor U1131 (N_1131,In_782,In_2018);
nor U1132 (N_1132,In_2026,In_2115);
and U1133 (N_1133,In_450,In_1542);
xnor U1134 (N_1134,In_61,In_2754);
nor U1135 (N_1135,In_979,In_407);
nor U1136 (N_1136,In_2951,In_836);
nand U1137 (N_1137,In_1356,In_1268);
xnor U1138 (N_1138,In_1165,In_1724);
nand U1139 (N_1139,In_1079,In_896);
nand U1140 (N_1140,In_1806,In_2691);
nand U1141 (N_1141,In_236,In_599);
nand U1142 (N_1142,In_1137,In_840);
xor U1143 (N_1143,In_2885,In_2696);
and U1144 (N_1144,In_499,In_665);
xnor U1145 (N_1145,In_2520,In_2038);
nor U1146 (N_1146,In_576,In_2627);
and U1147 (N_1147,In_2127,In_101);
nor U1148 (N_1148,In_1929,In_784);
nor U1149 (N_1149,In_2200,In_1260);
and U1150 (N_1150,In_2047,In_2092);
and U1151 (N_1151,In_410,In_815);
xnor U1152 (N_1152,In_2559,In_634);
nand U1153 (N_1153,In_2077,In_479);
and U1154 (N_1154,In_823,In_2658);
nand U1155 (N_1155,In_1285,In_2908);
xnor U1156 (N_1156,In_2965,In_1849);
nand U1157 (N_1157,In_1632,In_1063);
nor U1158 (N_1158,In_2043,In_949);
nor U1159 (N_1159,In_2614,In_1169);
nand U1160 (N_1160,In_279,In_1427);
nand U1161 (N_1161,In_2735,In_741);
nor U1162 (N_1162,In_2690,In_1414);
or U1163 (N_1163,In_1470,In_1730);
nand U1164 (N_1164,In_21,In_2195);
nor U1165 (N_1165,In_1370,In_95);
nand U1166 (N_1166,In_2285,In_1069);
nand U1167 (N_1167,In_363,In_2284);
and U1168 (N_1168,In_2918,In_1584);
nor U1169 (N_1169,In_570,In_1420);
or U1170 (N_1170,In_2704,In_2713);
and U1171 (N_1171,In_2238,In_629);
xnor U1172 (N_1172,In_1057,In_2068);
nor U1173 (N_1173,In_2662,In_56);
and U1174 (N_1174,In_612,In_464);
nand U1175 (N_1175,In_2441,In_165);
and U1176 (N_1176,In_310,In_2219);
and U1177 (N_1177,In_89,In_1792);
nand U1178 (N_1178,In_1519,In_885);
xnor U1179 (N_1179,In_1182,In_47);
or U1180 (N_1180,In_581,In_132);
xor U1181 (N_1181,In_2245,In_1075);
xnor U1182 (N_1182,In_2708,In_1153);
or U1183 (N_1183,In_2678,In_2322);
or U1184 (N_1184,In_2787,In_226);
or U1185 (N_1185,In_2979,In_2171);
nand U1186 (N_1186,In_1879,In_2711);
and U1187 (N_1187,In_174,In_989);
xnor U1188 (N_1188,In_1978,In_600);
xnor U1189 (N_1189,In_588,In_1329);
nor U1190 (N_1190,In_822,In_711);
xor U1191 (N_1191,In_1352,In_1750);
nor U1192 (N_1192,In_1522,In_801);
xnor U1193 (N_1193,In_2542,In_1316);
nor U1194 (N_1194,In_2769,In_2148);
and U1195 (N_1195,In_2764,In_2008);
or U1196 (N_1196,In_73,In_477);
and U1197 (N_1197,In_1318,In_2303);
xor U1198 (N_1198,In_191,In_1173);
xor U1199 (N_1199,In_2074,In_2413);
and U1200 (N_1200,In_1682,In_1392);
and U1201 (N_1201,In_942,In_2211);
nand U1202 (N_1202,In_328,In_1839);
and U1203 (N_1203,In_693,In_1353);
or U1204 (N_1204,In_1696,In_2548);
nor U1205 (N_1205,In_172,In_716);
xnor U1206 (N_1206,In_1036,In_399);
and U1207 (N_1207,In_420,In_1418);
xnor U1208 (N_1208,In_137,In_205);
nor U1209 (N_1209,In_2101,In_2896);
xor U1210 (N_1210,In_1873,In_2417);
or U1211 (N_1211,In_1688,In_232);
xnor U1212 (N_1212,In_40,In_34);
nand U1213 (N_1213,In_1596,In_860);
nand U1214 (N_1214,In_2633,In_867);
and U1215 (N_1215,In_1477,In_593);
and U1216 (N_1216,In_2450,In_1383);
nor U1217 (N_1217,In_2509,In_12);
and U1218 (N_1218,In_2145,In_870);
nor U1219 (N_1219,In_427,In_2456);
and U1220 (N_1220,In_422,In_738);
nand U1221 (N_1221,In_1054,In_2420);
and U1222 (N_1222,In_2525,In_983);
or U1223 (N_1223,In_1797,In_319);
and U1224 (N_1224,In_2668,In_2733);
nand U1225 (N_1225,In_2558,In_1752);
nand U1226 (N_1226,In_1040,In_1917);
or U1227 (N_1227,In_661,In_2085);
or U1228 (N_1228,In_2153,In_2129);
xor U1229 (N_1229,In_1878,In_90);
and U1230 (N_1230,In_2870,In_2969);
or U1231 (N_1231,In_2621,In_404);
and U1232 (N_1232,In_2981,In_2022);
nor U1233 (N_1233,In_910,In_648);
or U1234 (N_1234,In_736,In_394);
nand U1235 (N_1235,In_2755,In_2204);
or U1236 (N_1236,In_794,In_590);
xnor U1237 (N_1237,In_1771,In_2434);
nor U1238 (N_1238,In_1705,In_11);
xor U1239 (N_1239,In_1908,In_2818);
nor U1240 (N_1240,In_640,In_1005);
nand U1241 (N_1241,In_2256,In_1469);
xnor U1242 (N_1242,In_2514,In_2702);
xor U1243 (N_1243,In_423,In_2717);
xnor U1244 (N_1244,In_2687,In_1143);
and U1245 (N_1245,In_189,In_182);
xnor U1246 (N_1246,In_2850,In_2237);
nand U1247 (N_1247,In_2618,In_2957);
nor U1248 (N_1248,In_2269,In_1208);
and U1249 (N_1249,In_1600,In_2804);
or U1250 (N_1250,In_83,In_808);
and U1251 (N_1251,In_1312,In_338);
xor U1252 (N_1252,In_1255,In_1313);
and U1253 (N_1253,In_918,In_1769);
nor U1254 (N_1254,In_1055,In_157);
nor U1255 (N_1255,In_582,In_763);
or U1256 (N_1256,In_638,In_2037);
and U1257 (N_1257,In_758,In_718);
nor U1258 (N_1258,In_100,In_1248);
or U1259 (N_1259,In_2937,In_2213);
or U1260 (N_1260,In_2223,In_2142);
nor U1261 (N_1261,In_1773,In_620);
and U1262 (N_1262,In_596,In_2508);
or U1263 (N_1263,In_2436,In_212);
xor U1264 (N_1264,In_257,In_635);
and U1265 (N_1265,In_1784,In_861);
xor U1266 (N_1266,In_1056,In_1119);
xnor U1267 (N_1267,In_1101,In_2535);
nor U1268 (N_1268,In_935,In_2268);
xor U1269 (N_1269,In_1053,In_691);
and U1270 (N_1270,In_1280,In_488);
nor U1271 (N_1271,In_745,In_2538);
and U1272 (N_1272,In_759,In_1960);
nor U1273 (N_1273,In_585,In_2591);
xor U1274 (N_1274,In_1431,In_2946);
nand U1275 (N_1275,In_2689,In_1229);
xnor U1276 (N_1276,In_2472,In_2470);
nor U1277 (N_1277,In_2025,In_2676);
or U1278 (N_1278,In_2823,In_2088);
or U1279 (N_1279,In_2465,In_2406);
nor U1280 (N_1280,In_704,In_2748);
nor U1281 (N_1281,In_2821,In_800);
nand U1282 (N_1282,In_1659,In_2063);
and U1283 (N_1283,In_2189,In_2607);
or U1284 (N_1284,In_2724,In_602);
xor U1285 (N_1285,In_177,In_1374);
or U1286 (N_1286,In_686,In_2384);
and U1287 (N_1287,In_1959,In_2867);
or U1288 (N_1288,In_2966,In_2317);
xnor U1289 (N_1289,In_298,In_2597);
nand U1290 (N_1290,In_545,In_566);
xor U1291 (N_1291,In_2140,In_1686);
nand U1292 (N_1292,In_1015,In_2901);
nand U1293 (N_1293,In_2916,In_1209);
nand U1294 (N_1294,In_334,In_1898);
or U1295 (N_1295,In_330,In_2051);
or U1296 (N_1296,In_1007,In_2862);
nor U1297 (N_1297,In_361,In_1072);
and U1298 (N_1298,In_1650,In_2433);
nand U1299 (N_1299,In_1410,In_2910);
or U1300 (N_1300,In_354,In_1843);
or U1301 (N_1301,In_270,In_970);
and U1302 (N_1302,In_9,In_458);
nand U1303 (N_1303,In_2575,In_771);
xor U1304 (N_1304,In_1925,In_1340);
and U1305 (N_1305,In_510,In_529);
nand U1306 (N_1306,In_1448,In_2346);
or U1307 (N_1307,In_6,In_2226);
nand U1308 (N_1308,In_2797,In_2292);
and U1309 (N_1309,In_1346,In_1645);
and U1310 (N_1310,In_663,In_626);
and U1311 (N_1311,In_1387,In_1361);
nand U1312 (N_1312,In_1160,In_1284);
or U1313 (N_1313,In_2396,In_1758);
nor U1314 (N_1314,In_326,In_2589);
or U1315 (N_1315,In_1451,In_1746);
nor U1316 (N_1316,In_2278,In_1385);
and U1317 (N_1317,In_1171,In_2927);
or U1318 (N_1318,In_2829,In_2144);
and U1319 (N_1319,In_2184,In_329);
nor U1320 (N_1320,In_2576,In_449);
nor U1321 (N_1321,In_36,In_206);
nand U1322 (N_1322,In_1945,In_1707);
and U1323 (N_1323,In_1599,In_1855);
nand U1324 (N_1324,In_695,In_2107);
or U1325 (N_1325,In_1439,In_2352);
or U1326 (N_1326,In_847,In_414);
nand U1327 (N_1327,In_333,In_2746);
or U1328 (N_1328,In_2073,In_480);
or U1329 (N_1329,In_783,In_2296);
and U1330 (N_1330,In_1550,In_812);
nand U1331 (N_1331,In_2763,In_2837);
xor U1332 (N_1332,In_1780,In_742);
or U1333 (N_1333,In_1911,In_2265);
xnor U1334 (N_1334,In_2122,In_1627);
or U1335 (N_1335,In_2192,In_1971);
and U1336 (N_1336,In_231,In_2185);
nor U1337 (N_1337,In_26,In_1305);
nor U1338 (N_1338,In_2224,In_1434);
nor U1339 (N_1339,In_1282,In_1748);
nor U1340 (N_1340,In_497,In_1674);
or U1341 (N_1341,In_2579,In_1506);
xnor U1342 (N_1342,In_647,In_549);
nand U1343 (N_1343,In_788,In_863);
nor U1344 (N_1344,In_2651,In_1287);
nor U1345 (N_1345,In_1281,In_967);
or U1346 (N_1346,In_211,In_2326);
and U1347 (N_1347,In_1496,In_1198);
nand U1348 (N_1348,In_266,In_462);
or U1349 (N_1349,In_295,In_1892);
nand U1350 (N_1350,In_1927,In_1826);
nand U1351 (N_1351,In_1492,In_2050);
or U1352 (N_1352,In_2313,In_780);
and U1353 (N_1353,In_2975,In_2120);
or U1354 (N_1354,In_1365,In_2625);
nor U1355 (N_1355,In_1887,In_560);
xor U1356 (N_1356,In_1191,In_1619);
xnor U1357 (N_1357,In_1421,In_269);
nor U1358 (N_1358,In_2793,In_1274);
or U1359 (N_1359,In_2599,In_2149);
nor U1360 (N_1360,In_2093,In_2906);
nor U1361 (N_1361,In_1653,In_1167);
or U1362 (N_1362,In_2555,In_2283);
or U1363 (N_1363,In_283,In_2761);
xor U1364 (N_1364,In_1744,In_2197);
nand U1365 (N_1365,In_2000,In_1120);
and U1366 (N_1366,In_1719,In_1417);
or U1367 (N_1367,In_2998,In_685);
xor U1368 (N_1368,In_1013,In_22);
and U1369 (N_1369,In_2792,In_2974);
nor U1370 (N_1370,In_2826,In_234);
nor U1371 (N_1371,In_2976,In_2675);
or U1372 (N_1372,In_2498,In_251);
nor U1373 (N_1373,In_645,In_2639);
or U1374 (N_1374,In_1338,In_1944);
nor U1375 (N_1375,In_1077,In_2035);
nor U1376 (N_1376,In_2736,In_1513);
and U1377 (N_1377,In_1663,In_1243);
and U1378 (N_1378,In_245,In_511);
and U1379 (N_1379,In_104,In_2831);
nand U1380 (N_1380,In_1180,In_2947);
or U1381 (N_1381,In_317,In_1794);
nor U1382 (N_1382,In_2494,In_302);
or U1383 (N_1383,In_2742,In_2427);
nor U1384 (N_1384,In_1831,In_1038);
and U1385 (N_1385,In_1965,In_1590);
nand U1386 (N_1386,In_1265,In_874);
xor U1387 (N_1387,In_94,In_1422);
nand U1388 (N_1388,In_832,In_2469);
nor U1389 (N_1389,In_2522,In_850);
xnor U1390 (N_1390,In_513,In_1066);
nor U1391 (N_1391,In_1145,In_1973);
xnor U1392 (N_1392,In_1206,In_1258);
nor U1393 (N_1393,In_1442,In_1092);
and U1394 (N_1394,In_1985,In_2928);
xor U1395 (N_1395,In_753,In_887);
xnor U1396 (N_1396,In_904,In_2531);
and U1397 (N_1397,In_1090,In_2011);
and U1398 (N_1398,In_1246,In_1671);
nor U1399 (N_1399,In_1564,In_1568);
nand U1400 (N_1400,In_525,In_2956);
nand U1401 (N_1401,In_2314,In_358);
and U1402 (N_1402,In_2941,In_2378);
and U1403 (N_1403,In_1241,In_1335);
nand U1404 (N_1404,In_2231,In_548);
nor U1405 (N_1405,In_369,In_1216);
and U1406 (N_1406,In_2049,In_2914);
and U1407 (N_1407,In_2341,In_937);
xor U1408 (N_1408,In_1288,In_1097);
or U1409 (N_1409,In_597,In_2166);
or U1410 (N_1410,In_1106,In_2971);
and U1411 (N_1411,In_1093,In_2447);
and U1412 (N_1412,In_587,In_258);
nand U1413 (N_1413,In_2418,In_119);
nand U1414 (N_1414,In_1049,In_180);
and U1415 (N_1415,In_2393,In_2871);
nor U1416 (N_1416,In_2130,In_517);
or U1417 (N_1417,In_2873,In_2653);
and U1418 (N_1418,In_76,In_335);
nand U1419 (N_1419,In_2233,In_2006);
nand U1420 (N_1420,In_1011,In_1292);
xnor U1421 (N_1421,In_776,In_439);
or U1422 (N_1422,In_1399,In_2423);
xnor U1423 (N_1423,In_792,In_2900);
or U1424 (N_1424,In_161,In_163);
and U1425 (N_1425,In_2820,In_819);
or U1426 (N_1426,In_52,In_1603);
or U1427 (N_1427,In_1302,In_2132);
nor U1428 (N_1428,In_327,In_2110);
and U1429 (N_1429,In_779,In_84);
nor U1430 (N_1430,In_408,In_1870);
nand U1431 (N_1431,In_17,In_1272);
nor U1432 (N_1432,In_2731,In_2935);
xor U1433 (N_1433,In_1184,In_1869);
nand U1434 (N_1434,In_2790,In_868);
and U1435 (N_1435,In_1332,In_699);
nand U1436 (N_1436,In_2895,In_2994);
nand U1437 (N_1437,In_687,In_2286);
and U1438 (N_1438,In_1149,In_1088);
nand U1439 (N_1439,In_248,In_2774);
nand U1440 (N_1440,In_1264,In_2095);
and U1441 (N_1441,In_2194,In_2064);
xor U1442 (N_1442,In_1656,In_149);
nor U1443 (N_1443,In_1733,In_1692);
or U1444 (N_1444,In_1616,In_133);
and U1445 (N_1445,In_2933,In_948);
nor U1446 (N_1446,In_514,In_1183);
xnor U1447 (N_1447,In_1987,In_1060);
and U1448 (N_1448,In_2501,In_239);
nand U1449 (N_1449,In_2921,In_353);
nor U1450 (N_1450,In_2320,In_1956);
or U1451 (N_1451,In_2487,In_2349);
xnor U1452 (N_1452,In_737,In_1856);
xor U1453 (N_1453,In_2425,In_884);
nand U1454 (N_1454,In_1860,In_49);
and U1455 (N_1455,In_2949,In_2654);
xnor U1456 (N_1456,In_1468,In_1569);
nor U1457 (N_1457,In_1813,In_2361);
and U1458 (N_1458,In_1117,In_2169);
nand U1459 (N_1459,In_2669,In_2387);
nor U1460 (N_1460,In_43,In_482);
and U1461 (N_1461,In_2424,In_2617);
or U1462 (N_1462,In_1114,In_2721);
nor U1463 (N_1463,In_1795,In_2547);
and U1464 (N_1464,In_1321,In_1718);
xnor U1465 (N_1465,In_2066,In_2681);
and U1466 (N_1466,In_1296,In_2611);
or U1467 (N_1467,In_431,In_2806);
or U1468 (N_1468,In_1930,In_622);
or U1469 (N_1469,In_2505,In_1732);
nand U1470 (N_1470,In_838,In_19);
nor U1471 (N_1471,In_2355,In_1444);
nand U1472 (N_1472,In_627,In_1002);
xnor U1473 (N_1473,In_91,In_415);
xor U1474 (N_1474,In_1555,In_1495);
and U1475 (N_1475,In_639,In_2167);
nor U1476 (N_1476,In_2262,In_2100);
nor U1477 (N_1477,In_2594,In_1966);
nor U1478 (N_1478,In_484,In_271);
nor U1479 (N_1479,In_1765,In_1742);
and U1480 (N_1480,In_1805,In_2486);
nor U1481 (N_1481,In_2121,In_917);
and U1482 (N_1482,In_1516,In_2869);
or U1483 (N_1483,In_2055,In_1115);
and U1484 (N_1484,In_409,In_2833);
xnor U1485 (N_1485,In_2328,In_1665);
nand U1486 (N_1486,In_1331,In_1783);
or U1487 (N_1487,In_1689,In_268);
xnor U1488 (N_1488,In_692,In_1740);
and U1489 (N_1489,In_2452,In_2729);
nand U1490 (N_1490,In_2398,In_1012);
nand U1491 (N_1491,In_2123,In_2108);
or U1492 (N_1492,In_2032,In_1904);
xor U1493 (N_1493,In_2816,In_1997);
xor U1494 (N_1494,In_901,In_2305);
xor U1495 (N_1495,In_1278,In_2751);
nor U1496 (N_1496,In_2106,In_1975);
nor U1497 (N_1497,In_2638,In_2577);
xor U1498 (N_1498,In_2996,In_1071);
or U1499 (N_1499,In_2784,In_1202);
nor U1500 (N_1500,In_785,In_2433);
nand U1501 (N_1501,In_2149,In_385);
nand U1502 (N_1502,In_413,In_1195);
and U1503 (N_1503,In_2223,In_423);
nand U1504 (N_1504,In_2510,In_2280);
nand U1505 (N_1505,In_1102,In_2423);
and U1506 (N_1506,In_2442,In_2990);
and U1507 (N_1507,In_2529,In_363);
xnor U1508 (N_1508,In_497,In_1855);
nand U1509 (N_1509,In_160,In_1866);
and U1510 (N_1510,In_648,In_1271);
and U1511 (N_1511,In_853,In_1958);
nand U1512 (N_1512,In_2717,In_2957);
and U1513 (N_1513,In_198,In_579);
xor U1514 (N_1514,In_1826,In_1618);
or U1515 (N_1515,In_838,In_112);
and U1516 (N_1516,In_886,In_1489);
nor U1517 (N_1517,In_602,In_2685);
or U1518 (N_1518,In_2343,In_324);
nor U1519 (N_1519,In_1590,In_1080);
and U1520 (N_1520,In_1327,In_2663);
xor U1521 (N_1521,In_1039,In_1742);
xor U1522 (N_1522,In_584,In_2165);
and U1523 (N_1523,In_2702,In_708);
xnor U1524 (N_1524,In_2669,In_1440);
xor U1525 (N_1525,In_2907,In_578);
or U1526 (N_1526,In_2933,In_16);
and U1527 (N_1527,In_2986,In_2475);
xnor U1528 (N_1528,In_1778,In_1501);
nor U1529 (N_1529,In_1559,In_225);
nand U1530 (N_1530,In_2095,In_701);
xor U1531 (N_1531,In_2314,In_1368);
xnor U1532 (N_1532,In_1677,In_1004);
nand U1533 (N_1533,In_2477,In_1068);
xor U1534 (N_1534,In_183,In_840);
or U1535 (N_1535,In_2855,In_2292);
nor U1536 (N_1536,In_326,In_1893);
nand U1537 (N_1537,In_2089,In_516);
xnor U1538 (N_1538,In_1,In_1001);
xnor U1539 (N_1539,In_1668,In_222);
xnor U1540 (N_1540,In_319,In_1838);
xor U1541 (N_1541,In_1704,In_925);
nor U1542 (N_1542,In_917,In_1987);
and U1543 (N_1543,In_436,In_2475);
nand U1544 (N_1544,In_1013,In_2544);
or U1545 (N_1545,In_627,In_1261);
or U1546 (N_1546,In_2187,In_59);
nand U1547 (N_1547,In_1371,In_2102);
nor U1548 (N_1548,In_2911,In_1311);
xnor U1549 (N_1549,In_2840,In_2966);
nor U1550 (N_1550,In_893,In_968);
or U1551 (N_1551,In_707,In_1461);
nor U1552 (N_1552,In_2592,In_916);
nor U1553 (N_1553,In_2019,In_2994);
xnor U1554 (N_1554,In_240,In_2078);
xnor U1555 (N_1555,In_353,In_2568);
or U1556 (N_1556,In_473,In_750);
and U1557 (N_1557,In_833,In_324);
or U1558 (N_1558,In_1955,In_1209);
or U1559 (N_1559,In_170,In_2717);
xnor U1560 (N_1560,In_748,In_200);
or U1561 (N_1561,In_2524,In_31);
nor U1562 (N_1562,In_805,In_1006);
and U1563 (N_1563,In_711,In_308);
or U1564 (N_1564,In_2867,In_1886);
xnor U1565 (N_1565,In_2519,In_2908);
and U1566 (N_1566,In_327,In_1749);
xnor U1567 (N_1567,In_500,In_2886);
or U1568 (N_1568,In_1779,In_2459);
and U1569 (N_1569,In_1462,In_185);
or U1570 (N_1570,In_0,In_261);
nor U1571 (N_1571,In_2920,In_2064);
nand U1572 (N_1572,In_2595,In_2262);
or U1573 (N_1573,In_2882,In_2134);
nor U1574 (N_1574,In_998,In_822);
and U1575 (N_1575,In_517,In_1861);
and U1576 (N_1576,In_461,In_1532);
and U1577 (N_1577,In_2956,In_1651);
xor U1578 (N_1578,In_2322,In_1354);
xor U1579 (N_1579,In_1116,In_1879);
nor U1580 (N_1580,In_928,In_2424);
nand U1581 (N_1581,In_1957,In_1286);
and U1582 (N_1582,In_2094,In_591);
or U1583 (N_1583,In_784,In_2717);
or U1584 (N_1584,In_2833,In_1974);
and U1585 (N_1585,In_913,In_1286);
and U1586 (N_1586,In_1497,In_1229);
xnor U1587 (N_1587,In_1413,In_392);
nand U1588 (N_1588,In_2332,In_1686);
xor U1589 (N_1589,In_2665,In_2821);
xnor U1590 (N_1590,In_2199,In_2890);
and U1591 (N_1591,In_2368,In_2460);
nor U1592 (N_1592,In_217,In_2473);
nand U1593 (N_1593,In_1587,In_651);
or U1594 (N_1594,In_955,In_1055);
and U1595 (N_1595,In_966,In_1360);
nand U1596 (N_1596,In_10,In_1043);
xnor U1597 (N_1597,In_1627,In_2838);
nand U1598 (N_1598,In_2947,In_1903);
nand U1599 (N_1599,In_2350,In_1808);
xnor U1600 (N_1600,In_1729,In_1191);
xnor U1601 (N_1601,In_279,In_328);
or U1602 (N_1602,In_2728,In_1058);
and U1603 (N_1603,In_258,In_1337);
nand U1604 (N_1604,In_461,In_878);
or U1605 (N_1605,In_609,In_113);
or U1606 (N_1606,In_2229,In_692);
or U1607 (N_1607,In_2872,In_1657);
nand U1608 (N_1608,In_2043,In_2277);
or U1609 (N_1609,In_824,In_2069);
nand U1610 (N_1610,In_2194,In_1796);
or U1611 (N_1611,In_1989,In_1446);
nand U1612 (N_1612,In_164,In_1459);
xnor U1613 (N_1613,In_754,In_2675);
or U1614 (N_1614,In_2564,In_2463);
and U1615 (N_1615,In_386,In_1695);
nor U1616 (N_1616,In_1796,In_2934);
or U1617 (N_1617,In_263,In_1617);
or U1618 (N_1618,In_2010,In_2413);
nor U1619 (N_1619,In_2671,In_2854);
nand U1620 (N_1620,In_2759,In_1379);
and U1621 (N_1621,In_204,In_2304);
nor U1622 (N_1622,In_122,In_1435);
nand U1623 (N_1623,In_377,In_2461);
nor U1624 (N_1624,In_1943,In_1022);
nand U1625 (N_1625,In_1587,In_2486);
xnor U1626 (N_1626,In_2783,In_2399);
and U1627 (N_1627,In_2572,In_1957);
nor U1628 (N_1628,In_2057,In_2605);
nor U1629 (N_1629,In_110,In_540);
xnor U1630 (N_1630,In_2285,In_1610);
nand U1631 (N_1631,In_2791,In_396);
or U1632 (N_1632,In_675,In_829);
or U1633 (N_1633,In_2352,In_1811);
nor U1634 (N_1634,In_339,In_393);
xnor U1635 (N_1635,In_1052,In_1698);
or U1636 (N_1636,In_2693,In_429);
and U1637 (N_1637,In_1633,In_1427);
or U1638 (N_1638,In_815,In_2554);
nand U1639 (N_1639,In_492,In_518);
nor U1640 (N_1640,In_1506,In_2798);
nor U1641 (N_1641,In_2681,In_17);
and U1642 (N_1642,In_2874,In_2342);
nand U1643 (N_1643,In_1544,In_984);
nand U1644 (N_1644,In_1066,In_2630);
nor U1645 (N_1645,In_337,In_1812);
nor U1646 (N_1646,In_282,In_720);
or U1647 (N_1647,In_8,In_2757);
nand U1648 (N_1648,In_1030,In_1981);
nor U1649 (N_1649,In_2149,In_2873);
nor U1650 (N_1650,In_2438,In_71);
nand U1651 (N_1651,In_2259,In_1476);
and U1652 (N_1652,In_750,In_2973);
xnor U1653 (N_1653,In_1607,In_1831);
xor U1654 (N_1654,In_2048,In_2575);
nor U1655 (N_1655,In_108,In_391);
or U1656 (N_1656,In_1663,In_2712);
and U1657 (N_1657,In_848,In_2206);
nand U1658 (N_1658,In_713,In_201);
or U1659 (N_1659,In_1776,In_2316);
nor U1660 (N_1660,In_1285,In_618);
or U1661 (N_1661,In_538,In_1960);
or U1662 (N_1662,In_154,In_2519);
or U1663 (N_1663,In_2307,In_1812);
and U1664 (N_1664,In_2703,In_1161);
xor U1665 (N_1665,In_425,In_2819);
and U1666 (N_1666,In_1854,In_2313);
nand U1667 (N_1667,In_1916,In_989);
nor U1668 (N_1668,In_377,In_2697);
xor U1669 (N_1669,In_390,In_242);
xor U1670 (N_1670,In_1658,In_1448);
xor U1671 (N_1671,In_1265,In_1041);
nor U1672 (N_1672,In_2793,In_803);
nor U1673 (N_1673,In_1512,In_2950);
nor U1674 (N_1674,In_2147,In_886);
nor U1675 (N_1675,In_929,In_851);
or U1676 (N_1676,In_621,In_1974);
nor U1677 (N_1677,In_545,In_190);
and U1678 (N_1678,In_1510,In_2794);
nor U1679 (N_1679,In_1810,In_1966);
nor U1680 (N_1680,In_1912,In_661);
nand U1681 (N_1681,In_1639,In_2000);
xnor U1682 (N_1682,In_691,In_2173);
and U1683 (N_1683,In_1266,In_1858);
nand U1684 (N_1684,In_2112,In_991);
or U1685 (N_1685,In_2752,In_2841);
or U1686 (N_1686,In_1627,In_2912);
xnor U1687 (N_1687,In_342,In_6);
or U1688 (N_1688,In_1538,In_2634);
nor U1689 (N_1689,In_2333,In_91);
nor U1690 (N_1690,In_2537,In_1115);
nand U1691 (N_1691,In_730,In_2376);
xnor U1692 (N_1692,In_452,In_767);
nand U1693 (N_1693,In_200,In_2842);
nor U1694 (N_1694,In_649,In_1021);
and U1695 (N_1695,In_513,In_2284);
nor U1696 (N_1696,In_2185,In_277);
nand U1697 (N_1697,In_1377,In_544);
nand U1698 (N_1698,In_1226,In_1027);
xnor U1699 (N_1699,In_2117,In_2061);
or U1700 (N_1700,In_1971,In_2425);
or U1701 (N_1701,In_2154,In_2588);
xor U1702 (N_1702,In_1300,In_725);
nor U1703 (N_1703,In_1681,In_145);
nand U1704 (N_1704,In_1258,In_1635);
and U1705 (N_1705,In_2619,In_355);
xor U1706 (N_1706,In_405,In_1263);
and U1707 (N_1707,In_1689,In_1209);
xor U1708 (N_1708,In_1474,In_1488);
and U1709 (N_1709,In_100,In_1285);
nand U1710 (N_1710,In_1166,In_1343);
xnor U1711 (N_1711,In_2480,In_679);
xnor U1712 (N_1712,In_429,In_509);
nor U1713 (N_1713,In_2553,In_1041);
or U1714 (N_1714,In_261,In_1531);
nor U1715 (N_1715,In_211,In_2033);
or U1716 (N_1716,In_802,In_2706);
or U1717 (N_1717,In_2081,In_1865);
nor U1718 (N_1718,In_1001,In_1420);
or U1719 (N_1719,In_1105,In_416);
and U1720 (N_1720,In_1609,In_696);
nor U1721 (N_1721,In_258,In_1462);
nor U1722 (N_1722,In_365,In_1026);
or U1723 (N_1723,In_2557,In_95);
or U1724 (N_1724,In_1415,In_2099);
nor U1725 (N_1725,In_1094,In_861);
xnor U1726 (N_1726,In_1230,In_2875);
nor U1727 (N_1727,In_1511,In_2381);
or U1728 (N_1728,In_2823,In_2260);
nor U1729 (N_1729,In_1820,In_1531);
or U1730 (N_1730,In_1180,In_888);
and U1731 (N_1731,In_274,In_286);
and U1732 (N_1732,In_2558,In_886);
nand U1733 (N_1733,In_2437,In_200);
or U1734 (N_1734,In_1163,In_85);
and U1735 (N_1735,In_645,In_1060);
and U1736 (N_1736,In_470,In_913);
xnor U1737 (N_1737,In_2005,In_2917);
nand U1738 (N_1738,In_2995,In_1502);
xor U1739 (N_1739,In_663,In_1784);
nor U1740 (N_1740,In_188,In_1403);
and U1741 (N_1741,In_1489,In_627);
nor U1742 (N_1742,In_626,In_579);
or U1743 (N_1743,In_1429,In_440);
xor U1744 (N_1744,In_1659,In_2951);
nor U1745 (N_1745,In_17,In_1023);
xnor U1746 (N_1746,In_2279,In_313);
nor U1747 (N_1747,In_148,In_1798);
xnor U1748 (N_1748,In_1120,In_1150);
nor U1749 (N_1749,In_1567,In_615);
and U1750 (N_1750,In_1,In_419);
and U1751 (N_1751,In_839,In_2044);
and U1752 (N_1752,In_1355,In_901);
or U1753 (N_1753,In_2861,In_702);
and U1754 (N_1754,In_2650,In_365);
xnor U1755 (N_1755,In_1885,In_541);
xor U1756 (N_1756,In_1659,In_2243);
nor U1757 (N_1757,In_2339,In_1694);
or U1758 (N_1758,In_995,In_1347);
and U1759 (N_1759,In_686,In_133);
nand U1760 (N_1760,In_1813,In_2682);
nor U1761 (N_1761,In_227,In_1364);
or U1762 (N_1762,In_886,In_2038);
nand U1763 (N_1763,In_1542,In_2827);
xnor U1764 (N_1764,In_877,In_2521);
and U1765 (N_1765,In_815,In_2419);
nand U1766 (N_1766,In_1356,In_72);
nor U1767 (N_1767,In_1156,In_953);
or U1768 (N_1768,In_1887,In_1514);
nor U1769 (N_1769,In_1976,In_697);
xor U1770 (N_1770,In_1315,In_1207);
xnor U1771 (N_1771,In_1616,In_1688);
nand U1772 (N_1772,In_906,In_921);
or U1773 (N_1773,In_1160,In_2950);
xnor U1774 (N_1774,In_2613,In_2913);
or U1775 (N_1775,In_2976,In_1084);
xnor U1776 (N_1776,In_2246,In_1805);
or U1777 (N_1777,In_2520,In_2118);
and U1778 (N_1778,In_2908,In_773);
nand U1779 (N_1779,In_1162,In_2757);
nand U1780 (N_1780,In_2581,In_2683);
nand U1781 (N_1781,In_2133,In_2937);
xor U1782 (N_1782,In_2183,In_824);
nor U1783 (N_1783,In_2153,In_2268);
nand U1784 (N_1784,In_1868,In_1934);
or U1785 (N_1785,In_2076,In_1204);
nand U1786 (N_1786,In_301,In_1714);
xnor U1787 (N_1787,In_825,In_70);
nor U1788 (N_1788,In_174,In_815);
nor U1789 (N_1789,In_386,In_1121);
or U1790 (N_1790,In_744,In_1344);
nor U1791 (N_1791,In_2700,In_731);
or U1792 (N_1792,In_1319,In_28);
and U1793 (N_1793,In_1493,In_1172);
and U1794 (N_1794,In_2070,In_794);
nor U1795 (N_1795,In_2035,In_2313);
and U1796 (N_1796,In_2856,In_2203);
or U1797 (N_1797,In_1170,In_2807);
nand U1798 (N_1798,In_2414,In_1903);
nor U1799 (N_1799,In_1533,In_62);
nand U1800 (N_1800,In_1091,In_1655);
nor U1801 (N_1801,In_1077,In_2490);
and U1802 (N_1802,In_2988,In_934);
nand U1803 (N_1803,In_2557,In_1642);
or U1804 (N_1804,In_1254,In_7);
nor U1805 (N_1805,In_633,In_2878);
nor U1806 (N_1806,In_2113,In_721);
nor U1807 (N_1807,In_2046,In_988);
and U1808 (N_1808,In_2758,In_2443);
xor U1809 (N_1809,In_2388,In_444);
xor U1810 (N_1810,In_2180,In_2426);
xnor U1811 (N_1811,In_23,In_2362);
xor U1812 (N_1812,In_1618,In_2285);
xor U1813 (N_1813,In_2084,In_2293);
and U1814 (N_1814,In_799,In_1749);
nand U1815 (N_1815,In_2252,In_2579);
nand U1816 (N_1816,In_2451,In_541);
nand U1817 (N_1817,In_1201,In_890);
nand U1818 (N_1818,In_563,In_2415);
xor U1819 (N_1819,In_1430,In_1793);
nor U1820 (N_1820,In_2555,In_673);
nor U1821 (N_1821,In_2581,In_2540);
nand U1822 (N_1822,In_156,In_1328);
xor U1823 (N_1823,In_2898,In_979);
or U1824 (N_1824,In_120,In_462);
nand U1825 (N_1825,In_764,In_2966);
and U1826 (N_1826,In_1323,In_1479);
xor U1827 (N_1827,In_2639,In_2776);
nand U1828 (N_1828,In_1111,In_316);
nor U1829 (N_1829,In_424,In_2238);
nor U1830 (N_1830,In_46,In_601);
and U1831 (N_1831,In_44,In_2827);
nand U1832 (N_1832,In_674,In_2575);
nor U1833 (N_1833,In_1092,In_668);
and U1834 (N_1834,In_2637,In_1924);
nor U1835 (N_1835,In_38,In_250);
nand U1836 (N_1836,In_2437,In_1157);
nand U1837 (N_1837,In_2384,In_2003);
nand U1838 (N_1838,In_2923,In_1510);
or U1839 (N_1839,In_1236,In_1815);
and U1840 (N_1840,In_551,In_141);
and U1841 (N_1841,In_1594,In_1633);
xnor U1842 (N_1842,In_204,In_1280);
xor U1843 (N_1843,In_1759,In_2945);
xnor U1844 (N_1844,In_581,In_2700);
xor U1845 (N_1845,In_325,In_578);
and U1846 (N_1846,In_1981,In_2417);
or U1847 (N_1847,In_2354,In_2847);
and U1848 (N_1848,In_2788,In_2118);
xnor U1849 (N_1849,In_2005,In_696);
nor U1850 (N_1850,In_493,In_124);
nand U1851 (N_1851,In_865,In_1423);
and U1852 (N_1852,In_1604,In_72);
xor U1853 (N_1853,In_1928,In_482);
or U1854 (N_1854,In_2603,In_1236);
nand U1855 (N_1855,In_867,In_354);
nand U1856 (N_1856,In_1044,In_748);
nor U1857 (N_1857,In_316,In_610);
nor U1858 (N_1858,In_758,In_2588);
nor U1859 (N_1859,In_724,In_2087);
nor U1860 (N_1860,In_2819,In_2996);
and U1861 (N_1861,In_494,In_1575);
nand U1862 (N_1862,In_2260,In_778);
nor U1863 (N_1863,In_681,In_1664);
and U1864 (N_1864,In_2764,In_1110);
nand U1865 (N_1865,In_990,In_2933);
nor U1866 (N_1866,In_2925,In_1108);
nor U1867 (N_1867,In_2917,In_294);
or U1868 (N_1868,In_2819,In_2857);
xor U1869 (N_1869,In_1733,In_93);
nand U1870 (N_1870,In_160,In_516);
nor U1871 (N_1871,In_1024,In_1518);
nor U1872 (N_1872,In_214,In_2721);
or U1873 (N_1873,In_899,In_1270);
xor U1874 (N_1874,In_1048,In_1034);
nor U1875 (N_1875,In_2060,In_2047);
xor U1876 (N_1876,In_2,In_2551);
or U1877 (N_1877,In_1405,In_1483);
and U1878 (N_1878,In_2041,In_2495);
nor U1879 (N_1879,In_2517,In_745);
nand U1880 (N_1880,In_501,In_1736);
or U1881 (N_1881,In_1319,In_1873);
nor U1882 (N_1882,In_2598,In_808);
xor U1883 (N_1883,In_470,In_327);
nand U1884 (N_1884,In_1964,In_2389);
or U1885 (N_1885,In_2338,In_1116);
xor U1886 (N_1886,In_2276,In_335);
or U1887 (N_1887,In_1356,In_1160);
nand U1888 (N_1888,In_2296,In_1520);
and U1889 (N_1889,In_1199,In_2108);
and U1890 (N_1890,In_1289,In_114);
or U1891 (N_1891,In_136,In_576);
and U1892 (N_1892,In_1728,In_2488);
nor U1893 (N_1893,In_2309,In_1084);
nand U1894 (N_1894,In_586,In_567);
nor U1895 (N_1895,In_72,In_85);
nor U1896 (N_1896,In_137,In_2993);
xor U1897 (N_1897,In_955,In_1568);
nor U1898 (N_1898,In_2054,In_1010);
and U1899 (N_1899,In_2938,In_635);
xnor U1900 (N_1900,In_2611,In_2555);
or U1901 (N_1901,In_1252,In_18);
or U1902 (N_1902,In_1726,In_476);
xor U1903 (N_1903,In_713,In_2351);
nor U1904 (N_1904,In_395,In_2580);
xor U1905 (N_1905,In_1008,In_1480);
or U1906 (N_1906,In_177,In_1641);
nand U1907 (N_1907,In_2971,In_820);
and U1908 (N_1908,In_711,In_490);
nor U1909 (N_1909,In_1500,In_323);
xor U1910 (N_1910,In_1593,In_1057);
and U1911 (N_1911,In_98,In_1765);
or U1912 (N_1912,In_505,In_1921);
nand U1913 (N_1913,In_688,In_211);
nand U1914 (N_1914,In_1833,In_747);
and U1915 (N_1915,In_1159,In_478);
xor U1916 (N_1916,In_2441,In_2655);
and U1917 (N_1917,In_2003,In_802);
or U1918 (N_1918,In_2071,In_1965);
xor U1919 (N_1919,In_2957,In_1244);
or U1920 (N_1920,In_568,In_1657);
xor U1921 (N_1921,In_2416,In_497);
xnor U1922 (N_1922,In_1298,In_1635);
nand U1923 (N_1923,In_166,In_438);
or U1924 (N_1924,In_659,In_2966);
xor U1925 (N_1925,In_801,In_2082);
nor U1926 (N_1926,In_1541,In_1511);
and U1927 (N_1927,In_291,In_2310);
or U1928 (N_1928,In_2250,In_1321);
xnor U1929 (N_1929,In_2138,In_702);
or U1930 (N_1930,In_984,In_1348);
nor U1931 (N_1931,In_99,In_2745);
xnor U1932 (N_1932,In_2856,In_929);
xnor U1933 (N_1933,In_2014,In_1777);
and U1934 (N_1934,In_2130,In_277);
xnor U1935 (N_1935,In_881,In_2269);
nand U1936 (N_1936,In_775,In_219);
xor U1937 (N_1937,In_513,In_2952);
nor U1938 (N_1938,In_2200,In_588);
and U1939 (N_1939,In_1808,In_1843);
or U1940 (N_1940,In_2876,In_752);
and U1941 (N_1941,In_1714,In_820);
xor U1942 (N_1942,In_382,In_1601);
and U1943 (N_1943,In_833,In_1445);
nor U1944 (N_1944,In_409,In_2857);
or U1945 (N_1945,In_1344,In_86);
and U1946 (N_1946,In_2581,In_2405);
nor U1947 (N_1947,In_1068,In_1468);
and U1948 (N_1948,In_2574,In_2474);
xor U1949 (N_1949,In_487,In_262);
nor U1950 (N_1950,In_228,In_1130);
xor U1951 (N_1951,In_1102,In_1634);
or U1952 (N_1952,In_1836,In_946);
or U1953 (N_1953,In_2741,In_214);
nor U1954 (N_1954,In_2296,In_2140);
or U1955 (N_1955,In_146,In_1312);
and U1956 (N_1956,In_278,In_2162);
xnor U1957 (N_1957,In_1429,In_2395);
and U1958 (N_1958,In_691,In_1315);
and U1959 (N_1959,In_2351,In_2164);
nand U1960 (N_1960,In_2131,In_2533);
nand U1961 (N_1961,In_2370,In_453);
and U1962 (N_1962,In_712,In_1518);
or U1963 (N_1963,In_2438,In_795);
xor U1964 (N_1964,In_1395,In_2729);
nor U1965 (N_1965,In_1342,In_1185);
xnor U1966 (N_1966,In_1043,In_1463);
or U1967 (N_1967,In_347,In_2772);
and U1968 (N_1968,In_708,In_234);
nand U1969 (N_1969,In_1090,In_836);
nor U1970 (N_1970,In_1107,In_2704);
or U1971 (N_1971,In_1461,In_2806);
or U1972 (N_1972,In_2010,In_84);
xor U1973 (N_1973,In_320,In_2361);
and U1974 (N_1974,In_606,In_1514);
and U1975 (N_1975,In_128,In_2965);
and U1976 (N_1976,In_1480,In_72);
xor U1977 (N_1977,In_354,In_521);
or U1978 (N_1978,In_1289,In_1684);
or U1979 (N_1979,In_1945,In_2506);
nand U1980 (N_1980,In_1422,In_2754);
xor U1981 (N_1981,In_911,In_2571);
nor U1982 (N_1982,In_130,In_2591);
or U1983 (N_1983,In_2267,In_632);
nor U1984 (N_1984,In_2551,In_373);
and U1985 (N_1985,In_2808,In_531);
or U1986 (N_1986,In_595,In_526);
nand U1987 (N_1987,In_1741,In_234);
nand U1988 (N_1988,In_2728,In_1590);
and U1989 (N_1989,In_2115,In_1761);
nor U1990 (N_1990,In_1837,In_1611);
or U1991 (N_1991,In_258,In_2706);
xnor U1992 (N_1992,In_449,In_341);
and U1993 (N_1993,In_168,In_445);
xnor U1994 (N_1994,In_1523,In_3);
nor U1995 (N_1995,In_2202,In_1192);
or U1996 (N_1996,In_2197,In_2593);
xor U1997 (N_1997,In_2498,In_1361);
nand U1998 (N_1998,In_1745,In_1490);
xnor U1999 (N_1999,In_1690,In_2534);
nor U2000 (N_2000,In_1554,In_2153);
nand U2001 (N_2001,In_515,In_2588);
nand U2002 (N_2002,In_1926,In_2301);
xor U2003 (N_2003,In_453,In_980);
nor U2004 (N_2004,In_2089,In_108);
nor U2005 (N_2005,In_1936,In_1246);
nor U2006 (N_2006,In_2338,In_2599);
and U2007 (N_2007,In_462,In_2856);
or U2008 (N_2008,In_2949,In_2065);
xnor U2009 (N_2009,In_1974,In_2074);
nor U2010 (N_2010,In_1343,In_638);
or U2011 (N_2011,In_2404,In_2982);
and U2012 (N_2012,In_2364,In_481);
xor U2013 (N_2013,In_1070,In_1622);
and U2014 (N_2014,In_1278,In_1363);
or U2015 (N_2015,In_1821,In_2584);
or U2016 (N_2016,In_1084,In_229);
nand U2017 (N_2017,In_1158,In_1324);
and U2018 (N_2018,In_1961,In_593);
and U2019 (N_2019,In_1152,In_627);
or U2020 (N_2020,In_268,In_540);
nand U2021 (N_2021,In_1033,In_1134);
xnor U2022 (N_2022,In_2975,In_878);
nand U2023 (N_2023,In_994,In_2174);
and U2024 (N_2024,In_1500,In_2008);
nand U2025 (N_2025,In_889,In_2636);
nand U2026 (N_2026,In_2485,In_1140);
xnor U2027 (N_2027,In_45,In_282);
nor U2028 (N_2028,In_2144,In_2941);
nand U2029 (N_2029,In_2563,In_1498);
nand U2030 (N_2030,In_751,In_2581);
and U2031 (N_2031,In_1180,In_1790);
nand U2032 (N_2032,In_1132,In_2228);
nor U2033 (N_2033,In_1555,In_209);
nor U2034 (N_2034,In_386,In_2428);
and U2035 (N_2035,In_962,In_2353);
or U2036 (N_2036,In_1232,In_1086);
and U2037 (N_2037,In_781,In_775);
and U2038 (N_2038,In_1289,In_2247);
nand U2039 (N_2039,In_1218,In_2950);
nor U2040 (N_2040,In_569,In_2415);
xnor U2041 (N_2041,In_2004,In_891);
or U2042 (N_2042,In_971,In_2069);
and U2043 (N_2043,In_2899,In_2411);
xor U2044 (N_2044,In_2789,In_2303);
or U2045 (N_2045,In_1794,In_1132);
nor U2046 (N_2046,In_369,In_2244);
xor U2047 (N_2047,In_680,In_2332);
nor U2048 (N_2048,In_2208,In_1372);
xnor U2049 (N_2049,In_980,In_1774);
nor U2050 (N_2050,In_1701,In_336);
xnor U2051 (N_2051,In_2070,In_722);
xor U2052 (N_2052,In_959,In_1667);
nand U2053 (N_2053,In_141,In_806);
or U2054 (N_2054,In_2515,In_2613);
and U2055 (N_2055,In_303,In_1313);
nor U2056 (N_2056,In_104,In_1471);
or U2057 (N_2057,In_241,In_1211);
and U2058 (N_2058,In_1049,In_2328);
and U2059 (N_2059,In_954,In_1012);
or U2060 (N_2060,In_2543,In_1893);
xor U2061 (N_2061,In_1652,In_2976);
nand U2062 (N_2062,In_1376,In_2896);
nand U2063 (N_2063,In_2698,In_2562);
nor U2064 (N_2064,In_2541,In_1110);
and U2065 (N_2065,In_37,In_1543);
xnor U2066 (N_2066,In_389,In_645);
or U2067 (N_2067,In_2180,In_979);
nand U2068 (N_2068,In_57,In_1773);
xor U2069 (N_2069,In_1070,In_2360);
and U2070 (N_2070,In_720,In_2418);
xor U2071 (N_2071,In_941,In_1897);
and U2072 (N_2072,In_1786,In_1484);
nor U2073 (N_2073,In_651,In_501);
xor U2074 (N_2074,In_1893,In_814);
xnor U2075 (N_2075,In_722,In_2670);
nor U2076 (N_2076,In_103,In_2367);
nor U2077 (N_2077,In_1426,In_1422);
nor U2078 (N_2078,In_1295,In_2704);
xor U2079 (N_2079,In_382,In_1419);
nand U2080 (N_2080,In_1272,In_854);
and U2081 (N_2081,In_2972,In_2642);
and U2082 (N_2082,In_2496,In_2974);
nand U2083 (N_2083,In_676,In_2637);
nor U2084 (N_2084,In_1083,In_1106);
nor U2085 (N_2085,In_236,In_18);
and U2086 (N_2086,In_2364,In_1492);
nand U2087 (N_2087,In_2309,In_314);
and U2088 (N_2088,In_469,In_2781);
and U2089 (N_2089,In_170,In_1471);
nand U2090 (N_2090,In_295,In_2517);
and U2091 (N_2091,In_1621,In_105);
xnor U2092 (N_2092,In_1587,In_913);
or U2093 (N_2093,In_654,In_2349);
xor U2094 (N_2094,In_2476,In_1439);
nand U2095 (N_2095,In_2670,In_563);
or U2096 (N_2096,In_2191,In_2010);
xor U2097 (N_2097,In_2184,In_870);
xnor U2098 (N_2098,In_692,In_1257);
or U2099 (N_2099,In_1541,In_2565);
nand U2100 (N_2100,In_860,In_2039);
and U2101 (N_2101,In_2096,In_534);
or U2102 (N_2102,In_2742,In_1068);
and U2103 (N_2103,In_857,In_2276);
or U2104 (N_2104,In_1051,In_2889);
nor U2105 (N_2105,In_2322,In_728);
nand U2106 (N_2106,In_1175,In_922);
nor U2107 (N_2107,In_955,In_1957);
nand U2108 (N_2108,In_1927,In_1278);
nor U2109 (N_2109,In_159,In_2549);
nand U2110 (N_2110,In_1218,In_2187);
nand U2111 (N_2111,In_1376,In_1234);
or U2112 (N_2112,In_224,In_755);
nand U2113 (N_2113,In_1603,In_214);
nand U2114 (N_2114,In_2650,In_1472);
or U2115 (N_2115,In_2421,In_2105);
nand U2116 (N_2116,In_2919,In_510);
nor U2117 (N_2117,In_1340,In_1047);
or U2118 (N_2118,In_1390,In_833);
xnor U2119 (N_2119,In_1250,In_908);
xnor U2120 (N_2120,In_1467,In_2588);
nand U2121 (N_2121,In_106,In_785);
and U2122 (N_2122,In_212,In_2840);
nand U2123 (N_2123,In_2708,In_10);
nor U2124 (N_2124,In_1646,In_2968);
or U2125 (N_2125,In_1038,In_312);
or U2126 (N_2126,In_2012,In_918);
or U2127 (N_2127,In_2314,In_775);
nor U2128 (N_2128,In_510,In_642);
or U2129 (N_2129,In_1200,In_918);
nor U2130 (N_2130,In_1585,In_2653);
or U2131 (N_2131,In_1056,In_2560);
nand U2132 (N_2132,In_2510,In_2742);
and U2133 (N_2133,In_541,In_2644);
xnor U2134 (N_2134,In_1032,In_2834);
or U2135 (N_2135,In_38,In_2794);
nor U2136 (N_2136,In_2678,In_1641);
nand U2137 (N_2137,In_1491,In_1870);
and U2138 (N_2138,In_1536,In_1501);
nand U2139 (N_2139,In_2159,In_2141);
nor U2140 (N_2140,In_459,In_503);
or U2141 (N_2141,In_1799,In_2726);
or U2142 (N_2142,In_2943,In_2013);
or U2143 (N_2143,In_2438,In_2762);
or U2144 (N_2144,In_297,In_1437);
or U2145 (N_2145,In_2158,In_1152);
nand U2146 (N_2146,In_454,In_1838);
and U2147 (N_2147,In_2280,In_2552);
nand U2148 (N_2148,In_2033,In_2802);
nand U2149 (N_2149,In_840,In_2693);
nor U2150 (N_2150,In_1997,In_1310);
nand U2151 (N_2151,In_2689,In_1688);
xnor U2152 (N_2152,In_1821,In_1069);
or U2153 (N_2153,In_1496,In_2417);
or U2154 (N_2154,In_148,In_118);
or U2155 (N_2155,In_2825,In_2244);
nand U2156 (N_2156,In_1982,In_2413);
or U2157 (N_2157,In_1139,In_978);
xor U2158 (N_2158,In_1818,In_1257);
and U2159 (N_2159,In_1438,In_965);
and U2160 (N_2160,In_2230,In_2693);
xor U2161 (N_2161,In_948,In_415);
xor U2162 (N_2162,In_2137,In_2916);
nand U2163 (N_2163,In_358,In_426);
xor U2164 (N_2164,In_2494,In_2562);
xnor U2165 (N_2165,In_1901,In_814);
xor U2166 (N_2166,In_2576,In_2387);
xnor U2167 (N_2167,In_267,In_1650);
and U2168 (N_2168,In_1235,In_2114);
xnor U2169 (N_2169,In_1808,In_1868);
xnor U2170 (N_2170,In_1504,In_2557);
or U2171 (N_2171,In_1856,In_1719);
nor U2172 (N_2172,In_797,In_60);
or U2173 (N_2173,In_972,In_2738);
xnor U2174 (N_2174,In_2665,In_2739);
xnor U2175 (N_2175,In_353,In_1179);
nand U2176 (N_2176,In_375,In_1937);
and U2177 (N_2177,In_2347,In_464);
nor U2178 (N_2178,In_2612,In_1983);
nand U2179 (N_2179,In_154,In_2619);
nand U2180 (N_2180,In_1423,In_1480);
xor U2181 (N_2181,In_269,In_2467);
xnor U2182 (N_2182,In_902,In_2940);
nand U2183 (N_2183,In_1267,In_1541);
or U2184 (N_2184,In_1634,In_1076);
nand U2185 (N_2185,In_1410,In_2705);
nand U2186 (N_2186,In_799,In_2876);
nand U2187 (N_2187,In_1606,In_1113);
or U2188 (N_2188,In_1048,In_2445);
nand U2189 (N_2189,In_347,In_1974);
and U2190 (N_2190,In_1879,In_1345);
nand U2191 (N_2191,In_1182,In_1255);
nor U2192 (N_2192,In_1577,In_1223);
nor U2193 (N_2193,In_1867,In_386);
and U2194 (N_2194,In_1982,In_454);
and U2195 (N_2195,In_563,In_615);
xor U2196 (N_2196,In_945,In_104);
or U2197 (N_2197,In_1111,In_2834);
or U2198 (N_2198,In_2103,In_996);
or U2199 (N_2199,In_1204,In_1284);
xnor U2200 (N_2200,In_652,In_943);
nand U2201 (N_2201,In_1323,In_2094);
and U2202 (N_2202,In_2323,In_2489);
or U2203 (N_2203,In_920,In_1128);
nor U2204 (N_2204,In_2362,In_271);
xor U2205 (N_2205,In_2771,In_2849);
nand U2206 (N_2206,In_2440,In_2376);
nor U2207 (N_2207,In_786,In_1296);
and U2208 (N_2208,In_1722,In_876);
nand U2209 (N_2209,In_2363,In_143);
and U2210 (N_2210,In_2182,In_1076);
nor U2211 (N_2211,In_2654,In_56);
nor U2212 (N_2212,In_1123,In_2231);
nand U2213 (N_2213,In_2809,In_948);
nand U2214 (N_2214,In_2132,In_2559);
or U2215 (N_2215,In_1905,In_57);
or U2216 (N_2216,In_1308,In_695);
nand U2217 (N_2217,In_2233,In_552);
nor U2218 (N_2218,In_1586,In_1043);
and U2219 (N_2219,In_1563,In_1637);
and U2220 (N_2220,In_1999,In_2245);
nor U2221 (N_2221,In_579,In_723);
nand U2222 (N_2222,In_2535,In_1595);
nor U2223 (N_2223,In_399,In_1903);
xnor U2224 (N_2224,In_2963,In_2568);
or U2225 (N_2225,In_2053,In_492);
xnor U2226 (N_2226,In_1834,In_243);
xor U2227 (N_2227,In_2268,In_1068);
or U2228 (N_2228,In_2305,In_620);
or U2229 (N_2229,In_2405,In_2681);
or U2230 (N_2230,In_1243,In_873);
xor U2231 (N_2231,In_1921,In_1168);
nor U2232 (N_2232,In_1658,In_1427);
xnor U2233 (N_2233,In_2880,In_1555);
xor U2234 (N_2234,In_81,In_1826);
nor U2235 (N_2235,In_356,In_596);
and U2236 (N_2236,In_121,In_1005);
nand U2237 (N_2237,In_883,In_122);
nor U2238 (N_2238,In_2099,In_2773);
nor U2239 (N_2239,In_822,In_2636);
nand U2240 (N_2240,In_750,In_436);
nand U2241 (N_2241,In_259,In_2842);
nor U2242 (N_2242,In_812,In_2948);
and U2243 (N_2243,In_1807,In_665);
and U2244 (N_2244,In_1952,In_113);
or U2245 (N_2245,In_2495,In_231);
nand U2246 (N_2246,In_2081,In_184);
or U2247 (N_2247,In_1162,In_2617);
xor U2248 (N_2248,In_2266,In_1501);
or U2249 (N_2249,In_2913,In_2363);
or U2250 (N_2250,In_364,In_1360);
nor U2251 (N_2251,In_1751,In_2755);
and U2252 (N_2252,In_2930,In_1248);
nor U2253 (N_2253,In_2901,In_1317);
nor U2254 (N_2254,In_2830,In_1359);
and U2255 (N_2255,In_419,In_1183);
nand U2256 (N_2256,In_1232,In_8);
and U2257 (N_2257,In_2258,In_1105);
xor U2258 (N_2258,In_2888,In_2918);
and U2259 (N_2259,In_829,In_1104);
and U2260 (N_2260,In_681,In_2374);
and U2261 (N_2261,In_2682,In_1844);
nand U2262 (N_2262,In_2290,In_690);
xnor U2263 (N_2263,In_1680,In_1468);
and U2264 (N_2264,In_1672,In_593);
and U2265 (N_2265,In_2900,In_2320);
nor U2266 (N_2266,In_2152,In_2655);
xnor U2267 (N_2267,In_308,In_929);
nor U2268 (N_2268,In_589,In_1598);
nand U2269 (N_2269,In_1274,In_2387);
and U2270 (N_2270,In_460,In_1940);
nand U2271 (N_2271,In_1097,In_1710);
nor U2272 (N_2272,In_41,In_2073);
or U2273 (N_2273,In_2092,In_716);
nor U2274 (N_2274,In_1394,In_2804);
nor U2275 (N_2275,In_1818,In_1688);
nand U2276 (N_2276,In_1111,In_1734);
nand U2277 (N_2277,In_1426,In_679);
nand U2278 (N_2278,In_1980,In_1399);
xnor U2279 (N_2279,In_2909,In_2988);
or U2280 (N_2280,In_2491,In_2661);
or U2281 (N_2281,In_116,In_2436);
and U2282 (N_2282,In_828,In_1099);
xor U2283 (N_2283,In_2236,In_2055);
nor U2284 (N_2284,In_58,In_1872);
nand U2285 (N_2285,In_1134,In_1761);
or U2286 (N_2286,In_2173,In_1365);
or U2287 (N_2287,In_158,In_840);
or U2288 (N_2288,In_2324,In_2075);
and U2289 (N_2289,In_527,In_794);
and U2290 (N_2290,In_1392,In_1218);
xor U2291 (N_2291,In_2271,In_2939);
xnor U2292 (N_2292,In_1680,In_1563);
xnor U2293 (N_2293,In_1785,In_801);
nor U2294 (N_2294,In_1974,In_1457);
or U2295 (N_2295,In_1614,In_1685);
or U2296 (N_2296,In_852,In_1101);
and U2297 (N_2297,In_873,In_647);
nand U2298 (N_2298,In_1448,In_1543);
xnor U2299 (N_2299,In_2561,In_951);
xnor U2300 (N_2300,In_2585,In_349);
nand U2301 (N_2301,In_129,In_2240);
or U2302 (N_2302,In_2080,In_90);
nor U2303 (N_2303,In_842,In_2042);
nand U2304 (N_2304,In_2842,In_1678);
xor U2305 (N_2305,In_2666,In_383);
nand U2306 (N_2306,In_1172,In_2820);
nor U2307 (N_2307,In_2651,In_724);
nor U2308 (N_2308,In_2873,In_837);
or U2309 (N_2309,In_1847,In_103);
and U2310 (N_2310,In_2109,In_2436);
and U2311 (N_2311,In_1962,In_2019);
nor U2312 (N_2312,In_2618,In_2944);
nor U2313 (N_2313,In_804,In_13);
or U2314 (N_2314,In_2614,In_499);
nand U2315 (N_2315,In_1969,In_2222);
or U2316 (N_2316,In_1220,In_65);
or U2317 (N_2317,In_1947,In_1932);
and U2318 (N_2318,In_972,In_452);
nand U2319 (N_2319,In_603,In_584);
nand U2320 (N_2320,In_2458,In_2540);
xnor U2321 (N_2321,In_1094,In_1513);
and U2322 (N_2322,In_335,In_1639);
or U2323 (N_2323,In_1096,In_4);
or U2324 (N_2324,In_1951,In_2247);
nor U2325 (N_2325,In_851,In_2039);
or U2326 (N_2326,In_494,In_1011);
and U2327 (N_2327,In_1763,In_523);
and U2328 (N_2328,In_820,In_359);
xor U2329 (N_2329,In_436,In_2183);
xnor U2330 (N_2330,In_1140,In_1468);
nor U2331 (N_2331,In_1727,In_2004);
and U2332 (N_2332,In_2058,In_793);
nor U2333 (N_2333,In_620,In_1679);
and U2334 (N_2334,In_2127,In_1925);
and U2335 (N_2335,In_264,In_1214);
nand U2336 (N_2336,In_2642,In_324);
or U2337 (N_2337,In_1633,In_2645);
nand U2338 (N_2338,In_1641,In_1914);
and U2339 (N_2339,In_2566,In_932);
xnor U2340 (N_2340,In_1827,In_1138);
and U2341 (N_2341,In_2888,In_2439);
xnor U2342 (N_2342,In_666,In_2763);
and U2343 (N_2343,In_1627,In_1992);
or U2344 (N_2344,In_487,In_439);
nor U2345 (N_2345,In_1283,In_303);
xnor U2346 (N_2346,In_2657,In_213);
xor U2347 (N_2347,In_1825,In_1271);
xor U2348 (N_2348,In_1337,In_25);
nand U2349 (N_2349,In_1101,In_2783);
nand U2350 (N_2350,In_2746,In_2647);
nor U2351 (N_2351,In_2667,In_2037);
or U2352 (N_2352,In_1069,In_461);
nand U2353 (N_2353,In_2747,In_2572);
xnor U2354 (N_2354,In_1360,In_2361);
nand U2355 (N_2355,In_1325,In_1573);
nand U2356 (N_2356,In_2324,In_1479);
or U2357 (N_2357,In_1387,In_2686);
nor U2358 (N_2358,In_2886,In_626);
xnor U2359 (N_2359,In_2281,In_2182);
and U2360 (N_2360,In_1298,In_1299);
or U2361 (N_2361,In_1835,In_655);
nand U2362 (N_2362,In_2766,In_1329);
nand U2363 (N_2363,In_2419,In_2864);
nand U2364 (N_2364,In_2646,In_473);
or U2365 (N_2365,In_1326,In_1012);
nor U2366 (N_2366,In_2458,In_2726);
or U2367 (N_2367,In_737,In_1884);
nor U2368 (N_2368,In_1474,In_1436);
xor U2369 (N_2369,In_734,In_402);
xnor U2370 (N_2370,In_2483,In_716);
or U2371 (N_2371,In_1119,In_166);
nor U2372 (N_2372,In_1032,In_221);
nor U2373 (N_2373,In_2201,In_2170);
nand U2374 (N_2374,In_2997,In_950);
xor U2375 (N_2375,In_87,In_1882);
and U2376 (N_2376,In_2255,In_2227);
nor U2377 (N_2377,In_473,In_2079);
nand U2378 (N_2378,In_483,In_1058);
xnor U2379 (N_2379,In_978,In_781);
nand U2380 (N_2380,In_1189,In_1969);
xnor U2381 (N_2381,In_2445,In_1263);
xor U2382 (N_2382,In_977,In_1184);
and U2383 (N_2383,In_1228,In_846);
or U2384 (N_2384,In_833,In_2528);
nand U2385 (N_2385,In_1960,In_2809);
nor U2386 (N_2386,In_2903,In_2589);
or U2387 (N_2387,In_1139,In_2645);
nor U2388 (N_2388,In_1762,In_2983);
or U2389 (N_2389,In_612,In_1852);
nor U2390 (N_2390,In_510,In_1526);
nand U2391 (N_2391,In_1752,In_1709);
or U2392 (N_2392,In_2772,In_2981);
or U2393 (N_2393,In_815,In_275);
nor U2394 (N_2394,In_1309,In_59);
xor U2395 (N_2395,In_57,In_2240);
nand U2396 (N_2396,In_2740,In_2587);
and U2397 (N_2397,In_754,In_119);
nor U2398 (N_2398,In_1662,In_2066);
nor U2399 (N_2399,In_1810,In_43);
or U2400 (N_2400,In_1359,In_2878);
and U2401 (N_2401,In_2322,In_93);
or U2402 (N_2402,In_2375,In_2181);
nand U2403 (N_2403,In_2675,In_2172);
nor U2404 (N_2404,In_1713,In_1161);
nor U2405 (N_2405,In_1058,In_913);
nor U2406 (N_2406,In_2719,In_2839);
or U2407 (N_2407,In_1698,In_1763);
and U2408 (N_2408,In_351,In_2225);
xor U2409 (N_2409,In_2986,In_554);
nor U2410 (N_2410,In_2955,In_2749);
or U2411 (N_2411,In_510,In_2400);
or U2412 (N_2412,In_2338,In_238);
and U2413 (N_2413,In_777,In_933);
nand U2414 (N_2414,In_2519,In_910);
or U2415 (N_2415,In_1293,In_2544);
nor U2416 (N_2416,In_2358,In_2192);
xnor U2417 (N_2417,In_2227,In_1476);
and U2418 (N_2418,In_573,In_332);
xor U2419 (N_2419,In_1582,In_1802);
xor U2420 (N_2420,In_2187,In_1830);
xor U2421 (N_2421,In_593,In_240);
nand U2422 (N_2422,In_1397,In_856);
xor U2423 (N_2423,In_1488,In_2941);
xor U2424 (N_2424,In_2705,In_1912);
and U2425 (N_2425,In_2518,In_417);
and U2426 (N_2426,In_2455,In_359);
xnor U2427 (N_2427,In_2961,In_2786);
and U2428 (N_2428,In_388,In_2524);
and U2429 (N_2429,In_2494,In_2361);
and U2430 (N_2430,In_2421,In_1626);
or U2431 (N_2431,In_135,In_2227);
nor U2432 (N_2432,In_2649,In_1827);
xnor U2433 (N_2433,In_1133,In_507);
or U2434 (N_2434,In_1206,In_1697);
or U2435 (N_2435,In_1256,In_678);
xnor U2436 (N_2436,In_1549,In_457);
xnor U2437 (N_2437,In_2071,In_1637);
or U2438 (N_2438,In_770,In_249);
nor U2439 (N_2439,In_2491,In_316);
and U2440 (N_2440,In_1471,In_1868);
xor U2441 (N_2441,In_2568,In_1952);
and U2442 (N_2442,In_1985,In_3);
nand U2443 (N_2443,In_323,In_911);
nand U2444 (N_2444,In_660,In_380);
xnor U2445 (N_2445,In_1149,In_2808);
nand U2446 (N_2446,In_1862,In_193);
nand U2447 (N_2447,In_1847,In_6);
nor U2448 (N_2448,In_803,In_1664);
and U2449 (N_2449,In_2547,In_188);
xor U2450 (N_2450,In_2587,In_2038);
nor U2451 (N_2451,In_278,In_2542);
nand U2452 (N_2452,In_223,In_1247);
nand U2453 (N_2453,In_19,In_438);
nand U2454 (N_2454,In_1119,In_1084);
xor U2455 (N_2455,In_1800,In_924);
xnor U2456 (N_2456,In_1154,In_2810);
nor U2457 (N_2457,In_904,In_1342);
nand U2458 (N_2458,In_10,In_1177);
nand U2459 (N_2459,In_1586,In_2664);
xnor U2460 (N_2460,In_2488,In_2931);
nand U2461 (N_2461,In_2678,In_223);
and U2462 (N_2462,In_717,In_777);
nand U2463 (N_2463,In_322,In_2534);
nor U2464 (N_2464,In_125,In_405);
nand U2465 (N_2465,In_1342,In_490);
and U2466 (N_2466,In_862,In_1932);
nand U2467 (N_2467,In_2442,In_1452);
nand U2468 (N_2468,In_1439,In_645);
nor U2469 (N_2469,In_311,In_485);
xnor U2470 (N_2470,In_1286,In_2238);
nand U2471 (N_2471,In_1810,In_2984);
nor U2472 (N_2472,In_2398,In_1977);
xor U2473 (N_2473,In_2510,In_278);
and U2474 (N_2474,In_2338,In_833);
or U2475 (N_2475,In_942,In_2598);
and U2476 (N_2476,In_314,In_1677);
or U2477 (N_2477,In_1588,In_1072);
xor U2478 (N_2478,In_2618,In_496);
nor U2479 (N_2479,In_2662,In_2343);
and U2480 (N_2480,In_25,In_1199);
nor U2481 (N_2481,In_2194,In_83);
nor U2482 (N_2482,In_1054,In_149);
nand U2483 (N_2483,In_380,In_431);
nor U2484 (N_2484,In_213,In_278);
or U2485 (N_2485,In_2202,In_2762);
or U2486 (N_2486,In_2808,In_2883);
nor U2487 (N_2487,In_2431,In_2087);
nand U2488 (N_2488,In_849,In_1229);
nor U2489 (N_2489,In_2565,In_411);
nand U2490 (N_2490,In_2238,In_2115);
nor U2491 (N_2491,In_1112,In_2907);
or U2492 (N_2492,In_186,In_2504);
nor U2493 (N_2493,In_1477,In_2380);
nor U2494 (N_2494,In_883,In_1408);
or U2495 (N_2495,In_699,In_2739);
nand U2496 (N_2496,In_2046,In_2927);
xnor U2497 (N_2497,In_1690,In_2968);
nand U2498 (N_2498,In_1109,In_249);
nand U2499 (N_2499,In_804,In_1150);
xnor U2500 (N_2500,In_2037,In_1420);
nor U2501 (N_2501,In_2108,In_1405);
xor U2502 (N_2502,In_1248,In_1521);
nand U2503 (N_2503,In_1722,In_554);
and U2504 (N_2504,In_1826,In_2255);
and U2505 (N_2505,In_2639,In_680);
nand U2506 (N_2506,In_1771,In_43);
or U2507 (N_2507,In_1224,In_498);
and U2508 (N_2508,In_1041,In_327);
or U2509 (N_2509,In_774,In_2681);
or U2510 (N_2510,In_2159,In_2797);
and U2511 (N_2511,In_2526,In_892);
and U2512 (N_2512,In_2295,In_2687);
and U2513 (N_2513,In_1257,In_857);
nand U2514 (N_2514,In_1001,In_69);
xnor U2515 (N_2515,In_1997,In_338);
xnor U2516 (N_2516,In_2430,In_522);
or U2517 (N_2517,In_175,In_65);
or U2518 (N_2518,In_2306,In_2064);
or U2519 (N_2519,In_1427,In_596);
nor U2520 (N_2520,In_1462,In_1038);
nor U2521 (N_2521,In_969,In_910);
xor U2522 (N_2522,In_2953,In_1418);
nand U2523 (N_2523,In_1639,In_447);
nor U2524 (N_2524,In_2311,In_2230);
xnor U2525 (N_2525,In_2015,In_1201);
and U2526 (N_2526,In_2574,In_1955);
nand U2527 (N_2527,In_929,In_1556);
or U2528 (N_2528,In_946,In_26);
xnor U2529 (N_2529,In_2464,In_598);
nand U2530 (N_2530,In_1907,In_1016);
or U2531 (N_2531,In_2940,In_880);
xnor U2532 (N_2532,In_2308,In_2995);
or U2533 (N_2533,In_659,In_2167);
xor U2534 (N_2534,In_1256,In_2075);
xnor U2535 (N_2535,In_760,In_2194);
nor U2536 (N_2536,In_2772,In_671);
nand U2537 (N_2537,In_1128,In_2966);
or U2538 (N_2538,In_1398,In_507);
nor U2539 (N_2539,In_1065,In_1868);
nor U2540 (N_2540,In_1267,In_1427);
nand U2541 (N_2541,In_335,In_117);
xor U2542 (N_2542,In_475,In_112);
nand U2543 (N_2543,In_2166,In_2326);
nor U2544 (N_2544,In_2238,In_2917);
and U2545 (N_2545,In_2835,In_790);
nand U2546 (N_2546,In_1686,In_427);
and U2547 (N_2547,In_2730,In_2130);
or U2548 (N_2548,In_1713,In_2632);
xnor U2549 (N_2549,In_2793,In_2526);
nand U2550 (N_2550,In_991,In_967);
or U2551 (N_2551,In_510,In_2702);
xnor U2552 (N_2552,In_1196,In_1660);
xnor U2553 (N_2553,In_456,In_2431);
xnor U2554 (N_2554,In_1850,In_1784);
nor U2555 (N_2555,In_989,In_2387);
nor U2556 (N_2556,In_1545,In_1255);
and U2557 (N_2557,In_2235,In_2598);
xor U2558 (N_2558,In_776,In_2966);
nor U2559 (N_2559,In_108,In_1976);
and U2560 (N_2560,In_1465,In_1689);
nor U2561 (N_2561,In_2993,In_1733);
xnor U2562 (N_2562,In_469,In_825);
or U2563 (N_2563,In_2775,In_1723);
and U2564 (N_2564,In_791,In_1990);
and U2565 (N_2565,In_1386,In_2169);
and U2566 (N_2566,In_2428,In_2963);
or U2567 (N_2567,In_1404,In_850);
nor U2568 (N_2568,In_2082,In_400);
xnor U2569 (N_2569,In_1372,In_205);
and U2570 (N_2570,In_1159,In_1970);
nor U2571 (N_2571,In_2604,In_2839);
xnor U2572 (N_2572,In_264,In_1988);
xor U2573 (N_2573,In_732,In_1214);
nand U2574 (N_2574,In_1880,In_514);
or U2575 (N_2575,In_1124,In_2907);
or U2576 (N_2576,In_367,In_326);
and U2577 (N_2577,In_2100,In_2028);
or U2578 (N_2578,In_2422,In_6);
and U2579 (N_2579,In_1682,In_2321);
xor U2580 (N_2580,In_49,In_887);
nand U2581 (N_2581,In_2180,In_2750);
or U2582 (N_2582,In_2566,In_38);
nor U2583 (N_2583,In_143,In_42);
and U2584 (N_2584,In_1180,In_2212);
nand U2585 (N_2585,In_2834,In_2985);
nor U2586 (N_2586,In_1094,In_1961);
xor U2587 (N_2587,In_1586,In_1721);
xnor U2588 (N_2588,In_1675,In_2872);
or U2589 (N_2589,In_2181,In_2840);
xnor U2590 (N_2590,In_404,In_2574);
nor U2591 (N_2591,In_2281,In_2593);
xor U2592 (N_2592,In_285,In_2020);
nand U2593 (N_2593,In_923,In_248);
xor U2594 (N_2594,In_2188,In_916);
or U2595 (N_2595,In_980,In_702);
nor U2596 (N_2596,In_1574,In_4);
and U2597 (N_2597,In_552,In_2358);
nand U2598 (N_2598,In_2968,In_2866);
and U2599 (N_2599,In_2635,In_1994);
xnor U2600 (N_2600,In_2570,In_2093);
and U2601 (N_2601,In_819,In_2579);
and U2602 (N_2602,In_38,In_2465);
and U2603 (N_2603,In_1576,In_363);
or U2604 (N_2604,In_942,In_152);
and U2605 (N_2605,In_2122,In_322);
nand U2606 (N_2606,In_430,In_540);
and U2607 (N_2607,In_1171,In_1209);
or U2608 (N_2608,In_1265,In_2594);
nand U2609 (N_2609,In_1812,In_878);
xnor U2610 (N_2610,In_2794,In_573);
nor U2611 (N_2611,In_425,In_1081);
nand U2612 (N_2612,In_1400,In_2356);
nand U2613 (N_2613,In_169,In_2215);
and U2614 (N_2614,In_184,In_661);
nor U2615 (N_2615,In_132,In_2471);
nand U2616 (N_2616,In_743,In_2953);
or U2617 (N_2617,In_1294,In_2956);
and U2618 (N_2618,In_1725,In_2097);
or U2619 (N_2619,In_1519,In_1591);
and U2620 (N_2620,In_648,In_134);
xnor U2621 (N_2621,In_520,In_1000);
and U2622 (N_2622,In_2942,In_1350);
nor U2623 (N_2623,In_1206,In_2479);
nor U2624 (N_2624,In_575,In_2826);
or U2625 (N_2625,In_1836,In_388);
xnor U2626 (N_2626,In_2342,In_322);
nand U2627 (N_2627,In_183,In_1730);
nor U2628 (N_2628,In_536,In_1333);
and U2629 (N_2629,In_2597,In_1884);
nand U2630 (N_2630,In_1619,In_1458);
or U2631 (N_2631,In_2032,In_2026);
nand U2632 (N_2632,In_2166,In_2607);
or U2633 (N_2633,In_1969,In_1032);
nor U2634 (N_2634,In_1403,In_715);
or U2635 (N_2635,In_2355,In_2795);
and U2636 (N_2636,In_1300,In_630);
nand U2637 (N_2637,In_1380,In_842);
nand U2638 (N_2638,In_2283,In_2440);
or U2639 (N_2639,In_706,In_820);
xnor U2640 (N_2640,In_2000,In_2154);
nor U2641 (N_2641,In_516,In_1398);
xor U2642 (N_2642,In_299,In_568);
nand U2643 (N_2643,In_2372,In_527);
or U2644 (N_2644,In_2120,In_2869);
xnor U2645 (N_2645,In_435,In_1164);
xnor U2646 (N_2646,In_868,In_2838);
xor U2647 (N_2647,In_654,In_2906);
nor U2648 (N_2648,In_1265,In_1996);
nand U2649 (N_2649,In_2627,In_1287);
and U2650 (N_2650,In_886,In_1757);
xnor U2651 (N_2651,In_879,In_1570);
nor U2652 (N_2652,In_2099,In_2242);
nor U2653 (N_2653,In_294,In_1431);
xnor U2654 (N_2654,In_2055,In_763);
xor U2655 (N_2655,In_2962,In_1433);
nand U2656 (N_2656,In_2050,In_2391);
or U2657 (N_2657,In_150,In_4);
or U2658 (N_2658,In_240,In_19);
or U2659 (N_2659,In_2820,In_889);
xnor U2660 (N_2660,In_521,In_20);
nand U2661 (N_2661,In_2009,In_523);
and U2662 (N_2662,In_2484,In_330);
and U2663 (N_2663,In_2683,In_341);
or U2664 (N_2664,In_2800,In_1304);
nor U2665 (N_2665,In_1713,In_728);
or U2666 (N_2666,In_1127,In_2587);
or U2667 (N_2667,In_1882,In_727);
and U2668 (N_2668,In_89,In_831);
nand U2669 (N_2669,In_2541,In_1344);
and U2670 (N_2670,In_2552,In_410);
nor U2671 (N_2671,In_2301,In_2533);
nand U2672 (N_2672,In_1752,In_430);
and U2673 (N_2673,In_332,In_2327);
nor U2674 (N_2674,In_432,In_1738);
xnor U2675 (N_2675,In_116,In_582);
nor U2676 (N_2676,In_2710,In_1999);
nand U2677 (N_2677,In_1866,In_1063);
xnor U2678 (N_2678,In_424,In_289);
nor U2679 (N_2679,In_656,In_1158);
xnor U2680 (N_2680,In_1467,In_2751);
or U2681 (N_2681,In_2833,In_531);
nor U2682 (N_2682,In_2378,In_2793);
nand U2683 (N_2683,In_1239,In_1610);
nor U2684 (N_2684,In_256,In_665);
and U2685 (N_2685,In_372,In_2758);
or U2686 (N_2686,In_2174,In_2379);
and U2687 (N_2687,In_2846,In_1066);
or U2688 (N_2688,In_1005,In_459);
xor U2689 (N_2689,In_840,In_1035);
or U2690 (N_2690,In_2639,In_2680);
nand U2691 (N_2691,In_976,In_971);
or U2692 (N_2692,In_1034,In_1409);
and U2693 (N_2693,In_1574,In_1169);
nor U2694 (N_2694,In_2787,In_1317);
nand U2695 (N_2695,In_2935,In_469);
nor U2696 (N_2696,In_2415,In_834);
or U2697 (N_2697,In_1427,In_1282);
and U2698 (N_2698,In_2974,In_11);
and U2699 (N_2699,In_2576,In_1649);
xor U2700 (N_2700,In_1294,In_465);
and U2701 (N_2701,In_641,In_1590);
nor U2702 (N_2702,In_100,In_478);
xor U2703 (N_2703,In_483,In_2721);
nand U2704 (N_2704,In_2790,In_1043);
xnor U2705 (N_2705,In_1954,In_696);
and U2706 (N_2706,In_818,In_1829);
or U2707 (N_2707,In_904,In_2707);
nand U2708 (N_2708,In_1962,In_337);
and U2709 (N_2709,In_2766,In_928);
xnor U2710 (N_2710,In_1773,In_452);
and U2711 (N_2711,In_1707,In_1276);
and U2712 (N_2712,In_2739,In_142);
xor U2713 (N_2713,In_927,In_1316);
nor U2714 (N_2714,In_2820,In_2083);
xnor U2715 (N_2715,In_526,In_842);
or U2716 (N_2716,In_416,In_2177);
xnor U2717 (N_2717,In_680,In_568);
xnor U2718 (N_2718,In_2627,In_238);
nor U2719 (N_2719,In_618,In_169);
nand U2720 (N_2720,In_1534,In_2659);
nor U2721 (N_2721,In_891,In_2636);
nor U2722 (N_2722,In_2479,In_1474);
xnor U2723 (N_2723,In_2585,In_1360);
nor U2724 (N_2724,In_79,In_2256);
xnor U2725 (N_2725,In_926,In_1831);
or U2726 (N_2726,In_2799,In_1580);
nand U2727 (N_2727,In_2259,In_909);
nand U2728 (N_2728,In_1539,In_2105);
xnor U2729 (N_2729,In_2805,In_1114);
nand U2730 (N_2730,In_1692,In_1426);
nor U2731 (N_2731,In_1210,In_935);
nor U2732 (N_2732,In_604,In_1112);
nand U2733 (N_2733,In_308,In_280);
nor U2734 (N_2734,In_2861,In_834);
or U2735 (N_2735,In_1198,In_170);
or U2736 (N_2736,In_1797,In_2918);
nand U2737 (N_2737,In_2714,In_711);
nor U2738 (N_2738,In_2359,In_1404);
or U2739 (N_2739,In_1818,In_547);
or U2740 (N_2740,In_1896,In_978);
and U2741 (N_2741,In_546,In_415);
nand U2742 (N_2742,In_368,In_606);
nor U2743 (N_2743,In_836,In_83);
nand U2744 (N_2744,In_989,In_1444);
or U2745 (N_2745,In_957,In_1564);
and U2746 (N_2746,In_585,In_21);
nand U2747 (N_2747,In_540,In_880);
nor U2748 (N_2748,In_367,In_1920);
and U2749 (N_2749,In_2563,In_1282);
nor U2750 (N_2750,In_2484,In_915);
xnor U2751 (N_2751,In_2855,In_579);
nor U2752 (N_2752,In_902,In_1688);
or U2753 (N_2753,In_2401,In_1647);
and U2754 (N_2754,In_225,In_2868);
xor U2755 (N_2755,In_1990,In_921);
or U2756 (N_2756,In_332,In_1934);
or U2757 (N_2757,In_1804,In_1392);
nand U2758 (N_2758,In_1449,In_2509);
xor U2759 (N_2759,In_741,In_1932);
or U2760 (N_2760,In_1391,In_2732);
nor U2761 (N_2761,In_2294,In_278);
xor U2762 (N_2762,In_288,In_1056);
and U2763 (N_2763,In_957,In_819);
nor U2764 (N_2764,In_1474,In_2860);
xor U2765 (N_2765,In_1061,In_2400);
or U2766 (N_2766,In_339,In_522);
nor U2767 (N_2767,In_1659,In_2622);
nand U2768 (N_2768,In_1025,In_886);
or U2769 (N_2769,In_1964,In_2671);
xnor U2770 (N_2770,In_1409,In_1494);
nor U2771 (N_2771,In_2560,In_2984);
xor U2772 (N_2772,In_2208,In_1321);
nand U2773 (N_2773,In_574,In_375);
nor U2774 (N_2774,In_495,In_2973);
nand U2775 (N_2775,In_2142,In_2402);
or U2776 (N_2776,In_652,In_2715);
nand U2777 (N_2777,In_1048,In_459);
nor U2778 (N_2778,In_1624,In_576);
nand U2779 (N_2779,In_2893,In_2321);
nor U2780 (N_2780,In_1076,In_192);
nand U2781 (N_2781,In_1464,In_224);
or U2782 (N_2782,In_1377,In_2122);
nand U2783 (N_2783,In_1805,In_2135);
nor U2784 (N_2784,In_1669,In_1901);
or U2785 (N_2785,In_795,In_1952);
and U2786 (N_2786,In_2883,In_1436);
and U2787 (N_2787,In_1661,In_2898);
xnor U2788 (N_2788,In_1706,In_786);
xor U2789 (N_2789,In_1724,In_1158);
xnor U2790 (N_2790,In_2798,In_1076);
nand U2791 (N_2791,In_1141,In_2471);
or U2792 (N_2792,In_357,In_2476);
and U2793 (N_2793,In_1971,In_1648);
or U2794 (N_2794,In_1096,In_1470);
nor U2795 (N_2795,In_1443,In_2141);
xnor U2796 (N_2796,In_309,In_1413);
nand U2797 (N_2797,In_2243,In_1645);
and U2798 (N_2798,In_77,In_1979);
or U2799 (N_2799,In_1878,In_2863);
nand U2800 (N_2800,In_380,In_916);
or U2801 (N_2801,In_883,In_793);
nor U2802 (N_2802,In_2701,In_603);
or U2803 (N_2803,In_2687,In_2621);
xor U2804 (N_2804,In_787,In_2767);
and U2805 (N_2805,In_1369,In_2932);
xor U2806 (N_2806,In_1230,In_634);
nor U2807 (N_2807,In_2633,In_2075);
and U2808 (N_2808,In_1432,In_2753);
nand U2809 (N_2809,In_2368,In_1098);
nand U2810 (N_2810,In_1222,In_874);
or U2811 (N_2811,In_1987,In_257);
xnor U2812 (N_2812,In_2171,In_1863);
nand U2813 (N_2813,In_1342,In_1384);
and U2814 (N_2814,In_2678,In_838);
nor U2815 (N_2815,In_1995,In_1712);
nand U2816 (N_2816,In_1304,In_2288);
nand U2817 (N_2817,In_1944,In_1362);
or U2818 (N_2818,In_1464,In_2525);
nor U2819 (N_2819,In_296,In_837);
nand U2820 (N_2820,In_740,In_1609);
nand U2821 (N_2821,In_982,In_2963);
nor U2822 (N_2822,In_1646,In_755);
nand U2823 (N_2823,In_493,In_2463);
xnor U2824 (N_2824,In_1065,In_2777);
and U2825 (N_2825,In_2584,In_2346);
nand U2826 (N_2826,In_1219,In_2462);
xnor U2827 (N_2827,In_183,In_1518);
or U2828 (N_2828,In_2111,In_612);
xor U2829 (N_2829,In_1618,In_804);
nand U2830 (N_2830,In_331,In_2805);
xor U2831 (N_2831,In_1282,In_2538);
xor U2832 (N_2832,In_2377,In_2795);
and U2833 (N_2833,In_12,In_1185);
nand U2834 (N_2834,In_12,In_2672);
nand U2835 (N_2835,In_2470,In_457);
nand U2836 (N_2836,In_2168,In_374);
xor U2837 (N_2837,In_2203,In_900);
nand U2838 (N_2838,In_884,In_408);
xnor U2839 (N_2839,In_1039,In_121);
or U2840 (N_2840,In_2267,In_1961);
or U2841 (N_2841,In_2958,In_630);
nand U2842 (N_2842,In_2452,In_1680);
xor U2843 (N_2843,In_1724,In_1692);
and U2844 (N_2844,In_130,In_664);
and U2845 (N_2845,In_2004,In_1726);
xor U2846 (N_2846,In_1252,In_2402);
and U2847 (N_2847,In_1587,In_2740);
nand U2848 (N_2848,In_1628,In_487);
nand U2849 (N_2849,In_2894,In_418);
xnor U2850 (N_2850,In_1247,In_2416);
and U2851 (N_2851,In_1626,In_1144);
nor U2852 (N_2852,In_513,In_910);
and U2853 (N_2853,In_2725,In_908);
xnor U2854 (N_2854,In_1915,In_977);
nand U2855 (N_2855,In_1561,In_669);
and U2856 (N_2856,In_178,In_577);
or U2857 (N_2857,In_122,In_1354);
nor U2858 (N_2858,In_1600,In_488);
xnor U2859 (N_2859,In_288,In_775);
or U2860 (N_2860,In_1587,In_2582);
and U2861 (N_2861,In_17,In_2808);
nor U2862 (N_2862,In_504,In_1836);
and U2863 (N_2863,In_187,In_43);
or U2864 (N_2864,In_2168,In_1919);
or U2865 (N_2865,In_1472,In_952);
and U2866 (N_2866,In_2681,In_1886);
xor U2867 (N_2867,In_2537,In_589);
nor U2868 (N_2868,In_1733,In_51);
xor U2869 (N_2869,In_1255,In_961);
xnor U2870 (N_2870,In_1661,In_2354);
and U2871 (N_2871,In_2219,In_840);
or U2872 (N_2872,In_605,In_971);
nor U2873 (N_2873,In_1815,In_447);
nor U2874 (N_2874,In_1110,In_293);
and U2875 (N_2875,In_1200,In_1930);
nand U2876 (N_2876,In_779,In_2165);
xor U2877 (N_2877,In_2621,In_2034);
nor U2878 (N_2878,In_2447,In_1578);
and U2879 (N_2879,In_1674,In_1552);
nor U2880 (N_2880,In_550,In_1379);
or U2881 (N_2881,In_2977,In_287);
nand U2882 (N_2882,In_2139,In_1841);
or U2883 (N_2883,In_33,In_1334);
or U2884 (N_2884,In_2734,In_1046);
nor U2885 (N_2885,In_262,In_185);
and U2886 (N_2886,In_1959,In_2302);
xnor U2887 (N_2887,In_784,In_2585);
nand U2888 (N_2888,In_2090,In_1040);
nand U2889 (N_2889,In_49,In_296);
nand U2890 (N_2890,In_1283,In_552);
and U2891 (N_2891,In_1358,In_50);
nor U2892 (N_2892,In_2940,In_971);
nand U2893 (N_2893,In_2583,In_777);
or U2894 (N_2894,In_465,In_1058);
and U2895 (N_2895,In_2539,In_1835);
nand U2896 (N_2896,In_2623,In_2527);
xor U2897 (N_2897,In_553,In_1432);
or U2898 (N_2898,In_1788,In_1528);
nor U2899 (N_2899,In_799,In_743);
nor U2900 (N_2900,In_2122,In_1907);
nand U2901 (N_2901,In_768,In_1968);
nor U2902 (N_2902,In_729,In_442);
xor U2903 (N_2903,In_792,In_1367);
nand U2904 (N_2904,In_992,In_1181);
and U2905 (N_2905,In_1238,In_1948);
and U2906 (N_2906,In_1715,In_2198);
xnor U2907 (N_2907,In_428,In_1625);
nor U2908 (N_2908,In_154,In_569);
and U2909 (N_2909,In_293,In_829);
nor U2910 (N_2910,In_2715,In_408);
xnor U2911 (N_2911,In_2208,In_563);
or U2912 (N_2912,In_2080,In_811);
nor U2913 (N_2913,In_722,In_1952);
and U2914 (N_2914,In_139,In_1954);
nand U2915 (N_2915,In_1872,In_322);
nor U2916 (N_2916,In_2802,In_1279);
nor U2917 (N_2917,In_2444,In_1109);
or U2918 (N_2918,In_2020,In_2183);
and U2919 (N_2919,In_284,In_2009);
nand U2920 (N_2920,In_925,In_2633);
and U2921 (N_2921,In_2759,In_378);
nor U2922 (N_2922,In_1352,In_2336);
and U2923 (N_2923,In_105,In_1417);
xnor U2924 (N_2924,In_2241,In_2497);
and U2925 (N_2925,In_2855,In_900);
and U2926 (N_2926,In_2026,In_2875);
xnor U2927 (N_2927,In_877,In_1710);
xor U2928 (N_2928,In_184,In_2927);
and U2929 (N_2929,In_230,In_2858);
nand U2930 (N_2930,In_2590,In_323);
xnor U2931 (N_2931,In_868,In_841);
and U2932 (N_2932,In_2573,In_378);
or U2933 (N_2933,In_578,In_1129);
nand U2934 (N_2934,In_906,In_2149);
nor U2935 (N_2935,In_1273,In_1163);
xnor U2936 (N_2936,In_2274,In_1465);
or U2937 (N_2937,In_701,In_1285);
xor U2938 (N_2938,In_744,In_1264);
xor U2939 (N_2939,In_1120,In_2608);
and U2940 (N_2940,In_122,In_736);
nor U2941 (N_2941,In_593,In_971);
and U2942 (N_2942,In_907,In_1042);
nor U2943 (N_2943,In_1515,In_1734);
nand U2944 (N_2944,In_1048,In_2086);
nand U2945 (N_2945,In_1038,In_58);
nor U2946 (N_2946,In_495,In_2185);
and U2947 (N_2947,In_20,In_2761);
and U2948 (N_2948,In_1539,In_1603);
or U2949 (N_2949,In_1020,In_2931);
nand U2950 (N_2950,In_590,In_1721);
or U2951 (N_2951,In_2192,In_589);
nand U2952 (N_2952,In_888,In_1212);
xnor U2953 (N_2953,In_2335,In_168);
and U2954 (N_2954,In_1352,In_1877);
xor U2955 (N_2955,In_701,In_2788);
nor U2956 (N_2956,In_2357,In_243);
nand U2957 (N_2957,In_2251,In_1022);
nor U2958 (N_2958,In_154,In_2938);
xor U2959 (N_2959,In_1092,In_1403);
nand U2960 (N_2960,In_674,In_508);
xor U2961 (N_2961,In_2193,In_86);
or U2962 (N_2962,In_2480,In_2514);
and U2963 (N_2963,In_2286,In_2770);
and U2964 (N_2964,In_1784,In_2283);
nor U2965 (N_2965,In_1399,In_2523);
xnor U2966 (N_2966,In_1532,In_491);
and U2967 (N_2967,In_1751,In_381);
xnor U2968 (N_2968,In_2687,In_51);
nor U2969 (N_2969,In_253,In_1346);
nand U2970 (N_2970,In_1582,In_2533);
and U2971 (N_2971,In_477,In_324);
and U2972 (N_2972,In_1582,In_395);
xor U2973 (N_2973,In_36,In_2780);
xor U2974 (N_2974,In_2177,In_1219);
or U2975 (N_2975,In_1673,In_1384);
nor U2976 (N_2976,In_2511,In_455);
nor U2977 (N_2977,In_415,In_2987);
nor U2978 (N_2978,In_773,In_343);
or U2979 (N_2979,In_2830,In_193);
xnor U2980 (N_2980,In_988,In_2479);
xor U2981 (N_2981,In_15,In_779);
or U2982 (N_2982,In_496,In_555);
nand U2983 (N_2983,In_2041,In_533);
nor U2984 (N_2984,In_399,In_936);
nor U2985 (N_2985,In_2943,In_1224);
nor U2986 (N_2986,In_47,In_2800);
nand U2987 (N_2987,In_559,In_1870);
xnor U2988 (N_2988,In_746,In_281);
xnor U2989 (N_2989,In_1175,In_1781);
and U2990 (N_2990,In_658,In_1569);
nand U2991 (N_2991,In_1622,In_1494);
xnor U2992 (N_2992,In_2691,In_2041);
or U2993 (N_2993,In_2143,In_195);
and U2994 (N_2994,In_804,In_1977);
or U2995 (N_2995,In_2835,In_521);
and U2996 (N_2996,In_2748,In_1694);
or U2997 (N_2997,In_2733,In_2199);
nand U2998 (N_2998,In_2344,In_197);
or U2999 (N_2999,In_1201,In_2612);
or U3000 (N_3000,In_507,In_2898);
nor U3001 (N_3001,In_241,In_360);
or U3002 (N_3002,In_1807,In_2631);
or U3003 (N_3003,In_1566,In_484);
nor U3004 (N_3004,In_2029,In_2636);
xor U3005 (N_3005,In_1530,In_344);
and U3006 (N_3006,In_271,In_2900);
nand U3007 (N_3007,In_974,In_555);
or U3008 (N_3008,In_2419,In_1336);
xnor U3009 (N_3009,In_2991,In_986);
nor U3010 (N_3010,In_1826,In_1749);
nand U3011 (N_3011,In_1529,In_1016);
and U3012 (N_3012,In_932,In_2240);
or U3013 (N_3013,In_2106,In_2347);
nor U3014 (N_3014,In_2574,In_819);
nand U3015 (N_3015,In_105,In_1525);
nand U3016 (N_3016,In_1214,In_825);
or U3017 (N_3017,In_1355,In_2409);
nor U3018 (N_3018,In_1605,In_1102);
and U3019 (N_3019,In_472,In_687);
or U3020 (N_3020,In_1081,In_2129);
xnor U3021 (N_3021,In_324,In_921);
nand U3022 (N_3022,In_1541,In_863);
and U3023 (N_3023,In_1791,In_2644);
and U3024 (N_3024,In_1755,In_246);
nor U3025 (N_3025,In_1610,In_577);
and U3026 (N_3026,In_2969,In_1387);
nor U3027 (N_3027,In_458,In_2322);
nand U3028 (N_3028,In_170,In_2400);
or U3029 (N_3029,In_161,In_2781);
xor U3030 (N_3030,In_2127,In_2623);
nand U3031 (N_3031,In_1093,In_2765);
or U3032 (N_3032,In_2761,In_867);
or U3033 (N_3033,In_2624,In_1201);
or U3034 (N_3034,In_1077,In_789);
or U3035 (N_3035,In_1705,In_1033);
and U3036 (N_3036,In_2994,In_1619);
or U3037 (N_3037,In_108,In_2497);
and U3038 (N_3038,In_2625,In_2595);
and U3039 (N_3039,In_2814,In_967);
and U3040 (N_3040,In_2962,In_918);
xnor U3041 (N_3041,In_1133,In_2147);
xor U3042 (N_3042,In_810,In_408);
and U3043 (N_3043,In_2542,In_1366);
xnor U3044 (N_3044,In_674,In_2062);
nand U3045 (N_3045,In_1389,In_2795);
nand U3046 (N_3046,In_113,In_285);
and U3047 (N_3047,In_1411,In_269);
or U3048 (N_3048,In_1301,In_2568);
nand U3049 (N_3049,In_2981,In_1183);
nand U3050 (N_3050,In_1559,In_2707);
and U3051 (N_3051,In_1602,In_2877);
nor U3052 (N_3052,In_1892,In_1428);
and U3053 (N_3053,In_40,In_2629);
or U3054 (N_3054,In_1837,In_608);
nor U3055 (N_3055,In_2673,In_993);
nand U3056 (N_3056,In_523,In_279);
xnor U3057 (N_3057,In_865,In_478);
nor U3058 (N_3058,In_600,In_2138);
and U3059 (N_3059,In_2922,In_826);
nor U3060 (N_3060,In_691,In_2163);
and U3061 (N_3061,In_2250,In_1373);
or U3062 (N_3062,In_396,In_435);
and U3063 (N_3063,In_2838,In_361);
nor U3064 (N_3064,In_1610,In_2005);
xnor U3065 (N_3065,In_314,In_2003);
and U3066 (N_3066,In_2939,In_1574);
or U3067 (N_3067,In_1810,In_1958);
or U3068 (N_3068,In_1231,In_315);
and U3069 (N_3069,In_2894,In_2024);
xor U3070 (N_3070,In_2394,In_2157);
and U3071 (N_3071,In_2027,In_137);
nand U3072 (N_3072,In_2004,In_457);
nor U3073 (N_3073,In_2913,In_1210);
xor U3074 (N_3074,In_2650,In_703);
nor U3075 (N_3075,In_1795,In_571);
and U3076 (N_3076,In_533,In_2046);
or U3077 (N_3077,In_853,In_769);
or U3078 (N_3078,In_2735,In_2216);
nand U3079 (N_3079,In_182,In_425);
or U3080 (N_3080,In_368,In_509);
and U3081 (N_3081,In_2066,In_710);
nand U3082 (N_3082,In_1633,In_2736);
and U3083 (N_3083,In_1146,In_1598);
nand U3084 (N_3084,In_1441,In_2677);
and U3085 (N_3085,In_478,In_2488);
or U3086 (N_3086,In_809,In_2980);
nor U3087 (N_3087,In_2187,In_2591);
or U3088 (N_3088,In_2874,In_1575);
or U3089 (N_3089,In_2017,In_337);
and U3090 (N_3090,In_1527,In_2876);
nor U3091 (N_3091,In_2220,In_856);
xnor U3092 (N_3092,In_1423,In_1116);
or U3093 (N_3093,In_706,In_244);
nor U3094 (N_3094,In_446,In_2885);
and U3095 (N_3095,In_2653,In_267);
and U3096 (N_3096,In_704,In_2722);
and U3097 (N_3097,In_743,In_2295);
nand U3098 (N_3098,In_311,In_2825);
xnor U3099 (N_3099,In_2138,In_2142);
nand U3100 (N_3100,In_2117,In_447);
nand U3101 (N_3101,In_2877,In_757);
xnor U3102 (N_3102,In_771,In_137);
or U3103 (N_3103,In_1645,In_1779);
nor U3104 (N_3104,In_1877,In_2181);
nor U3105 (N_3105,In_871,In_1263);
nor U3106 (N_3106,In_2504,In_1038);
xnor U3107 (N_3107,In_551,In_1072);
and U3108 (N_3108,In_161,In_1193);
or U3109 (N_3109,In_1799,In_722);
xor U3110 (N_3110,In_1782,In_2265);
xor U3111 (N_3111,In_352,In_1954);
nor U3112 (N_3112,In_1741,In_2778);
xor U3113 (N_3113,In_2033,In_44);
nand U3114 (N_3114,In_110,In_300);
and U3115 (N_3115,In_902,In_2934);
nor U3116 (N_3116,In_698,In_80);
and U3117 (N_3117,In_1414,In_1324);
and U3118 (N_3118,In_28,In_1565);
or U3119 (N_3119,In_2860,In_1337);
nand U3120 (N_3120,In_244,In_2663);
nor U3121 (N_3121,In_1936,In_1729);
nand U3122 (N_3122,In_1212,In_2270);
and U3123 (N_3123,In_2354,In_1280);
nand U3124 (N_3124,In_2291,In_597);
xnor U3125 (N_3125,In_2239,In_2606);
or U3126 (N_3126,In_541,In_663);
and U3127 (N_3127,In_746,In_2608);
or U3128 (N_3128,In_1121,In_1052);
nor U3129 (N_3129,In_108,In_446);
nor U3130 (N_3130,In_1111,In_630);
and U3131 (N_3131,In_2894,In_2090);
xor U3132 (N_3132,In_2910,In_2529);
nand U3133 (N_3133,In_553,In_2161);
or U3134 (N_3134,In_1568,In_2951);
nor U3135 (N_3135,In_1742,In_2068);
and U3136 (N_3136,In_2490,In_1326);
xor U3137 (N_3137,In_1433,In_887);
nand U3138 (N_3138,In_1628,In_2648);
or U3139 (N_3139,In_2137,In_102);
or U3140 (N_3140,In_1278,In_1763);
nand U3141 (N_3141,In_1870,In_2927);
or U3142 (N_3142,In_1843,In_405);
or U3143 (N_3143,In_1804,In_1049);
and U3144 (N_3144,In_2519,In_532);
nand U3145 (N_3145,In_1113,In_1373);
and U3146 (N_3146,In_1071,In_2834);
xnor U3147 (N_3147,In_2360,In_1722);
and U3148 (N_3148,In_1919,In_1676);
xnor U3149 (N_3149,In_2590,In_2195);
xnor U3150 (N_3150,In_2322,In_992);
xnor U3151 (N_3151,In_935,In_1762);
nor U3152 (N_3152,In_758,In_1354);
and U3153 (N_3153,In_522,In_914);
xor U3154 (N_3154,In_1800,In_1448);
xnor U3155 (N_3155,In_934,In_1461);
nand U3156 (N_3156,In_1839,In_628);
nand U3157 (N_3157,In_2483,In_2755);
and U3158 (N_3158,In_1759,In_2070);
xor U3159 (N_3159,In_2112,In_1752);
nor U3160 (N_3160,In_363,In_681);
and U3161 (N_3161,In_2189,In_1309);
nand U3162 (N_3162,In_1049,In_487);
or U3163 (N_3163,In_99,In_2242);
or U3164 (N_3164,In_487,In_536);
xor U3165 (N_3165,In_1099,In_472);
and U3166 (N_3166,In_1081,In_460);
nor U3167 (N_3167,In_284,In_796);
or U3168 (N_3168,In_2260,In_767);
nand U3169 (N_3169,In_2283,In_1613);
or U3170 (N_3170,In_440,In_1238);
and U3171 (N_3171,In_759,In_2564);
nor U3172 (N_3172,In_2392,In_1628);
or U3173 (N_3173,In_576,In_2670);
and U3174 (N_3174,In_1158,In_2213);
and U3175 (N_3175,In_1841,In_1380);
xnor U3176 (N_3176,In_1806,In_623);
or U3177 (N_3177,In_285,In_2075);
xor U3178 (N_3178,In_1836,In_2507);
and U3179 (N_3179,In_2850,In_2874);
nor U3180 (N_3180,In_2045,In_570);
and U3181 (N_3181,In_1388,In_389);
nand U3182 (N_3182,In_1276,In_300);
xor U3183 (N_3183,In_988,In_1248);
nor U3184 (N_3184,In_1948,In_755);
nand U3185 (N_3185,In_1802,In_1110);
nand U3186 (N_3186,In_2089,In_1485);
and U3187 (N_3187,In_294,In_2759);
or U3188 (N_3188,In_1154,In_2266);
nand U3189 (N_3189,In_1630,In_817);
xnor U3190 (N_3190,In_2163,In_951);
nor U3191 (N_3191,In_243,In_2760);
and U3192 (N_3192,In_1164,In_2549);
nand U3193 (N_3193,In_1088,In_1471);
and U3194 (N_3194,In_2602,In_2711);
nor U3195 (N_3195,In_650,In_368);
and U3196 (N_3196,In_694,In_1084);
nand U3197 (N_3197,In_906,In_2822);
xor U3198 (N_3198,In_2936,In_349);
nand U3199 (N_3199,In_311,In_2254);
nor U3200 (N_3200,In_1185,In_818);
xnor U3201 (N_3201,In_1357,In_1444);
and U3202 (N_3202,In_2780,In_2452);
xnor U3203 (N_3203,In_1784,In_2762);
nand U3204 (N_3204,In_2568,In_2931);
and U3205 (N_3205,In_1441,In_1282);
and U3206 (N_3206,In_2711,In_729);
xnor U3207 (N_3207,In_2579,In_2661);
nand U3208 (N_3208,In_1558,In_1146);
nor U3209 (N_3209,In_1507,In_1272);
xor U3210 (N_3210,In_1098,In_1736);
xnor U3211 (N_3211,In_108,In_783);
and U3212 (N_3212,In_1749,In_1870);
xnor U3213 (N_3213,In_774,In_1585);
nand U3214 (N_3214,In_1526,In_1468);
nor U3215 (N_3215,In_2373,In_1155);
xnor U3216 (N_3216,In_208,In_704);
or U3217 (N_3217,In_2082,In_2946);
nor U3218 (N_3218,In_1553,In_508);
nand U3219 (N_3219,In_1830,In_2541);
or U3220 (N_3220,In_1462,In_1223);
xor U3221 (N_3221,In_2789,In_2848);
nor U3222 (N_3222,In_1999,In_344);
or U3223 (N_3223,In_2539,In_1190);
and U3224 (N_3224,In_391,In_1084);
nand U3225 (N_3225,In_1228,In_1955);
nor U3226 (N_3226,In_1626,In_1705);
nand U3227 (N_3227,In_2169,In_2134);
nand U3228 (N_3228,In_2377,In_1277);
or U3229 (N_3229,In_480,In_616);
xnor U3230 (N_3230,In_1469,In_1805);
nor U3231 (N_3231,In_1374,In_2978);
nand U3232 (N_3232,In_2011,In_571);
nand U3233 (N_3233,In_1901,In_129);
and U3234 (N_3234,In_1533,In_353);
or U3235 (N_3235,In_2369,In_1715);
xor U3236 (N_3236,In_1209,In_1413);
and U3237 (N_3237,In_869,In_127);
xor U3238 (N_3238,In_849,In_2932);
and U3239 (N_3239,In_1894,In_1297);
and U3240 (N_3240,In_476,In_1775);
xor U3241 (N_3241,In_744,In_1509);
or U3242 (N_3242,In_1556,In_2073);
xor U3243 (N_3243,In_1820,In_719);
nor U3244 (N_3244,In_149,In_1855);
nor U3245 (N_3245,In_2683,In_2900);
and U3246 (N_3246,In_1942,In_1405);
and U3247 (N_3247,In_1562,In_1991);
and U3248 (N_3248,In_934,In_1345);
and U3249 (N_3249,In_1299,In_1919);
xor U3250 (N_3250,In_2196,In_2260);
or U3251 (N_3251,In_536,In_1437);
and U3252 (N_3252,In_1193,In_1079);
xor U3253 (N_3253,In_1600,In_2630);
nand U3254 (N_3254,In_356,In_2506);
nor U3255 (N_3255,In_2657,In_1795);
or U3256 (N_3256,In_804,In_370);
or U3257 (N_3257,In_786,In_653);
or U3258 (N_3258,In_206,In_2629);
nor U3259 (N_3259,In_995,In_2174);
nand U3260 (N_3260,In_588,In_1010);
xor U3261 (N_3261,In_2468,In_876);
xor U3262 (N_3262,In_1044,In_2748);
nand U3263 (N_3263,In_908,In_1654);
and U3264 (N_3264,In_2780,In_1269);
nor U3265 (N_3265,In_137,In_2241);
nor U3266 (N_3266,In_1503,In_1232);
or U3267 (N_3267,In_2163,In_574);
and U3268 (N_3268,In_359,In_2389);
xor U3269 (N_3269,In_1830,In_2624);
nand U3270 (N_3270,In_122,In_945);
nor U3271 (N_3271,In_1690,In_1743);
and U3272 (N_3272,In_1850,In_1759);
and U3273 (N_3273,In_1147,In_1906);
and U3274 (N_3274,In_2166,In_486);
xnor U3275 (N_3275,In_1166,In_1618);
and U3276 (N_3276,In_1936,In_2238);
and U3277 (N_3277,In_1742,In_1878);
nand U3278 (N_3278,In_965,In_2230);
xor U3279 (N_3279,In_2714,In_2337);
nor U3280 (N_3280,In_2357,In_1014);
nand U3281 (N_3281,In_1318,In_142);
and U3282 (N_3282,In_147,In_1882);
and U3283 (N_3283,In_2870,In_1384);
xor U3284 (N_3284,In_2038,In_1264);
and U3285 (N_3285,In_1699,In_684);
or U3286 (N_3286,In_685,In_782);
xnor U3287 (N_3287,In_1493,In_2982);
and U3288 (N_3288,In_1684,In_487);
xor U3289 (N_3289,In_1672,In_2995);
and U3290 (N_3290,In_1232,In_1750);
and U3291 (N_3291,In_867,In_2270);
xor U3292 (N_3292,In_2008,In_1213);
xnor U3293 (N_3293,In_1085,In_708);
and U3294 (N_3294,In_1851,In_2874);
or U3295 (N_3295,In_981,In_2062);
nand U3296 (N_3296,In_1729,In_2402);
xnor U3297 (N_3297,In_1491,In_1323);
or U3298 (N_3298,In_2772,In_1167);
xor U3299 (N_3299,In_2524,In_1976);
xor U3300 (N_3300,In_630,In_220);
xnor U3301 (N_3301,In_1563,In_272);
xor U3302 (N_3302,In_2406,In_1762);
xor U3303 (N_3303,In_1602,In_1881);
xor U3304 (N_3304,In_1987,In_1121);
nor U3305 (N_3305,In_158,In_534);
nand U3306 (N_3306,In_534,In_1700);
or U3307 (N_3307,In_2498,In_1267);
xor U3308 (N_3308,In_1859,In_1674);
and U3309 (N_3309,In_945,In_962);
xor U3310 (N_3310,In_1526,In_792);
nor U3311 (N_3311,In_1862,In_473);
or U3312 (N_3312,In_728,In_1239);
or U3313 (N_3313,In_1287,In_350);
or U3314 (N_3314,In_2561,In_716);
nor U3315 (N_3315,In_1861,In_1608);
or U3316 (N_3316,In_2944,In_2665);
nor U3317 (N_3317,In_1197,In_269);
nor U3318 (N_3318,In_2117,In_1602);
nand U3319 (N_3319,In_1827,In_105);
or U3320 (N_3320,In_2590,In_2248);
nor U3321 (N_3321,In_2750,In_726);
and U3322 (N_3322,In_169,In_599);
nor U3323 (N_3323,In_2501,In_1995);
nand U3324 (N_3324,In_1664,In_2188);
nor U3325 (N_3325,In_324,In_2157);
nand U3326 (N_3326,In_2332,In_2659);
nor U3327 (N_3327,In_143,In_2311);
or U3328 (N_3328,In_369,In_1393);
or U3329 (N_3329,In_1967,In_2940);
and U3330 (N_3330,In_1758,In_626);
or U3331 (N_3331,In_2074,In_509);
nor U3332 (N_3332,In_2717,In_1371);
nand U3333 (N_3333,In_1480,In_286);
nand U3334 (N_3334,In_2691,In_287);
and U3335 (N_3335,In_2604,In_2178);
or U3336 (N_3336,In_1735,In_2675);
or U3337 (N_3337,In_2236,In_1815);
and U3338 (N_3338,In_597,In_2146);
xnor U3339 (N_3339,In_2978,In_1719);
xnor U3340 (N_3340,In_686,In_2164);
and U3341 (N_3341,In_369,In_1636);
nor U3342 (N_3342,In_563,In_1273);
nor U3343 (N_3343,In_35,In_1714);
or U3344 (N_3344,In_2723,In_1995);
and U3345 (N_3345,In_766,In_2390);
or U3346 (N_3346,In_649,In_574);
nand U3347 (N_3347,In_877,In_185);
or U3348 (N_3348,In_1382,In_2276);
nor U3349 (N_3349,In_100,In_2243);
nor U3350 (N_3350,In_74,In_2282);
and U3351 (N_3351,In_941,In_2773);
or U3352 (N_3352,In_208,In_1325);
xor U3353 (N_3353,In_2464,In_94);
or U3354 (N_3354,In_2582,In_359);
nand U3355 (N_3355,In_735,In_2285);
and U3356 (N_3356,In_2329,In_997);
and U3357 (N_3357,In_1955,In_1760);
nor U3358 (N_3358,In_1355,In_2711);
and U3359 (N_3359,In_1439,In_2619);
nor U3360 (N_3360,In_1958,In_835);
nand U3361 (N_3361,In_1944,In_1983);
nand U3362 (N_3362,In_1932,In_2547);
nor U3363 (N_3363,In_1627,In_2459);
xnor U3364 (N_3364,In_385,In_2761);
xnor U3365 (N_3365,In_217,In_953);
xor U3366 (N_3366,In_70,In_1018);
or U3367 (N_3367,In_294,In_1669);
xor U3368 (N_3368,In_50,In_391);
nor U3369 (N_3369,In_1621,In_388);
nand U3370 (N_3370,In_2676,In_2022);
xor U3371 (N_3371,In_2483,In_787);
xnor U3372 (N_3372,In_2578,In_120);
nand U3373 (N_3373,In_2614,In_805);
nor U3374 (N_3374,In_2185,In_475);
nor U3375 (N_3375,In_1418,In_1740);
and U3376 (N_3376,In_2716,In_1602);
nor U3377 (N_3377,In_1643,In_578);
and U3378 (N_3378,In_1619,In_319);
and U3379 (N_3379,In_1678,In_2751);
nand U3380 (N_3380,In_2428,In_854);
and U3381 (N_3381,In_126,In_1179);
nand U3382 (N_3382,In_2667,In_2646);
or U3383 (N_3383,In_379,In_53);
or U3384 (N_3384,In_2868,In_2830);
nand U3385 (N_3385,In_2692,In_2348);
or U3386 (N_3386,In_1828,In_247);
and U3387 (N_3387,In_956,In_723);
and U3388 (N_3388,In_1329,In_1902);
xnor U3389 (N_3389,In_2168,In_1659);
xnor U3390 (N_3390,In_321,In_1987);
or U3391 (N_3391,In_1552,In_1922);
xnor U3392 (N_3392,In_72,In_1212);
or U3393 (N_3393,In_407,In_797);
nand U3394 (N_3394,In_2923,In_2112);
and U3395 (N_3395,In_690,In_1632);
nor U3396 (N_3396,In_967,In_464);
or U3397 (N_3397,In_504,In_1515);
nand U3398 (N_3398,In_2436,In_1267);
nor U3399 (N_3399,In_1393,In_1997);
nand U3400 (N_3400,In_2716,In_2662);
or U3401 (N_3401,In_2421,In_2397);
or U3402 (N_3402,In_434,In_135);
nand U3403 (N_3403,In_1432,In_2385);
xnor U3404 (N_3404,In_1060,In_1786);
or U3405 (N_3405,In_992,In_2618);
or U3406 (N_3406,In_749,In_1635);
or U3407 (N_3407,In_2025,In_16);
and U3408 (N_3408,In_2712,In_1341);
xnor U3409 (N_3409,In_2214,In_229);
and U3410 (N_3410,In_522,In_2172);
and U3411 (N_3411,In_2135,In_2302);
or U3412 (N_3412,In_2120,In_1534);
and U3413 (N_3413,In_2848,In_831);
or U3414 (N_3414,In_23,In_2929);
and U3415 (N_3415,In_2305,In_294);
xnor U3416 (N_3416,In_2468,In_2019);
or U3417 (N_3417,In_44,In_2498);
xor U3418 (N_3418,In_84,In_239);
xor U3419 (N_3419,In_1190,In_1974);
nand U3420 (N_3420,In_480,In_1406);
nand U3421 (N_3421,In_285,In_1290);
nor U3422 (N_3422,In_2238,In_2956);
nand U3423 (N_3423,In_1028,In_2104);
nor U3424 (N_3424,In_2492,In_316);
nor U3425 (N_3425,In_345,In_1748);
or U3426 (N_3426,In_1973,In_1512);
nand U3427 (N_3427,In_2853,In_866);
and U3428 (N_3428,In_1068,In_2397);
and U3429 (N_3429,In_2273,In_622);
nor U3430 (N_3430,In_2628,In_462);
and U3431 (N_3431,In_230,In_296);
or U3432 (N_3432,In_598,In_818);
and U3433 (N_3433,In_2623,In_1527);
xnor U3434 (N_3434,In_1585,In_1624);
nand U3435 (N_3435,In_939,In_168);
nand U3436 (N_3436,In_2909,In_989);
nor U3437 (N_3437,In_2063,In_280);
nand U3438 (N_3438,In_992,In_1040);
and U3439 (N_3439,In_2443,In_2703);
and U3440 (N_3440,In_39,In_1052);
nand U3441 (N_3441,In_2650,In_2436);
xor U3442 (N_3442,In_1142,In_2123);
or U3443 (N_3443,In_1244,In_1655);
xor U3444 (N_3444,In_2825,In_2482);
nor U3445 (N_3445,In_785,In_465);
or U3446 (N_3446,In_1768,In_1614);
and U3447 (N_3447,In_250,In_1303);
xor U3448 (N_3448,In_1058,In_439);
nand U3449 (N_3449,In_2738,In_2156);
nand U3450 (N_3450,In_713,In_2287);
and U3451 (N_3451,In_356,In_1222);
nor U3452 (N_3452,In_147,In_2235);
nor U3453 (N_3453,In_2672,In_1453);
nand U3454 (N_3454,In_2692,In_339);
nor U3455 (N_3455,In_2614,In_164);
nand U3456 (N_3456,In_965,In_540);
and U3457 (N_3457,In_1495,In_112);
and U3458 (N_3458,In_2185,In_2422);
nand U3459 (N_3459,In_918,In_2302);
or U3460 (N_3460,In_558,In_2323);
xor U3461 (N_3461,In_2457,In_2015);
nand U3462 (N_3462,In_2923,In_2890);
and U3463 (N_3463,In_268,In_682);
or U3464 (N_3464,In_2774,In_2990);
nor U3465 (N_3465,In_1475,In_2320);
nor U3466 (N_3466,In_145,In_707);
xnor U3467 (N_3467,In_689,In_2876);
nor U3468 (N_3468,In_1362,In_2084);
nor U3469 (N_3469,In_2664,In_1311);
and U3470 (N_3470,In_2662,In_2002);
xor U3471 (N_3471,In_1629,In_1226);
nand U3472 (N_3472,In_2276,In_1034);
nor U3473 (N_3473,In_683,In_460);
xnor U3474 (N_3474,In_265,In_1637);
and U3475 (N_3475,In_2040,In_1500);
nand U3476 (N_3476,In_717,In_396);
nand U3477 (N_3477,In_1268,In_1990);
or U3478 (N_3478,In_577,In_1886);
xnor U3479 (N_3479,In_2725,In_2317);
nand U3480 (N_3480,In_1759,In_1298);
nor U3481 (N_3481,In_221,In_2001);
or U3482 (N_3482,In_2728,In_2367);
nand U3483 (N_3483,In_2488,In_2344);
and U3484 (N_3484,In_861,In_2900);
nor U3485 (N_3485,In_1022,In_553);
xnor U3486 (N_3486,In_843,In_344);
nor U3487 (N_3487,In_1065,In_2499);
and U3488 (N_3488,In_1239,In_2780);
or U3489 (N_3489,In_2180,In_2980);
nand U3490 (N_3490,In_2902,In_63);
xnor U3491 (N_3491,In_611,In_2126);
nand U3492 (N_3492,In_108,In_562);
or U3493 (N_3493,In_769,In_2699);
or U3494 (N_3494,In_624,In_446);
nand U3495 (N_3495,In_2928,In_663);
or U3496 (N_3496,In_2851,In_2140);
nand U3497 (N_3497,In_1385,In_1406);
xor U3498 (N_3498,In_472,In_171);
xor U3499 (N_3499,In_142,In_2054);
or U3500 (N_3500,In_2382,In_1352);
nor U3501 (N_3501,In_2275,In_367);
nand U3502 (N_3502,In_1635,In_2197);
nor U3503 (N_3503,In_502,In_2629);
xnor U3504 (N_3504,In_352,In_1855);
xor U3505 (N_3505,In_520,In_2073);
nand U3506 (N_3506,In_409,In_1843);
xnor U3507 (N_3507,In_2037,In_1939);
or U3508 (N_3508,In_2228,In_2080);
and U3509 (N_3509,In_1820,In_2970);
and U3510 (N_3510,In_2031,In_2254);
nor U3511 (N_3511,In_157,In_1071);
nor U3512 (N_3512,In_1679,In_936);
and U3513 (N_3513,In_1718,In_641);
and U3514 (N_3514,In_490,In_2971);
or U3515 (N_3515,In_695,In_391);
and U3516 (N_3516,In_1375,In_2382);
nor U3517 (N_3517,In_1841,In_360);
nor U3518 (N_3518,In_2678,In_1327);
and U3519 (N_3519,In_226,In_1234);
xnor U3520 (N_3520,In_2838,In_2494);
and U3521 (N_3521,In_1226,In_672);
nand U3522 (N_3522,In_2938,In_2405);
xnor U3523 (N_3523,In_1563,In_2322);
xnor U3524 (N_3524,In_2779,In_2232);
nor U3525 (N_3525,In_1857,In_1219);
xnor U3526 (N_3526,In_2750,In_2147);
or U3527 (N_3527,In_1484,In_1527);
and U3528 (N_3528,In_967,In_1636);
nand U3529 (N_3529,In_1697,In_880);
nand U3530 (N_3530,In_96,In_1711);
nand U3531 (N_3531,In_2686,In_1063);
and U3532 (N_3532,In_1735,In_293);
and U3533 (N_3533,In_2203,In_2147);
or U3534 (N_3534,In_1388,In_832);
nor U3535 (N_3535,In_1136,In_695);
nand U3536 (N_3536,In_2053,In_424);
nand U3537 (N_3537,In_2942,In_51);
nor U3538 (N_3538,In_2036,In_757);
or U3539 (N_3539,In_889,In_1078);
and U3540 (N_3540,In_1224,In_313);
nand U3541 (N_3541,In_1675,In_2627);
and U3542 (N_3542,In_209,In_1162);
or U3543 (N_3543,In_2155,In_1870);
nand U3544 (N_3544,In_1865,In_1552);
xor U3545 (N_3545,In_404,In_2077);
and U3546 (N_3546,In_1874,In_2912);
nor U3547 (N_3547,In_2765,In_431);
nor U3548 (N_3548,In_1174,In_2884);
xor U3549 (N_3549,In_207,In_2965);
xnor U3550 (N_3550,In_2797,In_1350);
or U3551 (N_3551,In_723,In_2368);
or U3552 (N_3552,In_190,In_191);
nor U3553 (N_3553,In_1625,In_1901);
and U3554 (N_3554,In_846,In_29);
nor U3555 (N_3555,In_2662,In_2305);
xor U3556 (N_3556,In_898,In_2438);
nor U3557 (N_3557,In_2041,In_2999);
nor U3558 (N_3558,In_1402,In_2469);
and U3559 (N_3559,In_2216,In_2440);
xnor U3560 (N_3560,In_2983,In_882);
nand U3561 (N_3561,In_2509,In_2523);
xnor U3562 (N_3562,In_176,In_2989);
nor U3563 (N_3563,In_1509,In_1182);
nor U3564 (N_3564,In_1969,In_2197);
or U3565 (N_3565,In_1391,In_869);
xnor U3566 (N_3566,In_579,In_232);
or U3567 (N_3567,In_840,In_2831);
xor U3568 (N_3568,In_354,In_2222);
and U3569 (N_3569,In_1324,In_298);
nor U3570 (N_3570,In_2036,In_868);
nand U3571 (N_3571,In_1715,In_2331);
nor U3572 (N_3572,In_2089,In_306);
and U3573 (N_3573,In_427,In_1283);
xor U3574 (N_3574,In_654,In_1348);
or U3575 (N_3575,In_1787,In_2745);
nor U3576 (N_3576,In_2825,In_212);
or U3577 (N_3577,In_1799,In_354);
xnor U3578 (N_3578,In_433,In_1663);
xnor U3579 (N_3579,In_542,In_2899);
nor U3580 (N_3580,In_129,In_289);
or U3581 (N_3581,In_2502,In_2243);
nand U3582 (N_3582,In_2257,In_1094);
nor U3583 (N_3583,In_1530,In_544);
and U3584 (N_3584,In_2511,In_929);
nor U3585 (N_3585,In_219,In_2342);
or U3586 (N_3586,In_2179,In_1287);
nand U3587 (N_3587,In_2308,In_2803);
or U3588 (N_3588,In_2133,In_2768);
xnor U3589 (N_3589,In_2839,In_2864);
or U3590 (N_3590,In_1471,In_2224);
or U3591 (N_3591,In_2790,In_1368);
nor U3592 (N_3592,In_368,In_1012);
and U3593 (N_3593,In_2892,In_1363);
and U3594 (N_3594,In_2213,In_821);
or U3595 (N_3595,In_1220,In_1842);
nand U3596 (N_3596,In_399,In_1837);
xor U3597 (N_3597,In_2933,In_980);
xnor U3598 (N_3598,In_998,In_2889);
xnor U3599 (N_3599,In_601,In_120);
nand U3600 (N_3600,In_2849,In_1183);
and U3601 (N_3601,In_589,In_639);
nand U3602 (N_3602,In_1625,In_471);
and U3603 (N_3603,In_2090,In_1193);
and U3604 (N_3604,In_117,In_2934);
nor U3605 (N_3605,In_2895,In_401);
or U3606 (N_3606,In_2061,In_1741);
and U3607 (N_3607,In_1715,In_37);
nor U3608 (N_3608,In_2717,In_2732);
nand U3609 (N_3609,In_2685,In_2859);
nor U3610 (N_3610,In_2563,In_2072);
nor U3611 (N_3611,In_2372,In_1731);
and U3612 (N_3612,In_2788,In_884);
nor U3613 (N_3613,In_2916,In_1239);
nand U3614 (N_3614,In_320,In_804);
nand U3615 (N_3615,In_2171,In_2574);
xor U3616 (N_3616,In_2969,In_749);
and U3617 (N_3617,In_1725,In_151);
nand U3618 (N_3618,In_2175,In_2276);
or U3619 (N_3619,In_2983,In_2289);
or U3620 (N_3620,In_1412,In_1798);
and U3621 (N_3621,In_1508,In_2072);
or U3622 (N_3622,In_1757,In_1805);
xnor U3623 (N_3623,In_353,In_325);
and U3624 (N_3624,In_89,In_610);
nor U3625 (N_3625,In_1435,In_1080);
and U3626 (N_3626,In_1729,In_2263);
xor U3627 (N_3627,In_2991,In_1121);
xnor U3628 (N_3628,In_544,In_1294);
xor U3629 (N_3629,In_2709,In_1400);
xnor U3630 (N_3630,In_56,In_2782);
xor U3631 (N_3631,In_161,In_1478);
xor U3632 (N_3632,In_1121,In_1257);
xor U3633 (N_3633,In_2207,In_2926);
and U3634 (N_3634,In_2385,In_1515);
and U3635 (N_3635,In_29,In_2523);
and U3636 (N_3636,In_2969,In_2822);
nor U3637 (N_3637,In_1891,In_2044);
xnor U3638 (N_3638,In_1813,In_861);
nor U3639 (N_3639,In_2524,In_415);
or U3640 (N_3640,In_760,In_2326);
nor U3641 (N_3641,In_223,In_1902);
nor U3642 (N_3642,In_2587,In_1453);
nor U3643 (N_3643,In_1510,In_1549);
nand U3644 (N_3644,In_581,In_988);
xor U3645 (N_3645,In_1940,In_175);
nand U3646 (N_3646,In_2388,In_1731);
nor U3647 (N_3647,In_1240,In_2020);
or U3648 (N_3648,In_639,In_1146);
or U3649 (N_3649,In_2413,In_598);
xor U3650 (N_3650,In_287,In_2596);
and U3651 (N_3651,In_96,In_917);
nor U3652 (N_3652,In_1093,In_1950);
nand U3653 (N_3653,In_1044,In_179);
nor U3654 (N_3654,In_689,In_2166);
xnor U3655 (N_3655,In_1106,In_543);
nor U3656 (N_3656,In_605,In_2844);
or U3657 (N_3657,In_1503,In_1447);
nand U3658 (N_3658,In_1117,In_2904);
or U3659 (N_3659,In_329,In_1523);
nand U3660 (N_3660,In_1126,In_1748);
nor U3661 (N_3661,In_1387,In_1804);
nor U3662 (N_3662,In_1703,In_102);
and U3663 (N_3663,In_2129,In_1900);
nor U3664 (N_3664,In_2242,In_149);
and U3665 (N_3665,In_530,In_632);
and U3666 (N_3666,In_1668,In_1435);
xnor U3667 (N_3667,In_1475,In_1575);
or U3668 (N_3668,In_2035,In_2135);
or U3669 (N_3669,In_1559,In_2760);
xnor U3670 (N_3670,In_15,In_1701);
and U3671 (N_3671,In_869,In_1413);
or U3672 (N_3672,In_916,In_1207);
nor U3673 (N_3673,In_2459,In_2491);
and U3674 (N_3674,In_1918,In_2881);
or U3675 (N_3675,In_498,In_1205);
or U3676 (N_3676,In_659,In_806);
xor U3677 (N_3677,In_1857,In_1144);
nor U3678 (N_3678,In_577,In_459);
and U3679 (N_3679,In_445,In_2393);
xor U3680 (N_3680,In_423,In_281);
nand U3681 (N_3681,In_2097,In_595);
and U3682 (N_3682,In_2487,In_1093);
or U3683 (N_3683,In_2359,In_975);
nand U3684 (N_3684,In_354,In_1183);
nor U3685 (N_3685,In_417,In_1208);
or U3686 (N_3686,In_1899,In_1129);
and U3687 (N_3687,In_2767,In_1701);
nor U3688 (N_3688,In_993,In_114);
nor U3689 (N_3689,In_2515,In_2296);
nand U3690 (N_3690,In_1008,In_111);
or U3691 (N_3691,In_2707,In_171);
nor U3692 (N_3692,In_2658,In_283);
xnor U3693 (N_3693,In_442,In_453);
and U3694 (N_3694,In_2212,In_1148);
xnor U3695 (N_3695,In_804,In_1002);
and U3696 (N_3696,In_2294,In_2612);
or U3697 (N_3697,In_1433,In_337);
nor U3698 (N_3698,In_1525,In_2789);
nor U3699 (N_3699,In_2855,In_1398);
and U3700 (N_3700,In_1528,In_1473);
nor U3701 (N_3701,In_235,In_630);
or U3702 (N_3702,In_1318,In_2421);
or U3703 (N_3703,In_1476,In_2184);
xnor U3704 (N_3704,In_515,In_125);
and U3705 (N_3705,In_526,In_2472);
nor U3706 (N_3706,In_2417,In_670);
and U3707 (N_3707,In_2270,In_1235);
and U3708 (N_3708,In_1354,In_479);
and U3709 (N_3709,In_1706,In_1565);
nand U3710 (N_3710,In_811,In_133);
xor U3711 (N_3711,In_2568,In_2240);
and U3712 (N_3712,In_2688,In_1157);
and U3713 (N_3713,In_1282,In_1509);
or U3714 (N_3714,In_927,In_2831);
and U3715 (N_3715,In_2643,In_381);
nor U3716 (N_3716,In_2935,In_2939);
and U3717 (N_3717,In_40,In_1636);
and U3718 (N_3718,In_2091,In_1870);
or U3719 (N_3719,In_815,In_2067);
or U3720 (N_3720,In_2728,In_1005);
and U3721 (N_3721,In_1562,In_306);
xor U3722 (N_3722,In_1467,In_2732);
and U3723 (N_3723,In_2566,In_1243);
nand U3724 (N_3724,In_51,In_2145);
nand U3725 (N_3725,In_936,In_1939);
or U3726 (N_3726,In_1823,In_2761);
xor U3727 (N_3727,In_2465,In_838);
and U3728 (N_3728,In_888,In_498);
xnor U3729 (N_3729,In_1841,In_272);
nand U3730 (N_3730,In_2863,In_1121);
xnor U3731 (N_3731,In_1409,In_692);
and U3732 (N_3732,In_2320,In_2871);
xnor U3733 (N_3733,In_1017,In_1977);
nor U3734 (N_3734,In_2310,In_1392);
xnor U3735 (N_3735,In_1954,In_2213);
nand U3736 (N_3736,In_684,In_2871);
and U3737 (N_3737,In_1949,In_162);
and U3738 (N_3738,In_1607,In_1376);
nand U3739 (N_3739,In_2923,In_1945);
and U3740 (N_3740,In_2671,In_245);
xor U3741 (N_3741,In_1540,In_2429);
nand U3742 (N_3742,In_2173,In_201);
or U3743 (N_3743,In_710,In_2213);
and U3744 (N_3744,In_1958,In_2709);
and U3745 (N_3745,In_1645,In_2726);
xor U3746 (N_3746,In_1513,In_1810);
and U3747 (N_3747,In_1507,In_538);
and U3748 (N_3748,In_2804,In_1430);
nand U3749 (N_3749,In_2131,In_1183);
and U3750 (N_3750,In_2083,In_2290);
nand U3751 (N_3751,In_1494,In_2747);
nand U3752 (N_3752,In_613,In_1054);
xnor U3753 (N_3753,In_2911,In_655);
or U3754 (N_3754,In_222,In_2055);
or U3755 (N_3755,In_1082,In_2313);
and U3756 (N_3756,In_437,In_1346);
and U3757 (N_3757,In_1220,In_1915);
nor U3758 (N_3758,In_2816,In_2200);
xnor U3759 (N_3759,In_2644,In_466);
xnor U3760 (N_3760,In_1699,In_2993);
nor U3761 (N_3761,In_2800,In_1699);
and U3762 (N_3762,In_1106,In_782);
and U3763 (N_3763,In_1966,In_1283);
nand U3764 (N_3764,In_2663,In_336);
nand U3765 (N_3765,In_51,In_867);
nor U3766 (N_3766,In_392,In_2495);
or U3767 (N_3767,In_2990,In_797);
xor U3768 (N_3768,In_1687,In_270);
nand U3769 (N_3769,In_1442,In_541);
and U3770 (N_3770,In_1934,In_244);
or U3771 (N_3771,In_71,In_2719);
and U3772 (N_3772,In_61,In_1488);
nand U3773 (N_3773,In_2849,In_930);
nor U3774 (N_3774,In_96,In_1898);
nand U3775 (N_3775,In_2346,In_227);
or U3776 (N_3776,In_1394,In_1753);
nor U3777 (N_3777,In_2651,In_2293);
or U3778 (N_3778,In_2798,In_280);
or U3779 (N_3779,In_1884,In_2449);
nor U3780 (N_3780,In_111,In_372);
nor U3781 (N_3781,In_1860,In_725);
nand U3782 (N_3782,In_926,In_2055);
nor U3783 (N_3783,In_2882,In_2311);
nand U3784 (N_3784,In_2814,In_1215);
nand U3785 (N_3785,In_2377,In_2934);
or U3786 (N_3786,In_2777,In_1338);
nand U3787 (N_3787,In_2426,In_710);
xnor U3788 (N_3788,In_2544,In_2315);
and U3789 (N_3789,In_2968,In_155);
nand U3790 (N_3790,In_751,In_2468);
nand U3791 (N_3791,In_2477,In_497);
nand U3792 (N_3792,In_2191,In_1151);
or U3793 (N_3793,In_1768,In_2981);
nand U3794 (N_3794,In_1998,In_2235);
or U3795 (N_3795,In_526,In_1400);
nor U3796 (N_3796,In_2437,In_1591);
xnor U3797 (N_3797,In_1134,In_1108);
nand U3798 (N_3798,In_1991,In_1877);
xor U3799 (N_3799,In_1500,In_714);
nor U3800 (N_3800,In_2571,In_1281);
and U3801 (N_3801,In_2009,In_1491);
xnor U3802 (N_3802,In_939,In_589);
xnor U3803 (N_3803,In_1373,In_1147);
nand U3804 (N_3804,In_2067,In_424);
xor U3805 (N_3805,In_2676,In_1939);
and U3806 (N_3806,In_1573,In_187);
nand U3807 (N_3807,In_1614,In_437);
nand U3808 (N_3808,In_2179,In_533);
nand U3809 (N_3809,In_595,In_2773);
and U3810 (N_3810,In_198,In_634);
nand U3811 (N_3811,In_2984,In_1740);
or U3812 (N_3812,In_2840,In_329);
or U3813 (N_3813,In_47,In_1658);
or U3814 (N_3814,In_730,In_1069);
or U3815 (N_3815,In_2186,In_987);
nand U3816 (N_3816,In_1992,In_1301);
nand U3817 (N_3817,In_2399,In_2678);
nand U3818 (N_3818,In_2582,In_1599);
nor U3819 (N_3819,In_841,In_2516);
xor U3820 (N_3820,In_899,In_691);
xor U3821 (N_3821,In_1362,In_1856);
xor U3822 (N_3822,In_657,In_1476);
and U3823 (N_3823,In_203,In_694);
xnor U3824 (N_3824,In_1634,In_960);
and U3825 (N_3825,In_2975,In_1246);
nor U3826 (N_3826,In_193,In_943);
or U3827 (N_3827,In_674,In_258);
nand U3828 (N_3828,In_1850,In_34);
xnor U3829 (N_3829,In_2912,In_1520);
xor U3830 (N_3830,In_1977,In_1009);
xnor U3831 (N_3831,In_2364,In_422);
and U3832 (N_3832,In_670,In_7);
and U3833 (N_3833,In_2556,In_1527);
or U3834 (N_3834,In_1567,In_52);
nor U3835 (N_3835,In_1221,In_2759);
nor U3836 (N_3836,In_1759,In_1877);
xnor U3837 (N_3837,In_1967,In_76);
nor U3838 (N_3838,In_894,In_332);
nor U3839 (N_3839,In_706,In_1959);
nor U3840 (N_3840,In_1778,In_2600);
nor U3841 (N_3841,In_808,In_1632);
nand U3842 (N_3842,In_2197,In_964);
or U3843 (N_3843,In_2821,In_1626);
nor U3844 (N_3844,In_2339,In_761);
xnor U3845 (N_3845,In_1554,In_612);
nand U3846 (N_3846,In_2775,In_2356);
or U3847 (N_3847,In_2321,In_1214);
nand U3848 (N_3848,In_2295,In_1376);
xor U3849 (N_3849,In_2613,In_2283);
and U3850 (N_3850,In_897,In_2555);
or U3851 (N_3851,In_508,In_1774);
or U3852 (N_3852,In_2892,In_1277);
xnor U3853 (N_3853,In_320,In_2996);
or U3854 (N_3854,In_2667,In_1808);
xor U3855 (N_3855,In_104,In_2280);
nor U3856 (N_3856,In_2785,In_883);
or U3857 (N_3857,In_1923,In_2944);
xor U3858 (N_3858,In_1932,In_1137);
nand U3859 (N_3859,In_103,In_2812);
and U3860 (N_3860,In_1588,In_2726);
xor U3861 (N_3861,In_127,In_877);
xnor U3862 (N_3862,In_1469,In_1026);
or U3863 (N_3863,In_2236,In_915);
or U3864 (N_3864,In_1657,In_251);
nor U3865 (N_3865,In_2774,In_2833);
nand U3866 (N_3866,In_485,In_2384);
nand U3867 (N_3867,In_2508,In_897);
nand U3868 (N_3868,In_1853,In_757);
nor U3869 (N_3869,In_2316,In_2710);
nand U3870 (N_3870,In_2427,In_1139);
and U3871 (N_3871,In_1084,In_2002);
or U3872 (N_3872,In_2378,In_512);
nand U3873 (N_3873,In_565,In_931);
nand U3874 (N_3874,In_1453,In_2080);
nor U3875 (N_3875,In_1572,In_1447);
or U3876 (N_3876,In_595,In_1729);
and U3877 (N_3877,In_378,In_1801);
xnor U3878 (N_3878,In_2857,In_525);
and U3879 (N_3879,In_1032,In_1957);
or U3880 (N_3880,In_743,In_2275);
or U3881 (N_3881,In_371,In_2497);
nor U3882 (N_3882,In_2777,In_616);
xor U3883 (N_3883,In_2525,In_964);
nand U3884 (N_3884,In_146,In_990);
or U3885 (N_3885,In_2083,In_2646);
xor U3886 (N_3886,In_599,In_2596);
nor U3887 (N_3887,In_852,In_2589);
xnor U3888 (N_3888,In_944,In_1468);
and U3889 (N_3889,In_2864,In_2979);
nand U3890 (N_3890,In_2032,In_2341);
nand U3891 (N_3891,In_2042,In_2330);
nor U3892 (N_3892,In_344,In_2004);
or U3893 (N_3893,In_970,In_1090);
or U3894 (N_3894,In_2771,In_1233);
and U3895 (N_3895,In_2467,In_1692);
xor U3896 (N_3896,In_1151,In_2152);
xor U3897 (N_3897,In_2964,In_813);
xnor U3898 (N_3898,In_109,In_2787);
and U3899 (N_3899,In_70,In_1954);
xnor U3900 (N_3900,In_2431,In_581);
nand U3901 (N_3901,In_1762,In_1412);
nand U3902 (N_3902,In_1985,In_1933);
nand U3903 (N_3903,In_2751,In_2535);
and U3904 (N_3904,In_1264,In_2396);
nand U3905 (N_3905,In_1252,In_1819);
xor U3906 (N_3906,In_2102,In_749);
or U3907 (N_3907,In_1254,In_2111);
and U3908 (N_3908,In_333,In_776);
or U3909 (N_3909,In_43,In_905);
nand U3910 (N_3910,In_1990,In_709);
nor U3911 (N_3911,In_1330,In_447);
xnor U3912 (N_3912,In_494,In_2547);
nor U3913 (N_3913,In_2373,In_2029);
and U3914 (N_3914,In_1986,In_1333);
or U3915 (N_3915,In_1650,In_1190);
nand U3916 (N_3916,In_2348,In_1029);
or U3917 (N_3917,In_2667,In_2502);
or U3918 (N_3918,In_2700,In_2374);
or U3919 (N_3919,In_1010,In_535);
or U3920 (N_3920,In_1944,In_38);
or U3921 (N_3921,In_2485,In_500);
xnor U3922 (N_3922,In_554,In_581);
nand U3923 (N_3923,In_2854,In_1192);
nor U3924 (N_3924,In_407,In_1250);
or U3925 (N_3925,In_1432,In_2373);
nor U3926 (N_3926,In_1951,In_471);
nand U3927 (N_3927,In_2353,In_805);
nor U3928 (N_3928,In_2952,In_521);
nor U3929 (N_3929,In_2541,In_2614);
nand U3930 (N_3930,In_2426,In_1179);
nor U3931 (N_3931,In_2260,In_2811);
xor U3932 (N_3932,In_1153,In_1798);
nand U3933 (N_3933,In_949,In_2327);
and U3934 (N_3934,In_1276,In_2577);
or U3935 (N_3935,In_2785,In_2047);
nor U3936 (N_3936,In_2195,In_2952);
or U3937 (N_3937,In_2625,In_935);
xnor U3938 (N_3938,In_1887,In_571);
xnor U3939 (N_3939,In_260,In_2556);
xor U3940 (N_3940,In_219,In_2358);
and U3941 (N_3941,In_2982,In_888);
nand U3942 (N_3942,In_1842,In_797);
and U3943 (N_3943,In_2577,In_47);
xor U3944 (N_3944,In_250,In_982);
nand U3945 (N_3945,In_2458,In_1620);
or U3946 (N_3946,In_411,In_1624);
nand U3947 (N_3947,In_1204,In_1004);
nor U3948 (N_3948,In_2795,In_2010);
nand U3949 (N_3949,In_1867,In_1140);
nand U3950 (N_3950,In_2094,In_1306);
and U3951 (N_3951,In_2398,In_2285);
nor U3952 (N_3952,In_1689,In_2372);
or U3953 (N_3953,In_839,In_1270);
nor U3954 (N_3954,In_386,In_2907);
or U3955 (N_3955,In_520,In_2338);
nor U3956 (N_3956,In_1255,In_1498);
nor U3957 (N_3957,In_2108,In_2118);
or U3958 (N_3958,In_354,In_1013);
and U3959 (N_3959,In_2838,In_2084);
nand U3960 (N_3960,In_1892,In_279);
nand U3961 (N_3961,In_2054,In_229);
and U3962 (N_3962,In_2151,In_2433);
nor U3963 (N_3963,In_75,In_441);
or U3964 (N_3964,In_197,In_951);
xnor U3965 (N_3965,In_283,In_1744);
or U3966 (N_3966,In_2062,In_1428);
xor U3967 (N_3967,In_1127,In_2623);
nand U3968 (N_3968,In_2289,In_839);
or U3969 (N_3969,In_1322,In_1771);
xnor U3970 (N_3970,In_383,In_2357);
nand U3971 (N_3971,In_503,In_137);
or U3972 (N_3972,In_453,In_975);
nor U3973 (N_3973,In_1956,In_1460);
nor U3974 (N_3974,In_1878,In_152);
and U3975 (N_3975,In_83,In_570);
nor U3976 (N_3976,In_166,In_1579);
nand U3977 (N_3977,In_2379,In_2646);
nor U3978 (N_3978,In_1184,In_1733);
xor U3979 (N_3979,In_2087,In_2182);
nor U3980 (N_3980,In_1534,In_331);
and U3981 (N_3981,In_1198,In_362);
nand U3982 (N_3982,In_1020,In_2529);
xor U3983 (N_3983,In_1342,In_2453);
and U3984 (N_3984,In_2962,In_387);
and U3985 (N_3985,In_1226,In_1915);
and U3986 (N_3986,In_815,In_1866);
and U3987 (N_3987,In_1868,In_2606);
and U3988 (N_3988,In_2565,In_2381);
nand U3989 (N_3989,In_91,In_1069);
or U3990 (N_3990,In_2454,In_1790);
nor U3991 (N_3991,In_2637,In_1016);
nand U3992 (N_3992,In_2339,In_2126);
nor U3993 (N_3993,In_1655,In_108);
and U3994 (N_3994,In_129,In_1691);
or U3995 (N_3995,In_124,In_2771);
or U3996 (N_3996,In_2923,In_1416);
or U3997 (N_3997,In_748,In_2380);
nand U3998 (N_3998,In_2429,In_1326);
or U3999 (N_3999,In_525,In_1892);
and U4000 (N_4000,In_602,In_2740);
nand U4001 (N_4001,In_448,In_762);
xnor U4002 (N_4002,In_2263,In_2567);
nor U4003 (N_4003,In_342,In_2359);
or U4004 (N_4004,In_388,In_1026);
xor U4005 (N_4005,In_1559,In_2901);
xnor U4006 (N_4006,In_681,In_1894);
and U4007 (N_4007,In_180,In_57);
nor U4008 (N_4008,In_2741,In_404);
and U4009 (N_4009,In_1436,In_1252);
and U4010 (N_4010,In_1671,In_2099);
and U4011 (N_4011,In_1584,In_839);
nand U4012 (N_4012,In_1352,In_1194);
or U4013 (N_4013,In_2019,In_1412);
or U4014 (N_4014,In_130,In_2714);
nor U4015 (N_4015,In_1313,In_2140);
and U4016 (N_4016,In_2426,In_574);
nor U4017 (N_4017,In_658,In_55);
nor U4018 (N_4018,In_706,In_1266);
and U4019 (N_4019,In_1897,In_1376);
and U4020 (N_4020,In_1900,In_756);
nor U4021 (N_4021,In_1252,In_2463);
nor U4022 (N_4022,In_852,In_1447);
xnor U4023 (N_4023,In_1038,In_370);
or U4024 (N_4024,In_580,In_985);
or U4025 (N_4025,In_1684,In_2597);
xor U4026 (N_4026,In_2776,In_1646);
and U4027 (N_4027,In_2709,In_1793);
and U4028 (N_4028,In_181,In_331);
nand U4029 (N_4029,In_1970,In_1436);
and U4030 (N_4030,In_1815,In_266);
and U4031 (N_4031,In_409,In_1251);
and U4032 (N_4032,In_915,In_374);
or U4033 (N_4033,In_1871,In_1944);
nand U4034 (N_4034,In_2371,In_2812);
and U4035 (N_4035,In_2455,In_530);
and U4036 (N_4036,In_2854,In_2668);
xor U4037 (N_4037,In_1325,In_1031);
nor U4038 (N_4038,In_1057,In_1956);
nand U4039 (N_4039,In_992,In_2819);
and U4040 (N_4040,In_2057,In_1255);
nor U4041 (N_4041,In_1266,In_1602);
or U4042 (N_4042,In_632,In_709);
nor U4043 (N_4043,In_1901,In_2409);
or U4044 (N_4044,In_43,In_2504);
nand U4045 (N_4045,In_394,In_2972);
nor U4046 (N_4046,In_1819,In_2569);
xor U4047 (N_4047,In_2970,In_565);
xnor U4048 (N_4048,In_1298,In_2014);
and U4049 (N_4049,In_1642,In_2184);
xnor U4050 (N_4050,In_894,In_1204);
nor U4051 (N_4051,In_2836,In_1040);
nand U4052 (N_4052,In_2025,In_2308);
nand U4053 (N_4053,In_2957,In_2723);
or U4054 (N_4054,In_1888,In_2391);
nor U4055 (N_4055,In_487,In_1156);
or U4056 (N_4056,In_2983,In_1712);
and U4057 (N_4057,In_1334,In_2767);
nand U4058 (N_4058,In_843,In_433);
and U4059 (N_4059,In_764,In_2668);
and U4060 (N_4060,In_2339,In_2708);
or U4061 (N_4061,In_1472,In_1750);
or U4062 (N_4062,In_2217,In_35);
and U4063 (N_4063,In_1955,In_2778);
nand U4064 (N_4064,In_2505,In_1103);
or U4065 (N_4065,In_1477,In_841);
and U4066 (N_4066,In_2347,In_1451);
and U4067 (N_4067,In_923,In_879);
xnor U4068 (N_4068,In_728,In_2227);
xor U4069 (N_4069,In_280,In_63);
nand U4070 (N_4070,In_976,In_454);
and U4071 (N_4071,In_2162,In_995);
xor U4072 (N_4072,In_128,In_2532);
xor U4073 (N_4073,In_2741,In_1332);
or U4074 (N_4074,In_459,In_10);
nor U4075 (N_4075,In_2811,In_702);
xnor U4076 (N_4076,In_516,In_2118);
nor U4077 (N_4077,In_346,In_2819);
xnor U4078 (N_4078,In_1312,In_418);
or U4079 (N_4079,In_1113,In_385);
nand U4080 (N_4080,In_1209,In_895);
and U4081 (N_4081,In_2407,In_2676);
nor U4082 (N_4082,In_1075,In_934);
and U4083 (N_4083,In_2040,In_2581);
or U4084 (N_4084,In_1738,In_787);
xnor U4085 (N_4085,In_555,In_332);
nor U4086 (N_4086,In_2258,In_1996);
xor U4087 (N_4087,In_2026,In_2999);
nor U4088 (N_4088,In_1896,In_2369);
xnor U4089 (N_4089,In_2489,In_499);
nor U4090 (N_4090,In_1903,In_2574);
or U4091 (N_4091,In_2710,In_2511);
or U4092 (N_4092,In_415,In_1576);
xnor U4093 (N_4093,In_2230,In_1030);
or U4094 (N_4094,In_1701,In_2593);
nor U4095 (N_4095,In_2839,In_795);
nor U4096 (N_4096,In_1924,In_2287);
or U4097 (N_4097,In_2437,In_428);
and U4098 (N_4098,In_1625,In_1212);
xnor U4099 (N_4099,In_1237,In_1382);
and U4100 (N_4100,In_1354,In_2448);
xnor U4101 (N_4101,In_1271,In_1555);
and U4102 (N_4102,In_2539,In_335);
xor U4103 (N_4103,In_1752,In_2876);
nand U4104 (N_4104,In_1440,In_537);
xnor U4105 (N_4105,In_1676,In_2191);
nand U4106 (N_4106,In_2505,In_2261);
nor U4107 (N_4107,In_2634,In_647);
xnor U4108 (N_4108,In_13,In_392);
xnor U4109 (N_4109,In_1392,In_977);
xnor U4110 (N_4110,In_500,In_700);
nor U4111 (N_4111,In_2955,In_1103);
nor U4112 (N_4112,In_402,In_1063);
nand U4113 (N_4113,In_240,In_1738);
xnor U4114 (N_4114,In_1453,In_548);
and U4115 (N_4115,In_1330,In_2722);
or U4116 (N_4116,In_1208,In_763);
and U4117 (N_4117,In_1434,In_1287);
nand U4118 (N_4118,In_1430,In_1596);
xor U4119 (N_4119,In_1764,In_1430);
and U4120 (N_4120,In_2773,In_1887);
or U4121 (N_4121,In_170,In_1995);
and U4122 (N_4122,In_531,In_465);
or U4123 (N_4123,In_1665,In_1920);
xor U4124 (N_4124,In_120,In_2875);
or U4125 (N_4125,In_1640,In_46);
nand U4126 (N_4126,In_1033,In_1564);
and U4127 (N_4127,In_1940,In_1571);
nand U4128 (N_4128,In_749,In_1179);
nor U4129 (N_4129,In_2904,In_238);
and U4130 (N_4130,In_666,In_2514);
or U4131 (N_4131,In_2421,In_333);
nor U4132 (N_4132,In_249,In_1540);
nor U4133 (N_4133,In_1695,In_1602);
xor U4134 (N_4134,In_493,In_2995);
xor U4135 (N_4135,In_351,In_848);
nor U4136 (N_4136,In_2736,In_2892);
and U4137 (N_4137,In_227,In_1100);
and U4138 (N_4138,In_1980,In_960);
xor U4139 (N_4139,In_2028,In_1863);
nor U4140 (N_4140,In_2926,In_1972);
nor U4141 (N_4141,In_1600,In_2553);
nor U4142 (N_4142,In_2776,In_1619);
nand U4143 (N_4143,In_208,In_1570);
and U4144 (N_4144,In_1120,In_2709);
and U4145 (N_4145,In_2896,In_2504);
nor U4146 (N_4146,In_288,In_674);
nor U4147 (N_4147,In_2485,In_863);
or U4148 (N_4148,In_2770,In_2966);
nand U4149 (N_4149,In_2268,In_789);
and U4150 (N_4150,In_970,In_2130);
nand U4151 (N_4151,In_41,In_1139);
or U4152 (N_4152,In_1289,In_2041);
xor U4153 (N_4153,In_2364,In_924);
nor U4154 (N_4154,In_1250,In_2501);
and U4155 (N_4155,In_1259,In_2238);
nand U4156 (N_4156,In_1729,In_241);
nand U4157 (N_4157,In_1473,In_2031);
or U4158 (N_4158,In_1576,In_451);
xor U4159 (N_4159,In_605,In_2199);
and U4160 (N_4160,In_2142,In_1250);
nand U4161 (N_4161,In_2488,In_2916);
xnor U4162 (N_4162,In_2082,In_2318);
nor U4163 (N_4163,In_2377,In_2517);
nand U4164 (N_4164,In_2910,In_461);
xnor U4165 (N_4165,In_1890,In_885);
or U4166 (N_4166,In_1091,In_915);
nand U4167 (N_4167,In_2307,In_1135);
and U4168 (N_4168,In_1208,In_107);
nor U4169 (N_4169,In_629,In_1628);
and U4170 (N_4170,In_1598,In_2244);
nand U4171 (N_4171,In_1728,In_2917);
nor U4172 (N_4172,In_181,In_298);
nand U4173 (N_4173,In_1494,In_2159);
nand U4174 (N_4174,In_438,In_709);
nor U4175 (N_4175,In_960,In_959);
xnor U4176 (N_4176,In_2259,In_1703);
or U4177 (N_4177,In_2154,In_2108);
xor U4178 (N_4178,In_2852,In_2681);
xor U4179 (N_4179,In_1993,In_2469);
xnor U4180 (N_4180,In_2799,In_2994);
nand U4181 (N_4181,In_301,In_606);
nor U4182 (N_4182,In_818,In_2212);
and U4183 (N_4183,In_1478,In_2982);
and U4184 (N_4184,In_140,In_1564);
nand U4185 (N_4185,In_1151,In_2002);
xnor U4186 (N_4186,In_1390,In_2302);
and U4187 (N_4187,In_516,In_1972);
or U4188 (N_4188,In_26,In_1283);
or U4189 (N_4189,In_73,In_2062);
nand U4190 (N_4190,In_1238,In_1655);
xnor U4191 (N_4191,In_2632,In_54);
and U4192 (N_4192,In_619,In_2066);
nor U4193 (N_4193,In_23,In_2280);
nand U4194 (N_4194,In_2476,In_2900);
nand U4195 (N_4195,In_1783,In_258);
or U4196 (N_4196,In_881,In_1032);
nor U4197 (N_4197,In_1860,In_1846);
or U4198 (N_4198,In_2180,In_2235);
or U4199 (N_4199,In_1706,In_1763);
and U4200 (N_4200,In_368,In_2597);
nor U4201 (N_4201,In_1107,In_2288);
nor U4202 (N_4202,In_247,In_1752);
or U4203 (N_4203,In_2010,In_922);
nand U4204 (N_4204,In_2658,In_1051);
or U4205 (N_4205,In_880,In_2538);
nand U4206 (N_4206,In_1991,In_2765);
xor U4207 (N_4207,In_462,In_2899);
xor U4208 (N_4208,In_2512,In_1908);
or U4209 (N_4209,In_1810,In_901);
and U4210 (N_4210,In_1553,In_2856);
xnor U4211 (N_4211,In_743,In_1429);
nor U4212 (N_4212,In_2754,In_489);
xor U4213 (N_4213,In_2013,In_1920);
xor U4214 (N_4214,In_1107,In_2294);
xor U4215 (N_4215,In_683,In_2237);
nand U4216 (N_4216,In_2729,In_687);
nor U4217 (N_4217,In_2800,In_2656);
nor U4218 (N_4218,In_111,In_576);
xnor U4219 (N_4219,In_111,In_1109);
xnor U4220 (N_4220,In_1829,In_1108);
and U4221 (N_4221,In_565,In_2812);
nor U4222 (N_4222,In_1598,In_1061);
nand U4223 (N_4223,In_592,In_1209);
nor U4224 (N_4224,In_2562,In_2458);
nor U4225 (N_4225,In_2595,In_1551);
xnor U4226 (N_4226,In_1890,In_2836);
xnor U4227 (N_4227,In_632,In_751);
xnor U4228 (N_4228,In_247,In_1793);
or U4229 (N_4229,In_845,In_2435);
nor U4230 (N_4230,In_2472,In_2587);
xnor U4231 (N_4231,In_8,In_1758);
nor U4232 (N_4232,In_391,In_1029);
and U4233 (N_4233,In_675,In_140);
xor U4234 (N_4234,In_2405,In_871);
nor U4235 (N_4235,In_2026,In_120);
and U4236 (N_4236,In_400,In_1131);
xnor U4237 (N_4237,In_1545,In_2967);
nand U4238 (N_4238,In_1235,In_406);
or U4239 (N_4239,In_1665,In_276);
xnor U4240 (N_4240,In_2258,In_2530);
and U4241 (N_4241,In_1102,In_1480);
nor U4242 (N_4242,In_1186,In_379);
nand U4243 (N_4243,In_1974,In_1655);
xor U4244 (N_4244,In_393,In_1660);
nand U4245 (N_4245,In_799,In_457);
nand U4246 (N_4246,In_1580,In_384);
and U4247 (N_4247,In_1037,In_2534);
xor U4248 (N_4248,In_2876,In_46);
and U4249 (N_4249,In_2872,In_701);
xor U4250 (N_4250,In_1483,In_999);
or U4251 (N_4251,In_1767,In_421);
or U4252 (N_4252,In_2939,In_210);
or U4253 (N_4253,In_458,In_2437);
and U4254 (N_4254,In_39,In_2574);
nor U4255 (N_4255,In_890,In_175);
nand U4256 (N_4256,In_1196,In_1175);
and U4257 (N_4257,In_2443,In_1009);
and U4258 (N_4258,In_685,In_944);
nor U4259 (N_4259,In_1498,In_1256);
or U4260 (N_4260,In_2478,In_1271);
xnor U4261 (N_4261,In_2818,In_2621);
or U4262 (N_4262,In_887,In_1391);
xnor U4263 (N_4263,In_2069,In_1865);
nand U4264 (N_4264,In_2283,In_242);
xor U4265 (N_4265,In_1434,In_1474);
nand U4266 (N_4266,In_396,In_619);
nand U4267 (N_4267,In_1283,In_222);
xor U4268 (N_4268,In_2712,In_2331);
nor U4269 (N_4269,In_1526,In_2574);
nand U4270 (N_4270,In_962,In_1661);
and U4271 (N_4271,In_1595,In_2799);
xor U4272 (N_4272,In_2041,In_130);
and U4273 (N_4273,In_303,In_376);
or U4274 (N_4274,In_1361,In_634);
or U4275 (N_4275,In_2523,In_418);
xor U4276 (N_4276,In_2684,In_157);
nand U4277 (N_4277,In_1672,In_1052);
or U4278 (N_4278,In_2921,In_512);
nor U4279 (N_4279,In_1076,In_55);
and U4280 (N_4280,In_1943,In_674);
or U4281 (N_4281,In_143,In_2749);
or U4282 (N_4282,In_133,In_1852);
nand U4283 (N_4283,In_542,In_357);
nor U4284 (N_4284,In_1962,In_543);
or U4285 (N_4285,In_2532,In_16);
xnor U4286 (N_4286,In_2899,In_670);
or U4287 (N_4287,In_2434,In_1482);
xnor U4288 (N_4288,In_748,In_2873);
xor U4289 (N_4289,In_2951,In_1222);
nand U4290 (N_4290,In_824,In_1681);
nand U4291 (N_4291,In_2714,In_1621);
or U4292 (N_4292,In_2033,In_667);
and U4293 (N_4293,In_2807,In_2190);
or U4294 (N_4294,In_374,In_1888);
and U4295 (N_4295,In_293,In_1247);
nand U4296 (N_4296,In_1840,In_57);
nand U4297 (N_4297,In_67,In_5);
or U4298 (N_4298,In_1904,In_2195);
nand U4299 (N_4299,In_1205,In_833);
xor U4300 (N_4300,In_237,In_1758);
and U4301 (N_4301,In_2614,In_286);
and U4302 (N_4302,In_1988,In_2548);
nand U4303 (N_4303,In_1470,In_2891);
nand U4304 (N_4304,In_240,In_1637);
and U4305 (N_4305,In_1422,In_1771);
and U4306 (N_4306,In_945,In_661);
nand U4307 (N_4307,In_893,In_1404);
or U4308 (N_4308,In_2847,In_150);
nor U4309 (N_4309,In_543,In_626);
xor U4310 (N_4310,In_499,In_111);
nor U4311 (N_4311,In_1051,In_215);
nor U4312 (N_4312,In_151,In_1397);
xnor U4313 (N_4313,In_1293,In_1995);
nand U4314 (N_4314,In_2781,In_2421);
and U4315 (N_4315,In_1046,In_417);
or U4316 (N_4316,In_2605,In_2786);
nor U4317 (N_4317,In_2430,In_79);
and U4318 (N_4318,In_470,In_1745);
xnor U4319 (N_4319,In_156,In_676);
and U4320 (N_4320,In_2315,In_2375);
or U4321 (N_4321,In_268,In_215);
and U4322 (N_4322,In_967,In_376);
and U4323 (N_4323,In_272,In_2373);
and U4324 (N_4324,In_1905,In_99);
nand U4325 (N_4325,In_2824,In_2541);
and U4326 (N_4326,In_926,In_776);
or U4327 (N_4327,In_226,In_2865);
or U4328 (N_4328,In_693,In_1367);
nor U4329 (N_4329,In_2253,In_1983);
nor U4330 (N_4330,In_720,In_320);
xnor U4331 (N_4331,In_1414,In_941);
nand U4332 (N_4332,In_287,In_1014);
xnor U4333 (N_4333,In_7,In_2716);
nand U4334 (N_4334,In_1456,In_2251);
nor U4335 (N_4335,In_891,In_2098);
nor U4336 (N_4336,In_1461,In_2966);
or U4337 (N_4337,In_1183,In_1156);
xor U4338 (N_4338,In_691,In_2500);
nand U4339 (N_4339,In_219,In_964);
nand U4340 (N_4340,In_712,In_1486);
and U4341 (N_4341,In_702,In_1474);
or U4342 (N_4342,In_1989,In_803);
xnor U4343 (N_4343,In_1428,In_1046);
nor U4344 (N_4344,In_2651,In_2831);
nand U4345 (N_4345,In_1181,In_2389);
and U4346 (N_4346,In_2774,In_284);
or U4347 (N_4347,In_2150,In_218);
nor U4348 (N_4348,In_1382,In_2957);
or U4349 (N_4349,In_550,In_361);
and U4350 (N_4350,In_2362,In_1367);
and U4351 (N_4351,In_2261,In_2902);
nand U4352 (N_4352,In_994,In_5);
and U4353 (N_4353,In_1590,In_784);
xor U4354 (N_4354,In_2600,In_839);
nor U4355 (N_4355,In_216,In_2463);
xnor U4356 (N_4356,In_192,In_1304);
nor U4357 (N_4357,In_1390,In_2272);
and U4358 (N_4358,In_1721,In_163);
xor U4359 (N_4359,In_2857,In_2999);
nand U4360 (N_4360,In_1804,In_610);
and U4361 (N_4361,In_1644,In_1371);
nor U4362 (N_4362,In_905,In_1615);
nand U4363 (N_4363,In_1821,In_650);
and U4364 (N_4364,In_857,In_1821);
nor U4365 (N_4365,In_2880,In_1180);
and U4366 (N_4366,In_487,In_2478);
nand U4367 (N_4367,In_1772,In_2319);
nor U4368 (N_4368,In_42,In_1934);
nor U4369 (N_4369,In_1229,In_1013);
or U4370 (N_4370,In_526,In_965);
or U4371 (N_4371,In_2169,In_1583);
and U4372 (N_4372,In_827,In_1647);
and U4373 (N_4373,In_1261,In_813);
and U4374 (N_4374,In_1362,In_2757);
xor U4375 (N_4375,In_2679,In_728);
xor U4376 (N_4376,In_1925,In_907);
and U4377 (N_4377,In_1121,In_950);
nor U4378 (N_4378,In_2241,In_2771);
xor U4379 (N_4379,In_224,In_1477);
xor U4380 (N_4380,In_2411,In_2530);
nor U4381 (N_4381,In_581,In_2744);
nand U4382 (N_4382,In_2914,In_989);
or U4383 (N_4383,In_2662,In_428);
and U4384 (N_4384,In_804,In_1160);
or U4385 (N_4385,In_640,In_2781);
or U4386 (N_4386,In_2358,In_317);
nand U4387 (N_4387,In_91,In_717);
nor U4388 (N_4388,In_2097,In_1323);
xnor U4389 (N_4389,In_1192,In_1913);
nor U4390 (N_4390,In_400,In_9);
xor U4391 (N_4391,In_1256,In_933);
xnor U4392 (N_4392,In_523,In_804);
nand U4393 (N_4393,In_2886,In_450);
xor U4394 (N_4394,In_2511,In_1245);
or U4395 (N_4395,In_1362,In_1165);
or U4396 (N_4396,In_1238,In_2805);
nor U4397 (N_4397,In_2560,In_1767);
or U4398 (N_4398,In_2431,In_2253);
xnor U4399 (N_4399,In_34,In_1031);
nand U4400 (N_4400,In_2439,In_2856);
xnor U4401 (N_4401,In_2886,In_2282);
nor U4402 (N_4402,In_1502,In_928);
and U4403 (N_4403,In_710,In_235);
and U4404 (N_4404,In_705,In_1349);
nand U4405 (N_4405,In_130,In_2649);
nor U4406 (N_4406,In_389,In_1625);
xor U4407 (N_4407,In_1218,In_2622);
nor U4408 (N_4408,In_1318,In_257);
and U4409 (N_4409,In_2470,In_1984);
xor U4410 (N_4410,In_2885,In_1068);
nand U4411 (N_4411,In_1340,In_218);
and U4412 (N_4412,In_70,In_228);
and U4413 (N_4413,In_1772,In_919);
xnor U4414 (N_4414,In_2847,In_1432);
or U4415 (N_4415,In_2622,In_2851);
xnor U4416 (N_4416,In_860,In_280);
and U4417 (N_4417,In_1125,In_369);
and U4418 (N_4418,In_710,In_1440);
or U4419 (N_4419,In_1328,In_1816);
xnor U4420 (N_4420,In_1869,In_1116);
or U4421 (N_4421,In_2248,In_384);
or U4422 (N_4422,In_365,In_190);
nor U4423 (N_4423,In_2094,In_2316);
or U4424 (N_4424,In_58,In_2250);
nand U4425 (N_4425,In_1365,In_2410);
or U4426 (N_4426,In_1750,In_1542);
and U4427 (N_4427,In_705,In_1291);
nor U4428 (N_4428,In_1284,In_2739);
and U4429 (N_4429,In_930,In_61);
xor U4430 (N_4430,In_623,In_1650);
nor U4431 (N_4431,In_1183,In_1194);
nor U4432 (N_4432,In_1211,In_2188);
and U4433 (N_4433,In_2791,In_1213);
xnor U4434 (N_4434,In_2446,In_341);
or U4435 (N_4435,In_1745,In_455);
or U4436 (N_4436,In_1514,In_2163);
and U4437 (N_4437,In_2100,In_1202);
and U4438 (N_4438,In_350,In_1555);
xor U4439 (N_4439,In_2069,In_1502);
xnor U4440 (N_4440,In_2153,In_1449);
xor U4441 (N_4441,In_1506,In_1805);
nor U4442 (N_4442,In_1377,In_1543);
nor U4443 (N_4443,In_119,In_2272);
nand U4444 (N_4444,In_1994,In_2975);
nand U4445 (N_4445,In_1169,In_1170);
or U4446 (N_4446,In_910,In_2079);
nand U4447 (N_4447,In_2539,In_750);
xnor U4448 (N_4448,In_1731,In_509);
or U4449 (N_4449,In_180,In_2140);
xor U4450 (N_4450,In_996,In_1076);
nor U4451 (N_4451,In_2080,In_1091);
nand U4452 (N_4452,In_1076,In_384);
nand U4453 (N_4453,In_119,In_1157);
and U4454 (N_4454,In_440,In_2067);
and U4455 (N_4455,In_1485,In_1883);
nor U4456 (N_4456,In_825,In_1483);
nand U4457 (N_4457,In_1032,In_760);
nor U4458 (N_4458,In_1300,In_2746);
nand U4459 (N_4459,In_209,In_2529);
nand U4460 (N_4460,In_1175,In_1199);
and U4461 (N_4461,In_1628,In_277);
nor U4462 (N_4462,In_2897,In_1466);
or U4463 (N_4463,In_1640,In_1390);
and U4464 (N_4464,In_1823,In_2739);
or U4465 (N_4465,In_859,In_1572);
and U4466 (N_4466,In_1473,In_2983);
nand U4467 (N_4467,In_2580,In_162);
and U4468 (N_4468,In_394,In_739);
and U4469 (N_4469,In_387,In_1408);
xnor U4470 (N_4470,In_2596,In_1006);
xnor U4471 (N_4471,In_1340,In_1391);
or U4472 (N_4472,In_2952,In_1829);
xnor U4473 (N_4473,In_451,In_1159);
xor U4474 (N_4474,In_1460,In_1875);
or U4475 (N_4475,In_349,In_2306);
nand U4476 (N_4476,In_2994,In_1637);
nor U4477 (N_4477,In_2105,In_1399);
xor U4478 (N_4478,In_1554,In_1998);
and U4479 (N_4479,In_2310,In_1685);
nor U4480 (N_4480,In_2328,In_2332);
and U4481 (N_4481,In_27,In_541);
xor U4482 (N_4482,In_1951,In_2333);
or U4483 (N_4483,In_2733,In_1544);
and U4484 (N_4484,In_1136,In_2057);
nor U4485 (N_4485,In_1965,In_2702);
xnor U4486 (N_4486,In_1316,In_1892);
xor U4487 (N_4487,In_496,In_300);
xnor U4488 (N_4488,In_1724,In_2887);
or U4489 (N_4489,In_2703,In_2817);
nor U4490 (N_4490,In_14,In_2428);
xnor U4491 (N_4491,In_1761,In_1352);
xor U4492 (N_4492,In_2903,In_181);
or U4493 (N_4493,In_2637,In_1740);
and U4494 (N_4494,In_2219,In_2034);
or U4495 (N_4495,In_520,In_624);
nor U4496 (N_4496,In_1031,In_2617);
nand U4497 (N_4497,In_194,In_131);
nor U4498 (N_4498,In_1600,In_2621);
xnor U4499 (N_4499,In_1709,In_2879);
and U4500 (N_4500,In_2725,In_654);
nor U4501 (N_4501,In_73,In_7);
nand U4502 (N_4502,In_1122,In_1371);
and U4503 (N_4503,In_1135,In_699);
and U4504 (N_4504,In_1814,In_2361);
and U4505 (N_4505,In_2466,In_904);
nor U4506 (N_4506,In_1646,In_2468);
nand U4507 (N_4507,In_2553,In_2562);
and U4508 (N_4508,In_457,In_2760);
or U4509 (N_4509,In_2238,In_2863);
xnor U4510 (N_4510,In_2430,In_1042);
xnor U4511 (N_4511,In_2758,In_2092);
nand U4512 (N_4512,In_2703,In_1004);
nand U4513 (N_4513,In_1349,In_1339);
nor U4514 (N_4514,In_584,In_2709);
nand U4515 (N_4515,In_522,In_1121);
nand U4516 (N_4516,In_780,In_1959);
xor U4517 (N_4517,In_2370,In_2876);
nor U4518 (N_4518,In_1616,In_234);
nor U4519 (N_4519,In_1493,In_308);
or U4520 (N_4520,In_2145,In_827);
nor U4521 (N_4521,In_738,In_1911);
nand U4522 (N_4522,In_184,In_1656);
and U4523 (N_4523,In_1181,In_1141);
and U4524 (N_4524,In_1242,In_1065);
or U4525 (N_4525,In_2281,In_1632);
or U4526 (N_4526,In_97,In_321);
and U4527 (N_4527,In_1126,In_2612);
and U4528 (N_4528,In_1006,In_2558);
or U4529 (N_4529,In_1739,In_2864);
nor U4530 (N_4530,In_1795,In_1488);
or U4531 (N_4531,In_302,In_1900);
or U4532 (N_4532,In_1734,In_2450);
nor U4533 (N_4533,In_2677,In_2273);
and U4534 (N_4534,In_2161,In_2831);
nand U4535 (N_4535,In_2369,In_173);
or U4536 (N_4536,In_1971,In_84);
and U4537 (N_4537,In_1185,In_109);
nand U4538 (N_4538,In_2689,In_1475);
and U4539 (N_4539,In_1878,In_758);
or U4540 (N_4540,In_1745,In_1713);
nor U4541 (N_4541,In_1881,In_811);
nand U4542 (N_4542,In_873,In_2383);
and U4543 (N_4543,In_2722,In_2552);
or U4544 (N_4544,In_2518,In_2079);
or U4545 (N_4545,In_2690,In_1463);
nor U4546 (N_4546,In_458,In_741);
nor U4547 (N_4547,In_1596,In_2410);
nand U4548 (N_4548,In_491,In_1791);
xnor U4549 (N_4549,In_2521,In_465);
nand U4550 (N_4550,In_1445,In_2374);
or U4551 (N_4551,In_1531,In_587);
or U4552 (N_4552,In_232,In_2051);
xor U4553 (N_4553,In_2905,In_1878);
or U4554 (N_4554,In_1488,In_393);
or U4555 (N_4555,In_825,In_554);
xor U4556 (N_4556,In_315,In_2784);
and U4557 (N_4557,In_1437,In_112);
nor U4558 (N_4558,In_245,In_2260);
and U4559 (N_4559,In_376,In_982);
and U4560 (N_4560,In_967,In_24);
nand U4561 (N_4561,In_1041,In_1423);
nand U4562 (N_4562,In_2152,In_154);
or U4563 (N_4563,In_617,In_2175);
xnor U4564 (N_4564,In_2113,In_1459);
nand U4565 (N_4565,In_1335,In_1307);
and U4566 (N_4566,In_1084,In_106);
nor U4567 (N_4567,In_2853,In_2577);
and U4568 (N_4568,In_2439,In_1920);
nor U4569 (N_4569,In_2858,In_314);
nand U4570 (N_4570,In_1921,In_833);
nand U4571 (N_4571,In_1452,In_401);
nand U4572 (N_4572,In_951,In_2188);
or U4573 (N_4573,In_1114,In_320);
nand U4574 (N_4574,In_1147,In_2317);
or U4575 (N_4575,In_2493,In_2204);
and U4576 (N_4576,In_1542,In_1197);
nor U4577 (N_4577,In_619,In_2054);
xnor U4578 (N_4578,In_695,In_748);
and U4579 (N_4579,In_1583,In_741);
and U4580 (N_4580,In_1843,In_1617);
nor U4581 (N_4581,In_2746,In_655);
and U4582 (N_4582,In_1114,In_1117);
and U4583 (N_4583,In_2920,In_398);
or U4584 (N_4584,In_2439,In_1182);
nand U4585 (N_4585,In_983,In_40);
nor U4586 (N_4586,In_475,In_642);
or U4587 (N_4587,In_1888,In_1029);
nand U4588 (N_4588,In_1541,In_1191);
and U4589 (N_4589,In_797,In_2900);
nand U4590 (N_4590,In_2162,In_2147);
or U4591 (N_4591,In_2877,In_532);
or U4592 (N_4592,In_1437,In_2401);
nand U4593 (N_4593,In_2481,In_1526);
nand U4594 (N_4594,In_1868,In_1228);
and U4595 (N_4595,In_2508,In_792);
xnor U4596 (N_4596,In_2516,In_2871);
xor U4597 (N_4597,In_1817,In_2364);
or U4598 (N_4598,In_147,In_44);
or U4599 (N_4599,In_2947,In_2675);
nand U4600 (N_4600,In_2569,In_1124);
nor U4601 (N_4601,In_212,In_294);
nand U4602 (N_4602,In_115,In_1549);
or U4603 (N_4603,In_2046,In_1553);
xor U4604 (N_4604,In_42,In_656);
or U4605 (N_4605,In_2494,In_1751);
xnor U4606 (N_4606,In_758,In_1747);
nand U4607 (N_4607,In_1618,In_2088);
xor U4608 (N_4608,In_2410,In_130);
nand U4609 (N_4609,In_1524,In_1993);
xor U4610 (N_4610,In_84,In_1160);
or U4611 (N_4611,In_898,In_700);
nand U4612 (N_4612,In_2639,In_1656);
or U4613 (N_4613,In_120,In_1951);
and U4614 (N_4614,In_988,In_479);
nor U4615 (N_4615,In_1076,In_521);
xnor U4616 (N_4616,In_236,In_336);
or U4617 (N_4617,In_1567,In_604);
and U4618 (N_4618,In_2765,In_1886);
and U4619 (N_4619,In_2290,In_1063);
or U4620 (N_4620,In_1087,In_2615);
xnor U4621 (N_4621,In_1622,In_2460);
xor U4622 (N_4622,In_2899,In_931);
nand U4623 (N_4623,In_1119,In_2621);
nor U4624 (N_4624,In_295,In_240);
or U4625 (N_4625,In_2990,In_1380);
xnor U4626 (N_4626,In_965,In_1523);
and U4627 (N_4627,In_953,In_1898);
and U4628 (N_4628,In_2282,In_1744);
or U4629 (N_4629,In_448,In_641);
nand U4630 (N_4630,In_2591,In_1102);
and U4631 (N_4631,In_54,In_1940);
and U4632 (N_4632,In_2248,In_2733);
nand U4633 (N_4633,In_152,In_1663);
xnor U4634 (N_4634,In_1826,In_1760);
nand U4635 (N_4635,In_2616,In_1743);
and U4636 (N_4636,In_2060,In_1312);
or U4637 (N_4637,In_1530,In_455);
and U4638 (N_4638,In_1467,In_1827);
and U4639 (N_4639,In_2143,In_2720);
nor U4640 (N_4640,In_2927,In_941);
or U4641 (N_4641,In_1332,In_1377);
and U4642 (N_4642,In_956,In_1637);
nor U4643 (N_4643,In_767,In_1662);
or U4644 (N_4644,In_1574,In_2961);
xnor U4645 (N_4645,In_2404,In_1318);
nand U4646 (N_4646,In_2689,In_1366);
nor U4647 (N_4647,In_838,In_202);
xnor U4648 (N_4648,In_1032,In_2422);
xnor U4649 (N_4649,In_688,In_254);
xor U4650 (N_4650,In_1428,In_1522);
and U4651 (N_4651,In_1388,In_1281);
nand U4652 (N_4652,In_1727,In_1406);
and U4653 (N_4653,In_2540,In_1790);
nor U4654 (N_4654,In_1028,In_2410);
nand U4655 (N_4655,In_355,In_2133);
nand U4656 (N_4656,In_914,In_1304);
nand U4657 (N_4657,In_791,In_2308);
nor U4658 (N_4658,In_1466,In_1602);
nand U4659 (N_4659,In_253,In_2817);
and U4660 (N_4660,In_1402,In_2765);
and U4661 (N_4661,In_2320,In_115);
nor U4662 (N_4662,In_1167,In_2988);
and U4663 (N_4663,In_610,In_680);
nand U4664 (N_4664,In_2446,In_2006);
nand U4665 (N_4665,In_881,In_2480);
and U4666 (N_4666,In_462,In_1175);
nand U4667 (N_4667,In_2252,In_1142);
or U4668 (N_4668,In_1594,In_1982);
and U4669 (N_4669,In_886,In_2778);
nand U4670 (N_4670,In_329,In_1410);
or U4671 (N_4671,In_1917,In_2129);
nand U4672 (N_4672,In_2105,In_2681);
xnor U4673 (N_4673,In_871,In_2173);
or U4674 (N_4674,In_2035,In_2443);
or U4675 (N_4675,In_2399,In_1399);
xnor U4676 (N_4676,In_431,In_2155);
and U4677 (N_4677,In_1061,In_2524);
nand U4678 (N_4678,In_172,In_2736);
or U4679 (N_4679,In_1331,In_1398);
xor U4680 (N_4680,In_2769,In_684);
nor U4681 (N_4681,In_2632,In_1156);
or U4682 (N_4682,In_298,In_2784);
xor U4683 (N_4683,In_338,In_921);
or U4684 (N_4684,In_1108,In_95);
nand U4685 (N_4685,In_99,In_541);
xor U4686 (N_4686,In_852,In_242);
or U4687 (N_4687,In_166,In_171);
nor U4688 (N_4688,In_2578,In_285);
or U4689 (N_4689,In_1130,In_1131);
nand U4690 (N_4690,In_1248,In_2146);
xor U4691 (N_4691,In_938,In_2503);
nor U4692 (N_4692,In_2561,In_1489);
nand U4693 (N_4693,In_2377,In_2904);
or U4694 (N_4694,In_2652,In_423);
and U4695 (N_4695,In_15,In_81);
nor U4696 (N_4696,In_741,In_1259);
nor U4697 (N_4697,In_1800,In_262);
nor U4698 (N_4698,In_598,In_902);
nor U4699 (N_4699,In_1083,In_894);
nand U4700 (N_4700,In_729,In_812);
xor U4701 (N_4701,In_2566,In_525);
and U4702 (N_4702,In_951,In_83);
xor U4703 (N_4703,In_1792,In_2111);
and U4704 (N_4704,In_1061,In_95);
xor U4705 (N_4705,In_2663,In_1795);
or U4706 (N_4706,In_903,In_1130);
and U4707 (N_4707,In_1806,In_1483);
or U4708 (N_4708,In_243,In_2856);
nand U4709 (N_4709,In_1990,In_2017);
or U4710 (N_4710,In_352,In_1679);
nor U4711 (N_4711,In_2728,In_2303);
or U4712 (N_4712,In_2064,In_2);
nor U4713 (N_4713,In_1059,In_2466);
xor U4714 (N_4714,In_284,In_2328);
xor U4715 (N_4715,In_2227,In_1137);
nor U4716 (N_4716,In_2732,In_2468);
nand U4717 (N_4717,In_831,In_2730);
nand U4718 (N_4718,In_1149,In_189);
or U4719 (N_4719,In_1566,In_2534);
or U4720 (N_4720,In_394,In_2197);
nor U4721 (N_4721,In_1395,In_2990);
or U4722 (N_4722,In_498,In_72);
and U4723 (N_4723,In_2762,In_2178);
nand U4724 (N_4724,In_228,In_2869);
nand U4725 (N_4725,In_219,In_913);
or U4726 (N_4726,In_151,In_2381);
xnor U4727 (N_4727,In_749,In_816);
or U4728 (N_4728,In_2383,In_208);
or U4729 (N_4729,In_669,In_508);
xor U4730 (N_4730,In_2015,In_1426);
and U4731 (N_4731,In_1741,In_305);
or U4732 (N_4732,In_1906,In_456);
xor U4733 (N_4733,In_2809,In_1861);
xnor U4734 (N_4734,In_2538,In_1644);
xor U4735 (N_4735,In_1057,In_2232);
nor U4736 (N_4736,In_2912,In_2973);
xor U4737 (N_4737,In_2794,In_2145);
or U4738 (N_4738,In_1685,In_1246);
xnor U4739 (N_4739,In_1735,In_443);
nor U4740 (N_4740,In_2167,In_2938);
xnor U4741 (N_4741,In_955,In_1766);
xor U4742 (N_4742,In_375,In_2732);
or U4743 (N_4743,In_1478,In_2178);
nand U4744 (N_4744,In_536,In_897);
and U4745 (N_4745,In_1622,In_1747);
and U4746 (N_4746,In_1290,In_613);
or U4747 (N_4747,In_345,In_1667);
nor U4748 (N_4748,In_1792,In_516);
nor U4749 (N_4749,In_1017,In_2962);
or U4750 (N_4750,In_54,In_1327);
xnor U4751 (N_4751,In_561,In_1732);
xor U4752 (N_4752,In_1698,In_1789);
xor U4753 (N_4753,In_2642,In_1628);
and U4754 (N_4754,In_101,In_1620);
xnor U4755 (N_4755,In_1528,In_550);
xor U4756 (N_4756,In_1091,In_1675);
nand U4757 (N_4757,In_242,In_2380);
nand U4758 (N_4758,In_305,In_2971);
nand U4759 (N_4759,In_1946,In_2335);
nor U4760 (N_4760,In_785,In_159);
or U4761 (N_4761,In_414,In_2284);
and U4762 (N_4762,In_335,In_2688);
and U4763 (N_4763,In_461,In_163);
or U4764 (N_4764,In_2242,In_822);
nor U4765 (N_4765,In_2948,In_2383);
nand U4766 (N_4766,In_2170,In_1301);
xnor U4767 (N_4767,In_1156,In_402);
and U4768 (N_4768,In_165,In_898);
xnor U4769 (N_4769,In_1179,In_2551);
nand U4770 (N_4770,In_785,In_2162);
and U4771 (N_4771,In_1315,In_2361);
and U4772 (N_4772,In_747,In_2247);
nand U4773 (N_4773,In_1774,In_2296);
nor U4774 (N_4774,In_2421,In_798);
nor U4775 (N_4775,In_555,In_2406);
nor U4776 (N_4776,In_151,In_497);
and U4777 (N_4777,In_355,In_2252);
and U4778 (N_4778,In_2042,In_1785);
or U4779 (N_4779,In_1475,In_2847);
nand U4780 (N_4780,In_1920,In_732);
and U4781 (N_4781,In_39,In_1984);
nor U4782 (N_4782,In_2224,In_1092);
nand U4783 (N_4783,In_903,In_2147);
xor U4784 (N_4784,In_1013,In_2077);
or U4785 (N_4785,In_180,In_2109);
or U4786 (N_4786,In_775,In_1808);
and U4787 (N_4787,In_911,In_1114);
nor U4788 (N_4788,In_424,In_2806);
and U4789 (N_4789,In_820,In_2933);
xnor U4790 (N_4790,In_630,In_1403);
and U4791 (N_4791,In_2488,In_1356);
or U4792 (N_4792,In_1811,In_1659);
xnor U4793 (N_4793,In_648,In_2397);
nand U4794 (N_4794,In_2146,In_962);
and U4795 (N_4795,In_844,In_1081);
nand U4796 (N_4796,In_1154,In_363);
nor U4797 (N_4797,In_6,In_33);
nor U4798 (N_4798,In_1318,In_1908);
nor U4799 (N_4799,In_1347,In_1932);
nor U4800 (N_4800,In_793,In_721);
and U4801 (N_4801,In_1590,In_2386);
nand U4802 (N_4802,In_461,In_1915);
nand U4803 (N_4803,In_2630,In_2287);
xor U4804 (N_4804,In_1297,In_1586);
or U4805 (N_4805,In_441,In_2915);
or U4806 (N_4806,In_2750,In_1555);
and U4807 (N_4807,In_1083,In_352);
nand U4808 (N_4808,In_1020,In_2271);
or U4809 (N_4809,In_1429,In_1828);
and U4810 (N_4810,In_2842,In_1435);
nor U4811 (N_4811,In_1465,In_1594);
nand U4812 (N_4812,In_396,In_1882);
and U4813 (N_4813,In_636,In_1909);
nor U4814 (N_4814,In_1309,In_1551);
xnor U4815 (N_4815,In_253,In_1783);
and U4816 (N_4816,In_2621,In_2832);
nand U4817 (N_4817,In_2644,In_389);
xor U4818 (N_4818,In_495,In_1118);
xnor U4819 (N_4819,In_2476,In_914);
xnor U4820 (N_4820,In_2890,In_1458);
xor U4821 (N_4821,In_742,In_515);
xor U4822 (N_4822,In_1459,In_2098);
nand U4823 (N_4823,In_2509,In_1174);
nor U4824 (N_4824,In_1538,In_2137);
xnor U4825 (N_4825,In_2019,In_1273);
or U4826 (N_4826,In_2256,In_2027);
nand U4827 (N_4827,In_2138,In_1018);
xor U4828 (N_4828,In_2593,In_2498);
nor U4829 (N_4829,In_1449,In_2092);
or U4830 (N_4830,In_2791,In_2993);
or U4831 (N_4831,In_1179,In_2275);
xor U4832 (N_4832,In_964,In_65);
and U4833 (N_4833,In_222,In_2586);
and U4834 (N_4834,In_1111,In_714);
and U4835 (N_4835,In_1851,In_2199);
nor U4836 (N_4836,In_2058,In_417);
nor U4837 (N_4837,In_2623,In_1001);
or U4838 (N_4838,In_2526,In_2238);
and U4839 (N_4839,In_377,In_1147);
or U4840 (N_4840,In_450,In_1059);
nand U4841 (N_4841,In_222,In_263);
xor U4842 (N_4842,In_279,In_2282);
nor U4843 (N_4843,In_341,In_999);
or U4844 (N_4844,In_2890,In_1446);
nand U4845 (N_4845,In_1398,In_1737);
and U4846 (N_4846,In_1246,In_2308);
xnor U4847 (N_4847,In_2289,In_2410);
and U4848 (N_4848,In_2136,In_2453);
xor U4849 (N_4849,In_893,In_1671);
and U4850 (N_4850,In_1736,In_2755);
or U4851 (N_4851,In_903,In_1114);
and U4852 (N_4852,In_1067,In_1974);
and U4853 (N_4853,In_144,In_2898);
or U4854 (N_4854,In_648,In_378);
or U4855 (N_4855,In_2161,In_2657);
nor U4856 (N_4856,In_1253,In_1958);
and U4857 (N_4857,In_536,In_1078);
nand U4858 (N_4858,In_863,In_1979);
or U4859 (N_4859,In_1564,In_2308);
xor U4860 (N_4860,In_2056,In_822);
nor U4861 (N_4861,In_2965,In_1411);
or U4862 (N_4862,In_808,In_1856);
nor U4863 (N_4863,In_1243,In_1208);
xor U4864 (N_4864,In_349,In_2631);
or U4865 (N_4865,In_98,In_1461);
xor U4866 (N_4866,In_2250,In_2957);
nor U4867 (N_4867,In_735,In_2732);
or U4868 (N_4868,In_1062,In_1827);
xnor U4869 (N_4869,In_967,In_539);
or U4870 (N_4870,In_2117,In_1029);
and U4871 (N_4871,In_1367,In_480);
or U4872 (N_4872,In_719,In_2212);
or U4873 (N_4873,In_2248,In_2786);
and U4874 (N_4874,In_2762,In_622);
xnor U4875 (N_4875,In_2824,In_716);
nor U4876 (N_4876,In_1635,In_377);
nor U4877 (N_4877,In_1451,In_57);
nand U4878 (N_4878,In_2148,In_2770);
xnor U4879 (N_4879,In_2826,In_264);
or U4880 (N_4880,In_1811,In_1398);
xnor U4881 (N_4881,In_2156,In_28);
nor U4882 (N_4882,In_2902,In_564);
nand U4883 (N_4883,In_2011,In_135);
and U4884 (N_4884,In_539,In_2531);
xnor U4885 (N_4885,In_162,In_1960);
or U4886 (N_4886,In_1189,In_29);
xor U4887 (N_4887,In_787,In_312);
or U4888 (N_4888,In_335,In_2325);
and U4889 (N_4889,In_2323,In_1718);
xnor U4890 (N_4890,In_277,In_2949);
nor U4891 (N_4891,In_1058,In_1411);
nor U4892 (N_4892,In_671,In_1727);
nor U4893 (N_4893,In_2908,In_1912);
xor U4894 (N_4894,In_631,In_2335);
and U4895 (N_4895,In_1791,In_2623);
xor U4896 (N_4896,In_1321,In_1403);
nand U4897 (N_4897,In_1389,In_2807);
xor U4898 (N_4898,In_2319,In_182);
nand U4899 (N_4899,In_928,In_2858);
or U4900 (N_4900,In_588,In_2825);
nor U4901 (N_4901,In_1680,In_169);
or U4902 (N_4902,In_156,In_2802);
xnor U4903 (N_4903,In_1585,In_2582);
or U4904 (N_4904,In_1898,In_2831);
nand U4905 (N_4905,In_1405,In_454);
nand U4906 (N_4906,In_2016,In_735);
nand U4907 (N_4907,In_2458,In_2090);
xor U4908 (N_4908,In_869,In_2492);
nand U4909 (N_4909,In_2251,In_1469);
and U4910 (N_4910,In_2562,In_1034);
or U4911 (N_4911,In_1997,In_2042);
xor U4912 (N_4912,In_2291,In_1305);
and U4913 (N_4913,In_1477,In_2550);
xnor U4914 (N_4914,In_1122,In_286);
and U4915 (N_4915,In_1641,In_1445);
xnor U4916 (N_4916,In_1001,In_1884);
or U4917 (N_4917,In_2154,In_2079);
xor U4918 (N_4918,In_776,In_92);
nor U4919 (N_4919,In_2880,In_808);
nand U4920 (N_4920,In_941,In_771);
or U4921 (N_4921,In_947,In_690);
xnor U4922 (N_4922,In_1868,In_2816);
and U4923 (N_4923,In_1529,In_1438);
nand U4924 (N_4924,In_56,In_1910);
nand U4925 (N_4925,In_1361,In_1294);
or U4926 (N_4926,In_2512,In_841);
xor U4927 (N_4927,In_1405,In_2255);
nand U4928 (N_4928,In_2380,In_1653);
and U4929 (N_4929,In_1330,In_2144);
nor U4930 (N_4930,In_589,In_1542);
and U4931 (N_4931,In_1478,In_450);
xnor U4932 (N_4932,In_627,In_1531);
nor U4933 (N_4933,In_306,In_1162);
or U4934 (N_4934,In_2069,In_389);
nor U4935 (N_4935,In_1031,In_1900);
and U4936 (N_4936,In_1215,In_1781);
nand U4937 (N_4937,In_1659,In_1082);
nor U4938 (N_4938,In_2737,In_715);
nor U4939 (N_4939,In_822,In_2530);
nand U4940 (N_4940,In_2811,In_2582);
nor U4941 (N_4941,In_367,In_955);
nor U4942 (N_4942,In_2126,In_2758);
nand U4943 (N_4943,In_1044,In_1175);
nand U4944 (N_4944,In_657,In_1631);
nand U4945 (N_4945,In_1560,In_1343);
xnor U4946 (N_4946,In_1577,In_504);
xor U4947 (N_4947,In_395,In_545);
or U4948 (N_4948,In_1920,In_495);
and U4949 (N_4949,In_196,In_2872);
and U4950 (N_4950,In_1470,In_589);
xnor U4951 (N_4951,In_1866,In_686);
or U4952 (N_4952,In_1491,In_1058);
nand U4953 (N_4953,In_2578,In_2374);
and U4954 (N_4954,In_778,In_2937);
nand U4955 (N_4955,In_379,In_734);
nor U4956 (N_4956,In_2429,In_1943);
nand U4957 (N_4957,In_2498,In_1701);
or U4958 (N_4958,In_2514,In_1860);
xor U4959 (N_4959,In_2510,In_1578);
nor U4960 (N_4960,In_1521,In_2252);
xnor U4961 (N_4961,In_2110,In_2635);
nand U4962 (N_4962,In_2247,In_2959);
xor U4963 (N_4963,In_1658,In_1390);
or U4964 (N_4964,In_1626,In_1407);
and U4965 (N_4965,In_2319,In_2059);
nand U4966 (N_4966,In_54,In_1023);
or U4967 (N_4967,In_2219,In_2811);
or U4968 (N_4968,In_2732,In_2951);
xnor U4969 (N_4969,In_420,In_2068);
and U4970 (N_4970,In_10,In_1936);
or U4971 (N_4971,In_713,In_582);
or U4972 (N_4972,In_1222,In_2798);
xor U4973 (N_4973,In_2145,In_2878);
xnor U4974 (N_4974,In_1565,In_1571);
nor U4975 (N_4975,In_1316,In_211);
nor U4976 (N_4976,In_1540,In_2671);
xnor U4977 (N_4977,In_1947,In_1342);
xor U4978 (N_4978,In_538,In_2226);
or U4979 (N_4979,In_2981,In_998);
or U4980 (N_4980,In_2197,In_2010);
or U4981 (N_4981,In_2522,In_2447);
xor U4982 (N_4982,In_2561,In_1584);
xor U4983 (N_4983,In_443,In_982);
or U4984 (N_4984,In_2820,In_2690);
and U4985 (N_4985,In_2500,In_16);
nand U4986 (N_4986,In_107,In_1381);
or U4987 (N_4987,In_2268,In_503);
or U4988 (N_4988,In_410,In_689);
xnor U4989 (N_4989,In_1122,In_2551);
and U4990 (N_4990,In_2091,In_2196);
or U4991 (N_4991,In_1743,In_586);
xor U4992 (N_4992,In_715,In_2955);
or U4993 (N_4993,In_1140,In_2075);
xor U4994 (N_4994,In_2309,In_899);
nand U4995 (N_4995,In_996,In_2225);
and U4996 (N_4996,In_2684,In_1863);
xnor U4997 (N_4997,In_500,In_637);
nor U4998 (N_4998,In_822,In_275);
xnor U4999 (N_4999,In_2812,In_1723);
xor U5000 (N_5000,N_1401,N_4998);
nor U5001 (N_5001,N_826,N_4314);
or U5002 (N_5002,N_2904,N_302);
xor U5003 (N_5003,N_4458,N_2130);
nand U5004 (N_5004,N_625,N_1289);
or U5005 (N_5005,N_4124,N_3369);
and U5006 (N_5006,N_3930,N_2282);
and U5007 (N_5007,N_3036,N_4944);
and U5008 (N_5008,N_3512,N_1492);
xor U5009 (N_5009,N_1516,N_3042);
and U5010 (N_5010,N_3406,N_1660);
and U5011 (N_5011,N_2422,N_1298);
or U5012 (N_5012,N_92,N_1274);
or U5013 (N_5013,N_4699,N_2240);
nor U5014 (N_5014,N_845,N_1471);
nand U5015 (N_5015,N_3198,N_3920);
nand U5016 (N_5016,N_1390,N_3854);
and U5017 (N_5017,N_878,N_291);
nor U5018 (N_5018,N_4920,N_4993);
nor U5019 (N_5019,N_2480,N_1669);
nor U5020 (N_5020,N_1322,N_2857);
xor U5021 (N_5021,N_2464,N_333);
nor U5022 (N_5022,N_1002,N_4760);
and U5023 (N_5023,N_4239,N_2592);
or U5024 (N_5024,N_3657,N_4295);
or U5025 (N_5025,N_4764,N_19);
nor U5026 (N_5026,N_4834,N_2897);
and U5027 (N_5027,N_142,N_3517);
xnor U5028 (N_5028,N_2060,N_3342);
and U5029 (N_5029,N_1070,N_1798);
nor U5030 (N_5030,N_1803,N_1490);
or U5031 (N_5031,N_3394,N_3646);
nor U5032 (N_5032,N_3858,N_236);
or U5033 (N_5033,N_4700,N_1383);
nor U5034 (N_5034,N_4554,N_4604);
and U5035 (N_5035,N_2767,N_155);
nor U5036 (N_5036,N_4877,N_400);
xnor U5037 (N_5037,N_3054,N_321);
xnor U5038 (N_5038,N_4070,N_4446);
and U5039 (N_5039,N_2334,N_2917);
nand U5040 (N_5040,N_1578,N_935);
xnor U5041 (N_5041,N_860,N_2074);
nor U5042 (N_5042,N_1221,N_2026);
and U5043 (N_5043,N_732,N_186);
nor U5044 (N_5044,N_4532,N_4394);
nor U5045 (N_5045,N_3612,N_4845);
and U5046 (N_5046,N_4423,N_4876);
xnor U5047 (N_5047,N_1863,N_366);
nor U5048 (N_5048,N_112,N_4254);
and U5049 (N_5049,N_4456,N_1139);
and U5050 (N_5050,N_4260,N_825);
nor U5051 (N_5051,N_3067,N_4478);
nor U5052 (N_5052,N_1642,N_3549);
nand U5053 (N_5053,N_497,N_235);
or U5054 (N_5054,N_4015,N_990);
xor U5055 (N_5055,N_2698,N_4242);
or U5056 (N_5056,N_4636,N_829);
nand U5057 (N_5057,N_3941,N_328);
nor U5058 (N_5058,N_1657,N_4722);
xor U5059 (N_5059,N_2736,N_1891);
nand U5060 (N_5060,N_3360,N_3960);
nor U5061 (N_5061,N_311,N_2233);
and U5062 (N_5062,N_4237,N_1852);
and U5063 (N_5063,N_3053,N_871);
and U5064 (N_5064,N_13,N_307);
and U5065 (N_5065,N_481,N_74);
and U5066 (N_5066,N_1150,N_4795);
and U5067 (N_5067,N_1443,N_1498);
and U5068 (N_5068,N_2291,N_4529);
and U5069 (N_5069,N_4880,N_618);
nand U5070 (N_5070,N_2387,N_853);
nand U5071 (N_5071,N_2571,N_863);
xnor U5072 (N_5072,N_2088,N_4819);
nor U5073 (N_5073,N_2192,N_2431);
and U5074 (N_5074,N_538,N_3939);
nor U5075 (N_5075,N_554,N_2093);
xnor U5076 (N_5076,N_3983,N_2327);
nor U5077 (N_5077,N_4471,N_4563);
xor U5078 (N_5078,N_940,N_2153);
nand U5079 (N_5079,N_3090,N_694);
xnor U5080 (N_5080,N_2593,N_2944);
nor U5081 (N_5081,N_3463,N_4008);
or U5082 (N_5082,N_573,N_2568);
nor U5083 (N_5083,N_4747,N_2353);
nor U5084 (N_5084,N_3702,N_2475);
or U5085 (N_5085,N_4249,N_2670);
nand U5086 (N_5086,N_4621,N_4995);
nand U5087 (N_5087,N_458,N_815);
xor U5088 (N_5088,N_1271,N_2655);
nor U5089 (N_5089,N_3382,N_4550);
xnor U5090 (N_5090,N_2034,N_1215);
xor U5091 (N_5091,N_474,N_4957);
and U5092 (N_5092,N_3759,N_1908);
xor U5093 (N_5093,N_313,N_2357);
nor U5094 (N_5094,N_3353,N_2631);
and U5095 (N_5095,N_2530,N_2288);
nand U5096 (N_5096,N_3482,N_3004);
and U5097 (N_5097,N_3459,N_537);
or U5098 (N_5098,N_763,N_1413);
and U5099 (N_5099,N_2172,N_3308);
nand U5100 (N_5100,N_94,N_1685);
and U5101 (N_5101,N_4964,N_957);
nand U5102 (N_5102,N_4972,N_396);
nor U5103 (N_5103,N_4858,N_2924);
nand U5104 (N_5104,N_375,N_373);
nand U5105 (N_5105,N_4727,N_643);
nand U5106 (N_5106,N_1086,N_2636);
or U5107 (N_5107,N_3486,N_4890);
nand U5108 (N_5108,N_2190,N_1698);
xor U5109 (N_5109,N_3423,N_4041);
nand U5110 (N_5110,N_3837,N_3079);
or U5111 (N_5111,N_3431,N_1427);
and U5112 (N_5112,N_46,N_240);
nand U5113 (N_5113,N_4047,N_2829);
nor U5114 (N_5114,N_1889,N_819);
xor U5115 (N_5115,N_591,N_4064);
nand U5116 (N_5116,N_250,N_1946);
or U5117 (N_5117,N_2094,N_475);
xor U5118 (N_5118,N_3648,N_2117);
nand U5119 (N_5119,N_3921,N_2833);
nor U5120 (N_5120,N_3900,N_3650);
or U5121 (N_5121,N_2788,N_3598);
nor U5122 (N_5122,N_2004,N_2125);
nor U5123 (N_5123,N_3516,N_4734);
xor U5124 (N_5124,N_294,N_1209);
xnor U5125 (N_5125,N_2477,N_3021);
and U5126 (N_5126,N_524,N_2906);
nand U5127 (N_5127,N_4870,N_663);
and U5128 (N_5128,N_4716,N_424);
nand U5129 (N_5129,N_2802,N_3807);
or U5130 (N_5130,N_1522,N_1104);
and U5131 (N_5131,N_3851,N_2169);
or U5132 (N_5132,N_2341,N_203);
nand U5133 (N_5133,N_551,N_858);
nor U5134 (N_5134,N_2145,N_2392);
and U5135 (N_5135,N_1124,N_2438);
nor U5136 (N_5136,N_1069,N_2359);
nand U5137 (N_5137,N_2209,N_3962);
nand U5138 (N_5138,N_3870,N_4552);
xor U5139 (N_5139,N_3362,N_3754);
or U5140 (N_5140,N_4414,N_3562);
or U5141 (N_5141,N_2067,N_2517);
or U5142 (N_5142,N_3465,N_4489);
and U5143 (N_5143,N_4386,N_4322);
xor U5144 (N_5144,N_4472,N_1621);
xor U5145 (N_5145,N_1109,N_1297);
xor U5146 (N_5146,N_2007,N_4987);
or U5147 (N_5147,N_4925,N_2379);
xnor U5148 (N_5148,N_2985,N_4428);
and U5149 (N_5149,N_2030,N_2828);
nand U5150 (N_5150,N_1461,N_331);
or U5151 (N_5151,N_4167,N_547);
or U5152 (N_5152,N_3952,N_4939);
xor U5153 (N_5153,N_1268,N_4777);
nand U5154 (N_5154,N_4039,N_803);
xnor U5155 (N_5155,N_3306,N_1965);
xor U5156 (N_5156,N_4686,N_3554);
nand U5157 (N_5157,N_2051,N_429);
or U5158 (N_5158,N_3520,N_4588);
and U5159 (N_5159,N_2160,N_4931);
nor U5160 (N_5160,N_1746,N_2149);
or U5161 (N_5161,N_965,N_4492);
xnor U5162 (N_5162,N_2785,N_371);
nand U5163 (N_5163,N_2968,N_3985);
nor U5164 (N_5164,N_2812,N_1005);
xnor U5165 (N_5165,N_427,N_3893);
xnor U5166 (N_5166,N_1904,N_1003);
or U5167 (N_5167,N_3092,N_1821);
or U5168 (N_5168,N_2402,N_2086);
nand U5169 (N_5169,N_4664,N_3584);
nand U5170 (N_5170,N_1447,N_692);
and U5171 (N_5171,N_987,N_2586);
nand U5172 (N_5172,N_1098,N_281);
xor U5173 (N_5173,N_939,N_1906);
or U5174 (N_5174,N_1633,N_4671);
and U5175 (N_5175,N_639,N_387);
nand U5176 (N_5176,N_2346,N_3157);
or U5177 (N_5177,N_1396,N_696);
nand U5178 (N_5178,N_2385,N_3064);
xnor U5179 (N_5179,N_2869,N_1812);
nor U5180 (N_5180,N_4932,N_3179);
nor U5181 (N_5181,N_3386,N_4882);
nand U5182 (N_5182,N_964,N_1778);
nand U5183 (N_5183,N_992,N_4348);
nand U5184 (N_5184,N_757,N_504);
and U5185 (N_5185,N_1591,N_39);
and U5186 (N_5186,N_2619,N_2782);
or U5187 (N_5187,N_4329,N_3329);
and U5188 (N_5188,N_4036,N_946);
nand U5189 (N_5189,N_4682,N_943);
nor U5190 (N_5190,N_1974,N_640);
nand U5191 (N_5191,N_2315,N_4754);
and U5192 (N_5192,N_3785,N_4571);
xor U5193 (N_5193,N_391,N_2537);
nor U5194 (N_5194,N_4048,N_509);
xor U5195 (N_5195,N_2338,N_336);
nor U5196 (N_5196,N_4004,N_469);
or U5197 (N_5197,N_1488,N_1800);
nor U5198 (N_5198,N_1795,N_386);
nor U5199 (N_5199,N_4137,N_3180);
or U5200 (N_5200,N_1476,N_3168);
nand U5201 (N_5201,N_3031,N_4000);
nor U5202 (N_5202,N_3300,N_3999);
and U5203 (N_5203,N_329,N_4017);
or U5204 (N_5204,N_1329,N_367);
xnor U5205 (N_5205,N_1761,N_1638);
and U5206 (N_5206,N_4152,N_2069);
or U5207 (N_5207,N_3736,N_3048);
and U5208 (N_5208,N_4518,N_3847);
xor U5209 (N_5209,N_4328,N_1049);
nand U5210 (N_5210,N_1239,N_2099);
nor U5211 (N_5211,N_4283,N_3396);
or U5212 (N_5212,N_4705,N_4991);
xor U5213 (N_5213,N_4191,N_178);
or U5214 (N_5214,N_141,N_2747);
and U5215 (N_5215,N_3832,N_1814);
or U5216 (N_5216,N_4038,N_1593);
or U5217 (N_5217,N_1682,N_3816);
nand U5218 (N_5218,N_3532,N_4079);
nand U5219 (N_5219,N_471,N_744);
nand U5220 (N_5220,N_108,N_1900);
and U5221 (N_5221,N_192,N_2707);
xnor U5222 (N_5222,N_2333,N_4466);
or U5223 (N_5223,N_1464,N_2428);
nor U5224 (N_5224,N_1818,N_1115);
nand U5225 (N_5225,N_1910,N_2432);
and U5226 (N_5226,N_2588,N_64);
and U5227 (N_5227,N_928,N_4633);
nand U5228 (N_5228,N_593,N_4872);
nor U5229 (N_5229,N_699,N_796);
nand U5230 (N_5230,N_2276,N_4339);
and U5231 (N_5231,N_365,N_2755);
nand U5232 (N_5232,N_4483,N_3641);
nor U5233 (N_5233,N_3364,N_90);
xnor U5234 (N_5234,N_3522,N_1075);
nor U5235 (N_5235,N_3901,N_4797);
nand U5236 (N_5236,N_2625,N_4127);
and U5237 (N_5237,N_2349,N_1792);
or U5238 (N_5238,N_65,N_2495);
or U5239 (N_5239,N_3447,N_4413);
nor U5240 (N_5240,N_298,N_4303);
xor U5241 (N_5241,N_569,N_4580);
nor U5242 (N_5242,N_434,N_3393);
nor U5243 (N_5243,N_4334,N_2649);
xnor U5244 (N_5244,N_4353,N_1984);
or U5245 (N_5245,N_2515,N_886);
or U5246 (N_5246,N_3005,N_2876);
nor U5247 (N_5247,N_4293,N_2621);
xor U5248 (N_5248,N_2470,N_1035);
nand U5249 (N_5249,N_4647,N_283);
xnor U5250 (N_5250,N_4337,N_1467);
nand U5251 (N_5251,N_4893,N_3931);
xor U5252 (N_5252,N_2957,N_4468);
xor U5253 (N_5253,N_659,N_3487);
nor U5254 (N_5254,N_4990,N_1376);
xnor U5255 (N_5255,N_4556,N_3194);
xor U5256 (N_5256,N_4406,N_1280);
xor U5257 (N_5257,N_405,N_648);
or U5258 (N_5258,N_1809,N_4172);
nand U5259 (N_5259,N_1892,N_4397);
nand U5260 (N_5260,N_1112,N_2771);
nor U5261 (N_5261,N_4775,N_3170);
or U5262 (N_5262,N_3305,N_2436);
and U5263 (N_5263,N_4591,N_4440);
or U5264 (N_5264,N_4356,N_1072);
nand U5265 (N_5265,N_2865,N_2448);
and U5266 (N_5266,N_4497,N_3122);
nor U5267 (N_5267,N_4698,N_2966);
nor U5268 (N_5268,N_4097,N_3683);
nor U5269 (N_5269,N_2692,N_3221);
or U5270 (N_5270,N_2182,N_285);
or U5271 (N_5271,N_702,N_4573);
and U5272 (N_5272,N_50,N_808);
nor U5273 (N_5273,N_1597,N_559);
xnor U5274 (N_5274,N_635,N_3793);
nor U5275 (N_5275,N_1225,N_1439);
or U5276 (N_5276,N_827,N_3343);
or U5277 (N_5277,N_2560,N_2245);
nor U5278 (N_5278,N_3859,N_3006);
or U5279 (N_5279,N_4966,N_2573);
xor U5280 (N_5280,N_4728,N_288);
nand U5281 (N_5281,N_1008,N_1941);
and U5282 (N_5282,N_2241,N_3615);
and U5283 (N_5283,N_3917,N_185);
or U5284 (N_5284,N_2010,N_3104);
or U5285 (N_5285,N_2710,N_4275);
and U5286 (N_5286,N_3226,N_2599);
and U5287 (N_5287,N_929,N_2708);
nor U5288 (N_5288,N_1631,N_4016);
nand U5289 (N_5289,N_29,N_1874);
or U5290 (N_5290,N_806,N_954);
and U5291 (N_5291,N_2919,N_2734);
nand U5292 (N_5292,N_3632,N_4973);
xor U5293 (N_5293,N_4520,N_2330);
nand U5294 (N_5294,N_1056,N_440);
and U5295 (N_5295,N_3440,N_3223);
or U5296 (N_5296,N_2574,N_4619);
or U5297 (N_5297,N_2668,N_125);
or U5298 (N_5298,N_3315,N_3553);
nand U5299 (N_5299,N_2119,N_444);
or U5300 (N_5300,N_2453,N_2055);
nand U5301 (N_5301,N_4197,N_3032);
xnor U5302 (N_5302,N_4343,N_1202);
and U5303 (N_5303,N_1048,N_4557);
and U5304 (N_5304,N_4480,N_4342);
and U5305 (N_5305,N_2723,N_2971);
nor U5306 (N_5306,N_491,N_1846);
and U5307 (N_5307,N_2663,N_4945);
nand U5308 (N_5308,N_1006,N_1480);
nor U5309 (N_5309,N_2285,N_4);
nand U5310 (N_5310,N_2711,N_1875);
nor U5311 (N_5311,N_3167,N_4702);
and U5312 (N_5312,N_1304,N_4357);
nand U5313 (N_5313,N_4188,N_3942);
xnor U5314 (N_5314,N_1102,N_1200);
and U5315 (N_5315,N_2694,N_2725);
nor U5316 (N_5316,N_1884,N_3768);
and U5317 (N_5317,N_42,N_4838);
and U5318 (N_5318,N_2909,N_4474);
and U5319 (N_5319,N_1911,N_3703);
or U5320 (N_5320,N_3762,N_2926);
or U5321 (N_5321,N_4364,N_2665);
or U5322 (N_5322,N_3594,N_54);
nor U5323 (N_5323,N_3891,N_3550);
and U5324 (N_5324,N_3746,N_1106);
nand U5325 (N_5325,N_4380,N_3622);
nor U5326 (N_5326,N_996,N_270);
and U5327 (N_5327,N_4831,N_2974);
and U5328 (N_5328,N_2916,N_613);
and U5329 (N_5329,N_87,N_3506);
nor U5330 (N_5330,N_79,N_4323);
or U5331 (N_5331,N_1815,N_4156);
nand U5332 (N_5332,N_3923,N_337);
or U5333 (N_5333,N_2684,N_588);
nand U5334 (N_5334,N_655,N_78);
xnor U5335 (N_5335,N_3298,N_4222);
or U5336 (N_5336,N_3260,N_1615);
or U5337 (N_5337,N_4436,N_1773);
or U5338 (N_5338,N_3016,N_2662);
or U5339 (N_5339,N_969,N_1090);
or U5340 (N_5340,N_2270,N_3576);
nand U5341 (N_5341,N_1136,N_1001);
xnor U5342 (N_5342,N_4219,N_2351);
nor U5343 (N_5343,N_1777,N_196);
nor U5344 (N_5344,N_1142,N_4154);
or U5345 (N_5345,N_342,N_1402);
xnor U5346 (N_5346,N_4128,N_582);
nor U5347 (N_5347,N_2607,N_565);
nand U5348 (N_5348,N_2445,N_604);
and U5349 (N_5349,N_1211,N_2577);
or U5350 (N_5350,N_3402,N_4926);
or U5351 (N_5351,N_1170,N_2693);
nor U5352 (N_5352,N_4980,N_4684);
nand U5353 (N_5353,N_1629,N_4543);
and U5354 (N_5354,N_2195,N_731);
or U5355 (N_5355,N_2413,N_2439);
xnor U5356 (N_5356,N_363,N_1757);
xnor U5357 (N_5357,N_3137,N_1559);
xor U5358 (N_5358,N_4799,N_4692);
xor U5359 (N_5359,N_2491,N_892);
nand U5360 (N_5360,N_1061,N_652);
nand U5361 (N_5361,N_1405,N_4642);
nor U5362 (N_5362,N_1585,N_900);
nor U5363 (N_5363,N_4798,N_798);
nor U5364 (N_5364,N_1720,N_3907);
nor U5365 (N_5365,N_70,N_718);
nand U5366 (N_5366,N_2699,N_2637);
nor U5367 (N_5367,N_1357,N_1607);
or U5368 (N_5368,N_3581,N_1704);
and U5369 (N_5369,N_4791,N_4788);
nand U5370 (N_5370,N_693,N_1080);
nand U5371 (N_5371,N_37,N_2307);
nand U5372 (N_5372,N_1716,N_3264);
nand U5373 (N_5373,N_1713,N_77);
or U5374 (N_5374,N_72,N_3103);
or U5375 (N_5375,N_890,N_2215);
and U5376 (N_5376,N_3346,N_3833);
and U5377 (N_5377,N_1347,N_2123);
or U5378 (N_5378,N_595,N_1625);
or U5379 (N_5379,N_1616,N_1389);
nand U5380 (N_5380,N_2814,N_4246);
xor U5381 (N_5381,N_608,N_4919);
nand U5382 (N_5382,N_113,N_1921);
nor U5383 (N_5383,N_3685,N_4978);
nor U5384 (N_5384,N_4632,N_3593);
nand U5385 (N_5385,N_952,N_3670);
nor U5386 (N_5386,N_2446,N_4068);
and U5387 (N_5387,N_4052,N_3799);
or U5388 (N_5388,N_1861,N_1101);
or U5389 (N_5389,N_2612,N_2221);
nand U5390 (N_5390,N_4132,N_1132);
nand U5391 (N_5391,N_418,N_2035);
nor U5392 (N_5392,N_2513,N_1417);
xnor U5393 (N_5393,N_465,N_1886);
and U5394 (N_5394,N_466,N_207);
nor U5395 (N_5395,N_678,N_3937);
nor U5396 (N_5396,N_3184,N_3496);
nand U5397 (N_5397,N_2648,N_1753);
or U5398 (N_5398,N_167,N_525);
nor U5399 (N_5399,N_4617,N_3959);
and U5400 (N_5400,N_907,N_1866);
and U5401 (N_5401,N_3716,N_1934);
nor U5402 (N_5402,N_1572,N_1764);
or U5403 (N_5403,N_310,N_3780);
nand U5404 (N_5404,N_1515,N_4538);
or U5405 (N_5405,N_1362,N_4950);
xor U5406 (N_5406,N_1917,N_2680);
or U5407 (N_5407,N_4594,N_1549);
or U5408 (N_5408,N_3708,N_4826);
nand U5409 (N_5409,N_2984,N_238);
or U5410 (N_5410,N_1703,N_4104);
xor U5411 (N_5411,N_3233,N_144);
and U5412 (N_5412,N_3915,N_3741);
nor U5413 (N_5413,N_308,N_1025);
nand U5414 (N_5414,N_1084,N_2382);
nor U5415 (N_5415,N_1611,N_2766);
nand U5416 (N_5416,N_2242,N_380);
xnor U5417 (N_5417,N_3250,N_423);
nor U5418 (N_5418,N_4326,N_1656);
or U5419 (N_5419,N_1442,N_1395);
xor U5420 (N_5420,N_1228,N_3188);
or U5421 (N_5421,N_3230,N_980);
and U5422 (N_5422,N_2959,N_406);
nor U5423 (N_5423,N_2809,N_847);
or U5424 (N_5424,N_1979,N_1734);
or U5425 (N_5425,N_2146,N_179);
or U5426 (N_5426,N_2675,N_2765);
nand U5427 (N_5427,N_3357,N_4042);
xor U5428 (N_5428,N_3081,N_2690);
nor U5429 (N_5429,N_895,N_1010);
nand U5430 (N_5430,N_2572,N_1269);
and U5431 (N_5431,N_2014,N_1530);
or U5432 (N_5432,N_2548,N_4315);
and U5433 (N_5433,N_4994,N_1975);
or U5434 (N_5434,N_2360,N_4895);
and U5435 (N_5435,N_4110,N_1301);
nand U5436 (N_5436,N_482,N_2481);
or U5437 (N_5437,N_4861,N_495);
nand U5438 (N_5438,N_2556,N_975);
nor U5439 (N_5439,N_2462,N_2009);
and U5440 (N_5440,N_2133,N_1896);
or U5441 (N_5441,N_4680,N_528);
or U5442 (N_5442,N_4714,N_1368);
xnor U5443 (N_5443,N_356,N_3257);
or U5444 (N_5444,N_1775,N_3153);
xnor U5445 (N_5445,N_403,N_2310);
nand U5446 (N_5446,N_4886,N_2264);
and U5447 (N_5447,N_2908,N_426);
or U5448 (N_5448,N_2664,N_917);
xnor U5449 (N_5449,N_268,N_4400);
nand U5450 (N_5450,N_4765,N_2156);
nor U5451 (N_5451,N_884,N_3424);
nor U5452 (N_5452,N_4013,N_1054);
nor U5453 (N_5453,N_2188,N_2033);
and U5454 (N_5454,N_289,N_1730);
or U5455 (N_5455,N_1945,N_3609);
and U5456 (N_5456,N_1365,N_4613);
and U5457 (N_5457,N_3659,N_3152);
nand U5458 (N_5458,N_1253,N_1412);
nand U5459 (N_5459,N_1248,N_4007);
or U5460 (N_5460,N_736,N_4860);
and U5461 (N_5461,N_4969,N_161);
and U5462 (N_5462,N_4731,N_3126);
xor U5463 (N_5463,N_3484,N_850);
nor U5464 (N_5464,N_489,N_2293);
and U5465 (N_5465,N_4245,N_4928);
or U5466 (N_5466,N_3753,N_4215);
or U5467 (N_5467,N_3478,N_4953);
or U5468 (N_5468,N_3892,N_412);
nand U5469 (N_5469,N_4997,N_4310);
and U5470 (N_5470,N_256,N_1738);
nor U5471 (N_5471,N_1157,N_2021);
nor U5472 (N_5472,N_3093,N_431);
xnor U5473 (N_5473,N_2229,N_4581);
nor U5474 (N_5474,N_667,N_1888);
and U5475 (N_5475,N_1919,N_4740);
nand U5476 (N_5476,N_194,N_1811);
or U5477 (N_5477,N_2442,N_4486);
nor U5478 (N_5478,N_735,N_775);
nor U5479 (N_5479,N_1292,N_20);
nor U5480 (N_5480,N_3065,N_2611);
nand U5481 (N_5481,N_2744,N_3987);
or U5482 (N_5482,N_4030,N_637);
nand U5483 (N_5483,N_3926,N_2669);
or U5484 (N_5484,N_4076,N_3840);
or U5485 (N_5485,N_3990,N_3503);
and U5486 (N_5486,N_3139,N_4832);
xnor U5487 (N_5487,N_86,N_2580);
or U5488 (N_5488,N_3715,N_360);
and U5489 (N_5489,N_485,N_2620);
xnor U5490 (N_5490,N_4843,N_4541);
xor U5491 (N_5491,N_4421,N_786);
or U5492 (N_5492,N_2411,N_202);
nor U5493 (N_5493,N_753,N_4629);
or U5494 (N_5494,N_2296,N_2352);
or U5495 (N_5495,N_3313,N_4217);
or U5496 (N_5496,N_3825,N_4874);
xnor U5497 (N_5497,N_1839,N_1398);
or U5498 (N_5498,N_4018,N_4719);
nor U5499 (N_5499,N_4084,N_452);
and U5500 (N_5500,N_2280,N_1050);
or U5501 (N_5501,N_3631,N_876);
nand U5502 (N_5502,N_3451,N_190);
or U5503 (N_5503,N_4238,N_3432);
or U5504 (N_5504,N_249,N_3884);
or U5505 (N_5505,N_2271,N_3585);
or U5506 (N_5506,N_1172,N_2032);
and U5507 (N_5507,N_114,N_1756);
nor U5508 (N_5508,N_3196,N_1835);
nand U5509 (N_5509,N_576,N_377);
nand U5510 (N_5510,N_960,N_123);
xnor U5511 (N_5511,N_4507,N_3117);
nor U5512 (N_5512,N_733,N_4578);
nor U5513 (N_5513,N_2498,N_3675);
nand U5514 (N_5514,N_2103,N_1586);
or U5515 (N_5515,N_2724,N_4417);
nand U5516 (N_5516,N_483,N_1475);
xnor U5517 (N_5517,N_544,N_2923);
xnor U5518 (N_5518,N_1240,N_326);
and U5519 (N_5519,N_2518,N_1197);
or U5520 (N_5520,N_3980,N_1193);
and U5521 (N_5521,N_2819,N_4090);
and U5522 (N_5522,N_877,N_4531);
xnor U5523 (N_5523,N_2507,N_299);
xor U5524 (N_5524,N_4770,N_2206);
nand U5525 (N_5525,N_4307,N_2022);
and U5526 (N_5526,N_956,N_1717);
and U5527 (N_5527,N_728,N_2967);
nor U5528 (N_5528,N_2098,N_2654);
nand U5529 (N_5529,N_2721,N_3311);
or U5530 (N_5530,N_1511,N_2780);
xnor U5531 (N_5531,N_2479,N_1797);
or U5532 (N_5532,N_1535,N_166);
nor U5533 (N_5533,N_3166,N_3597);
nor U5534 (N_5534,N_1354,N_1971);
and U5535 (N_5535,N_1146,N_4635);
and U5536 (N_5536,N_4151,N_2787);
nor U5537 (N_5537,N_3192,N_3763);
and U5538 (N_5538,N_2197,N_3037);
nand U5539 (N_5539,N_4091,N_55);
nand U5540 (N_5540,N_149,N_2294);
nand U5541 (N_5541,N_3637,N_3208);
xnor U5542 (N_5542,N_3205,N_512);
nand U5543 (N_5543,N_701,N_2309);
xor U5544 (N_5544,N_4190,N_1319);
xnor U5545 (N_5545,N_823,N_3469);
nor U5546 (N_5546,N_4372,N_2313);
and U5547 (N_5547,N_3896,N_3395);
nand U5548 (N_5548,N_2505,N_4349);
and U5549 (N_5549,N_902,N_16);
nor U5550 (N_5550,N_1794,N_4450);
nor U5551 (N_5551,N_1181,N_4164);
or U5552 (N_5552,N_4028,N_2111);
nor U5553 (N_5553,N_4726,N_137);
xor U5554 (N_5554,N_2375,N_4582);
and U5555 (N_5555,N_260,N_227);
or U5556 (N_5556,N_2143,N_932);
nand U5557 (N_5557,N_1899,N_1725);
nand U5558 (N_5558,N_3204,N_397);
or U5559 (N_5559,N_4235,N_2597);
xor U5560 (N_5560,N_2316,N_817);
nand U5561 (N_5561,N_2799,N_2440);
nand U5562 (N_5562,N_706,N_4107);
nand U5563 (N_5563,N_1046,N_1739);
nor U5564 (N_5564,N_3460,N_3420);
nand U5565 (N_5565,N_1022,N_1321);
nand U5566 (N_5566,N_1440,N_315);
or U5567 (N_5567,N_3671,N_3665);
and U5568 (N_5568,N_930,N_1627);
or U5569 (N_5569,N_3710,N_880);
xnor U5570 (N_5570,N_4652,N_4675);
xnor U5571 (N_5571,N_3038,N_3240);
nor U5572 (N_5572,N_2536,N_382);
nand U5573 (N_5573,N_3797,N_1692);
nor U5574 (N_5574,N_91,N_109);
and U5575 (N_5575,N_3815,N_874);
xor U5576 (N_5576,N_4817,N_2317);
nor U5577 (N_5577,N_3696,N_2458);
xor U5578 (N_5578,N_1068,N_104);
or U5579 (N_5579,N_2656,N_2714);
or U5580 (N_5580,N_330,N_2992);
xor U5581 (N_5581,N_3601,N_3388);
nor U5582 (N_5582,N_3112,N_501);
and U5583 (N_5583,N_4109,N_1957);
or U5584 (N_5584,N_3413,N_1767);
nand U5585 (N_5585,N_1843,N_1708);
or U5586 (N_5586,N_2871,N_1219);
xnor U5587 (N_5587,N_3863,N_3245);
nor U5588 (N_5588,N_4024,N_717);
nor U5589 (N_5589,N_3146,N_2743);
or U5590 (N_5590,N_133,N_4053);
or U5591 (N_5591,N_4772,N_3161);
nor U5592 (N_5592,N_683,N_2039);
or U5593 (N_5593,N_3748,N_1528);
nand U5594 (N_5594,N_3495,N_2682);
nand U5595 (N_5595,N_2575,N_441);
or U5596 (N_5596,N_650,N_855);
nor U5597 (N_5597,N_3389,N_1521);
nand U5598 (N_5598,N_2938,N_1600);
nand U5599 (N_5599,N_3181,N_2841);
and U5600 (N_5600,N_4300,N_1147);
or U5601 (N_5601,N_1438,N_916);
xor U5602 (N_5602,N_3573,N_27);
nor U5603 (N_5603,N_4981,N_3849);
nand U5604 (N_5604,N_1609,N_4503);
and U5605 (N_5605,N_3689,N_1632);
xnor U5606 (N_5606,N_1596,N_2838);
nor U5607 (N_5607,N_3371,N_2527);
xnor U5608 (N_5608,N_3569,N_53);
and U5609 (N_5609,N_1386,N_3835);
and U5610 (N_5610,N_1416,N_3491);
and U5611 (N_5611,N_3529,N_4330);
nor U5612 (N_5612,N_4029,N_4947);
or U5613 (N_5613,N_1370,N_3446);
or U5614 (N_5614,N_3663,N_1373);
nor U5615 (N_5615,N_3616,N_1599);
nor U5616 (N_5616,N_25,N_3730);
nand U5617 (N_5617,N_2947,N_782);
and U5618 (N_5618,N_2396,N_195);
and U5619 (N_5619,N_84,N_4899);
nor U5620 (N_5620,N_2362,N_3203);
nor U5621 (N_5621,N_4294,N_2753);
nor U5622 (N_5622,N_2384,N_3975);
nand U5623 (N_5623,N_1444,N_4424);
xnor U5624 (N_5624,N_784,N_619);
xnor U5625 (N_5625,N_2210,N_2914);
nor U5626 (N_5626,N_4495,N_2627);
nand U5627 (N_5627,N_1701,N_2849);
and U5628 (N_5628,N_4936,N_857);
nand U5629 (N_5629,N_1133,N_494);
xnor U5630 (N_5630,N_3418,N_1374);
and U5631 (N_5631,N_2377,N_4463);
nor U5632 (N_5632,N_1564,N_1279);
nor U5633 (N_5633,N_4871,N_1740);
xor U5634 (N_5634,N_3932,N_3225);
nor U5635 (N_5635,N_3261,N_2681);
nand U5636 (N_5636,N_3427,N_4888);
and U5637 (N_5637,N_4251,N_2488);
xor U5638 (N_5638,N_4756,N_2120);
and U5639 (N_5639,N_2061,N_3377);
nor U5640 (N_5640,N_3903,N_3739);
nor U5641 (N_5641,N_4317,N_2482);
xnor U5642 (N_5642,N_1643,N_698);
and U5643 (N_5643,N_2772,N_1305);
and U5644 (N_5644,N_4968,N_3239);
nor U5645 (N_5645,N_3448,N_154);
or U5646 (N_5646,N_4766,N_1624);
nor U5647 (N_5647,N_2265,N_4083);
or U5648 (N_5648,N_2695,N_3902);
xor U5649 (N_5649,N_3376,N_3283);
nor U5650 (N_5650,N_173,N_767);
xor U5651 (N_5651,N_4949,N_2894);
xnor U5652 (N_5652,N_3398,N_164);
xnor U5653 (N_5653,N_1714,N_4513);
nor U5654 (N_5654,N_2100,N_1577);
xor U5655 (N_5655,N_82,N_2171);
or U5656 (N_5656,N_402,N_4351);
nor U5657 (N_5657,N_3624,N_1697);
nand U5658 (N_5658,N_1503,N_3162);
xor U5659 (N_5659,N_938,N_3163);
or U5660 (N_5660,N_2152,N_1569);
xnor U5661 (N_5661,N_3246,N_3777);
xor U5662 (N_5662,N_3297,N_3984);
nor U5663 (N_5663,N_4984,N_925);
and U5664 (N_5664,N_1188,N_3148);
xnor U5665 (N_5665,N_3220,N_1184);
or U5666 (N_5666,N_4589,N_2269);
and U5667 (N_5667,N_4192,N_3524);
nand U5668 (N_5668,N_3583,N_4252);
nor U5669 (N_5669,N_3497,N_4427);
or U5670 (N_5670,N_4033,N_3784);
nor U5671 (N_5671,N_673,N_358);
xnor U5672 (N_5672,N_2842,N_533);
and U5673 (N_5673,N_2383,N_1071);
nand U5674 (N_5674,N_2332,N_561);
or U5675 (N_5675,N_278,N_1450);
nor U5676 (N_5676,N_3025,N_1817);
nand U5677 (N_5677,N_1786,N_1993);
or U5678 (N_5678,N_1426,N_2875);
and U5679 (N_5679,N_3434,N_1636);
xor U5680 (N_5680,N_4277,N_4549);
and U5681 (N_5681,N_4546,N_1759);
xor U5682 (N_5682,N_2151,N_4381);
nor U5683 (N_5683,N_3639,N_3526);
nor U5684 (N_5684,N_4390,N_3227);
or U5685 (N_5685,N_4751,N_340);
or U5686 (N_5686,N_1343,N_4697);
nor U5687 (N_5687,N_4490,N_68);
or U5688 (N_5688,N_3026,N_3077);
nand U5689 (N_5689,N_2493,N_2183);
or U5690 (N_5690,N_69,N_924);
nor U5691 (N_5691,N_1243,N_1897);
xnor U5692 (N_5692,N_1176,N_245);
nand U5693 (N_5693,N_1463,N_661);
xnor U5694 (N_5694,N_1042,N_2371);
or U5695 (N_5695,N_3435,N_2905);
and U5696 (N_5696,N_4670,N_3519);
or U5697 (N_5697,N_3229,N_891);
xnor U5698 (N_5698,N_3327,N_2256);
xnor U5699 (N_5699,N_413,N_1695);
nor U5700 (N_5700,N_743,N_10);
or U5701 (N_5701,N_2979,N_4934);
nor U5702 (N_5702,N_2414,N_4410);
xor U5703 (N_5703,N_746,N_2419);
nor U5704 (N_5704,N_3862,N_2948);
or U5705 (N_5705,N_4142,N_357);
nand U5706 (N_5706,N_4889,N_4452);
nor U5707 (N_5707,N_4290,N_351);
xnor U5708 (N_5708,N_2642,N_1885);
xnor U5709 (N_5709,N_2716,N_395);
or U5710 (N_5710,N_1159,N_3372);
nor U5711 (N_5711,N_60,N_1415);
nand U5712 (N_5712,N_740,N_4111);
and U5713 (N_5713,N_2685,N_2750);
nor U5714 (N_5714,N_1195,N_1785);
nand U5715 (N_5715,N_1399,N_3410);
nor U5716 (N_5716,N_4340,N_4355);
nor U5717 (N_5717,N_1529,N_3792);
xnor U5718 (N_5718,N_3108,N_2216);
nand U5719 (N_5719,N_1340,N_3488);
nor U5720 (N_5720,N_148,N_4547);
and U5721 (N_5721,N_1363,N_1690);
xor U5722 (N_5722,N_4202,N_844);
xor U5723 (N_5723,N_811,N_993);
and U5724 (N_5724,N_3578,N_1640);
or U5725 (N_5725,N_3071,N_1959);
nor U5726 (N_5726,N_3699,N_531);
nand U5727 (N_5727,N_18,N_4327);
nand U5728 (N_5728,N_4416,N_28);
xnor U5729 (N_5729,N_4638,N_4115);
or U5730 (N_5730,N_513,N_3176);
and U5731 (N_5731,N_4767,N_75);
and U5732 (N_5732,N_115,N_4046);
nor U5733 (N_5733,N_2127,N_4536);
xnor U5734 (N_5734,N_2388,N_338);
nor U5735 (N_5735,N_1244,N_4268);
and U5736 (N_5736,N_1742,N_392);
nand U5737 (N_5737,N_1560,N_1988);
and U5738 (N_5738,N_4544,N_3544);
nand U5739 (N_5739,N_4473,N_4710);
xor U5740 (N_5740,N_4712,N_1127);
or U5741 (N_5741,N_3102,N_4049);
nor U5742 (N_5742,N_2025,N_3348);
or U5743 (N_5743,N_100,N_2175);
or U5744 (N_5744,N_3979,N_626);
nor U5745 (N_5745,N_1358,N_638);
nand U5746 (N_5746,N_787,N_3737);
and U5747 (N_5747,N_2246,N_792);
and U5748 (N_5748,N_2134,N_48);
nor U5749 (N_5749,N_246,N_2826);
and U5750 (N_5750,N_1153,N_2298);
xor U5751 (N_5751,N_146,N_555);
and U5752 (N_5752,N_3256,N_4240);
nand U5753 (N_5753,N_1902,N_3557);
xnor U5754 (N_5754,N_1576,N_3978);
nor U5755 (N_5755,N_4901,N_4358);
xor U5756 (N_5756,N_4181,N_1448);
or U5757 (N_5757,N_3127,N_4433);
xnor U5758 (N_5758,N_4600,N_2077);
xor U5759 (N_5759,N_1065,N_1937);
or U5760 (N_5760,N_4979,N_3531);
or U5761 (N_5761,N_600,N_254);
nor U5762 (N_5762,N_3149,N_4779);
or U5763 (N_5763,N_4158,N_1610);
and U5764 (N_5764,N_2847,N_4614);
nand U5765 (N_5765,N_3001,N_725);
nand U5766 (N_5766,N_4316,N_2510);
and U5767 (N_5767,N_3087,N_1360);
nor U5768 (N_5768,N_36,N_1603);
nand U5769 (N_5769,N_1518,N_1381);
nor U5770 (N_5770,N_2506,N_2590);
or U5771 (N_5771,N_1391,N_61);
nand U5772 (N_5772,N_2102,N_4644);
nor U5773 (N_5773,N_3213,N_2639);
nand U5774 (N_5774,N_1089,N_1458);
or U5775 (N_5775,N_2987,N_1755);
and U5776 (N_5776,N_3613,N_253);
xnor U5777 (N_5777,N_1232,N_4607);
and U5778 (N_5778,N_4833,N_468);
xor U5779 (N_5779,N_4502,N_1198);
and U5780 (N_5780,N_2457,N_3951);
or U5781 (N_5781,N_1710,N_3928);
and U5782 (N_5782,N_3135,N_4796);
nand U5783 (N_5783,N_1051,N_1663);
or U5784 (N_5784,N_248,N_2236);
or U5785 (N_5785,N_1825,N_1588);
nor U5786 (N_5786,N_1404,N_2892);
nand U5787 (N_5787,N_266,N_3177);
or U5788 (N_5788,N_4432,N_4599);
and U5789 (N_5789,N_3528,N_4391);
or U5790 (N_5790,N_385,N_589);
xnor U5791 (N_5791,N_2818,N_4545);
and U5792 (N_5792,N_1533,N_1486);
nand U5793 (N_5793,N_4034,N_3235);
and U5794 (N_5794,N_224,N_1247);
or U5795 (N_5795,N_3326,N_4462);
and U5796 (N_5796,N_4196,N_4376);
nand U5797 (N_5797,N_4850,N_726);
or U5798 (N_5798,N_163,N_998);
xor U5799 (N_5799,N_4723,N_5);
nor U5800 (N_5800,N_4902,N_1234);
xor U5801 (N_5801,N_222,N_2012);
nand U5802 (N_5802,N_4141,N_1750);
or U5803 (N_5803,N_4521,N_44);
and U5804 (N_5804,N_2113,N_887);
and U5805 (N_5805,N_257,N_3141);
and U5806 (N_5806,N_3705,N_3697);
and U5807 (N_5807,N_3336,N_4078);
or U5808 (N_5808,N_4288,N_4244);
nor U5809 (N_5809,N_2002,N_4441);
nor U5810 (N_5810,N_4927,N_1420);
or U5811 (N_5811,N_4499,N_3592);
and U5812 (N_5812,N_4067,N_721);
nand U5813 (N_5813,N_1947,N_820);
and U5814 (N_5814,N_3559,N_4941);
nand U5815 (N_5815,N_2822,N_1302);
nor U5816 (N_5816,N_3591,N_4840);
nand U5817 (N_5817,N_1250,N_4512);
nor U5818 (N_5818,N_1326,N_1114);
or U5819 (N_5819,N_1392,N_2399);
or U5820 (N_5820,N_4086,N_2408);
or U5821 (N_5821,N_3344,N_3356);
and U5822 (N_5822,N_4040,N_1294);
nand U5823 (N_5823,N_4469,N_4274);
nor U5824 (N_5824,N_1548,N_2940);
or U5825 (N_5825,N_991,N_3222);
or U5826 (N_5826,N_1497,N_3493);
xor U5827 (N_5827,N_934,N_3426);
nor U5828 (N_5828,N_1849,N_4367);
or U5829 (N_5829,N_33,N_708);
nand U5830 (N_5830,N_3664,N_1023);
and U5831 (N_5831,N_3265,N_1964);
nand U5832 (N_5832,N_1478,N_677);
xor U5833 (N_5833,N_2658,N_4952);
or U5834 (N_5834,N_1081,N_783);
xnor U5835 (N_5835,N_3575,N_4241);
and U5836 (N_5836,N_4820,N_4975);
nand U5837 (N_5837,N_1323,N_1477);
xor U5838 (N_5838,N_2528,N_3477);
nand U5839 (N_5839,N_2539,N_2118);
and U5840 (N_5840,N_98,N_3338);
or U5841 (N_5841,N_4308,N_479);
and U5842 (N_5842,N_4587,N_3212);
nor U5843 (N_5843,N_3686,N_450);
xnor U5844 (N_5844,N_4672,N_4135);
and U5845 (N_5845,N_4257,N_4551);
xor U5846 (N_5846,N_4725,N_671);
nor U5847 (N_5847,N_4803,N_2777);
nor U5848 (N_5848,N_3537,N_1397);
or U5849 (N_5849,N_4575,N_3846);
nand U5850 (N_5850,N_1987,N_4977);
nor U5851 (N_5851,N_2041,N_197);
and U5852 (N_5852,N_1182,N_3651);
nor U5853 (N_5853,N_665,N_4509);
nor U5854 (N_5854,N_4163,N_1862);
and U5855 (N_5855,N_3211,N_4938);
and U5856 (N_5856,N_218,N_1233);
nand U5857 (N_5857,N_2832,N_1465);
and U5858 (N_5858,N_704,N_4718);
xor U5859 (N_5859,N_3099,N_2040);
nand U5860 (N_5860,N_1912,N_2509);
nor U5861 (N_5861,N_2023,N_119);
and U5862 (N_5862,N_3050,N_984);
nand U5863 (N_5863,N_921,N_2101);
xnor U5864 (N_5864,N_1665,N_2232);
xnor U5865 (N_5865,N_4569,N_3844);
nor U5866 (N_5866,N_1033,N_4361);
nand U5867 (N_5867,N_1013,N_1410);
nor U5868 (N_5868,N_4106,N_2804);
nor U5869 (N_5869,N_1421,N_3656);
and U5870 (N_5870,N_3317,N_1748);
xnor U5871 (N_5871,N_4379,N_3252);
or U5872 (N_5872,N_1838,N_2544);
and U5873 (N_5873,N_4553,N_824);
nand U5874 (N_5874,N_1460,N_1864);
xnor U5875 (N_5875,N_4112,N_752);
and U5876 (N_5876,N_3009,N_1016);
xor U5877 (N_5877,N_2796,N_3151);
nor U5878 (N_5878,N_2712,N_3069);
xnor U5879 (N_5879,N_498,N_3514);
nand U5880 (N_5880,N_3732,N_3857);
nand U5881 (N_5881,N_4062,N_562);
nand U5882 (N_5882,N_1681,N_4023);
nand U5883 (N_5883,N_4144,N_682);
xnor U5884 (N_5884,N_809,N_3567);
nand U5885 (N_5885,N_211,N_4218);
and U5886 (N_5886,N_3944,N_2299);
and U5887 (N_5887,N_2728,N_1870);
nand U5888 (N_5888,N_2472,N_1539);
xnor U5889 (N_5889,N_4388,N_97);
nand U5890 (N_5890,N_2706,N_1138);
nor U5891 (N_5891,N_3820,N_4857);
nand U5892 (N_5892,N_598,N_3132);
xnor U5893 (N_5893,N_1029,N_3119);
or U5894 (N_5894,N_4804,N_3778);
and U5895 (N_5895,N_4606,N_2017);
or U5896 (N_5896,N_244,N_3072);
xor U5897 (N_5897,N_1163,N_4405);
and U5898 (N_5898,N_2844,N_1920);
and U5899 (N_5899,N_4855,N_4050);
nand U5900 (N_5900,N_4967,N_1385);
xnor U5901 (N_5901,N_1808,N_325);
or U5902 (N_5902,N_4001,N_1691);
nand U5903 (N_5903,N_2884,N_2460);
and U5904 (N_5904,N_462,N_4913);
or U5905 (N_5905,N_3655,N_3726);
and U5906 (N_5906,N_297,N_1093);
nor U5907 (N_5907,N_4072,N_1052);
or U5908 (N_5908,N_1948,N_797);
xnor U5909 (N_5909,N_2720,N_4085);
xor U5910 (N_5910,N_1097,N_4384);
xnor U5911 (N_5911,N_3121,N_259);
nor U5912 (N_5912,N_2551,N_4627);
or U5913 (N_5913,N_649,N_159);
nand U5914 (N_5914,N_1185,N_1254);
nor U5915 (N_5915,N_1587,N_3713);
nor U5916 (N_5916,N_3676,N_2461);
nor U5917 (N_5917,N_2601,N_1251);
xor U5918 (N_5918,N_1787,N_4171);
or U5919 (N_5919,N_1732,N_2775);
nor U5920 (N_5920,N_2281,N_4264);
nor U5921 (N_5921,N_2645,N_305);
and U5922 (N_5922,N_2566,N_1949);
or U5923 (N_5923,N_2687,N_3994);
xor U5924 (N_5924,N_2585,N_3725);
nand U5925 (N_5925,N_1283,N_1160);
and U5926 (N_5926,N_4732,N_3234);
nor U5927 (N_5927,N_4570,N_3672);
nor U5928 (N_5928,N_4721,N_2993);
or U5929 (N_5929,N_4476,N_110);
nand U5930 (N_5930,N_612,N_1451);
xor U5931 (N_5931,N_4527,N_546);
xor U5932 (N_5932,N_2110,N_1806);
xor U5933 (N_5933,N_862,N_1938);
and U5934 (N_5934,N_2087,N_1793);
xor U5935 (N_5935,N_4270,N_2511);
nand U5936 (N_5936,N_3906,N_140);
nor U5937 (N_5937,N_3110,N_745);
xnor U5938 (N_5938,N_4762,N_1520);
nand U5939 (N_5939,N_463,N_2303);
xnor U5940 (N_5940,N_2758,N_1880);
nand U5941 (N_5941,N_1400,N_4138);
nand U5942 (N_5942,N_2562,N_2870);
xor U5943 (N_5943,N_1224,N_1236);
xor U5944 (N_5944,N_3023,N_514);
nor U5945 (N_5945,N_1939,N_2354);
nor U5946 (N_5946,N_4273,N_4759);
or U5947 (N_5947,N_2186,N_3425);
and U5948 (N_5948,N_243,N_38);
and U5949 (N_5949,N_748,N_3094);
and U5950 (N_5950,N_3367,N_4116);
nand U5951 (N_5951,N_2049,N_1446);
nand U5952 (N_5952,N_2456,N_4065);
nand U5953 (N_5953,N_1265,N_4624);
nor U5954 (N_5954,N_2779,N_59);
nand U5955 (N_5955,N_4500,N_936);
nand U5956 (N_5956,N_2144,N_711);
xnor U5957 (N_5957,N_926,N_4813);
nand U5958 (N_5958,N_3000,N_3134);
nor U5959 (N_5959,N_3450,N_4689);
nand U5960 (N_5960,N_1647,N_1903);
nand U5961 (N_5961,N_2650,N_3055);
xnor U5962 (N_5962,N_4055,N_1320);
xnor U5963 (N_5963,N_3277,N_2561);
xor U5964 (N_5964,N_1914,N_962);
xor U5965 (N_5965,N_4645,N_3075);
nand U5966 (N_5966,N_2170,N_881);
or U5967 (N_5967,N_3172,N_4236);
or U5968 (N_5968,N_1776,N_4906);
or U5969 (N_5969,N_723,N_3345);
xnor U5970 (N_5970,N_3749,N_1589);
or U5971 (N_5971,N_606,N_3536);
and U5972 (N_5972,N_904,N_3946);
and U5973 (N_5973,N_1612,N_1393);
nor U5974 (N_5974,N_4656,N_3351);
or U5975 (N_5975,N_2218,N_4641);
xnor U5976 (N_5976,N_4296,N_2981);
nor U5977 (N_5977,N_4976,N_3242);
nor U5978 (N_5978,N_3105,N_3666);
nor U5979 (N_5979,N_410,N_4411);
or U5980 (N_5980,N_2792,N_4131);
nand U5981 (N_5981,N_515,N_3237);
or U5982 (N_5982,N_1562,N_4108);
and U5983 (N_5983,N_1645,N_601);
nand U5984 (N_5984,N_3325,N_4637);
or U5985 (N_5985,N_4226,N_4324);
nand U5986 (N_5986,N_1334,N_4148);
nand U5987 (N_5987,N_3904,N_3218);
and U5988 (N_5988,N_1799,N_1418);
nor U5989 (N_5989,N_1288,N_2465);
nor U5990 (N_5990,N_2808,N_3680);
nand U5991 (N_5991,N_1007,N_1423);
nor U5992 (N_5992,N_2578,N_3924);
nor U5993 (N_5993,N_534,N_3888);
nand U5994 (N_5994,N_4059,N_3988);
nor U5995 (N_5995,N_2435,N_617);
and U5996 (N_5996,N_1951,N_2277);
and U5997 (N_5997,N_2891,N_4263);
nor U5998 (N_5998,N_317,N_951);
and U5999 (N_5999,N_4567,N_2651);
xor U6000 (N_6000,N_3814,N_1952);
nor U6001 (N_6001,N_1648,N_1989);
and U6002 (N_6002,N_3627,N_680);
nor U6003 (N_6003,N_496,N_3143);
nand U6004 (N_6004,N_1099,N_765);
nor U6005 (N_6005,N_116,N_777);
and U6006 (N_6006,N_1216,N_1053);
or U6007 (N_6007,N_1403,N_1711);
nand U6008 (N_6008,N_4212,N_1928);
nand U6009 (N_6009,N_2048,N_4649);
xnor U6010 (N_6010,N_3913,N_3236);
xor U6011 (N_6011,N_3190,N_3621);
or U6012 (N_6012,N_781,N_199);
or U6013 (N_6013,N_4063,N_2609);
and U6014 (N_6014,N_3786,N_3045);
nor U6015 (N_6015,N_3996,N_3605);
nand U6016 (N_6016,N_584,N_1190);
nor U6017 (N_6017,N_3078,N_3850);
or U6018 (N_6018,N_4459,N_3625);
or U6019 (N_6019,N_181,N_1456);
nand U6020 (N_6020,N_3404,N_3533);
xnor U6021 (N_6021,N_4418,N_3992);
or U6022 (N_6022,N_4359,N_3076);
and U6023 (N_6023,N_4454,N_1506);
nor U6024 (N_6024,N_3678,N_1223);
nor U6025 (N_6025,N_1833,N_1327);
and U6026 (N_6026,N_205,N_4352);
or U6027 (N_6027,N_4200,N_4465);
nor U6028 (N_6028,N_1335,N_3457);
and U6029 (N_6029,N_4434,N_4835);
and U6030 (N_6030,N_4933,N_3468);
nor U6031 (N_6031,N_1032,N_73);
and U6032 (N_6032,N_2052,N_1226);
xnor U6033 (N_6033,N_3588,N_4921);
nor U6034 (N_6034,N_2394,N_2634);
nand U6035 (N_6035,N_1258,N_2858);
and U6036 (N_6036,N_2784,N_3466);
nand U6037 (N_6037,N_2433,N_3019);
xor U6038 (N_6038,N_4003,N_187);
nor U6039 (N_6039,N_420,N_3733);
nor U6040 (N_6040,N_2204,N_1871);
nand U6041 (N_6041,N_3940,N_791);
nand U6042 (N_6042,N_1116,N_3614);
or U6043 (N_6043,N_3579,N_2056);
nand U6044 (N_6044,N_3895,N_818);
nor U6045 (N_6045,N_4146,N_3320);
xnor U6046 (N_6046,N_3216,N_2602);
nand U6047 (N_6047,N_4566,N_1943);
or U6048 (N_6048,N_4477,N_995);
xor U6049 (N_6049,N_3669,N_3288);
nand U6050 (N_6050,N_3541,N_3922);
or U6051 (N_6051,N_3339,N_3948);
xnor U6052 (N_6052,N_67,N_1161);
xor U6053 (N_6053,N_1955,N_4847);
xor U6054 (N_6054,N_4382,N_215);
xor U6055 (N_6055,N_3443,N_1601);
nor U6056 (N_6056,N_1019,N_443);
and U6057 (N_6057,N_4808,N_3219);
nor U6058 (N_6058,N_2013,N_2390);
or U6059 (N_6059,N_1967,N_2786);
and U6060 (N_6060,N_3599,N_399);
and U6061 (N_6061,N_2806,N_4530);
nand U6062 (N_6062,N_4558,N_4811);
nor U6063 (N_6063,N_2532,N_2168);
and U6064 (N_6064,N_3096,N_320);
and U6065 (N_6065,N_2260,N_530);
xnor U6066 (N_6066,N_3603,N_376);
xnor U6067 (N_6067,N_2042,N_622);
and U6068 (N_6068,N_3270,N_3024);
nor U6069 (N_6069,N_232,N_2554);
xnor U6070 (N_6070,N_3534,N_1664);
or U6071 (N_6071,N_419,N_3885);
nor U6072 (N_6072,N_893,N_986);
or U6073 (N_6073,N_1659,N_2279);
and U6074 (N_6074,N_511,N_4147);
nand U6075 (N_6075,N_3774,N_4736);
nand U6076 (N_6076,N_2348,N_1230);
xnor U6077 (N_6077,N_3390,N_906);
or U6078 (N_6078,N_2258,N_1639);
nand U6079 (N_6079,N_3408,N_1918);
or U6080 (N_6080,N_2198,N_319);
xor U6081 (N_6081,N_210,N_3285);
nor U6082 (N_6082,N_2356,N_3886);
xnor U6083 (N_6083,N_1653,N_2810);
or U6084 (N_6084,N_362,N_2719);
or U6085 (N_6085,N_4881,N_4255);
and U6086 (N_6086,N_988,N_3361);
or U6087 (N_6087,N_2641,N_920);
and U6088 (N_6088,N_1905,N_550);
xor U6089 (N_6089,N_2717,N_4501);
or U6090 (N_6090,N_3296,N_1201);
and U6091 (N_6091,N_3991,N_306);
xnor U6092 (N_6092,N_2485,N_2165);
and U6093 (N_6093,N_4665,N_3142);
xor U6094 (N_6094,N_4073,N_1873);
nor U6095 (N_6095,N_3982,N_4301);
or U6096 (N_6096,N_3756,N_571);
nand U6097 (N_6097,N_3545,N_1637);
nand U6098 (N_6098,N_277,N_364);
and U6099 (N_6099,N_4139,N_3008);
nor U6100 (N_6100,N_4409,N_4309);
or U6101 (N_6101,N_3855,N_3114);
nand U6102 (N_6102,N_2305,N_3540);
or U6103 (N_6103,N_3860,N_2868);
nor U6104 (N_6104,N_4660,N_611);
nor U6105 (N_6105,N_1096,N_945);
nand U6106 (N_6106,N_1898,N_3262);
and U6107 (N_6107,N_1369,N_265);
and U6108 (N_6108,N_3518,N_3030);
and U6109 (N_6109,N_3363,N_1105);
xor U6110 (N_6110,N_1194,N_1981);
xor U6111 (N_6111,N_4837,N_3823);
xnor U6112 (N_6112,N_3414,N_252);
nand U6113 (N_6113,N_843,N_4077);
nor U6114 (N_6114,N_129,N_4020);
xnor U6115 (N_6115,N_171,N_1125);
nand U6116 (N_6116,N_3400,N_1893);
nand U6117 (N_6117,N_3643,N_2557);
and U6118 (N_6118,N_2001,N_3243);
and U6119 (N_6119,N_3073,N_2003);
nand U6120 (N_6120,N_344,N_3610);
nand U6121 (N_6121,N_2107,N_3131);
nand U6122 (N_6122,N_2018,N_4103);
and U6123 (N_6123,N_3020,N_3811);
nand U6124 (N_6124,N_2473,N_4298);
xnor U6125 (N_6125,N_1306,N_691);
xnor U6126 (N_6126,N_408,N_3501);
nand U6127 (N_6127,N_1807,N_4408);
nor U6128 (N_6128,N_3861,N_3740);
nor U6129 (N_6129,N_3813,N_2109);
nand U6130 (N_6130,N_4345,N_3934);
nor U6131 (N_6131,N_2084,N_4211);
nand U6132 (N_6132,N_2468,N_4333);
nor U6133 (N_6133,N_822,N_2881);
nor U6134 (N_6134,N_165,N_3821);
or U6135 (N_6135,N_3539,N_1953);
or U6136 (N_6136,N_1337,N_2768);
nand U6137 (N_6137,N_1262,N_1509);
nand U6138 (N_6138,N_394,N_833);
or U6139 (N_6139,N_1345,N_4677);
nor U6140 (N_6140,N_1213,N_3674);
and U6141 (N_6141,N_2946,N_2463);
or U6142 (N_6142,N_2666,N_1094);
xnor U6143 (N_6143,N_1273,N_4866);
xor U6144 (N_6144,N_2735,N_3841);
and U6145 (N_6145,N_1141,N_2550);
and U6146 (N_6146,N_3304,N_944);
nor U6147 (N_6147,N_2370,N_3735);
and U6148 (N_6148,N_1479,N_1118);
nor U6149 (N_6149,N_2688,N_12);
or U6150 (N_6150,N_1173,N_3826);
nor U6151 (N_6151,N_2274,N_3761);
and U6152 (N_6152,N_4203,N_3029);
nor U6153 (N_6153,N_1579,N_4590);
or U6154 (N_6154,N_2024,N_3039);
or U6155 (N_6155,N_1339,N_4346);
or U6156 (N_6156,N_3215,N_4806);
or U6157 (N_6157,N_4258,N_4959);
xnor U6158 (N_6158,N_2982,N_415);
xor U6159 (N_6159,N_1552,N_3224);
nor U6160 (N_6160,N_4031,N_428);
nor U6161 (N_6161,N_2273,N_2126);
xor U6162 (N_6162,N_1445,N_1760);
nand U6163 (N_6163,N_1854,N_2252);
nor U6164 (N_6164,N_2389,N_1960);
nor U6165 (N_6165,N_1557,N_4768);
xor U6166 (N_6166,N_2268,N_4170);
xnor U6167 (N_6167,N_669,N_2860);
xnor U6168 (N_6168,N_918,N_2825);
nor U6169 (N_6169,N_1850,N_764);
or U6170 (N_6170,N_2104,N_4485);
xnor U6171 (N_6171,N_1956,N_1651);
or U6172 (N_6172,N_126,N_3120);
and U6173 (N_6173,N_2555,N_2016);
or U6174 (N_6174,N_4622,N_2683);
and U6175 (N_6175,N_2492,N_2400);
and U6176 (N_6176,N_2363,N_106);
xnor U6177 (N_6177,N_2028,N_1754);
or U6178 (N_6178,N_2738,N_4113);
nor U6179 (N_6179,N_1045,N_101);
xor U6180 (N_6180,N_3040,N_3043);
nor U6181 (N_6181,N_922,N_23);
xor U6182 (N_6182,N_2989,N_2701);
or U6183 (N_6183,N_2836,N_3416);
nor U6184 (N_6184,N_656,N_1264);
xnor U6185 (N_6185,N_851,N_486);
xnor U6186 (N_6186,N_2671,N_4233);
or U6187 (N_6187,N_3852,N_4362);
or U6188 (N_6188,N_172,N_4201);
or U6189 (N_6189,N_3681,N_4709);
and U6190 (N_6190,N_2969,N_3560);
nor U6191 (N_6191,N_11,N_3138);
nor U6192 (N_6192,N_1220,N_3286);
xor U6193 (N_6193,N_2235,N_1344);
xor U6194 (N_6194,N_1617,N_1205);
xnor U6195 (N_6195,N_3028,N_1573);
and U6196 (N_6196,N_700,N_293);
and U6197 (N_6197,N_2219,N_2194);
or U6198 (N_6198,N_3111,N_4189);
nor U6199 (N_6199,N_912,N_1848);
or U6200 (N_6200,N_4827,N_416);
xnor U6201 (N_6201,N_3255,N_63);
nand U6202 (N_6202,N_467,N_3822);
nor U6203 (N_6203,N_4336,N_3331);
nor U6204 (N_6204,N_4102,N_2867);
nor U6205 (N_6205,N_2798,N_2078);
xor U6206 (N_6206,N_4815,N_660);
xnor U6207 (N_6207,N_3717,N_2494);
xor U6208 (N_6208,N_1041,N_2855);
nor U6209 (N_6209,N_3510,N_4560);
and U6210 (N_6210,N_3866,N_2076);
nor U6211 (N_6211,N_4746,N_2830);
nand U6212 (N_6212,N_4688,N_4666);
nand U6213 (N_6213,N_2583,N_2136);
or U6214 (N_6214,N_21,N_492);
nand U6215 (N_6215,N_2591,N_3281);
nand U6216 (N_6216,N_2325,N_2623);
xnor U6217 (N_6217,N_276,N_1167);
and U6218 (N_6218,N_4193,N_756);
nor U6219 (N_6219,N_103,N_438);
nor U6220 (N_6220,N_4125,N_3961);
and U6221 (N_6221,N_3375,N_343);
nor U6222 (N_6222,N_4937,N_3525);
nand U6223 (N_6223,N_2606,N_2769);
and U6224 (N_6224,N_4679,N_2350);
nor U6225 (N_6225,N_3049,N_1568);
nor U6226 (N_6226,N_1721,N_170);
nand U6227 (N_6227,N_4099,N_4220);
and U6228 (N_6228,N_804,N_953);
nor U6229 (N_6229,N_1020,N_2942);
xnor U6230 (N_6230,N_4313,N_4402);
xor U6231 (N_6231,N_3314,N_3742);
and U6232 (N_6232,N_470,N_540);
and U6233 (N_6233,N_1709,N_3033);
xnor U6234 (N_6234,N_4586,N_3810);
xor U6235 (N_6235,N_4745,N_2312);
xor U6236 (N_6236,N_3546,N_1378);
xnor U6237 (N_6237,N_4206,N_7);
or U6238 (N_6238,N_3461,N_3136);
nor U6239 (N_6239,N_2702,N_4250);
or U6240 (N_6240,N_647,N_856);
xnor U6241 (N_6241,N_174,N_4058);
and U6242 (N_6242,N_3658,N_1245);
or U6243 (N_6243,N_773,N_1976);
nand U6244 (N_6244,N_4319,N_2995);
nor U6245 (N_6245,N_3724,N_1038);
xnor U6246 (N_6246,N_2713,N_1282);
nor U6247 (N_6247,N_2208,N_977);
and U6248 (N_6248,N_2976,N_645);
or U6249 (N_6249,N_2911,N_2608);
nand U6250 (N_6250,N_2815,N_2913);
or U6251 (N_6251,N_3279,N_707);
nand U6252 (N_6252,N_4574,N_636);
and U6253 (N_6253,N_1671,N_670);
xnor U6254 (N_6254,N_2187,N_2295);
nor U6255 (N_6255,N_772,N_136);
nand U6256 (N_6256,N_314,N_1731);
or U6257 (N_6257,N_602,N_3661);
or U6258 (N_6258,N_2395,N_4909);
xnor U6259 (N_6259,N_4848,N_1366);
xnor U6260 (N_6260,N_2287,N_1531);
nor U6261 (N_6261,N_716,N_3989);
and U6262 (N_6262,N_3515,N_948);
xor U6263 (N_6263,N_1485,N_1567);
or U6264 (N_6264,N_1148,N_903);
or U6265 (N_6265,N_3611,N_3623);
nand U6266 (N_6266,N_3925,N_1134);
xor U6267 (N_6267,N_2581,N_4515);
nand U6268 (N_6268,N_2217,N_2225);
nor U6269 (N_6269,N_4282,N_2862);
xor U6270 (N_6270,N_2941,N_651);
or U6271 (N_6271,N_34,N_4805);
nand U6272 (N_6272,N_830,N_2063);
nor U6273 (N_6273,N_1350,N_1878);
xor U6274 (N_6274,N_2314,N_2418);
and U6275 (N_6275,N_4100,N_2705);
nor U6276 (N_6276,N_4366,N_2434);
or U6277 (N_6277,N_3804,N_1468);
or U6278 (N_6278,N_147,N_4996);
nor U6279 (N_6279,N_1083,N_4066);
nand U6280 (N_6280,N_2781,N_2467);
and U6281 (N_6281,N_1085,N_3289);
or U6282 (N_6282,N_111,N_4460);
or U6283 (N_6283,N_4054,N_586);
nand U6284 (N_6284,N_1628,N_4663);
and U6285 (N_6285,N_841,N_4626);
xor U6286 (N_6286,N_3017,N_3535);
xnor U6287 (N_6287,N_1541,N_3640);
nor U6288 (N_6288,N_134,N_2524);
nand U6289 (N_6289,N_83,N_1276);
nand U6290 (N_6290,N_3323,N_4865);
or U6291 (N_6291,N_4595,N_4232);
nor U6292 (N_6292,N_3022,N_457);
nand U6293 (N_6293,N_2579,N_738);
or U6294 (N_6294,N_4519,N_870);
nand U6295 (N_6295,N_3719,N_1729);
or U6296 (N_6296,N_4178,N_720);
nand U6297 (N_6297,N_3965,N_145);
and U6298 (N_6298,N_1977,N_3210);
and U6299 (N_6299,N_2008,N_3502);
nor U6300 (N_6300,N_3098,N_4616);
nor U6301 (N_6301,N_435,N_1441);
nor U6302 (N_6302,N_642,N_3333);
xnor U6303 (N_6303,N_1687,N_2324);
nor U6304 (N_6304,N_687,N_2543);
xnor U6305 (N_6305,N_2930,N_3462);
and U6306 (N_6306,N_1261,N_4265);
xnor U6307 (N_6307,N_1907,N_4809);
xnor U6308 (N_6308,N_138,N_3771);
and U6309 (N_6309,N_4630,N_3258);
or U6310 (N_6310,N_1672,N_3379);
nor U6311 (N_6311,N_9,N_2361);
xor U6312 (N_6312,N_4773,N_2839);
or U6313 (N_6313,N_4044,N_1171);
nand U6314 (N_6314,N_4674,N_1330);
nand U6315 (N_6315,N_4706,N_2254);
or U6316 (N_6316,N_1425,N_3890);
and U6317 (N_6317,N_3189,N_564);
xnor U6318 (N_6318,N_805,N_749);
xor U6319 (N_6319,N_790,N_2406);
nor U6320 (N_6320,N_449,N_4306);
nand U6321 (N_6321,N_3407,N_1249);
and U6322 (N_6322,N_2403,N_2478);
or U6323 (N_6323,N_3399,N_579);
nor U6324 (N_6324,N_3801,N_153);
nor U6325 (N_6325,N_1598,N_2490);
nor U6326 (N_6326,N_4204,N_499);
nor U6327 (N_6327,N_828,N_615);
xor U6328 (N_6328,N_3391,N_432);
nor U6329 (N_6329,N_2386,N_2686);
nor U6330 (N_6330,N_1341,N_1291);
nand U6331 (N_6331,N_4253,N_3267);
nor U6332 (N_6332,N_821,N_761);
nand U6333 (N_6333,N_1823,N_1113);
or U6334 (N_6334,N_2628,N_2154);
nand U6335 (N_6335,N_3595,N_1154);
nand U6336 (N_6336,N_1144,N_3590);
or U6337 (N_6337,N_4183,N_674);
xor U6338 (N_6338,N_3731,N_2471);
xnor U6339 (N_6339,N_3034,N_1351);
or U6340 (N_6340,N_724,N_162);
and U6341 (N_6341,N_955,N_4912);
and U6342 (N_6342,N_2570,N_1107);
or U6343 (N_6343,N_4923,N_3626);
xnor U6344 (N_6344,N_4829,N_814);
nand U6345 (N_6345,N_898,N_2797);
nor U6346 (N_6346,N_566,N_1429);
and U6347 (N_6347,N_4922,N_1342);
or U6348 (N_6348,N_3751,N_2973);
nor U6349 (N_6349,N_1108,N_3074);
xnor U6350 (N_6350,N_2124,N_1702);
or U6351 (N_6351,N_2988,N_4121);
nand U6352 (N_6352,N_1678,N_1832);
nand U6353 (N_6353,N_1204,N_2963);
or U6354 (N_6354,N_4230,N_2843);
nor U6355 (N_6355,N_1837,N_3769);
nor U6356 (N_6356,N_2140,N_4825);
nor U6357 (N_6357,N_3898,N_4510);
nor U6358 (N_6358,N_2880,N_3186);
nor U6359 (N_6359,N_2831,N_4730);
or U6360 (N_6360,N_2220,N_2057);
and U6361 (N_6361,N_1992,N_4694);
xnor U6362 (N_6362,N_1705,N_2304);
xor U6363 (N_6363,N_2500,N_1788);
and U6364 (N_6364,N_2037,N_4199);
or U6365 (N_6365,N_1883,N_2020);
or U6366 (N_6366,N_2538,N_3011);
nor U6367 (N_6367,N_3819,N_4269);
nand U6368 (N_6368,N_2595,N_1859);
xor U6369 (N_6369,N_4118,N_4092);
and U6370 (N_6370,N_3874,N_1834);
nor U6371 (N_6371,N_1313,N_4640);
nor U6372 (N_6372,N_2089,N_2082);
nor U6373 (N_6373,N_4784,N_384);
nand U6374 (N_6374,N_1187,N_1017);
or U6375 (N_6375,N_2364,N_4453);
nand U6376 (N_6376,N_4869,N_4961);
xnor U6377 (N_6377,N_3956,N_3779);
xor U6378 (N_6378,N_4075,N_3066);
nand U6379 (N_6379,N_4910,N_2005);
nand U6380 (N_6380,N_1728,N_3494);
and U6381 (N_6381,N_575,N_1380);
nor U6382 (N_6382,N_2856,N_4213);
and U6383 (N_6383,N_2956,N_4037);
nor U6384 (N_6384,N_4305,N_865);
xnor U6385 (N_6385,N_6,N_1166);
and U6386 (N_6386,N_3842,N_967);
xor U6387 (N_6387,N_755,N_1409);
or U6388 (N_6388,N_3709,N_578);
xor U6389 (N_6389,N_1674,N_864);
or U6390 (N_6390,N_41,N_2821);
nor U6391 (N_6391,N_2824,N_2239);
nor U6392 (N_6392,N_4291,N_3088);
nor U6393 (N_6393,N_1758,N_519);
nand U6394 (N_6394,N_2722,N_2328);
or U6395 (N_6395,N_535,N_1266);
xnor U6396 (N_6396,N_4615,N_1571);
nand U6397 (N_6397,N_4528,N_2228);
nor U6398 (N_6398,N_1165,N_2547);
nor U6399 (N_6399,N_4435,N_213);
nor U6400 (N_6400,N_3543,N_958);
or U6401 (N_6401,N_1751,N_3839);
and U6402 (N_6402,N_4320,N_2817);
nand U6403 (N_6403,N_45,N_801);
xor U6404 (N_6404,N_2696,N_2945);
nand U6405 (N_6405,N_968,N_258);
nor U6406 (N_6406,N_1551,N_2541);
and U6407 (N_6407,N_4445,N_4643);
xor U6408 (N_6408,N_3263,N_2823);
nand U6409 (N_6409,N_2311,N_4375);
nor U6410 (N_6410,N_230,N_4533);
or U6411 (N_6411,N_2553,N_2980);
and U6412 (N_6412,N_1074,N_1689);
or U6413 (N_6413,N_2955,N_2223);
and U6414 (N_6414,N_628,N_688);
or U6415 (N_6415,N_1040,N_1570);
nand U6416 (N_6416,N_372,N_493);
or U6417 (N_6417,N_130,N_2635);
or U6418 (N_6418,N_388,N_3911);
nand U6419 (N_6419,N_989,N_3781);
nor U6420 (N_6420,N_228,N_1021);
xnor U6421 (N_6421,N_1359,N_703);
nor U6422 (N_6422,N_3368,N_3764);
xnor U6423 (N_6423,N_2466,N_1064);
nor U6424 (N_6424,N_1158,N_2846);
nor U6425 (N_6425,N_2678,N_2000);
nand U6426 (N_6426,N_3303,N_4517);
xnor U6427 (N_6427,N_3971,N_1028);
or U6428 (N_6428,N_383,N_3770);
or U6429 (N_6429,N_941,N_662);
nor U6430 (N_6430,N_304,N_4415);
nor U6431 (N_6431,N_3542,N_2297);
xor U6432 (N_6432,N_2097,N_1462);
nand U6433 (N_6433,N_3647,N_3322);
or U6434 (N_6434,N_2667,N_3945);
nor U6435 (N_6435,N_184,N_2890);
xor U6436 (N_6436,N_4194,N_4789);
xor U6437 (N_6437,N_1545,N_2672);
and U6438 (N_6438,N_401,N_1432);
nor U6439 (N_6439,N_1810,N_2523);
nand U6440 (N_6440,N_1719,N_4344);
nand U6441 (N_6441,N_4444,N_1581);
or U6442 (N_6442,N_3010,N_1367);
xnor U6443 (N_6443,N_2928,N_2953);
xor U6444 (N_6444,N_4713,N_2733);
xnor U6445 (N_6445,N_2741,N_523);
nand U6446 (N_6446,N_1338,N_1853);
nor U6447 (N_6447,N_4467,N_3195);
nand U6448 (N_6448,N_3100,N_3472);
and U6449 (N_6449,N_838,N_47);
xor U6450 (N_6450,N_1747,N_2673);
and U6451 (N_6451,N_4378,N_3967);
nor U6452 (N_6452,N_85,N_2047);
nor U6453 (N_6453,N_1267,N_927);
nor U6454 (N_6454,N_4071,N_2476);
nand U6455 (N_6455,N_4043,N_2065);
nor U6456 (N_6456,N_572,N_1466);
nand U6457 (N_6457,N_3409,N_4954);
nor U6458 (N_6458,N_3827,N_762);
nand U6459 (N_6459,N_4360,N_4958);
or U6460 (N_6460,N_1030,N_970);
and U6461 (N_6461,N_1770,N_1517);
xnor U6462 (N_6462,N_507,N_2429);
nor U6463 (N_6463,N_558,N_4354);
nand U6464 (N_6464,N_4828,N_4101);
nor U6465 (N_6465,N_574,N_3505);
xor U6466 (N_6466,N_1679,N_1844);
nor U6467 (N_6467,N_3145,N_1079);
nor U6468 (N_6468,N_4579,N_2138);
nor U6469 (N_6469,N_4782,N_1372);
xor U6470 (N_6470,N_2300,N_3062);
nor U6471 (N_6471,N_280,N_3405);
xor U6472 (N_6472,N_2879,N_2412);
nor U6473 (N_6473,N_4403,N_2046);
xnor U6474 (N_6474,N_1328,N_3115);
and U6475 (N_6475,N_3438,N_4304);
nand U6476 (N_6476,N_3909,N_3182);
xnor U6477 (N_6477,N_526,N_1972);
xnor U6478 (N_6478,N_369,N_2202);
nand U6479 (N_6479,N_2783,N_3894);
or U6480 (N_6480,N_2998,N_2629);
or U6481 (N_6481,N_4155,N_3474);
xnor U6482 (N_6482,N_2925,N_1088);
nor U6483 (N_6483,N_2986,N_2816);
and U6484 (N_6484,N_4836,N_3660);
nand U6485 (N_6485,N_3292,N_352);
or U6486 (N_6486,N_2563,N_1826);
nand U6487 (N_6487,N_1210,N_4286);
and U6488 (N_6488,N_370,N_3101);
nand U6489 (N_6489,N_4577,N_237);
nand U6490 (N_6490,N_3691,N_2756);
nand U6491 (N_6491,N_1180,N_1459);
nor U6492 (N_6492,N_3720,N_1169);
and U6493 (N_6493,N_908,N_4160);
nor U6494 (N_6494,N_3957,N_4389);
nand U6495 (N_6495,N_2624,N_1024);
xor U6496 (N_6496,N_3086,N_300);
xnor U6497 (N_6497,N_4598,N_3383);
nor U6498 (N_6498,N_3480,N_3500);
nor U6499 (N_6499,N_2739,N_1666);
nor U6500 (N_6500,N_2740,N_899);
nand U6501 (N_6501,N_3794,N_448);
nand U6502 (N_6502,N_3013,N_4650);
nand U6503 (N_6503,N_3744,N_4209);
or U6504 (N_6504,N_2653,N_3745);
and U6505 (N_6505,N_105,N_334);
or U6506 (N_6506,N_3007,N_1499);
nor U6507 (N_6507,N_2259,N_3596);
xnor U6508 (N_6508,N_4917,N_2230);
and U6509 (N_6509,N_2596,N_1707);
xor U6510 (N_6510,N_1982,N_263);
nand U6511 (N_6511,N_3251,N_2019);
or U6512 (N_6512,N_3003,N_4601);
and U6513 (N_6513,N_3981,N_4437);
nand U6514 (N_6514,N_345,N_1532);
and U6515 (N_6515,N_1783,N_4859);
or U6516 (N_6516,N_3986,N_4383);
or U6517 (N_6517,N_1857,N_3113);
xnor U6518 (N_6518,N_2115,N_1352);
nand U6519 (N_6519,N_1487,N_1962);
nand U6520 (N_6520,N_3760,N_3116);
nand U6521 (N_6521,N_2062,N_2972);
xor U6522 (N_6522,N_2343,N_2199);
and U6523 (N_6523,N_1575,N_4778);
nand U6524 (N_6524,N_4248,N_1936);
or U6525 (N_6525,N_1481,N_869);
and U6526 (N_6526,N_4412,N_4449);
nor U6527 (N_6527,N_2486,N_4149);
nand U6528 (N_6528,N_3974,N_905);
nor U6529 (N_6529,N_4982,N_322);
nor U6530 (N_6530,N_983,N_124);
nand U6531 (N_6531,N_2514,N_3644);
nor U6532 (N_6532,N_2778,N_4634);
and U6533 (N_6533,N_120,N_4842);
nand U6534 (N_6534,N_4687,N_979);
nand U6535 (N_6535,N_2423,N_3458);
nor U6536 (N_6536,N_4027,N_4174);
or U6537 (N_6537,N_2071,N_1969);
xor U6538 (N_6538,N_4153,N_1333);
nand U6539 (N_6539,N_1177,N_2730);
nand U6540 (N_6540,N_1435,N_1454);
nand U6541 (N_6541,N_1315,N_4989);
or U6542 (N_6542,N_854,N_191);
or U6543 (N_6543,N_2920,N_368);
xor U6544 (N_6544,N_785,N_1514);
nor U6545 (N_6545,N_4186,N_3244);
and U6546 (N_6546,N_1931,N_734);
nand U6547 (N_6547,N_4005,N_3538);
or U6548 (N_6548,N_2106,N_3701);
nand U6549 (N_6549,N_272,N_3679);
nor U6550 (N_6550,N_807,N_1259);
nand U6551 (N_6551,N_2179,N_4143);
nor U6552 (N_6552,N_2450,N_1382);
nand U6553 (N_6553,N_624,N_2749);
xor U6554 (N_6554,N_684,N_4231);
nand U6555 (N_6555,N_152,N_1375);
xnor U6556 (N_6556,N_3106,N_2159);
nand U6557 (N_6557,N_4214,N_2659);
xor U6558 (N_6558,N_3266,N_1940);
or U6559 (N_6559,N_2837,N_472);
and U6560 (N_6560,N_4457,N_4735);
nand U6561 (N_6561,N_189,N_3905);
xor U6562 (N_6562,N_2569,N_3773);
xor U6563 (N_6563,N_911,N_4771);
and U6564 (N_6564,N_751,N_541);
xor U6565 (N_6565,N_2405,N_3798);
and U6566 (N_6566,N_2212,N_4061);
and U6567 (N_6567,N_193,N_1978);
nor U6568 (N_6568,N_290,N_759);
xnor U6569 (N_6569,N_3566,N_411);
nor U6570 (N_6570,N_747,N_3453);
nor U6571 (N_6571,N_4704,N_156);
and U6572 (N_6572,N_1331,N_3848);
nand U6573 (N_6573,N_2272,N_3082);
xnor U6574 (N_6574,N_2776,N_4562);
or U6575 (N_6575,N_2676,N_568);
xor U6576 (N_6576,N_1431,N_2512);
or U6577 (N_6577,N_570,N_3428);
nand U6578 (N_6578,N_271,N_520);
and U6579 (N_6579,N_390,N_2760);
or U6580 (N_6580,N_2795,N_2603);
nand U6581 (N_6581,N_1145,N_3747);
and U6582 (N_6582,N_2617,N_3958);
or U6583 (N_6583,N_1966,N_433);
and U6584 (N_6584,N_2234,N_710);
or U6585 (N_6585,N_831,N_2546);
and U6586 (N_6586,N_1111,N_2080);
xor U6587 (N_6587,N_2803,N_1349);
xnor U6588 (N_6588,N_500,N_3437);
and U6589 (N_6589,N_3809,N_897);
and U6590 (N_6590,N_2660,N_3160);
xor U6591 (N_6591,N_2746,N_879);
nor U6592 (N_6592,N_1473,N_3649);
or U6593 (N_6593,N_2358,N_3324);
nand U6594 (N_6594,N_2533,N_3097);
or U6595 (N_6595,N_2751,N_3963);
nor U6596 (N_6596,N_1769,N_4347);
or U6597 (N_6597,N_4377,N_1724);
and U6598 (N_6598,N_4514,N_4903);
nand U6599 (N_6599,N_2489,N_3565);
and U6600 (N_6600,N_1470,N_4035);
xnor U6601 (N_6601,N_872,N_2727);
nand U6602 (N_6602,N_1168,N_4187);
nor U6603 (N_6603,N_4885,N_4914);
or U6604 (N_6604,N_3953,N_3479);
and U6605 (N_6605,N_2709,N_4711);
and U6606 (N_6606,N_2426,N_2864);
or U6607 (N_6607,N_2582,N_1619);
and U6608 (N_6608,N_1212,N_873);
nand U6609 (N_6609,N_1502,N_2337);
nand U6610 (N_6610,N_2424,N_1067);
nand U6611 (N_6611,N_3634,N_1543);
xor U6612 (N_6612,N_4180,N_2887);
nand U6613 (N_6613,N_361,N_404);
or U6614 (N_6614,N_1063,N_1676);
or U6615 (N_6615,N_1869,N_2150);
or U6616 (N_6616,N_4757,N_4585);
or U6617 (N_6617,N_947,N_3973);
nand U6618 (N_6618,N_139,N_1290);
nor U6619 (N_6619,N_309,N_2638);
or U6620 (N_6620,N_778,N_4082);
nand U6621 (N_6621,N_35,N_3997);
or U6622 (N_6622,N_1556,N_839);
xnor U6623 (N_6623,N_552,N_4897);
xnor U6624 (N_6624,N_3275,N_3635);
nand U6625 (N_6625,N_417,N_1218);
nand U6626 (N_6626,N_1152,N_3403);
xnor U6627 (N_6627,N_1424,N_2960);
nor U6628 (N_6628,N_3899,N_1428);
xnor U6629 (N_6629,N_4184,N_3287);
and U6630 (N_6630,N_517,N_2257);
and U6631 (N_6631,N_3919,N_4491);
xnor U6632 (N_6632,N_56,N_1820);
nand U6633 (N_6633,N_2794,N_2290);
or U6634 (N_6634,N_4896,N_3319);
and U6635 (N_6635,N_1189,N_3600);
nand U6636 (N_6636,N_976,N_30);
and U6637 (N_6637,N_3767,N_4299);
nand U6638 (N_6638,N_1,N_1324);
or U6639 (N_6639,N_4742,N_3586);
and U6640 (N_6640,N_1733,N_2283);
nand U6641 (N_6641,N_389,N_1059);
nor U6642 (N_6642,N_4854,N_2243);
nand U6643 (N_6643,N_527,N_3046);
nand U6644 (N_6644,N_2247,N_107);
or U6645 (N_6645,N_3417,N_3787);
nor U6646 (N_6646,N_327,N_122);
and U6647 (N_6647,N_4287,N_4243);
and U6648 (N_6648,N_209,N_255);
nor U6649 (N_6649,N_1840,N_4695);
xnor U6650 (N_6650,N_4285,N_4907);
xnor U6651 (N_6651,N_633,N_4168);
xor U6652 (N_6652,N_3254,N_4852);
nand U6653 (N_6653,N_712,N_3178);
nor U6654 (N_6654,N_1246,N_2754);
xor U6655 (N_6655,N_2284,N_1235);
xor U6656 (N_6656,N_1658,N_2302);
nor U6657 (N_6657,N_1422,N_1062);
nor U6658 (N_6658,N_3966,N_3412);
or U6659 (N_6659,N_3164,N_4602);
nand U6660 (N_6660,N_3397,N_3274);
or U6661 (N_6661,N_1087,N_1882);
xnor U6662 (N_6662,N_4368,N_1784);
and U6663 (N_6663,N_2703,N_4006);
xor U6664 (N_6664,N_2854,N_2962);
and U6665 (N_6665,N_2226,N_629);
xor U6666 (N_6666,N_2301,N_287);
nand U6667 (N_6667,N_2949,N_2893);
nor U6668 (N_6668,N_1847,N_1434);
and U6669 (N_6669,N_4701,N_4690);
xnor U6670 (N_6670,N_3452,N_1688);
xor U6671 (N_6671,N_3129,N_3673);
nor U6672 (N_6672,N_4525,N_3818);
or U6673 (N_6673,N_3355,N_1241);
or U6674 (N_6674,N_350,N_2644);
nand U6675 (N_6675,N_3059,N_1915);
and U6676 (N_6676,N_2943,N_2834);
or U6677 (N_6677,N_267,N_398);
and U6678 (N_6678,N_2529,N_4161);
nand U6679 (N_6679,N_1696,N_446);
and U6680 (N_6680,N_456,N_1500);
nand U6681 (N_6681,N_3687,N_4266);
or U6682 (N_6682,N_4134,N_1095);
or U6683 (N_6683,N_668,N_279);
and U6684 (N_6684,N_208,N_2996);
nand U6685 (N_6685,N_233,N_454);
or U6686 (N_6686,N_620,N_1973);
xor U6687 (N_6687,N_2487,N_3734);
nand U6688 (N_6688,N_585,N_2452);
nor U6689 (N_6689,N_1765,N_3483);
nor U6690 (N_6690,N_3570,N_4278);
nor U6691 (N_6691,N_4523,N_2345);
nand U6692 (N_6692,N_4793,N_4060);
nand U6693 (N_6693,N_1310,N_587);
nor U6694 (N_6694,N_2253,N_583);
xor U6695 (N_6695,N_1238,N_1252);
nand U6696 (N_6696,N_22,N_1512);
xor U6697 (N_6697,N_4157,N_1805);
nand U6698 (N_6698,N_234,N_4371);
or U6699 (N_6699,N_4892,N_66);
xnor U6700 (N_6700,N_3564,N_3556);
and U6701 (N_6701,N_1121,N_3209);
xor U6702 (N_6702,N_1044,N_2335);
and U6703 (N_6703,N_1140,N_4117);
or U6704 (N_6704,N_3738,N_1295);
and U6705 (N_6705,N_1667,N_959);
and U6706 (N_6706,N_1641,N_713);
and U6707 (N_6707,N_3197,N_1384);
and U6708 (N_6708,N_3551,N_3422);
nand U6709 (N_6709,N_971,N_2369);
or U6710 (N_6710,N_62,N_889);
and U6711 (N_6711,N_1155,N_4387);
nor U6712 (N_6712,N_3419,N_4908);
xnor U6713 (N_6713,N_2011,N_1590);
or U6714 (N_6714,N_4341,N_1901);
and U6715 (N_6715,N_348,N_4438);
nand U6716 (N_6716,N_972,N_3964);
and U6717 (N_6717,N_4289,N_480);
nor U6718 (N_6718,N_4216,N_4755);
nand U6719 (N_6719,N_1303,N_4605);
nor U6720 (N_6720,N_518,N_1483);
xor U6721 (N_6721,N_2326,N_4584);
or U6722 (N_6722,N_3758,N_1909);
and U6723 (N_6723,N_1229,N_1018);
nand U6724 (N_6724,N_1836,N_2927);
or U6725 (N_6725,N_1237,N_599);
and U6726 (N_6726,N_2632,N_2878);
xnor U6727 (N_6727,N_239,N_241);
nand U6728 (N_6728,N_3247,N_2213);
and U6729 (N_6729,N_2250,N_2912);
nor U6730 (N_6730,N_3193,N_4974);
nor U6731 (N_6731,N_201,N_2757);
nand U6732 (N_6732,N_1526,N_93);
and U6733 (N_6733,N_4801,N_1309);
or U6734 (N_6734,N_2991,N_3548);
or U6735 (N_6735,N_641,N_2135);
and U6736 (N_6736,N_3684,N_810);
xnor U6737 (N_6737,N_919,N_1501);
nor U6738 (N_6738,N_4748,N_2576);
nor U6739 (N_6739,N_609,N_3829);
nor U6740 (N_6740,N_264,N_4259);
nor U6741 (N_6741,N_2211,N_1566);
and U6742 (N_6742,N_3523,N_1078);
or U6743 (N_6743,N_4841,N_1855);
or U6744 (N_6744,N_1510,N_4653);
xor U6745 (N_6745,N_3173,N_4839);
nor U6746 (N_6746,N_3035,N_3147);
nor U6747 (N_6747,N_2921,N_1314);
nand U6748 (N_6748,N_3436,N_1037);
nand U6749 (N_6749,N_1998,N_2374);
and U6750 (N_6750,N_3248,N_2789);
nor U6751 (N_6751,N_437,N_188);
or U6752 (N_6752,N_1986,N_1000);
xor U6753 (N_6753,N_657,N_2347);
or U6754 (N_6754,N_4363,N_3790);
xnor U6755 (N_6755,N_1482,N_3698);
nor U6756 (N_6756,N_1287,N_1255);
xor U6757 (N_6757,N_223,N_175);
nand U6758 (N_6758,N_4776,N_346);
nand U6759 (N_6759,N_4864,N_1635);
nor U6760 (N_6760,N_1723,N_3411);
nor U6761 (N_6761,N_1060,N_1789);
nor U6762 (N_6762,N_1743,N_4696);
and U6763 (N_6763,N_634,N_2910);
and U6764 (N_6764,N_2410,N_220);
and U6765 (N_6765,N_597,N_43);
and U6766 (N_6766,N_4133,N_1505);
and U6767 (N_6767,N_2372,N_4894);
or U6768 (N_6768,N_3949,N_4089);
nand U6769 (N_6769,N_3018,N_1926);
or U6770 (N_6770,N_4875,N_2306);
and U6771 (N_6771,N_1100,N_2430);
or U6772 (N_6772,N_1047,N_1196);
or U6773 (N_6773,N_1684,N_1540);
and U6774 (N_6774,N_1727,N_4448);
or U6775 (N_6775,N_453,N_4752);
xor U6776 (N_6776,N_275,N_3877);
and U6777 (N_6777,N_2409,N_2139);
nand U6778 (N_6778,N_2129,N_3433);
nor U6779 (N_6779,N_1214,N_4657);
nand U6780 (N_6780,N_96,N_2508);
or U6781 (N_6781,N_4904,N_2558);
and U6782 (N_6782,N_4943,N_3707);
and U6783 (N_6783,N_1580,N_3232);
nand U6784 (N_6784,N_3401,N_4093);
nor U6785 (N_6785,N_644,N_1766);
nand U6786 (N_6786,N_4014,N_539);
nor U6787 (N_6787,N_630,N_1231);
nor U6788 (N_6788,N_4786,N_4526);
xor U6789 (N_6789,N_909,N_2064);
and U6790 (N_6790,N_1652,N_3508);
xnor U6791 (N_6791,N_2594,N_2950);
nor U6792 (N_6792,N_760,N_3712);
xor U6793 (N_6793,N_3441,N_2085);
or U6794 (N_6794,N_766,N_888);
or U6795 (N_6795,N_4658,N_2933);
or U6796 (N_6796,N_1036,N_2148);
or U6797 (N_6797,N_521,N_3869);
xor U6798 (N_6798,N_200,N_2811);
and U6799 (N_6799,N_2244,N_4988);
nand U6800 (N_6800,N_381,N_89);
and U6801 (N_6801,N_4074,N_4783);
and U6802 (N_6802,N_4572,N_3695);
xnor U6803 (N_6803,N_2661,N_1990);
xor U6804 (N_6804,N_4661,N_1110);
or U6805 (N_6805,N_1622,N_1525);
or U6806 (N_6806,N_1277,N_2203);
nand U6807 (N_6807,N_4281,N_3743);
xor U6808 (N_6808,N_49,N_2559);
nand U6809 (N_6809,N_2540,N_4608);
and U6810 (N_6810,N_2454,N_455);
or U6811 (N_6811,N_1618,N_769);
xor U6812 (N_6812,N_2397,N_3202);
nor U6813 (N_6813,N_2525,N_2763);
xnor U6814 (N_6814,N_621,N_3284);
nand U6815 (N_6815,N_1860,N_2163);
or U6816 (N_6816,N_4942,N_3109);
and U6817 (N_6817,N_378,N_2072);
and U6818 (N_6818,N_4185,N_3384);
nand U6819 (N_6819,N_4816,N_510);
nor U6820 (N_6820,N_1829,N_3571);
and U6821 (N_6821,N_2737,N_1484);
xnor U6822 (N_6822,N_4321,N_4210);
or U6823 (N_6823,N_4461,N_2091);
xnor U6824 (N_6824,N_1527,N_3352);
nor U6825 (N_6825,N_2549,N_4398);
and U6826 (N_6826,N_3341,N_4884);
or U6827 (N_6827,N_3563,N_231);
xnor U6828 (N_6828,N_503,N_4470);
or U6829 (N_6829,N_3445,N_2748);
and U6830 (N_6830,N_2936,N_563);
and U6831 (N_6831,N_4130,N_212);
xor U6832 (N_6832,N_4983,N_4623);
nand U6833 (N_6833,N_2531,N_852);
nor U6834 (N_6834,N_2526,N_2715);
xor U6835 (N_6835,N_2318,N_3155);
nor U6836 (N_6836,N_4176,N_1968);
or U6837 (N_6837,N_2437,N_169);
and U6838 (N_6838,N_2997,N_4395);
nor U6839 (N_6839,N_4818,N_2774);
and U6840 (N_6840,N_3056,N_1411);
nand U6841 (N_6841,N_4401,N_2614);
and U6842 (N_6842,N_3897,N_3490);
or U6843 (N_6843,N_4535,N_4971);
xor U6844 (N_6844,N_2255,N_4420);
nor U6845 (N_6845,N_1772,N_2045);
and U6846 (N_6846,N_4179,N_730);
or U6847 (N_6847,N_4790,N_2068);
nor U6848 (N_6848,N_1227,N_1872);
nor U6849 (N_6849,N_2367,N_4195);
and U6850 (N_6850,N_4272,N_799);
xnor U6851 (N_6851,N_3241,N_1256);
or U6852 (N_6852,N_3969,N_2610);
nor U6853 (N_6853,N_2983,N_4708);
nand U6854 (N_6854,N_1779,N_4451);
xnor U6855 (N_6855,N_2848,N_2813);
nor U6856 (N_6856,N_476,N_868);
nand U6857 (N_6857,N_543,N_3636);
or U6858 (N_6858,N_4399,N_2630);
and U6859 (N_6859,N_1299,N_3334);
nor U6860 (N_6860,N_1922,N_1474);
or U6861 (N_6861,N_1452,N_3014);
nor U6862 (N_6862,N_875,N_901);
nor U6863 (N_6863,N_2227,N_117);
xnor U6864 (N_6864,N_3060,N_780);
and U6865 (N_6865,N_2278,N_3700);
xor U6866 (N_6866,N_1842,N_4673);
nor U6867 (N_6867,N_2275,N_4429);
nor U6868 (N_6868,N_3140,N_658);
xor U6869 (N_6869,N_1151,N_3527);
or U6870 (N_6870,N_596,N_4960);
and U6871 (N_6871,N_2147,N_4221);
xnor U6872 (N_6872,N_3366,N_1673);
or U6873 (N_6873,N_529,N_2447);
nor U6874 (N_6874,N_490,N_1156);
and U6875 (N_6875,N_1655,N_3070);
and U6876 (N_6876,N_3873,N_422);
xnor U6877 (N_6877,N_295,N_4537);
nor U6878 (N_6878,N_1661,N_2054);
nor U6879 (N_6879,N_2373,N_2970);
xor U6880 (N_6880,N_1845,N_4879);
nand U6881 (N_6881,N_3765,N_3791);
and U6882 (N_6882,N_24,N_4935);
and U6883 (N_6883,N_3187,N_1286);
xor U6884 (N_6884,N_3128,N_2105);
nand U6885 (N_6885,N_4724,N_4603);
xor U6886 (N_6886,N_3509,N_4887);
nor U6887 (N_6887,N_1980,N_1741);
and U6888 (N_6888,N_3373,N_4484);
nand U6889 (N_6889,N_1662,N_2801);
or U6890 (N_6890,N_1623,N_4129);
xor U6891 (N_6891,N_4019,N_4844);
or U6892 (N_6892,N_4114,N_151);
or U6893 (N_6893,N_488,N_1715);
and U6894 (N_6894,N_3872,N_1542);
and U6895 (N_6895,N_477,N_1999);
nor U6896 (N_6896,N_1865,N_4853);
xnor U6897 (N_6897,N_459,N_1128);
nor U6898 (N_6898,N_58,N_3429);
nor U6899 (N_6899,N_542,N_3752);
and U6900 (N_6900,N_3845,N_3347);
xnor U6901 (N_6901,N_1394,N_689);
and U6902 (N_6902,N_0,N_2732);
or U6903 (N_6903,N_3199,N_323);
nor U6904 (N_6904,N_2866,N_379);
nand U6905 (N_6905,N_961,N_2918);
nand U6906 (N_6906,N_4262,N_3993);
nor U6907 (N_6907,N_3430,N_1524);
nor U6908 (N_6908,N_3,N_705);
and U6909 (N_6909,N_4487,N_1813);
or U6910 (N_6910,N_883,N_4056);
nand U6911 (N_6911,N_2496,N_3159);
and U6912 (N_6912,N_131,N_2053);
or U6913 (N_6913,N_4891,N_407);
and U6914 (N_6914,N_4539,N_556);
and U6915 (N_6915,N_3378,N_4830);
xor U6916 (N_6916,N_882,N_3662);
xor U6917 (N_6917,N_157,N_1550);
nand U6918 (N_6918,N_3507,N_607);
nor U6919 (N_6919,N_1749,N_3868);
xor U6920 (N_6920,N_3977,N_2598);
xor U6921 (N_6921,N_3972,N_3727);
nand U6922 (N_6922,N_1675,N_4516);
or U6923 (N_6923,N_2932,N_4668);
nor U6924 (N_6924,N_719,N_4373);
nor U6925 (N_6925,N_3335,N_2121);
nand U6926 (N_6926,N_2237,N_1830);
or U6927 (N_6927,N_4396,N_4900);
nor U6928 (N_6928,N_1819,N_2840);
nand U6929 (N_6929,N_4753,N_950);
and U6930 (N_6930,N_3282,N_1991);
and U6931 (N_6931,N_1816,N_3253);
or U6932 (N_6932,N_2167,N_894);
and U6933 (N_6933,N_553,N_1469);
nand U6934 (N_6934,N_4955,N_168);
nor U6935 (N_6935,N_3200,N_4227);
nor U6936 (N_6936,N_3340,N_3206);
and U6937 (N_6937,N_3677,N_2132);
xor U6938 (N_6938,N_3095,N_1924);
nand U6939 (N_6939,N_1790,N_2083);
and U6940 (N_6940,N_3107,N_3444);
or U6941 (N_6941,N_284,N_2604);
or U6942 (N_6942,N_204,N_1544);
xnor U6943 (N_6943,N_770,N_4426);
or U6944 (N_6944,N_31,N_3089);
nor U6945 (N_6945,N_3936,N_1388);
or U6946 (N_6946,N_2901,N_1076);
xnor U6947 (N_6947,N_1706,N_994);
or U6948 (N_6948,N_1507,N_2922);
and U6949 (N_6949,N_739,N_2378);
and U6950 (N_6950,N_2564,N_2677);
and U6951 (N_6951,N_3299,N_1867);
xnor U6952 (N_6952,N_937,N_4867);
nor U6953 (N_6953,N_447,N_1630);
nand U6954 (N_6954,N_473,N_4948);
or U6955 (N_6955,N_2861,N_2185);
and U6956 (N_6956,N_3853,N_2131);
nor U6957 (N_6957,N_4026,N_464);
nor U6958 (N_6958,N_1718,N_2455);
and U6959 (N_6959,N_3830,N_2029);
xnor U6960 (N_6960,N_393,N_4165);
nor U6961 (N_6961,N_2761,N_1881);
and U6962 (N_6962,N_2584,N_2142);
xnor U6963 (N_6963,N_3158,N_1077);
and U6964 (N_6964,N_461,N_1174);
nand U6965 (N_6965,N_1620,N_4481);
xor U6966 (N_6966,N_2177,N_57);
nand U6967 (N_6967,N_2266,N_2155);
nand U6968 (N_6968,N_4750,N_3714);
or U6969 (N_6969,N_3123,N_1736);
nand U6970 (N_6970,N_4057,N_4986);
nor U6971 (N_6971,N_4823,N_1781);
nand U6972 (N_6972,N_3169,N_3133);
nor U6973 (N_6973,N_1752,N_1311);
xnor U6974 (N_6974,N_1183,N_3668);
and U6975 (N_6975,N_4625,N_2415);
xor U6976 (N_6976,N_4175,N_3530);
nand U6977 (N_6977,N_3052,N_1164);
or U6978 (N_6978,N_180,N_1963);
xnor U6979 (N_6979,N_359,N_4488);
nand U6980 (N_6980,N_842,N_158);
xnor U6981 (N_6981,N_627,N_414);
nor U6982 (N_6982,N_4496,N_567);
or U6983 (N_6983,N_2114,N_4628);
and U6984 (N_6984,N_1851,N_999);
and U6985 (N_6985,N_226,N_4098);
or U6986 (N_6986,N_4785,N_2200);
or U6987 (N_6987,N_198,N_505);
xnor U6988 (N_6988,N_4962,N_1997);
or U6989 (N_6989,N_679,N_1876);
or U6990 (N_6990,N_548,N_4749);
nand U6991 (N_6991,N_4392,N_3380);
and U6992 (N_6992,N_1536,N_4703);
or U6993 (N_6993,N_247,N_487);
and U6994 (N_6994,N_2368,N_3795);
xor U6995 (N_6995,N_132,N_4868);
or U6996 (N_6996,N_779,N_1012);
and U6997 (N_6997,N_3574,N_2329);
nor U6998 (N_6998,N_3201,N_95);
and U6999 (N_6999,N_4370,N_1546);
nor U7000 (N_7000,N_296,N_2161);
nand U7001 (N_7001,N_2176,N_4648);
xor U7002 (N_7002,N_2951,N_4812);
nor U7003 (N_7003,N_4929,N_14);
xor U7004 (N_7004,N_2958,N_15);
nor U7005 (N_7005,N_4810,N_2773);
and U7006 (N_7006,N_1574,N_610);
nor U7007 (N_7007,N_2978,N_3806);
nand U7008 (N_7008,N_3871,N_1203);
nand U7009 (N_7009,N_1011,N_768);
xor U7010 (N_7010,N_2059,N_3789);
nor U7011 (N_7011,N_3629,N_4646);
xnor U7012 (N_7012,N_1592,N_1565);
or U7013 (N_7013,N_1260,N_3058);
nor U7014 (N_7014,N_502,N_4522);
nor U7015 (N_7015,N_3047,N_2616);
nor U7016 (N_7016,N_1824,N_1361);
and U7017 (N_7017,N_3834,N_1744);
xnor U7018 (N_7018,N_1646,N_3552);
nand U7019 (N_7019,N_4565,N_3587);
nand U7020 (N_7020,N_3910,N_1336);
xnor U7021 (N_7021,N_2398,N_1950);
nand U7022 (N_7022,N_4173,N_2729);
nand U7023 (N_7023,N_409,N_3882);
and U7024 (N_7024,N_2567,N_3415);
nand U7025 (N_7025,N_4256,N_1712);
nand U7026 (N_7026,N_3918,N_4407);
nand U7027 (N_7027,N_672,N_4069);
nor U7028 (N_7028,N_3864,N_3887);
or U7029 (N_7029,N_2339,N_2907);
and U7030 (N_7030,N_4374,N_1457);
xnor U7031 (N_7031,N_2961,N_4849);
and U7032 (N_7032,N_2344,N_1407);
xnor U7033 (N_7033,N_1558,N_1495);
xnor U7034 (N_7034,N_2070,N_1602);
or U7035 (N_7035,N_316,N_3476);
and U7036 (N_7036,N_3489,N_771);
or U7037 (N_7037,N_242,N_776);
nand U7038 (N_7038,N_508,N_4548);
nand U7039 (N_7039,N_1827,N_1763);
xnor U7040 (N_7040,N_966,N_3294);
nor U7041 (N_7041,N_2096,N_3555);
nor U7042 (N_7042,N_3608,N_4225);
nand U7043 (N_7043,N_1377,N_1191);
and U7044 (N_7044,N_3068,N_913);
or U7045 (N_7045,N_2036,N_160);
and U7046 (N_7046,N_2073,N_1039);
nor U7047 (N_7047,N_3704,N_4229);
nand U7048 (N_7048,N_374,N_1308);
xor U7049 (N_7049,N_2965,N_4596);
xor U7050 (N_7050,N_2323,N_1414);
xor U7051 (N_7051,N_2193,N_3968);
xor U7052 (N_7052,N_4965,N_1317);
nand U7053 (N_7053,N_2340,N_2162);
or U7054 (N_7054,N_2863,N_1683);
nor U7055 (N_7055,N_4678,N_51);
nor U7056 (N_7056,N_1356,N_3513);
and U7057 (N_7057,N_1649,N_3301);
nand U7058 (N_7058,N_2365,N_274);
nor U7059 (N_7059,N_269,N_675);
nor U7060 (N_7060,N_4095,N_1175);
and U7061 (N_7061,N_3259,N_2157);
or U7062 (N_7062,N_3268,N_3976);
nand U7063 (N_7063,N_2939,N_3723);
and U7064 (N_7064,N_261,N_1994);
and U7065 (N_7065,N_451,N_1737);
or U7066 (N_7066,N_3577,N_3955);
or U7067 (N_7067,N_1082,N_3504);
xor U7068 (N_7068,N_2376,N_3694);
nand U7069 (N_7069,N_1538,N_3511);
xor U7070 (N_7070,N_1547,N_1015);
nor U7071 (N_7071,N_2626,N_603);
and U7072 (N_7072,N_354,N_3083);
or U7073 (N_7073,N_1768,N_3276);
and U7074 (N_7074,N_1353,N_3118);
nor U7075 (N_7075,N_3309,N_4284);
or U7076 (N_7076,N_581,N_2718);
xnor U7077 (N_7077,N_3278,N_3467);
or U7078 (N_7078,N_1120,N_4824);
or U7079 (N_7079,N_3602,N_3310);
xor U7080 (N_7080,N_1561,N_1419);
nand U7081 (N_7081,N_3711,N_99);
nand U7082 (N_7082,N_2173,N_3290);
nand U7083 (N_7083,N_1123,N_80);
nor U7084 (N_7084,N_1284,N_2935);
nand U7085 (N_7085,N_3908,N_1073);
nand U7086 (N_7086,N_923,N_974);
nor U7087 (N_7087,N_3085,N_4787);
nor U7088 (N_7088,N_4576,N_3027);
nor U7089 (N_7089,N_3645,N_4136);
and U7090 (N_7090,N_3249,N_3933);
nand U7091 (N_7091,N_2700,N_695);
or U7092 (N_7092,N_1762,N_3929);
xor U7093 (N_7093,N_1014,N_2622);
and U7094 (N_7094,N_1455,N_1877);
xnor U7095 (N_7095,N_4720,N_4905);
xnor U7096 (N_7096,N_3456,N_4999);
xor U7097 (N_7097,N_4318,N_1894);
nand U7098 (N_7098,N_3582,N_1828);
nor U7099 (N_7099,N_3063,N_1325);
nor U7100 (N_7100,N_1437,N_3231);
and U7101 (N_7101,N_2497,N_2474);
nor U7102 (N_7102,N_4911,N_4609);
nand U7103 (N_7103,N_2964,N_4655);
or U7104 (N_7104,N_183,N_4583);
xor U7105 (N_7105,N_697,N_1563);
nor U7106 (N_7106,N_182,N_931);
xor U7107 (N_7107,N_1379,N_4970);
nor U7108 (N_7108,N_1091,N_3998);
xor U7109 (N_7109,N_1626,N_742);
nor U7110 (N_7110,N_3867,N_788);
or U7111 (N_7111,N_2552,N_2516);
xor U7112 (N_7112,N_557,N_2286);
and U7113 (N_7113,N_2308,N_4631);
nand U7114 (N_7114,N_4930,N_1130);
and U7115 (N_7115,N_3080,N_1119);
and U7116 (N_7116,N_1996,N_1092);
or U7117 (N_7117,N_1143,N_997);
or U7118 (N_7118,N_3125,N_2900);
nand U7119 (N_7119,N_3766,N_2164);
and U7120 (N_7120,N_981,N_709);
xor U7121 (N_7121,N_3881,N_592);
nor U7122 (N_7122,N_2319,N_1606);
or U7123 (N_7123,N_229,N_2112);
and U7124 (N_7124,N_3174,N_4792);
nand U7125 (N_7125,N_1406,N_2331);
xor U7126 (N_7126,N_722,N_3175);
and U7127 (N_7127,N_2081,N_3812);
nand U7128 (N_7128,N_560,N_1491);
nor U7129 (N_7129,N_3914,N_3927);
or U7130 (N_7130,N_1613,N_2520);
or U7131 (N_7131,N_221,N_3358);
nor U7132 (N_7132,N_3318,N_3938);
or U7133 (N_7133,N_2689,N_1583);
or U7134 (N_7134,N_2851,N_4247);
nand U7135 (N_7135,N_3607,N_2589);
nor U7136 (N_7136,N_3652,N_4685);
nand U7137 (N_7137,N_4561,N_4918);
or U7138 (N_7138,N_2790,N_3473);
nor U7139 (N_7139,N_3619,N_292);
nor U7140 (N_7140,N_1722,N_4087);
xor U7141 (N_7141,N_2896,N_4568);
and U7142 (N_7142,N_2108,N_442);
and U7143 (N_7143,N_2320,N_1162);
or U7144 (N_7144,N_632,N_4506);
nor U7145 (N_7145,N_1930,N_143);
nand U7146 (N_7146,N_4761,N_1206);
or U7147 (N_7147,N_4032,N_2420);
nor U7148 (N_7148,N_2427,N_1553);
nor U7149 (N_7149,N_2499,N_1026);
or U7150 (N_7150,N_1433,N_177);
xor U7151 (N_7151,N_861,N_425);
or U7152 (N_7152,N_3498,N_3935);
or U7153 (N_7153,N_4177,N_910);
and U7154 (N_7154,N_4419,N_2770);
and U7155 (N_7155,N_3824,N_1608);
or U7156 (N_7156,N_251,N_949);
nand U7157 (N_7157,N_2745,N_1970);
and U7158 (N_7158,N_812,N_2166);
or U7159 (N_7159,N_1913,N_3617);
nand U7160 (N_7160,N_3185,N_2647);
nor U7161 (N_7161,N_973,N_2214);
nand U7162 (N_7162,N_332,N_4464);
nand U7163 (N_7163,N_2643,N_445);
and U7164 (N_7164,N_3653,N_1879);
and U7165 (N_7165,N_4088,N_654);
or U7166 (N_7166,N_4802,N_3630);
or U7167 (N_7167,N_2292,N_816);
nand U7168 (N_7168,N_4651,N_4369);
nand U7169 (N_7169,N_4851,N_4166);
nor U7170 (N_7170,N_835,N_4331);
and U7171 (N_7171,N_1534,N_2902);
nand U7172 (N_7172,N_4140,N_1208);
and U7173 (N_7173,N_754,N_2793);
nor U7174 (N_7174,N_2401,N_1644);
nor U7175 (N_7175,N_1222,N_2289);
nor U7176 (N_7176,N_4493,N_3572);
and U7177 (N_7177,N_3916,N_2931);
nand U7178 (N_7178,N_4611,N_2613);
nand U7179 (N_7179,N_1929,N_2903);
or U7180 (N_7180,N_4404,N_631);
and U7181 (N_7181,N_3589,N_3293);
or U7182 (N_7182,N_2469,N_1296);
nand U7183 (N_7183,N_2178,N_4878);
xor U7184 (N_7184,N_813,N_1371);
or U7185 (N_7185,N_3757,N_3350);
xnor U7186 (N_7186,N_4224,N_26);
xor U7187 (N_7187,N_2835,N_102);
nand U7188 (N_7188,N_4425,N_3316);
nor U7189 (N_7189,N_2504,N_2615);
or U7190 (N_7190,N_3878,N_4555);
and U7191 (N_7191,N_1387,N_2534);
xnor U7192 (N_7192,N_436,N_623);
xor U7193 (N_7193,N_206,N_549);
and U7194 (N_7194,N_4297,N_729);
or U7195 (N_7195,N_1472,N_4963);
or U7196 (N_7196,N_40,N_1293);
or U7197 (N_7197,N_4011,N_1027);
nand U7198 (N_7198,N_605,N_676);
or U7199 (N_7199,N_2231,N_4769);
xnor U7200 (N_7200,N_4743,N_3312);
nor U7201 (N_7201,N_3091,N_3620);
nor U7202 (N_7202,N_4228,N_2443);
nor U7203 (N_7203,N_577,N_2248);
nand U7204 (N_7204,N_4447,N_3808);
nor U7205 (N_7205,N_3349,N_3856);
nand U7206 (N_7206,N_2058,N_2852);
xor U7207 (N_7207,N_2882,N_686);
nor U7208 (N_7208,N_2895,N_594);
nor U7209 (N_7209,N_1364,N_3692);
xnor U7210 (N_7210,N_522,N_2174);
or U7211 (N_7211,N_2742,N_1554);
or U7212 (N_7212,N_318,N_1668);
xor U7213 (N_7213,N_4915,N_914);
nand U7214 (N_7214,N_4691,N_849);
nor U7215 (N_7215,N_4593,N_2322);
nor U7216 (N_7216,N_2027,N_1217);
nor U7217 (N_7217,N_4542,N_4223);
and U7218 (N_7218,N_2196,N_1831);
xnor U7219 (N_7219,N_1307,N_355);
xnor U7220 (N_7220,N_2417,N_2404);
xnor U7221 (N_7221,N_1700,N_3755);
nand U7222 (N_7222,N_4763,N_4781);
xnor U7223 (N_7223,N_3547,N_1841);
nor U7224 (N_7224,N_3654,N_3828);
and U7225 (N_7225,N_866,N_1004);
xnor U7226 (N_7226,N_4350,N_3718);
xnor U7227 (N_7227,N_439,N_4120);
and U7228 (N_7228,N_1263,N_664);
nand U7229 (N_7229,N_3947,N_3269);
nor U7230 (N_7230,N_2181,N_81);
or U7231 (N_7231,N_335,N_3332);
and U7232 (N_7232,N_1043,N_2889);
xnor U7233 (N_7233,N_1272,N_4620);
nand U7234 (N_7234,N_836,N_4012);
nor U7235 (N_7235,N_4094,N_1332);
nand U7236 (N_7236,N_715,N_3805);
xor U7237 (N_7237,N_2449,N_4683);
and U7238 (N_7238,N_3492,N_3387);
and U7239 (N_7239,N_1983,N_1346);
xnor U7240 (N_7240,N_3271,N_2137);
nor U7241 (N_7241,N_4123,N_4280);
nand U7242 (N_7242,N_1449,N_758);
xnor U7243 (N_7243,N_3273,N_4335);
or U7244 (N_7244,N_2238,N_3722);
xor U7245 (N_7245,N_859,N_3706);
xor U7246 (N_7246,N_2657,N_653);
and U7247 (N_7247,N_3481,N_3130);
nor U7248 (N_7248,N_4271,N_3012);
or U7249 (N_7249,N_3144,N_3330);
nand U7250 (N_7250,N_3950,N_3783);
or U7251 (N_7251,N_4505,N_1670);
or U7252 (N_7252,N_1270,N_347);
and U7253 (N_7253,N_4758,N_3280);
nand U7254 (N_7254,N_3165,N_1726);
or U7255 (N_7255,N_4511,N_1822);
nor U7256 (N_7256,N_2535,N_1771);
and U7257 (N_7257,N_1614,N_2128);
or U7258 (N_7258,N_2451,N_216);
or U7259 (N_7259,N_4856,N_3359);
and U7260 (N_7260,N_750,N_1207);
xor U7261 (N_7261,N_128,N_963);
and U7262 (N_7262,N_1944,N_3521);
or U7263 (N_7263,N_614,N_2251);
and U7264 (N_7264,N_2267,N_3970);
or U7265 (N_7265,N_4045,N_4096);
xnor U7266 (N_7266,N_4182,N_32);
or U7267 (N_7267,N_2542,N_3638);
nand U7268 (N_7268,N_3889,N_1318);
nor U7269 (N_7269,N_4311,N_4051);
or U7270 (N_7270,N_4814,N_2006);
or U7271 (N_7271,N_3328,N_3485);
nor U7272 (N_7272,N_832,N_341);
xor U7273 (N_7273,N_2646,N_1802);
xnor U7274 (N_7274,N_1135,N_532);
nor U7275 (N_7275,N_4821,N_3124);
or U7276 (N_7276,N_3321,N_1594);
and U7277 (N_7277,N_1493,N_3464);
nor U7278 (N_7278,N_3875,N_2764);
nor U7279 (N_7279,N_4739,N_478);
and U7280 (N_7280,N_2521,N_1513);
and U7281 (N_7281,N_896,N_4741);
or U7282 (N_7282,N_4780,N_3191);
nand U7283 (N_7283,N_933,N_4717);
or U7284 (N_7284,N_312,N_4159);
or U7285 (N_7285,N_2459,N_685);
xor U7286 (N_7286,N_2899,N_1537);
or U7287 (N_7287,N_1680,N_273);
xor U7288 (N_7288,N_1858,N_3272);
nor U7289 (N_7289,N_4916,N_2441);
nand U7290 (N_7290,N_3455,N_2640);
nor U7291 (N_7291,N_4150,N_2381);
nand U7292 (N_7292,N_2180,N_4385);
nand U7293 (N_7293,N_303,N_3690);
or U7294 (N_7294,N_4312,N_3214);
xor U7295 (N_7295,N_2380,N_135);
nor U7296 (N_7296,N_4393,N_2122);
nand U7297 (N_7297,N_4302,N_4940);
or U7298 (N_7298,N_3381,N_2031);
and U7299 (N_7299,N_2885,N_3337);
xor U7300 (N_7300,N_4021,N_1801);
nand U7301 (N_7301,N_2691,N_3943);
and U7302 (N_7302,N_2336,N_1489);
and U7303 (N_7303,N_3802,N_2999);
or U7304 (N_7304,N_2874,N_2342);
and U7305 (N_7305,N_4431,N_1942);
and U7306 (N_7306,N_1923,N_3392);
xor U7307 (N_7307,N_2207,N_1179);
or U7308 (N_7308,N_2805,N_324);
xnor U7309 (N_7309,N_4618,N_4883);
xor U7310 (N_7310,N_846,N_484);
and U7311 (N_7311,N_1281,N_1508);
xnor U7312 (N_7312,N_2859,N_1604);
nand U7313 (N_7313,N_3883,N_1300);
xnor U7314 (N_7314,N_2391,N_4332);
nand U7315 (N_7315,N_460,N_2845);
nand U7316 (N_7316,N_4002,N_4774);
and U7317 (N_7317,N_2934,N_2184);
nand U7318 (N_7318,N_794,N_4325);
and U7319 (N_7319,N_1285,N_985);
and U7320 (N_7320,N_516,N_4807);
or U7321 (N_7321,N_2421,N_1103);
xnor U7322 (N_7322,N_2416,N_1745);
xor U7323 (N_7323,N_1932,N_2222);
or U7324 (N_7324,N_1958,N_2038);
and U7325 (N_7325,N_4081,N_1916);
nand U7326 (N_7326,N_3633,N_4985);
nand U7327 (N_7327,N_4009,N_1453);
nand U7328 (N_7328,N_4676,N_1782);
nand U7329 (N_7329,N_1436,N_2366);
xor U7330 (N_7330,N_1494,N_4862);
or U7331 (N_7331,N_3775,N_2886);
nor U7332 (N_7332,N_2827,N_2201);
nor U7333 (N_7333,N_4207,N_1595);
or U7334 (N_7334,N_2731,N_4422);
nand U7335 (N_7335,N_3171,N_4126);
xor U7336 (N_7336,N_848,N_2425);
xnor U7337 (N_7337,N_1735,N_2263);
and U7338 (N_7338,N_3295,N_3370);
nand U7339 (N_7339,N_3568,N_4508);
xnor U7340 (N_7340,N_4693,N_2618);
nand U7341 (N_7341,N_2116,N_1257);
nor U7342 (N_7342,N_214,N_1055);
and U7343 (N_7343,N_3307,N_2952);
xor U7344 (N_7344,N_3803,N_2850);
nand U7345 (N_7345,N_4234,N_1693);
nor U7346 (N_7346,N_3688,N_1780);
nand U7347 (N_7347,N_3015,N_2807);
and U7348 (N_7348,N_1504,N_176);
xnor U7349 (N_7349,N_3061,N_3002);
and U7350 (N_7350,N_1408,N_3385);
nand U7351 (N_7351,N_71,N_1791);
nor U7352 (N_7352,N_3750,N_286);
or U7353 (N_7353,N_1985,N_1677);
and U7354 (N_7354,N_8,N_3365);
xor U7355 (N_7355,N_76,N_3831);
nor U7356 (N_7356,N_4025,N_3796);
nor U7357 (N_7357,N_3374,N_3475);
and U7358 (N_7358,N_4737,N_4681);
nor U7359 (N_7359,N_4873,N_430);
and U7360 (N_7360,N_1584,N_4800);
nor U7361 (N_7361,N_3150,N_17);
and U7362 (N_7362,N_1856,N_3207);
or U7363 (N_7363,N_4105,N_1935);
xnor U7364 (N_7364,N_4442,N_2883);
nor U7365 (N_7365,N_1555,N_2075);
xor U7366 (N_7366,N_3561,N_3041);
nand U7367 (N_7367,N_2261,N_2092);
xnor U7368 (N_7368,N_3156,N_3667);
xnor U7369 (N_7369,N_2407,N_1961);
and U7370 (N_7370,N_4639,N_219);
or U7371 (N_7371,N_2393,N_3470);
xor U7372 (N_7372,N_982,N_2444);
xnor U7373 (N_7373,N_2484,N_793);
nor U7374 (N_7374,N_1523,N_1895);
or U7375 (N_7375,N_1009,N_2502);
nor U7376 (N_7376,N_3471,N_2249);
nand U7377 (N_7377,N_2994,N_2355);
xnor U7378 (N_7378,N_4610,N_885);
xnor U7379 (N_7379,N_802,N_4822);
nand U7380 (N_7380,N_1137,N_3912);
nor U7381 (N_7381,N_3044,N_1355);
nand U7382 (N_7382,N_1686,N_2820);
xor U7383 (N_7383,N_2321,N_3788);
xor U7384 (N_7384,N_1699,N_1634);
xnor U7385 (N_7385,N_4119,N_2090);
or U7386 (N_7386,N_3879,N_2501);
xnor U7387 (N_7387,N_4430,N_2877);
and U7388 (N_7388,N_2600,N_1149);
nor U7389 (N_7389,N_2937,N_4540);
and U7390 (N_7390,N_2522,N_1126);
nand U7391 (N_7391,N_3183,N_118);
nor U7392 (N_7392,N_4564,N_4846);
or U7393 (N_7393,N_536,N_3291);
or U7394 (N_7394,N_2726,N_789);
nand U7395 (N_7395,N_3782,N_837);
nand U7396 (N_7396,N_88,N_421);
xor U7397 (N_7397,N_2652,N_1694);
or U7398 (N_7398,N_3628,N_2545);
or U7399 (N_7399,N_4956,N_3499);
or U7400 (N_7400,N_666,N_978);
xnor U7401 (N_7401,N_545,N_225);
nand U7402 (N_7402,N_3154,N_1582);
nand U7403 (N_7403,N_2519,N_3580);
xor U7404 (N_7404,N_1275,N_4654);
nand U7405 (N_7405,N_4198,N_3642);
xor U7406 (N_7406,N_4276,N_4898);
or U7407 (N_7407,N_4205,N_1057);
nand U7408 (N_7408,N_4145,N_840);
nor U7409 (N_7409,N_580,N_1650);
or U7410 (N_7410,N_2605,N_4946);
and U7411 (N_7411,N_3354,N_4667);
or U7412 (N_7412,N_646,N_2674);
or U7413 (N_7413,N_1995,N_4524);
or U7414 (N_7414,N_3876,N_4494);
nor U7415 (N_7415,N_506,N_3051);
nor U7416 (N_7416,N_339,N_2791);
nand U7417 (N_7417,N_727,N_1654);
and U7418 (N_7418,N_2191,N_3682);
or U7419 (N_7419,N_1242,N_741);
xor U7420 (N_7420,N_127,N_4479);
xnor U7421 (N_7421,N_3454,N_3238);
or U7422 (N_7422,N_3721,N_1496);
nor U7423 (N_7423,N_4733,N_1430);
xnor U7424 (N_7424,N_4443,N_690);
xor U7425 (N_7425,N_3843,N_3439);
or U7426 (N_7426,N_3865,N_2954);
nor U7427 (N_7427,N_262,N_4794);
or U7428 (N_7428,N_3729,N_1034);
xor U7429 (N_7429,N_1316,N_4162);
or U7430 (N_7430,N_800,N_1058);
nand U7431 (N_7431,N_2915,N_4022);
and U7432 (N_7432,N_2224,N_4122);
nor U7433 (N_7433,N_4338,N_3817);
nor U7434 (N_7434,N_4992,N_942);
or U7435 (N_7435,N_4559,N_1312);
and U7436 (N_7436,N_3217,N_3606);
and U7437 (N_7437,N_150,N_3558);
and U7438 (N_7438,N_3421,N_4279);
xnor U7439 (N_7439,N_1348,N_4010);
nor U7440 (N_7440,N_2800,N_3880);
and U7441 (N_7441,N_2565,N_1954);
or U7442 (N_7442,N_4738,N_4662);
nor U7443 (N_7443,N_590,N_1804);
or U7444 (N_7444,N_1131,N_834);
nand U7445 (N_7445,N_301,N_3693);
xor U7446 (N_7446,N_3449,N_3838);
or U7447 (N_7447,N_3954,N_2043);
or U7448 (N_7448,N_2095,N_3618);
nand U7449 (N_7449,N_2262,N_2762);
nor U7450 (N_7450,N_4863,N_1192);
nor U7451 (N_7451,N_2141,N_3728);
xnor U7452 (N_7452,N_3302,N_121);
nand U7453 (N_7453,N_2929,N_1925);
xor U7454 (N_7454,N_2853,N_2079);
nor U7455 (N_7455,N_4267,N_2990);
nor U7456 (N_7456,N_2704,N_1031);
xnor U7457 (N_7457,N_4498,N_4659);
nand U7458 (N_7458,N_3228,N_1186);
or U7459 (N_7459,N_2205,N_2975);
or U7460 (N_7460,N_2633,N_2679);
and U7461 (N_7461,N_867,N_2697);
and U7462 (N_7462,N_3604,N_1887);
or U7463 (N_7463,N_4715,N_2587);
nor U7464 (N_7464,N_2503,N_3084);
nand U7465 (N_7465,N_2044,N_52);
and U7466 (N_7466,N_4534,N_1199);
and U7467 (N_7467,N_4365,N_2050);
xnor U7468 (N_7468,N_2158,N_2898);
and U7469 (N_7469,N_4475,N_3995);
and U7470 (N_7470,N_795,N_282);
nor U7471 (N_7471,N_4439,N_2872);
xor U7472 (N_7472,N_1129,N_4504);
nor U7473 (N_7473,N_915,N_774);
nor U7474 (N_7474,N_4292,N_4707);
and U7475 (N_7475,N_2977,N_3800);
xnor U7476 (N_7476,N_2189,N_217);
and U7477 (N_7477,N_3776,N_1890);
or U7478 (N_7478,N_2,N_353);
xnor U7479 (N_7479,N_4592,N_616);
or U7480 (N_7480,N_1117,N_1178);
and U7481 (N_7481,N_714,N_4729);
nor U7482 (N_7482,N_3057,N_681);
xor U7483 (N_7483,N_1933,N_4597);
and U7484 (N_7484,N_4744,N_1066);
nand U7485 (N_7485,N_1774,N_2752);
or U7486 (N_7486,N_2015,N_4208);
or U7487 (N_7487,N_1868,N_3442);
and U7488 (N_7488,N_4669,N_3836);
nor U7489 (N_7489,N_2888,N_2066);
and U7490 (N_7490,N_1605,N_4169);
or U7491 (N_7491,N_737,N_1796);
and U7492 (N_7492,N_4455,N_1519);
and U7493 (N_7493,N_4261,N_2873);
and U7494 (N_7494,N_1122,N_4612);
nand U7495 (N_7495,N_4482,N_1927);
xor U7496 (N_7496,N_2483,N_4951);
and U7497 (N_7497,N_2759,N_3772);
and U7498 (N_7498,N_4924,N_349);
nand U7499 (N_7499,N_4080,N_1278);
or U7500 (N_7500,N_2633,N_4518);
nand U7501 (N_7501,N_2465,N_4170);
nand U7502 (N_7502,N_1737,N_4133);
nand U7503 (N_7503,N_4679,N_248);
or U7504 (N_7504,N_1821,N_3353);
or U7505 (N_7505,N_2330,N_1534);
nor U7506 (N_7506,N_3430,N_1983);
nand U7507 (N_7507,N_1280,N_3703);
xnor U7508 (N_7508,N_1732,N_1005);
nor U7509 (N_7509,N_2837,N_348);
nor U7510 (N_7510,N_4262,N_3478);
xnor U7511 (N_7511,N_3210,N_1637);
nor U7512 (N_7512,N_4472,N_530);
and U7513 (N_7513,N_2024,N_4496);
nor U7514 (N_7514,N_315,N_909);
xor U7515 (N_7515,N_3988,N_4202);
and U7516 (N_7516,N_4315,N_410);
and U7517 (N_7517,N_1832,N_3202);
and U7518 (N_7518,N_4823,N_1184);
nor U7519 (N_7519,N_4048,N_3809);
or U7520 (N_7520,N_4071,N_3317);
and U7521 (N_7521,N_4980,N_973);
nor U7522 (N_7522,N_1036,N_1106);
or U7523 (N_7523,N_4039,N_4182);
and U7524 (N_7524,N_1487,N_1549);
nor U7525 (N_7525,N_942,N_1239);
xor U7526 (N_7526,N_92,N_4999);
xor U7527 (N_7527,N_4195,N_4338);
xor U7528 (N_7528,N_2324,N_989);
xor U7529 (N_7529,N_2104,N_757);
or U7530 (N_7530,N_4618,N_112);
nand U7531 (N_7531,N_1366,N_3358);
or U7532 (N_7532,N_3667,N_4450);
nand U7533 (N_7533,N_1473,N_2076);
xor U7534 (N_7534,N_4571,N_3901);
xnor U7535 (N_7535,N_397,N_169);
xnor U7536 (N_7536,N_3575,N_2000);
nand U7537 (N_7537,N_2381,N_201);
xnor U7538 (N_7538,N_2656,N_4895);
and U7539 (N_7539,N_4479,N_2847);
and U7540 (N_7540,N_2265,N_530);
nor U7541 (N_7541,N_3359,N_258);
nand U7542 (N_7542,N_154,N_1048);
nor U7543 (N_7543,N_2988,N_1446);
and U7544 (N_7544,N_1064,N_3190);
nand U7545 (N_7545,N_4827,N_3133);
nor U7546 (N_7546,N_2471,N_3390);
or U7547 (N_7547,N_3130,N_4212);
or U7548 (N_7548,N_514,N_3473);
or U7549 (N_7549,N_1058,N_2522);
nand U7550 (N_7550,N_1201,N_2413);
nand U7551 (N_7551,N_116,N_4137);
nand U7552 (N_7552,N_4186,N_1123);
and U7553 (N_7553,N_610,N_3167);
and U7554 (N_7554,N_3958,N_1431);
nor U7555 (N_7555,N_903,N_2542);
or U7556 (N_7556,N_2041,N_1583);
nand U7557 (N_7557,N_716,N_2630);
xor U7558 (N_7558,N_3570,N_1973);
nand U7559 (N_7559,N_3420,N_309);
nor U7560 (N_7560,N_4948,N_3181);
nand U7561 (N_7561,N_1937,N_824);
and U7562 (N_7562,N_2957,N_4607);
nand U7563 (N_7563,N_3843,N_2585);
nand U7564 (N_7564,N_2617,N_2573);
nor U7565 (N_7565,N_3364,N_2613);
and U7566 (N_7566,N_3127,N_777);
or U7567 (N_7567,N_2386,N_1207);
nand U7568 (N_7568,N_1677,N_1711);
nand U7569 (N_7569,N_1544,N_3671);
nor U7570 (N_7570,N_4755,N_1623);
and U7571 (N_7571,N_3669,N_4040);
nor U7572 (N_7572,N_2295,N_3544);
xnor U7573 (N_7573,N_2439,N_1833);
nor U7574 (N_7574,N_3898,N_3118);
xnor U7575 (N_7575,N_150,N_225);
and U7576 (N_7576,N_3904,N_566);
nand U7577 (N_7577,N_3350,N_719);
or U7578 (N_7578,N_1451,N_3972);
nor U7579 (N_7579,N_773,N_1461);
or U7580 (N_7580,N_4384,N_163);
nand U7581 (N_7581,N_3157,N_819);
xor U7582 (N_7582,N_2110,N_290);
nand U7583 (N_7583,N_1185,N_2207);
and U7584 (N_7584,N_2543,N_975);
or U7585 (N_7585,N_1001,N_2481);
and U7586 (N_7586,N_185,N_557);
nor U7587 (N_7587,N_457,N_4485);
xnor U7588 (N_7588,N_2208,N_4285);
xor U7589 (N_7589,N_3184,N_4625);
xnor U7590 (N_7590,N_1498,N_3167);
or U7591 (N_7591,N_349,N_417);
nor U7592 (N_7592,N_2132,N_3809);
xor U7593 (N_7593,N_2186,N_554);
or U7594 (N_7594,N_3696,N_87);
and U7595 (N_7595,N_1678,N_3883);
and U7596 (N_7596,N_4092,N_3503);
nor U7597 (N_7597,N_3982,N_984);
and U7598 (N_7598,N_4512,N_2554);
and U7599 (N_7599,N_2622,N_3746);
nor U7600 (N_7600,N_2470,N_2895);
nand U7601 (N_7601,N_1329,N_3854);
xnor U7602 (N_7602,N_4990,N_596);
nor U7603 (N_7603,N_3163,N_1502);
xnor U7604 (N_7604,N_4662,N_1244);
nor U7605 (N_7605,N_3212,N_1657);
nand U7606 (N_7606,N_1016,N_3109);
and U7607 (N_7607,N_3223,N_1301);
nand U7608 (N_7608,N_1218,N_2442);
and U7609 (N_7609,N_2431,N_4105);
nor U7610 (N_7610,N_4651,N_4983);
nor U7611 (N_7611,N_4295,N_3938);
xnor U7612 (N_7612,N_1975,N_4863);
or U7613 (N_7613,N_4476,N_3936);
xnor U7614 (N_7614,N_2538,N_3234);
nand U7615 (N_7615,N_2867,N_1752);
xnor U7616 (N_7616,N_1554,N_1696);
and U7617 (N_7617,N_811,N_1016);
xor U7618 (N_7618,N_4556,N_2054);
or U7619 (N_7619,N_3200,N_587);
and U7620 (N_7620,N_739,N_393);
and U7621 (N_7621,N_1802,N_408);
or U7622 (N_7622,N_1302,N_1358);
or U7623 (N_7623,N_2403,N_4930);
nand U7624 (N_7624,N_1438,N_3744);
and U7625 (N_7625,N_4049,N_2431);
nand U7626 (N_7626,N_2164,N_4728);
xnor U7627 (N_7627,N_2958,N_3501);
nand U7628 (N_7628,N_4061,N_877);
xor U7629 (N_7629,N_2932,N_1837);
xnor U7630 (N_7630,N_4306,N_2516);
xor U7631 (N_7631,N_3245,N_3282);
and U7632 (N_7632,N_2706,N_3660);
xor U7633 (N_7633,N_3710,N_3712);
and U7634 (N_7634,N_4319,N_4470);
xnor U7635 (N_7635,N_3753,N_2572);
nand U7636 (N_7636,N_3454,N_2010);
nand U7637 (N_7637,N_3805,N_2067);
and U7638 (N_7638,N_3663,N_4407);
and U7639 (N_7639,N_2517,N_3495);
nand U7640 (N_7640,N_2898,N_808);
or U7641 (N_7641,N_1615,N_109);
nor U7642 (N_7642,N_2764,N_4107);
or U7643 (N_7643,N_2703,N_1144);
xnor U7644 (N_7644,N_4871,N_3798);
xnor U7645 (N_7645,N_3937,N_2108);
or U7646 (N_7646,N_1437,N_2654);
nand U7647 (N_7647,N_671,N_3600);
xor U7648 (N_7648,N_1528,N_1896);
nor U7649 (N_7649,N_1308,N_2513);
and U7650 (N_7650,N_1057,N_108);
nor U7651 (N_7651,N_562,N_358);
nand U7652 (N_7652,N_1413,N_141);
nand U7653 (N_7653,N_187,N_1536);
and U7654 (N_7654,N_3444,N_1602);
xnor U7655 (N_7655,N_4128,N_860);
xnor U7656 (N_7656,N_537,N_2502);
or U7657 (N_7657,N_3070,N_877);
nor U7658 (N_7658,N_873,N_2256);
and U7659 (N_7659,N_296,N_3923);
xnor U7660 (N_7660,N_448,N_3956);
and U7661 (N_7661,N_4262,N_1245);
nor U7662 (N_7662,N_4132,N_1743);
xor U7663 (N_7663,N_411,N_465);
xnor U7664 (N_7664,N_3400,N_2796);
nor U7665 (N_7665,N_2975,N_242);
or U7666 (N_7666,N_4194,N_1286);
nand U7667 (N_7667,N_460,N_4065);
xnor U7668 (N_7668,N_3727,N_2876);
or U7669 (N_7669,N_1177,N_617);
xor U7670 (N_7670,N_10,N_171);
or U7671 (N_7671,N_1859,N_1565);
nand U7672 (N_7672,N_4563,N_4375);
xnor U7673 (N_7673,N_2977,N_1097);
nand U7674 (N_7674,N_4018,N_1188);
xor U7675 (N_7675,N_4911,N_2903);
xor U7676 (N_7676,N_4792,N_2732);
nand U7677 (N_7677,N_911,N_3252);
and U7678 (N_7678,N_1456,N_4548);
nand U7679 (N_7679,N_3021,N_2276);
xnor U7680 (N_7680,N_4215,N_2891);
or U7681 (N_7681,N_2057,N_529);
nor U7682 (N_7682,N_4419,N_322);
xnor U7683 (N_7683,N_2979,N_2459);
or U7684 (N_7684,N_833,N_4413);
and U7685 (N_7685,N_4639,N_3806);
nor U7686 (N_7686,N_1064,N_1101);
and U7687 (N_7687,N_3356,N_3243);
and U7688 (N_7688,N_1917,N_1670);
and U7689 (N_7689,N_3889,N_2765);
and U7690 (N_7690,N_938,N_4628);
and U7691 (N_7691,N_1458,N_2842);
and U7692 (N_7692,N_2478,N_4572);
nand U7693 (N_7693,N_220,N_2991);
nor U7694 (N_7694,N_3792,N_2811);
nor U7695 (N_7695,N_1646,N_2344);
or U7696 (N_7696,N_855,N_1799);
nand U7697 (N_7697,N_1089,N_1272);
nor U7698 (N_7698,N_2557,N_3372);
or U7699 (N_7699,N_136,N_1806);
xor U7700 (N_7700,N_1202,N_3007);
xor U7701 (N_7701,N_2551,N_2727);
nor U7702 (N_7702,N_1425,N_885);
nand U7703 (N_7703,N_937,N_515);
nor U7704 (N_7704,N_1175,N_1910);
and U7705 (N_7705,N_2616,N_4390);
nor U7706 (N_7706,N_2448,N_4509);
xnor U7707 (N_7707,N_4517,N_4257);
nor U7708 (N_7708,N_4353,N_2327);
or U7709 (N_7709,N_2806,N_3939);
nor U7710 (N_7710,N_2554,N_278);
nor U7711 (N_7711,N_4391,N_586);
xor U7712 (N_7712,N_4029,N_1776);
or U7713 (N_7713,N_342,N_4159);
nand U7714 (N_7714,N_3179,N_1349);
or U7715 (N_7715,N_2212,N_2026);
nor U7716 (N_7716,N_3285,N_788);
and U7717 (N_7717,N_424,N_4371);
nand U7718 (N_7718,N_3968,N_3686);
nand U7719 (N_7719,N_2444,N_2322);
xor U7720 (N_7720,N_1280,N_4500);
or U7721 (N_7721,N_3701,N_300);
xnor U7722 (N_7722,N_447,N_2881);
or U7723 (N_7723,N_867,N_3448);
nor U7724 (N_7724,N_3409,N_4991);
nor U7725 (N_7725,N_3609,N_4721);
or U7726 (N_7726,N_818,N_3465);
xor U7727 (N_7727,N_3842,N_604);
xor U7728 (N_7728,N_805,N_1461);
or U7729 (N_7729,N_2904,N_870);
or U7730 (N_7730,N_889,N_3715);
nand U7731 (N_7731,N_4431,N_3293);
or U7732 (N_7732,N_3947,N_2160);
nand U7733 (N_7733,N_1933,N_4976);
or U7734 (N_7734,N_4089,N_260);
nand U7735 (N_7735,N_3953,N_2063);
nand U7736 (N_7736,N_4390,N_4995);
and U7737 (N_7737,N_3989,N_3539);
or U7738 (N_7738,N_961,N_4980);
xor U7739 (N_7739,N_2642,N_3050);
and U7740 (N_7740,N_4752,N_274);
xnor U7741 (N_7741,N_1694,N_33);
nand U7742 (N_7742,N_4004,N_3296);
or U7743 (N_7743,N_362,N_1464);
nand U7744 (N_7744,N_4824,N_1342);
nand U7745 (N_7745,N_83,N_853);
xnor U7746 (N_7746,N_493,N_820);
and U7747 (N_7747,N_1420,N_4698);
nand U7748 (N_7748,N_3467,N_2780);
nor U7749 (N_7749,N_2381,N_4931);
or U7750 (N_7750,N_4987,N_236);
nor U7751 (N_7751,N_1237,N_1620);
nor U7752 (N_7752,N_4114,N_1116);
and U7753 (N_7753,N_1060,N_1034);
or U7754 (N_7754,N_4662,N_3684);
nor U7755 (N_7755,N_1615,N_1214);
nor U7756 (N_7756,N_2966,N_4978);
nand U7757 (N_7757,N_723,N_4383);
xnor U7758 (N_7758,N_2803,N_3854);
xnor U7759 (N_7759,N_3695,N_1698);
or U7760 (N_7760,N_1074,N_684);
and U7761 (N_7761,N_1232,N_2579);
and U7762 (N_7762,N_2821,N_1245);
xnor U7763 (N_7763,N_1852,N_4920);
nor U7764 (N_7764,N_405,N_4967);
and U7765 (N_7765,N_1449,N_712);
nor U7766 (N_7766,N_3424,N_4499);
and U7767 (N_7767,N_4200,N_1463);
or U7768 (N_7768,N_3485,N_4744);
nand U7769 (N_7769,N_895,N_4859);
xnor U7770 (N_7770,N_3131,N_2925);
nor U7771 (N_7771,N_58,N_2873);
or U7772 (N_7772,N_3043,N_953);
xnor U7773 (N_7773,N_1353,N_495);
xor U7774 (N_7774,N_4923,N_3193);
nand U7775 (N_7775,N_1130,N_1029);
xor U7776 (N_7776,N_1684,N_3847);
nand U7777 (N_7777,N_1687,N_1943);
xnor U7778 (N_7778,N_2234,N_4748);
nor U7779 (N_7779,N_3859,N_2018);
or U7780 (N_7780,N_3408,N_1481);
xor U7781 (N_7781,N_2198,N_4762);
and U7782 (N_7782,N_3940,N_2350);
nand U7783 (N_7783,N_2553,N_2290);
or U7784 (N_7784,N_3269,N_1267);
and U7785 (N_7785,N_1635,N_2140);
nand U7786 (N_7786,N_4620,N_1979);
or U7787 (N_7787,N_3756,N_3555);
nor U7788 (N_7788,N_3109,N_259);
nor U7789 (N_7789,N_3206,N_2512);
or U7790 (N_7790,N_3032,N_4537);
xnor U7791 (N_7791,N_543,N_4811);
or U7792 (N_7792,N_3912,N_35);
xor U7793 (N_7793,N_3290,N_4889);
nor U7794 (N_7794,N_3016,N_2132);
xor U7795 (N_7795,N_3752,N_198);
or U7796 (N_7796,N_4600,N_2641);
nand U7797 (N_7797,N_1796,N_3174);
and U7798 (N_7798,N_3215,N_552);
and U7799 (N_7799,N_4331,N_1318);
xor U7800 (N_7800,N_1444,N_883);
nor U7801 (N_7801,N_1446,N_1221);
xor U7802 (N_7802,N_4012,N_1617);
nor U7803 (N_7803,N_237,N_4553);
or U7804 (N_7804,N_3529,N_4995);
or U7805 (N_7805,N_874,N_4670);
and U7806 (N_7806,N_3776,N_2569);
and U7807 (N_7807,N_4799,N_2895);
and U7808 (N_7808,N_4114,N_3063);
nand U7809 (N_7809,N_685,N_385);
nand U7810 (N_7810,N_1477,N_3442);
nor U7811 (N_7811,N_4872,N_4147);
nand U7812 (N_7812,N_207,N_4517);
nor U7813 (N_7813,N_2366,N_2923);
nor U7814 (N_7814,N_4950,N_3214);
or U7815 (N_7815,N_1498,N_4476);
nand U7816 (N_7816,N_3029,N_42);
nor U7817 (N_7817,N_1625,N_817);
and U7818 (N_7818,N_4216,N_4781);
nand U7819 (N_7819,N_215,N_1878);
and U7820 (N_7820,N_967,N_3915);
and U7821 (N_7821,N_2804,N_3320);
nor U7822 (N_7822,N_4477,N_1507);
nor U7823 (N_7823,N_2603,N_3185);
and U7824 (N_7824,N_2430,N_3567);
xor U7825 (N_7825,N_4030,N_4732);
and U7826 (N_7826,N_1969,N_2752);
nand U7827 (N_7827,N_3642,N_4463);
or U7828 (N_7828,N_746,N_3787);
and U7829 (N_7829,N_3870,N_2001);
xor U7830 (N_7830,N_4203,N_3256);
nor U7831 (N_7831,N_4282,N_3313);
nand U7832 (N_7832,N_4505,N_841);
xnor U7833 (N_7833,N_591,N_1598);
or U7834 (N_7834,N_3964,N_1524);
nor U7835 (N_7835,N_2443,N_4529);
nor U7836 (N_7836,N_1271,N_3537);
or U7837 (N_7837,N_118,N_3289);
or U7838 (N_7838,N_1488,N_3924);
and U7839 (N_7839,N_2364,N_1009);
or U7840 (N_7840,N_1778,N_4174);
nand U7841 (N_7841,N_2780,N_56);
nand U7842 (N_7842,N_4337,N_3979);
nand U7843 (N_7843,N_3421,N_3228);
and U7844 (N_7844,N_3912,N_1439);
nand U7845 (N_7845,N_255,N_4381);
or U7846 (N_7846,N_1201,N_1599);
and U7847 (N_7847,N_3042,N_2365);
nand U7848 (N_7848,N_530,N_278);
xor U7849 (N_7849,N_2473,N_3263);
nor U7850 (N_7850,N_2057,N_749);
nor U7851 (N_7851,N_1066,N_1689);
xor U7852 (N_7852,N_422,N_4801);
and U7853 (N_7853,N_3934,N_4193);
nand U7854 (N_7854,N_3450,N_79);
and U7855 (N_7855,N_70,N_4785);
or U7856 (N_7856,N_2345,N_0);
nor U7857 (N_7857,N_4503,N_964);
and U7858 (N_7858,N_3716,N_671);
xnor U7859 (N_7859,N_1990,N_3508);
xor U7860 (N_7860,N_2079,N_961);
nor U7861 (N_7861,N_3245,N_724);
or U7862 (N_7862,N_3271,N_2792);
nand U7863 (N_7863,N_3588,N_4153);
nor U7864 (N_7864,N_3480,N_4923);
and U7865 (N_7865,N_454,N_1309);
or U7866 (N_7866,N_4498,N_63);
xor U7867 (N_7867,N_879,N_3847);
nor U7868 (N_7868,N_2161,N_2532);
nand U7869 (N_7869,N_4690,N_4001);
nand U7870 (N_7870,N_2603,N_2062);
and U7871 (N_7871,N_613,N_1600);
nor U7872 (N_7872,N_1392,N_3590);
nor U7873 (N_7873,N_3454,N_3047);
and U7874 (N_7874,N_547,N_4473);
nor U7875 (N_7875,N_4987,N_1739);
or U7876 (N_7876,N_884,N_4147);
nand U7877 (N_7877,N_1506,N_3754);
nand U7878 (N_7878,N_2219,N_3902);
or U7879 (N_7879,N_686,N_3882);
nor U7880 (N_7880,N_277,N_3565);
or U7881 (N_7881,N_1699,N_4724);
nor U7882 (N_7882,N_4102,N_2712);
or U7883 (N_7883,N_3092,N_3533);
or U7884 (N_7884,N_4072,N_562);
xor U7885 (N_7885,N_1701,N_3037);
nand U7886 (N_7886,N_3882,N_3294);
xor U7887 (N_7887,N_2493,N_139);
and U7888 (N_7888,N_3790,N_160);
and U7889 (N_7889,N_2534,N_3847);
and U7890 (N_7890,N_999,N_1671);
nor U7891 (N_7891,N_810,N_4302);
nor U7892 (N_7892,N_3288,N_1294);
or U7893 (N_7893,N_449,N_1508);
and U7894 (N_7894,N_2157,N_2236);
nor U7895 (N_7895,N_2313,N_1079);
or U7896 (N_7896,N_4559,N_2108);
nor U7897 (N_7897,N_45,N_1721);
and U7898 (N_7898,N_2486,N_4048);
and U7899 (N_7899,N_3713,N_1155);
or U7900 (N_7900,N_818,N_4584);
nor U7901 (N_7901,N_4804,N_2210);
and U7902 (N_7902,N_3867,N_168);
and U7903 (N_7903,N_4794,N_2195);
xnor U7904 (N_7904,N_2166,N_670);
nor U7905 (N_7905,N_680,N_875);
xor U7906 (N_7906,N_819,N_1178);
nand U7907 (N_7907,N_1800,N_4778);
nor U7908 (N_7908,N_2182,N_2152);
xor U7909 (N_7909,N_22,N_4876);
or U7910 (N_7910,N_816,N_2293);
nand U7911 (N_7911,N_2488,N_3771);
xnor U7912 (N_7912,N_2321,N_606);
xor U7913 (N_7913,N_907,N_4796);
nand U7914 (N_7914,N_2967,N_1832);
nor U7915 (N_7915,N_3972,N_4930);
xor U7916 (N_7916,N_2024,N_3317);
xnor U7917 (N_7917,N_1863,N_173);
nor U7918 (N_7918,N_4290,N_2040);
nor U7919 (N_7919,N_2080,N_2507);
xor U7920 (N_7920,N_401,N_3781);
xnor U7921 (N_7921,N_927,N_4941);
nand U7922 (N_7922,N_4563,N_2331);
or U7923 (N_7923,N_2130,N_1665);
and U7924 (N_7924,N_3874,N_4504);
xnor U7925 (N_7925,N_595,N_1049);
or U7926 (N_7926,N_2272,N_1093);
nor U7927 (N_7927,N_2666,N_4015);
xor U7928 (N_7928,N_2400,N_4384);
nor U7929 (N_7929,N_101,N_1098);
nand U7930 (N_7930,N_489,N_2259);
nand U7931 (N_7931,N_2596,N_3754);
xnor U7932 (N_7932,N_4302,N_4499);
or U7933 (N_7933,N_1084,N_4515);
nor U7934 (N_7934,N_1973,N_4683);
or U7935 (N_7935,N_2779,N_703);
and U7936 (N_7936,N_4591,N_4222);
and U7937 (N_7937,N_686,N_124);
and U7938 (N_7938,N_3878,N_1735);
or U7939 (N_7939,N_1038,N_3893);
nand U7940 (N_7940,N_2412,N_4196);
nand U7941 (N_7941,N_943,N_242);
nor U7942 (N_7942,N_3516,N_4547);
nand U7943 (N_7943,N_4990,N_2897);
nor U7944 (N_7944,N_3639,N_901);
and U7945 (N_7945,N_625,N_4154);
and U7946 (N_7946,N_2515,N_2030);
nor U7947 (N_7947,N_4198,N_48);
and U7948 (N_7948,N_2294,N_356);
xor U7949 (N_7949,N_2218,N_1275);
nand U7950 (N_7950,N_756,N_2622);
xor U7951 (N_7951,N_4449,N_356);
xor U7952 (N_7952,N_2200,N_2662);
nand U7953 (N_7953,N_2852,N_4748);
or U7954 (N_7954,N_4883,N_1860);
xnor U7955 (N_7955,N_3967,N_2486);
nor U7956 (N_7956,N_3261,N_4978);
or U7957 (N_7957,N_4135,N_431);
or U7958 (N_7958,N_1302,N_2188);
and U7959 (N_7959,N_1744,N_3800);
and U7960 (N_7960,N_1073,N_1957);
nand U7961 (N_7961,N_836,N_3794);
or U7962 (N_7962,N_529,N_2286);
nor U7963 (N_7963,N_2851,N_1404);
nand U7964 (N_7964,N_3431,N_4171);
nand U7965 (N_7965,N_4822,N_3060);
or U7966 (N_7966,N_1819,N_456);
xor U7967 (N_7967,N_3915,N_1131);
nand U7968 (N_7968,N_3757,N_1719);
and U7969 (N_7969,N_18,N_3795);
nor U7970 (N_7970,N_9,N_792);
or U7971 (N_7971,N_4434,N_4594);
nor U7972 (N_7972,N_4115,N_1247);
and U7973 (N_7973,N_3742,N_4505);
and U7974 (N_7974,N_3875,N_4056);
or U7975 (N_7975,N_4494,N_1670);
xor U7976 (N_7976,N_4490,N_3982);
nor U7977 (N_7977,N_3995,N_2041);
xor U7978 (N_7978,N_4785,N_4717);
or U7979 (N_7979,N_2978,N_4209);
nor U7980 (N_7980,N_1666,N_2802);
and U7981 (N_7981,N_4068,N_159);
and U7982 (N_7982,N_2593,N_4256);
or U7983 (N_7983,N_3251,N_1264);
nand U7984 (N_7984,N_1548,N_2528);
nor U7985 (N_7985,N_828,N_3036);
nand U7986 (N_7986,N_229,N_1538);
or U7987 (N_7987,N_108,N_289);
xor U7988 (N_7988,N_487,N_3138);
nand U7989 (N_7989,N_4114,N_1906);
or U7990 (N_7990,N_1105,N_530);
nor U7991 (N_7991,N_2137,N_3500);
nand U7992 (N_7992,N_1930,N_222);
xor U7993 (N_7993,N_324,N_67);
nand U7994 (N_7994,N_1110,N_374);
nand U7995 (N_7995,N_2495,N_2563);
xnor U7996 (N_7996,N_3909,N_1029);
nand U7997 (N_7997,N_2837,N_3292);
nor U7998 (N_7998,N_908,N_2912);
or U7999 (N_7999,N_2652,N_4853);
or U8000 (N_8000,N_2146,N_4366);
and U8001 (N_8001,N_4294,N_3711);
xor U8002 (N_8002,N_1577,N_41);
nor U8003 (N_8003,N_1974,N_4969);
xnor U8004 (N_8004,N_1439,N_2046);
xor U8005 (N_8005,N_3997,N_666);
nand U8006 (N_8006,N_2465,N_3152);
nor U8007 (N_8007,N_986,N_2034);
or U8008 (N_8008,N_4799,N_4405);
or U8009 (N_8009,N_2462,N_3383);
nor U8010 (N_8010,N_1819,N_4438);
nand U8011 (N_8011,N_2408,N_3793);
xnor U8012 (N_8012,N_438,N_3340);
nor U8013 (N_8013,N_4970,N_424);
nor U8014 (N_8014,N_4780,N_4378);
xor U8015 (N_8015,N_588,N_1467);
nand U8016 (N_8016,N_4411,N_2688);
nor U8017 (N_8017,N_3862,N_2317);
nand U8018 (N_8018,N_2522,N_2268);
or U8019 (N_8019,N_955,N_1939);
and U8020 (N_8020,N_3888,N_4493);
nand U8021 (N_8021,N_2912,N_3062);
nand U8022 (N_8022,N_2084,N_2250);
nor U8023 (N_8023,N_4690,N_665);
and U8024 (N_8024,N_2261,N_717);
xnor U8025 (N_8025,N_3803,N_1343);
nor U8026 (N_8026,N_833,N_3217);
nor U8027 (N_8027,N_2602,N_490);
nand U8028 (N_8028,N_4505,N_1073);
and U8029 (N_8029,N_779,N_1533);
xor U8030 (N_8030,N_1511,N_673);
or U8031 (N_8031,N_3501,N_4304);
xnor U8032 (N_8032,N_2599,N_3402);
xor U8033 (N_8033,N_4092,N_214);
xor U8034 (N_8034,N_713,N_3127);
nand U8035 (N_8035,N_965,N_4989);
nand U8036 (N_8036,N_4552,N_1187);
xnor U8037 (N_8037,N_2634,N_4657);
nor U8038 (N_8038,N_3747,N_2272);
xnor U8039 (N_8039,N_2183,N_2430);
nand U8040 (N_8040,N_3381,N_259);
or U8041 (N_8041,N_4740,N_306);
and U8042 (N_8042,N_1060,N_1360);
nand U8043 (N_8043,N_1135,N_3533);
nor U8044 (N_8044,N_2834,N_3685);
and U8045 (N_8045,N_1813,N_1468);
nor U8046 (N_8046,N_700,N_3429);
and U8047 (N_8047,N_2148,N_3633);
nor U8048 (N_8048,N_3048,N_4220);
nand U8049 (N_8049,N_1122,N_2604);
nand U8050 (N_8050,N_2468,N_3836);
nor U8051 (N_8051,N_4177,N_487);
xor U8052 (N_8052,N_2238,N_4010);
and U8053 (N_8053,N_2814,N_544);
or U8054 (N_8054,N_3882,N_3562);
nand U8055 (N_8055,N_501,N_1583);
and U8056 (N_8056,N_1464,N_2481);
or U8057 (N_8057,N_4127,N_3978);
nor U8058 (N_8058,N_2625,N_4008);
and U8059 (N_8059,N_3998,N_297);
xnor U8060 (N_8060,N_171,N_1001);
nand U8061 (N_8061,N_3792,N_3998);
and U8062 (N_8062,N_3590,N_3565);
xnor U8063 (N_8063,N_3546,N_2548);
nor U8064 (N_8064,N_4406,N_3024);
xnor U8065 (N_8065,N_2435,N_623);
or U8066 (N_8066,N_4694,N_413);
and U8067 (N_8067,N_2423,N_3526);
nor U8068 (N_8068,N_308,N_3050);
nor U8069 (N_8069,N_1621,N_1433);
nor U8070 (N_8070,N_2335,N_721);
nor U8071 (N_8071,N_869,N_918);
nor U8072 (N_8072,N_3332,N_4545);
or U8073 (N_8073,N_656,N_4930);
or U8074 (N_8074,N_1716,N_80);
nor U8075 (N_8075,N_2112,N_858);
nor U8076 (N_8076,N_4126,N_763);
nor U8077 (N_8077,N_2720,N_2364);
xor U8078 (N_8078,N_3951,N_4827);
nor U8079 (N_8079,N_1342,N_113);
or U8080 (N_8080,N_2487,N_2316);
xor U8081 (N_8081,N_1017,N_4873);
and U8082 (N_8082,N_2793,N_286);
xor U8083 (N_8083,N_963,N_3299);
nand U8084 (N_8084,N_1469,N_4676);
nand U8085 (N_8085,N_3423,N_1404);
and U8086 (N_8086,N_3182,N_2400);
or U8087 (N_8087,N_4243,N_530);
xnor U8088 (N_8088,N_1030,N_2756);
or U8089 (N_8089,N_3093,N_4770);
and U8090 (N_8090,N_1030,N_2780);
xor U8091 (N_8091,N_4758,N_837);
or U8092 (N_8092,N_2244,N_2650);
nand U8093 (N_8093,N_3871,N_3081);
and U8094 (N_8094,N_3236,N_1672);
xor U8095 (N_8095,N_534,N_2121);
xor U8096 (N_8096,N_1776,N_4888);
nor U8097 (N_8097,N_873,N_3409);
nor U8098 (N_8098,N_4407,N_4162);
nor U8099 (N_8099,N_4779,N_1469);
or U8100 (N_8100,N_3934,N_2825);
and U8101 (N_8101,N_2221,N_1370);
xor U8102 (N_8102,N_4379,N_2854);
nor U8103 (N_8103,N_767,N_2327);
nor U8104 (N_8104,N_1288,N_3941);
xor U8105 (N_8105,N_2352,N_3332);
nand U8106 (N_8106,N_4436,N_2851);
nand U8107 (N_8107,N_731,N_758);
and U8108 (N_8108,N_657,N_3841);
xnor U8109 (N_8109,N_412,N_4851);
nor U8110 (N_8110,N_753,N_4874);
nor U8111 (N_8111,N_1291,N_34);
nor U8112 (N_8112,N_3365,N_2401);
nor U8113 (N_8113,N_3243,N_4460);
nand U8114 (N_8114,N_1511,N_165);
and U8115 (N_8115,N_4817,N_2869);
xnor U8116 (N_8116,N_4473,N_2598);
or U8117 (N_8117,N_2750,N_2583);
and U8118 (N_8118,N_1603,N_2237);
nand U8119 (N_8119,N_3667,N_688);
or U8120 (N_8120,N_466,N_1054);
nor U8121 (N_8121,N_2747,N_2063);
nor U8122 (N_8122,N_1363,N_3497);
and U8123 (N_8123,N_2917,N_2025);
and U8124 (N_8124,N_2972,N_1169);
and U8125 (N_8125,N_2243,N_2861);
nand U8126 (N_8126,N_296,N_3847);
or U8127 (N_8127,N_2849,N_2514);
nor U8128 (N_8128,N_2937,N_1860);
or U8129 (N_8129,N_3235,N_4518);
xor U8130 (N_8130,N_1417,N_3283);
nor U8131 (N_8131,N_2935,N_2931);
nand U8132 (N_8132,N_3904,N_4244);
nand U8133 (N_8133,N_3049,N_1685);
nand U8134 (N_8134,N_1456,N_2145);
or U8135 (N_8135,N_3846,N_2953);
nor U8136 (N_8136,N_4641,N_2830);
or U8137 (N_8137,N_4382,N_571);
nor U8138 (N_8138,N_496,N_2809);
or U8139 (N_8139,N_4465,N_3661);
and U8140 (N_8140,N_2552,N_2363);
nor U8141 (N_8141,N_3952,N_3614);
or U8142 (N_8142,N_3917,N_317);
nor U8143 (N_8143,N_1323,N_1855);
nor U8144 (N_8144,N_4588,N_2725);
and U8145 (N_8145,N_1829,N_1693);
xnor U8146 (N_8146,N_1619,N_491);
xnor U8147 (N_8147,N_2505,N_3922);
or U8148 (N_8148,N_4967,N_311);
nor U8149 (N_8149,N_4241,N_1690);
or U8150 (N_8150,N_1315,N_3361);
nand U8151 (N_8151,N_2060,N_2203);
nand U8152 (N_8152,N_4086,N_270);
nor U8153 (N_8153,N_3758,N_985);
nor U8154 (N_8154,N_2176,N_4490);
and U8155 (N_8155,N_345,N_648);
nor U8156 (N_8156,N_2452,N_3878);
xnor U8157 (N_8157,N_808,N_2425);
and U8158 (N_8158,N_3131,N_1242);
nor U8159 (N_8159,N_2261,N_3049);
nand U8160 (N_8160,N_393,N_1107);
and U8161 (N_8161,N_937,N_2976);
xor U8162 (N_8162,N_3890,N_2578);
nor U8163 (N_8163,N_365,N_2558);
xnor U8164 (N_8164,N_699,N_1572);
nor U8165 (N_8165,N_3376,N_4394);
xor U8166 (N_8166,N_2453,N_4947);
nor U8167 (N_8167,N_2696,N_2216);
nor U8168 (N_8168,N_839,N_2634);
nand U8169 (N_8169,N_1821,N_2715);
or U8170 (N_8170,N_542,N_2223);
or U8171 (N_8171,N_884,N_2773);
or U8172 (N_8172,N_1470,N_697);
and U8173 (N_8173,N_2335,N_3724);
and U8174 (N_8174,N_1026,N_3847);
xnor U8175 (N_8175,N_3034,N_4957);
xor U8176 (N_8176,N_2713,N_4890);
or U8177 (N_8177,N_143,N_359);
or U8178 (N_8178,N_4519,N_1561);
nand U8179 (N_8179,N_4376,N_1779);
nand U8180 (N_8180,N_2234,N_4691);
xnor U8181 (N_8181,N_850,N_830);
nand U8182 (N_8182,N_1846,N_4054);
xnor U8183 (N_8183,N_1348,N_2009);
or U8184 (N_8184,N_4243,N_1861);
xnor U8185 (N_8185,N_2132,N_4812);
nand U8186 (N_8186,N_92,N_2700);
xor U8187 (N_8187,N_705,N_1850);
nand U8188 (N_8188,N_3720,N_1684);
nor U8189 (N_8189,N_1183,N_1750);
nor U8190 (N_8190,N_2390,N_83);
and U8191 (N_8191,N_4257,N_1225);
and U8192 (N_8192,N_378,N_934);
nand U8193 (N_8193,N_3064,N_3146);
or U8194 (N_8194,N_4826,N_963);
nor U8195 (N_8195,N_3433,N_250);
and U8196 (N_8196,N_1020,N_646);
nand U8197 (N_8197,N_3044,N_1572);
xnor U8198 (N_8198,N_1684,N_2654);
nor U8199 (N_8199,N_3244,N_4598);
nand U8200 (N_8200,N_4111,N_1950);
xnor U8201 (N_8201,N_1303,N_1479);
or U8202 (N_8202,N_2314,N_2546);
or U8203 (N_8203,N_3355,N_4125);
nor U8204 (N_8204,N_1749,N_4349);
and U8205 (N_8205,N_3938,N_3723);
or U8206 (N_8206,N_3419,N_2544);
xnor U8207 (N_8207,N_2915,N_4065);
or U8208 (N_8208,N_4559,N_4056);
nor U8209 (N_8209,N_3660,N_1903);
nor U8210 (N_8210,N_2777,N_4610);
nand U8211 (N_8211,N_2064,N_4914);
nor U8212 (N_8212,N_1525,N_689);
nor U8213 (N_8213,N_3573,N_2657);
and U8214 (N_8214,N_1399,N_4726);
or U8215 (N_8215,N_99,N_2753);
or U8216 (N_8216,N_3248,N_3625);
nor U8217 (N_8217,N_2126,N_1119);
xnor U8218 (N_8218,N_3775,N_290);
and U8219 (N_8219,N_2606,N_3718);
nor U8220 (N_8220,N_1588,N_1828);
xor U8221 (N_8221,N_4097,N_3255);
or U8222 (N_8222,N_4985,N_548);
nand U8223 (N_8223,N_3172,N_4294);
xor U8224 (N_8224,N_4505,N_1150);
nand U8225 (N_8225,N_2001,N_40);
nand U8226 (N_8226,N_4112,N_1403);
xnor U8227 (N_8227,N_4264,N_2472);
or U8228 (N_8228,N_2562,N_2949);
xnor U8229 (N_8229,N_1600,N_739);
xnor U8230 (N_8230,N_2061,N_816);
and U8231 (N_8231,N_1865,N_2107);
and U8232 (N_8232,N_2110,N_3489);
or U8233 (N_8233,N_538,N_513);
and U8234 (N_8234,N_3037,N_4429);
or U8235 (N_8235,N_4634,N_3587);
and U8236 (N_8236,N_3009,N_3851);
nor U8237 (N_8237,N_3649,N_4285);
nor U8238 (N_8238,N_2102,N_3126);
or U8239 (N_8239,N_1498,N_448);
xnor U8240 (N_8240,N_4864,N_989);
nor U8241 (N_8241,N_3255,N_1869);
xnor U8242 (N_8242,N_3086,N_795);
nand U8243 (N_8243,N_268,N_2975);
nor U8244 (N_8244,N_3036,N_3343);
nand U8245 (N_8245,N_3826,N_3861);
nor U8246 (N_8246,N_1700,N_1418);
xor U8247 (N_8247,N_3847,N_2451);
or U8248 (N_8248,N_1970,N_908);
nand U8249 (N_8249,N_1066,N_2435);
nand U8250 (N_8250,N_1208,N_1078);
nor U8251 (N_8251,N_2216,N_1447);
or U8252 (N_8252,N_4795,N_2214);
xor U8253 (N_8253,N_37,N_2913);
and U8254 (N_8254,N_3824,N_3417);
and U8255 (N_8255,N_4404,N_4558);
or U8256 (N_8256,N_3543,N_4512);
or U8257 (N_8257,N_1825,N_1627);
and U8258 (N_8258,N_4393,N_4992);
xor U8259 (N_8259,N_2836,N_3283);
or U8260 (N_8260,N_2844,N_4428);
xor U8261 (N_8261,N_2302,N_4755);
nand U8262 (N_8262,N_4225,N_364);
or U8263 (N_8263,N_1163,N_572);
nor U8264 (N_8264,N_4342,N_2568);
or U8265 (N_8265,N_987,N_306);
nor U8266 (N_8266,N_2319,N_1486);
nor U8267 (N_8267,N_929,N_1695);
nor U8268 (N_8268,N_1138,N_4207);
xnor U8269 (N_8269,N_3996,N_334);
nor U8270 (N_8270,N_2186,N_2570);
and U8271 (N_8271,N_829,N_1896);
nand U8272 (N_8272,N_2700,N_2567);
and U8273 (N_8273,N_2064,N_4809);
or U8274 (N_8274,N_155,N_4989);
nand U8275 (N_8275,N_3730,N_2155);
nand U8276 (N_8276,N_2732,N_2035);
nand U8277 (N_8277,N_4078,N_4607);
and U8278 (N_8278,N_34,N_2536);
nand U8279 (N_8279,N_3046,N_2557);
xnor U8280 (N_8280,N_3884,N_831);
xor U8281 (N_8281,N_135,N_1481);
or U8282 (N_8282,N_3575,N_1307);
or U8283 (N_8283,N_1091,N_1799);
nor U8284 (N_8284,N_1902,N_929);
nand U8285 (N_8285,N_39,N_2606);
and U8286 (N_8286,N_2168,N_2545);
nor U8287 (N_8287,N_4855,N_4440);
nor U8288 (N_8288,N_2586,N_3215);
nor U8289 (N_8289,N_2673,N_1279);
nand U8290 (N_8290,N_4189,N_2232);
nor U8291 (N_8291,N_1747,N_250);
nor U8292 (N_8292,N_787,N_4027);
nand U8293 (N_8293,N_38,N_2305);
xor U8294 (N_8294,N_1421,N_3209);
nor U8295 (N_8295,N_3164,N_309);
and U8296 (N_8296,N_3599,N_1140);
or U8297 (N_8297,N_459,N_145);
and U8298 (N_8298,N_376,N_4503);
and U8299 (N_8299,N_4171,N_789);
xnor U8300 (N_8300,N_4247,N_1982);
nand U8301 (N_8301,N_276,N_4336);
and U8302 (N_8302,N_2795,N_1276);
or U8303 (N_8303,N_4143,N_3537);
nand U8304 (N_8304,N_497,N_3319);
nand U8305 (N_8305,N_1171,N_2906);
or U8306 (N_8306,N_1032,N_1428);
and U8307 (N_8307,N_3343,N_1965);
nand U8308 (N_8308,N_2302,N_325);
or U8309 (N_8309,N_2798,N_2316);
nor U8310 (N_8310,N_3222,N_1011);
or U8311 (N_8311,N_4552,N_2057);
and U8312 (N_8312,N_2984,N_4876);
and U8313 (N_8313,N_4641,N_1033);
nand U8314 (N_8314,N_2492,N_174);
or U8315 (N_8315,N_2485,N_1557);
xor U8316 (N_8316,N_46,N_3778);
xor U8317 (N_8317,N_2327,N_2040);
nand U8318 (N_8318,N_1168,N_2230);
nand U8319 (N_8319,N_634,N_237);
or U8320 (N_8320,N_2524,N_754);
nor U8321 (N_8321,N_1071,N_464);
or U8322 (N_8322,N_3524,N_326);
xnor U8323 (N_8323,N_2517,N_2009);
xor U8324 (N_8324,N_4353,N_1418);
xnor U8325 (N_8325,N_4883,N_712);
or U8326 (N_8326,N_1256,N_3601);
nor U8327 (N_8327,N_97,N_4334);
or U8328 (N_8328,N_4185,N_1346);
or U8329 (N_8329,N_1590,N_1722);
and U8330 (N_8330,N_1590,N_3755);
nand U8331 (N_8331,N_2749,N_1028);
nand U8332 (N_8332,N_4537,N_480);
nand U8333 (N_8333,N_1103,N_2073);
nand U8334 (N_8334,N_2326,N_2120);
and U8335 (N_8335,N_4008,N_1578);
or U8336 (N_8336,N_1565,N_3563);
and U8337 (N_8337,N_3214,N_4386);
and U8338 (N_8338,N_4381,N_3576);
and U8339 (N_8339,N_2659,N_1231);
and U8340 (N_8340,N_4935,N_2941);
nor U8341 (N_8341,N_1085,N_3468);
nand U8342 (N_8342,N_549,N_3325);
nand U8343 (N_8343,N_4146,N_2625);
xnor U8344 (N_8344,N_4880,N_3891);
nand U8345 (N_8345,N_537,N_2553);
nor U8346 (N_8346,N_4148,N_2181);
xor U8347 (N_8347,N_765,N_2679);
or U8348 (N_8348,N_251,N_2289);
xnor U8349 (N_8349,N_3279,N_2713);
or U8350 (N_8350,N_4131,N_1670);
or U8351 (N_8351,N_653,N_76);
or U8352 (N_8352,N_2381,N_124);
and U8353 (N_8353,N_2757,N_4858);
and U8354 (N_8354,N_4513,N_2884);
nand U8355 (N_8355,N_3606,N_3439);
nor U8356 (N_8356,N_1547,N_242);
and U8357 (N_8357,N_3008,N_1886);
nand U8358 (N_8358,N_3604,N_158);
and U8359 (N_8359,N_3015,N_3099);
or U8360 (N_8360,N_928,N_2308);
and U8361 (N_8361,N_26,N_3100);
nor U8362 (N_8362,N_892,N_1164);
nand U8363 (N_8363,N_571,N_2479);
xor U8364 (N_8364,N_1525,N_3589);
and U8365 (N_8365,N_3719,N_2642);
xnor U8366 (N_8366,N_4584,N_107);
nand U8367 (N_8367,N_3256,N_2532);
nand U8368 (N_8368,N_734,N_4180);
nand U8369 (N_8369,N_1002,N_4998);
and U8370 (N_8370,N_2916,N_3903);
xnor U8371 (N_8371,N_544,N_1831);
or U8372 (N_8372,N_2830,N_386);
nor U8373 (N_8373,N_954,N_600);
or U8374 (N_8374,N_2457,N_1407);
nand U8375 (N_8375,N_2822,N_1383);
or U8376 (N_8376,N_400,N_2592);
or U8377 (N_8377,N_1804,N_563);
xor U8378 (N_8378,N_2978,N_1806);
xor U8379 (N_8379,N_1728,N_4461);
and U8380 (N_8380,N_1427,N_3896);
nor U8381 (N_8381,N_4216,N_2386);
xnor U8382 (N_8382,N_3277,N_886);
and U8383 (N_8383,N_4369,N_620);
xor U8384 (N_8384,N_1983,N_4673);
xor U8385 (N_8385,N_1677,N_2687);
nand U8386 (N_8386,N_1828,N_986);
or U8387 (N_8387,N_557,N_884);
nand U8388 (N_8388,N_1366,N_2223);
nand U8389 (N_8389,N_2176,N_360);
nor U8390 (N_8390,N_4417,N_4747);
nand U8391 (N_8391,N_2122,N_1950);
xnor U8392 (N_8392,N_1778,N_4578);
and U8393 (N_8393,N_692,N_4498);
nor U8394 (N_8394,N_1130,N_1228);
xor U8395 (N_8395,N_4373,N_2951);
or U8396 (N_8396,N_874,N_1506);
nor U8397 (N_8397,N_1118,N_1619);
and U8398 (N_8398,N_1535,N_3589);
and U8399 (N_8399,N_1832,N_1953);
nand U8400 (N_8400,N_4874,N_4730);
nand U8401 (N_8401,N_2492,N_2809);
and U8402 (N_8402,N_2466,N_1849);
nor U8403 (N_8403,N_1191,N_3712);
or U8404 (N_8404,N_3518,N_3284);
or U8405 (N_8405,N_26,N_1851);
nand U8406 (N_8406,N_4314,N_1615);
and U8407 (N_8407,N_3858,N_4618);
nor U8408 (N_8408,N_947,N_4976);
nor U8409 (N_8409,N_4371,N_4549);
or U8410 (N_8410,N_220,N_4781);
nand U8411 (N_8411,N_4988,N_296);
nand U8412 (N_8412,N_3298,N_3140);
xnor U8413 (N_8413,N_784,N_1022);
nor U8414 (N_8414,N_3152,N_3473);
and U8415 (N_8415,N_2144,N_2816);
and U8416 (N_8416,N_4326,N_4168);
nand U8417 (N_8417,N_4995,N_2215);
nor U8418 (N_8418,N_4410,N_4685);
nand U8419 (N_8419,N_3222,N_622);
nor U8420 (N_8420,N_723,N_799);
nor U8421 (N_8421,N_4351,N_4007);
or U8422 (N_8422,N_827,N_817);
or U8423 (N_8423,N_4698,N_4721);
nor U8424 (N_8424,N_2296,N_416);
nor U8425 (N_8425,N_1019,N_799);
nand U8426 (N_8426,N_4978,N_3836);
and U8427 (N_8427,N_3310,N_2484);
or U8428 (N_8428,N_4190,N_3512);
and U8429 (N_8429,N_2687,N_3293);
nand U8430 (N_8430,N_2809,N_1352);
xnor U8431 (N_8431,N_4166,N_543);
xnor U8432 (N_8432,N_2977,N_2983);
nor U8433 (N_8433,N_2934,N_193);
xnor U8434 (N_8434,N_3100,N_3371);
and U8435 (N_8435,N_3131,N_2072);
or U8436 (N_8436,N_1044,N_4495);
and U8437 (N_8437,N_3002,N_2395);
nor U8438 (N_8438,N_4629,N_4742);
and U8439 (N_8439,N_3153,N_4611);
xor U8440 (N_8440,N_3021,N_4023);
and U8441 (N_8441,N_3552,N_3008);
or U8442 (N_8442,N_1765,N_2797);
xor U8443 (N_8443,N_1304,N_1048);
or U8444 (N_8444,N_3366,N_2550);
or U8445 (N_8445,N_4449,N_3554);
xor U8446 (N_8446,N_3661,N_2653);
nand U8447 (N_8447,N_2400,N_1034);
nor U8448 (N_8448,N_4920,N_4959);
nor U8449 (N_8449,N_4696,N_4900);
and U8450 (N_8450,N_1904,N_1403);
nand U8451 (N_8451,N_819,N_2911);
or U8452 (N_8452,N_4194,N_1329);
xor U8453 (N_8453,N_1096,N_4480);
xnor U8454 (N_8454,N_50,N_329);
xor U8455 (N_8455,N_741,N_4135);
and U8456 (N_8456,N_1645,N_2975);
and U8457 (N_8457,N_3930,N_3517);
nand U8458 (N_8458,N_685,N_1575);
and U8459 (N_8459,N_632,N_4549);
and U8460 (N_8460,N_1050,N_3370);
or U8461 (N_8461,N_1269,N_628);
nor U8462 (N_8462,N_2767,N_2847);
or U8463 (N_8463,N_1274,N_2879);
and U8464 (N_8464,N_3505,N_418);
nand U8465 (N_8465,N_1375,N_2456);
nor U8466 (N_8466,N_4039,N_1856);
or U8467 (N_8467,N_520,N_3496);
and U8468 (N_8468,N_1941,N_2232);
or U8469 (N_8469,N_2144,N_3895);
nor U8470 (N_8470,N_4201,N_2928);
nand U8471 (N_8471,N_694,N_610);
or U8472 (N_8472,N_3636,N_673);
nand U8473 (N_8473,N_2394,N_2850);
and U8474 (N_8474,N_3615,N_4313);
and U8475 (N_8475,N_2826,N_2427);
xnor U8476 (N_8476,N_1014,N_2310);
xor U8477 (N_8477,N_2672,N_340);
nand U8478 (N_8478,N_3448,N_4062);
or U8479 (N_8479,N_3228,N_2032);
or U8480 (N_8480,N_2538,N_2046);
nand U8481 (N_8481,N_2991,N_1505);
xor U8482 (N_8482,N_1327,N_2050);
xnor U8483 (N_8483,N_2581,N_4797);
nand U8484 (N_8484,N_447,N_1601);
or U8485 (N_8485,N_440,N_894);
xnor U8486 (N_8486,N_4914,N_3089);
nand U8487 (N_8487,N_3508,N_3404);
xor U8488 (N_8488,N_864,N_2032);
nand U8489 (N_8489,N_2242,N_2231);
or U8490 (N_8490,N_4908,N_4077);
nor U8491 (N_8491,N_14,N_3472);
or U8492 (N_8492,N_135,N_3811);
xnor U8493 (N_8493,N_4953,N_3317);
nor U8494 (N_8494,N_94,N_1626);
xnor U8495 (N_8495,N_1150,N_612);
nor U8496 (N_8496,N_3457,N_605);
xnor U8497 (N_8497,N_1713,N_3971);
xnor U8498 (N_8498,N_4776,N_945);
xnor U8499 (N_8499,N_1069,N_342);
or U8500 (N_8500,N_500,N_2637);
xor U8501 (N_8501,N_611,N_130);
nand U8502 (N_8502,N_3046,N_2843);
nor U8503 (N_8503,N_2605,N_1588);
nor U8504 (N_8504,N_1382,N_4144);
nor U8505 (N_8505,N_822,N_2549);
xor U8506 (N_8506,N_4258,N_2100);
and U8507 (N_8507,N_3049,N_2346);
xnor U8508 (N_8508,N_1228,N_123);
xnor U8509 (N_8509,N_4437,N_904);
xnor U8510 (N_8510,N_4564,N_1341);
nor U8511 (N_8511,N_4336,N_4477);
and U8512 (N_8512,N_4517,N_421);
nor U8513 (N_8513,N_4437,N_346);
xnor U8514 (N_8514,N_4125,N_4695);
or U8515 (N_8515,N_1587,N_2151);
and U8516 (N_8516,N_262,N_1544);
nand U8517 (N_8517,N_4407,N_3109);
or U8518 (N_8518,N_3975,N_2131);
xor U8519 (N_8519,N_3652,N_4058);
and U8520 (N_8520,N_3434,N_2260);
and U8521 (N_8521,N_4664,N_1574);
nand U8522 (N_8522,N_2977,N_908);
nand U8523 (N_8523,N_3236,N_2084);
nand U8524 (N_8524,N_3351,N_1797);
and U8525 (N_8525,N_1014,N_2094);
and U8526 (N_8526,N_3927,N_3417);
and U8527 (N_8527,N_2687,N_3866);
or U8528 (N_8528,N_1244,N_4401);
nand U8529 (N_8529,N_1780,N_1977);
xnor U8530 (N_8530,N_1882,N_2555);
and U8531 (N_8531,N_3941,N_4543);
xor U8532 (N_8532,N_2845,N_664);
or U8533 (N_8533,N_179,N_574);
xnor U8534 (N_8534,N_426,N_2372);
and U8535 (N_8535,N_2555,N_2968);
nand U8536 (N_8536,N_1119,N_4209);
nor U8537 (N_8537,N_4959,N_1938);
or U8538 (N_8538,N_13,N_4252);
and U8539 (N_8539,N_2996,N_4716);
nor U8540 (N_8540,N_987,N_1568);
xnor U8541 (N_8541,N_2872,N_1463);
nand U8542 (N_8542,N_1602,N_1775);
nand U8543 (N_8543,N_4240,N_2150);
xor U8544 (N_8544,N_4205,N_4152);
and U8545 (N_8545,N_4434,N_276);
xnor U8546 (N_8546,N_3742,N_1289);
nand U8547 (N_8547,N_2652,N_4650);
and U8548 (N_8548,N_2538,N_3080);
and U8549 (N_8549,N_3405,N_1976);
nor U8550 (N_8550,N_2982,N_3188);
xnor U8551 (N_8551,N_1104,N_1132);
xor U8552 (N_8552,N_3620,N_727);
xor U8553 (N_8553,N_707,N_4783);
and U8554 (N_8554,N_1775,N_726);
or U8555 (N_8555,N_3305,N_4772);
nand U8556 (N_8556,N_257,N_578);
xor U8557 (N_8557,N_2991,N_534);
or U8558 (N_8558,N_2452,N_2610);
or U8559 (N_8559,N_3028,N_1064);
xnor U8560 (N_8560,N_4968,N_2959);
or U8561 (N_8561,N_4569,N_231);
nand U8562 (N_8562,N_1091,N_1830);
nor U8563 (N_8563,N_4320,N_4330);
nor U8564 (N_8564,N_2879,N_1862);
and U8565 (N_8565,N_1837,N_333);
xnor U8566 (N_8566,N_1236,N_4313);
nor U8567 (N_8567,N_1327,N_532);
nand U8568 (N_8568,N_2186,N_942);
and U8569 (N_8569,N_3112,N_2410);
nand U8570 (N_8570,N_2766,N_396);
or U8571 (N_8571,N_2027,N_1626);
or U8572 (N_8572,N_486,N_309);
and U8573 (N_8573,N_787,N_605);
and U8574 (N_8574,N_4484,N_2598);
and U8575 (N_8575,N_3213,N_3911);
or U8576 (N_8576,N_1435,N_4960);
or U8577 (N_8577,N_142,N_4382);
xnor U8578 (N_8578,N_144,N_1524);
nor U8579 (N_8579,N_2188,N_3176);
nor U8580 (N_8580,N_4173,N_455);
nand U8581 (N_8581,N_4744,N_3349);
or U8582 (N_8582,N_3558,N_2227);
or U8583 (N_8583,N_1211,N_334);
xnor U8584 (N_8584,N_4715,N_262);
nand U8585 (N_8585,N_1253,N_4311);
xnor U8586 (N_8586,N_4652,N_3041);
nor U8587 (N_8587,N_890,N_2136);
nor U8588 (N_8588,N_2661,N_4796);
xnor U8589 (N_8589,N_2858,N_4190);
and U8590 (N_8590,N_322,N_1612);
nor U8591 (N_8591,N_4243,N_3788);
xor U8592 (N_8592,N_3390,N_136);
nand U8593 (N_8593,N_4390,N_1481);
nor U8594 (N_8594,N_1038,N_4111);
or U8595 (N_8595,N_3621,N_3883);
or U8596 (N_8596,N_1456,N_4652);
nand U8597 (N_8597,N_2205,N_3118);
xnor U8598 (N_8598,N_4373,N_2823);
or U8599 (N_8599,N_856,N_4396);
and U8600 (N_8600,N_326,N_1372);
and U8601 (N_8601,N_1608,N_1462);
and U8602 (N_8602,N_2111,N_1595);
nor U8603 (N_8603,N_3588,N_437);
nand U8604 (N_8604,N_4633,N_1308);
and U8605 (N_8605,N_3895,N_4432);
xor U8606 (N_8606,N_3490,N_1256);
nand U8607 (N_8607,N_3873,N_3307);
and U8608 (N_8608,N_1766,N_935);
and U8609 (N_8609,N_1239,N_3024);
nand U8610 (N_8610,N_2116,N_4675);
nand U8611 (N_8611,N_2018,N_815);
xnor U8612 (N_8612,N_3534,N_667);
nand U8613 (N_8613,N_4824,N_3032);
and U8614 (N_8614,N_4382,N_1376);
or U8615 (N_8615,N_64,N_1733);
and U8616 (N_8616,N_4177,N_111);
xnor U8617 (N_8617,N_2865,N_3227);
nor U8618 (N_8618,N_2091,N_3276);
and U8619 (N_8619,N_1266,N_83);
nor U8620 (N_8620,N_806,N_2324);
and U8621 (N_8621,N_4255,N_4005);
or U8622 (N_8622,N_53,N_4529);
xor U8623 (N_8623,N_1828,N_1415);
nand U8624 (N_8624,N_3191,N_3125);
or U8625 (N_8625,N_1510,N_469);
nor U8626 (N_8626,N_2223,N_2620);
xor U8627 (N_8627,N_3597,N_373);
xnor U8628 (N_8628,N_2777,N_3367);
and U8629 (N_8629,N_4637,N_3250);
or U8630 (N_8630,N_2053,N_74);
and U8631 (N_8631,N_2687,N_3037);
and U8632 (N_8632,N_840,N_689);
xor U8633 (N_8633,N_703,N_4312);
or U8634 (N_8634,N_2695,N_4299);
and U8635 (N_8635,N_2492,N_57);
nand U8636 (N_8636,N_494,N_1358);
nor U8637 (N_8637,N_2573,N_3777);
and U8638 (N_8638,N_1207,N_2530);
or U8639 (N_8639,N_1923,N_3669);
nand U8640 (N_8640,N_4665,N_4212);
xnor U8641 (N_8641,N_717,N_4441);
or U8642 (N_8642,N_4698,N_542);
nor U8643 (N_8643,N_1547,N_513);
nand U8644 (N_8644,N_1177,N_2607);
nor U8645 (N_8645,N_4532,N_1379);
nand U8646 (N_8646,N_357,N_1324);
nor U8647 (N_8647,N_886,N_4699);
nand U8648 (N_8648,N_2695,N_2748);
xor U8649 (N_8649,N_4119,N_135);
and U8650 (N_8650,N_1421,N_3567);
or U8651 (N_8651,N_612,N_2232);
xnor U8652 (N_8652,N_3649,N_839);
nor U8653 (N_8653,N_2571,N_2378);
xor U8654 (N_8654,N_1772,N_308);
and U8655 (N_8655,N_969,N_1801);
or U8656 (N_8656,N_3146,N_76);
and U8657 (N_8657,N_2227,N_1209);
nor U8658 (N_8658,N_1235,N_1136);
or U8659 (N_8659,N_4932,N_1144);
nor U8660 (N_8660,N_4869,N_1643);
and U8661 (N_8661,N_997,N_2674);
nand U8662 (N_8662,N_1059,N_401);
or U8663 (N_8663,N_3044,N_4418);
nor U8664 (N_8664,N_146,N_2617);
nor U8665 (N_8665,N_2248,N_20);
xor U8666 (N_8666,N_1674,N_2951);
nand U8667 (N_8667,N_4787,N_3236);
nand U8668 (N_8668,N_4206,N_112);
xnor U8669 (N_8669,N_478,N_1683);
nor U8670 (N_8670,N_936,N_2771);
nand U8671 (N_8671,N_4483,N_1970);
nor U8672 (N_8672,N_1637,N_1425);
xnor U8673 (N_8673,N_1937,N_2270);
and U8674 (N_8674,N_1218,N_523);
nand U8675 (N_8675,N_409,N_1734);
and U8676 (N_8676,N_2761,N_334);
or U8677 (N_8677,N_3087,N_780);
xnor U8678 (N_8678,N_1577,N_2587);
nand U8679 (N_8679,N_3989,N_3084);
nor U8680 (N_8680,N_1164,N_1556);
nor U8681 (N_8681,N_599,N_4777);
and U8682 (N_8682,N_405,N_4229);
nor U8683 (N_8683,N_765,N_2064);
and U8684 (N_8684,N_4453,N_1576);
nand U8685 (N_8685,N_3297,N_3749);
nor U8686 (N_8686,N_3609,N_4684);
or U8687 (N_8687,N_3539,N_1007);
xor U8688 (N_8688,N_386,N_165);
nand U8689 (N_8689,N_1279,N_3839);
xnor U8690 (N_8690,N_2119,N_1799);
and U8691 (N_8691,N_1315,N_2408);
nand U8692 (N_8692,N_3399,N_707);
xnor U8693 (N_8693,N_2960,N_4628);
and U8694 (N_8694,N_714,N_3046);
and U8695 (N_8695,N_203,N_3353);
and U8696 (N_8696,N_4968,N_4339);
or U8697 (N_8697,N_960,N_3912);
nand U8698 (N_8698,N_3925,N_2406);
or U8699 (N_8699,N_854,N_2268);
or U8700 (N_8700,N_559,N_1182);
and U8701 (N_8701,N_4826,N_2215);
nand U8702 (N_8702,N_4499,N_4540);
xnor U8703 (N_8703,N_535,N_129);
or U8704 (N_8704,N_3751,N_953);
or U8705 (N_8705,N_2797,N_2432);
nand U8706 (N_8706,N_4349,N_3373);
nand U8707 (N_8707,N_4724,N_1212);
nor U8708 (N_8708,N_4996,N_2677);
and U8709 (N_8709,N_931,N_1759);
xor U8710 (N_8710,N_4336,N_318);
xnor U8711 (N_8711,N_3200,N_2501);
and U8712 (N_8712,N_3935,N_159);
nand U8713 (N_8713,N_4123,N_4128);
or U8714 (N_8714,N_1377,N_4662);
xor U8715 (N_8715,N_1739,N_4464);
and U8716 (N_8716,N_3586,N_2656);
nand U8717 (N_8717,N_4698,N_3710);
and U8718 (N_8718,N_2700,N_3481);
and U8719 (N_8719,N_4609,N_85);
and U8720 (N_8720,N_4825,N_1987);
nand U8721 (N_8721,N_4250,N_2734);
nand U8722 (N_8722,N_1662,N_2690);
nand U8723 (N_8723,N_1646,N_4647);
xnor U8724 (N_8724,N_2593,N_2014);
xnor U8725 (N_8725,N_4062,N_1463);
nand U8726 (N_8726,N_2623,N_2039);
xnor U8727 (N_8727,N_3338,N_1941);
nand U8728 (N_8728,N_2735,N_673);
or U8729 (N_8729,N_4975,N_4870);
nor U8730 (N_8730,N_1437,N_3184);
nand U8731 (N_8731,N_3669,N_726);
xnor U8732 (N_8732,N_1657,N_3138);
xnor U8733 (N_8733,N_3877,N_466);
xor U8734 (N_8734,N_483,N_4362);
xnor U8735 (N_8735,N_293,N_778);
nand U8736 (N_8736,N_892,N_2290);
nor U8737 (N_8737,N_3062,N_1206);
nor U8738 (N_8738,N_3961,N_4462);
xor U8739 (N_8739,N_3676,N_4656);
or U8740 (N_8740,N_4845,N_810);
nor U8741 (N_8741,N_2009,N_524);
or U8742 (N_8742,N_3409,N_1474);
or U8743 (N_8743,N_4401,N_1710);
nand U8744 (N_8744,N_557,N_4732);
or U8745 (N_8745,N_4678,N_107);
or U8746 (N_8746,N_1147,N_2960);
and U8747 (N_8747,N_2352,N_4167);
nor U8748 (N_8748,N_3445,N_354);
and U8749 (N_8749,N_2965,N_1872);
nor U8750 (N_8750,N_4381,N_3438);
or U8751 (N_8751,N_1283,N_3685);
nand U8752 (N_8752,N_2913,N_2686);
nand U8753 (N_8753,N_600,N_2815);
nor U8754 (N_8754,N_3390,N_3615);
nand U8755 (N_8755,N_4689,N_3758);
nor U8756 (N_8756,N_2255,N_2109);
or U8757 (N_8757,N_558,N_864);
xor U8758 (N_8758,N_1658,N_2979);
nor U8759 (N_8759,N_3214,N_3504);
and U8760 (N_8760,N_637,N_1735);
and U8761 (N_8761,N_177,N_1682);
xnor U8762 (N_8762,N_3794,N_1531);
xnor U8763 (N_8763,N_3519,N_2696);
nand U8764 (N_8764,N_4652,N_1334);
xor U8765 (N_8765,N_4057,N_766);
nor U8766 (N_8766,N_2697,N_1296);
or U8767 (N_8767,N_1586,N_1437);
nor U8768 (N_8768,N_1945,N_641);
and U8769 (N_8769,N_674,N_4717);
nand U8770 (N_8770,N_3510,N_1984);
xor U8771 (N_8771,N_1902,N_4360);
nor U8772 (N_8772,N_1371,N_1792);
or U8773 (N_8773,N_441,N_1610);
and U8774 (N_8774,N_2672,N_3991);
nor U8775 (N_8775,N_2565,N_3325);
nor U8776 (N_8776,N_619,N_953);
nor U8777 (N_8777,N_4390,N_525);
nand U8778 (N_8778,N_159,N_842);
and U8779 (N_8779,N_2402,N_1062);
nand U8780 (N_8780,N_2001,N_3641);
nor U8781 (N_8781,N_4750,N_3267);
nor U8782 (N_8782,N_4981,N_11);
and U8783 (N_8783,N_4120,N_678);
nand U8784 (N_8784,N_1939,N_3353);
nor U8785 (N_8785,N_28,N_1057);
or U8786 (N_8786,N_4921,N_1051);
nand U8787 (N_8787,N_3867,N_774);
or U8788 (N_8788,N_296,N_259);
or U8789 (N_8789,N_4755,N_4006);
and U8790 (N_8790,N_2690,N_3118);
nand U8791 (N_8791,N_1510,N_1442);
nand U8792 (N_8792,N_4688,N_2590);
or U8793 (N_8793,N_729,N_1449);
or U8794 (N_8794,N_3461,N_2817);
nor U8795 (N_8795,N_1259,N_313);
nand U8796 (N_8796,N_489,N_119);
nor U8797 (N_8797,N_3404,N_1851);
nor U8798 (N_8798,N_4361,N_3778);
nand U8799 (N_8799,N_2848,N_4935);
nor U8800 (N_8800,N_2822,N_4638);
and U8801 (N_8801,N_1752,N_1418);
or U8802 (N_8802,N_1730,N_2761);
or U8803 (N_8803,N_840,N_3267);
and U8804 (N_8804,N_757,N_2474);
nand U8805 (N_8805,N_4505,N_1088);
and U8806 (N_8806,N_2164,N_275);
nand U8807 (N_8807,N_2468,N_102);
nor U8808 (N_8808,N_1518,N_1630);
nand U8809 (N_8809,N_4926,N_888);
nand U8810 (N_8810,N_3245,N_3045);
or U8811 (N_8811,N_1042,N_2675);
nor U8812 (N_8812,N_3073,N_4341);
xnor U8813 (N_8813,N_4367,N_3219);
nand U8814 (N_8814,N_2596,N_826);
or U8815 (N_8815,N_750,N_3870);
and U8816 (N_8816,N_893,N_819);
or U8817 (N_8817,N_622,N_1564);
xnor U8818 (N_8818,N_1518,N_4717);
nor U8819 (N_8819,N_678,N_4487);
xnor U8820 (N_8820,N_4965,N_4549);
nor U8821 (N_8821,N_4581,N_1361);
or U8822 (N_8822,N_3469,N_3893);
xnor U8823 (N_8823,N_3517,N_4385);
and U8824 (N_8824,N_1732,N_4931);
nor U8825 (N_8825,N_2502,N_884);
nor U8826 (N_8826,N_2704,N_2594);
xnor U8827 (N_8827,N_2666,N_3191);
nor U8828 (N_8828,N_1852,N_2387);
nor U8829 (N_8829,N_3958,N_2414);
nor U8830 (N_8830,N_2016,N_2257);
and U8831 (N_8831,N_4537,N_1634);
nand U8832 (N_8832,N_592,N_390);
and U8833 (N_8833,N_1512,N_1265);
or U8834 (N_8834,N_3059,N_1069);
and U8835 (N_8835,N_3437,N_4479);
or U8836 (N_8836,N_297,N_2623);
nor U8837 (N_8837,N_4990,N_3550);
nand U8838 (N_8838,N_1403,N_4257);
nand U8839 (N_8839,N_1173,N_1141);
and U8840 (N_8840,N_169,N_1165);
nand U8841 (N_8841,N_1435,N_49);
nor U8842 (N_8842,N_296,N_3435);
xnor U8843 (N_8843,N_624,N_2876);
nand U8844 (N_8844,N_3985,N_2693);
or U8845 (N_8845,N_2371,N_2713);
or U8846 (N_8846,N_1916,N_614);
nor U8847 (N_8847,N_4522,N_2176);
and U8848 (N_8848,N_3827,N_2389);
nand U8849 (N_8849,N_3156,N_3745);
or U8850 (N_8850,N_3493,N_1208);
xor U8851 (N_8851,N_1074,N_4685);
nor U8852 (N_8852,N_1535,N_3937);
nor U8853 (N_8853,N_2650,N_4068);
nand U8854 (N_8854,N_3616,N_4274);
and U8855 (N_8855,N_1517,N_2547);
and U8856 (N_8856,N_1956,N_2297);
nor U8857 (N_8857,N_385,N_4422);
nand U8858 (N_8858,N_2549,N_4986);
nand U8859 (N_8859,N_3860,N_879);
and U8860 (N_8860,N_6,N_1283);
or U8861 (N_8861,N_3591,N_3036);
nand U8862 (N_8862,N_4319,N_4441);
nand U8863 (N_8863,N_2748,N_4805);
and U8864 (N_8864,N_1439,N_34);
nor U8865 (N_8865,N_3813,N_3855);
nand U8866 (N_8866,N_314,N_2805);
xnor U8867 (N_8867,N_2473,N_1193);
xor U8868 (N_8868,N_3190,N_1848);
nor U8869 (N_8869,N_3269,N_2808);
and U8870 (N_8870,N_4224,N_506);
xor U8871 (N_8871,N_2361,N_1069);
or U8872 (N_8872,N_2873,N_1979);
and U8873 (N_8873,N_2178,N_3005);
xnor U8874 (N_8874,N_3945,N_1648);
and U8875 (N_8875,N_1365,N_2526);
or U8876 (N_8876,N_2906,N_620);
and U8877 (N_8877,N_2009,N_4469);
nand U8878 (N_8878,N_916,N_3761);
nand U8879 (N_8879,N_2210,N_1460);
xor U8880 (N_8880,N_3976,N_1954);
or U8881 (N_8881,N_16,N_1214);
nand U8882 (N_8882,N_1915,N_4791);
nand U8883 (N_8883,N_85,N_4446);
nor U8884 (N_8884,N_3246,N_4665);
nand U8885 (N_8885,N_892,N_1397);
nor U8886 (N_8886,N_2791,N_3787);
xor U8887 (N_8887,N_1416,N_4800);
or U8888 (N_8888,N_1509,N_1204);
xor U8889 (N_8889,N_2859,N_1632);
and U8890 (N_8890,N_4199,N_593);
or U8891 (N_8891,N_2799,N_605);
nor U8892 (N_8892,N_2631,N_1505);
nand U8893 (N_8893,N_4781,N_962);
xnor U8894 (N_8894,N_1920,N_489);
xor U8895 (N_8895,N_2558,N_269);
or U8896 (N_8896,N_1896,N_1693);
xnor U8897 (N_8897,N_412,N_4844);
nand U8898 (N_8898,N_2380,N_1476);
nand U8899 (N_8899,N_2509,N_543);
nor U8900 (N_8900,N_3804,N_137);
xor U8901 (N_8901,N_2590,N_1529);
nor U8902 (N_8902,N_920,N_1156);
or U8903 (N_8903,N_2975,N_2689);
and U8904 (N_8904,N_65,N_4064);
and U8905 (N_8905,N_197,N_2233);
and U8906 (N_8906,N_358,N_1360);
nand U8907 (N_8907,N_3252,N_4944);
nand U8908 (N_8908,N_436,N_1304);
and U8909 (N_8909,N_1874,N_3125);
nor U8910 (N_8910,N_191,N_4456);
nor U8911 (N_8911,N_2900,N_2451);
and U8912 (N_8912,N_3715,N_4703);
or U8913 (N_8913,N_2282,N_3499);
or U8914 (N_8914,N_2330,N_96);
or U8915 (N_8915,N_4159,N_1703);
or U8916 (N_8916,N_3003,N_4689);
nor U8917 (N_8917,N_4173,N_1867);
nand U8918 (N_8918,N_2295,N_4172);
nor U8919 (N_8919,N_189,N_1755);
and U8920 (N_8920,N_603,N_596);
nor U8921 (N_8921,N_2846,N_158);
nor U8922 (N_8922,N_669,N_988);
nand U8923 (N_8923,N_3287,N_3680);
or U8924 (N_8924,N_4919,N_1190);
xnor U8925 (N_8925,N_3876,N_815);
xor U8926 (N_8926,N_4381,N_3117);
nor U8927 (N_8927,N_4152,N_923);
nand U8928 (N_8928,N_3108,N_4670);
or U8929 (N_8929,N_2581,N_780);
xor U8930 (N_8930,N_293,N_226);
xnor U8931 (N_8931,N_857,N_9);
nand U8932 (N_8932,N_3592,N_1505);
nor U8933 (N_8933,N_3291,N_4448);
nor U8934 (N_8934,N_3271,N_153);
nand U8935 (N_8935,N_1521,N_4791);
xnor U8936 (N_8936,N_4495,N_1933);
or U8937 (N_8937,N_3277,N_1910);
or U8938 (N_8938,N_3122,N_4166);
nor U8939 (N_8939,N_530,N_3080);
nand U8940 (N_8940,N_334,N_1609);
nor U8941 (N_8941,N_1068,N_407);
or U8942 (N_8942,N_923,N_3284);
nor U8943 (N_8943,N_2748,N_3795);
and U8944 (N_8944,N_4344,N_4864);
or U8945 (N_8945,N_1933,N_1164);
xor U8946 (N_8946,N_3217,N_545);
xor U8947 (N_8947,N_315,N_1490);
or U8948 (N_8948,N_885,N_4034);
or U8949 (N_8949,N_2223,N_659);
nand U8950 (N_8950,N_1868,N_2184);
xor U8951 (N_8951,N_4262,N_4837);
xnor U8952 (N_8952,N_3427,N_1499);
nand U8953 (N_8953,N_4833,N_3980);
or U8954 (N_8954,N_4925,N_2606);
xnor U8955 (N_8955,N_4667,N_2007);
or U8956 (N_8956,N_3785,N_4677);
or U8957 (N_8957,N_1374,N_4503);
and U8958 (N_8958,N_671,N_4129);
nand U8959 (N_8959,N_4971,N_647);
nand U8960 (N_8960,N_1190,N_390);
nand U8961 (N_8961,N_3425,N_939);
and U8962 (N_8962,N_2985,N_4243);
xor U8963 (N_8963,N_276,N_4835);
xnor U8964 (N_8964,N_1956,N_4734);
or U8965 (N_8965,N_4960,N_1514);
or U8966 (N_8966,N_1466,N_4653);
nor U8967 (N_8967,N_2844,N_1733);
or U8968 (N_8968,N_4793,N_325);
nor U8969 (N_8969,N_4697,N_4828);
xor U8970 (N_8970,N_706,N_164);
and U8971 (N_8971,N_1910,N_392);
xnor U8972 (N_8972,N_611,N_3573);
or U8973 (N_8973,N_4234,N_2118);
xnor U8974 (N_8974,N_1123,N_1228);
xor U8975 (N_8975,N_1114,N_3401);
xor U8976 (N_8976,N_2268,N_56);
nor U8977 (N_8977,N_3322,N_1569);
nor U8978 (N_8978,N_1656,N_2182);
or U8979 (N_8979,N_3483,N_1344);
nand U8980 (N_8980,N_4466,N_4838);
or U8981 (N_8981,N_3555,N_4212);
nand U8982 (N_8982,N_1487,N_4188);
nor U8983 (N_8983,N_2269,N_4329);
nor U8984 (N_8984,N_1011,N_4119);
nand U8985 (N_8985,N_1362,N_2738);
xor U8986 (N_8986,N_660,N_2136);
nand U8987 (N_8987,N_517,N_4254);
nor U8988 (N_8988,N_822,N_2651);
nor U8989 (N_8989,N_1271,N_1398);
nand U8990 (N_8990,N_3049,N_3685);
xor U8991 (N_8991,N_4356,N_4702);
nand U8992 (N_8992,N_1955,N_843);
xor U8993 (N_8993,N_3235,N_211);
nand U8994 (N_8994,N_2473,N_3383);
nand U8995 (N_8995,N_2505,N_4023);
nand U8996 (N_8996,N_4515,N_3273);
nor U8997 (N_8997,N_4433,N_2568);
or U8998 (N_8998,N_2393,N_1823);
or U8999 (N_8999,N_596,N_3391);
and U9000 (N_9000,N_2019,N_1375);
xor U9001 (N_9001,N_941,N_3850);
nand U9002 (N_9002,N_4784,N_4485);
nand U9003 (N_9003,N_2901,N_3135);
nor U9004 (N_9004,N_4385,N_953);
nor U9005 (N_9005,N_3022,N_85);
nor U9006 (N_9006,N_2712,N_3478);
nor U9007 (N_9007,N_1411,N_2212);
and U9008 (N_9008,N_1687,N_2645);
xnor U9009 (N_9009,N_3771,N_3325);
or U9010 (N_9010,N_3375,N_306);
xnor U9011 (N_9011,N_1688,N_3694);
xor U9012 (N_9012,N_1131,N_734);
nor U9013 (N_9013,N_2882,N_935);
nand U9014 (N_9014,N_971,N_391);
or U9015 (N_9015,N_4073,N_2555);
or U9016 (N_9016,N_843,N_3884);
nor U9017 (N_9017,N_4370,N_3640);
nor U9018 (N_9018,N_91,N_288);
or U9019 (N_9019,N_425,N_2487);
and U9020 (N_9020,N_442,N_3107);
and U9021 (N_9021,N_1509,N_508);
xor U9022 (N_9022,N_124,N_3672);
nor U9023 (N_9023,N_1956,N_1361);
nor U9024 (N_9024,N_1843,N_4476);
nor U9025 (N_9025,N_2563,N_1243);
nand U9026 (N_9026,N_2625,N_1715);
xnor U9027 (N_9027,N_3795,N_3586);
or U9028 (N_9028,N_2225,N_2792);
and U9029 (N_9029,N_3922,N_4804);
nand U9030 (N_9030,N_1839,N_2510);
or U9031 (N_9031,N_2161,N_3963);
nand U9032 (N_9032,N_4653,N_3216);
or U9033 (N_9033,N_1002,N_3328);
nand U9034 (N_9034,N_3331,N_4507);
nand U9035 (N_9035,N_4487,N_785);
or U9036 (N_9036,N_2091,N_2173);
or U9037 (N_9037,N_2681,N_1198);
and U9038 (N_9038,N_1089,N_2227);
nor U9039 (N_9039,N_2513,N_4420);
and U9040 (N_9040,N_3234,N_657);
xnor U9041 (N_9041,N_2561,N_1170);
nor U9042 (N_9042,N_1109,N_3900);
xor U9043 (N_9043,N_3174,N_4675);
nor U9044 (N_9044,N_2909,N_4415);
or U9045 (N_9045,N_3334,N_324);
nor U9046 (N_9046,N_1223,N_1797);
xor U9047 (N_9047,N_1111,N_1884);
xnor U9048 (N_9048,N_411,N_3590);
and U9049 (N_9049,N_3600,N_3405);
nand U9050 (N_9050,N_3787,N_3144);
and U9051 (N_9051,N_4817,N_4728);
and U9052 (N_9052,N_2491,N_1624);
nand U9053 (N_9053,N_4642,N_2786);
or U9054 (N_9054,N_3790,N_1946);
or U9055 (N_9055,N_4837,N_3709);
nor U9056 (N_9056,N_1849,N_508);
or U9057 (N_9057,N_2434,N_2533);
xor U9058 (N_9058,N_51,N_687);
nor U9059 (N_9059,N_1717,N_3405);
nor U9060 (N_9060,N_2117,N_3741);
or U9061 (N_9061,N_1216,N_1851);
nand U9062 (N_9062,N_4544,N_4057);
xnor U9063 (N_9063,N_2945,N_3143);
xor U9064 (N_9064,N_214,N_3406);
and U9065 (N_9065,N_3211,N_455);
or U9066 (N_9066,N_3563,N_1048);
and U9067 (N_9067,N_2722,N_1803);
or U9068 (N_9068,N_3329,N_3557);
and U9069 (N_9069,N_1167,N_18);
nand U9070 (N_9070,N_1452,N_2165);
nand U9071 (N_9071,N_274,N_507);
xnor U9072 (N_9072,N_2490,N_3768);
or U9073 (N_9073,N_3171,N_4626);
nand U9074 (N_9074,N_3838,N_519);
nor U9075 (N_9075,N_111,N_3746);
or U9076 (N_9076,N_1104,N_3296);
nor U9077 (N_9077,N_827,N_3119);
or U9078 (N_9078,N_2830,N_4836);
and U9079 (N_9079,N_4081,N_2058);
nor U9080 (N_9080,N_31,N_2601);
nand U9081 (N_9081,N_1187,N_98);
xor U9082 (N_9082,N_2688,N_2129);
and U9083 (N_9083,N_4238,N_4267);
xnor U9084 (N_9084,N_2867,N_4551);
nor U9085 (N_9085,N_3149,N_681);
and U9086 (N_9086,N_4351,N_245);
nor U9087 (N_9087,N_242,N_4571);
and U9088 (N_9088,N_3387,N_3907);
or U9089 (N_9089,N_3726,N_2322);
or U9090 (N_9090,N_433,N_2584);
xnor U9091 (N_9091,N_4608,N_2267);
or U9092 (N_9092,N_3166,N_4540);
and U9093 (N_9093,N_815,N_2310);
nand U9094 (N_9094,N_2328,N_3617);
nand U9095 (N_9095,N_617,N_135);
nand U9096 (N_9096,N_4899,N_2483);
nand U9097 (N_9097,N_3851,N_1172);
nor U9098 (N_9098,N_3352,N_4332);
or U9099 (N_9099,N_2853,N_2199);
or U9100 (N_9100,N_3069,N_945);
nor U9101 (N_9101,N_3762,N_39);
nor U9102 (N_9102,N_4945,N_3200);
nor U9103 (N_9103,N_4586,N_1922);
xor U9104 (N_9104,N_143,N_20);
or U9105 (N_9105,N_3467,N_1255);
xor U9106 (N_9106,N_541,N_1781);
and U9107 (N_9107,N_3624,N_603);
or U9108 (N_9108,N_1134,N_855);
and U9109 (N_9109,N_4591,N_2282);
and U9110 (N_9110,N_504,N_1672);
nor U9111 (N_9111,N_3231,N_279);
xnor U9112 (N_9112,N_65,N_2853);
nand U9113 (N_9113,N_3178,N_2921);
xor U9114 (N_9114,N_4169,N_2343);
nand U9115 (N_9115,N_3701,N_713);
xor U9116 (N_9116,N_3864,N_642);
or U9117 (N_9117,N_3809,N_554);
and U9118 (N_9118,N_1277,N_4286);
xor U9119 (N_9119,N_681,N_2500);
nor U9120 (N_9120,N_4058,N_3648);
or U9121 (N_9121,N_604,N_1519);
or U9122 (N_9122,N_1548,N_3043);
nand U9123 (N_9123,N_501,N_1880);
or U9124 (N_9124,N_3200,N_4175);
and U9125 (N_9125,N_3105,N_1197);
and U9126 (N_9126,N_3364,N_2105);
nor U9127 (N_9127,N_888,N_2827);
nor U9128 (N_9128,N_1462,N_546);
or U9129 (N_9129,N_3969,N_3943);
nand U9130 (N_9130,N_2805,N_2215);
or U9131 (N_9131,N_3385,N_1231);
xor U9132 (N_9132,N_2862,N_2645);
nor U9133 (N_9133,N_4674,N_1310);
and U9134 (N_9134,N_4406,N_2099);
or U9135 (N_9135,N_3622,N_1227);
nor U9136 (N_9136,N_4630,N_279);
nand U9137 (N_9137,N_3354,N_2021);
xor U9138 (N_9138,N_4632,N_1271);
and U9139 (N_9139,N_248,N_1769);
xor U9140 (N_9140,N_2014,N_3505);
and U9141 (N_9141,N_605,N_2947);
and U9142 (N_9142,N_4711,N_532);
or U9143 (N_9143,N_837,N_4675);
or U9144 (N_9144,N_3147,N_3301);
or U9145 (N_9145,N_2648,N_3865);
or U9146 (N_9146,N_1331,N_4888);
or U9147 (N_9147,N_1510,N_4799);
xor U9148 (N_9148,N_684,N_4787);
xor U9149 (N_9149,N_19,N_209);
nor U9150 (N_9150,N_4266,N_4407);
nand U9151 (N_9151,N_3609,N_1658);
nor U9152 (N_9152,N_1458,N_1466);
nor U9153 (N_9153,N_1949,N_2400);
and U9154 (N_9154,N_4457,N_1547);
nor U9155 (N_9155,N_4479,N_4604);
nor U9156 (N_9156,N_654,N_2252);
nand U9157 (N_9157,N_3903,N_1944);
and U9158 (N_9158,N_4605,N_2378);
and U9159 (N_9159,N_2464,N_1314);
or U9160 (N_9160,N_4831,N_2246);
and U9161 (N_9161,N_2339,N_2221);
nor U9162 (N_9162,N_3794,N_371);
xnor U9163 (N_9163,N_4733,N_4265);
or U9164 (N_9164,N_2097,N_4337);
or U9165 (N_9165,N_637,N_2502);
and U9166 (N_9166,N_4037,N_2298);
xnor U9167 (N_9167,N_4016,N_210);
nand U9168 (N_9168,N_23,N_874);
nor U9169 (N_9169,N_0,N_4997);
xnor U9170 (N_9170,N_2029,N_4440);
and U9171 (N_9171,N_3545,N_1774);
xnor U9172 (N_9172,N_1578,N_1630);
nor U9173 (N_9173,N_3770,N_3486);
and U9174 (N_9174,N_82,N_789);
xor U9175 (N_9175,N_4527,N_4314);
xor U9176 (N_9176,N_1332,N_2771);
nor U9177 (N_9177,N_623,N_2757);
or U9178 (N_9178,N_3105,N_4767);
nand U9179 (N_9179,N_1684,N_3723);
nor U9180 (N_9180,N_2172,N_2019);
or U9181 (N_9181,N_2339,N_1092);
nor U9182 (N_9182,N_4109,N_1329);
and U9183 (N_9183,N_2682,N_1114);
nand U9184 (N_9184,N_2825,N_3256);
xnor U9185 (N_9185,N_922,N_4445);
or U9186 (N_9186,N_584,N_2263);
nor U9187 (N_9187,N_736,N_2532);
xor U9188 (N_9188,N_4679,N_3506);
and U9189 (N_9189,N_4764,N_1193);
nor U9190 (N_9190,N_3982,N_2711);
nand U9191 (N_9191,N_3460,N_2932);
or U9192 (N_9192,N_370,N_2163);
and U9193 (N_9193,N_1197,N_1616);
nand U9194 (N_9194,N_1263,N_2348);
and U9195 (N_9195,N_774,N_957);
and U9196 (N_9196,N_2022,N_3630);
xor U9197 (N_9197,N_579,N_2857);
nor U9198 (N_9198,N_690,N_2639);
xnor U9199 (N_9199,N_144,N_3160);
or U9200 (N_9200,N_3774,N_4622);
nand U9201 (N_9201,N_852,N_3264);
nor U9202 (N_9202,N_822,N_3931);
or U9203 (N_9203,N_3247,N_3206);
or U9204 (N_9204,N_4415,N_2914);
and U9205 (N_9205,N_1331,N_3250);
and U9206 (N_9206,N_1488,N_1872);
and U9207 (N_9207,N_624,N_1955);
nor U9208 (N_9208,N_127,N_3497);
or U9209 (N_9209,N_4156,N_4381);
nor U9210 (N_9210,N_1269,N_4547);
nand U9211 (N_9211,N_3486,N_4091);
nor U9212 (N_9212,N_3252,N_1256);
nand U9213 (N_9213,N_3851,N_3685);
or U9214 (N_9214,N_2146,N_4867);
nor U9215 (N_9215,N_2103,N_4300);
nor U9216 (N_9216,N_2034,N_3909);
xor U9217 (N_9217,N_2006,N_4985);
or U9218 (N_9218,N_2277,N_1952);
nand U9219 (N_9219,N_1819,N_1617);
xor U9220 (N_9220,N_3193,N_788);
or U9221 (N_9221,N_3322,N_2322);
nor U9222 (N_9222,N_970,N_1776);
and U9223 (N_9223,N_1577,N_3533);
and U9224 (N_9224,N_455,N_4694);
nand U9225 (N_9225,N_618,N_2924);
or U9226 (N_9226,N_2853,N_4489);
and U9227 (N_9227,N_892,N_2708);
xnor U9228 (N_9228,N_2571,N_2691);
nor U9229 (N_9229,N_1084,N_2056);
and U9230 (N_9230,N_376,N_3449);
nor U9231 (N_9231,N_3277,N_2084);
nand U9232 (N_9232,N_219,N_4269);
nand U9233 (N_9233,N_4102,N_2756);
nand U9234 (N_9234,N_2575,N_4315);
and U9235 (N_9235,N_2410,N_1149);
xor U9236 (N_9236,N_129,N_4993);
nand U9237 (N_9237,N_4789,N_2316);
or U9238 (N_9238,N_2384,N_4190);
nand U9239 (N_9239,N_1840,N_1423);
xor U9240 (N_9240,N_1881,N_3018);
or U9241 (N_9241,N_3064,N_2204);
or U9242 (N_9242,N_1216,N_2334);
nor U9243 (N_9243,N_432,N_1641);
xnor U9244 (N_9244,N_735,N_2236);
xor U9245 (N_9245,N_4008,N_1301);
or U9246 (N_9246,N_3809,N_1936);
xor U9247 (N_9247,N_3026,N_4780);
xnor U9248 (N_9248,N_2693,N_3280);
or U9249 (N_9249,N_2991,N_1648);
or U9250 (N_9250,N_2583,N_4045);
nor U9251 (N_9251,N_3985,N_3819);
nand U9252 (N_9252,N_3677,N_2240);
or U9253 (N_9253,N_4308,N_923);
nor U9254 (N_9254,N_182,N_4109);
nor U9255 (N_9255,N_1697,N_2531);
nor U9256 (N_9256,N_4160,N_4652);
or U9257 (N_9257,N_2046,N_3226);
nand U9258 (N_9258,N_2794,N_2245);
or U9259 (N_9259,N_2603,N_4433);
and U9260 (N_9260,N_2160,N_4709);
or U9261 (N_9261,N_4013,N_3981);
xnor U9262 (N_9262,N_388,N_1664);
and U9263 (N_9263,N_946,N_374);
nor U9264 (N_9264,N_2640,N_4138);
nand U9265 (N_9265,N_699,N_4538);
xor U9266 (N_9266,N_2675,N_4276);
nand U9267 (N_9267,N_3760,N_1988);
nor U9268 (N_9268,N_2938,N_3238);
nor U9269 (N_9269,N_2512,N_4777);
or U9270 (N_9270,N_4338,N_3450);
and U9271 (N_9271,N_1261,N_1684);
or U9272 (N_9272,N_3851,N_2705);
xor U9273 (N_9273,N_4275,N_998);
nor U9274 (N_9274,N_877,N_1887);
xor U9275 (N_9275,N_2893,N_3620);
xor U9276 (N_9276,N_657,N_1822);
or U9277 (N_9277,N_3311,N_4598);
nand U9278 (N_9278,N_365,N_728);
and U9279 (N_9279,N_101,N_3539);
nand U9280 (N_9280,N_1961,N_4351);
and U9281 (N_9281,N_4020,N_3198);
nand U9282 (N_9282,N_692,N_3045);
or U9283 (N_9283,N_2736,N_4192);
xor U9284 (N_9284,N_15,N_1563);
and U9285 (N_9285,N_2992,N_32);
or U9286 (N_9286,N_604,N_2015);
nand U9287 (N_9287,N_3230,N_3288);
and U9288 (N_9288,N_1927,N_1223);
and U9289 (N_9289,N_2225,N_3172);
nor U9290 (N_9290,N_4831,N_1087);
or U9291 (N_9291,N_2748,N_4787);
xor U9292 (N_9292,N_626,N_2161);
or U9293 (N_9293,N_2282,N_1559);
or U9294 (N_9294,N_2527,N_1817);
or U9295 (N_9295,N_52,N_119);
or U9296 (N_9296,N_2627,N_2553);
nor U9297 (N_9297,N_4871,N_2799);
or U9298 (N_9298,N_4252,N_2962);
nand U9299 (N_9299,N_1539,N_4610);
or U9300 (N_9300,N_2959,N_258);
xnor U9301 (N_9301,N_3381,N_650);
and U9302 (N_9302,N_4828,N_571);
xor U9303 (N_9303,N_3067,N_3070);
or U9304 (N_9304,N_208,N_2643);
or U9305 (N_9305,N_240,N_4935);
nor U9306 (N_9306,N_398,N_1045);
nand U9307 (N_9307,N_4488,N_443);
nand U9308 (N_9308,N_169,N_2023);
nand U9309 (N_9309,N_4898,N_794);
nand U9310 (N_9310,N_3312,N_4179);
nand U9311 (N_9311,N_869,N_3870);
xor U9312 (N_9312,N_2321,N_4733);
nand U9313 (N_9313,N_3200,N_2887);
nor U9314 (N_9314,N_4204,N_736);
xor U9315 (N_9315,N_882,N_436);
or U9316 (N_9316,N_3135,N_2508);
nand U9317 (N_9317,N_3183,N_2361);
nor U9318 (N_9318,N_1951,N_4344);
xnor U9319 (N_9319,N_770,N_2760);
or U9320 (N_9320,N_88,N_566);
xor U9321 (N_9321,N_249,N_1312);
and U9322 (N_9322,N_3175,N_4742);
and U9323 (N_9323,N_4470,N_642);
nand U9324 (N_9324,N_3172,N_3323);
nor U9325 (N_9325,N_349,N_380);
and U9326 (N_9326,N_104,N_1302);
and U9327 (N_9327,N_58,N_4109);
and U9328 (N_9328,N_2975,N_1725);
or U9329 (N_9329,N_1373,N_4836);
nand U9330 (N_9330,N_3345,N_3185);
nor U9331 (N_9331,N_4855,N_3274);
nor U9332 (N_9332,N_532,N_1672);
xor U9333 (N_9333,N_2230,N_1392);
or U9334 (N_9334,N_3903,N_3105);
xnor U9335 (N_9335,N_1495,N_3440);
nand U9336 (N_9336,N_1113,N_578);
and U9337 (N_9337,N_2199,N_4197);
and U9338 (N_9338,N_4364,N_4028);
nor U9339 (N_9339,N_3243,N_802);
or U9340 (N_9340,N_3246,N_499);
or U9341 (N_9341,N_4834,N_342);
or U9342 (N_9342,N_2429,N_3476);
or U9343 (N_9343,N_297,N_3115);
xnor U9344 (N_9344,N_562,N_3949);
or U9345 (N_9345,N_4567,N_4094);
and U9346 (N_9346,N_1930,N_2746);
nor U9347 (N_9347,N_2347,N_3666);
or U9348 (N_9348,N_3810,N_4397);
nor U9349 (N_9349,N_1386,N_3511);
and U9350 (N_9350,N_950,N_140);
xor U9351 (N_9351,N_3205,N_1485);
nand U9352 (N_9352,N_3222,N_2244);
nand U9353 (N_9353,N_797,N_1840);
nor U9354 (N_9354,N_2168,N_4254);
nor U9355 (N_9355,N_2130,N_4258);
nor U9356 (N_9356,N_6,N_2636);
and U9357 (N_9357,N_122,N_419);
and U9358 (N_9358,N_2690,N_1213);
nand U9359 (N_9359,N_4722,N_4546);
nor U9360 (N_9360,N_4189,N_4079);
xnor U9361 (N_9361,N_2055,N_1889);
nand U9362 (N_9362,N_4256,N_2697);
xnor U9363 (N_9363,N_4157,N_4691);
nor U9364 (N_9364,N_4084,N_1466);
or U9365 (N_9365,N_4986,N_188);
xnor U9366 (N_9366,N_388,N_2403);
nand U9367 (N_9367,N_4011,N_1235);
nand U9368 (N_9368,N_2012,N_540);
xor U9369 (N_9369,N_4728,N_2082);
and U9370 (N_9370,N_1221,N_1913);
nand U9371 (N_9371,N_2202,N_1074);
and U9372 (N_9372,N_1339,N_4497);
nand U9373 (N_9373,N_3075,N_4075);
nand U9374 (N_9374,N_2604,N_989);
nor U9375 (N_9375,N_4430,N_523);
nand U9376 (N_9376,N_1121,N_3102);
nand U9377 (N_9377,N_4707,N_3992);
xnor U9378 (N_9378,N_4253,N_1963);
nand U9379 (N_9379,N_10,N_4088);
xnor U9380 (N_9380,N_4343,N_295);
xor U9381 (N_9381,N_2567,N_3909);
nand U9382 (N_9382,N_1220,N_2000);
and U9383 (N_9383,N_2151,N_1402);
or U9384 (N_9384,N_2394,N_3097);
nand U9385 (N_9385,N_1938,N_3756);
xnor U9386 (N_9386,N_2441,N_1860);
nor U9387 (N_9387,N_1814,N_1051);
nor U9388 (N_9388,N_796,N_1281);
and U9389 (N_9389,N_4539,N_1702);
nand U9390 (N_9390,N_2674,N_3842);
or U9391 (N_9391,N_3605,N_1652);
and U9392 (N_9392,N_1691,N_518);
nand U9393 (N_9393,N_646,N_4254);
xor U9394 (N_9394,N_77,N_2722);
xor U9395 (N_9395,N_395,N_1646);
xnor U9396 (N_9396,N_3250,N_1344);
nor U9397 (N_9397,N_1989,N_713);
and U9398 (N_9398,N_1665,N_2615);
xnor U9399 (N_9399,N_727,N_200);
or U9400 (N_9400,N_3731,N_1696);
nand U9401 (N_9401,N_613,N_42);
or U9402 (N_9402,N_2606,N_1907);
or U9403 (N_9403,N_4831,N_2796);
nand U9404 (N_9404,N_2863,N_3502);
nand U9405 (N_9405,N_4057,N_3059);
xor U9406 (N_9406,N_3777,N_1118);
nand U9407 (N_9407,N_88,N_1226);
nor U9408 (N_9408,N_4532,N_241);
or U9409 (N_9409,N_2334,N_3548);
nand U9410 (N_9410,N_3438,N_2754);
xnor U9411 (N_9411,N_2472,N_3860);
xor U9412 (N_9412,N_3370,N_3395);
or U9413 (N_9413,N_2777,N_14);
xnor U9414 (N_9414,N_4144,N_4293);
nand U9415 (N_9415,N_1393,N_2723);
nor U9416 (N_9416,N_87,N_501);
nand U9417 (N_9417,N_4220,N_1621);
or U9418 (N_9418,N_4261,N_1218);
nor U9419 (N_9419,N_3562,N_681);
and U9420 (N_9420,N_2134,N_225);
nor U9421 (N_9421,N_3366,N_4470);
and U9422 (N_9422,N_4978,N_2921);
and U9423 (N_9423,N_269,N_2130);
nor U9424 (N_9424,N_2155,N_238);
nand U9425 (N_9425,N_3777,N_4844);
nand U9426 (N_9426,N_50,N_1227);
nor U9427 (N_9427,N_3685,N_544);
nor U9428 (N_9428,N_270,N_4543);
nor U9429 (N_9429,N_2269,N_195);
nand U9430 (N_9430,N_452,N_373);
xor U9431 (N_9431,N_574,N_350);
or U9432 (N_9432,N_2204,N_2589);
or U9433 (N_9433,N_4655,N_1745);
nand U9434 (N_9434,N_2246,N_48);
xnor U9435 (N_9435,N_290,N_1670);
and U9436 (N_9436,N_158,N_4255);
and U9437 (N_9437,N_3516,N_1584);
or U9438 (N_9438,N_1486,N_1738);
and U9439 (N_9439,N_3735,N_3601);
nand U9440 (N_9440,N_4464,N_3109);
nor U9441 (N_9441,N_3501,N_3548);
xnor U9442 (N_9442,N_3421,N_735);
xnor U9443 (N_9443,N_4933,N_138);
or U9444 (N_9444,N_3459,N_2931);
and U9445 (N_9445,N_4015,N_3304);
nand U9446 (N_9446,N_647,N_3591);
xnor U9447 (N_9447,N_1618,N_1562);
or U9448 (N_9448,N_2395,N_2739);
xnor U9449 (N_9449,N_2452,N_1358);
nand U9450 (N_9450,N_4538,N_1003);
nand U9451 (N_9451,N_2721,N_4223);
and U9452 (N_9452,N_3167,N_3308);
nor U9453 (N_9453,N_12,N_989);
xor U9454 (N_9454,N_4397,N_862);
and U9455 (N_9455,N_400,N_3658);
xnor U9456 (N_9456,N_2730,N_2818);
nor U9457 (N_9457,N_1354,N_1609);
nor U9458 (N_9458,N_471,N_2437);
or U9459 (N_9459,N_4620,N_2020);
nor U9460 (N_9460,N_4005,N_712);
nor U9461 (N_9461,N_4560,N_1140);
nand U9462 (N_9462,N_2387,N_819);
nand U9463 (N_9463,N_1031,N_3474);
nand U9464 (N_9464,N_1406,N_2420);
nand U9465 (N_9465,N_4252,N_1585);
xor U9466 (N_9466,N_1651,N_138);
nand U9467 (N_9467,N_2548,N_4545);
nor U9468 (N_9468,N_557,N_2428);
nor U9469 (N_9469,N_2004,N_2094);
nand U9470 (N_9470,N_3328,N_4710);
and U9471 (N_9471,N_3757,N_1159);
and U9472 (N_9472,N_1878,N_4045);
and U9473 (N_9473,N_374,N_2635);
nor U9474 (N_9474,N_3672,N_737);
and U9475 (N_9475,N_13,N_4896);
and U9476 (N_9476,N_4711,N_2029);
nand U9477 (N_9477,N_791,N_3095);
and U9478 (N_9478,N_4045,N_2801);
or U9479 (N_9479,N_2838,N_2475);
xor U9480 (N_9480,N_289,N_3674);
nor U9481 (N_9481,N_3581,N_2264);
nand U9482 (N_9482,N_836,N_974);
nand U9483 (N_9483,N_3932,N_2791);
nor U9484 (N_9484,N_4648,N_4364);
nand U9485 (N_9485,N_3859,N_4318);
nand U9486 (N_9486,N_1910,N_1290);
or U9487 (N_9487,N_4818,N_1063);
nand U9488 (N_9488,N_260,N_2003);
nand U9489 (N_9489,N_1085,N_4025);
nand U9490 (N_9490,N_2122,N_2989);
nand U9491 (N_9491,N_202,N_4938);
and U9492 (N_9492,N_1848,N_2732);
nor U9493 (N_9493,N_2486,N_2698);
xor U9494 (N_9494,N_1051,N_2938);
nor U9495 (N_9495,N_1639,N_4724);
or U9496 (N_9496,N_559,N_1018);
nor U9497 (N_9497,N_1491,N_88);
or U9498 (N_9498,N_2860,N_1587);
or U9499 (N_9499,N_4091,N_3851);
and U9500 (N_9500,N_369,N_4815);
xnor U9501 (N_9501,N_529,N_1974);
and U9502 (N_9502,N_1633,N_149);
or U9503 (N_9503,N_312,N_748);
xnor U9504 (N_9504,N_99,N_3306);
or U9505 (N_9505,N_3069,N_4853);
nor U9506 (N_9506,N_3511,N_602);
nor U9507 (N_9507,N_1307,N_691);
nor U9508 (N_9508,N_2904,N_110);
nand U9509 (N_9509,N_1083,N_4341);
or U9510 (N_9510,N_1010,N_1106);
nor U9511 (N_9511,N_1376,N_4872);
xnor U9512 (N_9512,N_152,N_600);
nand U9513 (N_9513,N_4746,N_1424);
and U9514 (N_9514,N_2631,N_3567);
nand U9515 (N_9515,N_100,N_4581);
and U9516 (N_9516,N_4705,N_3117);
nand U9517 (N_9517,N_3297,N_4243);
and U9518 (N_9518,N_183,N_1068);
nor U9519 (N_9519,N_1827,N_3734);
or U9520 (N_9520,N_4834,N_3383);
nand U9521 (N_9521,N_2241,N_4412);
or U9522 (N_9522,N_620,N_808);
or U9523 (N_9523,N_301,N_1794);
and U9524 (N_9524,N_2523,N_4803);
xor U9525 (N_9525,N_603,N_1855);
and U9526 (N_9526,N_4113,N_3921);
or U9527 (N_9527,N_2486,N_1380);
nor U9528 (N_9528,N_2070,N_91);
and U9529 (N_9529,N_41,N_3295);
nand U9530 (N_9530,N_4995,N_381);
nand U9531 (N_9531,N_4667,N_2409);
or U9532 (N_9532,N_2106,N_1337);
xor U9533 (N_9533,N_3314,N_2341);
xnor U9534 (N_9534,N_16,N_1614);
and U9535 (N_9535,N_4706,N_3640);
nand U9536 (N_9536,N_1067,N_303);
and U9537 (N_9537,N_22,N_3384);
nor U9538 (N_9538,N_94,N_1749);
and U9539 (N_9539,N_3406,N_1013);
and U9540 (N_9540,N_3622,N_2976);
or U9541 (N_9541,N_3888,N_1806);
nand U9542 (N_9542,N_251,N_1203);
nor U9543 (N_9543,N_2962,N_3041);
nand U9544 (N_9544,N_145,N_3812);
and U9545 (N_9545,N_2802,N_2248);
and U9546 (N_9546,N_4139,N_1741);
or U9547 (N_9547,N_811,N_2576);
or U9548 (N_9548,N_2910,N_843);
and U9549 (N_9549,N_2215,N_3001);
xor U9550 (N_9550,N_3132,N_2027);
or U9551 (N_9551,N_405,N_4644);
nand U9552 (N_9552,N_2805,N_4014);
nor U9553 (N_9553,N_430,N_839);
nand U9554 (N_9554,N_1237,N_4897);
nand U9555 (N_9555,N_1655,N_4274);
nor U9556 (N_9556,N_1584,N_2261);
or U9557 (N_9557,N_1245,N_2606);
nor U9558 (N_9558,N_66,N_4526);
nand U9559 (N_9559,N_4096,N_4967);
xor U9560 (N_9560,N_1889,N_1610);
xor U9561 (N_9561,N_1292,N_4546);
nand U9562 (N_9562,N_2894,N_1595);
or U9563 (N_9563,N_3897,N_4383);
and U9564 (N_9564,N_1336,N_3440);
nor U9565 (N_9565,N_3094,N_4105);
nand U9566 (N_9566,N_1598,N_1825);
and U9567 (N_9567,N_356,N_1417);
nor U9568 (N_9568,N_4524,N_1469);
xor U9569 (N_9569,N_2555,N_1939);
and U9570 (N_9570,N_1238,N_2236);
nand U9571 (N_9571,N_2944,N_1053);
or U9572 (N_9572,N_2891,N_3415);
nand U9573 (N_9573,N_3695,N_4092);
xnor U9574 (N_9574,N_2714,N_1453);
nor U9575 (N_9575,N_3185,N_753);
nor U9576 (N_9576,N_3749,N_2206);
or U9577 (N_9577,N_4093,N_4619);
nor U9578 (N_9578,N_4382,N_1446);
and U9579 (N_9579,N_4113,N_817);
xor U9580 (N_9580,N_2153,N_2838);
xor U9581 (N_9581,N_3728,N_4333);
or U9582 (N_9582,N_2730,N_739);
nor U9583 (N_9583,N_1115,N_4915);
xor U9584 (N_9584,N_2146,N_4638);
and U9585 (N_9585,N_2299,N_1373);
xnor U9586 (N_9586,N_4773,N_1656);
and U9587 (N_9587,N_1885,N_1247);
or U9588 (N_9588,N_3369,N_2354);
and U9589 (N_9589,N_7,N_344);
nor U9590 (N_9590,N_4893,N_4017);
or U9591 (N_9591,N_3837,N_3460);
nand U9592 (N_9592,N_3462,N_438);
or U9593 (N_9593,N_4412,N_4238);
xor U9594 (N_9594,N_4635,N_4556);
nor U9595 (N_9595,N_1827,N_4485);
nor U9596 (N_9596,N_447,N_4029);
nand U9597 (N_9597,N_4634,N_727);
nand U9598 (N_9598,N_3507,N_2419);
and U9599 (N_9599,N_2594,N_1509);
xor U9600 (N_9600,N_1195,N_1764);
nor U9601 (N_9601,N_4315,N_4993);
xnor U9602 (N_9602,N_4405,N_597);
or U9603 (N_9603,N_4913,N_3956);
nor U9604 (N_9604,N_2516,N_1131);
and U9605 (N_9605,N_4930,N_2958);
or U9606 (N_9606,N_274,N_3882);
and U9607 (N_9607,N_3773,N_4188);
or U9608 (N_9608,N_2301,N_3556);
nand U9609 (N_9609,N_4416,N_1889);
nor U9610 (N_9610,N_2682,N_2771);
nand U9611 (N_9611,N_4266,N_2235);
or U9612 (N_9612,N_777,N_1250);
nand U9613 (N_9613,N_4653,N_2309);
and U9614 (N_9614,N_3843,N_742);
xor U9615 (N_9615,N_2275,N_4053);
or U9616 (N_9616,N_2259,N_2539);
nand U9617 (N_9617,N_2215,N_3822);
and U9618 (N_9618,N_2915,N_14);
or U9619 (N_9619,N_2906,N_2663);
nand U9620 (N_9620,N_1172,N_4326);
xnor U9621 (N_9621,N_2048,N_2527);
and U9622 (N_9622,N_534,N_2278);
and U9623 (N_9623,N_3827,N_2482);
xnor U9624 (N_9624,N_679,N_445);
and U9625 (N_9625,N_1374,N_997);
and U9626 (N_9626,N_2868,N_4428);
nor U9627 (N_9627,N_214,N_3480);
xor U9628 (N_9628,N_1832,N_680);
and U9629 (N_9629,N_1881,N_782);
or U9630 (N_9630,N_2106,N_2778);
and U9631 (N_9631,N_3864,N_4753);
xnor U9632 (N_9632,N_2199,N_487);
nand U9633 (N_9633,N_590,N_2683);
nor U9634 (N_9634,N_2003,N_2656);
or U9635 (N_9635,N_2676,N_3135);
nor U9636 (N_9636,N_1169,N_724);
xnor U9637 (N_9637,N_400,N_1017);
or U9638 (N_9638,N_4071,N_1305);
nand U9639 (N_9639,N_4094,N_2063);
and U9640 (N_9640,N_4517,N_3698);
or U9641 (N_9641,N_4464,N_2847);
nand U9642 (N_9642,N_1416,N_2514);
nor U9643 (N_9643,N_96,N_4098);
nor U9644 (N_9644,N_4187,N_992);
and U9645 (N_9645,N_3267,N_3629);
and U9646 (N_9646,N_2976,N_2033);
nand U9647 (N_9647,N_3747,N_3632);
xnor U9648 (N_9648,N_2889,N_4252);
or U9649 (N_9649,N_3987,N_3162);
nand U9650 (N_9650,N_702,N_1320);
nor U9651 (N_9651,N_2364,N_2738);
or U9652 (N_9652,N_849,N_2600);
nand U9653 (N_9653,N_4360,N_310);
and U9654 (N_9654,N_462,N_222);
xor U9655 (N_9655,N_2179,N_614);
and U9656 (N_9656,N_2494,N_1769);
nor U9657 (N_9657,N_977,N_4168);
or U9658 (N_9658,N_229,N_2904);
nor U9659 (N_9659,N_4954,N_1337);
xor U9660 (N_9660,N_854,N_839);
xor U9661 (N_9661,N_2112,N_1110);
or U9662 (N_9662,N_1484,N_2672);
nand U9663 (N_9663,N_2353,N_3921);
or U9664 (N_9664,N_2976,N_2863);
xor U9665 (N_9665,N_3561,N_96);
and U9666 (N_9666,N_3143,N_2464);
nand U9667 (N_9667,N_2498,N_3118);
or U9668 (N_9668,N_2202,N_4320);
nand U9669 (N_9669,N_435,N_4876);
xnor U9670 (N_9670,N_4508,N_4438);
nand U9671 (N_9671,N_4227,N_4690);
or U9672 (N_9672,N_1043,N_4517);
nand U9673 (N_9673,N_4944,N_522);
and U9674 (N_9674,N_3025,N_4569);
or U9675 (N_9675,N_2600,N_2885);
and U9676 (N_9676,N_1560,N_3096);
xnor U9677 (N_9677,N_3620,N_954);
or U9678 (N_9678,N_3418,N_389);
nor U9679 (N_9679,N_1138,N_3833);
xnor U9680 (N_9680,N_2842,N_801);
xor U9681 (N_9681,N_4995,N_1041);
xor U9682 (N_9682,N_4166,N_34);
and U9683 (N_9683,N_1286,N_791);
and U9684 (N_9684,N_4264,N_202);
and U9685 (N_9685,N_2709,N_1437);
and U9686 (N_9686,N_4948,N_2800);
xor U9687 (N_9687,N_3998,N_1112);
and U9688 (N_9688,N_3568,N_1432);
nor U9689 (N_9689,N_3123,N_4994);
and U9690 (N_9690,N_3138,N_1705);
nand U9691 (N_9691,N_1445,N_1398);
or U9692 (N_9692,N_2915,N_3444);
xor U9693 (N_9693,N_4451,N_3123);
or U9694 (N_9694,N_2438,N_340);
nor U9695 (N_9695,N_368,N_4730);
and U9696 (N_9696,N_1132,N_3554);
or U9697 (N_9697,N_4871,N_3770);
and U9698 (N_9698,N_1000,N_758);
nand U9699 (N_9699,N_1171,N_4676);
xor U9700 (N_9700,N_868,N_1718);
nand U9701 (N_9701,N_2696,N_2062);
or U9702 (N_9702,N_4958,N_4212);
xnor U9703 (N_9703,N_1880,N_4878);
and U9704 (N_9704,N_1401,N_2309);
and U9705 (N_9705,N_2000,N_79);
or U9706 (N_9706,N_1068,N_4041);
or U9707 (N_9707,N_2349,N_460);
and U9708 (N_9708,N_2097,N_425);
nand U9709 (N_9709,N_1258,N_1025);
xnor U9710 (N_9710,N_4377,N_1009);
nor U9711 (N_9711,N_773,N_667);
or U9712 (N_9712,N_2649,N_2646);
nand U9713 (N_9713,N_3544,N_4296);
xor U9714 (N_9714,N_2800,N_847);
nand U9715 (N_9715,N_2623,N_4003);
and U9716 (N_9716,N_611,N_3950);
or U9717 (N_9717,N_853,N_4045);
xnor U9718 (N_9718,N_3833,N_2801);
nand U9719 (N_9719,N_2179,N_2033);
nand U9720 (N_9720,N_3550,N_144);
and U9721 (N_9721,N_3150,N_780);
nor U9722 (N_9722,N_1657,N_4317);
or U9723 (N_9723,N_4508,N_3155);
nand U9724 (N_9724,N_48,N_2715);
or U9725 (N_9725,N_2814,N_3806);
xor U9726 (N_9726,N_344,N_2773);
or U9727 (N_9727,N_1598,N_1260);
and U9728 (N_9728,N_1609,N_450);
nor U9729 (N_9729,N_2119,N_1729);
xnor U9730 (N_9730,N_3062,N_3974);
nor U9731 (N_9731,N_1552,N_3456);
nor U9732 (N_9732,N_451,N_3080);
and U9733 (N_9733,N_1873,N_347);
or U9734 (N_9734,N_3954,N_2480);
and U9735 (N_9735,N_2400,N_1492);
xnor U9736 (N_9736,N_2462,N_4774);
nand U9737 (N_9737,N_991,N_534);
and U9738 (N_9738,N_4560,N_515);
nor U9739 (N_9739,N_3602,N_3822);
nor U9740 (N_9740,N_659,N_2630);
nor U9741 (N_9741,N_1370,N_1091);
xnor U9742 (N_9742,N_3869,N_1856);
or U9743 (N_9743,N_4859,N_308);
xor U9744 (N_9744,N_3736,N_4633);
xor U9745 (N_9745,N_741,N_4891);
xnor U9746 (N_9746,N_1297,N_2375);
xnor U9747 (N_9747,N_3625,N_463);
xnor U9748 (N_9748,N_4021,N_2479);
nor U9749 (N_9749,N_4965,N_1258);
xnor U9750 (N_9750,N_2653,N_936);
xnor U9751 (N_9751,N_3952,N_284);
xor U9752 (N_9752,N_3858,N_970);
nand U9753 (N_9753,N_3867,N_2952);
or U9754 (N_9754,N_4797,N_3407);
nor U9755 (N_9755,N_4405,N_1076);
nand U9756 (N_9756,N_4484,N_2186);
nor U9757 (N_9757,N_1136,N_3411);
nand U9758 (N_9758,N_4264,N_4478);
nor U9759 (N_9759,N_2679,N_4962);
xor U9760 (N_9760,N_2750,N_696);
nor U9761 (N_9761,N_1934,N_2189);
nor U9762 (N_9762,N_1689,N_2816);
and U9763 (N_9763,N_172,N_3109);
nand U9764 (N_9764,N_1856,N_4543);
or U9765 (N_9765,N_2361,N_2105);
nand U9766 (N_9766,N_4755,N_3427);
nand U9767 (N_9767,N_1198,N_2285);
nand U9768 (N_9768,N_484,N_1927);
or U9769 (N_9769,N_1142,N_1607);
xor U9770 (N_9770,N_4115,N_229);
and U9771 (N_9771,N_4988,N_412);
or U9772 (N_9772,N_2329,N_3025);
and U9773 (N_9773,N_3119,N_4919);
and U9774 (N_9774,N_897,N_2709);
nand U9775 (N_9775,N_3947,N_1596);
nand U9776 (N_9776,N_3594,N_4351);
and U9777 (N_9777,N_84,N_4117);
or U9778 (N_9778,N_159,N_3621);
or U9779 (N_9779,N_971,N_4660);
or U9780 (N_9780,N_4862,N_111);
or U9781 (N_9781,N_4542,N_4235);
nand U9782 (N_9782,N_4954,N_1015);
or U9783 (N_9783,N_4428,N_1472);
nor U9784 (N_9784,N_1389,N_4405);
or U9785 (N_9785,N_2162,N_3723);
nand U9786 (N_9786,N_658,N_613);
xnor U9787 (N_9787,N_2965,N_4185);
and U9788 (N_9788,N_641,N_2199);
or U9789 (N_9789,N_993,N_1303);
xor U9790 (N_9790,N_92,N_1748);
or U9791 (N_9791,N_1821,N_4666);
nor U9792 (N_9792,N_2104,N_4338);
nor U9793 (N_9793,N_1107,N_1944);
xnor U9794 (N_9794,N_1360,N_3510);
and U9795 (N_9795,N_4946,N_3506);
and U9796 (N_9796,N_1706,N_3817);
nand U9797 (N_9797,N_1799,N_2410);
xor U9798 (N_9798,N_2020,N_1856);
or U9799 (N_9799,N_4093,N_3679);
and U9800 (N_9800,N_2145,N_3490);
or U9801 (N_9801,N_2024,N_417);
xor U9802 (N_9802,N_2811,N_1211);
xor U9803 (N_9803,N_3149,N_3790);
xor U9804 (N_9804,N_2005,N_6);
nand U9805 (N_9805,N_3143,N_4685);
and U9806 (N_9806,N_3972,N_3737);
or U9807 (N_9807,N_3784,N_1590);
xor U9808 (N_9808,N_2801,N_3449);
xor U9809 (N_9809,N_2935,N_64);
nand U9810 (N_9810,N_1536,N_2025);
xnor U9811 (N_9811,N_556,N_3596);
xor U9812 (N_9812,N_3471,N_749);
nor U9813 (N_9813,N_3419,N_1694);
or U9814 (N_9814,N_264,N_2530);
nor U9815 (N_9815,N_2185,N_2513);
and U9816 (N_9816,N_4470,N_3238);
xnor U9817 (N_9817,N_565,N_4343);
xnor U9818 (N_9818,N_4444,N_3278);
and U9819 (N_9819,N_1381,N_737);
or U9820 (N_9820,N_3694,N_3204);
and U9821 (N_9821,N_4956,N_1425);
or U9822 (N_9822,N_1243,N_3747);
and U9823 (N_9823,N_2378,N_2172);
nor U9824 (N_9824,N_967,N_1557);
xor U9825 (N_9825,N_3208,N_2370);
nand U9826 (N_9826,N_4062,N_1164);
nor U9827 (N_9827,N_1462,N_1452);
xor U9828 (N_9828,N_3217,N_4180);
or U9829 (N_9829,N_4768,N_4973);
or U9830 (N_9830,N_967,N_3375);
and U9831 (N_9831,N_4867,N_2570);
and U9832 (N_9832,N_1630,N_743);
xnor U9833 (N_9833,N_954,N_3664);
and U9834 (N_9834,N_2538,N_3629);
nor U9835 (N_9835,N_3209,N_651);
nor U9836 (N_9836,N_619,N_1543);
and U9837 (N_9837,N_3986,N_2881);
or U9838 (N_9838,N_1637,N_391);
and U9839 (N_9839,N_1267,N_4549);
and U9840 (N_9840,N_3800,N_2379);
and U9841 (N_9841,N_1252,N_860);
and U9842 (N_9842,N_1593,N_1375);
and U9843 (N_9843,N_3300,N_1478);
or U9844 (N_9844,N_3144,N_823);
and U9845 (N_9845,N_4239,N_4187);
or U9846 (N_9846,N_4227,N_3201);
and U9847 (N_9847,N_3800,N_4917);
xor U9848 (N_9848,N_1105,N_269);
nand U9849 (N_9849,N_2913,N_3554);
nand U9850 (N_9850,N_1288,N_1025);
and U9851 (N_9851,N_3379,N_2325);
nand U9852 (N_9852,N_4961,N_1489);
nor U9853 (N_9853,N_2946,N_354);
nor U9854 (N_9854,N_4138,N_4482);
nand U9855 (N_9855,N_4439,N_43);
and U9856 (N_9856,N_3006,N_3029);
nor U9857 (N_9857,N_1697,N_1258);
or U9858 (N_9858,N_1744,N_1675);
and U9859 (N_9859,N_3295,N_1503);
nand U9860 (N_9860,N_4081,N_1961);
or U9861 (N_9861,N_958,N_903);
or U9862 (N_9862,N_2049,N_3704);
nor U9863 (N_9863,N_4066,N_3596);
nand U9864 (N_9864,N_3675,N_1164);
or U9865 (N_9865,N_224,N_2562);
and U9866 (N_9866,N_4225,N_4855);
nand U9867 (N_9867,N_199,N_1696);
nand U9868 (N_9868,N_1349,N_484);
xor U9869 (N_9869,N_2947,N_3273);
or U9870 (N_9870,N_572,N_2634);
and U9871 (N_9871,N_4397,N_699);
nor U9872 (N_9872,N_97,N_152);
or U9873 (N_9873,N_166,N_445);
nor U9874 (N_9874,N_899,N_4047);
xor U9875 (N_9875,N_917,N_1068);
or U9876 (N_9876,N_3191,N_4065);
nor U9877 (N_9877,N_1505,N_4355);
and U9878 (N_9878,N_2834,N_227);
or U9879 (N_9879,N_2649,N_2057);
nor U9880 (N_9880,N_3164,N_4987);
xor U9881 (N_9881,N_4007,N_1537);
xnor U9882 (N_9882,N_527,N_2904);
nor U9883 (N_9883,N_3758,N_2387);
xor U9884 (N_9884,N_1707,N_4240);
nand U9885 (N_9885,N_60,N_4212);
nand U9886 (N_9886,N_2488,N_2698);
or U9887 (N_9887,N_531,N_4258);
nor U9888 (N_9888,N_2183,N_214);
and U9889 (N_9889,N_1115,N_3244);
and U9890 (N_9890,N_3959,N_3884);
nor U9891 (N_9891,N_3978,N_1992);
xnor U9892 (N_9892,N_2432,N_3983);
or U9893 (N_9893,N_3355,N_3995);
xnor U9894 (N_9894,N_1561,N_2965);
and U9895 (N_9895,N_3046,N_4797);
nand U9896 (N_9896,N_2034,N_2237);
or U9897 (N_9897,N_3580,N_4931);
nor U9898 (N_9898,N_4008,N_1479);
nor U9899 (N_9899,N_2701,N_2527);
nor U9900 (N_9900,N_2752,N_4583);
nand U9901 (N_9901,N_3870,N_290);
nand U9902 (N_9902,N_801,N_2097);
nand U9903 (N_9903,N_4434,N_3434);
and U9904 (N_9904,N_3117,N_2554);
or U9905 (N_9905,N_3905,N_287);
and U9906 (N_9906,N_2451,N_3658);
xor U9907 (N_9907,N_347,N_2436);
or U9908 (N_9908,N_1228,N_1709);
or U9909 (N_9909,N_4389,N_430);
or U9910 (N_9910,N_842,N_4602);
or U9911 (N_9911,N_4723,N_1643);
xnor U9912 (N_9912,N_3042,N_3006);
xor U9913 (N_9913,N_332,N_2092);
or U9914 (N_9914,N_2531,N_1519);
and U9915 (N_9915,N_1247,N_2600);
or U9916 (N_9916,N_4519,N_1852);
nand U9917 (N_9917,N_3555,N_2001);
nand U9918 (N_9918,N_1232,N_899);
and U9919 (N_9919,N_1005,N_929);
nand U9920 (N_9920,N_4718,N_4472);
and U9921 (N_9921,N_1290,N_81);
or U9922 (N_9922,N_685,N_1469);
nand U9923 (N_9923,N_1206,N_621);
and U9924 (N_9924,N_2311,N_101);
nor U9925 (N_9925,N_4401,N_3061);
or U9926 (N_9926,N_188,N_1501);
and U9927 (N_9927,N_3248,N_3467);
nand U9928 (N_9928,N_4817,N_4904);
xor U9929 (N_9929,N_4645,N_142);
xor U9930 (N_9930,N_4792,N_2689);
nor U9931 (N_9931,N_2949,N_498);
xor U9932 (N_9932,N_3135,N_927);
or U9933 (N_9933,N_2462,N_4048);
nor U9934 (N_9934,N_4004,N_2606);
nor U9935 (N_9935,N_2800,N_2336);
xor U9936 (N_9936,N_1947,N_4435);
and U9937 (N_9937,N_2451,N_742);
and U9938 (N_9938,N_424,N_4997);
xnor U9939 (N_9939,N_4891,N_3429);
xnor U9940 (N_9940,N_3127,N_3824);
xnor U9941 (N_9941,N_4925,N_2184);
nor U9942 (N_9942,N_3699,N_2042);
or U9943 (N_9943,N_4717,N_1630);
nor U9944 (N_9944,N_3181,N_1755);
nor U9945 (N_9945,N_564,N_2740);
nand U9946 (N_9946,N_4068,N_2981);
xor U9947 (N_9947,N_1615,N_4094);
nand U9948 (N_9948,N_3251,N_2097);
and U9949 (N_9949,N_3874,N_2816);
xnor U9950 (N_9950,N_3205,N_3017);
xor U9951 (N_9951,N_2449,N_3348);
nor U9952 (N_9952,N_2965,N_1053);
and U9953 (N_9953,N_4338,N_2115);
nand U9954 (N_9954,N_2056,N_620);
nand U9955 (N_9955,N_1051,N_4261);
nor U9956 (N_9956,N_4786,N_829);
and U9957 (N_9957,N_156,N_2967);
xor U9958 (N_9958,N_3053,N_877);
or U9959 (N_9959,N_1722,N_4751);
nor U9960 (N_9960,N_1338,N_1400);
or U9961 (N_9961,N_3453,N_4347);
nand U9962 (N_9962,N_707,N_3084);
xor U9963 (N_9963,N_4207,N_1335);
and U9964 (N_9964,N_2578,N_3914);
nand U9965 (N_9965,N_1519,N_4922);
nor U9966 (N_9966,N_4234,N_4040);
and U9967 (N_9967,N_3199,N_3645);
nand U9968 (N_9968,N_484,N_4696);
nor U9969 (N_9969,N_3040,N_554);
or U9970 (N_9970,N_4040,N_3923);
and U9971 (N_9971,N_676,N_4825);
and U9972 (N_9972,N_1615,N_3326);
xor U9973 (N_9973,N_2844,N_3733);
xnor U9974 (N_9974,N_1296,N_2199);
and U9975 (N_9975,N_2496,N_4856);
nand U9976 (N_9976,N_822,N_1767);
nor U9977 (N_9977,N_3084,N_1310);
nand U9978 (N_9978,N_4329,N_2194);
or U9979 (N_9979,N_672,N_539);
nand U9980 (N_9980,N_952,N_487);
or U9981 (N_9981,N_3072,N_1968);
xor U9982 (N_9982,N_4202,N_3138);
and U9983 (N_9983,N_4340,N_673);
and U9984 (N_9984,N_1431,N_540);
or U9985 (N_9985,N_1160,N_3750);
xor U9986 (N_9986,N_1061,N_2013);
or U9987 (N_9987,N_1244,N_3324);
nor U9988 (N_9988,N_4254,N_1632);
xnor U9989 (N_9989,N_3922,N_2003);
nand U9990 (N_9990,N_863,N_1048);
or U9991 (N_9991,N_1874,N_335);
nor U9992 (N_9992,N_1313,N_1894);
and U9993 (N_9993,N_4774,N_2967);
or U9994 (N_9994,N_3348,N_2531);
or U9995 (N_9995,N_3913,N_1746);
and U9996 (N_9996,N_4412,N_3906);
or U9997 (N_9997,N_4646,N_4038);
and U9998 (N_9998,N_4046,N_431);
nand U9999 (N_9999,N_191,N_3686);
and U10000 (N_10000,N_5439,N_6910);
nor U10001 (N_10001,N_5065,N_8690);
or U10002 (N_10002,N_5720,N_6163);
xor U10003 (N_10003,N_6267,N_7046);
and U10004 (N_10004,N_6593,N_6509);
or U10005 (N_10005,N_8846,N_5420);
or U10006 (N_10006,N_5651,N_8128);
nor U10007 (N_10007,N_6051,N_6662);
xor U10008 (N_10008,N_9285,N_8401);
xnor U10009 (N_10009,N_5454,N_5832);
nand U10010 (N_10010,N_6191,N_8938);
nand U10011 (N_10011,N_5629,N_8209);
and U10012 (N_10012,N_6245,N_7304);
xnor U10013 (N_10013,N_6804,N_7763);
xnor U10014 (N_10014,N_5884,N_8254);
nor U10015 (N_10015,N_9408,N_7322);
or U10016 (N_10016,N_8032,N_5365);
xor U10017 (N_10017,N_9592,N_8957);
or U10018 (N_10018,N_6115,N_6428);
nor U10019 (N_10019,N_5422,N_6471);
nor U10020 (N_10020,N_7145,N_6969);
and U10021 (N_10021,N_6608,N_6644);
or U10022 (N_10022,N_8852,N_9126);
or U10023 (N_10023,N_6948,N_7937);
or U10024 (N_10024,N_8115,N_8969);
nor U10025 (N_10025,N_8974,N_5627);
or U10026 (N_10026,N_7952,N_5515);
nor U10027 (N_10027,N_6551,N_9044);
and U10028 (N_10028,N_5687,N_5797);
and U10029 (N_10029,N_8861,N_5142);
and U10030 (N_10030,N_8179,N_8421);
and U10031 (N_10031,N_5663,N_6974);
or U10032 (N_10032,N_9920,N_9003);
xnor U10033 (N_10033,N_6415,N_9441);
nor U10034 (N_10034,N_9498,N_8737);
or U10035 (N_10035,N_9307,N_7930);
or U10036 (N_10036,N_8781,N_7258);
nor U10037 (N_10037,N_6376,N_5685);
nand U10038 (N_10038,N_9131,N_5602);
nand U10039 (N_10039,N_9090,N_6702);
xor U10040 (N_10040,N_9310,N_6556);
and U10041 (N_10041,N_9554,N_9296);
nand U10042 (N_10042,N_6962,N_8892);
nor U10043 (N_10043,N_5985,N_7005);
or U10044 (N_10044,N_8831,N_7629);
nor U10045 (N_10045,N_6324,N_5398);
nor U10046 (N_10046,N_6041,N_7080);
and U10047 (N_10047,N_5689,N_6583);
nand U10048 (N_10048,N_8211,N_9020);
or U10049 (N_10049,N_7924,N_7075);
and U10050 (N_10050,N_7237,N_8809);
nand U10051 (N_10051,N_5086,N_9396);
or U10052 (N_10052,N_6027,N_8444);
or U10053 (N_10053,N_6176,N_6648);
nor U10054 (N_10054,N_7708,N_9968);
nor U10055 (N_10055,N_8180,N_8662);
and U10056 (N_10056,N_8870,N_5928);
and U10057 (N_10057,N_6894,N_9382);
nand U10058 (N_10058,N_9555,N_6122);
and U10059 (N_10059,N_6280,N_7283);
nor U10060 (N_10060,N_6299,N_9801);
nor U10061 (N_10061,N_8124,N_5566);
nor U10062 (N_10062,N_5227,N_6769);
and U10063 (N_10063,N_6255,N_8789);
or U10064 (N_10064,N_7895,N_6935);
nor U10065 (N_10065,N_8205,N_8986);
or U10066 (N_10066,N_9717,N_5939);
xor U10067 (N_10067,N_9085,N_6628);
nand U10068 (N_10068,N_9014,N_5618);
or U10069 (N_10069,N_8497,N_9141);
nand U10070 (N_10070,N_9199,N_9488);
xor U10071 (N_10071,N_8890,N_9982);
or U10072 (N_10072,N_5571,N_8730);
nor U10073 (N_10073,N_5081,N_5074);
or U10074 (N_10074,N_8388,N_7058);
xor U10075 (N_10075,N_9144,N_7712);
xor U10076 (N_10076,N_7330,N_7940);
nand U10077 (N_10077,N_5414,N_6683);
nor U10078 (N_10078,N_7262,N_8677);
or U10079 (N_10079,N_5171,N_8481);
or U10080 (N_10080,N_8150,N_7980);
xnor U10081 (N_10081,N_8098,N_8676);
xor U10082 (N_10082,N_9526,N_9262);
nand U10083 (N_10083,N_8556,N_6486);
and U10084 (N_10084,N_8782,N_6447);
nor U10085 (N_10085,N_9768,N_8772);
nor U10086 (N_10086,N_8377,N_5197);
or U10087 (N_10087,N_8891,N_9933);
and U10088 (N_10088,N_9538,N_7527);
and U10089 (N_10089,N_6800,N_7321);
xor U10090 (N_10090,N_6254,N_7383);
and U10091 (N_10091,N_5528,N_6754);
nand U10092 (N_10092,N_6738,N_7843);
xnor U10093 (N_10093,N_9814,N_7561);
or U10094 (N_10094,N_7280,N_8470);
and U10095 (N_10095,N_8322,N_9347);
xor U10096 (N_10096,N_5290,N_6316);
nor U10097 (N_10097,N_8043,N_5781);
nor U10098 (N_10098,N_5619,N_8167);
nand U10099 (N_10099,N_9461,N_7423);
nand U10100 (N_10100,N_7549,N_9688);
xor U10101 (N_10101,N_5851,N_9989);
and U10102 (N_10102,N_9708,N_9251);
or U10103 (N_10103,N_8999,N_5683);
and U10104 (N_10104,N_6923,N_7025);
and U10105 (N_10105,N_5043,N_5057);
xor U10106 (N_10106,N_7996,N_7380);
nor U10107 (N_10107,N_8888,N_5843);
or U10108 (N_10108,N_5117,N_7488);
and U10109 (N_10109,N_6806,N_5765);
and U10110 (N_10110,N_9980,N_6523);
or U10111 (N_10111,N_6525,N_7516);
xnor U10112 (N_10112,N_8199,N_5662);
xnor U10113 (N_10113,N_5527,N_5650);
xnor U10114 (N_10114,N_8825,N_7230);
nor U10115 (N_10115,N_9107,N_9115);
and U10116 (N_10116,N_8183,N_8193);
nor U10117 (N_10117,N_7818,N_9692);
xnor U10118 (N_10118,N_9274,N_7781);
xor U10119 (N_10119,N_9471,N_8044);
nand U10120 (N_10120,N_8505,N_5927);
xnor U10121 (N_10121,N_6646,N_8758);
nor U10122 (N_10122,N_6013,N_6076);
xnor U10123 (N_10123,N_8403,N_7071);
nor U10124 (N_10124,N_5854,N_6421);
or U10125 (N_10125,N_6217,N_9777);
nand U10126 (N_10126,N_8640,N_7081);
nor U10127 (N_10127,N_8534,N_5358);
or U10128 (N_10128,N_9237,N_9084);
nand U10129 (N_10129,N_9186,N_7630);
or U10130 (N_10130,N_9765,N_8268);
xnor U10131 (N_10131,N_8887,N_7426);
nand U10132 (N_10132,N_6364,N_8682);
and U10133 (N_10133,N_5071,N_7251);
and U10134 (N_10134,N_6949,N_8227);
nor U10135 (N_10135,N_6695,N_7395);
xnor U10136 (N_10136,N_9574,N_6391);
or U10137 (N_10137,N_5277,N_8422);
or U10138 (N_10138,N_8568,N_5763);
and U10139 (N_10139,N_7185,N_6272);
nand U10140 (N_10140,N_7337,N_6141);
or U10141 (N_10141,N_8394,N_7389);
nor U10142 (N_10142,N_7663,N_9962);
and U10143 (N_10143,N_6188,N_9176);
nand U10144 (N_10144,N_9532,N_5611);
nand U10145 (N_10145,N_6452,N_7319);
or U10146 (N_10146,N_5542,N_8415);
nand U10147 (N_10147,N_8151,N_8427);
nor U10148 (N_10148,N_8702,N_6566);
or U10149 (N_10149,N_5078,N_9293);
and U10150 (N_10150,N_5333,N_5586);
nor U10151 (N_10151,N_8363,N_7816);
nor U10152 (N_10152,N_7370,N_8159);
nor U10153 (N_10153,N_6340,N_8023);
nor U10154 (N_10154,N_7770,N_8406);
or U10155 (N_10155,N_8712,N_9501);
nor U10156 (N_10156,N_6855,N_6393);
or U10157 (N_10157,N_8583,N_8095);
xor U10158 (N_10158,N_6463,N_6507);
and U10159 (N_10159,N_6327,N_5091);
and U10160 (N_10160,N_8136,N_7248);
and U10161 (N_10161,N_5319,N_7520);
nand U10162 (N_10162,N_6331,N_7933);
and U10163 (N_10163,N_7963,N_7265);
xor U10164 (N_10164,N_5001,N_8450);
xnor U10165 (N_10165,N_6614,N_8101);
and U10166 (N_10166,N_8373,N_5433);
nor U10167 (N_10167,N_8121,N_5355);
nand U10168 (N_10168,N_5579,N_8826);
nand U10169 (N_10169,N_9507,N_7635);
xor U10170 (N_10170,N_6479,N_5730);
nand U10171 (N_10171,N_8350,N_8441);
and U10172 (N_10172,N_9531,N_9702);
and U10173 (N_10173,N_7580,N_8691);
nand U10174 (N_10174,N_5581,N_7351);
nor U10175 (N_10175,N_5232,N_8141);
xor U10176 (N_10176,N_9178,N_5608);
and U10177 (N_10177,N_7827,N_8483);
or U10178 (N_10178,N_5200,N_6968);
xor U10179 (N_10179,N_8577,N_7259);
or U10180 (N_10180,N_7226,N_7915);
nand U10181 (N_10181,N_9650,N_8219);
and U10182 (N_10182,N_7539,N_7212);
xor U10183 (N_10183,N_7674,N_8968);
or U10184 (N_10184,N_6901,N_9972);
and U10185 (N_10185,N_7774,N_5309);
xnor U10186 (N_10186,N_5080,N_5140);
nor U10187 (N_10187,N_8975,N_6124);
nand U10188 (N_10188,N_5953,N_9052);
or U10189 (N_10189,N_9660,N_7345);
or U10190 (N_10190,N_9550,N_6559);
and U10191 (N_10191,N_7027,N_5759);
or U10192 (N_10192,N_5762,N_6953);
and U10193 (N_10193,N_8244,N_6455);
and U10194 (N_10194,N_9529,N_6836);
nand U10195 (N_10195,N_7907,N_8645);
or U10196 (N_10196,N_7585,N_7067);
nand U10197 (N_10197,N_9418,N_6419);
or U10198 (N_10198,N_8019,N_6030);
or U10199 (N_10199,N_6519,N_6462);
and U10200 (N_10200,N_8879,N_9102);
or U10201 (N_10201,N_7317,N_9258);
nor U10202 (N_10202,N_8500,N_6793);
and U10203 (N_10203,N_8941,N_6997);
nand U10204 (N_10204,N_7333,N_5338);
or U10205 (N_10205,N_6920,N_9716);
and U10206 (N_10206,N_9887,N_5130);
nand U10207 (N_10207,N_9250,N_8531);
nor U10208 (N_10208,N_6043,N_9598);
xor U10209 (N_10209,N_7161,N_8566);
or U10210 (N_10210,N_7773,N_8960);
nor U10211 (N_10211,N_9425,N_8228);
or U10212 (N_10212,N_8082,N_8426);
or U10213 (N_10213,N_7695,N_9913);
nor U10214 (N_10214,N_5003,N_7335);
and U10215 (N_10215,N_8232,N_6190);
nand U10216 (N_10216,N_8686,N_9436);
or U10217 (N_10217,N_5752,N_7328);
nand U10218 (N_10218,N_9832,N_6125);
xor U10219 (N_10219,N_7641,N_6323);
or U10220 (N_10220,N_8512,N_5942);
xor U10221 (N_10221,N_8806,N_9205);
or U10222 (N_10222,N_5559,N_7332);
xor U10223 (N_10223,N_6232,N_6528);
nor U10224 (N_10224,N_7518,N_6199);
xnor U10225 (N_10225,N_8765,N_5554);
or U10226 (N_10226,N_6240,N_5501);
and U10227 (N_10227,N_7495,N_8718);
nor U10228 (N_10228,N_7702,N_6771);
xnor U10229 (N_10229,N_9698,N_6829);
xnor U10230 (N_10230,N_5099,N_6412);
and U10231 (N_10231,N_9034,N_9482);
and U10232 (N_10232,N_8587,N_5899);
xor U10233 (N_10233,N_7989,N_5361);
and U10234 (N_10234,N_8489,N_6165);
nand U10235 (N_10235,N_6145,N_6161);
nor U10236 (N_10236,N_7897,N_5273);
and U10237 (N_10237,N_5042,N_5263);
or U10238 (N_10238,N_6065,N_7010);
and U10239 (N_10239,N_5346,N_5222);
or U10240 (N_10240,N_9624,N_9076);
nor U10241 (N_10241,N_9192,N_8631);
and U10242 (N_10242,N_6639,N_7078);
xor U10243 (N_10243,N_7448,N_7074);
nand U10244 (N_10244,N_7633,N_6616);
or U10245 (N_10245,N_5745,N_6397);
nand U10246 (N_10246,N_8907,N_9257);
or U10247 (N_10247,N_9451,N_7172);
xnor U10248 (N_10248,N_9625,N_8818);
and U10249 (N_10249,N_8955,N_5183);
nor U10250 (N_10250,N_7888,N_8911);
and U10251 (N_10251,N_5894,N_5029);
or U10252 (N_10252,N_6694,N_8003);
nor U10253 (N_10253,N_9757,N_7961);
nand U10254 (N_10254,N_6404,N_5739);
xnor U10255 (N_10255,N_9934,N_9087);
xnor U10256 (N_10256,N_5425,N_8001);
nand U10257 (N_10257,N_7724,N_8886);
and U10258 (N_10258,N_5727,N_7443);
nand U10259 (N_10259,N_6674,N_7603);
xnor U10260 (N_10260,N_7812,N_7195);
nand U10261 (N_10261,N_8191,N_5865);
nand U10262 (N_10262,N_8139,N_7146);
nand U10263 (N_10263,N_9955,N_7419);
xnor U10264 (N_10264,N_6164,N_6396);
nand U10265 (N_10265,N_7032,N_7284);
and U10266 (N_10266,N_7087,N_7538);
nand U10267 (N_10267,N_7048,N_9630);
and U10268 (N_10268,N_8605,N_9750);
or U10269 (N_10269,N_9118,N_7289);
and U10270 (N_10270,N_9135,N_6685);
nand U10271 (N_10271,N_9764,N_7750);
nor U10272 (N_10272,N_8632,N_7797);
and U10273 (N_10273,N_5858,N_5316);
or U10274 (N_10274,N_6120,N_9782);
nor U10275 (N_10275,N_7662,N_7084);
nand U10276 (N_10276,N_6579,N_8935);
and U10277 (N_10277,N_8466,N_9100);
or U10278 (N_10278,N_5728,N_7036);
nor U10279 (N_10279,N_7642,N_6736);
or U10280 (N_10280,N_5275,N_9416);
or U10281 (N_10281,N_6353,N_7233);
or U10282 (N_10282,N_8693,N_8995);
nor U10283 (N_10283,N_8327,N_9690);
xnor U10284 (N_10284,N_6242,N_9859);
xor U10285 (N_10285,N_7955,N_7399);
xor U10286 (N_10286,N_6945,N_9539);
xor U10287 (N_10287,N_6727,N_9305);
and U10288 (N_10288,N_7679,N_9122);
or U10289 (N_10289,N_9886,N_5421);
and U10290 (N_10290,N_7820,N_7831);
nand U10291 (N_10291,N_7397,N_9220);
nand U10292 (N_10292,N_6664,N_8592);
nand U10293 (N_10293,N_9618,N_7503);
xor U10294 (N_10294,N_6576,N_8787);
nor U10295 (N_10295,N_7623,N_8252);
xor U10296 (N_10296,N_5061,N_5516);
nand U10297 (N_10297,N_9754,N_8759);
or U10298 (N_10298,N_7892,N_7444);
nand U10299 (N_10299,N_8778,N_7649);
nand U10300 (N_10300,N_7061,N_6541);
nor U10301 (N_10301,N_7135,N_9283);
xnor U10302 (N_10302,N_5392,N_9393);
xnor U10303 (N_10303,N_7184,N_8937);
nor U10304 (N_10304,N_5032,N_5005);
nor U10305 (N_10305,N_9064,N_5401);
nor U10306 (N_10306,N_9331,N_7745);
nand U10307 (N_10307,N_9313,N_9224);
nor U10308 (N_10308,N_6655,N_6786);
xnor U10309 (N_10309,N_5610,N_5758);
nand U10310 (N_10310,N_5167,N_6869);
nor U10311 (N_10311,N_7865,N_9039);
and U10312 (N_10312,N_9005,N_7205);
nor U10313 (N_10313,N_5966,N_6842);
nor U10314 (N_10314,N_9234,N_7835);
xor U10315 (N_10315,N_6742,N_7311);
and U10316 (N_10316,N_8522,N_7502);
xnor U10317 (N_10317,N_5850,N_9926);
nor U10318 (N_10318,N_5933,N_5960);
nand U10319 (N_10319,N_5264,N_8075);
nor U10320 (N_10320,N_6632,N_8142);
or U10321 (N_10321,N_5257,N_5203);
nor U10322 (N_10322,N_9734,N_6365);
or U10323 (N_10323,N_5537,N_8336);
xor U10324 (N_10324,N_5213,N_5779);
nor U10325 (N_10325,N_8253,N_9993);
xor U10326 (N_10326,N_9036,N_7846);
or U10327 (N_10327,N_7267,N_6056);
nand U10328 (N_10328,N_7929,N_6435);
or U10329 (N_10329,N_8635,N_7524);
or U10330 (N_10330,N_7007,N_9735);
and U10331 (N_10331,N_8680,N_5457);
nand U10332 (N_10332,N_8832,N_8041);
or U10333 (N_10333,N_8595,N_9540);
nand U10334 (N_10334,N_6863,N_7686);
and U10335 (N_10335,N_8959,N_6864);
or U10336 (N_10336,N_7992,N_6673);
nand U10337 (N_10337,N_7990,N_9156);
nand U10338 (N_10338,N_9429,N_5702);
or U10339 (N_10339,N_7646,N_5216);
or U10340 (N_10340,N_8212,N_5934);
xnor U10341 (N_10341,N_8794,N_7017);
and U10342 (N_10342,N_8777,N_5048);
nand U10343 (N_10343,N_5922,N_6357);
and U10344 (N_10344,N_8103,N_5652);
and U10345 (N_10345,N_6976,N_9965);
and U10346 (N_10346,N_8520,N_9541);
or U10347 (N_10347,N_8695,N_6814);
and U10348 (N_10348,N_7290,N_5382);
or U10349 (N_10349,N_8611,N_8696);
nor U10350 (N_10350,N_8462,N_5754);
and U10351 (N_10351,N_7204,N_5009);
or U10352 (N_10352,N_6631,N_8857);
nor U10353 (N_10353,N_7090,N_7936);
xnor U10354 (N_10354,N_8560,N_7971);
nand U10355 (N_10355,N_9763,N_6466);
nor U10356 (N_10356,N_8018,N_6368);
and U10357 (N_10357,N_8613,N_9902);
and U10358 (N_10358,N_6290,N_8352);
xor U10359 (N_10359,N_7805,N_5707);
and U10360 (N_10360,N_8515,N_7782);
nor U10361 (N_10361,N_7566,N_6385);
nor U10362 (N_10362,N_6606,N_7749);
xnor U10363 (N_10363,N_7210,N_6483);
nor U10364 (N_10364,N_8882,N_6715);
nor U10365 (N_10365,N_8576,N_6690);
nor U10366 (N_10366,N_6813,N_8815);
or U10367 (N_10367,N_6066,N_9678);
or U10368 (N_10368,N_6339,N_6809);
and U10369 (N_10369,N_7377,N_7747);
nand U10370 (N_10370,N_9970,N_7093);
or U10371 (N_10371,N_6747,N_9861);
nand U10372 (N_10372,N_9204,N_7542);
xor U10373 (N_10373,N_8620,N_8055);
and U10374 (N_10374,N_9974,N_5533);
or U10375 (N_10375,N_8034,N_7769);
nor U10376 (N_10376,N_5569,N_6060);
nor U10377 (N_10377,N_6048,N_7949);
or U10378 (N_10378,N_5380,N_8182);
and U10379 (N_10379,N_5822,N_8865);
nand U10380 (N_10380,N_6828,N_9465);
nand U10381 (N_10381,N_8126,N_7301);
and U10382 (N_10382,N_6511,N_6315);
nor U10383 (N_10383,N_9255,N_5390);
nand U10384 (N_10384,N_9202,N_8723);
or U10385 (N_10385,N_9981,N_7789);
xnor U10386 (N_10386,N_9086,N_8598);
nand U10387 (N_10387,N_8623,N_9196);
or U10388 (N_10388,N_6237,N_8221);
nand U10389 (N_10389,N_8654,N_9149);
nor U10390 (N_10390,N_5228,N_9895);
and U10391 (N_10391,N_6886,N_8156);
or U10392 (N_10392,N_8346,N_6832);
xnor U10393 (N_10393,N_7224,N_6524);
nor U10394 (N_10394,N_5393,N_9388);
or U10395 (N_10395,N_8912,N_9029);
or U10396 (N_10396,N_8056,N_9843);
nor U10397 (N_10397,N_5241,N_5475);
or U10398 (N_10398,N_8049,N_9159);
or U10399 (N_10399,N_5294,N_8436);
nand U10400 (N_10400,N_9997,N_5090);
and U10401 (N_10401,N_9365,N_8451);
xnor U10402 (N_10402,N_8321,N_8864);
or U10403 (N_10403,N_8769,N_7256);
nor U10404 (N_10404,N_9281,N_8954);
and U10405 (N_10405,N_6967,N_7836);
xor U10406 (N_10406,N_8575,N_9627);
or U10407 (N_10407,N_6868,N_7742);
or U10408 (N_10408,N_5963,N_5345);
nand U10409 (N_10409,N_8965,N_8347);
or U10410 (N_10410,N_9506,N_8485);
xor U10411 (N_10411,N_8978,N_9807);
or U10412 (N_10412,N_5468,N_7575);
or U10413 (N_10413,N_9935,N_6436);
nand U10414 (N_10414,N_8302,N_7858);
xnor U10415 (N_10415,N_7018,N_6273);
nor U10416 (N_10416,N_7367,N_7615);
nor U10417 (N_10417,N_5235,N_7719);
xor U10418 (N_10418,N_9417,N_5062);
nand U10419 (N_10419,N_6221,N_5244);
or U10420 (N_10420,N_9367,N_7736);
or U10421 (N_10421,N_5255,N_9710);
and U10422 (N_10422,N_6169,N_8086);
nor U10423 (N_10423,N_6582,N_5943);
xnor U10424 (N_10424,N_6142,N_5357);
nand U10425 (N_10425,N_6209,N_8543);
or U10426 (N_10426,N_8675,N_6815);
nand U10427 (N_10427,N_8549,N_9447);
xor U10428 (N_10428,N_8823,N_5037);
and U10429 (N_10429,N_6629,N_6568);
nor U10430 (N_10430,N_9083,N_5848);
nand U10431 (N_10431,N_7407,N_6244);
or U10432 (N_10432,N_6478,N_5525);
or U10433 (N_10433,N_9444,N_8755);
or U10434 (N_10434,N_5478,N_8646);
or U10435 (N_10435,N_8349,N_7920);
or U10436 (N_10436,N_8154,N_8684);
xnor U10437 (N_10437,N_5761,N_7612);
and U10438 (N_10438,N_6902,N_7703);
nor U10439 (N_10439,N_6856,N_6440);
and U10440 (N_10440,N_8474,N_8816);
nor U10441 (N_10441,N_7178,N_6563);
nor U10442 (N_10442,N_6197,N_8192);
nor U10443 (N_10443,N_8259,N_8107);
and U10444 (N_10444,N_5070,N_7097);
or U10445 (N_10445,N_7449,N_8165);
and U10446 (N_10446,N_9586,N_6883);
or U10447 (N_10447,N_5512,N_8314);
and U10448 (N_10448,N_7182,N_7751);
xor U10449 (N_10449,N_7348,N_5718);
or U10450 (N_10450,N_7501,N_8571);
nor U10451 (N_10451,N_7456,N_8929);
nand U10452 (N_10452,N_9909,N_5455);
xor U10453 (N_10453,N_6805,N_5523);
nand U10454 (N_10454,N_9691,N_5407);
xnor U10455 (N_10455,N_9495,N_6584);
nand U10456 (N_10456,N_5535,N_6140);
nand U10457 (N_10457,N_8973,N_7141);
xor U10458 (N_10458,N_9760,N_7899);
nor U10459 (N_10459,N_9905,N_5448);
xor U10460 (N_10460,N_8710,N_8344);
or U10461 (N_10461,N_7547,N_5281);
xnor U10462 (N_10462,N_8389,N_8842);
nor U10463 (N_10463,N_9259,N_6653);
and U10464 (N_10464,N_7540,N_5064);
or U10465 (N_10465,N_7794,N_6206);
nor U10466 (N_10466,N_8651,N_6726);
nor U10467 (N_10467,N_8801,N_6229);
and U10468 (N_10468,N_6291,N_5202);
and U10469 (N_10469,N_7645,N_7203);
or U10470 (N_10470,N_7880,N_8223);
xnor U10471 (N_10471,N_8392,N_8883);
or U10472 (N_10472,N_6959,N_5946);
xor U10473 (N_10473,N_8129,N_9221);
or U10474 (N_10474,N_9023,N_7130);
and U10475 (N_10475,N_7513,N_8033);
nand U10476 (N_10476,N_5019,N_7414);
nand U10477 (N_10477,N_6908,N_9336);
and U10478 (N_10478,N_6493,N_8355);
xnor U10479 (N_10479,N_6045,N_7126);
nand U10480 (N_10480,N_9235,N_6624);
xnor U10481 (N_10481,N_9600,N_9892);
nor U10482 (N_10482,N_7602,N_9629);
or U10483 (N_10483,N_9751,N_9510);
or U10484 (N_10484,N_6116,N_5853);
nor U10485 (N_10485,N_5013,N_8046);
xnor U10486 (N_10486,N_9143,N_9991);
nand U10487 (N_10487,N_9286,N_5354);
nor U10488 (N_10488,N_6348,N_7632);
and U10489 (N_10489,N_8459,N_9079);
xnor U10490 (N_10490,N_5396,N_6363);
nor U10491 (N_10491,N_9707,N_8301);
or U10492 (N_10492,N_5695,N_9016);
nor U10493 (N_10493,N_6947,N_8962);
or U10494 (N_10494,N_7475,N_8734);
nand U10495 (N_10495,N_6377,N_8849);
nand U10496 (N_10496,N_7365,N_9037);
nor U10497 (N_10497,N_5729,N_7510);
or U10498 (N_10498,N_7604,N_9676);
and U10499 (N_10499,N_7478,N_8261);
xor U10500 (N_10500,N_7096,N_7038);
or U10501 (N_10501,N_9622,N_5502);
or U10502 (N_10502,N_9045,N_6835);
and U10503 (N_10503,N_8926,N_6993);
nand U10504 (N_10504,N_6933,N_9999);
and U10505 (N_10505,N_9929,N_8855);
xor U10506 (N_10506,N_5570,N_8503);
and U10507 (N_10507,N_8557,N_6474);
xnor U10508 (N_10508,N_6888,N_8454);
nor U10509 (N_10509,N_5187,N_8925);
or U10510 (N_10510,N_5163,N_9494);
nor U10511 (N_10511,N_9386,N_7016);
and U10512 (N_10512,N_6172,N_8834);
nor U10513 (N_10513,N_8091,N_7023);
or U10514 (N_10514,N_7064,N_6335);
xnor U10515 (N_10515,N_9577,N_6047);
xnor U10516 (N_10516,N_7785,N_5323);
or U10517 (N_10517,N_9848,N_6871);
nand U10518 (N_10518,N_9613,N_8145);
or U10519 (N_10519,N_8707,N_6767);
nand U10520 (N_10520,N_8114,N_6382);
nor U10521 (N_10521,N_7637,N_8633);
and U10522 (N_10522,N_7647,N_5118);
nand U10523 (N_10523,N_9928,N_9051);
nor U10524 (N_10524,N_5840,N_9210);
nor U10525 (N_10525,N_7960,N_9213);
and U10526 (N_10526,N_8365,N_8565);
xnor U10527 (N_10527,N_8811,N_9106);
or U10528 (N_10528,N_7969,N_9065);
nor U10529 (N_10529,N_7600,N_6079);
and U10530 (N_10530,N_6181,N_5616);
nand U10531 (N_10531,N_8771,N_5679);
or U10532 (N_10532,N_9947,N_9219);
or U10533 (N_10533,N_6344,N_7721);
nand U10534 (N_10534,N_6074,N_8936);
or U10535 (N_10535,N_8553,N_7410);
or U10536 (N_10536,N_6884,N_5381);
and U10537 (N_10537,N_7806,N_5336);
or U10538 (N_10538,N_8040,N_6213);
nor U10539 (N_10539,N_8536,N_7558);
xor U10540 (N_10540,N_7504,N_6709);
and U10541 (N_10541,N_7400,N_5092);
and U10542 (N_10542,N_9864,N_6345);
xnor U10543 (N_10543,N_9544,N_6892);
or U10544 (N_10544,N_6126,N_6495);
or U10545 (N_10545,N_7271,N_5482);
nand U10546 (N_10546,N_7134,N_6862);
and U10547 (N_10547,N_9558,N_6442);
and U10548 (N_10548,N_5684,N_5819);
and U10549 (N_10549,N_8653,N_8196);
xnor U10550 (N_10550,N_6007,N_5524);
nor U10551 (N_10551,N_5208,N_8366);
nor U10552 (N_10552,N_7882,N_6505);
xnor U10553 (N_10553,N_8597,N_8468);
nor U10554 (N_10554,N_6227,N_9930);
nor U10555 (N_10555,N_8881,N_7531);
nor U10556 (N_10556,N_5807,N_5987);
nor U10557 (N_10557,N_8814,N_6729);
xor U10558 (N_10558,N_5322,N_7404);
xor U10559 (N_10559,N_8669,N_9546);
and U10560 (N_10560,N_6241,N_9440);
or U10561 (N_10561,N_9802,N_7393);
nand U10562 (N_10562,N_5359,N_7457);
nand U10563 (N_10563,N_7698,N_8053);
xor U10564 (N_10564,N_5760,N_7533);
or U10565 (N_10565,N_5680,N_9756);
nor U10566 (N_10566,N_6668,N_6373);
nand U10567 (N_10567,N_8780,N_6033);
or U10568 (N_10568,N_7593,N_5996);
nand U10569 (N_10569,N_8335,N_6473);
or U10570 (N_10570,N_8324,N_7076);
nor U10571 (N_10571,N_9959,N_5245);
nand U10572 (N_10572,N_5994,N_7834);
nor U10573 (N_10573,N_7759,N_6825);
xnor U10574 (N_10574,N_9428,N_8279);
nand U10575 (N_10575,N_5108,N_8721);
or U10576 (N_10576,N_7254,N_5368);
xor U10577 (N_10577,N_5153,N_8715);
xor U10578 (N_10578,N_8616,N_9123);
or U10579 (N_10579,N_9871,N_5282);
and U10580 (N_10580,N_8094,N_9024);
xnor U10581 (N_10581,N_8703,N_6602);
or U10582 (N_10582,N_5697,N_6641);
xor U10583 (N_10583,N_5367,N_7077);
and U10584 (N_10584,N_8368,N_7993);
and U10585 (N_10585,N_6087,N_8548);
nand U10586 (N_10586,N_9128,N_5017);
nand U10587 (N_10587,N_9781,N_5757);
xnor U10588 (N_10588,N_6789,N_9327);
nor U10589 (N_10589,N_7274,N_5543);
or U10590 (N_10590,N_8650,N_8902);
and U10591 (N_10591,N_9198,N_7034);
nor U10592 (N_10592,N_7136,N_6349);
nand U10593 (N_10593,N_6459,N_8494);
nor U10594 (N_10594,N_6454,N_7166);
nand U10595 (N_10595,N_5806,N_8972);
nor U10596 (N_10596,N_7595,N_7903);
xnor U10597 (N_10597,N_5519,N_8862);
and U10598 (N_10598,N_7236,N_5386);
and U10599 (N_10599,N_5673,N_7906);
and U10600 (N_10600,N_9744,N_9356);
xor U10601 (N_10601,N_8078,N_7838);
xor U10602 (N_10602,N_5376,N_8184);
nor U10603 (N_10603,N_9239,N_5240);
nand U10604 (N_10604,N_7310,N_5647);
or U10605 (N_10605,N_7133,N_7942);
nor U10606 (N_10606,N_6731,N_9177);
and U10607 (N_10607,N_8100,N_6055);
and U10608 (N_10608,N_5385,N_6739);
or U10609 (N_10609,N_8160,N_5112);
xnor U10610 (N_10610,N_5756,N_5585);
nand U10611 (N_10611,N_6380,N_9889);
or U10612 (N_10612,N_8027,N_9987);
xor U10613 (N_10613,N_7716,N_8950);
nor U10614 (N_10614,N_6256,N_9111);
or U10615 (N_10615,N_6261,N_8342);
xor U10616 (N_10616,N_6547,N_7896);
or U10617 (N_10617,N_9458,N_9661);
nand U10618 (N_10618,N_8385,N_6354);
or U10619 (N_10619,N_7546,N_5937);
or U10620 (N_10620,N_9851,N_7544);
nand U10621 (N_10621,N_9653,N_6305);
or U10622 (N_10622,N_9522,N_9432);
nand U10623 (N_10623,N_6481,N_7201);
nor U10624 (N_10624,N_5236,N_9256);
and U10625 (N_10625,N_7589,N_7356);
nand U10626 (N_10626,N_7854,N_8070);
or U10627 (N_10627,N_5489,N_9479);
nor U10628 (N_10628,N_7591,N_8367);
xor U10629 (N_10629,N_6167,N_9469);
or U10630 (N_10630,N_5866,N_6220);
nand U10631 (N_10631,N_7729,N_8666);
nor U10632 (N_10632,N_7306,N_6930);
xnor U10633 (N_10633,N_9354,N_7024);
and U10634 (N_10634,N_9116,N_6134);
or U10635 (N_10635,N_6831,N_8511);
xor U10636 (N_10636,N_7187,N_6306);
xnor U10637 (N_10637,N_8994,N_8641);
xor U10638 (N_10638,N_7878,N_9026);
xor U10639 (N_10639,N_9197,N_9923);
or U10640 (N_10640,N_5696,N_6956);
xor U10641 (N_10641,N_5830,N_5746);
and U10642 (N_10642,N_6238,N_9438);
nor U10643 (N_10643,N_8764,N_9172);
and U10644 (N_10644,N_5270,N_8178);
and U10645 (N_10645,N_8146,N_8079);
nor U10646 (N_10646,N_9130,N_6392);
nor U10647 (N_10647,N_7140,N_7432);
or U10648 (N_10648,N_6801,N_8148);
or U10649 (N_10649,N_6557,N_8628);
nand U10650 (N_10650,N_9519,N_5377);
xnor U10651 (N_10651,N_8762,N_6932);
nand U10652 (N_10652,N_5159,N_7900);
nand U10653 (N_10653,N_5201,N_8237);
nor U10654 (N_10654,N_5311,N_9637);
nor U10655 (N_10655,N_5341,N_9236);
nor U10656 (N_10656,N_9780,N_9105);
and U10657 (N_10657,N_6489,N_5636);
and U10658 (N_10658,N_9723,N_6542);
nand U10659 (N_10659,N_7167,N_7273);
xor U10660 (N_10660,N_5052,N_8619);
nor U10661 (N_10661,N_5094,N_6311);
nand U10662 (N_10662,N_7360,N_8819);
nand U10663 (N_10663,N_6317,N_8527);
nor U10664 (N_10664,N_9837,N_9903);
and U10665 (N_10665,N_7582,N_6654);
and U10666 (N_10666,N_5633,N_9092);
or U10667 (N_10667,N_7859,N_6925);
or U10668 (N_10668,N_8797,N_7033);
nand U10669 (N_10669,N_9809,N_9145);
or U10670 (N_10670,N_5045,N_5628);
nand U10671 (N_10671,N_8609,N_6746);
nand U10672 (N_10672,N_7327,N_8269);
nor U10673 (N_10673,N_9373,N_7743);
or U10674 (N_10674,N_9978,N_7853);
and U10675 (N_10675,N_5531,N_8442);
nand U10676 (N_10676,N_6420,N_6081);
nand U10677 (N_10677,N_9641,N_5484);
or U10678 (N_10678,N_9437,N_8706);
xnor U10679 (N_10679,N_7492,N_8051);
or U10680 (N_10680,N_9509,N_7092);
or U10681 (N_10681,N_9511,N_7581);
and U10682 (N_10682,N_7294,N_5638);
xor U10683 (N_10683,N_6979,N_9667);
or U10684 (N_10684,N_8333,N_8660);
and U10685 (N_10685,N_5330,N_9927);
or U10686 (N_10686,N_7627,N_9914);
or U10687 (N_10687,N_5488,N_7638);
and U10688 (N_10688,N_7707,N_9820);
or U10689 (N_10689,N_8267,N_8899);
xor U10690 (N_10690,N_7514,N_6994);
nor U10691 (N_10691,N_5470,N_8222);
or U10692 (N_10692,N_7644,N_6413);
xnor U10693 (N_10693,N_7215,N_5266);
xor U10694 (N_10694,N_6405,N_8750);
nand U10695 (N_10695,N_7144,N_8256);
or U10696 (N_10696,N_5423,N_5378);
nor U10697 (N_10697,N_7129,N_8170);
xor U10698 (N_10698,N_5947,N_7013);
and U10699 (N_10699,N_8917,N_8353);
and U10700 (N_10700,N_5150,N_7998);
nand U10701 (N_10701,N_9175,N_9395);
nor U10702 (N_10702,N_7654,N_8021);
and U10703 (N_10703,N_7694,N_6592);
nand U10704 (N_10704,N_6623,N_9477);
and U10705 (N_10705,N_5852,N_7386);
and U10706 (N_10706,N_5741,N_7039);
nor U10707 (N_10707,N_8638,N_5021);
or U10708 (N_10708,N_9340,N_8585);
nand U10709 (N_10709,N_5212,N_8533);
nor U10710 (N_10710,N_9769,N_6781);
or U10711 (N_10711,N_5643,N_8860);
xnor U10712 (N_10712,N_5181,N_6268);
and U10713 (N_10713,N_8538,N_8988);
nand U10714 (N_10714,N_7652,N_9487);
or U10715 (N_10715,N_5220,N_5540);
xnor U10716 (N_10716,N_8251,N_9869);
and U10717 (N_10717,N_5541,N_8306);
and U10718 (N_10718,N_5750,N_5480);
xnor U10719 (N_10719,N_5347,N_9747);
xor U10720 (N_10720,N_6395,N_8473);
xor U10721 (N_10721,N_9761,N_9505);
nor U10722 (N_10722,N_7031,N_8249);
and U10723 (N_10723,N_6418,N_6890);
nand U10724 (N_10724,N_6239,N_6940);
and U10725 (N_10725,N_8140,N_9740);
nor U10726 (N_10726,N_8803,N_8667);
and U10727 (N_10727,N_7800,N_7188);
nor U10728 (N_10728,N_7814,N_6588);
nand U10729 (N_10729,N_6723,N_5940);
and U10730 (N_10730,N_7622,N_9243);
or U10731 (N_10731,N_7270,N_8130);
xor U10732 (N_10732,N_7728,N_9160);
nand U10733 (N_10733,N_7278,N_6617);
nand U10734 (N_10734,N_8812,N_6995);
xor U10735 (N_10735,N_6110,N_8326);
and U10736 (N_10736,N_6515,N_8395);
or U10737 (N_10737,N_9404,N_8671);
xnor U10738 (N_10738,N_9081,N_6475);
xor U10739 (N_10739,N_5780,N_5878);
and U10740 (N_10740,N_6130,N_6274);
and U10741 (N_10741,N_8977,N_5509);
nor U10742 (N_10742,N_8478,N_7434);
xor U10743 (N_10743,N_5621,N_9308);
nand U10744 (N_10744,N_5698,N_5962);
and U10745 (N_10745,N_7499,N_9025);
nor U10746 (N_10746,N_7947,N_5796);
xnor U10747 (N_10747,N_7131,N_8447);
nor U10748 (N_10748,N_8069,N_6875);
and U10749 (N_10749,N_6411,N_9454);
xnor U10750 (N_10750,N_7091,N_8800);
and U10751 (N_10751,N_7889,N_6445);
xnor U10752 (N_10752,N_8841,N_9595);
nand U10753 (N_10753,N_8015,N_6704);
or U10754 (N_10754,N_8687,N_9486);
and U10755 (N_10755,N_9167,N_7682);
and U10756 (N_10756,N_9392,N_5205);
or U10757 (N_10757,N_5556,N_9391);
nand U10758 (N_10758,N_7338,N_9941);
nor U10759 (N_10759,N_8827,N_6898);
and U10760 (N_10760,N_8491,N_7948);
or U10761 (N_10761,N_8898,N_7821);
and U10762 (N_10762,N_5284,N_7692);
and U10763 (N_10763,N_8195,N_7158);
nor U10764 (N_10764,N_8603,N_7494);
nand U10765 (N_10765,N_6594,N_5795);
xor U10766 (N_10766,N_8746,N_8093);
nor U10767 (N_10767,N_9866,N_8513);
xor U10768 (N_10768,N_5664,N_7235);
nor U10769 (N_10769,N_6879,N_6841);
and U10770 (N_10770,N_5151,N_5428);
xor U10771 (N_10771,N_6882,N_5460);
nand U10772 (N_10772,N_7101,N_8991);
or U10773 (N_10773,N_5644,N_7748);
nor U10774 (N_10774,N_6136,N_9685);
and U10775 (N_10775,N_6210,N_5095);
nor U10776 (N_10776,N_7072,N_5442);
nand U10777 (N_10777,N_9986,N_5364);
nor U10778 (N_10778,N_6375,N_5514);
nand U10779 (N_10779,N_8697,N_9028);
nor U10780 (N_10780,N_8655,N_5902);
xor U10781 (N_10781,N_6722,N_6494);
or U10782 (N_10782,N_8594,N_6681);
or U10783 (N_10783,N_8958,N_8604);
nor U10784 (N_10784,N_9733,N_8031);
or U10785 (N_10785,N_8922,N_5885);
and U10786 (N_10786,N_8934,N_8283);
or U10787 (N_10787,N_6024,N_5230);
xor U10788 (N_10788,N_7511,N_5737);
or U10789 (N_10789,N_9535,N_5265);
xor U10790 (N_10790,N_9271,N_7496);
nand U10791 (N_10791,N_6670,N_8396);
and U10792 (N_10792,N_6538,N_8203);
xnor U10793 (N_10793,N_9748,N_9652);
nand U10794 (N_10794,N_6379,N_5911);
and U10795 (N_10795,N_9767,N_5794);
and U10796 (N_10796,N_5555,N_8795);
and U10797 (N_10797,N_8429,N_8545);
xnor U10798 (N_10798,N_5861,N_8309);
and U10799 (N_10799,N_9288,N_9041);
or U10800 (N_10800,N_6460,N_8743);
nor U10801 (N_10801,N_9215,N_7257);
or U10802 (N_10802,N_5552,N_5659);
or U10803 (N_10803,N_7918,N_6362);
or U10804 (N_10804,N_8471,N_5302);
nor U10805 (N_10805,N_7875,N_5024);
or U10806 (N_10806,N_8218,N_8544);
or U10807 (N_10807,N_9610,N_9449);
xnor U10808 (N_10808,N_8084,N_6577);
or U10809 (N_10809,N_5995,N_6330);
and U10810 (N_10810,N_5574,N_8009);
or U10811 (N_10811,N_5379,N_5298);
and U10812 (N_10812,N_7299,N_9969);
or U10813 (N_10813,N_5184,N_8417);
nand U10814 (N_10814,N_6794,N_8085);
nand U10815 (N_10815,N_7326,N_8312);
xor U10816 (N_10816,N_9325,N_9353);
xor U10817 (N_10817,N_6591,N_9317);
xnor U10818 (N_10818,N_8551,N_7775);
nor U10819 (N_10819,N_6889,N_7463);
or U10820 (N_10820,N_9975,N_5660);
nor U10821 (N_10821,N_6605,N_9739);
nand U10822 (N_10822,N_7760,N_9015);
or U10823 (N_10823,N_7590,N_5199);
and U10824 (N_10824,N_5211,N_6613);
or U10825 (N_10825,N_7320,N_5825);
or U10826 (N_10826,N_5646,N_9341);
and U10827 (N_10827,N_6009,N_7490);
nand U10828 (N_10828,N_7636,N_8134);
nor U10829 (N_10829,N_9158,N_6015);
or U10830 (N_10830,N_8998,N_5492);
nand U10831 (N_10831,N_8554,N_5820);
xnor U10832 (N_10832,N_5495,N_5485);
xor U10833 (N_10833,N_5888,N_9431);
nand U10834 (N_10834,N_9548,N_5674);
or U10835 (N_10835,N_5609,N_7664);
or U10836 (N_10836,N_8050,N_6876);
or U10837 (N_10837,N_7379,N_5125);
or U10838 (N_10838,N_5753,N_7962);
nor U10839 (N_10839,N_5973,N_7628);
nand U10840 (N_10840,N_5011,N_8288);
or U10841 (N_10841,N_9602,N_6857);
nor U10842 (N_10842,N_5657,N_7479);
nand U10843 (N_10843,N_9265,N_9743);
nor U10844 (N_10844,N_9278,N_9896);
or U10845 (N_10845,N_6900,N_9709);
nand U10846 (N_10846,N_5267,N_6539);
xor U10847 (N_10847,N_9714,N_7199);
and U10848 (N_10848,N_6526,N_8807);
nand U10849 (N_10849,N_9593,N_6370);
and U10850 (N_10850,N_5164,N_6314);
and U10851 (N_10851,N_8952,N_5565);
nand U10852 (N_10852,N_7385,N_8745);
or U10853 (N_10853,N_8626,N_6019);
or U10854 (N_10854,N_5656,N_7939);
or U10855 (N_10855,N_9018,N_5534);
nand U10856 (N_10856,N_5466,N_9594);
nor U10857 (N_10857,N_8408,N_9225);
nand U10858 (N_10858,N_6783,N_5251);
and U10859 (N_10859,N_7825,N_5667);
nor U10860 (N_10860,N_9450,N_5047);
or U10861 (N_10861,N_5190,N_7282);
nand U10862 (N_10862,N_5711,N_6063);
nor U10863 (N_10863,N_5034,N_9699);
nor U10864 (N_10864,N_5287,N_9075);
nor U10865 (N_10865,N_5877,N_6378);
xnor U10866 (N_10866,N_5744,N_5049);
or U10867 (N_10867,N_7848,N_9556);
xor U10868 (N_10868,N_5809,N_8558);
xnor U10869 (N_10869,N_8407,N_6957);
xor U10870 (N_10870,N_7468,N_6907);
or U10871 (N_10871,N_6535,N_7678);
xnor U10872 (N_10872,N_7985,N_5941);
or U10873 (N_10873,N_6153,N_6470);
or U10874 (N_10874,N_6714,N_7656);
nand U10875 (N_10875,N_5821,N_6977);
nand U10876 (N_10876,N_7392,N_6999);
and U10877 (N_10877,N_6326,N_5847);
nor U10878 (N_10878,N_8610,N_8090);
or U10879 (N_10879,N_7507,N_9670);
nor U10880 (N_10880,N_7009,N_7170);
or U10881 (N_10881,N_6909,N_5483);
nand U10882 (N_10882,N_8246,N_7100);
and U10883 (N_10883,N_9038,N_8440);
nand U10884 (N_10884,N_6798,N_8016);
or U10885 (N_10885,N_7734,N_5289);
nor U10886 (N_10886,N_7482,N_5147);
nor U10887 (N_10887,N_6302,N_9700);
and U10888 (N_10888,N_8416,N_8542);
nor U10889 (N_10889,N_8670,N_9473);
nand U10890 (N_10890,N_5471,N_9880);
or U10891 (N_10891,N_9838,N_5063);
and U10892 (N_10892,N_5170,N_7657);
xnor U10893 (N_10893,N_7246,N_7022);
or U10894 (N_10894,N_8736,N_7738);
xnor U10895 (N_10895,N_9682,N_8636);
or U10896 (N_10896,N_7573,N_8752);
and U10897 (N_10897,N_9816,N_6457);
nand U10898 (N_10898,N_7964,N_9636);
or U10899 (N_10899,N_5770,N_6128);
nor U10900 (N_10900,N_5179,N_7352);
nand U10901 (N_10901,N_6797,N_6807);
nand U10902 (N_10902,N_9203,N_9906);
nor U10903 (N_10903,N_6854,N_7269);
nor U10904 (N_10904,N_7082,N_9725);
or U10905 (N_10905,N_7127,N_8711);
nor U10906 (N_10906,N_8304,N_9267);
and U10907 (N_10907,N_7497,N_5721);
nor U10908 (N_10908,N_8011,N_6057);
xor U10909 (N_10909,N_9453,N_9648);
nand U10910 (N_10910,N_9008,N_5473);
xor U10911 (N_10911,N_9642,N_8612);
or U10912 (N_10912,N_7840,N_9401);
or U10913 (N_10913,N_9104,N_5935);
nand U10914 (N_10914,N_7867,N_7681);
and U10915 (N_10915,N_8720,N_8933);
xnor U10916 (N_10916,N_8847,N_7218);
and U10917 (N_10917,N_9616,N_9800);
or U10918 (N_10918,N_5054,N_9212);
nand U10919 (N_10919,N_5624,N_7300);
xnor U10920 (N_10920,N_8836,N_7355);
or U10921 (N_10921,N_9068,N_9088);
or U10922 (N_10922,N_5613,N_5256);
nor U10923 (N_10923,N_8169,N_8698);
xor U10924 (N_10924,N_9589,N_8488);
or U10925 (N_10925,N_8089,N_9300);
xor U10926 (N_10926,N_5343,N_6992);
xnor U10927 (N_10927,N_8108,N_7714);
xnor U10928 (N_10928,N_9189,N_9095);
nand U10929 (N_10929,N_7966,N_9496);
and U10930 (N_10930,N_5837,N_5530);
or U10931 (N_10931,N_7469,N_5040);
nor U10932 (N_10932,N_7244,N_8217);
nand U10933 (N_10933,N_9294,N_7804);
or U10934 (N_10934,N_6661,N_5018);
or U10935 (N_10935,N_5315,N_5000);
nand U10936 (N_10936,N_5046,N_7279);
nand U10937 (N_10937,N_9319,N_6492);
and U10938 (N_10938,N_5447,N_6061);
and U10939 (N_10939,N_9246,N_9078);
or U10940 (N_10940,N_5399,N_9010);
or U10941 (N_10941,N_5157,N_5067);
nand U10942 (N_10942,N_9021,N_5453);
and U10943 (N_10943,N_6625,N_5954);
nor U10944 (N_10944,N_7342,N_6185);
and U10945 (N_10945,N_5429,N_7227);
nand U10946 (N_10946,N_9638,N_7556);
and U10947 (N_10947,N_7155,N_8161);
nor U10948 (N_10948,N_6601,N_8724);
xnor U10949 (N_10949,N_7677,N_9984);
xnor U10950 (N_10950,N_9994,N_9900);
nand U10951 (N_10951,N_7275,N_5736);
and U10952 (N_10952,N_7841,N_9979);
xor U10953 (N_10953,N_8299,N_6401);
or U10954 (N_10954,N_8492,N_8719);
and U10955 (N_10955,N_8260,N_8004);
xnor U10956 (N_10956,N_8679,N_6885);
xnor U10957 (N_10957,N_5445,N_8329);
xnor U10958 (N_10958,N_5261,N_7592);
nor U10959 (N_10959,N_8370,N_5373);
or U10960 (N_10960,N_7245,N_9050);
nand U10961 (N_10961,N_9094,N_6031);
and U10962 (N_10962,N_6071,N_8835);
xor U10963 (N_10963,N_8939,N_9966);
nand U10964 (N_10964,N_5620,N_8910);
nand U10965 (N_10965,N_6834,N_8030);
nand U10966 (N_10966,N_6725,N_7169);
or U10967 (N_10967,N_7713,N_6289);
nor U10968 (N_10968,N_8689,N_6325);
and U10969 (N_10969,N_7988,N_6294);
nor U10970 (N_10970,N_8580,N_5926);
nor U10971 (N_10971,N_9362,N_6508);
nor U10972 (N_10972,N_9074,N_8895);
xor U10973 (N_10973,N_9304,N_5560);
nand U10974 (N_10974,N_9995,N_5920);
nand U10975 (N_10975,N_6484,N_7701);
xnor U10976 (N_10976,N_5068,N_9377);
or U10977 (N_10977,N_7437,N_6899);
nor U10978 (N_10978,N_6913,N_5677);
nor U10979 (N_10979,N_7157,N_8399);
or U10980 (N_10980,N_9621,N_9983);
or U10981 (N_10981,N_5601,N_9492);
nand U10982 (N_10982,N_5437,N_6677);
xor U10983 (N_10983,N_6684,N_5709);
nand U10984 (N_10984,N_6711,N_5035);
and U10985 (N_10985,N_5893,N_9462);
xnor U10986 (N_10986,N_5771,N_9872);
nor U10987 (N_10987,N_9378,N_9402);
xnor U10988 (N_10988,N_7051,N_6387);
nand U10989 (N_10989,N_8357,N_5391);
and U10990 (N_10990,N_8379,N_8132);
or U10991 (N_10991,N_8263,N_8947);
or U10992 (N_10992,N_6282,N_8983);
or U10993 (N_10993,N_5440,N_6599);
xnor U10994 (N_10994,N_8204,N_8443);
or U10995 (N_10995,N_9435,N_9089);
nand U10996 (N_10996,N_8343,N_5444);
nand U10997 (N_10997,N_5945,N_5897);
or U10998 (N_10998,N_7151,N_6158);
and U10999 (N_10999,N_5755,N_9249);
or U11000 (N_11000,N_9863,N_7249);
xor U11001 (N_11001,N_5991,N_9680);
nand U11002 (N_11002,N_7726,N_9575);
nor U11003 (N_11003,N_7505,N_9001);
and U11004 (N_11004,N_9463,N_8971);
xor U11005 (N_11005,N_9264,N_5814);
nor U11006 (N_11006,N_7118,N_7491);
nand U11007 (N_11007,N_8414,N_8391);
and U11008 (N_11008,N_5592,N_9405);
and U11009 (N_11009,N_9985,N_6262);
nand U11010 (N_11010,N_6170,N_5023);
nand U11011 (N_11011,N_6808,N_5020);
nand U11012 (N_11012,N_7329,N_7314);
or U11013 (N_11013,N_7683,N_9165);
nand U11014 (N_11014,N_7845,N_5397);
xor U11015 (N_11015,N_8293,N_9268);
xor U11016 (N_11016,N_5909,N_5102);
xnor U11017 (N_11017,N_6521,N_5180);
xor U11018 (N_11018,N_5513,N_5431);
or U11019 (N_11019,N_5785,N_7200);
xnor U11020 (N_11020,N_6784,N_8133);
nor U11021 (N_11021,N_5615,N_7221);
or U11022 (N_11022,N_6860,N_9504);
xnor U11023 (N_11023,N_5701,N_6679);
nor U11024 (N_11024,N_9668,N_9536);
nor U11025 (N_11025,N_5551,N_9359);
or U11026 (N_11026,N_9957,N_9810);
or U11027 (N_11027,N_5938,N_5459);
nand U11028 (N_11028,N_6151,N_9711);
nor U11029 (N_11029,N_6034,N_6143);
nor U11030 (N_11030,N_6791,N_5841);
nand U11031 (N_11031,N_9583,N_9113);
nor U11032 (N_11032,N_9216,N_5913);
or U11033 (N_11033,N_9475,N_6980);
xnor U11034 (N_11034,N_7344,N_6590);
and U11035 (N_11035,N_8469,N_5073);
xor U11036 (N_11036,N_6958,N_9696);
xor U11037 (N_11037,N_8802,N_5128);
nand U11038 (N_11038,N_9276,N_8510);
nor U11039 (N_11039,N_5614,N_5635);
and U11040 (N_11040,N_6705,N_7852);
nor U11041 (N_11041,N_9672,N_8985);
and U11042 (N_11042,N_5712,N_9542);
nand U11043 (N_11043,N_6069,N_9032);
nand U11044 (N_11044,N_6246,N_9389);
nor U11045 (N_11045,N_8008,N_5980);
xor U11046 (N_11046,N_6432,N_5259);
nor U11047 (N_11047,N_5829,N_5237);
nand U11048 (N_11048,N_6843,N_5493);
nor U11049 (N_11049,N_8295,N_7371);
nor U11050 (N_11050,N_5196,N_6085);
or U11051 (N_11051,N_9604,N_5085);
nor U11052 (N_11052,N_8313,N_6837);
nor U11053 (N_11053,N_5400,N_5166);
nor U11054 (N_11054,N_8405,N_5007);
or U11055 (N_11055,N_6919,N_8318);
nor U11056 (N_11056,N_6838,N_7459);
nand U11057 (N_11057,N_6477,N_5452);
or U11058 (N_11058,N_7473,N_5949);
and U11059 (N_11059,N_6123,N_9823);
xor U11060 (N_11060,N_5059,N_5148);
xnor U11061 (N_11061,N_7791,N_5836);
nor U11062 (N_11062,N_7995,N_5109);
or U11063 (N_11063,N_9125,N_8976);
nand U11064 (N_11064,N_5139,N_9188);
or U11065 (N_11065,N_7108,N_8824);
and U11066 (N_11066,N_8315,N_9142);
xnor U11067 (N_11067,N_6490,N_9248);
and U11068 (N_11068,N_9977,N_5499);
xnor U11069 (N_11069,N_8817,N_8946);
or U11070 (N_11070,N_8942,N_5285);
nor U11071 (N_11071,N_9943,N_8567);
and U11072 (N_11072,N_5292,N_6211);
nand U11073 (N_11073,N_9207,N_9731);
nand U11074 (N_11074,N_5881,N_9776);
or U11075 (N_11075,N_7217,N_8428);
xnor U11076 (N_11076,N_6003,N_7250);
xor U11077 (N_11077,N_7228,N_9758);
and U11078 (N_11078,N_7307,N_9588);
nor U11079 (N_11079,N_8966,N_6394);
xor U11080 (N_11080,N_6426,N_6026);
xnor U11081 (N_11081,N_5704,N_9729);
nand U11082 (N_11082,N_7543,N_6574);
nand U11083 (N_11083,N_8799,N_8077);
xor U11084 (N_11084,N_7390,N_9919);
nand U11085 (N_11085,N_5532,N_7398);
and U11086 (N_11086,N_7762,N_5790);
or U11087 (N_11087,N_7119,N_6765);
xor U11088 (N_11088,N_7139,N_6148);
nor U11089 (N_11089,N_7725,N_9701);
nand U11090 (N_11090,N_7149,N_5491);
nand U11091 (N_11091,N_7665,N_7471);
nand U11092 (N_11092,N_5424,N_9963);
nand U11093 (N_11093,N_9818,N_8708);
or U11094 (N_11094,N_7884,N_7138);
nand U11095 (N_11095,N_5195,N_5767);
xor U11096 (N_11096,N_8206,N_5625);
nor U11097 (N_11097,N_5041,N_6050);
nor U11098 (N_11098,N_8903,N_9513);
xor U11099 (N_11099,N_9790,N_8798);
nand U11100 (N_11100,N_8796,N_6926);
nand U11101 (N_11101,N_5280,N_6098);
and U11102 (N_11102,N_7551,N_9164);
xnor U11103 (N_11103,N_5655,N_6156);
xor U11104 (N_11104,N_9380,N_7464);
and U11105 (N_11105,N_8390,N_6333);
and U11106 (N_11106,N_5469,N_7113);
nor U11107 (N_11107,N_6859,N_5079);
and U11108 (N_11108,N_5970,N_8289);
nor U11109 (N_11109,N_9066,N_7606);
xor U11110 (N_11110,N_7164,N_9415);
and U11111 (N_11111,N_8207,N_9324);
nand U11112 (N_11112,N_9715,N_8756);
xnor U11113 (N_11113,N_5127,N_9612);
xnor U11114 (N_11114,N_7109,N_5369);
xnor U11115 (N_11115,N_9819,N_5160);
nor U11116 (N_11116,N_8875,N_8384);
xnor U11117 (N_11117,N_8125,N_5605);
or U11118 (N_11118,N_7213,N_9534);
and U11119 (N_11119,N_5069,N_8286);
or U11120 (N_11120,N_9570,N_8005);
or U11121 (N_11121,N_8047,N_7349);
nor U11122 (N_11122,N_8339,N_7815);
nor U11123 (N_11123,N_6114,N_6298);
and U11124 (N_11124,N_6105,N_7353);
nor U11125 (N_11125,N_9883,N_9459);
nor U11126 (N_11126,N_5800,N_9794);
or U11127 (N_11127,N_9808,N_6016);
or U11128 (N_11128,N_8681,N_8705);
xnor U11129 (N_11129,N_6281,N_7776);
and U11130 (N_11130,N_5654,N_5027);
nor U11131 (N_11131,N_5811,N_9879);
and U11132 (N_11132,N_5572,N_5066);
nor U11133 (N_11133,N_8210,N_5719);
nor U11134 (N_11134,N_7584,N_9631);
nor U11135 (N_11135,N_5793,N_7026);
and U11136 (N_11136,N_8714,N_8419);
xnor U11137 (N_11137,N_8944,N_9806);
or U11138 (N_11138,N_9091,N_9241);
or U11139 (N_11139,N_5028,N_9852);
nor U11140 (N_11140,N_6011,N_6249);
and U11141 (N_11141,N_5782,N_5441);
nor U11142 (N_11142,N_6741,N_5912);
nor U11143 (N_11143,N_8837,N_7562);
nor U11144 (N_11144,N_8112,N_9321);
and U11145 (N_11145,N_7174,N_8155);
nor U11146 (N_11146,N_8006,N_6812);
xor U11147 (N_11147,N_6036,N_8239);
or U11148 (N_11148,N_8741,N_5479);
or U11149 (N_11149,N_6688,N_9446);
nand U11150 (N_11150,N_7576,N_7206);
or U11151 (N_11151,N_9077,N_6821);
nor U11152 (N_11152,N_6866,N_8067);
xnor U11153 (N_11153,N_9530,N_9150);
nor U11154 (N_11154,N_9420,N_8081);
or U11155 (N_11155,N_5792,N_7240);
nand U11156 (N_11156,N_9206,N_7438);
or U11157 (N_11157,N_8866,N_9136);
xnor U11158 (N_11158,N_5218,N_9557);
xnor U11159 (N_11159,N_5582,N_6975);
xnor U11160 (N_11160,N_5243,N_9882);
xor U11161 (N_11161,N_5327,N_9884);
nand U11162 (N_11162,N_7932,N_8378);
and U11163 (N_11163,N_8602,N_8749);
xnor U11164 (N_11164,N_6437,N_7225);
nand U11165 (N_11165,N_6342,N_9387);
and U11166 (N_11166,N_6403,N_9253);
or U11167 (N_11167,N_5464,N_6464);
and U11168 (N_11168,N_5015,N_8767);
and U11169 (N_11169,N_7945,N_6989);
or U11170 (N_11170,N_9328,N_9040);
nand U11171 (N_11171,N_7324,N_7266);
and U11172 (N_11172,N_9840,N_8863);
nand U11173 (N_11173,N_6622,N_9409);
nand U11174 (N_11174,N_5300,N_9858);
and U11175 (N_11175,N_6453,N_6954);
nor U11176 (N_11176,N_9591,N_7180);
nor U11177 (N_11177,N_5286,N_6929);
nor U11178 (N_11178,N_5250,N_6657);
xnor U11179 (N_11179,N_8829,N_5639);
xor U11180 (N_11180,N_9424,N_6005);
and U11181 (N_11181,N_5642,N_5006);
or U11182 (N_11182,N_5168,N_7413);
or U11183 (N_11183,N_6386,N_9951);
xor U11184 (N_11184,N_8455,N_9357);
and U11185 (N_11185,N_6133,N_9399);
xnor U11186 (N_11186,N_9894,N_8122);
xor U11187 (N_11187,N_8076,N_7004);
xnor U11188 (N_11188,N_5101,N_5486);
nand U11189 (N_11189,N_5818,N_7536);
nand U11190 (N_11190,N_6840,N_7611);
xor U11191 (N_11191,N_5906,N_6728);
nor U11192 (N_11192,N_6216,N_9990);
nor U11193 (N_11193,N_5670,N_8054);
or U11194 (N_11194,N_9430,N_6607);
nand U11195 (N_11195,N_9775,N_9523);
nor U11196 (N_11196,N_9623,N_8738);
or U11197 (N_11197,N_8052,N_8068);
or U11198 (N_11198,N_5272,N_9006);
and U11199 (N_11199,N_6971,N_7498);
nand U11200 (N_11200,N_7957,N_8643);
nor U11201 (N_11201,N_5904,N_5869);
nand U11202 (N_11202,N_8951,N_5476);
nand U11203 (N_11203,N_6283,N_8214);
and U11204 (N_11204,N_5849,N_6285);
xnor U11205 (N_11205,N_9601,N_6293);
nand U11206 (N_11206,N_6703,N_5742);
xor U11207 (N_11207,N_9907,N_7313);
nor U11208 (N_11208,N_6328,N_6219);
or U11209 (N_11209,N_9855,N_9870);
and U11210 (N_11210,N_9229,N_5271);
nand U11211 (N_11211,N_9762,N_6732);
nand U11212 (N_11212,N_9298,N_5313);
xor U11213 (N_11213,N_6035,N_8381);
or U11214 (N_11214,N_8908,N_7125);
and U11215 (N_11215,N_9551,N_8020);
and U11216 (N_11216,N_5033,N_6717);
and U11217 (N_11217,N_8294,N_8028);
nor U11218 (N_11218,N_6792,N_9411);
xor U11219 (N_11219,N_9371,N_5901);
and U11220 (N_11220,N_9960,N_9649);
xnor U11221 (N_11221,N_8880,N_8768);
and U11222 (N_11222,N_6388,N_7979);
and U11223 (N_11223,N_6660,N_7156);
or U11224 (N_11224,N_7922,N_9155);
nand U11225 (N_11225,N_7445,N_5388);
xor U11226 (N_11226,N_6687,N_7667);
nand U11227 (N_11227,N_9129,N_8647);
nand U11228 (N_11228,N_6645,N_9881);
xnor U11229 (N_11229,N_8038,N_9674);
nor U11230 (N_11230,N_8744,N_6359);
or U11231 (N_11231,N_9499,N_7088);
nor U11232 (N_11232,N_6516,N_8097);
xor U11233 (N_11233,N_7530,N_8423);
xor U11234 (N_11234,N_7477,N_7484);
and U11235 (N_11235,N_8546,N_8685);
or U11236 (N_11236,N_5306,N_8905);
nand U11237 (N_11237,N_8509,N_8773);
xor U11238 (N_11238,N_6865,N_9774);
nor U11239 (N_11239,N_8753,N_5339);
nor U11240 (N_11240,N_8430,N_5334);
and U11241 (N_11241,N_7085,N_7209);
xor U11242 (N_11242,N_8317,N_5842);
xnor U11243 (N_11243,N_5982,N_9915);
nor U11244 (N_11244,N_5249,N_8189);
nor U11245 (N_11245,N_6630,N_9201);
nor U11246 (N_11246,N_6561,N_8539);
xnor U11247 (N_11247,N_7697,N_5351);
nor U11248 (N_11248,N_7690,N_9528);
nand U11249 (N_11249,N_6358,N_6090);
and U11250 (N_11250,N_6044,N_6942);
nand U11251 (N_11251,N_5603,N_5215);
and U11252 (N_11252,N_8435,N_9706);
or U11253 (N_11253,N_7006,N_6787);
nor U11254 (N_11254,N_7451,N_5301);
or U11255 (N_11255,N_5456,N_7293);
or U11256 (N_11256,N_9004,N_6918);
and U11257 (N_11257,N_9644,N_7143);
and U11258 (N_11258,N_5239,N_8656);
or U11259 (N_11259,N_5846,N_8375);
nand U11260 (N_11260,N_8967,N_5496);
nor U11261 (N_11261,N_5773,N_7913);
xnor U11262 (N_11262,N_5008,N_9096);
and U11263 (N_11263,N_8739,N_5976);
or U11264 (N_11264,N_6827,N_7860);
and U11265 (N_11265,N_6195,N_8987);
nor U11266 (N_11266,N_7055,N_8694);
nor U11267 (N_11267,N_8808,N_6086);
nand U11268 (N_11268,N_9732,N_7953);
nand U11269 (N_11269,N_9942,N_7874);
and U11270 (N_11270,N_9233,N_5314);
or U11271 (N_11271,N_6425,N_8867);
and U11272 (N_11272,N_6059,N_8303);
xor U11273 (N_11273,N_7446,N_9584);
xnor U11274 (N_11274,N_9679,N_7020);
xor U11275 (N_11275,N_6234,N_5178);
xor U11276 (N_11276,N_9788,N_5823);
xor U11277 (N_11277,N_6922,N_6117);
nand U11278 (N_11278,N_9633,N_5889);
and U11279 (N_11279,N_9687,N_6973);
nor U11280 (N_11280,N_8508,N_9908);
or U11281 (N_11281,N_6077,N_9119);
nand U11282 (N_11282,N_7570,N_5964);
nor U11283 (N_11283,N_8569,N_7460);
or U11284 (N_11284,N_7925,N_9112);
or U11285 (N_11285,N_7285,N_8625);
or U11286 (N_11286,N_7669,N_7517);
and U11287 (N_11287,N_6018,N_7596);
nor U11288 (N_11288,N_8029,N_9403);
xor U11289 (N_11289,N_5223,N_7764);
nor U11290 (N_11290,N_6775,N_7733);
nand U11291 (N_11291,N_9543,N_8424);
nand U11292 (N_11292,N_6194,N_8964);
and U11293 (N_11293,N_5956,N_7234);
nand U11294 (N_11294,N_8916,N_6596);
and U11295 (N_11295,N_9860,N_9549);
nor U11296 (N_11296,N_9724,N_6310);
and U11297 (N_11297,N_9082,N_9244);
or U11298 (N_11298,N_6839,N_7506);
and U11299 (N_11299,N_7458,N_5111);
xor U11300 (N_11300,N_9057,N_7376);
and U11301 (N_11301,N_7798,N_7309);
and U11302 (N_11302,N_5100,N_8507);
nand U11303 (N_11303,N_9867,N_6083);
and U11304 (N_11304,N_6643,N_9897);
nand U11305 (N_11305,N_7063,N_9161);
or U11306 (N_11306,N_5504,N_6699);
or U11307 (N_11307,N_6652,N_7406);
xnor U11308 (N_11308,N_5961,N_7850);
nand U11309 (N_11309,N_5372,N_7911);
and U11310 (N_11310,N_5162,N_8731);
nor U11311 (N_11311,N_5060,N_9407);
or U11312 (N_11312,N_7107,N_6236);
xnor U11313 (N_11313,N_5668,N_7671);
or U11314 (N_11314,N_7208,N_5072);
nand U11315 (N_11315,N_6476,N_7706);
and U11316 (N_11316,N_5307,N_8590);
and U11317 (N_11317,N_6647,N_8113);
xor U11318 (N_11318,N_7035,N_6550);
xor U11319 (N_11319,N_6286,N_5748);
nand U11320 (N_11320,N_9247,N_9080);
nor U11321 (N_11321,N_9958,N_6270);
nand U11322 (N_11322,N_7650,N_9940);
xor U11323 (N_11323,N_7908,N_6580);
nor U11324 (N_11324,N_9665,N_8287);
or U11325 (N_11325,N_7651,N_5432);
nand U11326 (N_11326,N_8380,N_7114);
nor U11327 (N_11327,N_8901,N_6737);
and U11328 (N_11328,N_5723,N_6008);
nand U11329 (N_11329,N_6762,N_6168);
nor U11330 (N_11330,N_9410,N_7447);
or U11331 (N_11331,N_8578,N_6208);
nand U11332 (N_11332,N_8930,N_8664);
or U11333 (N_11333,N_6179,N_7196);
or U11334 (N_11334,N_7525,N_5304);
and U11335 (N_11335,N_6029,N_7626);
nand U11336 (N_11336,N_6970,N_9847);
nor U11337 (N_11337,N_8266,N_5449);
nor U11338 (N_11338,N_8106,N_6260);
or U11339 (N_11339,N_6701,N_5098);
nand U11340 (N_11340,N_5419,N_8446);
nand U11341 (N_11341,N_6159,N_8413);
nor U11342 (N_11342,N_6284,N_9611);
or U11343 (N_11343,N_6118,N_6295);
nand U11344 (N_11344,N_5798,N_7796);
and U11345 (N_11345,N_5138,N_6502);
nand U11346 (N_11346,N_6776,N_5577);
nor U11347 (N_11347,N_6228,N_9952);
and U11348 (N_11348,N_7811,N_7040);
xor U11349 (N_11349,N_7272,N_6297);
or U11350 (N_11350,N_5988,N_9138);
nor U11351 (N_11351,N_8258,N_7784);
nand U11352 (N_11352,N_6443,N_8354);
and U11353 (N_11353,N_7381,N_9152);
nand U11354 (N_11354,N_9179,N_8143);
nor U11355 (N_11355,N_7421,N_9101);
nor U11356 (N_11356,N_8138,N_6100);
nor U11357 (N_11357,N_7660,N_6755);
xnor U11358 (N_11358,N_5815,N_5119);
nor U11359 (N_11359,N_7975,N_9148);
nand U11360 (N_11360,N_6094,N_9103);
nand U11361 (N_11361,N_8541,N_9634);
xor U11362 (N_11362,N_6275,N_7943);
nand U11363 (N_11363,N_9419,N_7569);
nor U11364 (N_11364,N_8629,N_9888);
or U11365 (N_11365,N_6760,N_7159);
nor U11366 (N_11366,N_7976,N_7885);
and U11367 (N_11367,N_5362,N_8071);
nor U11368 (N_11368,N_6226,N_5584);
nand U11369 (N_11369,N_7439,N_9134);
and U11370 (N_11370,N_8482,N_6904);
and U11371 (N_11371,N_8393,N_7122);
xor U11372 (N_11372,N_5349,N_9109);
or U11373 (N_11373,N_7528,N_7177);
nor U11374 (N_11374,N_5864,N_7829);
or U11375 (N_11375,N_6039,N_5929);
nor U11376 (N_11376,N_9218,N_6817);
or U11377 (N_11377,N_6430,N_6678);
or U11378 (N_11378,N_8884,N_5141);
and U11379 (N_11379,N_8659,N_6046);
nand U11380 (N_11380,N_8621,N_8042);
or U11381 (N_11381,N_8465,N_7732);
nand U11382 (N_11382,N_7028,N_8168);
nor U11383 (N_11383,N_7965,N_5827);
or U11384 (N_11384,N_8776,N_5326);
nor U11385 (N_11385,N_5562,N_8552);
nand U11386 (N_11386,N_7470,N_8175);
xor U11387 (N_11387,N_5299,N_5691);
nor U11388 (N_11388,N_6184,N_9553);
nor U11389 (N_11389,N_5914,N_5389);
or U11390 (N_11390,N_9697,N_9846);
xnor U11391 (N_11391,N_6853,N_5353);
nand U11392 (N_11392,N_9269,N_6620);
nor U11393 (N_11393,N_8065,N_5356);
xnor U11394 (N_11394,N_7002,N_6322);
xnor U11395 (N_11395,N_9363,N_5844);
nand U11396 (N_11396,N_9854,N_9049);
and U11397 (N_11397,N_9314,N_8058);
and U11398 (N_11398,N_8296,N_9168);
nor U11399 (N_11399,N_6586,N_8490);
nand U11400 (N_11400,N_9673,N_7598);
or U11401 (N_11401,N_8102,N_8273);
nor U11402 (N_11402,N_8775,N_7050);
and U11403 (N_11403,N_5990,N_9275);
nand U11404 (N_11404,N_5623,N_8083);
or U11405 (N_11405,N_9669,N_7430);
nand U11406 (N_11406,N_6982,N_8732);
nand U11407 (N_11407,N_8037,N_8226);
xor U11408 (N_11408,N_6752,N_6569);
nor U11409 (N_11409,N_5776,N_8026);
nor U11410 (N_11410,N_8600,N_9208);
or U11411 (N_11411,N_6096,N_8688);
nand U11412 (N_11412,N_6598,N_6383);
xor U11413 (N_11413,N_8152,N_5944);
and U11414 (N_11414,N_7231,N_5234);
nor U11415 (N_11415,N_5873,N_6545);
or U11416 (N_11416,N_7191,N_5262);
or U11417 (N_11417,N_5458,N_9412);
and U11418 (N_11418,N_6429,N_8678);
nor U11419 (N_11419,N_7070,N_6111);
xor U11420 (N_11420,N_5172,N_6779);
or U11421 (N_11421,N_9876,N_7198);
and U11422 (N_11422,N_5144,N_5682);
and U11423 (N_11423,N_5706,N_8844);
or U11424 (N_11424,N_5189,N_9457);
xor U11425 (N_11425,N_5260,N_5871);
xor U11426 (N_11426,N_6456,N_7958);
nor U11427 (N_11427,N_6183,N_8665);
xnor U11428 (N_11428,N_5137,N_7639);
xnor U11429 (N_11429,N_7871,N_7462);
nand U11430 (N_11430,N_9400,N_9073);
or U11431 (N_11431,N_9295,N_6332);
xnor U11432 (N_11432,N_9182,N_9578);
and U11433 (N_11433,N_6423,N_9490);
nor U11434 (N_11434,N_5597,N_8555);
and U11435 (N_11435,N_8476,N_6287);
or U11436 (N_11436,N_5450,N_9626);
and U11437 (N_11437,N_8118,N_6640);
nand U11438 (N_11438,N_9918,N_8418);
nand U11439 (N_11439,N_8615,N_5305);
xnor U11440 (N_11440,N_8963,N_8297);
and U11441 (N_11441,N_8634,N_7803);
nand U11442 (N_11442,N_9749,N_8992);
nor U11443 (N_11443,N_7341,N_8200);
nor U11444 (N_11444,N_5589,N_9910);
nor U11445 (N_11445,N_7588,N_7830);
or U11446 (N_11446,N_5734,N_9576);
and U11447 (N_11447,N_7767,N_9703);
xnor U11448 (N_11448,N_8722,N_6135);
and U11449 (N_11449,N_5957,N_9485);
and U11450 (N_11450,N_5641,N_9922);
xnor U11451 (N_11451,N_7296,N_5896);
nand U11452 (N_11452,N_7431,N_7190);
xor U11453 (N_11453,N_9345,N_7053);
nor U11454 (N_11454,N_9727,N_8591);
or U11455 (N_11455,N_7535,N_9480);
xnor U11456 (N_11456,N_6266,N_7780);
xor U11457 (N_11457,N_7189,N_9829);
nand U11458 (N_11458,N_8270,N_7512);
and U11459 (N_11459,N_7959,N_6609);
nor U11460 (N_11460,N_6166,N_7617);
nor U11461 (N_11461,N_5268,N_8275);
nor U11462 (N_11462,N_5416,N_8518);
and U11463 (N_11463,N_7640,N_8550);
or U11464 (N_11464,N_9261,N_8498);
xnor U11465 (N_11465,N_6572,N_5772);
xnor U11466 (N_11466,N_7483,N_7037);
and U11467 (N_11467,N_8360,N_6078);
and U11468 (N_11468,N_5573,N_9796);
xnor U11469 (N_11469,N_8713,N_8761);
or U11470 (N_11470,N_7369,N_5824);
or U11471 (N_11471,N_9467,N_7672);
or U11472 (N_11472,N_7550,N_7557);
and U11473 (N_11473,N_5384,N_8495);
nor U11474 (N_11474,N_6215,N_8402);
xnor U11475 (N_11475,N_5669,N_5666);
xnor U11476 (N_11476,N_8022,N_7653);
nand U11477 (N_11477,N_8540,N_8692);
or U11478 (N_11478,N_6978,N_9527);
or U11479 (N_11479,N_9002,N_9055);
or U11480 (N_11480,N_7711,N_9445);
nor U11481 (N_11481,N_7357,N_7252);
xnor U11482 (N_11482,N_8943,N_8838);
nor U11483 (N_11483,N_6200,N_6092);
nand U11484 (N_11484,N_9834,N_7214);
and U11485 (N_11485,N_7150,N_8948);
nand U11486 (N_11486,N_5497,N_9456);
nor U11487 (N_11487,N_9133,N_9312);
or U11488 (N_11488,N_8045,N_6467);
xor U11489 (N_11489,N_9162,N_6131);
or U11490 (N_11490,N_5872,N_9793);
nor U11491 (N_11491,N_6002,N_6389);
nand U11492 (N_11492,N_9815,N_5631);
nand U11493 (N_11493,N_7723,N_7021);
and U11494 (N_11494,N_7102,N_8197);
nand U11495 (N_11495,N_7758,N_6384);
xor U11496 (N_11496,N_9620,N_6150);
and U11497 (N_11497,N_9043,N_9139);
xor U11498 (N_11498,N_5375,N_8701);
xor U11499 (N_11499,N_6749,N_6796);
nor U11500 (N_11500,N_6914,N_9804);
and U11501 (N_11501,N_6849,N_6951);
or U11502 (N_11502,N_5984,N_5722);
or U11503 (N_11503,N_9937,N_7842);
nor U11504 (N_11504,N_8072,N_5472);
nor U11505 (N_11505,N_7435,N_5892);
or U11506 (N_11506,N_8472,N_5747);
nand U11507 (N_11507,N_9169,N_6336);
and U11508 (N_11508,N_6109,N_5039);
and U11509 (N_11509,N_7000,N_5891);
and U11510 (N_11510,N_9525,N_8820);
nor U11511 (N_11511,N_6073,N_5194);
or U11512 (N_11512,N_5637,N_6730);
nor U11513 (N_11513,N_5520,N_8649);
nand U11514 (N_11514,N_5989,N_9120);
nand U11515 (N_11515,N_6707,N_9187);
xnor U11516 (N_11516,N_9263,N_5317);
or U11517 (N_11517,N_6906,N_6097);
nor U11518 (N_11518,N_8893,N_8087);
nor U11519 (N_11519,N_9339,N_6023);
or U11520 (N_11520,N_8111,N_8348);
and U11521 (N_11521,N_6816,N_5740);
and U11522 (N_11522,N_5903,N_8116);
or U11523 (N_11523,N_8900,N_9721);
nand U11524 (N_11524,N_8063,N_6318);
xor U11525 (N_11525,N_7116,N_9704);
nor U11526 (N_11526,N_9666,N_5548);
xnor U11527 (N_11527,N_7481,N_9033);
or U11528 (N_11528,N_9117,N_7222);
or U11529 (N_11529,N_6633,N_6589);
and U11530 (N_11530,N_5735,N_6891);
xor U11531 (N_11531,N_7905,N_8725);
or U11532 (N_11532,N_6845,N_5563);
xnor U11533 (N_11533,N_7849,N_6400);
nor U11534 (N_11534,N_9874,N_7132);
nor U11535 (N_11535,N_9337,N_5303);
nand U11536 (N_11536,N_5366,N_8923);
xnor U11537 (N_11537,N_7684,N_5538);
nand U11538 (N_11538,N_7670,N_7587);
and U11539 (N_11539,N_7675,N_9346);
xor U11540 (N_11540,N_5834,N_6517);
nor U11541 (N_11541,N_5916,N_6626);
nand U11542 (N_11542,N_7844,N_5134);
and U11543 (N_11543,N_8316,N_6458);
nand U11544 (N_11544,N_9797,N_6878);
or U11545 (N_11545,N_7689,N_8387);
nand U11546 (N_11546,N_5012,N_8162);
or U11547 (N_11547,N_6028,N_7705);
xor U11548 (N_11548,N_6198,N_7396);
nor U11549 (N_11549,N_5661,N_7727);
and U11550 (N_11550,N_8371,N_7624);
or U11551 (N_11551,N_8438,N_6672);
nor U11552 (N_11552,N_5983,N_6534);
or U11553 (N_11553,N_7658,N_5296);
and U11554 (N_11554,N_5705,N_8913);
nor U11555 (N_11555,N_6149,N_5436);
nor U11556 (N_11556,N_5907,N_7047);
and U11557 (N_11557,N_7921,N_5558);
and U11558 (N_11558,N_7866,N_7044);
nand U11559 (N_11559,N_6265,N_5998);
xor U11560 (N_11560,N_6663,N_9795);
or U11561 (N_11561,N_7334,N_9712);
and U11562 (N_11562,N_5105,N_7771);
or U11563 (N_11563,N_8291,N_5561);
nor U11564 (N_11564,N_7601,N_9277);
xnor U11565 (N_11565,N_7822,N_5731);
xor U11566 (N_11566,N_6300,N_5129);
and U11567 (N_11567,N_5868,N_5604);
nor U11568 (N_11568,N_7621,N_5743);
or U11569 (N_11569,N_5321,N_7253);
nand U11570 (N_11570,N_8181,N_5900);
or U11571 (N_11571,N_5645,N_9722);
nor U11572 (N_11572,N_9228,N_7401);
nor U11573 (N_11573,N_6560,N_9856);
nand U11574 (N_11574,N_8409,N_8897);
nand U11575 (N_11575,N_6848,N_7373);
nor U11576 (N_11576,N_9632,N_6928);
nand U11577 (N_11577,N_6247,N_5404);
and U11578 (N_11578,N_5590,N_8305);
and U11579 (N_11579,N_9132,N_5951);
xnor U11580 (N_11580,N_5536,N_5969);
xor U11581 (N_11581,N_9019,N_8949);
and U11582 (N_11582,N_8630,N_5113);
nand U11583 (N_11583,N_8171,N_5835);
xor U11584 (N_11584,N_5165,N_9379);
nor U11585 (N_11585,N_9736,N_7120);
nand U11586 (N_11586,N_9360,N_7315);
or U11587 (N_11587,N_6905,N_7255);
nor U11588 (N_11588,N_7526,N_7263);
and U11589 (N_11589,N_9301,N_9350);
or U11590 (N_11590,N_6996,N_7594);
nand U11591 (N_11591,N_8547,N_7910);
and U11592 (N_11592,N_6174,N_6527);
nand U11593 (N_11593,N_9681,N_9565);
and U11594 (N_11594,N_6972,N_5622);
nand U11595 (N_11595,N_9442,N_9056);
and U11596 (N_11596,N_9877,N_9988);
xor U11597 (N_11597,N_7981,N_9344);
and U11598 (N_11598,N_8073,N_9827);
xor U11599 (N_11599,N_5225,N_8300);
and U11600 (N_11600,N_7699,N_8584);
nor U11601 (N_11601,N_6189,N_8564);
or U11602 (N_11602,N_5252,N_9850);
and U11603 (N_11603,N_5833,N_8921);
nor U11604 (N_11604,N_8833,N_8074);
nor U11605 (N_11605,N_5231,N_6187);
and U11606 (N_11606,N_8060,N_8607);
or U11607 (N_11607,N_5676,N_9828);
and U11608 (N_11608,N_7405,N_5831);
xor U11609 (N_11609,N_7668,N_6367);
nor U11610 (N_11610,N_8224,N_5576);
xnor U11611 (N_11611,N_7466,N_6488);
xor U11612 (N_11612,N_9567,N_8173);
xor U11613 (N_11613,N_8109,N_7916);
nand U11614 (N_11614,N_8618,N_9647);
or U11615 (N_11615,N_9151,N_6113);
or U11616 (N_11616,N_8330,N_6716);
or U11617 (N_11617,N_6697,N_5875);
and U11618 (N_11618,N_7062,N_6850);
nand U11619 (N_11619,N_9383,N_7607);
nor U11620 (N_11620,N_7343,N_9491);
nand U11621 (N_11621,N_9617,N_6064);
nor U11622 (N_11622,N_8234,N_7186);
xor U11623 (N_11623,N_8572,N_9973);
xor U11624 (N_11624,N_5337,N_5591);
and U11625 (N_11625,N_6562,N_9366);
or U11626 (N_11626,N_6597,N_5044);
nor U11627 (N_11627,N_6500,N_7548);
and U11628 (N_11628,N_8673,N_6279);
and U11629 (N_11629,N_8588,N_6144);
and U11630 (N_11630,N_7777,N_9950);
nand U11631 (N_11631,N_9585,N_7731);
or U11632 (N_11632,N_9547,N_7824);
nand U11633 (N_11633,N_6233,N_9009);
nand U11634 (N_11634,N_9226,N_9901);
xor U11635 (N_11635,N_9826,N_6766);
xor U11636 (N_11636,N_6689,N_7868);
or U11637 (N_11637,N_8885,N_7179);
or U11638 (N_11638,N_5115,N_9476);
xnor U11639 (N_11639,N_6192,N_5055);
and U11640 (N_11640,N_6585,N_5075);
xnor U11641 (N_11641,N_7378,N_6099);
and U11642 (N_11642,N_6510,N_7354);
xor U11643 (N_11643,N_7065,N_5658);
or U11644 (N_11644,N_5169,N_8993);
or U11645 (N_11645,N_6675,N_6329);
nor U11646 (N_11646,N_6171,N_9580);
nor U11647 (N_11647,N_6182,N_9322);
nand U11648 (N_11648,N_9121,N_8727);
or U11649 (N_11649,N_5549,N_6529);
and U11650 (N_11650,N_8740,N_6966);
xnor U11651 (N_11651,N_7956,N_7433);
xnor U11652 (N_11652,N_7997,N_7509);
or U11653 (N_11653,N_5310,N_9349);
xor U11654 (N_11654,N_7162,N_7807);
xor U11655 (N_11655,N_6334,N_8822);
and U11656 (N_11656,N_8458,N_8247);
nand U11657 (N_11657,N_8400,N_9770);
xor U11658 (N_11658,N_9640,N_7362);
xnor U11659 (N_11659,N_8982,N_9342);
nor U11660 (N_11660,N_5968,N_7323);
xnor U11661 (N_11661,N_6146,N_7904);
nand U11662 (N_11662,N_5114,N_7121);
and U11663 (N_11663,N_6581,N_9358);
or U11664 (N_11664,N_5557,N_9282);
and U11665 (N_11665,N_5158,N_8931);
xnor U11666 (N_11666,N_7019,N_7238);
xnor U11667 (N_11667,N_5546,N_5931);
nand U11668 (N_11668,N_9996,N_6025);
nor U11669 (N_11669,N_6627,N_6991);
and U11670 (N_11670,N_9254,N_6222);
or U11671 (N_11671,N_7029,N_5924);
nor U11672 (N_11672,N_5498,N_8340);
nand U11673 (N_11673,N_8668,N_8608);
nand U11674 (N_11674,N_8310,N_5517);
and U11675 (N_11675,N_8779,N_5446);
or U11676 (N_11676,N_5182,N_9579);
xor U11677 (N_11677,N_6361,N_9917);
and U11678 (N_11678,N_8589,N_6852);
or U11679 (N_11679,N_7094,N_8785);
nand U11680 (N_11680,N_9443,N_6540);
xnor U11681 (N_11681,N_5161,N_5481);
nand U11682 (N_11682,N_9422,N_6160);
xnor U11683 (N_11683,N_5649,N_5717);
xnor U11684 (N_11684,N_5242,N_8586);
xnor U11685 (N_11685,N_5521,N_8039);
nand U11686 (N_11686,N_8233,N_5886);
xnor U11687 (N_11687,N_6491,N_7765);
nor U11688 (N_11688,N_5975,N_7350);
nand U11689 (N_11689,N_6564,N_5816);
nand U11690 (N_11690,N_9059,N_7450);
or U11691 (N_11691,N_5116,N_9607);
nand U11692 (N_11692,N_6292,N_7618);
nand U11693 (N_11693,N_6320,N_5508);
or U11694 (N_11694,N_8000,N_6698);
nor U11695 (N_11695,N_6012,N_8596);
nand U11696 (N_11696,N_9862,N_6518);
and U11697 (N_11697,N_6761,N_6422);
nor U11698 (N_11698,N_5783,N_5279);
and U11699 (N_11699,N_5617,N_7938);
and U11700 (N_11700,N_9656,N_8747);
or U11701 (N_11701,N_7761,N_8915);
and U11702 (N_11702,N_9998,N_5082);
xor U11703 (N_11703,N_9515,N_7752);
nand U11704 (N_11704,N_7493,N_9497);
and U11705 (N_11705,N_9070,N_9964);
xnor U11706 (N_11706,N_8290,N_7408);
nor U11707 (N_11707,N_9742,N_7577);
xnor U11708 (N_11708,N_5051,N_9831);
xor U11709 (N_11709,N_6180,N_7001);
xor U11710 (N_11710,N_6939,N_9745);
nand U11711 (N_11711,N_5329,N_8307);
and U11712 (N_11712,N_6634,N_5340);
and U11713 (N_11713,N_9726,N_5348);
or U11714 (N_11714,N_7291,N_8013);
or U11715 (N_11715,N_7813,N_5204);
xor U11716 (N_11716,N_9786,N_5828);
nand U11717 (N_11717,N_6127,N_8012);
nor U11718 (N_11718,N_8601,N_9569);
xor U11719 (N_11719,N_6851,N_6101);
nand U11720 (N_11720,N_9662,N_9223);
nor U11721 (N_11721,N_6313,N_8502);
xor U11722 (N_11722,N_6712,N_8163);
nor U11723 (N_11723,N_8876,N_7312);
or U11724 (N_11724,N_9521,N_9035);
xor U11725 (N_11725,N_7197,N_9309);
nor U11726 (N_11726,N_6139,N_6434);
nor U11727 (N_11727,N_9516,N_6847);
or U11728 (N_11728,N_8281,N_6881);
nor U11729 (N_11729,N_8748,N_7934);
nor U11730 (N_11730,N_9812,N_5089);
nand U11731 (N_11731,N_5870,N_9945);
xor U11732 (N_11732,N_5088,N_5350);
or U11733 (N_11733,N_8202,N_5258);
or U11734 (N_11734,N_7147,N_9174);
and U11735 (N_11735,N_7402,N_9671);
xnor U11736 (N_11736,N_7978,N_8277);
nand U11737 (N_11737,N_8186,N_6235);
nand U11738 (N_11738,N_8525,N_6565);
nand U11739 (N_11739,N_8532,N_6826);
nand U11740 (N_11740,N_7620,N_6858);
nand U11741 (N_11741,N_6612,N_8840);
xor U11742 (N_11742,N_8230,N_6264);
xnor U11743 (N_11743,N_9493,N_7308);
nor U11744 (N_11744,N_9124,N_5769);
and U11745 (N_11745,N_9306,N_7042);
or U11746 (N_11746,N_9976,N_8683);
or U11747 (N_11747,N_5693,N_5733);
nand U11748 (N_11748,N_7137,N_8080);
or U11749 (N_11749,N_9163,N_6764);
nor U11750 (N_11750,N_8434,N_5210);
nor U11751 (N_11751,N_9230,N_5409);
xnor U11752 (N_11752,N_5583,N_5191);
nor U11753 (N_11753,N_5344,N_9370);
and U11754 (N_11754,N_6823,N_5992);
or U11755 (N_11755,N_9470,N_7753);
and U11756 (N_11756,N_7873,N_7572);
nor U11757 (N_11757,N_7297,N_6319);
and U11758 (N_11758,N_7688,N_5568);
and U11759 (N_11759,N_8439,N_6638);
xnor U11760 (N_11760,N_7792,N_7303);
or U11761 (N_11761,N_7288,N_8519);
nor U11762 (N_11762,N_7687,N_5587);
nor U11763 (N_11763,N_5198,N_8726);
xor U11764 (N_11764,N_7487,N_8581);
or U11765 (N_11765,N_9635,N_6414);
and U11766 (N_11766,N_9663,N_6671);
xor U11767 (N_11767,N_5246,N_5595);
nand U11768 (N_11768,N_8928,N_8334);
and U11769 (N_11769,N_6485,N_5185);
xor U11770 (N_11770,N_9348,N_8521);
xnor U11771 (N_11771,N_5856,N_9332);
nand U11772 (N_11772,N_9791,N_8240);
xor U11773 (N_11773,N_7720,N_5413);
nand U11774 (N_11774,N_5545,N_7890);
xor U11775 (N_11775,N_7887,N_5030);
or U11776 (N_11776,N_6916,N_7931);
nand U11777 (N_11777,N_8984,N_9833);
and U11778 (N_11778,N_8331,N_8622);
nor U11779 (N_11779,N_6390,N_6912);
xor U11780 (N_11780,N_5640,N_8131);
and U11781 (N_11781,N_8904,N_6571);
or U11782 (N_11782,N_8262,N_8272);
nand U11783 (N_11783,N_9857,N_6022);
or U11784 (N_11784,N_6549,N_5887);
nor U11785 (N_11785,N_9916,N_7183);
nand U11786 (N_11786,N_8514,N_7427);
nor U11787 (N_11787,N_5716,N_6692);
or U11788 (N_11788,N_9114,N_6750);
xor U11789 (N_11789,N_5192,N_8792);
or U11790 (N_11790,N_7305,N_9489);
and U11791 (N_11791,N_5430,N_9011);
nand U11792 (N_11792,N_5135,N_8877);
or U11793 (N_11793,N_9836,N_5648);
nor U11794 (N_11794,N_7772,N_8099);
or U11795 (N_11795,N_5959,N_5671);
or U11796 (N_11796,N_8117,N_7648);
and U11797 (N_11797,N_7613,N_9830);
and U11798 (N_11798,N_5405,N_5578);
nor U11799 (N_11799,N_6089,N_7115);
nand U11800 (N_11800,N_6810,N_7316);
or U11801 (N_11801,N_5950,N_6296);
nor U11802 (N_11802,N_8255,N_5971);
and U11803 (N_11803,N_7098,N_9787);
xnor U11804 (N_11804,N_9484,N_7193);
nor U11805 (N_11805,N_5110,N_5494);
and U11806 (N_11806,N_8733,N_8372);
nor U11807 (N_11807,N_8425,N_8250);
nor U11808 (N_11808,N_9433,N_7565);
nand U11809 (N_11809,N_8320,N_7856);
nor U11810 (N_11810,N_6173,N_5490);
nor U11811 (N_11811,N_7066,N_7739);
xnor U11812 (N_11812,N_7801,N_9238);
xor U11813 (N_11813,N_6998,N_8804);
nand U11814 (N_11814,N_7898,N_7043);
nand U11815 (N_11815,N_5974,N_5149);
nor U11816 (N_11816,N_9414,N_9376);
or U11817 (N_11817,N_6321,N_9299);
nor U11818 (N_11818,N_8477,N_7912);
nor U11819 (N_11819,N_7826,N_6874);
xnor U11820 (N_11820,N_5714,N_9194);
nand U11821 (N_11821,N_9898,N_6984);
xnor U11822 (N_11822,N_8504,N_9384);
nand U11823 (N_11823,N_5226,N_6696);
or U11824 (N_11824,N_6288,N_9157);
nand U11825 (N_11825,N_5993,N_9839);
and U11826 (N_11826,N_5293,N_6250);
and U11827 (N_11827,N_7877,N_9657);
nand U11828 (N_11828,N_6543,N_7519);
xnor U11829 (N_11829,N_7142,N_5665);
xor U11830 (N_11830,N_7583,N_8850);
xor U11831 (N_11831,N_6309,N_9058);
or U11832 (N_11832,N_5010,N_9931);
and U11833 (N_11833,N_8376,N_7111);
nand U11834 (N_11834,N_8889,N_8461);
or U11835 (N_11835,N_9097,N_7967);
or U11836 (N_11836,N_5026,N_5156);
nand U11837 (N_11837,N_9245,N_5224);
xnor U11838 (N_11838,N_5503,N_9046);
nor U11839 (N_11839,N_8529,N_7268);
or U11840 (N_11840,N_9302,N_5672);
and U11841 (N_11841,N_7103,N_5867);
nand U11842 (N_11842,N_6873,N_6088);
xor U11843 (N_11843,N_9000,N_6259);
nor U11844 (N_11844,N_8766,N_5097);
nor U11845 (N_11845,N_5324,N_7069);
nor U11846 (N_11846,N_5276,N_7755);
or U11847 (N_11847,N_7346,N_5688);
nand U11848 (N_11848,N_8412,N_8526);
xnor U11849 (N_11849,N_5395,N_9368);
or U11850 (N_11850,N_7232,N_7741);
nand U11851 (N_11851,N_8751,N_9573);
or U11852 (N_11852,N_5173,N_5238);
or U11853 (N_11853,N_9398,N_8048);
and U11854 (N_11854,N_7717,N_7281);
or U11855 (N_11855,N_5986,N_8851);
nor U11856 (N_11856,N_5724,N_6768);
nor U11857 (N_11857,N_9885,N_9646);
nand U11858 (N_11858,N_9195,N_6520);
and U11859 (N_11859,N_8236,N_9266);
nand U11860 (N_11860,N_7735,N_7928);
nand U11861 (N_11861,N_7864,N_6777);
nor U11862 (N_11862,N_5371,N_6887);
nor U11863 (N_11863,N_8475,N_9875);
and U11864 (N_11864,N_7999,N_5859);
xor U11865 (N_11865,N_9394,N_8480);
and U11866 (N_11866,N_8914,N_7809);
xnor U11867 (N_11867,N_9741,N_9343);
and U11868 (N_11868,N_5839,N_6040);
or U11869 (N_11869,N_6903,N_7008);
xnor U11870 (N_11870,N_6371,N_5219);
xor U11871 (N_11871,N_5813,N_8153);
xor U11872 (N_11872,N_5426,N_9423);
or U11873 (N_11873,N_6402,N_6659);
xnor U11874 (N_11874,N_9813,N_5374);
and U11875 (N_11875,N_8709,N_7425);
xnor U11876 (N_11876,N_6431,N_5715);
nand U11877 (N_11877,N_8341,N_8868);
or U11878 (N_11878,N_8460,N_8953);
xor U11879 (N_11879,N_9953,N_8979);
nand U11880 (N_11880,N_8432,N_7117);
or U11881 (N_11881,N_6960,N_8410);
and U11882 (N_11882,N_8431,N_6224);
or U11883 (N_11883,N_9944,N_6600);
or U11884 (N_11884,N_9537,N_7223);
or U11885 (N_11885,N_9811,N_5146);
xor U11886 (N_11886,N_6931,N_8848);
xor U11887 (N_11887,N_5308,N_8499);
or U11888 (N_11888,N_8593,N_8839);
or U11889 (N_11889,N_5751,N_6713);
or U11890 (N_11890,N_6084,N_8002);
xor U11891 (N_11891,N_5477,N_5383);
xnor U11892 (N_11892,N_6917,N_6276);
xor U11893 (N_11893,N_6666,N_9222);
nor U11894 (N_11894,N_6441,N_7951);
and U11895 (N_11895,N_9824,N_5463);
xor U11896 (N_11896,N_8627,N_8274);
nand U11897 (N_11897,N_7411,N_6554);
xor U11898 (N_11898,N_7757,N_6570);
and U11899 (N_11899,N_9779,N_7124);
nor U11900 (N_11900,N_5768,N_7241);
and U11901 (N_11901,N_7112,N_7239);
nand U11902 (N_11902,N_7052,N_6872);
or U11903 (N_11903,N_7608,N_9289);
nand U11904 (N_11904,N_6360,N_8674);
or U11905 (N_11905,N_5539,N_7984);
xor U11906 (N_11906,N_6573,N_9568);
nor U11907 (N_11907,N_8920,N_5209);
xor U11908 (N_11908,N_7207,N_7673);
and U11909 (N_11909,N_9719,N_6637);
nand U11910 (N_11910,N_5370,N_8869);
and U11911 (N_11911,N_6381,N_6257);
nand U11912 (N_11912,N_7173,N_7730);
and U11913 (N_11913,N_9361,N_5217);
nor U11914 (N_11914,N_7318,N_5123);
nor U11915 (N_11915,N_8278,N_6307);
nor U11916 (N_11916,N_5789,N_9240);
nand U11917 (N_11917,N_9689,N_6480);
or U11918 (N_11918,N_5403,N_9939);
and U11919 (N_11919,N_6893,N_7941);
nor U11920 (N_11920,N_6514,N_9597);
nand U11921 (N_11921,N_6795,N_6820);
xnor U11922 (N_11922,N_8606,N_7718);
and U11923 (N_11923,N_7211,N_8092);
xnor U11924 (N_11924,N_5522,N_6861);
nand U11925 (N_11925,N_7919,N_8496);
nand U11926 (N_11926,N_7086,N_6214);
nor U11927 (N_11927,N_6068,N_9878);
xnor U11928 (N_11928,N_5084,N_9140);
or U11929 (N_11929,N_6721,N_7553);
or U11930 (N_11930,N_6410,N_8147);
or U11931 (N_11931,N_8411,N_9466);
or U11932 (N_11932,N_8213,N_8398);
nor U11933 (N_11933,N_5016,N_7012);
nor U11934 (N_11934,N_8177,N_6154);
nor U11935 (N_11935,N_5083,N_8639);
and U11936 (N_11936,N_5122,N_9645);
or U11937 (N_11937,N_6877,N_5810);
nor U11938 (N_11938,N_5544,N_5154);
nand U11939 (N_11939,N_6553,N_7857);
and U11940 (N_11940,N_9071,N_5176);
xor U11941 (N_11941,N_5553,N_9127);
and U11942 (N_11942,N_5764,N_5678);
nor U11943 (N_11943,N_9655,N_5526);
nor U11944 (N_11944,N_5269,N_7219);
nand U11945 (N_11945,N_8319,N_9517);
nor U11946 (N_11946,N_5860,N_5120);
nor U11947 (N_11947,N_7972,N_5106);
or U11948 (N_11948,N_5093,N_5777);
or U11949 (N_11949,N_6162,N_7986);
or U11950 (N_11950,N_6897,N_5708);
and U11951 (N_11951,N_8493,N_6075);
or U11952 (N_11952,N_5863,N_9478);
xor U11953 (N_11953,N_9773,N_6669);
nor U11954 (N_11954,N_6567,N_9533);
nand U11955 (N_11955,N_8537,N_6936);
nor U11956 (N_11956,N_7521,N_6155);
nor U11957 (N_11957,N_5955,N_7202);
xor U11958 (N_11958,N_9108,N_6587);
nor U11959 (N_11959,N_9587,N_7983);
or U11960 (N_11960,N_5700,N_8648);
nor U11961 (N_11961,N_6983,N_9242);
and U11962 (N_11962,N_7453,N_7486);
nor U11963 (N_11963,N_9868,N_5214);
nand U11964 (N_11964,N_7881,N_7902);
xor U11965 (N_11965,N_6773,N_9938);
and U11966 (N_11966,N_7823,N_8437);
or U11967 (N_11967,N_6830,N_9572);
nor U11968 (N_11968,N_5193,N_5905);
nor U11969 (N_11969,N_6439,N_6374);
and U11970 (N_11970,N_9606,N_9381);
nand U11971 (N_11971,N_6312,N_6175);
nand U11972 (N_11972,N_7923,N_5915);
xnor U11973 (N_11973,N_5675,N_9956);
xor U11974 (N_11974,N_5880,N_6990);
xnor U11975 (N_11975,N_8337,N_5787);
xnor U11976 (N_11976,N_6552,N_8292);
or U11977 (N_11977,N_6790,N_7476);
nand U11978 (N_11978,N_7894,N_8185);
nor U11979 (N_11979,N_8157,N_7099);
xor U11980 (N_11980,N_5580,N_9329);
or U11981 (N_11981,N_6223,N_8729);
nand U11982 (N_11982,N_9173,N_9211);
nor U11983 (N_11983,N_8932,N_9705);
or U11984 (N_11984,N_7793,N_9912);
or U11985 (N_11985,N_6686,N_5599);
xor U11986 (N_11986,N_5025,N_7586);
nand U11987 (N_11987,N_6658,N_6635);
and U11988 (N_11988,N_7474,N_7171);
nor U11989 (N_11989,N_6351,N_7737);
nor U11990 (N_11990,N_9686,N_8961);
nor U11991 (N_11991,N_6499,N_8463);
nor U11992 (N_11992,N_5022,N_6468);
or U11993 (N_11993,N_5600,N_7095);
xor U11994 (N_11994,N_8216,N_6347);
xnor U11995 (N_11995,N_9323,N_9921);
and U11996 (N_11996,N_5575,N_8035);
and U11997 (N_11997,N_8298,N_5981);
and U11998 (N_11998,N_7331,N_7276);
nand U11999 (N_11999,N_8637,N_7901);
or U12000 (N_12000,N_7610,N_5874);
nand U12001 (N_12001,N_6720,N_8453);
and U12002 (N_12002,N_8105,N_5174);
and U12003 (N_12003,N_5507,N_6802);
nand U12004 (N_12004,N_5890,N_6822);
and U12005 (N_12005,N_6230,N_6533);
nand U12006 (N_12006,N_6119,N_6196);
or U12007 (N_12007,N_6501,N_6733);
or U12008 (N_12008,N_7442,N_7508);
nor U12009 (N_12009,N_5511,N_7073);
xor U12010 (N_12010,N_7883,N_9899);
or U12011 (N_12011,N_6803,N_7740);
nor U12012 (N_12012,N_8528,N_8158);
nor U12013 (N_12013,N_5318,N_6961);
nor U12014 (N_12014,N_9738,N_8284);
nand U12015 (N_12015,N_5699,N_9561);
xor U12016 (N_12016,N_6965,N_8190);
nand U12017 (N_12017,N_8700,N_5206);
and U12018 (N_12018,N_6201,N_9562);
and U12019 (N_12019,N_5474,N_9911);
or U12020 (N_12020,N_6193,N_9421);
xnor U12021 (N_12021,N_7817,N_5248);
nand U12022 (N_12022,N_6512,N_7358);
xor U12023 (N_12023,N_9474,N_7563);
or U12024 (N_12024,N_8535,N_9564);
xnor U12025 (N_12025,N_6070,N_8793);
xor U12026 (N_12026,N_6137,N_9227);
nor U12027 (N_12027,N_6621,N_8699);
and U12028 (N_12028,N_6921,N_9481);
nor U12029 (N_12029,N_9759,N_6108);
nand U12030 (N_12030,N_6157,N_5410);
and U12031 (N_12031,N_6132,N_7110);
nand U12032 (N_12032,N_5031,N_6651);
and U12033 (N_12033,N_9110,N_6062);
nand U12034 (N_12034,N_5411,N_8658);
nand U12035 (N_12035,N_8856,N_6915);
and U12036 (N_12036,N_7372,N_7970);
and U12037 (N_12037,N_8220,N_6042);
nor U12038 (N_12038,N_6446,N_7944);
xnor U12039 (N_12039,N_6356,N_5876);
nand U12040 (N_12040,N_9552,N_7041);
nor U12041 (N_12041,N_7926,N_6575);
xnor U12042 (N_12042,N_8456,N_6369);
nand U12043 (N_12043,N_7364,N_8924);
and U12044 (N_12044,N_9746,N_6748);
or U12045 (N_12045,N_7676,N_6178);
and U12046 (N_12046,N_6152,N_8599);
and U12047 (N_12047,N_8282,N_6004);
nor U12048 (N_12048,N_8194,N_7160);
and U12049 (N_12049,N_9270,N_6785);
or U12050 (N_12050,N_8231,N_8672);
nand U12051 (N_12051,N_6017,N_6952);
nand U12052 (N_12052,N_7295,N_9472);
nor U12053 (N_12053,N_8166,N_9171);
and U12054 (N_12054,N_5749,N_7441);
nand U12055 (N_12055,N_9785,N_8784);
xor U12056 (N_12056,N_8854,N_5967);
or U12057 (N_12057,N_6757,N_8981);
and U12058 (N_12058,N_7163,N_5274);
and U12059 (N_12059,N_7083,N_7011);
nand U12060 (N_12060,N_8280,N_8338);
xnor U12061 (N_12061,N_5564,N_6082);
nand U12062 (N_12062,N_6513,N_9730);
and U12063 (N_12063,N_8457,N_5506);
or U12064 (N_12064,N_8717,N_6880);
nand U12065 (N_12065,N_9007,N_5518);
xor U12066 (N_12066,N_6693,N_7788);
and U12067 (N_12067,N_9413,N_6724);
or U12068 (N_12068,N_7216,N_6095);
and U12069 (N_12069,N_7537,N_9154);
xnor U12070 (N_12070,N_6337,N_5626);
or U12071 (N_12071,N_5977,N_9369);
nand U12072 (N_12072,N_6946,N_7982);
xor U12073 (N_12073,N_7260,N_6433);
or U12074 (N_12074,N_9651,N_7974);
nor U12075 (N_12075,N_5725,N_6753);
nand U12076 (N_12076,N_7605,N_9061);
or U12077 (N_12077,N_9720,N_8328);
nor U12078 (N_12078,N_9364,N_5342);
or U12079 (N_12079,N_7973,N_7634);
or U12080 (N_12080,N_7068,N_7054);
xnor U12081 (N_12081,N_8624,N_5775);
and U12082 (N_12082,N_7876,N_9694);
xnor U12083 (N_12083,N_8323,N_9924);
nand U12084 (N_12084,N_5186,N_6465);
nand U12085 (N_12085,N_9390,N_5288);
nor U12086 (N_12086,N_5726,N_7409);
and U12087 (N_12087,N_8066,N_8110);
nor U12088 (N_12088,N_7869,N_7057);
nand U12089 (N_12089,N_8989,N_9778);
xnor U12090 (N_12090,N_7060,N_5607);
xnor U12091 (N_12091,N_8813,N_7828);
xnor U12092 (N_12092,N_6778,N_8088);
nand U12093 (N_12093,N_9766,N_7833);
and U12094 (N_12094,N_7597,N_7003);
or U12095 (N_12095,N_7472,N_7783);
xor U12096 (N_12096,N_6981,N_7779);
and U12097 (N_12097,N_7104,N_9260);
nand U12098 (N_12098,N_9184,N_9566);
xor U12099 (N_12099,N_9335,N_6938);
or U12100 (N_12100,N_6038,N_7347);
xor U12101 (N_12101,N_7839,N_8229);
nand U12102 (N_12102,N_8420,N_5295);
nand U12103 (N_12103,N_7277,N_7927);
nand U12104 (N_12104,N_5175,N_9664);
or U12105 (N_12105,N_8464,N_6759);
or U12106 (N_12106,N_6407,N_8265);
xor U12107 (N_12107,N_7194,N_8062);
or U12108 (N_12108,N_6147,N_8790);
nand U12109 (N_12109,N_9434,N_6896);
nor U12110 (N_12110,N_9992,N_5435);
and U12111 (N_12111,N_9483,N_8119);
or U12112 (N_12112,N_6248,N_5788);
nand U12113 (N_12113,N_5247,N_8757);
or U12114 (N_12114,N_7661,N_7387);
and U12115 (N_12115,N_6636,N_6780);
or U12116 (N_12116,N_8176,N_9311);
xnor U12117 (N_12117,N_8945,N_5710);
xor U12118 (N_12118,N_7643,N_6986);
or U12119 (N_12119,N_9783,N_7181);
nand U12120 (N_12120,N_8872,N_8530);
xor U12121 (N_12121,N_5415,N_8345);
nor U12122 (N_12122,N_8704,N_8894);
xor U12123 (N_12123,N_9615,N_9273);
nand U12124 (N_12124,N_7168,N_5510);
nand U12125 (N_12125,N_9798,N_5703);
nand U12126 (N_12126,N_6927,N_9614);
xor U12127 (N_12127,N_6346,N_7709);
and U12128 (N_12128,N_5050,N_8754);
or U12129 (N_12129,N_5692,N_8644);
and U12130 (N_12130,N_7165,N_8810);
xor U12131 (N_12131,N_8276,N_6497);
nand U12132 (N_12132,N_6053,N_6718);
nor U12133 (N_12133,N_8238,N_7579);
nand U12134 (N_12134,N_5104,N_7452);
xor U12135 (N_12135,N_5550,N_6450);
xnor U12136 (N_12136,N_8770,N_9817);
or U12137 (N_12137,N_7625,N_6205);
or U12138 (N_12138,N_7176,N_8374);
nand U12139 (N_12139,N_5278,N_6021);
xnor U12140 (N_12140,N_5188,N_6398);
nand U12141 (N_12141,N_8061,N_6506);
nor U12142 (N_12142,N_6691,N_8573);
and U12143 (N_12143,N_7388,N_9385);
or U12144 (N_12144,N_9013,N_8308);
nor U12145 (N_12145,N_6818,N_7428);
and U12146 (N_12146,N_8248,N_9853);
xnor U12147 (N_12147,N_8449,N_9684);
or U12148 (N_12148,N_6708,N_6546);
xor U12149 (N_12149,N_8642,N_8828);
nor U12150 (N_12150,N_6619,N_7056);
nor U12151 (N_12151,N_9012,N_6941);
or U12152 (N_12152,N_8198,N_8760);
nand U12153 (N_12153,N_9190,N_8448);
xnor U12154 (N_12154,N_6530,N_5412);
or U12155 (N_12155,N_5124,N_8359);
or U12156 (N_12156,N_9789,N_7243);
nand U12157 (N_12157,N_8257,N_9821);
and U12158 (N_12158,N_7286,N_7403);
and U12159 (N_12159,N_9272,N_6058);
or U12160 (N_12160,N_8657,N_6416);
or U12161 (N_12161,N_5786,N_7366);
xnor U12162 (N_12162,N_5402,N_9067);
nor U12163 (N_12163,N_5121,N_9374);
or U12164 (N_12164,N_7292,N_9805);
or U12165 (N_12165,N_9280,N_7851);
nand U12166 (N_12166,N_9677,N_5320);
or U12167 (N_12167,N_6788,N_6104);
and U12168 (N_12168,N_5766,N_5862);
and U12169 (N_12169,N_6212,N_6824);
nor U12170 (N_12170,N_5594,N_6911);
nor U12171 (N_12171,N_6102,N_8096);
and U12172 (N_12172,N_8007,N_8235);
nor U12173 (N_12173,N_7545,N_8285);
nand U12174 (N_12174,N_7599,N_7049);
nor U12175 (N_12175,N_5919,N_5972);
xor U12176 (N_12176,N_6103,N_6107);
xnor U12177 (N_12177,N_6700,N_7786);
nand U12178 (N_12178,N_9799,N_5056);
nand U12179 (N_12179,N_5694,N_8871);
nand U12180 (N_12180,N_9599,N_7079);
or U12181 (N_12181,N_7500,N_8187);
nor U12182 (N_12182,N_8791,N_8059);
xnor U12183 (N_12183,N_6112,N_9654);
and U12184 (N_12184,N_5653,N_6129);
nand U12185 (N_12185,N_5221,N_7808);
nor U12186 (N_12186,N_5812,N_9406);
nor U12187 (N_12187,N_6269,N_9948);
nand U12188 (N_12188,N_9193,N_6650);
and U12189 (N_12189,N_7123,N_6225);
and U12190 (N_12190,N_6444,N_7917);
nand U12191 (N_12191,N_5004,N_7722);
nor U12192 (N_12192,N_5312,N_8024);
or U12193 (N_12193,N_9072,N_8120);
nand U12194 (N_12194,N_9967,N_6006);
and U12195 (N_12195,N_6706,N_7746);
xnor U12196 (N_12196,N_6448,N_5804);
xnor U12197 (N_12197,N_7991,N_7819);
xnor U12198 (N_12198,N_7302,N_9166);
and U12199 (N_12199,N_6498,N_7220);
or U12200 (N_12200,N_9326,N_8980);
or U12201 (N_12201,N_9590,N_6758);
nor U12202 (N_12202,N_6964,N_7417);
or U12203 (N_12203,N_9333,N_6427);
xor U12204 (N_12204,N_9559,N_6438);
nor U12205 (N_12205,N_6924,N_9502);
nor U12206 (N_12206,N_9520,N_9639);
xor U12207 (N_12207,N_8369,N_9825);
and U12208 (N_12208,N_7415,N_8996);
nor U12209 (N_12209,N_5434,N_8486);
or U12210 (N_12210,N_7578,N_7609);
nand U12211 (N_12211,N_6819,N_9460);
or U12212 (N_12212,N_7666,N_9822);
or U12213 (N_12213,N_6937,N_7374);
or U12214 (N_12214,N_8135,N_7946);
nand U12215 (N_12215,N_8036,N_7384);
and U12216 (N_12216,N_8927,N_5462);
xnor U12217 (N_12217,N_6177,N_5593);
nand U12218 (N_12218,N_9291,N_7339);
nand U12219 (N_12219,N_9946,N_6186);
xor U12220 (N_12220,N_9426,N_7893);
or U12221 (N_12221,N_6303,N_9844);
nor U12222 (N_12222,N_5596,N_6558);
nand U12223 (N_12223,N_9936,N_9137);
xnor U12224 (N_12224,N_8057,N_8452);
or U12225 (N_12225,N_9352,N_9063);
and U12226 (N_12226,N_7631,N_9099);
nor U12227 (N_12227,N_7436,N_8467);
xnor U12228 (N_12228,N_5784,N_7015);
and U12229 (N_12229,N_6001,N_5077);
or U12230 (N_12230,N_9022,N_7429);
xor U12231 (N_12231,N_7192,N_7247);
xor U12232 (N_12232,N_8788,N_7361);
xor U12233 (N_12233,N_8990,N_7148);
or U12234 (N_12234,N_7560,N_9893);
or U12235 (N_12235,N_9452,N_6032);
or U12236 (N_12236,N_9062,N_8361);
xor U12237 (N_12237,N_8010,N_5328);
and U12238 (N_12238,N_6496,N_5999);
and U12239 (N_12239,N_5418,N_9508);
nor U12240 (N_12240,N_6121,N_5803);
or U12241 (N_12241,N_5588,N_6350);
nand U12242 (N_12242,N_6744,N_6207);
xor U12243 (N_12243,N_9427,N_5801);
and U12244 (N_12244,N_7394,N_5438);
nand U12245 (N_12245,N_9971,N_9031);
and U12246 (N_12246,N_5918,N_9628);
xor U12247 (N_12247,N_5132,N_6988);
nand U12248 (N_12248,N_9017,N_9372);
nand U12249 (N_12249,N_5417,N_8241);
or U12250 (N_12250,N_7559,N_8364);
xnor U12251 (N_12251,N_9330,N_9279);
nor U12252 (N_12252,N_7696,N_5630);
xor U12253 (N_12253,N_9514,N_6472);
xor U12254 (N_12254,N_9448,N_5774);
xnor U12255 (N_12255,N_7363,N_5076);
nand U12256 (N_12256,N_8332,N_6603);
nor U12257 (N_12257,N_5952,N_8144);
xnor U12258 (N_12258,N_7552,N_8735);
nor U12259 (N_12259,N_7837,N_8215);
and U12260 (N_12260,N_7454,N_9252);
and U12261 (N_12261,N_8742,N_8896);
nand U12262 (N_12262,N_9455,N_6218);
and U12263 (N_12263,N_9784,N_6867);
and U12264 (N_12264,N_8970,N_5136);
xnor U12265 (N_12265,N_9232,N_6987);
and U12266 (N_12266,N_7375,N_9560);
nor U12267 (N_12267,N_6203,N_6665);
and U12268 (N_12268,N_9961,N_9728);
xnor U12269 (N_12269,N_7914,N_6469);
xor U12270 (N_12270,N_7522,N_6263);
xor U12271 (N_12271,N_5143,N_5883);
or U12272 (N_12272,N_8843,N_7264);
or U12273 (N_12273,N_5802,N_5461);
and U12274 (N_12274,N_7879,N_9695);
nand U12275 (N_12275,N_5567,N_6649);
or U12276 (N_12276,N_9849,N_8570);
and U12277 (N_12277,N_6985,N_8579);
and U12278 (N_12278,N_6595,N_5229);
or U12279 (N_12279,N_6399,N_9659);
nand U12280 (N_12280,N_8906,N_7424);
xnor U12281 (N_12281,N_7744,N_9563);
and U12282 (N_12282,N_6072,N_7412);
xor U12283 (N_12283,N_9772,N_9608);
and U12284 (N_12284,N_7778,N_7515);
and U12285 (N_12285,N_8164,N_5932);
and U12286 (N_12286,N_9755,N_7768);
nor U12287 (N_12287,N_9582,N_5427);
and U12288 (N_12288,N_8123,N_5791);
and U12289 (N_12289,N_8663,N_9675);
or U12290 (N_12290,N_5681,N_7685);
and U12291 (N_12291,N_6772,N_6366);
nor U12292 (N_12292,N_7287,N_9146);
xnor U12293 (N_12293,N_7691,N_8311);
nand U12294 (N_12294,N_5352,N_9180);
or U12295 (N_12295,N_8225,N_9865);
and U12296 (N_12296,N_9069,N_7325);
xnor U12297 (N_12297,N_9932,N_7422);
nand U12298 (N_12298,N_7440,N_9842);
nor U12299 (N_12299,N_7529,N_6277);
and U12300 (N_12300,N_6943,N_6308);
nand U12301 (N_12301,N_5253,N_8382);
nand U12302 (N_12302,N_6251,N_7872);
or U12303 (N_12303,N_6846,N_6417);
and U12304 (N_12304,N_9464,N_6682);
nor U12305 (N_12305,N_6372,N_9351);
or U12306 (N_12306,N_8325,N_7862);
or U12307 (N_12307,N_8845,N_7790);
nand U12308 (N_12308,N_9191,N_9518);
xnor U12309 (N_12309,N_7567,N_8614);
nor U12310 (N_12310,N_9693,N_5910);
nand U12311 (N_12311,N_7153,N_8397);
nand U12312 (N_12312,N_9891,N_9545);
or U12313 (N_12313,N_7700,N_8174);
and U12314 (N_12314,N_7467,N_6482);
and U12315 (N_12315,N_6080,N_5177);
and U12316 (N_12316,N_5036,N_8517);
or U12317 (N_12317,N_8445,N_7336);
nand U12318 (N_12318,N_6770,N_9752);
nand U12319 (N_12319,N_9303,N_6844);
nor U12320 (N_12320,N_8362,N_7532);
and U12321 (N_12321,N_7152,N_9290);
nor U12322 (N_12322,N_5087,N_5997);
nor U12323 (N_12323,N_7298,N_6774);
nor U12324 (N_12324,N_7480,N_5505);
xor U12325 (N_12325,N_5817,N_9030);
xor U12326 (N_12326,N_8484,N_7909);
nor U12327 (N_12327,N_9153,N_8404);
xor U12328 (N_12328,N_6049,N_5732);
nor U12329 (N_12329,N_8188,N_8661);
and U12330 (N_12330,N_5131,N_6243);
nor U12331 (N_12331,N_5331,N_6719);
or U12332 (N_12332,N_6763,N_7059);
xnor U12333 (N_12333,N_5598,N_6680);
xnor U12334 (N_12334,N_5002,N_7704);
or U12335 (N_12335,N_9027,N_6544);
and U12336 (N_12336,N_9048,N_7261);
and U12337 (N_12337,N_8858,N_8242);
xor U12338 (N_12338,N_8582,N_9297);
or U12339 (N_12339,N_9185,N_8716);
xnor U12340 (N_12340,N_6522,N_8559);
or U12341 (N_12341,N_6667,N_6710);
nor U12342 (N_12342,N_7994,N_5978);
or U12343 (N_12343,N_6536,N_9147);
and U12344 (N_12344,N_6604,N_5291);
nor U12345 (N_12345,N_5778,N_7619);
xor U12346 (N_12346,N_8479,N_5923);
xnor U12347 (N_12347,N_7455,N_6258);
and U12348 (N_12348,N_9397,N_7847);
nor U12349 (N_12349,N_7461,N_6799);
nor U12350 (N_12350,N_6743,N_6343);
and U12351 (N_12351,N_9500,N_6408);
nand U12352 (N_12352,N_5207,N_5805);
and U12353 (N_12353,N_8853,N_9718);
xnor U12354 (N_12354,N_5500,N_7616);
xnor U12355 (N_12355,N_9054,N_7045);
xor U12356 (N_12356,N_7614,N_7030);
or U12357 (N_12357,N_8763,N_5921);
and U12358 (N_12358,N_6963,N_5406);
and U12359 (N_12359,N_5936,N_6740);
or U12360 (N_12360,N_6341,N_9231);
xor U12361 (N_12361,N_8786,N_5686);
nand U12362 (N_12362,N_9468,N_8358);
nand U12363 (N_12363,N_9873,N_7693);
nand U12364 (N_12364,N_5965,N_6537);
xor U12365 (N_12365,N_7105,N_7554);
or U12366 (N_12366,N_8830,N_7555);
nand U12367 (N_12367,N_6014,N_5979);
or U12368 (N_12368,N_9771,N_6106);
or U12369 (N_12369,N_9334,N_5126);
xnor U12370 (N_12370,N_5898,N_8956);
xnor U12371 (N_12371,N_9316,N_5394);
nor U12372 (N_12372,N_7242,N_7541);
xnor U12373 (N_12373,N_7810,N_9954);
nand U12374 (N_12374,N_5014,N_5612);
nand U12375 (N_12375,N_5895,N_5325);
or U12376 (N_12376,N_8516,N_6615);
nand U12377 (N_12377,N_6000,N_6093);
nor U12378 (N_12378,N_6487,N_7659);
nor U12379 (N_12379,N_8918,N_6950);
or U12380 (N_12380,N_7861,N_7418);
nor U12381 (N_12381,N_7863,N_5335);
nand U12382 (N_12382,N_7420,N_5363);
nand U12383 (N_12383,N_6955,N_6252);
or U12384 (N_12384,N_7799,N_8356);
nor U12385 (N_12385,N_7229,N_9181);
or U12386 (N_12386,N_5857,N_8563);
nand U12387 (N_12387,N_9503,N_7855);
xnor U12388 (N_12388,N_6642,N_6782);
nand U12389 (N_12389,N_7950,N_8873);
or U12390 (N_12390,N_6304,N_5713);
xor U12391 (N_12391,N_6204,N_5332);
xnor U12392 (N_12392,N_7655,N_6271);
nand U12393 (N_12393,N_7756,N_9053);
nor U12394 (N_12394,N_7382,N_8127);
or U12395 (N_12395,N_8805,N_7954);
nand U12396 (N_12396,N_8506,N_9925);
nand U12397 (N_12397,N_7154,N_5925);
nand U12398 (N_12398,N_6503,N_9512);
nand U12399 (N_12399,N_9605,N_8383);
or U12400 (N_12400,N_7564,N_9287);
nand U12401 (N_12401,N_9315,N_8064);
or U12402 (N_12402,N_6406,N_5443);
or U12403 (N_12403,N_6424,N_8243);
or U12404 (N_12404,N_6010,N_8351);
or U12405 (N_12405,N_9753,N_7802);
xor U12406 (N_12406,N_8940,N_9792);
and U12407 (N_12407,N_8201,N_7935);
and U12408 (N_12408,N_7891,N_8562);
nand U12409 (N_12409,N_6020,N_7870);
nand U12410 (N_12410,N_9737,N_6656);
and U12411 (N_12411,N_5233,N_9200);
nand U12412 (N_12412,N_5826,N_5155);
xor U12413 (N_12413,N_6138,N_8245);
and U12414 (N_12414,N_6548,N_6578);
nand U12415 (N_12415,N_6461,N_8025);
nor U12416 (N_12416,N_9683,N_5096);
or U12417 (N_12417,N_9320,N_8919);
or U12418 (N_12418,N_5467,N_5908);
or U12419 (N_12419,N_6054,N_5283);
xor U12420 (N_12420,N_5855,N_9060);
and U12421 (N_12421,N_5408,N_7534);
nor U12422 (N_12422,N_6611,N_6037);
xnor U12423 (N_12423,N_7571,N_6532);
or U12424 (N_12424,N_7968,N_6253);
nor U12425 (N_12425,N_7368,N_6531);
nand U12426 (N_12426,N_9183,N_9658);
nor U12427 (N_12427,N_6504,N_9904);
and U12428 (N_12428,N_5948,N_8271);
and U12429 (N_12429,N_9596,N_9619);
xor U12430 (N_12430,N_8014,N_5451);
or U12431 (N_12431,N_7359,N_8172);
nor U12432 (N_12432,N_5547,N_9292);
and U12433 (N_12433,N_9093,N_9841);
xor U12434 (N_12434,N_6067,N_8524);
and U12435 (N_12435,N_8501,N_6734);
and U12436 (N_12436,N_8104,N_6735);
and U12437 (N_12437,N_6352,N_7987);
nor U12438 (N_12438,N_5465,N_8487);
and U12439 (N_12439,N_7766,N_6338);
or U12440 (N_12440,N_7489,N_7787);
nand U12441 (N_12441,N_7795,N_6833);
nor U12442 (N_12442,N_6278,N_6618);
nand U12443 (N_12443,N_7523,N_5387);
nand U12444 (N_12444,N_5882,N_8574);
nand U12445 (N_12445,N_5917,N_5808);
nor U12446 (N_12446,N_7886,N_9524);
nand U12447 (N_12447,N_6555,N_9047);
and U12448 (N_12448,N_5690,N_5958);
and U12449 (N_12449,N_8874,N_8859);
nor U12450 (N_12450,N_5103,N_8997);
or U12451 (N_12451,N_6610,N_7340);
nor U12452 (N_12452,N_7832,N_7715);
nor U12453 (N_12453,N_6301,N_7574);
xor U12454 (N_12454,N_8774,N_5058);
nand U12455 (N_12455,N_7106,N_9318);
or U12456 (N_12456,N_8137,N_7568);
and U12457 (N_12457,N_9209,N_5879);
and U12458 (N_12458,N_7416,N_8149);
nor U12459 (N_12459,N_5133,N_6934);
nor U12460 (N_12460,N_9439,N_6451);
nor U12461 (N_12461,N_9571,N_5529);
or U12462 (N_12462,N_9803,N_8523);
xnor U12463 (N_12463,N_6811,N_6895);
nand U12464 (N_12464,N_8208,N_7977);
xor U12465 (N_12465,N_7485,N_9355);
nor U12466 (N_12466,N_5145,N_5297);
and U12467 (N_12467,N_5799,N_5152);
nor U12468 (N_12468,N_7465,N_9603);
nand U12469 (N_12469,N_8821,N_7128);
and U12470 (N_12470,N_8652,N_5107);
xor U12471 (N_12471,N_5634,N_9375);
or U12472 (N_12472,N_8878,N_9098);
xor U12473 (N_12473,N_8386,N_5254);
nor U12474 (N_12474,N_5038,N_6202);
nor U12475 (N_12475,N_5487,N_9949);
nor U12476 (N_12476,N_5845,N_7680);
nor U12477 (N_12477,N_8264,N_9890);
or U12478 (N_12478,N_6745,N_9609);
nand U12479 (N_12479,N_6091,N_8728);
nand U12480 (N_12480,N_8433,N_6231);
or U12481 (N_12481,N_7175,N_6676);
and U12482 (N_12482,N_8783,N_6870);
or U12483 (N_12483,N_9713,N_9217);
and U12484 (N_12484,N_5838,N_7014);
nor U12485 (N_12485,N_7391,N_7754);
nand U12486 (N_12486,N_9845,N_7710);
nor U12487 (N_12487,N_5360,N_5930);
and U12488 (N_12488,N_9581,N_9214);
and U12489 (N_12489,N_6449,N_8617);
or U12490 (N_12490,N_8017,N_5606);
nand U12491 (N_12491,N_6355,N_6052);
nand U12492 (N_12492,N_9284,N_9170);
and U12493 (N_12493,N_6409,N_9835);
nand U12494 (N_12494,N_9338,N_5632);
and U12495 (N_12495,N_8909,N_5053);
nor U12496 (N_12496,N_9042,N_8561);
xor U12497 (N_12497,N_6944,N_7089);
nand U12498 (N_12498,N_5738,N_6756);
and U12499 (N_12499,N_9643,N_6751);
or U12500 (N_12500,N_8342,N_7992);
or U12501 (N_12501,N_6462,N_6868);
xor U12502 (N_12502,N_7396,N_8661);
nand U12503 (N_12503,N_9544,N_5088);
xor U12504 (N_12504,N_9723,N_7666);
nor U12505 (N_12505,N_9634,N_9078);
and U12506 (N_12506,N_9973,N_9487);
xor U12507 (N_12507,N_7593,N_9734);
nand U12508 (N_12508,N_5370,N_5058);
or U12509 (N_12509,N_7387,N_5638);
nand U12510 (N_12510,N_5347,N_5390);
nor U12511 (N_12511,N_6774,N_6878);
nor U12512 (N_12512,N_5975,N_8391);
nand U12513 (N_12513,N_7251,N_7421);
nor U12514 (N_12514,N_8916,N_7479);
or U12515 (N_12515,N_8571,N_9585);
nand U12516 (N_12516,N_9153,N_8179);
xor U12517 (N_12517,N_9567,N_6449);
nor U12518 (N_12518,N_8463,N_9551);
nand U12519 (N_12519,N_5804,N_5057);
nor U12520 (N_12520,N_7936,N_6783);
and U12521 (N_12521,N_8748,N_9293);
nor U12522 (N_12522,N_5082,N_9895);
or U12523 (N_12523,N_5830,N_8810);
nor U12524 (N_12524,N_8756,N_9564);
nor U12525 (N_12525,N_5198,N_7959);
and U12526 (N_12526,N_8869,N_6183);
or U12527 (N_12527,N_9746,N_9053);
nor U12528 (N_12528,N_6175,N_8910);
nand U12529 (N_12529,N_5918,N_9828);
or U12530 (N_12530,N_9554,N_6061);
nand U12531 (N_12531,N_9558,N_5220);
nand U12532 (N_12532,N_6773,N_9634);
xnor U12533 (N_12533,N_8550,N_7754);
and U12534 (N_12534,N_7359,N_6715);
and U12535 (N_12535,N_8596,N_5949);
nor U12536 (N_12536,N_6420,N_9645);
and U12537 (N_12537,N_5017,N_8740);
nand U12538 (N_12538,N_7349,N_6433);
nand U12539 (N_12539,N_6083,N_8831);
xnor U12540 (N_12540,N_7068,N_9997);
and U12541 (N_12541,N_6331,N_9050);
nand U12542 (N_12542,N_8281,N_7485);
nand U12543 (N_12543,N_8321,N_8727);
nor U12544 (N_12544,N_8739,N_9899);
xor U12545 (N_12545,N_6362,N_8543);
or U12546 (N_12546,N_6590,N_9026);
and U12547 (N_12547,N_5724,N_6561);
nand U12548 (N_12548,N_6070,N_9859);
nor U12549 (N_12549,N_6526,N_6140);
and U12550 (N_12550,N_8168,N_6349);
nand U12551 (N_12551,N_5842,N_6683);
xnor U12552 (N_12552,N_8990,N_8977);
or U12553 (N_12553,N_8838,N_6373);
or U12554 (N_12554,N_9846,N_9219);
or U12555 (N_12555,N_8474,N_7447);
or U12556 (N_12556,N_8362,N_9826);
nor U12557 (N_12557,N_7389,N_8821);
or U12558 (N_12558,N_8732,N_8429);
nand U12559 (N_12559,N_8573,N_7467);
xnor U12560 (N_12560,N_6618,N_5526);
or U12561 (N_12561,N_6360,N_7427);
and U12562 (N_12562,N_5318,N_5379);
and U12563 (N_12563,N_5677,N_6018);
xnor U12564 (N_12564,N_5366,N_5510);
nand U12565 (N_12565,N_9713,N_5633);
or U12566 (N_12566,N_9030,N_9306);
and U12567 (N_12567,N_6670,N_5338);
or U12568 (N_12568,N_8808,N_5745);
and U12569 (N_12569,N_6544,N_7639);
or U12570 (N_12570,N_7325,N_9616);
nand U12571 (N_12571,N_9394,N_9000);
or U12572 (N_12572,N_9845,N_5444);
or U12573 (N_12573,N_9630,N_7778);
nor U12574 (N_12574,N_5269,N_8901);
nor U12575 (N_12575,N_5093,N_5811);
or U12576 (N_12576,N_9251,N_9107);
and U12577 (N_12577,N_5805,N_7744);
nor U12578 (N_12578,N_8734,N_5606);
and U12579 (N_12579,N_8461,N_6092);
xnor U12580 (N_12580,N_8454,N_7655);
xnor U12581 (N_12581,N_8980,N_9040);
or U12582 (N_12582,N_6338,N_6214);
xnor U12583 (N_12583,N_7839,N_9229);
nor U12584 (N_12584,N_6953,N_7604);
xnor U12585 (N_12585,N_5623,N_8577);
or U12586 (N_12586,N_5588,N_7749);
nor U12587 (N_12587,N_8868,N_5521);
or U12588 (N_12588,N_7407,N_5013);
and U12589 (N_12589,N_9722,N_7947);
nor U12590 (N_12590,N_6015,N_9487);
nor U12591 (N_12591,N_5348,N_8676);
or U12592 (N_12592,N_7861,N_8970);
or U12593 (N_12593,N_5886,N_7967);
or U12594 (N_12594,N_6410,N_5107);
and U12595 (N_12595,N_5192,N_6616);
xnor U12596 (N_12596,N_9589,N_8026);
and U12597 (N_12597,N_9255,N_8994);
or U12598 (N_12598,N_6884,N_5009);
xor U12599 (N_12599,N_7572,N_7918);
nand U12600 (N_12600,N_5979,N_6571);
and U12601 (N_12601,N_6489,N_9231);
nor U12602 (N_12602,N_9722,N_5417);
nor U12603 (N_12603,N_5519,N_7741);
nor U12604 (N_12604,N_9067,N_5810);
or U12605 (N_12605,N_6497,N_5474);
and U12606 (N_12606,N_6793,N_7427);
or U12607 (N_12607,N_5656,N_5959);
nand U12608 (N_12608,N_9852,N_7411);
xor U12609 (N_12609,N_7116,N_5020);
xnor U12610 (N_12610,N_6109,N_9545);
xor U12611 (N_12611,N_7646,N_5079);
xor U12612 (N_12612,N_6183,N_6992);
or U12613 (N_12613,N_5087,N_7306);
or U12614 (N_12614,N_9103,N_8419);
xor U12615 (N_12615,N_6252,N_5746);
or U12616 (N_12616,N_5800,N_7198);
and U12617 (N_12617,N_5792,N_7562);
and U12618 (N_12618,N_9377,N_8680);
nor U12619 (N_12619,N_6961,N_7828);
nand U12620 (N_12620,N_9290,N_9419);
nand U12621 (N_12621,N_6350,N_8546);
and U12622 (N_12622,N_9106,N_6438);
xnor U12623 (N_12623,N_9662,N_7642);
or U12624 (N_12624,N_8602,N_5272);
and U12625 (N_12625,N_7181,N_8122);
or U12626 (N_12626,N_6316,N_7646);
or U12627 (N_12627,N_5622,N_9110);
and U12628 (N_12628,N_7491,N_8434);
nand U12629 (N_12629,N_8358,N_6155);
xnor U12630 (N_12630,N_7279,N_9327);
nor U12631 (N_12631,N_5625,N_7866);
nand U12632 (N_12632,N_5859,N_5715);
xnor U12633 (N_12633,N_5409,N_5522);
nand U12634 (N_12634,N_8719,N_5250);
or U12635 (N_12635,N_9304,N_7348);
nor U12636 (N_12636,N_5946,N_7699);
and U12637 (N_12637,N_5509,N_8309);
nand U12638 (N_12638,N_9561,N_6251);
xor U12639 (N_12639,N_8451,N_9400);
xnor U12640 (N_12640,N_7193,N_7138);
nor U12641 (N_12641,N_9206,N_5743);
or U12642 (N_12642,N_8812,N_8228);
xor U12643 (N_12643,N_5386,N_6806);
nor U12644 (N_12644,N_5736,N_9906);
xor U12645 (N_12645,N_5740,N_7943);
nor U12646 (N_12646,N_5700,N_9829);
xnor U12647 (N_12647,N_8721,N_6394);
xnor U12648 (N_12648,N_5538,N_9342);
xnor U12649 (N_12649,N_9243,N_5938);
xnor U12650 (N_12650,N_5977,N_7997);
nand U12651 (N_12651,N_7214,N_7852);
and U12652 (N_12652,N_9290,N_5564);
or U12653 (N_12653,N_8556,N_8853);
or U12654 (N_12654,N_5714,N_7163);
or U12655 (N_12655,N_9605,N_9686);
nand U12656 (N_12656,N_9704,N_9996);
xor U12657 (N_12657,N_7151,N_8246);
and U12658 (N_12658,N_5454,N_9279);
xor U12659 (N_12659,N_8906,N_5361);
or U12660 (N_12660,N_6051,N_7687);
xnor U12661 (N_12661,N_5787,N_9453);
and U12662 (N_12662,N_6390,N_8958);
xnor U12663 (N_12663,N_9738,N_6558);
or U12664 (N_12664,N_7721,N_8186);
nand U12665 (N_12665,N_6180,N_8189);
and U12666 (N_12666,N_8010,N_5701);
xnor U12667 (N_12667,N_8634,N_6637);
and U12668 (N_12668,N_9835,N_7060);
nand U12669 (N_12669,N_9787,N_6573);
or U12670 (N_12670,N_5986,N_9702);
nand U12671 (N_12671,N_9025,N_7082);
nor U12672 (N_12672,N_6330,N_9032);
and U12673 (N_12673,N_7552,N_7516);
and U12674 (N_12674,N_5955,N_5799);
and U12675 (N_12675,N_7418,N_5913);
nand U12676 (N_12676,N_9022,N_5617);
or U12677 (N_12677,N_5071,N_5857);
nor U12678 (N_12678,N_8144,N_5943);
nor U12679 (N_12679,N_9209,N_6260);
and U12680 (N_12680,N_8914,N_6336);
nand U12681 (N_12681,N_8851,N_7333);
nand U12682 (N_12682,N_5722,N_7409);
and U12683 (N_12683,N_8214,N_8090);
nand U12684 (N_12684,N_6189,N_8305);
or U12685 (N_12685,N_9313,N_8786);
nand U12686 (N_12686,N_6578,N_5706);
nor U12687 (N_12687,N_6570,N_9986);
nand U12688 (N_12688,N_9341,N_9657);
or U12689 (N_12689,N_6652,N_9048);
nand U12690 (N_12690,N_6084,N_5307);
nand U12691 (N_12691,N_8343,N_5012);
and U12692 (N_12692,N_7684,N_6019);
nor U12693 (N_12693,N_7075,N_9062);
nor U12694 (N_12694,N_5877,N_6370);
or U12695 (N_12695,N_6954,N_7743);
xor U12696 (N_12696,N_7938,N_8791);
or U12697 (N_12697,N_8978,N_5549);
or U12698 (N_12698,N_9114,N_6461);
and U12699 (N_12699,N_6161,N_5678);
and U12700 (N_12700,N_7778,N_8595);
or U12701 (N_12701,N_8417,N_8996);
or U12702 (N_12702,N_9541,N_9978);
nor U12703 (N_12703,N_5008,N_6505);
nand U12704 (N_12704,N_6205,N_8003);
nand U12705 (N_12705,N_6177,N_8523);
and U12706 (N_12706,N_9468,N_9622);
nand U12707 (N_12707,N_8326,N_6625);
nand U12708 (N_12708,N_9756,N_8761);
nor U12709 (N_12709,N_6623,N_8454);
nand U12710 (N_12710,N_8016,N_5421);
nor U12711 (N_12711,N_5413,N_5005);
nor U12712 (N_12712,N_5686,N_9016);
nand U12713 (N_12713,N_6007,N_9845);
xnor U12714 (N_12714,N_7503,N_9596);
or U12715 (N_12715,N_9160,N_5612);
and U12716 (N_12716,N_6038,N_5036);
nor U12717 (N_12717,N_6526,N_8490);
and U12718 (N_12718,N_8539,N_5607);
or U12719 (N_12719,N_8667,N_6524);
or U12720 (N_12720,N_5637,N_5592);
or U12721 (N_12721,N_6964,N_7808);
xor U12722 (N_12722,N_6992,N_8177);
or U12723 (N_12723,N_8610,N_7703);
nor U12724 (N_12724,N_9548,N_8687);
nand U12725 (N_12725,N_5444,N_6476);
xnor U12726 (N_12726,N_8814,N_7164);
xnor U12727 (N_12727,N_7038,N_8317);
or U12728 (N_12728,N_6828,N_9555);
or U12729 (N_12729,N_6759,N_8696);
nor U12730 (N_12730,N_7246,N_6117);
nor U12731 (N_12731,N_5658,N_9122);
or U12732 (N_12732,N_6858,N_7358);
and U12733 (N_12733,N_6920,N_8021);
or U12734 (N_12734,N_8427,N_5088);
nand U12735 (N_12735,N_5243,N_7439);
nand U12736 (N_12736,N_5450,N_7308);
and U12737 (N_12737,N_6774,N_6775);
xnor U12738 (N_12738,N_8740,N_5910);
nand U12739 (N_12739,N_5941,N_9104);
or U12740 (N_12740,N_8855,N_6617);
nor U12741 (N_12741,N_5166,N_8764);
nor U12742 (N_12742,N_6913,N_9429);
or U12743 (N_12743,N_6272,N_7362);
xor U12744 (N_12744,N_7391,N_9106);
or U12745 (N_12745,N_8407,N_5066);
nor U12746 (N_12746,N_8610,N_6611);
nor U12747 (N_12747,N_6930,N_5135);
and U12748 (N_12748,N_9520,N_9559);
xor U12749 (N_12749,N_9242,N_9084);
nor U12750 (N_12750,N_8567,N_7935);
or U12751 (N_12751,N_8658,N_9636);
or U12752 (N_12752,N_6641,N_5676);
xnor U12753 (N_12753,N_8318,N_7876);
nor U12754 (N_12754,N_9348,N_5923);
nand U12755 (N_12755,N_7252,N_9168);
xor U12756 (N_12756,N_9277,N_8520);
or U12757 (N_12757,N_7688,N_6542);
nor U12758 (N_12758,N_7912,N_8287);
or U12759 (N_12759,N_9256,N_9330);
or U12760 (N_12760,N_8105,N_9032);
or U12761 (N_12761,N_5194,N_7109);
nand U12762 (N_12762,N_8053,N_5866);
or U12763 (N_12763,N_7709,N_6757);
nand U12764 (N_12764,N_9230,N_9186);
xor U12765 (N_12765,N_5198,N_7023);
xnor U12766 (N_12766,N_9235,N_5523);
nand U12767 (N_12767,N_5969,N_8013);
nor U12768 (N_12768,N_9176,N_5454);
or U12769 (N_12769,N_5447,N_5953);
nand U12770 (N_12770,N_5391,N_6640);
nand U12771 (N_12771,N_5674,N_5210);
nand U12772 (N_12772,N_8095,N_6633);
nand U12773 (N_12773,N_7121,N_7008);
nor U12774 (N_12774,N_8909,N_6543);
xor U12775 (N_12775,N_5688,N_6972);
or U12776 (N_12776,N_5157,N_5464);
nor U12777 (N_12777,N_6173,N_5710);
and U12778 (N_12778,N_5299,N_5988);
or U12779 (N_12779,N_8780,N_5914);
nor U12780 (N_12780,N_6782,N_5013);
or U12781 (N_12781,N_9517,N_8576);
and U12782 (N_12782,N_9947,N_6763);
or U12783 (N_12783,N_8130,N_9889);
nand U12784 (N_12784,N_6055,N_5342);
nand U12785 (N_12785,N_6851,N_9335);
nor U12786 (N_12786,N_9683,N_9201);
and U12787 (N_12787,N_9785,N_5294);
and U12788 (N_12788,N_6424,N_9995);
or U12789 (N_12789,N_9664,N_5915);
and U12790 (N_12790,N_5682,N_7007);
nor U12791 (N_12791,N_9061,N_7027);
or U12792 (N_12792,N_6137,N_6072);
nand U12793 (N_12793,N_8415,N_7703);
nor U12794 (N_12794,N_9296,N_8510);
xor U12795 (N_12795,N_8725,N_9641);
and U12796 (N_12796,N_7639,N_8928);
nor U12797 (N_12797,N_7360,N_9666);
or U12798 (N_12798,N_6691,N_5179);
nand U12799 (N_12799,N_5929,N_8912);
and U12800 (N_12800,N_9142,N_8409);
and U12801 (N_12801,N_9785,N_8562);
nor U12802 (N_12802,N_8377,N_8686);
nor U12803 (N_12803,N_5129,N_9725);
and U12804 (N_12804,N_9501,N_6223);
and U12805 (N_12805,N_6138,N_8326);
or U12806 (N_12806,N_9197,N_7970);
and U12807 (N_12807,N_6269,N_6588);
nand U12808 (N_12808,N_6889,N_7926);
or U12809 (N_12809,N_7156,N_7007);
nand U12810 (N_12810,N_5653,N_8660);
or U12811 (N_12811,N_7922,N_9903);
xor U12812 (N_12812,N_9194,N_8790);
xor U12813 (N_12813,N_8509,N_5484);
xnor U12814 (N_12814,N_8751,N_5993);
xor U12815 (N_12815,N_6561,N_5630);
nor U12816 (N_12816,N_9637,N_5854);
and U12817 (N_12817,N_6327,N_6371);
xnor U12818 (N_12818,N_7618,N_9356);
and U12819 (N_12819,N_8699,N_5664);
xnor U12820 (N_12820,N_9651,N_6295);
or U12821 (N_12821,N_7448,N_6823);
xnor U12822 (N_12822,N_5227,N_5941);
or U12823 (N_12823,N_9480,N_7038);
nor U12824 (N_12824,N_5228,N_6160);
and U12825 (N_12825,N_9922,N_6821);
and U12826 (N_12826,N_5309,N_6844);
nand U12827 (N_12827,N_8493,N_9615);
nor U12828 (N_12828,N_7272,N_8894);
nand U12829 (N_12829,N_5712,N_8786);
or U12830 (N_12830,N_5025,N_5982);
nor U12831 (N_12831,N_8852,N_9848);
nand U12832 (N_12832,N_5322,N_6200);
nand U12833 (N_12833,N_6417,N_6306);
nor U12834 (N_12834,N_6160,N_6279);
nand U12835 (N_12835,N_8726,N_5344);
or U12836 (N_12836,N_6161,N_6587);
or U12837 (N_12837,N_7393,N_6460);
and U12838 (N_12838,N_8569,N_9219);
nand U12839 (N_12839,N_8773,N_6540);
nand U12840 (N_12840,N_7507,N_8395);
and U12841 (N_12841,N_9201,N_8590);
and U12842 (N_12842,N_6042,N_7209);
xor U12843 (N_12843,N_7419,N_7835);
xnor U12844 (N_12844,N_9772,N_7755);
and U12845 (N_12845,N_8951,N_8350);
xnor U12846 (N_12846,N_5092,N_8793);
and U12847 (N_12847,N_7154,N_7312);
or U12848 (N_12848,N_7072,N_5263);
and U12849 (N_12849,N_8794,N_6585);
xor U12850 (N_12850,N_7284,N_8060);
and U12851 (N_12851,N_8566,N_9117);
and U12852 (N_12852,N_8478,N_8814);
nand U12853 (N_12853,N_9003,N_8630);
and U12854 (N_12854,N_8146,N_6489);
nand U12855 (N_12855,N_8066,N_9266);
nor U12856 (N_12856,N_8229,N_7430);
or U12857 (N_12857,N_5186,N_7954);
xnor U12858 (N_12858,N_9872,N_6518);
or U12859 (N_12859,N_8874,N_6541);
nand U12860 (N_12860,N_9541,N_5426);
nor U12861 (N_12861,N_7722,N_6466);
nand U12862 (N_12862,N_7778,N_9558);
xor U12863 (N_12863,N_6518,N_7863);
or U12864 (N_12864,N_8349,N_8620);
nand U12865 (N_12865,N_8178,N_5665);
nand U12866 (N_12866,N_8012,N_8787);
and U12867 (N_12867,N_6041,N_7084);
nor U12868 (N_12868,N_6196,N_7784);
nand U12869 (N_12869,N_6557,N_9760);
xor U12870 (N_12870,N_6822,N_5245);
nor U12871 (N_12871,N_8830,N_5873);
nor U12872 (N_12872,N_6573,N_5621);
xnor U12873 (N_12873,N_6833,N_5083);
and U12874 (N_12874,N_7243,N_9617);
nor U12875 (N_12875,N_5342,N_5872);
or U12876 (N_12876,N_8517,N_6164);
nor U12877 (N_12877,N_6288,N_8353);
and U12878 (N_12878,N_9709,N_6219);
xnor U12879 (N_12879,N_6270,N_8166);
xor U12880 (N_12880,N_7906,N_8859);
and U12881 (N_12881,N_8931,N_9180);
or U12882 (N_12882,N_7008,N_6669);
nand U12883 (N_12883,N_9724,N_6833);
or U12884 (N_12884,N_9588,N_6718);
and U12885 (N_12885,N_7890,N_9390);
xnor U12886 (N_12886,N_5064,N_8291);
or U12887 (N_12887,N_8046,N_5348);
nand U12888 (N_12888,N_9851,N_6596);
or U12889 (N_12889,N_8613,N_6783);
or U12890 (N_12890,N_5454,N_8304);
and U12891 (N_12891,N_8039,N_5148);
nor U12892 (N_12892,N_7535,N_5874);
nor U12893 (N_12893,N_5880,N_5338);
nand U12894 (N_12894,N_5164,N_8818);
or U12895 (N_12895,N_8498,N_6867);
xor U12896 (N_12896,N_7103,N_7200);
and U12897 (N_12897,N_9275,N_9003);
nor U12898 (N_12898,N_7241,N_7046);
or U12899 (N_12899,N_6534,N_8102);
nand U12900 (N_12900,N_5045,N_6879);
or U12901 (N_12901,N_6291,N_5180);
and U12902 (N_12902,N_6501,N_7957);
xor U12903 (N_12903,N_7802,N_8141);
nand U12904 (N_12904,N_9690,N_8849);
xnor U12905 (N_12905,N_7106,N_9057);
nor U12906 (N_12906,N_5141,N_7384);
nand U12907 (N_12907,N_8706,N_7755);
xor U12908 (N_12908,N_8497,N_7097);
and U12909 (N_12909,N_7996,N_5724);
nor U12910 (N_12910,N_9038,N_5215);
nand U12911 (N_12911,N_9920,N_7778);
or U12912 (N_12912,N_5023,N_7157);
and U12913 (N_12913,N_5778,N_7120);
or U12914 (N_12914,N_6798,N_8627);
or U12915 (N_12915,N_6048,N_9166);
or U12916 (N_12916,N_6328,N_9113);
xor U12917 (N_12917,N_8443,N_8238);
nand U12918 (N_12918,N_8537,N_8478);
nor U12919 (N_12919,N_5212,N_7488);
and U12920 (N_12920,N_6755,N_8486);
xnor U12921 (N_12921,N_6815,N_7772);
nand U12922 (N_12922,N_9549,N_7333);
xnor U12923 (N_12923,N_5529,N_7903);
nor U12924 (N_12924,N_6141,N_6469);
nand U12925 (N_12925,N_5147,N_6452);
and U12926 (N_12926,N_7070,N_6795);
and U12927 (N_12927,N_6279,N_6445);
and U12928 (N_12928,N_7706,N_7686);
or U12929 (N_12929,N_7241,N_8472);
nor U12930 (N_12930,N_6527,N_7246);
nand U12931 (N_12931,N_9289,N_5342);
or U12932 (N_12932,N_6174,N_6760);
and U12933 (N_12933,N_9685,N_5114);
xnor U12934 (N_12934,N_6735,N_8863);
nand U12935 (N_12935,N_6225,N_8935);
or U12936 (N_12936,N_7744,N_5719);
xnor U12937 (N_12937,N_5677,N_5938);
nand U12938 (N_12938,N_5545,N_6207);
nand U12939 (N_12939,N_6899,N_9986);
nor U12940 (N_12940,N_6853,N_7907);
nand U12941 (N_12941,N_9034,N_7985);
and U12942 (N_12942,N_6452,N_8542);
or U12943 (N_12943,N_8657,N_9663);
nand U12944 (N_12944,N_6440,N_7439);
nand U12945 (N_12945,N_8335,N_9869);
and U12946 (N_12946,N_8927,N_8058);
nor U12947 (N_12947,N_5866,N_8560);
nand U12948 (N_12948,N_6973,N_7359);
or U12949 (N_12949,N_9172,N_5631);
nor U12950 (N_12950,N_9383,N_9313);
xor U12951 (N_12951,N_9247,N_5746);
nor U12952 (N_12952,N_8392,N_7787);
and U12953 (N_12953,N_9577,N_5619);
nor U12954 (N_12954,N_7965,N_7564);
and U12955 (N_12955,N_8992,N_6366);
xor U12956 (N_12956,N_9987,N_9684);
nor U12957 (N_12957,N_6808,N_7162);
or U12958 (N_12958,N_6412,N_5199);
or U12959 (N_12959,N_9626,N_8919);
nor U12960 (N_12960,N_8868,N_8936);
and U12961 (N_12961,N_7895,N_5209);
xnor U12962 (N_12962,N_9388,N_6972);
nor U12963 (N_12963,N_9939,N_9064);
or U12964 (N_12964,N_9437,N_7681);
nor U12965 (N_12965,N_8096,N_5954);
nand U12966 (N_12966,N_5533,N_8788);
xor U12967 (N_12967,N_7104,N_5292);
nor U12968 (N_12968,N_6775,N_5564);
nor U12969 (N_12969,N_7710,N_7085);
nand U12970 (N_12970,N_6028,N_6543);
xnor U12971 (N_12971,N_7055,N_7180);
nand U12972 (N_12972,N_6348,N_7541);
xor U12973 (N_12973,N_5687,N_6201);
nor U12974 (N_12974,N_5240,N_8351);
nor U12975 (N_12975,N_7600,N_9128);
nand U12976 (N_12976,N_7330,N_9454);
or U12977 (N_12977,N_9300,N_8450);
or U12978 (N_12978,N_8208,N_7620);
or U12979 (N_12979,N_6148,N_9846);
or U12980 (N_12980,N_9853,N_5714);
and U12981 (N_12981,N_6250,N_6916);
and U12982 (N_12982,N_9560,N_7987);
and U12983 (N_12983,N_8322,N_7469);
or U12984 (N_12984,N_9276,N_7643);
or U12985 (N_12985,N_8302,N_6596);
nor U12986 (N_12986,N_5399,N_8773);
nor U12987 (N_12987,N_9503,N_5255);
or U12988 (N_12988,N_9423,N_6137);
xnor U12989 (N_12989,N_5273,N_7891);
nand U12990 (N_12990,N_7154,N_9122);
nor U12991 (N_12991,N_9948,N_7168);
xor U12992 (N_12992,N_9821,N_9198);
nand U12993 (N_12993,N_5756,N_7246);
xor U12994 (N_12994,N_7635,N_7447);
xnor U12995 (N_12995,N_7942,N_6454);
nor U12996 (N_12996,N_5191,N_9653);
or U12997 (N_12997,N_7344,N_5756);
nor U12998 (N_12998,N_8641,N_7112);
nand U12999 (N_12999,N_7005,N_7600);
or U13000 (N_13000,N_7305,N_6936);
nand U13001 (N_13001,N_7737,N_9872);
xor U13002 (N_13002,N_8375,N_6869);
nor U13003 (N_13003,N_8190,N_9756);
nor U13004 (N_13004,N_6211,N_8455);
or U13005 (N_13005,N_6849,N_7713);
and U13006 (N_13006,N_7949,N_6167);
or U13007 (N_13007,N_8677,N_6170);
nor U13008 (N_13008,N_6095,N_9890);
xor U13009 (N_13009,N_7401,N_5532);
xor U13010 (N_13010,N_7807,N_6212);
nand U13011 (N_13011,N_8018,N_5243);
nand U13012 (N_13012,N_8927,N_8505);
nor U13013 (N_13013,N_9492,N_8969);
or U13014 (N_13014,N_8417,N_7383);
nor U13015 (N_13015,N_9924,N_9514);
nor U13016 (N_13016,N_9456,N_6965);
and U13017 (N_13017,N_6028,N_5465);
nand U13018 (N_13018,N_8634,N_9588);
xnor U13019 (N_13019,N_9015,N_9957);
nand U13020 (N_13020,N_5339,N_7946);
and U13021 (N_13021,N_9303,N_5865);
nor U13022 (N_13022,N_8524,N_9023);
xnor U13023 (N_13023,N_8224,N_8006);
xnor U13024 (N_13024,N_7112,N_5220);
nor U13025 (N_13025,N_6039,N_7175);
nand U13026 (N_13026,N_5009,N_9185);
and U13027 (N_13027,N_6147,N_9324);
and U13028 (N_13028,N_6631,N_8073);
nor U13029 (N_13029,N_5512,N_9767);
nand U13030 (N_13030,N_9346,N_6690);
nand U13031 (N_13031,N_5823,N_6151);
xor U13032 (N_13032,N_7786,N_7674);
nor U13033 (N_13033,N_6186,N_6347);
or U13034 (N_13034,N_5422,N_5085);
nor U13035 (N_13035,N_5893,N_6350);
or U13036 (N_13036,N_8235,N_9407);
nor U13037 (N_13037,N_8942,N_6141);
or U13038 (N_13038,N_6486,N_7327);
and U13039 (N_13039,N_8616,N_7916);
and U13040 (N_13040,N_5042,N_6230);
nor U13041 (N_13041,N_7960,N_7442);
and U13042 (N_13042,N_6592,N_6811);
nor U13043 (N_13043,N_5687,N_6742);
xnor U13044 (N_13044,N_5190,N_7586);
and U13045 (N_13045,N_7087,N_5603);
nor U13046 (N_13046,N_9767,N_8541);
nor U13047 (N_13047,N_8203,N_9688);
and U13048 (N_13048,N_8565,N_5447);
xor U13049 (N_13049,N_5017,N_8457);
xnor U13050 (N_13050,N_8719,N_9635);
and U13051 (N_13051,N_7200,N_7604);
nand U13052 (N_13052,N_7343,N_6769);
xor U13053 (N_13053,N_6386,N_7980);
or U13054 (N_13054,N_8195,N_6489);
nand U13055 (N_13055,N_6196,N_8490);
xor U13056 (N_13056,N_9789,N_7735);
xor U13057 (N_13057,N_8551,N_6856);
or U13058 (N_13058,N_6961,N_5341);
or U13059 (N_13059,N_6957,N_7267);
or U13060 (N_13060,N_6369,N_6681);
nand U13061 (N_13061,N_9166,N_5099);
nand U13062 (N_13062,N_6395,N_6837);
nand U13063 (N_13063,N_7499,N_6600);
nand U13064 (N_13064,N_7030,N_7388);
nand U13065 (N_13065,N_5350,N_9458);
xnor U13066 (N_13066,N_6736,N_8815);
nand U13067 (N_13067,N_7418,N_7112);
nand U13068 (N_13068,N_7075,N_5029);
nor U13069 (N_13069,N_6768,N_5217);
nor U13070 (N_13070,N_8918,N_9344);
and U13071 (N_13071,N_8024,N_9548);
or U13072 (N_13072,N_6602,N_5483);
nor U13073 (N_13073,N_8985,N_5373);
xor U13074 (N_13074,N_9909,N_7604);
or U13075 (N_13075,N_9552,N_8518);
nor U13076 (N_13076,N_7650,N_6738);
nand U13077 (N_13077,N_5476,N_5138);
nand U13078 (N_13078,N_7588,N_9782);
xor U13079 (N_13079,N_8475,N_5960);
nand U13080 (N_13080,N_9088,N_6030);
xnor U13081 (N_13081,N_7860,N_5574);
nor U13082 (N_13082,N_6895,N_6565);
and U13083 (N_13083,N_8289,N_8575);
nand U13084 (N_13084,N_5530,N_9317);
nand U13085 (N_13085,N_7618,N_5665);
or U13086 (N_13086,N_9041,N_5705);
nor U13087 (N_13087,N_9185,N_8219);
or U13088 (N_13088,N_7942,N_5702);
or U13089 (N_13089,N_5600,N_7593);
nand U13090 (N_13090,N_5860,N_9895);
and U13091 (N_13091,N_8347,N_9269);
or U13092 (N_13092,N_8858,N_8472);
and U13093 (N_13093,N_6009,N_6137);
and U13094 (N_13094,N_6498,N_8205);
and U13095 (N_13095,N_8819,N_8570);
nand U13096 (N_13096,N_8831,N_5572);
and U13097 (N_13097,N_7088,N_5225);
nand U13098 (N_13098,N_9733,N_6794);
xor U13099 (N_13099,N_8667,N_7192);
and U13100 (N_13100,N_8942,N_6129);
or U13101 (N_13101,N_9183,N_5383);
and U13102 (N_13102,N_5202,N_9048);
xnor U13103 (N_13103,N_9607,N_5063);
nand U13104 (N_13104,N_5694,N_8566);
xor U13105 (N_13105,N_7509,N_6293);
or U13106 (N_13106,N_9581,N_9377);
or U13107 (N_13107,N_8850,N_6212);
or U13108 (N_13108,N_6959,N_8418);
nor U13109 (N_13109,N_6181,N_8757);
and U13110 (N_13110,N_9696,N_5088);
and U13111 (N_13111,N_7168,N_6990);
nand U13112 (N_13112,N_6299,N_5081);
and U13113 (N_13113,N_7446,N_6426);
or U13114 (N_13114,N_9953,N_8972);
and U13115 (N_13115,N_6419,N_7915);
and U13116 (N_13116,N_8662,N_7622);
or U13117 (N_13117,N_9784,N_8713);
nor U13118 (N_13118,N_6424,N_7878);
nand U13119 (N_13119,N_8612,N_8106);
xnor U13120 (N_13120,N_9229,N_6003);
xor U13121 (N_13121,N_7825,N_5522);
and U13122 (N_13122,N_5066,N_7529);
or U13123 (N_13123,N_9073,N_8572);
xnor U13124 (N_13124,N_9603,N_8669);
and U13125 (N_13125,N_9667,N_6456);
xnor U13126 (N_13126,N_7799,N_6088);
or U13127 (N_13127,N_8165,N_8883);
nor U13128 (N_13128,N_8981,N_5193);
nor U13129 (N_13129,N_9008,N_5877);
nand U13130 (N_13130,N_8703,N_6268);
and U13131 (N_13131,N_9710,N_6334);
xor U13132 (N_13132,N_6482,N_7276);
nand U13133 (N_13133,N_5806,N_6673);
nor U13134 (N_13134,N_6136,N_8788);
xnor U13135 (N_13135,N_5039,N_6673);
and U13136 (N_13136,N_7947,N_6170);
or U13137 (N_13137,N_9709,N_7093);
xnor U13138 (N_13138,N_9998,N_7812);
xnor U13139 (N_13139,N_7234,N_7806);
or U13140 (N_13140,N_7996,N_6689);
or U13141 (N_13141,N_5973,N_5775);
or U13142 (N_13142,N_8452,N_5967);
xnor U13143 (N_13143,N_8947,N_6248);
xnor U13144 (N_13144,N_8311,N_6841);
nor U13145 (N_13145,N_7392,N_6067);
and U13146 (N_13146,N_8972,N_6065);
nor U13147 (N_13147,N_8508,N_7486);
nand U13148 (N_13148,N_6917,N_8247);
xnor U13149 (N_13149,N_7643,N_6829);
or U13150 (N_13150,N_6197,N_9726);
or U13151 (N_13151,N_8802,N_9276);
or U13152 (N_13152,N_7731,N_9852);
xor U13153 (N_13153,N_8142,N_6841);
nand U13154 (N_13154,N_7790,N_6610);
and U13155 (N_13155,N_6710,N_6960);
and U13156 (N_13156,N_5963,N_5056);
or U13157 (N_13157,N_8441,N_8960);
or U13158 (N_13158,N_9712,N_8677);
or U13159 (N_13159,N_9257,N_6892);
nand U13160 (N_13160,N_6999,N_7569);
nand U13161 (N_13161,N_9481,N_7851);
or U13162 (N_13162,N_5595,N_5463);
xnor U13163 (N_13163,N_6292,N_7989);
xor U13164 (N_13164,N_6562,N_8983);
and U13165 (N_13165,N_9621,N_6139);
nand U13166 (N_13166,N_9397,N_9897);
or U13167 (N_13167,N_7345,N_8624);
xnor U13168 (N_13168,N_6738,N_9326);
xor U13169 (N_13169,N_6039,N_6961);
nand U13170 (N_13170,N_5514,N_9664);
and U13171 (N_13171,N_6781,N_5014);
and U13172 (N_13172,N_9217,N_7882);
and U13173 (N_13173,N_7785,N_9445);
and U13174 (N_13174,N_5504,N_7067);
nor U13175 (N_13175,N_9973,N_5630);
nand U13176 (N_13176,N_5476,N_7896);
xnor U13177 (N_13177,N_7577,N_5634);
or U13178 (N_13178,N_9118,N_8579);
xor U13179 (N_13179,N_5443,N_7217);
nand U13180 (N_13180,N_9944,N_5964);
or U13181 (N_13181,N_6144,N_6702);
and U13182 (N_13182,N_5107,N_9444);
nor U13183 (N_13183,N_6116,N_7258);
nor U13184 (N_13184,N_8620,N_7459);
xnor U13185 (N_13185,N_8802,N_8266);
and U13186 (N_13186,N_7320,N_8356);
nor U13187 (N_13187,N_8546,N_9476);
nor U13188 (N_13188,N_9502,N_9778);
xnor U13189 (N_13189,N_5712,N_5340);
nor U13190 (N_13190,N_5059,N_8479);
nor U13191 (N_13191,N_9909,N_5002);
nand U13192 (N_13192,N_9372,N_9879);
and U13193 (N_13193,N_9991,N_5386);
or U13194 (N_13194,N_8257,N_6112);
nor U13195 (N_13195,N_7999,N_8649);
nand U13196 (N_13196,N_5482,N_9194);
xnor U13197 (N_13197,N_9713,N_6236);
or U13198 (N_13198,N_8302,N_9133);
or U13199 (N_13199,N_8924,N_9547);
nand U13200 (N_13200,N_7283,N_8754);
nor U13201 (N_13201,N_7053,N_9211);
and U13202 (N_13202,N_5190,N_8935);
xor U13203 (N_13203,N_8951,N_7373);
nor U13204 (N_13204,N_5461,N_8670);
or U13205 (N_13205,N_7849,N_5936);
nor U13206 (N_13206,N_9249,N_8593);
nand U13207 (N_13207,N_8024,N_8837);
nand U13208 (N_13208,N_7350,N_5108);
nand U13209 (N_13209,N_5037,N_6400);
xor U13210 (N_13210,N_6668,N_8696);
xnor U13211 (N_13211,N_6334,N_8453);
xnor U13212 (N_13212,N_5701,N_6496);
or U13213 (N_13213,N_9737,N_7255);
or U13214 (N_13214,N_9834,N_7448);
xor U13215 (N_13215,N_7744,N_8752);
nor U13216 (N_13216,N_5446,N_6275);
nor U13217 (N_13217,N_5566,N_5494);
nand U13218 (N_13218,N_5329,N_7858);
or U13219 (N_13219,N_8711,N_5768);
nand U13220 (N_13220,N_6638,N_7529);
nand U13221 (N_13221,N_5239,N_6939);
and U13222 (N_13222,N_8206,N_7797);
or U13223 (N_13223,N_6578,N_6152);
nand U13224 (N_13224,N_8633,N_5318);
or U13225 (N_13225,N_6240,N_8626);
nor U13226 (N_13226,N_7795,N_8572);
nor U13227 (N_13227,N_7110,N_7141);
nor U13228 (N_13228,N_8588,N_7804);
nand U13229 (N_13229,N_7504,N_7399);
nor U13230 (N_13230,N_8856,N_7531);
and U13231 (N_13231,N_7775,N_9926);
nor U13232 (N_13232,N_5561,N_7615);
xor U13233 (N_13233,N_7246,N_6961);
and U13234 (N_13234,N_7264,N_8459);
and U13235 (N_13235,N_9322,N_6593);
nand U13236 (N_13236,N_9126,N_5502);
xnor U13237 (N_13237,N_9601,N_9378);
and U13238 (N_13238,N_9884,N_6015);
or U13239 (N_13239,N_9346,N_8691);
nor U13240 (N_13240,N_8774,N_6938);
and U13241 (N_13241,N_5371,N_7029);
nand U13242 (N_13242,N_6244,N_7877);
or U13243 (N_13243,N_5991,N_7862);
or U13244 (N_13244,N_6032,N_7085);
nor U13245 (N_13245,N_6298,N_6245);
xnor U13246 (N_13246,N_9573,N_9425);
and U13247 (N_13247,N_6326,N_7874);
nand U13248 (N_13248,N_8609,N_6157);
or U13249 (N_13249,N_8877,N_9089);
xnor U13250 (N_13250,N_9979,N_5515);
nand U13251 (N_13251,N_7268,N_6080);
nor U13252 (N_13252,N_6968,N_5550);
xnor U13253 (N_13253,N_5135,N_5344);
nand U13254 (N_13254,N_6355,N_5133);
nor U13255 (N_13255,N_9324,N_9852);
nor U13256 (N_13256,N_5694,N_9912);
xor U13257 (N_13257,N_8189,N_7892);
xor U13258 (N_13258,N_7478,N_8021);
nand U13259 (N_13259,N_6870,N_6406);
nor U13260 (N_13260,N_6154,N_9035);
xor U13261 (N_13261,N_8178,N_8200);
nand U13262 (N_13262,N_8298,N_6344);
nand U13263 (N_13263,N_6767,N_6037);
or U13264 (N_13264,N_7251,N_6763);
and U13265 (N_13265,N_9020,N_7494);
nor U13266 (N_13266,N_5072,N_9158);
and U13267 (N_13267,N_7129,N_5915);
nand U13268 (N_13268,N_5183,N_7601);
nor U13269 (N_13269,N_8647,N_7321);
nand U13270 (N_13270,N_6161,N_5890);
or U13271 (N_13271,N_7060,N_9827);
nand U13272 (N_13272,N_6746,N_6508);
or U13273 (N_13273,N_8409,N_9693);
nand U13274 (N_13274,N_9493,N_9281);
nor U13275 (N_13275,N_5639,N_8289);
xor U13276 (N_13276,N_6081,N_7534);
or U13277 (N_13277,N_9552,N_6441);
xor U13278 (N_13278,N_7598,N_5184);
xnor U13279 (N_13279,N_9180,N_9524);
nand U13280 (N_13280,N_5993,N_6760);
or U13281 (N_13281,N_6873,N_5907);
nand U13282 (N_13282,N_6799,N_8228);
nor U13283 (N_13283,N_6151,N_5179);
xor U13284 (N_13284,N_8614,N_6787);
or U13285 (N_13285,N_5882,N_6378);
xnor U13286 (N_13286,N_5755,N_8284);
nor U13287 (N_13287,N_9680,N_8513);
nand U13288 (N_13288,N_5561,N_7955);
nor U13289 (N_13289,N_7163,N_8929);
or U13290 (N_13290,N_5001,N_6614);
xnor U13291 (N_13291,N_8685,N_8712);
nand U13292 (N_13292,N_7655,N_6051);
or U13293 (N_13293,N_8278,N_7881);
or U13294 (N_13294,N_9195,N_5668);
nand U13295 (N_13295,N_9512,N_9253);
and U13296 (N_13296,N_7585,N_6021);
xnor U13297 (N_13297,N_7894,N_7280);
and U13298 (N_13298,N_9845,N_7682);
nand U13299 (N_13299,N_8013,N_7212);
nor U13300 (N_13300,N_7073,N_5010);
or U13301 (N_13301,N_9290,N_7919);
and U13302 (N_13302,N_5924,N_7256);
xnor U13303 (N_13303,N_6090,N_7984);
nand U13304 (N_13304,N_8043,N_7538);
or U13305 (N_13305,N_5050,N_8460);
or U13306 (N_13306,N_6479,N_6343);
nor U13307 (N_13307,N_9527,N_9822);
or U13308 (N_13308,N_7330,N_6849);
or U13309 (N_13309,N_7427,N_9868);
and U13310 (N_13310,N_8863,N_9697);
or U13311 (N_13311,N_6736,N_7424);
xnor U13312 (N_13312,N_8852,N_9594);
or U13313 (N_13313,N_6300,N_5739);
or U13314 (N_13314,N_5117,N_5566);
xor U13315 (N_13315,N_5317,N_9663);
or U13316 (N_13316,N_7580,N_6813);
nor U13317 (N_13317,N_5488,N_7740);
or U13318 (N_13318,N_7597,N_6642);
and U13319 (N_13319,N_6850,N_6986);
nor U13320 (N_13320,N_5390,N_8698);
xor U13321 (N_13321,N_9772,N_7264);
or U13322 (N_13322,N_7272,N_5659);
nor U13323 (N_13323,N_5684,N_8736);
nand U13324 (N_13324,N_5976,N_8922);
nand U13325 (N_13325,N_7882,N_7370);
and U13326 (N_13326,N_5059,N_9422);
xor U13327 (N_13327,N_5480,N_6116);
or U13328 (N_13328,N_8452,N_9555);
nand U13329 (N_13329,N_9266,N_5917);
xor U13330 (N_13330,N_5876,N_9270);
nand U13331 (N_13331,N_9716,N_6897);
or U13332 (N_13332,N_5730,N_9005);
or U13333 (N_13333,N_8329,N_9378);
or U13334 (N_13334,N_9414,N_8695);
nand U13335 (N_13335,N_5836,N_9495);
nand U13336 (N_13336,N_6149,N_7356);
and U13337 (N_13337,N_9535,N_9183);
xnor U13338 (N_13338,N_6971,N_5189);
nor U13339 (N_13339,N_5003,N_6571);
xor U13340 (N_13340,N_8007,N_9631);
or U13341 (N_13341,N_9010,N_8733);
nor U13342 (N_13342,N_7382,N_7103);
or U13343 (N_13343,N_9694,N_6174);
or U13344 (N_13344,N_6974,N_7701);
and U13345 (N_13345,N_6234,N_7687);
xor U13346 (N_13346,N_6380,N_5340);
nor U13347 (N_13347,N_8377,N_7205);
and U13348 (N_13348,N_6137,N_7395);
or U13349 (N_13349,N_9255,N_7800);
nand U13350 (N_13350,N_5419,N_6701);
nand U13351 (N_13351,N_6940,N_6432);
nor U13352 (N_13352,N_9039,N_5953);
and U13353 (N_13353,N_5644,N_9985);
xnor U13354 (N_13354,N_5204,N_6403);
nand U13355 (N_13355,N_8201,N_7627);
or U13356 (N_13356,N_8077,N_9353);
nand U13357 (N_13357,N_8952,N_6769);
or U13358 (N_13358,N_9812,N_6563);
nor U13359 (N_13359,N_9170,N_9834);
nor U13360 (N_13360,N_6249,N_9864);
or U13361 (N_13361,N_8243,N_9219);
or U13362 (N_13362,N_5701,N_8716);
nor U13363 (N_13363,N_5802,N_5867);
and U13364 (N_13364,N_5053,N_8649);
and U13365 (N_13365,N_8151,N_9091);
xnor U13366 (N_13366,N_9751,N_5124);
xor U13367 (N_13367,N_7341,N_6071);
nor U13368 (N_13368,N_7854,N_8452);
nand U13369 (N_13369,N_8965,N_8006);
nor U13370 (N_13370,N_7683,N_5065);
nor U13371 (N_13371,N_6585,N_9602);
nor U13372 (N_13372,N_9316,N_6933);
and U13373 (N_13373,N_6329,N_5770);
or U13374 (N_13374,N_5142,N_6960);
and U13375 (N_13375,N_6400,N_7227);
or U13376 (N_13376,N_5144,N_8102);
nand U13377 (N_13377,N_8993,N_7547);
and U13378 (N_13378,N_8288,N_5048);
and U13379 (N_13379,N_7043,N_7072);
or U13380 (N_13380,N_5679,N_8870);
or U13381 (N_13381,N_7310,N_8456);
xnor U13382 (N_13382,N_9913,N_5390);
xor U13383 (N_13383,N_9681,N_8899);
nor U13384 (N_13384,N_5134,N_8824);
xnor U13385 (N_13385,N_8874,N_5207);
or U13386 (N_13386,N_5684,N_5512);
nand U13387 (N_13387,N_9532,N_8228);
and U13388 (N_13388,N_6464,N_8435);
nand U13389 (N_13389,N_7936,N_5673);
or U13390 (N_13390,N_9190,N_5958);
xor U13391 (N_13391,N_8372,N_7840);
nand U13392 (N_13392,N_8668,N_7662);
or U13393 (N_13393,N_9586,N_6380);
nor U13394 (N_13394,N_8325,N_5056);
nor U13395 (N_13395,N_5018,N_9193);
and U13396 (N_13396,N_5743,N_9331);
nor U13397 (N_13397,N_6145,N_9917);
xor U13398 (N_13398,N_5492,N_8113);
xor U13399 (N_13399,N_9883,N_7774);
and U13400 (N_13400,N_9758,N_5949);
xor U13401 (N_13401,N_9284,N_6973);
and U13402 (N_13402,N_9027,N_9316);
and U13403 (N_13403,N_8769,N_8996);
or U13404 (N_13404,N_8556,N_6083);
xor U13405 (N_13405,N_9755,N_5793);
nand U13406 (N_13406,N_7987,N_6773);
xnor U13407 (N_13407,N_6903,N_9901);
or U13408 (N_13408,N_6738,N_5981);
or U13409 (N_13409,N_5695,N_7864);
or U13410 (N_13410,N_9785,N_8400);
xor U13411 (N_13411,N_5210,N_7212);
xor U13412 (N_13412,N_7318,N_5564);
xor U13413 (N_13413,N_5616,N_8815);
nand U13414 (N_13414,N_5035,N_9015);
and U13415 (N_13415,N_7846,N_5176);
or U13416 (N_13416,N_6848,N_7639);
nand U13417 (N_13417,N_8308,N_6715);
nand U13418 (N_13418,N_7901,N_7163);
nand U13419 (N_13419,N_9097,N_7307);
nor U13420 (N_13420,N_5825,N_9353);
xnor U13421 (N_13421,N_7612,N_8504);
or U13422 (N_13422,N_6665,N_6296);
or U13423 (N_13423,N_7443,N_6476);
xor U13424 (N_13424,N_6357,N_6874);
or U13425 (N_13425,N_6433,N_8270);
xor U13426 (N_13426,N_9162,N_8681);
xnor U13427 (N_13427,N_9268,N_6956);
nand U13428 (N_13428,N_8445,N_5351);
or U13429 (N_13429,N_6047,N_7389);
nand U13430 (N_13430,N_7064,N_6955);
or U13431 (N_13431,N_8604,N_7821);
and U13432 (N_13432,N_8792,N_7883);
and U13433 (N_13433,N_7955,N_5076);
nand U13434 (N_13434,N_7643,N_9585);
and U13435 (N_13435,N_7918,N_6547);
nor U13436 (N_13436,N_5742,N_8497);
or U13437 (N_13437,N_8066,N_8221);
nand U13438 (N_13438,N_6463,N_9171);
or U13439 (N_13439,N_8823,N_8482);
xor U13440 (N_13440,N_6488,N_5304);
nor U13441 (N_13441,N_7143,N_9304);
and U13442 (N_13442,N_6412,N_6187);
and U13443 (N_13443,N_5083,N_6533);
or U13444 (N_13444,N_5507,N_6098);
xnor U13445 (N_13445,N_8242,N_8522);
xor U13446 (N_13446,N_7899,N_7530);
nand U13447 (N_13447,N_6134,N_5855);
xnor U13448 (N_13448,N_9428,N_9670);
and U13449 (N_13449,N_5882,N_9428);
xnor U13450 (N_13450,N_7691,N_7424);
or U13451 (N_13451,N_7483,N_9343);
nor U13452 (N_13452,N_6250,N_8286);
and U13453 (N_13453,N_7490,N_7086);
nand U13454 (N_13454,N_5305,N_7052);
nand U13455 (N_13455,N_8351,N_7459);
xnor U13456 (N_13456,N_5174,N_5381);
nor U13457 (N_13457,N_8051,N_8013);
and U13458 (N_13458,N_7172,N_5781);
or U13459 (N_13459,N_6388,N_8132);
xor U13460 (N_13460,N_6919,N_9896);
and U13461 (N_13461,N_6939,N_7160);
and U13462 (N_13462,N_8167,N_8402);
nor U13463 (N_13463,N_7714,N_6695);
nand U13464 (N_13464,N_5467,N_7165);
or U13465 (N_13465,N_7519,N_9132);
nand U13466 (N_13466,N_5952,N_7021);
and U13467 (N_13467,N_8532,N_9499);
or U13468 (N_13468,N_6098,N_7550);
and U13469 (N_13469,N_8651,N_8879);
nand U13470 (N_13470,N_8700,N_5422);
xnor U13471 (N_13471,N_9565,N_8943);
nand U13472 (N_13472,N_9051,N_5791);
xor U13473 (N_13473,N_5718,N_8315);
nor U13474 (N_13474,N_8659,N_7139);
xnor U13475 (N_13475,N_9098,N_8919);
and U13476 (N_13476,N_5941,N_9831);
nand U13477 (N_13477,N_8081,N_8235);
xnor U13478 (N_13478,N_6485,N_7276);
and U13479 (N_13479,N_5475,N_6648);
nand U13480 (N_13480,N_7329,N_7095);
or U13481 (N_13481,N_6954,N_8538);
or U13482 (N_13482,N_7454,N_8512);
and U13483 (N_13483,N_8607,N_7555);
nor U13484 (N_13484,N_7943,N_8216);
xor U13485 (N_13485,N_5231,N_8801);
and U13486 (N_13486,N_8126,N_5701);
nand U13487 (N_13487,N_5939,N_7014);
xor U13488 (N_13488,N_7263,N_7518);
and U13489 (N_13489,N_7638,N_6559);
xor U13490 (N_13490,N_9400,N_9003);
or U13491 (N_13491,N_5998,N_6778);
and U13492 (N_13492,N_6129,N_9184);
or U13493 (N_13493,N_5479,N_8485);
and U13494 (N_13494,N_8235,N_8445);
xnor U13495 (N_13495,N_6488,N_8222);
xor U13496 (N_13496,N_5225,N_8297);
nand U13497 (N_13497,N_6843,N_9425);
xnor U13498 (N_13498,N_6114,N_7981);
nor U13499 (N_13499,N_8544,N_6870);
nand U13500 (N_13500,N_7932,N_5349);
nor U13501 (N_13501,N_5308,N_8365);
nor U13502 (N_13502,N_7812,N_8649);
xor U13503 (N_13503,N_5240,N_8187);
and U13504 (N_13504,N_7823,N_9072);
nor U13505 (N_13505,N_6694,N_8296);
or U13506 (N_13506,N_6019,N_8642);
nand U13507 (N_13507,N_9799,N_8901);
nor U13508 (N_13508,N_7169,N_7253);
nand U13509 (N_13509,N_6565,N_5043);
and U13510 (N_13510,N_8221,N_5288);
nor U13511 (N_13511,N_7209,N_6981);
nand U13512 (N_13512,N_5758,N_7752);
xor U13513 (N_13513,N_7303,N_7689);
xnor U13514 (N_13514,N_6402,N_6414);
nand U13515 (N_13515,N_7955,N_6028);
xor U13516 (N_13516,N_8284,N_7411);
nor U13517 (N_13517,N_7487,N_9723);
and U13518 (N_13518,N_9126,N_7904);
xor U13519 (N_13519,N_8896,N_6846);
xor U13520 (N_13520,N_6780,N_9589);
nor U13521 (N_13521,N_6582,N_8177);
nor U13522 (N_13522,N_7748,N_7611);
nor U13523 (N_13523,N_5448,N_8909);
nand U13524 (N_13524,N_5462,N_5076);
nor U13525 (N_13525,N_9004,N_7089);
nor U13526 (N_13526,N_7837,N_7218);
and U13527 (N_13527,N_5131,N_5652);
or U13528 (N_13528,N_5158,N_9900);
nor U13529 (N_13529,N_9331,N_5780);
and U13530 (N_13530,N_6593,N_5720);
and U13531 (N_13531,N_9724,N_9630);
nor U13532 (N_13532,N_5963,N_5475);
nand U13533 (N_13533,N_5491,N_9771);
or U13534 (N_13534,N_8002,N_6346);
nand U13535 (N_13535,N_5627,N_6780);
xnor U13536 (N_13536,N_9387,N_8817);
or U13537 (N_13537,N_7899,N_7453);
nand U13538 (N_13538,N_9515,N_7704);
or U13539 (N_13539,N_5441,N_5007);
and U13540 (N_13540,N_9329,N_7926);
and U13541 (N_13541,N_8020,N_5708);
and U13542 (N_13542,N_7475,N_7830);
nand U13543 (N_13543,N_7025,N_8150);
or U13544 (N_13544,N_9062,N_7656);
or U13545 (N_13545,N_9182,N_5186);
nor U13546 (N_13546,N_8990,N_7784);
xor U13547 (N_13547,N_5390,N_9782);
nor U13548 (N_13548,N_5986,N_7329);
and U13549 (N_13549,N_7724,N_6284);
xnor U13550 (N_13550,N_9381,N_7522);
nand U13551 (N_13551,N_7899,N_7874);
nor U13552 (N_13552,N_8320,N_9319);
and U13553 (N_13553,N_6295,N_8679);
and U13554 (N_13554,N_9989,N_7003);
and U13555 (N_13555,N_6593,N_6213);
and U13556 (N_13556,N_6059,N_5725);
or U13557 (N_13557,N_8958,N_9890);
or U13558 (N_13558,N_5811,N_5112);
or U13559 (N_13559,N_8874,N_9737);
nor U13560 (N_13560,N_8209,N_9985);
nand U13561 (N_13561,N_5782,N_7263);
and U13562 (N_13562,N_6305,N_8811);
and U13563 (N_13563,N_7859,N_5959);
nor U13564 (N_13564,N_6405,N_7895);
nor U13565 (N_13565,N_9524,N_8535);
or U13566 (N_13566,N_6951,N_6776);
xor U13567 (N_13567,N_9301,N_9115);
nor U13568 (N_13568,N_9936,N_7650);
xor U13569 (N_13569,N_5203,N_6736);
nor U13570 (N_13570,N_5274,N_6471);
nor U13571 (N_13571,N_7192,N_9309);
or U13572 (N_13572,N_9673,N_8637);
nand U13573 (N_13573,N_5567,N_5261);
nor U13574 (N_13574,N_8334,N_8920);
or U13575 (N_13575,N_7468,N_6024);
xor U13576 (N_13576,N_5587,N_9768);
or U13577 (N_13577,N_5935,N_9606);
or U13578 (N_13578,N_5937,N_9868);
nor U13579 (N_13579,N_7966,N_9742);
or U13580 (N_13580,N_5479,N_9509);
and U13581 (N_13581,N_6848,N_5720);
or U13582 (N_13582,N_8332,N_8158);
nor U13583 (N_13583,N_5058,N_6072);
and U13584 (N_13584,N_8325,N_5352);
nor U13585 (N_13585,N_5687,N_9319);
or U13586 (N_13586,N_6152,N_9876);
nor U13587 (N_13587,N_7826,N_7709);
xor U13588 (N_13588,N_6952,N_6840);
and U13589 (N_13589,N_9267,N_9411);
nand U13590 (N_13590,N_6162,N_6303);
nand U13591 (N_13591,N_7752,N_7579);
nand U13592 (N_13592,N_7908,N_9003);
nor U13593 (N_13593,N_5451,N_9002);
and U13594 (N_13594,N_6580,N_9202);
xor U13595 (N_13595,N_9210,N_9141);
and U13596 (N_13596,N_6879,N_6674);
nand U13597 (N_13597,N_9887,N_9830);
nand U13598 (N_13598,N_6010,N_9828);
nand U13599 (N_13599,N_6254,N_8385);
or U13600 (N_13600,N_8821,N_7679);
and U13601 (N_13601,N_5034,N_8770);
or U13602 (N_13602,N_6691,N_7989);
or U13603 (N_13603,N_6908,N_7097);
nor U13604 (N_13604,N_9968,N_5696);
nand U13605 (N_13605,N_8980,N_9298);
nor U13606 (N_13606,N_7562,N_6920);
nand U13607 (N_13607,N_9106,N_6084);
xnor U13608 (N_13608,N_6863,N_6837);
and U13609 (N_13609,N_6829,N_6146);
nand U13610 (N_13610,N_6304,N_5326);
or U13611 (N_13611,N_6192,N_9415);
nand U13612 (N_13612,N_5520,N_6981);
or U13613 (N_13613,N_8443,N_9920);
nand U13614 (N_13614,N_5825,N_6183);
xnor U13615 (N_13615,N_7934,N_9679);
nor U13616 (N_13616,N_9972,N_7083);
or U13617 (N_13617,N_7578,N_7300);
and U13618 (N_13618,N_5270,N_9427);
xor U13619 (N_13619,N_7179,N_8366);
nor U13620 (N_13620,N_9380,N_9564);
xor U13621 (N_13621,N_7131,N_5661);
xor U13622 (N_13622,N_5741,N_6733);
and U13623 (N_13623,N_7787,N_9403);
or U13624 (N_13624,N_5071,N_8700);
nand U13625 (N_13625,N_5820,N_5208);
or U13626 (N_13626,N_6009,N_9377);
nor U13627 (N_13627,N_7119,N_5119);
and U13628 (N_13628,N_5365,N_8529);
or U13629 (N_13629,N_5100,N_7783);
and U13630 (N_13630,N_5049,N_7300);
xor U13631 (N_13631,N_5927,N_7443);
nand U13632 (N_13632,N_6028,N_7961);
nor U13633 (N_13633,N_9599,N_8077);
nand U13634 (N_13634,N_9901,N_8287);
nand U13635 (N_13635,N_9662,N_9265);
or U13636 (N_13636,N_7271,N_9009);
xnor U13637 (N_13637,N_7161,N_5312);
xor U13638 (N_13638,N_6861,N_5198);
xor U13639 (N_13639,N_9847,N_8047);
nand U13640 (N_13640,N_7480,N_7189);
nor U13641 (N_13641,N_5911,N_6775);
or U13642 (N_13642,N_5229,N_8041);
nor U13643 (N_13643,N_5565,N_6545);
nand U13644 (N_13644,N_6917,N_8238);
nor U13645 (N_13645,N_5411,N_9247);
xor U13646 (N_13646,N_8426,N_7709);
nand U13647 (N_13647,N_8546,N_5265);
nand U13648 (N_13648,N_5637,N_6441);
nor U13649 (N_13649,N_9280,N_9598);
xor U13650 (N_13650,N_5665,N_7897);
nand U13651 (N_13651,N_7071,N_7092);
nor U13652 (N_13652,N_9735,N_8708);
and U13653 (N_13653,N_7923,N_5260);
xor U13654 (N_13654,N_5676,N_6561);
and U13655 (N_13655,N_6922,N_6219);
and U13656 (N_13656,N_9564,N_8407);
xor U13657 (N_13657,N_6313,N_6837);
nand U13658 (N_13658,N_5060,N_9413);
nand U13659 (N_13659,N_7978,N_9978);
nor U13660 (N_13660,N_9332,N_7857);
xor U13661 (N_13661,N_6354,N_5800);
xor U13662 (N_13662,N_5052,N_6640);
nor U13663 (N_13663,N_6897,N_9819);
xnor U13664 (N_13664,N_5857,N_7225);
or U13665 (N_13665,N_8287,N_8266);
nand U13666 (N_13666,N_7279,N_8980);
nor U13667 (N_13667,N_9974,N_6924);
xnor U13668 (N_13668,N_6896,N_8310);
nor U13669 (N_13669,N_8113,N_6942);
nand U13670 (N_13670,N_8988,N_6247);
xnor U13671 (N_13671,N_9522,N_8870);
nor U13672 (N_13672,N_8895,N_5482);
nand U13673 (N_13673,N_5611,N_6292);
or U13674 (N_13674,N_6258,N_6920);
nand U13675 (N_13675,N_6078,N_5941);
and U13676 (N_13676,N_5131,N_9983);
nand U13677 (N_13677,N_8061,N_8976);
or U13678 (N_13678,N_8563,N_6221);
and U13679 (N_13679,N_8810,N_8219);
or U13680 (N_13680,N_7476,N_8998);
nand U13681 (N_13681,N_9703,N_5985);
nand U13682 (N_13682,N_6837,N_6252);
nor U13683 (N_13683,N_7096,N_8094);
nor U13684 (N_13684,N_9890,N_7030);
or U13685 (N_13685,N_8082,N_8623);
and U13686 (N_13686,N_8578,N_5413);
or U13687 (N_13687,N_5544,N_8104);
nand U13688 (N_13688,N_8715,N_9923);
and U13689 (N_13689,N_5159,N_8614);
and U13690 (N_13690,N_6931,N_9779);
or U13691 (N_13691,N_6463,N_8866);
xnor U13692 (N_13692,N_5036,N_9188);
or U13693 (N_13693,N_7560,N_7309);
xnor U13694 (N_13694,N_8267,N_7373);
and U13695 (N_13695,N_6658,N_7305);
or U13696 (N_13696,N_9487,N_7220);
nand U13697 (N_13697,N_5356,N_8193);
xor U13698 (N_13698,N_7716,N_7650);
nor U13699 (N_13699,N_7505,N_5825);
or U13700 (N_13700,N_8356,N_6073);
or U13701 (N_13701,N_9792,N_7243);
and U13702 (N_13702,N_6074,N_8741);
nand U13703 (N_13703,N_7897,N_9000);
nor U13704 (N_13704,N_8539,N_9526);
or U13705 (N_13705,N_6651,N_7224);
nand U13706 (N_13706,N_8605,N_6625);
xnor U13707 (N_13707,N_8262,N_7827);
xor U13708 (N_13708,N_8667,N_7548);
nor U13709 (N_13709,N_5355,N_7041);
nand U13710 (N_13710,N_8054,N_6045);
nand U13711 (N_13711,N_8860,N_7869);
nor U13712 (N_13712,N_9099,N_7456);
and U13713 (N_13713,N_7690,N_6367);
and U13714 (N_13714,N_7426,N_9487);
and U13715 (N_13715,N_7503,N_5478);
or U13716 (N_13716,N_8032,N_9640);
xor U13717 (N_13717,N_8917,N_5522);
xor U13718 (N_13718,N_8208,N_6241);
or U13719 (N_13719,N_9031,N_9496);
xnor U13720 (N_13720,N_7930,N_9698);
or U13721 (N_13721,N_7789,N_5708);
and U13722 (N_13722,N_8873,N_7558);
xnor U13723 (N_13723,N_5608,N_7938);
and U13724 (N_13724,N_5082,N_5432);
xor U13725 (N_13725,N_7483,N_6186);
and U13726 (N_13726,N_9036,N_8116);
nor U13727 (N_13727,N_7979,N_7128);
xnor U13728 (N_13728,N_8696,N_6154);
xor U13729 (N_13729,N_6227,N_5010);
nor U13730 (N_13730,N_7202,N_6842);
nand U13731 (N_13731,N_6196,N_7547);
nand U13732 (N_13732,N_7378,N_8164);
xnor U13733 (N_13733,N_6433,N_9569);
xor U13734 (N_13734,N_9986,N_9778);
or U13735 (N_13735,N_9061,N_8623);
xor U13736 (N_13736,N_9726,N_7412);
nor U13737 (N_13737,N_8124,N_5214);
nand U13738 (N_13738,N_6740,N_9206);
and U13739 (N_13739,N_8034,N_7189);
or U13740 (N_13740,N_7423,N_5363);
nor U13741 (N_13741,N_8787,N_5367);
or U13742 (N_13742,N_6198,N_7744);
or U13743 (N_13743,N_9748,N_8528);
xor U13744 (N_13744,N_7859,N_9756);
and U13745 (N_13745,N_8238,N_9935);
nor U13746 (N_13746,N_8136,N_9793);
and U13747 (N_13747,N_7268,N_8072);
nand U13748 (N_13748,N_5051,N_6023);
nor U13749 (N_13749,N_5467,N_5916);
or U13750 (N_13750,N_5658,N_7354);
or U13751 (N_13751,N_8824,N_7538);
nor U13752 (N_13752,N_7732,N_6420);
and U13753 (N_13753,N_6576,N_9831);
or U13754 (N_13754,N_6408,N_6821);
nand U13755 (N_13755,N_8616,N_7585);
or U13756 (N_13756,N_9644,N_9234);
nor U13757 (N_13757,N_8055,N_6612);
nor U13758 (N_13758,N_9558,N_5550);
xnor U13759 (N_13759,N_5202,N_9455);
and U13760 (N_13760,N_7235,N_8385);
nand U13761 (N_13761,N_6828,N_5656);
nand U13762 (N_13762,N_5704,N_7553);
and U13763 (N_13763,N_7189,N_9370);
nor U13764 (N_13764,N_7784,N_7932);
nor U13765 (N_13765,N_9099,N_6586);
and U13766 (N_13766,N_6251,N_7108);
xor U13767 (N_13767,N_8931,N_7482);
or U13768 (N_13768,N_7367,N_5119);
nand U13769 (N_13769,N_5225,N_8549);
or U13770 (N_13770,N_6741,N_6427);
nand U13771 (N_13771,N_8050,N_9962);
nor U13772 (N_13772,N_5745,N_9830);
xnor U13773 (N_13773,N_8228,N_6540);
xor U13774 (N_13774,N_7357,N_9649);
and U13775 (N_13775,N_5510,N_7898);
nor U13776 (N_13776,N_7781,N_8046);
nor U13777 (N_13777,N_7646,N_7369);
or U13778 (N_13778,N_8397,N_7061);
and U13779 (N_13779,N_6823,N_9908);
xnor U13780 (N_13780,N_7115,N_7497);
xor U13781 (N_13781,N_9225,N_8656);
xnor U13782 (N_13782,N_7810,N_6057);
or U13783 (N_13783,N_7857,N_8670);
xor U13784 (N_13784,N_9212,N_5289);
or U13785 (N_13785,N_9449,N_5572);
nor U13786 (N_13786,N_5955,N_9977);
and U13787 (N_13787,N_7471,N_8243);
nor U13788 (N_13788,N_5622,N_5077);
or U13789 (N_13789,N_8567,N_8696);
nand U13790 (N_13790,N_9509,N_8983);
nand U13791 (N_13791,N_9540,N_6972);
or U13792 (N_13792,N_8862,N_9870);
or U13793 (N_13793,N_7735,N_8181);
nor U13794 (N_13794,N_5654,N_9020);
or U13795 (N_13795,N_7476,N_7761);
nand U13796 (N_13796,N_6902,N_6997);
xor U13797 (N_13797,N_6265,N_8339);
xnor U13798 (N_13798,N_5461,N_6465);
and U13799 (N_13799,N_9640,N_8252);
and U13800 (N_13800,N_6072,N_9325);
nor U13801 (N_13801,N_8501,N_9322);
nor U13802 (N_13802,N_7136,N_5308);
nor U13803 (N_13803,N_7710,N_9612);
nor U13804 (N_13804,N_8094,N_5591);
nand U13805 (N_13805,N_5556,N_8816);
and U13806 (N_13806,N_5273,N_7592);
nand U13807 (N_13807,N_8662,N_7120);
nor U13808 (N_13808,N_5267,N_6404);
nor U13809 (N_13809,N_6325,N_9121);
or U13810 (N_13810,N_9220,N_8979);
and U13811 (N_13811,N_5547,N_9063);
and U13812 (N_13812,N_5258,N_8528);
and U13813 (N_13813,N_6272,N_6752);
xor U13814 (N_13814,N_8295,N_7302);
nand U13815 (N_13815,N_9326,N_6199);
xnor U13816 (N_13816,N_7479,N_7808);
or U13817 (N_13817,N_6976,N_9700);
nor U13818 (N_13818,N_5118,N_5588);
xnor U13819 (N_13819,N_7168,N_9178);
or U13820 (N_13820,N_9700,N_6482);
nor U13821 (N_13821,N_6765,N_6245);
or U13822 (N_13822,N_9277,N_8971);
xnor U13823 (N_13823,N_6149,N_6013);
nand U13824 (N_13824,N_5704,N_9373);
nor U13825 (N_13825,N_8877,N_6408);
nand U13826 (N_13826,N_9391,N_6671);
nand U13827 (N_13827,N_7225,N_8877);
nand U13828 (N_13828,N_5544,N_6809);
xnor U13829 (N_13829,N_6465,N_7946);
or U13830 (N_13830,N_9501,N_5532);
and U13831 (N_13831,N_7720,N_9535);
nand U13832 (N_13832,N_8489,N_7739);
xor U13833 (N_13833,N_9472,N_8867);
nor U13834 (N_13834,N_5360,N_7859);
xnor U13835 (N_13835,N_5793,N_7137);
nand U13836 (N_13836,N_5973,N_8701);
nand U13837 (N_13837,N_6601,N_8433);
xor U13838 (N_13838,N_9061,N_7731);
nand U13839 (N_13839,N_6804,N_6898);
xnor U13840 (N_13840,N_8211,N_9699);
nor U13841 (N_13841,N_8169,N_8068);
and U13842 (N_13842,N_6750,N_6293);
xor U13843 (N_13843,N_8714,N_5424);
xor U13844 (N_13844,N_5477,N_7338);
xnor U13845 (N_13845,N_9277,N_5964);
and U13846 (N_13846,N_8592,N_7758);
xor U13847 (N_13847,N_8310,N_8096);
nor U13848 (N_13848,N_7454,N_9165);
or U13849 (N_13849,N_9313,N_8780);
or U13850 (N_13850,N_8283,N_7992);
or U13851 (N_13851,N_5866,N_8461);
xor U13852 (N_13852,N_5713,N_9304);
or U13853 (N_13853,N_8850,N_7521);
nor U13854 (N_13854,N_6611,N_9641);
nand U13855 (N_13855,N_5244,N_9003);
nor U13856 (N_13856,N_8033,N_5003);
or U13857 (N_13857,N_7536,N_6614);
and U13858 (N_13858,N_6529,N_9814);
or U13859 (N_13859,N_7011,N_8770);
nand U13860 (N_13860,N_6703,N_7966);
xnor U13861 (N_13861,N_6950,N_8991);
nand U13862 (N_13862,N_7706,N_9708);
nand U13863 (N_13863,N_7020,N_5217);
xnor U13864 (N_13864,N_9807,N_6568);
nor U13865 (N_13865,N_8576,N_9547);
nor U13866 (N_13866,N_5146,N_8492);
nor U13867 (N_13867,N_8975,N_9814);
xnor U13868 (N_13868,N_7910,N_8837);
nor U13869 (N_13869,N_7760,N_9839);
and U13870 (N_13870,N_9895,N_7713);
nor U13871 (N_13871,N_5855,N_7120);
nand U13872 (N_13872,N_6879,N_6440);
or U13873 (N_13873,N_9271,N_9314);
and U13874 (N_13874,N_5841,N_9979);
or U13875 (N_13875,N_5246,N_7833);
nand U13876 (N_13876,N_5362,N_7369);
xor U13877 (N_13877,N_7733,N_9995);
nand U13878 (N_13878,N_6728,N_6855);
and U13879 (N_13879,N_8178,N_7764);
xnor U13880 (N_13880,N_8808,N_6101);
or U13881 (N_13881,N_8506,N_9652);
nor U13882 (N_13882,N_5935,N_7177);
or U13883 (N_13883,N_7117,N_6220);
nor U13884 (N_13884,N_8011,N_8559);
and U13885 (N_13885,N_9894,N_8318);
and U13886 (N_13886,N_5951,N_7371);
and U13887 (N_13887,N_5565,N_5869);
and U13888 (N_13888,N_5180,N_8668);
or U13889 (N_13889,N_9691,N_6067);
or U13890 (N_13890,N_8247,N_5006);
and U13891 (N_13891,N_6445,N_7123);
xnor U13892 (N_13892,N_9670,N_6084);
xnor U13893 (N_13893,N_7458,N_6398);
xor U13894 (N_13894,N_9378,N_7411);
or U13895 (N_13895,N_5302,N_9375);
and U13896 (N_13896,N_5779,N_8666);
nor U13897 (N_13897,N_7602,N_9069);
nor U13898 (N_13898,N_8489,N_8459);
and U13899 (N_13899,N_9167,N_9510);
and U13900 (N_13900,N_9760,N_7441);
or U13901 (N_13901,N_8275,N_6223);
nand U13902 (N_13902,N_7648,N_8892);
and U13903 (N_13903,N_8278,N_9879);
xnor U13904 (N_13904,N_8774,N_7925);
nand U13905 (N_13905,N_5787,N_7339);
or U13906 (N_13906,N_5999,N_7012);
xor U13907 (N_13907,N_7007,N_6069);
nand U13908 (N_13908,N_7978,N_9519);
and U13909 (N_13909,N_8676,N_5313);
and U13910 (N_13910,N_9936,N_6197);
or U13911 (N_13911,N_9789,N_9136);
nor U13912 (N_13912,N_6526,N_8678);
nor U13913 (N_13913,N_6689,N_8635);
xor U13914 (N_13914,N_9155,N_6889);
nor U13915 (N_13915,N_5617,N_9845);
nor U13916 (N_13916,N_6912,N_5987);
xnor U13917 (N_13917,N_6645,N_9467);
or U13918 (N_13918,N_7022,N_7726);
and U13919 (N_13919,N_6242,N_7408);
nor U13920 (N_13920,N_8094,N_8330);
nor U13921 (N_13921,N_6416,N_8210);
nand U13922 (N_13922,N_6163,N_6463);
nand U13923 (N_13923,N_9866,N_7539);
xnor U13924 (N_13924,N_7396,N_8922);
nor U13925 (N_13925,N_9329,N_7212);
nand U13926 (N_13926,N_5283,N_9550);
and U13927 (N_13927,N_6489,N_8921);
and U13928 (N_13928,N_5450,N_5957);
or U13929 (N_13929,N_5936,N_8224);
and U13930 (N_13930,N_6463,N_5433);
nand U13931 (N_13931,N_5285,N_7265);
nand U13932 (N_13932,N_9371,N_7275);
and U13933 (N_13933,N_7966,N_8376);
and U13934 (N_13934,N_8281,N_6218);
and U13935 (N_13935,N_7516,N_8987);
or U13936 (N_13936,N_6029,N_6771);
and U13937 (N_13937,N_5798,N_9887);
nand U13938 (N_13938,N_6618,N_6327);
or U13939 (N_13939,N_8880,N_6851);
or U13940 (N_13940,N_5091,N_6108);
and U13941 (N_13941,N_9084,N_8570);
and U13942 (N_13942,N_8705,N_9669);
or U13943 (N_13943,N_6757,N_9460);
nor U13944 (N_13944,N_5788,N_6501);
nor U13945 (N_13945,N_7910,N_9071);
and U13946 (N_13946,N_9953,N_5894);
or U13947 (N_13947,N_9734,N_8589);
or U13948 (N_13948,N_6402,N_8187);
and U13949 (N_13949,N_8173,N_6496);
nand U13950 (N_13950,N_9448,N_8038);
and U13951 (N_13951,N_7659,N_9848);
nand U13952 (N_13952,N_5039,N_9651);
nor U13953 (N_13953,N_7405,N_9042);
and U13954 (N_13954,N_7253,N_6712);
or U13955 (N_13955,N_5943,N_5421);
and U13956 (N_13956,N_6503,N_6274);
nand U13957 (N_13957,N_5366,N_9361);
nand U13958 (N_13958,N_6346,N_7163);
nor U13959 (N_13959,N_7440,N_7909);
or U13960 (N_13960,N_5420,N_9669);
nand U13961 (N_13961,N_5091,N_5556);
nand U13962 (N_13962,N_8743,N_5378);
xnor U13963 (N_13963,N_6992,N_6056);
and U13964 (N_13964,N_9447,N_5812);
xor U13965 (N_13965,N_6586,N_9770);
and U13966 (N_13966,N_9072,N_9254);
and U13967 (N_13967,N_9517,N_7523);
nor U13968 (N_13968,N_7004,N_8979);
nor U13969 (N_13969,N_9332,N_8931);
xnor U13970 (N_13970,N_8489,N_7900);
nor U13971 (N_13971,N_7589,N_5745);
and U13972 (N_13972,N_6926,N_5114);
or U13973 (N_13973,N_5033,N_6085);
xor U13974 (N_13974,N_5630,N_8183);
or U13975 (N_13975,N_5620,N_8113);
xor U13976 (N_13976,N_9011,N_7197);
and U13977 (N_13977,N_8033,N_5091);
nand U13978 (N_13978,N_9250,N_5050);
xor U13979 (N_13979,N_6206,N_7096);
or U13980 (N_13980,N_8966,N_9377);
and U13981 (N_13981,N_8959,N_6067);
xor U13982 (N_13982,N_7899,N_9154);
or U13983 (N_13983,N_6422,N_7471);
nand U13984 (N_13984,N_8842,N_5339);
nor U13985 (N_13985,N_5311,N_7577);
xor U13986 (N_13986,N_5830,N_7221);
xnor U13987 (N_13987,N_9557,N_8833);
nor U13988 (N_13988,N_9845,N_5920);
and U13989 (N_13989,N_6906,N_7304);
and U13990 (N_13990,N_8839,N_8607);
nand U13991 (N_13991,N_7785,N_5154);
nand U13992 (N_13992,N_5044,N_9794);
xnor U13993 (N_13993,N_9061,N_8244);
or U13994 (N_13994,N_6431,N_8173);
nor U13995 (N_13995,N_8935,N_6285);
xnor U13996 (N_13996,N_8857,N_5128);
xor U13997 (N_13997,N_8241,N_9689);
or U13998 (N_13998,N_9203,N_8659);
nor U13999 (N_13999,N_9861,N_5424);
nor U14000 (N_14000,N_6025,N_7517);
xor U14001 (N_14001,N_5207,N_7210);
or U14002 (N_14002,N_7496,N_9046);
and U14003 (N_14003,N_9388,N_9103);
nor U14004 (N_14004,N_6313,N_5141);
nand U14005 (N_14005,N_6012,N_7766);
xor U14006 (N_14006,N_6945,N_7307);
nor U14007 (N_14007,N_9712,N_8899);
and U14008 (N_14008,N_8677,N_6398);
xor U14009 (N_14009,N_5921,N_8744);
and U14010 (N_14010,N_5445,N_9451);
nor U14011 (N_14011,N_5516,N_9009);
or U14012 (N_14012,N_7489,N_7503);
or U14013 (N_14013,N_8456,N_6853);
xor U14014 (N_14014,N_8001,N_5930);
or U14015 (N_14015,N_8869,N_6783);
xnor U14016 (N_14016,N_9698,N_8975);
nand U14017 (N_14017,N_6996,N_9071);
nor U14018 (N_14018,N_6796,N_8720);
nand U14019 (N_14019,N_9737,N_9017);
nor U14020 (N_14020,N_9158,N_5182);
nand U14021 (N_14021,N_6135,N_7421);
nor U14022 (N_14022,N_7454,N_7081);
nand U14023 (N_14023,N_5605,N_7941);
nor U14024 (N_14024,N_5852,N_7917);
and U14025 (N_14025,N_8024,N_6724);
xnor U14026 (N_14026,N_7068,N_6076);
nor U14027 (N_14027,N_5423,N_8808);
nand U14028 (N_14028,N_6961,N_9936);
xnor U14029 (N_14029,N_9754,N_5753);
nor U14030 (N_14030,N_9803,N_7807);
and U14031 (N_14031,N_5950,N_8147);
or U14032 (N_14032,N_6468,N_8137);
nand U14033 (N_14033,N_6633,N_9496);
or U14034 (N_14034,N_7254,N_9195);
nor U14035 (N_14035,N_7108,N_6026);
nand U14036 (N_14036,N_6166,N_5934);
or U14037 (N_14037,N_8035,N_9345);
and U14038 (N_14038,N_9887,N_8248);
xor U14039 (N_14039,N_7662,N_7686);
nand U14040 (N_14040,N_7001,N_6843);
and U14041 (N_14041,N_8815,N_8787);
nand U14042 (N_14042,N_7275,N_5978);
nor U14043 (N_14043,N_9103,N_7138);
and U14044 (N_14044,N_8895,N_9944);
or U14045 (N_14045,N_7553,N_5586);
and U14046 (N_14046,N_7380,N_9529);
nand U14047 (N_14047,N_6461,N_8570);
xnor U14048 (N_14048,N_8705,N_8315);
nand U14049 (N_14049,N_8827,N_9748);
xor U14050 (N_14050,N_7010,N_7394);
xnor U14051 (N_14051,N_8750,N_7286);
nand U14052 (N_14052,N_8581,N_8802);
or U14053 (N_14053,N_6572,N_6010);
nor U14054 (N_14054,N_6123,N_8556);
and U14055 (N_14055,N_7524,N_6602);
or U14056 (N_14056,N_8723,N_7582);
or U14057 (N_14057,N_8100,N_7286);
xnor U14058 (N_14058,N_5068,N_5685);
xor U14059 (N_14059,N_9842,N_8514);
nand U14060 (N_14060,N_6568,N_5499);
and U14061 (N_14061,N_5318,N_6453);
and U14062 (N_14062,N_9705,N_7991);
or U14063 (N_14063,N_7771,N_7154);
and U14064 (N_14064,N_9500,N_9660);
nor U14065 (N_14065,N_6716,N_5258);
and U14066 (N_14066,N_8911,N_9672);
or U14067 (N_14067,N_7740,N_9092);
and U14068 (N_14068,N_7637,N_8147);
or U14069 (N_14069,N_8111,N_8693);
nand U14070 (N_14070,N_6538,N_8321);
nor U14071 (N_14071,N_7980,N_9087);
nand U14072 (N_14072,N_8642,N_6961);
or U14073 (N_14073,N_9424,N_8018);
or U14074 (N_14074,N_6517,N_6029);
nand U14075 (N_14075,N_9038,N_7691);
xnor U14076 (N_14076,N_6519,N_9111);
xnor U14077 (N_14077,N_7073,N_7183);
nand U14078 (N_14078,N_9723,N_8547);
or U14079 (N_14079,N_6934,N_5368);
or U14080 (N_14080,N_5421,N_6734);
or U14081 (N_14081,N_8731,N_6193);
xnor U14082 (N_14082,N_7378,N_6766);
or U14083 (N_14083,N_8615,N_5958);
nand U14084 (N_14084,N_5806,N_7360);
and U14085 (N_14085,N_7052,N_7712);
or U14086 (N_14086,N_8737,N_5413);
or U14087 (N_14087,N_7976,N_9569);
nand U14088 (N_14088,N_5858,N_5415);
xor U14089 (N_14089,N_8402,N_6309);
nor U14090 (N_14090,N_5695,N_5754);
nor U14091 (N_14091,N_5204,N_8574);
xor U14092 (N_14092,N_8484,N_5839);
or U14093 (N_14093,N_8200,N_6250);
or U14094 (N_14094,N_5045,N_8255);
nor U14095 (N_14095,N_5753,N_8502);
nor U14096 (N_14096,N_6167,N_7587);
and U14097 (N_14097,N_7410,N_7074);
xor U14098 (N_14098,N_8934,N_9721);
nor U14099 (N_14099,N_6636,N_7823);
nor U14100 (N_14100,N_5602,N_6536);
nand U14101 (N_14101,N_5377,N_5373);
nand U14102 (N_14102,N_9301,N_6156);
or U14103 (N_14103,N_8233,N_7199);
xnor U14104 (N_14104,N_8607,N_6336);
or U14105 (N_14105,N_9520,N_8178);
and U14106 (N_14106,N_6246,N_8752);
xor U14107 (N_14107,N_8390,N_5034);
nand U14108 (N_14108,N_9384,N_9610);
and U14109 (N_14109,N_7509,N_5916);
xnor U14110 (N_14110,N_7208,N_6532);
nand U14111 (N_14111,N_7282,N_8609);
xor U14112 (N_14112,N_9495,N_6038);
or U14113 (N_14113,N_5861,N_9452);
nor U14114 (N_14114,N_7707,N_9526);
xnor U14115 (N_14115,N_8395,N_9858);
xnor U14116 (N_14116,N_7098,N_6209);
nor U14117 (N_14117,N_8076,N_5926);
xor U14118 (N_14118,N_8340,N_7982);
xor U14119 (N_14119,N_9237,N_5968);
nor U14120 (N_14120,N_6182,N_5878);
or U14121 (N_14121,N_6840,N_8409);
nand U14122 (N_14122,N_5855,N_8185);
or U14123 (N_14123,N_8632,N_9049);
and U14124 (N_14124,N_7151,N_6482);
xor U14125 (N_14125,N_7565,N_5661);
nand U14126 (N_14126,N_5866,N_6661);
or U14127 (N_14127,N_9641,N_7954);
and U14128 (N_14128,N_6428,N_6139);
nor U14129 (N_14129,N_9174,N_9711);
xor U14130 (N_14130,N_5763,N_8776);
nand U14131 (N_14131,N_9120,N_5107);
nand U14132 (N_14132,N_9464,N_8550);
xnor U14133 (N_14133,N_5440,N_6144);
xnor U14134 (N_14134,N_6704,N_9459);
or U14135 (N_14135,N_6708,N_6291);
and U14136 (N_14136,N_6110,N_6528);
and U14137 (N_14137,N_6281,N_6402);
nor U14138 (N_14138,N_6967,N_5200);
and U14139 (N_14139,N_5000,N_7659);
xnor U14140 (N_14140,N_8695,N_9320);
nand U14141 (N_14141,N_5403,N_6920);
or U14142 (N_14142,N_7150,N_6641);
and U14143 (N_14143,N_6414,N_7402);
xnor U14144 (N_14144,N_9280,N_6165);
nand U14145 (N_14145,N_5521,N_5724);
xnor U14146 (N_14146,N_9120,N_6423);
nor U14147 (N_14147,N_8239,N_9771);
nand U14148 (N_14148,N_9027,N_5228);
and U14149 (N_14149,N_9171,N_9564);
or U14150 (N_14150,N_9199,N_5588);
nand U14151 (N_14151,N_7786,N_8013);
xnor U14152 (N_14152,N_8324,N_6023);
or U14153 (N_14153,N_9921,N_8175);
and U14154 (N_14154,N_9812,N_5957);
nand U14155 (N_14155,N_9761,N_5410);
xor U14156 (N_14156,N_7905,N_6293);
and U14157 (N_14157,N_9873,N_5953);
or U14158 (N_14158,N_6831,N_7451);
nor U14159 (N_14159,N_7231,N_5588);
or U14160 (N_14160,N_7825,N_7249);
and U14161 (N_14161,N_9941,N_8883);
or U14162 (N_14162,N_5788,N_8216);
xor U14163 (N_14163,N_9637,N_9616);
nor U14164 (N_14164,N_5984,N_5681);
nand U14165 (N_14165,N_6661,N_7907);
or U14166 (N_14166,N_5626,N_5089);
nor U14167 (N_14167,N_6270,N_8514);
and U14168 (N_14168,N_6325,N_5427);
or U14169 (N_14169,N_9079,N_8914);
nor U14170 (N_14170,N_6396,N_8883);
or U14171 (N_14171,N_8999,N_7666);
and U14172 (N_14172,N_5151,N_5919);
nor U14173 (N_14173,N_5800,N_9262);
or U14174 (N_14174,N_9469,N_9984);
nor U14175 (N_14175,N_8788,N_5164);
or U14176 (N_14176,N_6109,N_6015);
nor U14177 (N_14177,N_5356,N_8578);
nor U14178 (N_14178,N_8548,N_9147);
nor U14179 (N_14179,N_8524,N_5534);
nor U14180 (N_14180,N_7767,N_8100);
xnor U14181 (N_14181,N_6756,N_8929);
or U14182 (N_14182,N_8152,N_7026);
nor U14183 (N_14183,N_7995,N_7428);
nor U14184 (N_14184,N_6802,N_6672);
or U14185 (N_14185,N_9392,N_6258);
and U14186 (N_14186,N_9054,N_6124);
or U14187 (N_14187,N_5245,N_7994);
and U14188 (N_14188,N_5649,N_5159);
and U14189 (N_14189,N_6364,N_9723);
nor U14190 (N_14190,N_8046,N_5420);
or U14191 (N_14191,N_7158,N_9078);
and U14192 (N_14192,N_7699,N_9866);
or U14193 (N_14193,N_5878,N_9126);
and U14194 (N_14194,N_5465,N_9649);
or U14195 (N_14195,N_5988,N_6845);
or U14196 (N_14196,N_6790,N_6347);
or U14197 (N_14197,N_8779,N_6362);
or U14198 (N_14198,N_8636,N_6047);
nor U14199 (N_14199,N_6237,N_8709);
nand U14200 (N_14200,N_8186,N_8875);
xnor U14201 (N_14201,N_5331,N_5099);
xnor U14202 (N_14202,N_5006,N_6067);
xnor U14203 (N_14203,N_9521,N_5261);
nand U14204 (N_14204,N_8329,N_7625);
nand U14205 (N_14205,N_9664,N_8820);
xor U14206 (N_14206,N_9291,N_6238);
xor U14207 (N_14207,N_7434,N_7086);
nor U14208 (N_14208,N_9035,N_9241);
or U14209 (N_14209,N_5910,N_6656);
nand U14210 (N_14210,N_6009,N_5697);
xnor U14211 (N_14211,N_5311,N_9985);
nand U14212 (N_14212,N_5681,N_6446);
xor U14213 (N_14213,N_5277,N_7411);
and U14214 (N_14214,N_5596,N_5190);
or U14215 (N_14215,N_9377,N_8915);
or U14216 (N_14216,N_5482,N_5372);
or U14217 (N_14217,N_5666,N_6357);
nand U14218 (N_14218,N_7328,N_8116);
and U14219 (N_14219,N_5826,N_9140);
or U14220 (N_14220,N_7537,N_8561);
or U14221 (N_14221,N_5097,N_9863);
nor U14222 (N_14222,N_5013,N_6156);
and U14223 (N_14223,N_5552,N_7836);
nor U14224 (N_14224,N_9314,N_9309);
nand U14225 (N_14225,N_9479,N_6619);
and U14226 (N_14226,N_6068,N_8503);
nand U14227 (N_14227,N_7871,N_7451);
nor U14228 (N_14228,N_5644,N_6582);
xnor U14229 (N_14229,N_5800,N_7923);
nor U14230 (N_14230,N_7436,N_7222);
and U14231 (N_14231,N_7522,N_6361);
nor U14232 (N_14232,N_9981,N_6134);
nor U14233 (N_14233,N_6909,N_6912);
or U14234 (N_14234,N_9940,N_8229);
and U14235 (N_14235,N_9130,N_6692);
or U14236 (N_14236,N_6516,N_6362);
or U14237 (N_14237,N_8868,N_8184);
nor U14238 (N_14238,N_5965,N_5966);
nand U14239 (N_14239,N_9767,N_8324);
nand U14240 (N_14240,N_7773,N_7653);
or U14241 (N_14241,N_8783,N_9348);
nand U14242 (N_14242,N_7784,N_6359);
and U14243 (N_14243,N_9143,N_7678);
and U14244 (N_14244,N_9049,N_6826);
or U14245 (N_14245,N_5107,N_6011);
or U14246 (N_14246,N_8315,N_5771);
or U14247 (N_14247,N_9183,N_9813);
xor U14248 (N_14248,N_7362,N_5885);
nor U14249 (N_14249,N_5995,N_8455);
xnor U14250 (N_14250,N_7729,N_8950);
nand U14251 (N_14251,N_9797,N_6475);
nand U14252 (N_14252,N_8511,N_8852);
or U14253 (N_14253,N_5958,N_5406);
xnor U14254 (N_14254,N_9477,N_5863);
and U14255 (N_14255,N_5460,N_8999);
xnor U14256 (N_14256,N_7972,N_7867);
xnor U14257 (N_14257,N_9241,N_7852);
and U14258 (N_14258,N_7510,N_9368);
nand U14259 (N_14259,N_8617,N_7838);
nor U14260 (N_14260,N_5443,N_7636);
nor U14261 (N_14261,N_7507,N_8008);
nand U14262 (N_14262,N_9686,N_6996);
nand U14263 (N_14263,N_5946,N_7972);
xnor U14264 (N_14264,N_7692,N_6072);
or U14265 (N_14265,N_9311,N_5006);
and U14266 (N_14266,N_5987,N_7493);
nor U14267 (N_14267,N_7732,N_9872);
nand U14268 (N_14268,N_7072,N_6750);
and U14269 (N_14269,N_6166,N_5787);
xnor U14270 (N_14270,N_6265,N_9319);
xnor U14271 (N_14271,N_9502,N_6034);
nor U14272 (N_14272,N_6327,N_9039);
or U14273 (N_14273,N_7431,N_5104);
nor U14274 (N_14274,N_8901,N_7282);
nand U14275 (N_14275,N_8802,N_5798);
or U14276 (N_14276,N_6016,N_7738);
and U14277 (N_14277,N_6405,N_8476);
nor U14278 (N_14278,N_6204,N_9573);
nor U14279 (N_14279,N_7325,N_5767);
nand U14280 (N_14280,N_6829,N_7681);
xnor U14281 (N_14281,N_9014,N_8117);
nand U14282 (N_14282,N_7399,N_9709);
xnor U14283 (N_14283,N_8295,N_9956);
or U14284 (N_14284,N_8972,N_9927);
nand U14285 (N_14285,N_6697,N_6348);
nand U14286 (N_14286,N_6548,N_9727);
nand U14287 (N_14287,N_7822,N_9866);
or U14288 (N_14288,N_6678,N_6298);
xnor U14289 (N_14289,N_7643,N_8406);
and U14290 (N_14290,N_6217,N_5960);
xor U14291 (N_14291,N_6279,N_8007);
xor U14292 (N_14292,N_8597,N_7250);
xnor U14293 (N_14293,N_7443,N_5689);
nor U14294 (N_14294,N_6916,N_5042);
xnor U14295 (N_14295,N_7327,N_7970);
and U14296 (N_14296,N_5861,N_5728);
nand U14297 (N_14297,N_9587,N_5612);
and U14298 (N_14298,N_8293,N_7667);
or U14299 (N_14299,N_8517,N_6362);
nor U14300 (N_14300,N_7439,N_8792);
or U14301 (N_14301,N_8481,N_8119);
xor U14302 (N_14302,N_5985,N_5684);
and U14303 (N_14303,N_9578,N_9524);
and U14304 (N_14304,N_7679,N_5126);
nor U14305 (N_14305,N_7574,N_5369);
or U14306 (N_14306,N_6943,N_8144);
or U14307 (N_14307,N_7292,N_5031);
xor U14308 (N_14308,N_9515,N_9526);
nand U14309 (N_14309,N_9805,N_9771);
nor U14310 (N_14310,N_7713,N_5611);
nand U14311 (N_14311,N_5905,N_5008);
and U14312 (N_14312,N_8595,N_7600);
xor U14313 (N_14313,N_8812,N_9683);
nand U14314 (N_14314,N_9812,N_6865);
nand U14315 (N_14315,N_5156,N_8516);
or U14316 (N_14316,N_6523,N_7782);
or U14317 (N_14317,N_7574,N_5106);
or U14318 (N_14318,N_5383,N_7176);
or U14319 (N_14319,N_6558,N_8423);
nand U14320 (N_14320,N_5876,N_5324);
nor U14321 (N_14321,N_9400,N_7891);
nor U14322 (N_14322,N_7430,N_5851);
nand U14323 (N_14323,N_8802,N_5520);
nand U14324 (N_14324,N_9137,N_7835);
nand U14325 (N_14325,N_9215,N_8622);
nor U14326 (N_14326,N_9596,N_9463);
nand U14327 (N_14327,N_9264,N_6900);
xor U14328 (N_14328,N_7428,N_9329);
and U14329 (N_14329,N_8469,N_8266);
nor U14330 (N_14330,N_6815,N_9546);
nor U14331 (N_14331,N_8436,N_5567);
xnor U14332 (N_14332,N_5112,N_9654);
nor U14333 (N_14333,N_5738,N_7848);
nand U14334 (N_14334,N_6614,N_5495);
nand U14335 (N_14335,N_8360,N_8427);
and U14336 (N_14336,N_5029,N_7338);
xnor U14337 (N_14337,N_8015,N_5268);
and U14338 (N_14338,N_5265,N_9079);
nand U14339 (N_14339,N_5531,N_9796);
xnor U14340 (N_14340,N_5914,N_9139);
nand U14341 (N_14341,N_7913,N_9262);
and U14342 (N_14342,N_8947,N_7107);
xnor U14343 (N_14343,N_8325,N_8235);
and U14344 (N_14344,N_6569,N_5207);
and U14345 (N_14345,N_8489,N_8509);
nand U14346 (N_14346,N_9658,N_8832);
or U14347 (N_14347,N_8481,N_7614);
and U14348 (N_14348,N_5386,N_7175);
nor U14349 (N_14349,N_5511,N_7997);
and U14350 (N_14350,N_8551,N_8675);
or U14351 (N_14351,N_8229,N_9503);
and U14352 (N_14352,N_7892,N_5069);
nor U14353 (N_14353,N_7059,N_5461);
nand U14354 (N_14354,N_6912,N_9634);
and U14355 (N_14355,N_8968,N_7637);
nand U14356 (N_14356,N_8312,N_5543);
nand U14357 (N_14357,N_6051,N_9306);
and U14358 (N_14358,N_6813,N_7906);
xor U14359 (N_14359,N_9513,N_7802);
and U14360 (N_14360,N_6354,N_8452);
or U14361 (N_14361,N_6965,N_5629);
and U14362 (N_14362,N_6877,N_7868);
and U14363 (N_14363,N_8958,N_6936);
and U14364 (N_14364,N_7560,N_5438);
nor U14365 (N_14365,N_9652,N_6992);
nor U14366 (N_14366,N_8611,N_6006);
nor U14367 (N_14367,N_6490,N_8341);
nand U14368 (N_14368,N_7529,N_5246);
or U14369 (N_14369,N_7103,N_9229);
nand U14370 (N_14370,N_7057,N_5015);
or U14371 (N_14371,N_7048,N_9257);
or U14372 (N_14372,N_5734,N_6557);
and U14373 (N_14373,N_5353,N_8164);
and U14374 (N_14374,N_6467,N_9308);
xor U14375 (N_14375,N_9500,N_5643);
nand U14376 (N_14376,N_7672,N_6275);
nor U14377 (N_14377,N_9223,N_5052);
xor U14378 (N_14378,N_5672,N_7382);
nand U14379 (N_14379,N_5175,N_9106);
nand U14380 (N_14380,N_6547,N_6529);
nand U14381 (N_14381,N_9406,N_5519);
or U14382 (N_14382,N_5955,N_7402);
or U14383 (N_14383,N_8351,N_7201);
nand U14384 (N_14384,N_5025,N_9678);
nand U14385 (N_14385,N_5229,N_7655);
xnor U14386 (N_14386,N_6459,N_9375);
or U14387 (N_14387,N_6988,N_8669);
nand U14388 (N_14388,N_7475,N_5146);
nor U14389 (N_14389,N_5262,N_6707);
nand U14390 (N_14390,N_9813,N_9087);
and U14391 (N_14391,N_9157,N_7246);
or U14392 (N_14392,N_7682,N_5519);
nand U14393 (N_14393,N_7621,N_7027);
nor U14394 (N_14394,N_6075,N_7932);
or U14395 (N_14395,N_8832,N_8379);
and U14396 (N_14396,N_6184,N_5065);
and U14397 (N_14397,N_8650,N_6938);
nor U14398 (N_14398,N_6439,N_8477);
and U14399 (N_14399,N_8229,N_5039);
or U14400 (N_14400,N_7369,N_8165);
xnor U14401 (N_14401,N_7922,N_6711);
and U14402 (N_14402,N_9266,N_6719);
xor U14403 (N_14403,N_7121,N_6676);
xnor U14404 (N_14404,N_6508,N_7257);
nor U14405 (N_14405,N_5583,N_5868);
xnor U14406 (N_14406,N_7977,N_7807);
xor U14407 (N_14407,N_7279,N_7420);
nand U14408 (N_14408,N_5798,N_5726);
nand U14409 (N_14409,N_9382,N_9295);
xnor U14410 (N_14410,N_5639,N_9841);
and U14411 (N_14411,N_9545,N_6632);
xnor U14412 (N_14412,N_5109,N_7501);
or U14413 (N_14413,N_5690,N_8335);
nand U14414 (N_14414,N_7788,N_7837);
xnor U14415 (N_14415,N_5583,N_9275);
or U14416 (N_14416,N_6984,N_9848);
nand U14417 (N_14417,N_8187,N_9633);
nand U14418 (N_14418,N_8909,N_9578);
and U14419 (N_14419,N_5725,N_7625);
xnor U14420 (N_14420,N_7798,N_8300);
nor U14421 (N_14421,N_6272,N_6815);
nand U14422 (N_14422,N_6882,N_5009);
and U14423 (N_14423,N_7027,N_5311);
nor U14424 (N_14424,N_6196,N_5443);
xnor U14425 (N_14425,N_6824,N_7912);
or U14426 (N_14426,N_7368,N_8112);
nor U14427 (N_14427,N_5982,N_9459);
and U14428 (N_14428,N_7063,N_8188);
or U14429 (N_14429,N_9467,N_7430);
nor U14430 (N_14430,N_7662,N_7849);
xor U14431 (N_14431,N_8488,N_9368);
nand U14432 (N_14432,N_6050,N_5527);
nor U14433 (N_14433,N_8176,N_7734);
nand U14434 (N_14434,N_9680,N_6575);
or U14435 (N_14435,N_5126,N_8793);
xnor U14436 (N_14436,N_8688,N_7921);
xor U14437 (N_14437,N_6476,N_9252);
nor U14438 (N_14438,N_8542,N_5154);
and U14439 (N_14439,N_9168,N_5710);
or U14440 (N_14440,N_8968,N_7716);
nand U14441 (N_14441,N_7516,N_9268);
nand U14442 (N_14442,N_8740,N_6948);
xor U14443 (N_14443,N_7817,N_7320);
and U14444 (N_14444,N_6597,N_8275);
nand U14445 (N_14445,N_7370,N_6227);
and U14446 (N_14446,N_8119,N_6111);
nor U14447 (N_14447,N_5676,N_9959);
xor U14448 (N_14448,N_6984,N_9575);
xnor U14449 (N_14449,N_5059,N_9144);
and U14450 (N_14450,N_8051,N_6016);
nor U14451 (N_14451,N_6921,N_5301);
xor U14452 (N_14452,N_9290,N_7902);
and U14453 (N_14453,N_6126,N_7903);
xor U14454 (N_14454,N_7786,N_9184);
nor U14455 (N_14455,N_8018,N_9848);
and U14456 (N_14456,N_7525,N_6950);
or U14457 (N_14457,N_7323,N_5881);
xnor U14458 (N_14458,N_9318,N_9265);
xnor U14459 (N_14459,N_5348,N_9163);
or U14460 (N_14460,N_8862,N_5281);
and U14461 (N_14461,N_8460,N_7778);
nor U14462 (N_14462,N_7540,N_8216);
or U14463 (N_14463,N_7499,N_5000);
or U14464 (N_14464,N_8978,N_8322);
nand U14465 (N_14465,N_7570,N_5585);
or U14466 (N_14466,N_5163,N_7841);
and U14467 (N_14467,N_5584,N_5666);
nand U14468 (N_14468,N_7173,N_9723);
xnor U14469 (N_14469,N_7277,N_6786);
and U14470 (N_14470,N_8335,N_7591);
xor U14471 (N_14471,N_8166,N_9521);
or U14472 (N_14472,N_9260,N_6389);
xor U14473 (N_14473,N_9439,N_6323);
or U14474 (N_14474,N_5062,N_5428);
nand U14475 (N_14475,N_6062,N_5536);
xnor U14476 (N_14476,N_5522,N_8451);
or U14477 (N_14477,N_8201,N_6207);
nand U14478 (N_14478,N_6244,N_9826);
nor U14479 (N_14479,N_7288,N_9776);
nor U14480 (N_14480,N_6747,N_7267);
or U14481 (N_14481,N_6740,N_9999);
or U14482 (N_14482,N_9121,N_6363);
nor U14483 (N_14483,N_8154,N_8944);
nor U14484 (N_14484,N_8309,N_7182);
or U14485 (N_14485,N_9875,N_5924);
or U14486 (N_14486,N_5460,N_6896);
xnor U14487 (N_14487,N_7312,N_7548);
nor U14488 (N_14488,N_6187,N_5504);
nand U14489 (N_14489,N_8109,N_6841);
or U14490 (N_14490,N_6009,N_8432);
and U14491 (N_14491,N_7835,N_6652);
nand U14492 (N_14492,N_5370,N_8534);
nor U14493 (N_14493,N_5405,N_7431);
nand U14494 (N_14494,N_7024,N_9767);
nor U14495 (N_14495,N_6693,N_6180);
xnor U14496 (N_14496,N_7940,N_6822);
or U14497 (N_14497,N_8456,N_7649);
and U14498 (N_14498,N_8744,N_7159);
and U14499 (N_14499,N_7604,N_5269);
xor U14500 (N_14500,N_5063,N_9757);
and U14501 (N_14501,N_6744,N_6701);
nand U14502 (N_14502,N_8319,N_6331);
or U14503 (N_14503,N_9837,N_7068);
xor U14504 (N_14504,N_7400,N_7151);
nor U14505 (N_14505,N_7138,N_7406);
nor U14506 (N_14506,N_8399,N_5595);
xnor U14507 (N_14507,N_7357,N_9459);
nor U14508 (N_14508,N_5859,N_6814);
and U14509 (N_14509,N_7621,N_5332);
nor U14510 (N_14510,N_8548,N_5834);
nand U14511 (N_14511,N_8885,N_6855);
and U14512 (N_14512,N_7672,N_8406);
and U14513 (N_14513,N_5034,N_6644);
nor U14514 (N_14514,N_5408,N_7027);
nor U14515 (N_14515,N_5196,N_9608);
and U14516 (N_14516,N_6814,N_5644);
xor U14517 (N_14517,N_8936,N_6402);
nor U14518 (N_14518,N_7906,N_7048);
xnor U14519 (N_14519,N_5811,N_6247);
nor U14520 (N_14520,N_8355,N_6916);
or U14521 (N_14521,N_7044,N_6415);
xnor U14522 (N_14522,N_7448,N_8669);
nand U14523 (N_14523,N_9144,N_8111);
and U14524 (N_14524,N_5984,N_5761);
nand U14525 (N_14525,N_8215,N_6172);
nand U14526 (N_14526,N_8844,N_8947);
and U14527 (N_14527,N_6351,N_9970);
and U14528 (N_14528,N_5464,N_8016);
or U14529 (N_14529,N_5016,N_9894);
or U14530 (N_14530,N_5333,N_8421);
and U14531 (N_14531,N_6627,N_7223);
nor U14532 (N_14532,N_6776,N_5570);
or U14533 (N_14533,N_5025,N_8415);
nand U14534 (N_14534,N_5278,N_7188);
xor U14535 (N_14535,N_5568,N_7187);
and U14536 (N_14536,N_9033,N_9174);
xnor U14537 (N_14537,N_6628,N_5876);
and U14538 (N_14538,N_8324,N_5306);
nor U14539 (N_14539,N_7110,N_6812);
nor U14540 (N_14540,N_9564,N_8376);
nand U14541 (N_14541,N_9713,N_7513);
nor U14542 (N_14542,N_6092,N_7449);
xnor U14543 (N_14543,N_5474,N_7739);
nand U14544 (N_14544,N_5991,N_5894);
or U14545 (N_14545,N_9859,N_5913);
and U14546 (N_14546,N_9210,N_8426);
nor U14547 (N_14547,N_7707,N_6093);
or U14548 (N_14548,N_8530,N_5847);
nand U14549 (N_14549,N_9742,N_7020);
nand U14550 (N_14550,N_8662,N_6099);
or U14551 (N_14551,N_9107,N_6823);
and U14552 (N_14552,N_6899,N_9242);
xnor U14553 (N_14553,N_5802,N_9201);
and U14554 (N_14554,N_9559,N_7356);
and U14555 (N_14555,N_7180,N_7624);
and U14556 (N_14556,N_9986,N_8264);
xor U14557 (N_14557,N_5790,N_6773);
and U14558 (N_14558,N_5828,N_8958);
nor U14559 (N_14559,N_8209,N_8134);
nand U14560 (N_14560,N_8498,N_7474);
or U14561 (N_14561,N_9967,N_6987);
nand U14562 (N_14562,N_5244,N_8289);
nor U14563 (N_14563,N_6765,N_6920);
nand U14564 (N_14564,N_6487,N_5339);
xnor U14565 (N_14565,N_9258,N_8104);
or U14566 (N_14566,N_8278,N_8204);
nand U14567 (N_14567,N_9079,N_8788);
or U14568 (N_14568,N_6849,N_8635);
and U14569 (N_14569,N_9820,N_9199);
or U14570 (N_14570,N_9115,N_5058);
nor U14571 (N_14571,N_7414,N_7512);
and U14572 (N_14572,N_7098,N_7808);
nor U14573 (N_14573,N_6907,N_6562);
nand U14574 (N_14574,N_6912,N_8231);
nor U14575 (N_14575,N_5853,N_7574);
and U14576 (N_14576,N_5119,N_8392);
xor U14577 (N_14577,N_6734,N_6197);
or U14578 (N_14578,N_6201,N_9087);
or U14579 (N_14579,N_7010,N_6211);
and U14580 (N_14580,N_5565,N_6844);
nand U14581 (N_14581,N_5786,N_7698);
nand U14582 (N_14582,N_8348,N_9147);
and U14583 (N_14583,N_5852,N_8392);
nor U14584 (N_14584,N_9545,N_5897);
or U14585 (N_14585,N_8075,N_6651);
nand U14586 (N_14586,N_6329,N_7573);
and U14587 (N_14587,N_9651,N_7327);
and U14588 (N_14588,N_5072,N_9177);
or U14589 (N_14589,N_5456,N_6901);
xnor U14590 (N_14590,N_6224,N_5392);
nor U14591 (N_14591,N_9413,N_6372);
nor U14592 (N_14592,N_5769,N_7491);
xnor U14593 (N_14593,N_8468,N_9186);
and U14594 (N_14594,N_6040,N_6341);
nand U14595 (N_14595,N_5084,N_9891);
xor U14596 (N_14596,N_7885,N_7154);
nor U14597 (N_14597,N_7462,N_6810);
or U14598 (N_14598,N_5217,N_7980);
nand U14599 (N_14599,N_5867,N_7358);
or U14600 (N_14600,N_6981,N_9891);
nand U14601 (N_14601,N_9103,N_9608);
or U14602 (N_14602,N_7263,N_6207);
or U14603 (N_14603,N_6158,N_7665);
nor U14604 (N_14604,N_9059,N_7833);
xor U14605 (N_14605,N_5020,N_6815);
or U14606 (N_14606,N_8679,N_7734);
nand U14607 (N_14607,N_5571,N_8953);
and U14608 (N_14608,N_7049,N_6297);
nand U14609 (N_14609,N_7836,N_5941);
xnor U14610 (N_14610,N_7867,N_5090);
nand U14611 (N_14611,N_8049,N_6242);
and U14612 (N_14612,N_7806,N_8801);
nor U14613 (N_14613,N_7983,N_8127);
nand U14614 (N_14614,N_7677,N_8533);
nor U14615 (N_14615,N_9768,N_6758);
nand U14616 (N_14616,N_5515,N_8767);
xnor U14617 (N_14617,N_9079,N_5671);
or U14618 (N_14618,N_5295,N_5140);
xnor U14619 (N_14619,N_7799,N_8454);
xor U14620 (N_14620,N_7986,N_5281);
nand U14621 (N_14621,N_6810,N_9409);
nor U14622 (N_14622,N_5801,N_8240);
and U14623 (N_14623,N_9364,N_9251);
and U14624 (N_14624,N_6246,N_5218);
nor U14625 (N_14625,N_5869,N_9799);
xor U14626 (N_14626,N_7168,N_9812);
and U14627 (N_14627,N_6596,N_7477);
xnor U14628 (N_14628,N_5447,N_8410);
and U14629 (N_14629,N_6635,N_5288);
nor U14630 (N_14630,N_8730,N_5486);
and U14631 (N_14631,N_5631,N_7764);
or U14632 (N_14632,N_8885,N_9269);
and U14633 (N_14633,N_8102,N_6149);
nor U14634 (N_14634,N_8694,N_5973);
nor U14635 (N_14635,N_6624,N_7635);
and U14636 (N_14636,N_5212,N_8003);
xor U14637 (N_14637,N_7744,N_8596);
nor U14638 (N_14638,N_5102,N_7930);
nand U14639 (N_14639,N_5492,N_5279);
xor U14640 (N_14640,N_5142,N_9904);
or U14641 (N_14641,N_7579,N_8472);
nand U14642 (N_14642,N_6078,N_9020);
nand U14643 (N_14643,N_8002,N_7952);
or U14644 (N_14644,N_8132,N_9721);
nand U14645 (N_14645,N_6177,N_5297);
nor U14646 (N_14646,N_9167,N_9228);
xnor U14647 (N_14647,N_6593,N_7131);
nand U14648 (N_14648,N_6219,N_9367);
or U14649 (N_14649,N_8065,N_6928);
and U14650 (N_14650,N_5815,N_7186);
and U14651 (N_14651,N_8842,N_5610);
xor U14652 (N_14652,N_6167,N_9351);
or U14653 (N_14653,N_5657,N_8560);
nor U14654 (N_14654,N_5393,N_5228);
nand U14655 (N_14655,N_7979,N_9227);
xor U14656 (N_14656,N_6901,N_8363);
xor U14657 (N_14657,N_8240,N_6019);
nor U14658 (N_14658,N_5638,N_6724);
or U14659 (N_14659,N_7201,N_9502);
and U14660 (N_14660,N_7602,N_5304);
xor U14661 (N_14661,N_5550,N_8509);
and U14662 (N_14662,N_9953,N_5286);
nor U14663 (N_14663,N_7355,N_9492);
xor U14664 (N_14664,N_5946,N_6638);
and U14665 (N_14665,N_8068,N_9765);
and U14666 (N_14666,N_6726,N_5593);
nand U14667 (N_14667,N_5262,N_6073);
and U14668 (N_14668,N_9806,N_7300);
nand U14669 (N_14669,N_5777,N_8737);
nand U14670 (N_14670,N_7620,N_9632);
nand U14671 (N_14671,N_9111,N_9685);
nor U14672 (N_14672,N_5269,N_9414);
xnor U14673 (N_14673,N_9554,N_6943);
or U14674 (N_14674,N_9039,N_6692);
and U14675 (N_14675,N_5516,N_9001);
nand U14676 (N_14676,N_9900,N_5634);
nand U14677 (N_14677,N_9386,N_5655);
or U14678 (N_14678,N_6823,N_5953);
or U14679 (N_14679,N_7941,N_8359);
nand U14680 (N_14680,N_9051,N_9565);
nand U14681 (N_14681,N_6981,N_8165);
nor U14682 (N_14682,N_5195,N_8409);
nand U14683 (N_14683,N_7313,N_9914);
and U14684 (N_14684,N_6766,N_7264);
xnor U14685 (N_14685,N_8423,N_8187);
or U14686 (N_14686,N_5126,N_6872);
nor U14687 (N_14687,N_6366,N_9901);
and U14688 (N_14688,N_9539,N_5989);
nand U14689 (N_14689,N_8400,N_6992);
nand U14690 (N_14690,N_7720,N_7175);
or U14691 (N_14691,N_7774,N_8824);
xor U14692 (N_14692,N_9245,N_7072);
and U14693 (N_14693,N_9344,N_5390);
xnor U14694 (N_14694,N_6944,N_5454);
nand U14695 (N_14695,N_5299,N_7764);
xnor U14696 (N_14696,N_5767,N_9066);
nand U14697 (N_14697,N_7829,N_6984);
xor U14698 (N_14698,N_6679,N_9229);
and U14699 (N_14699,N_6420,N_7052);
nand U14700 (N_14700,N_5492,N_7080);
nor U14701 (N_14701,N_9334,N_9824);
and U14702 (N_14702,N_9490,N_7547);
or U14703 (N_14703,N_9229,N_9786);
or U14704 (N_14704,N_6053,N_7154);
nor U14705 (N_14705,N_7080,N_6346);
and U14706 (N_14706,N_9896,N_8409);
or U14707 (N_14707,N_7329,N_7488);
and U14708 (N_14708,N_6414,N_6148);
nor U14709 (N_14709,N_5947,N_9961);
xnor U14710 (N_14710,N_8549,N_9258);
or U14711 (N_14711,N_9791,N_8056);
or U14712 (N_14712,N_7216,N_9381);
nor U14713 (N_14713,N_9265,N_7417);
nand U14714 (N_14714,N_9967,N_8365);
xor U14715 (N_14715,N_5185,N_7410);
and U14716 (N_14716,N_5743,N_6423);
nor U14717 (N_14717,N_5310,N_7198);
xor U14718 (N_14718,N_9736,N_8532);
nand U14719 (N_14719,N_9830,N_5512);
xnor U14720 (N_14720,N_6459,N_7217);
nor U14721 (N_14721,N_7169,N_8536);
nand U14722 (N_14722,N_9386,N_9936);
or U14723 (N_14723,N_5498,N_9929);
nor U14724 (N_14724,N_5122,N_9755);
and U14725 (N_14725,N_7069,N_5828);
or U14726 (N_14726,N_7329,N_9348);
and U14727 (N_14727,N_9789,N_7068);
xor U14728 (N_14728,N_9420,N_7249);
and U14729 (N_14729,N_6190,N_7612);
nor U14730 (N_14730,N_8170,N_7341);
xor U14731 (N_14731,N_8319,N_6699);
and U14732 (N_14732,N_9378,N_5247);
nor U14733 (N_14733,N_7288,N_6260);
nand U14734 (N_14734,N_7168,N_5394);
and U14735 (N_14735,N_8891,N_6284);
xor U14736 (N_14736,N_6667,N_9397);
and U14737 (N_14737,N_7603,N_6489);
xnor U14738 (N_14738,N_6509,N_5551);
nand U14739 (N_14739,N_7806,N_6513);
nand U14740 (N_14740,N_6993,N_7438);
xor U14741 (N_14741,N_5435,N_8363);
xnor U14742 (N_14742,N_7186,N_5675);
nand U14743 (N_14743,N_6497,N_7904);
and U14744 (N_14744,N_9847,N_7964);
nand U14745 (N_14745,N_9960,N_9337);
xnor U14746 (N_14746,N_5834,N_9398);
nand U14747 (N_14747,N_8410,N_6919);
and U14748 (N_14748,N_5714,N_6116);
xnor U14749 (N_14749,N_7209,N_6318);
and U14750 (N_14750,N_7504,N_9155);
nor U14751 (N_14751,N_5994,N_9377);
xor U14752 (N_14752,N_6296,N_6689);
xnor U14753 (N_14753,N_9952,N_9455);
xor U14754 (N_14754,N_5481,N_8295);
xnor U14755 (N_14755,N_6496,N_7044);
and U14756 (N_14756,N_7267,N_6264);
nor U14757 (N_14757,N_9176,N_7095);
or U14758 (N_14758,N_9630,N_8892);
xor U14759 (N_14759,N_7493,N_5613);
nand U14760 (N_14760,N_6812,N_7325);
xor U14761 (N_14761,N_7960,N_7388);
or U14762 (N_14762,N_9891,N_9462);
or U14763 (N_14763,N_5777,N_9216);
xor U14764 (N_14764,N_7332,N_8616);
and U14765 (N_14765,N_6061,N_7010);
xor U14766 (N_14766,N_7476,N_9153);
and U14767 (N_14767,N_7768,N_6602);
nor U14768 (N_14768,N_6012,N_7756);
nand U14769 (N_14769,N_6872,N_9809);
or U14770 (N_14770,N_7184,N_5986);
xor U14771 (N_14771,N_5737,N_6947);
nand U14772 (N_14772,N_5672,N_5943);
or U14773 (N_14773,N_6517,N_8439);
xnor U14774 (N_14774,N_8633,N_8545);
nand U14775 (N_14775,N_6479,N_7773);
xnor U14776 (N_14776,N_7202,N_7339);
nand U14777 (N_14777,N_8621,N_7599);
nor U14778 (N_14778,N_6297,N_5450);
nand U14779 (N_14779,N_7939,N_8437);
or U14780 (N_14780,N_6994,N_8440);
or U14781 (N_14781,N_6699,N_5003);
or U14782 (N_14782,N_8870,N_7610);
nor U14783 (N_14783,N_7700,N_6754);
and U14784 (N_14784,N_6930,N_7642);
or U14785 (N_14785,N_6571,N_7238);
nand U14786 (N_14786,N_8486,N_6807);
nand U14787 (N_14787,N_9912,N_8480);
xnor U14788 (N_14788,N_6681,N_5296);
xor U14789 (N_14789,N_8061,N_5549);
nor U14790 (N_14790,N_6308,N_9948);
or U14791 (N_14791,N_8431,N_7649);
or U14792 (N_14792,N_6178,N_9794);
or U14793 (N_14793,N_6242,N_6930);
xnor U14794 (N_14794,N_8571,N_9298);
nor U14795 (N_14795,N_7606,N_7624);
and U14796 (N_14796,N_5120,N_7407);
xnor U14797 (N_14797,N_7011,N_6762);
or U14798 (N_14798,N_8361,N_8973);
xnor U14799 (N_14799,N_6601,N_9454);
nand U14800 (N_14800,N_5672,N_7006);
nand U14801 (N_14801,N_5119,N_6648);
and U14802 (N_14802,N_8576,N_6148);
nor U14803 (N_14803,N_8868,N_7801);
nor U14804 (N_14804,N_7216,N_7543);
xor U14805 (N_14805,N_6181,N_5820);
and U14806 (N_14806,N_8776,N_9568);
nor U14807 (N_14807,N_9283,N_8074);
or U14808 (N_14808,N_8230,N_8593);
xnor U14809 (N_14809,N_7132,N_8322);
xor U14810 (N_14810,N_9195,N_8983);
and U14811 (N_14811,N_6854,N_5136);
or U14812 (N_14812,N_8496,N_9827);
nor U14813 (N_14813,N_6087,N_5153);
xnor U14814 (N_14814,N_5620,N_7619);
nand U14815 (N_14815,N_8357,N_5353);
nand U14816 (N_14816,N_8065,N_9043);
nand U14817 (N_14817,N_6844,N_5660);
nand U14818 (N_14818,N_8423,N_5056);
nor U14819 (N_14819,N_9787,N_9871);
nor U14820 (N_14820,N_8997,N_9328);
xnor U14821 (N_14821,N_7720,N_9112);
and U14822 (N_14822,N_7892,N_6002);
nand U14823 (N_14823,N_5963,N_6310);
xnor U14824 (N_14824,N_7402,N_6989);
nand U14825 (N_14825,N_7648,N_8805);
and U14826 (N_14826,N_5604,N_9007);
xnor U14827 (N_14827,N_6301,N_8276);
nand U14828 (N_14828,N_9496,N_5376);
xor U14829 (N_14829,N_9995,N_9838);
nor U14830 (N_14830,N_6567,N_8847);
xor U14831 (N_14831,N_6242,N_7910);
or U14832 (N_14832,N_7350,N_6735);
nor U14833 (N_14833,N_6765,N_9317);
xor U14834 (N_14834,N_7051,N_9637);
nand U14835 (N_14835,N_9422,N_5108);
and U14836 (N_14836,N_5946,N_9427);
xnor U14837 (N_14837,N_6549,N_7712);
nand U14838 (N_14838,N_7773,N_9257);
xnor U14839 (N_14839,N_7375,N_8324);
nor U14840 (N_14840,N_8841,N_9718);
and U14841 (N_14841,N_5197,N_5486);
nor U14842 (N_14842,N_6304,N_6382);
and U14843 (N_14843,N_9340,N_6705);
nand U14844 (N_14844,N_9632,N_7765);
and U14845 (N_14845,N_8637,N_6016);
xnor U14846 (N_14846,N_6296,N_8636);
and U14847 (N_14847,N_6659,N_6698);
and U14848 (N_14848,N_7904,N_5881);
nor U14849 (N_14849,N_6947,N_7250);
and U14850 (N_14850,N_5095,N_7881);
nor U14851 (N_14851,N_6584,N_6165);
nor U14852 (N_14852,N_9134,N_6329);
nor U14853 (N_14853,N_7960,N_6385);
nand U14854 (N_14854,N_5198,N_9215);
nand U14855 (N_14855,N_9492,N_7599);
and U14856 (N_14856,N_8897,N_5085);
xor U14857 (N_14857,N_5504,N_6295);
xnor U14858 (N_14858,N_5450,N_8258);
nor U14859 (N_14859,N_7525,N_7722);
nor U14860 (N_14860,N_5392,N_9546);
xnor U14861 (N_14861,N_7456,N_8481);
or U14862 (N_14862,N_6392,N_9114);
xor U14863 (N_14863,N_6529,N_5588);
nor U14864 (N_14864,N_7176,N_9219);
or U14865 (N_14865,N_7790,N_6058);
nand U14866 (N_14866,N_9067,N_8856);
xnor U14867 (N_14867,N_9294,N_8787);
nor U14868 (N_14868,N_9058,N_7697);
nor U14869 (N_14869,N_7785,N_9485);
and U14870 (N_14870,N_7785,N_8210);
xor U14871 (N_14871,N_9288,N_7126);
nand U14872 (N_14872,N_8931,N_5819);
xnor U14873 (N_14873,N_6372,N_9407);
or U14874 (N_14874,N_7018,N_5687);
and U14875 (N_14875,N_8477,N_7668);
and U14876 (N_14876,N_9789,N_9179);
nor U14877 (N_14877,N_9343,N_5364);
nand U14878 (N_14878,N_7072,N_5704);
xor U14879 (N_14879,N_7398,N_9186);
xor U14880 (N_14880,N_7684,N_6749);
nand U14881 (N_14881,N_8342,N_9954);
nor U14882 (N_14882,N_8416,N_7204);
nand U14883 (N_14883,N_5670,N_9686);
xnor U14884 (N_14884,N_5415,N_9006);
nor U14885 (N_14885,N_6717,N_6446);
nor U14886 (N_14886,N_5203,N_7267);
nor U14887 (N_14887,N_6153,N_8723);
nor U14888 (N_14888,N_7361,N_7488);
or U14889 (N_14889,N_8999,N_6491);
nand U14890 (N_14890,N_7334,N_6766);
nand U14891 (N_14891,N_5979,N_7856);
nor U14892 (N_14892,N_9239,N_9616);
and U14893 (N_14893,N_6805,N_7717);
nor U14894 (N_14894,N_9700,N_7957);
or U14895 (N_14895,N_7085,N_6177);
nand U14896 (N_14896,N_9365,N_8045);
or U14897 (N_14897,N_5639,N_8165);
or U14898 (N_14898,N_5499,N_7886);
and U14899 (N_14899,N_6606,N_6192);
or U14900 (N_14900,N_6826,N_6054);
and U14901 (N_14901,N_8096,N_6117);
nor U14902 (N_14902,N_5543,N_5549);
or U14903 (N_14903,N_6648,N_8150);
or U14904 (N_14904,N_8379,N_8518);
nor U14905 (N_14905,N_6168,N_9907);
nand U14906 (N_14906,N_6504,N_8058);
xnor U14907 (N_14907,N_5008,N_6757);
and U14908 (N_14908,N_9069,N_9242);
xor U14909 (N_14909,N_9999,N_7429);
xor U14910 (N_14910,N_5109,N_9073);
or U14911 (N_14911,N_7011,N_7516);
nand U14912 (N_14912,N_5690,N_6877);
nand U14913 (N_14913,N_8846,N_9896);
or U14914 (N_14914,N_8868,N_9846);
and U14915 (N_14915,N_7804,N_9373);
nand U14916 (N_14916,N_7700,N_8487);
xnor U14917 (N_14917,N_8190,N_8119);
nand U14918 (N_14918,N_9809,N_8524);
and U14919 (N_14919,N_7181,N_7398);
nor U14920 (N_14920,N_6460,N_6450);
and U14921 (N_14921,N_6602,N_8683);
nor U14922 (N_14922,N_5189,N_5193);
and U14923 (N_14923,N_5677,N_7694);
nand U14924 (N_14924,N_5872,N_7109);
nand U14925 (N_14925,N_5773,N_8482);
and U14926 (N_14926,N_9006,N_5595);
xor U14927 (N_14927,N_8859,N_9341);
xnor U14928 (N_14928,N_7858,N_5922);
xnor U14929 (N_14929,N_6210,N_8213);
nor U14930 (N_14930,N_8460,N_7749);
xnor U14931 (N_14931,N_8443,N_5338);
xor U14932 (N_14932,N_5897,N_8981);
or U14933 (N_14933,N_8358,N_6791);
xnor U14934 (N_14934,N_9658,N_6926);
xor U14935 (N_14935,N_8816,N_9500);
or U14936 (N_14936,N_6053,N_6457);
and U14937 (N_14937,N_6663,N_8842);
xnor U14938 (N_14938,N_8083,N_5435);
nor U14939 (N_14939,N_7499,N_7055);
xor U14940 (N_14940,N_7859,N_6590);
or U14941 (N_14941,N_9025,N_6695);
or U14942 (N_14942,N_5662,N_6636);
or U14943 (N_14943,N_9179,N_5173);
or U14944 (N_14944,N_9763,N_7596);
and U14945 (N_14945,N_5421,N_9117);
nand U14946 (N_14946,N_8219,N_7747);
nor U14947 (N_14947,N_7313,N_6761);
xnor U14948 (N_14948,N_5382,N_6543);
nor U14949 (N_14949,N_8827,N_5104);
nand U14950 (N_14950,N_9635,N_6864);
nor U14951 (N_14951,N_5268,N_7186);
and U14952 (N_14952,N_8936,N_5566);
or U14953 (N_14953,N_7092,N_7072);
nand U14954 (N_14954,N_6320,N_9456);
xor U14955 (N_14955,N_7755,N_7528);
nand U14956 (N_14956,N_5503,N_8620);
xnor U14957 (N_14957,N_6588,N_9591);
or U14958 (N_14958,N_9355,N_6721);
and U14959 (N_14959,N_9759,N_5745);
or U14960 (N_14960,N_6764,N_6319);
nor U14961 (N_14961,N_9695,N_9242);
or U14962 (N_14962,N_8195,N_7659);
and U14963 (N_14963,N_9634,N_8126);
nand U14964 (N_14964,N_8983,N_9037);
and U14965 (N_14965,N_7083,N_9348);
nor U14966 (N_14966,N_6812,N_6115);
nand U14967 (N_14967,N_6381,N_7780);
or U14968 (N_14968,N_9032,N_7139);
or U14969 (N_14969,N_6985,N_9613);
xnor U14970 (N_14970,N_9022,N_6494);
nor U14971 (N_14971,N_6580,N_7192);
nand U14972 (N_14972,N_8675,N_7892);
and U14973 (N_14973,N_8302,N_5216);
or U14974 (N_14974,N_8945,N_7155);
and U14975 (N_14975,N_5450,N_5336);
xnor U14976 (N_14976,N_7723,N_8046);
nor U14977 (N_14977,N_6606,N_7373);
nand U14978 (N_14978,N_9438,N_5527);
nor U14979 (N_14979,N_7379,N_5599);
nand U14980 (N_14980,N_5940,N_8387);
and U14981 (N_14981,N_9639,N_6090);
and U14982 (N_14982,N_9403,N_8459);
and U14983 (N_14983,N_9123,N_7415);
nand U14984 (N_14984,N_8793,N_9302);
and U14985 (N_14985,N_6466,N_7083);
or U14986 (N_14986,N_6781,N_5799);
or U14987 (N_14987,N_5960,N_7827);
xor U14988 (N_14988,N_9465,N_6589);
nor U14989 (N_14989,N_6874,N_7082);
or U14990 (N_14990,N_7494,N_8680);
and U14991 (N_14991,N_9023,N_8768);
xor U14992 (N_14992,N_5182,N_8734);
xor U14993 (N_14993,N_9062,N_8003);
or U14994 (N_14994,N_8006,N_6695);
nand U14995 (N_14995,N_9804,N_8782);
nor U14996 (N_14996,N_6586,N_6474);
nor U14997 (N_14997,N_7494,N_9809);
or U14998 (N_14998,N_6465,N_6836);
xnor U14999 (N_14999,N_7669,N_7796);
xnor U15000 (N_15000,N_11922,N_13644);
and U15001 (N_15001,N_10599,N_11855);
xor U15002 (N_15002,N_10369,N_14285);
and U15003 (N_15003,N_13605,N_13778);
and U15004 (N_15004,N_11594,N_11972);
or U15005 (N_15005,N_11046,N_11042);
or U15006 (N_15006,N_13746,N_14405);
and U15007 (N_15007,N_14306,N_12722);
nor U15008 (N_15008,N_11707,N_10563);
and U15009 (N_15009,N_10005,N_12561);
nand U15010 (N_15010,N_12756,N_14483);
nand U15011 (N_15011,N_14169,N_12572);
and U15012 (N_15012,N_11664,N_14009);
or U15013 (N_15013,N_12611,N_10742);
xor U15014 (N_15014,N_10684,N_12869);
and U15015 (N_15015,N_11242,N_14017);
xor U15016 (N_15016,N_13054,N_14945);
or U15017 (N_15017,N_13362,N_12167);
or U15018 (N_15018,N_13081,N_11569);
or U15019 (N_15019,N_13999,N_10003);
xnor U15020 (N_15020,N_13516,N_14890);
or U15021 (N_15021,N_14880,N_11806);
or U15022 (N_15022,N_13522,N_10307);
xnor U15023 (N_15023,N_14246,N_13303);
xor U15024 (N_15024,N_12150,N_11198);
and U15025 (N_15025,N_13569,N_13821);
and U15026 (N_15026,N_12099,N_10553);
and U15027 (N_15027,N_13685,N_13373);
nor U15028 (N_15028,N_14682,N_14591);
xnor U15029 (N_15029,N_12841,N_14082);
nand U15030 (N_15030,N_12848,N_14923);
nand U15031 (N_15031,N_11607,N_11061);
nor U15032 (N_15032,N_13288,N_13940);
xnor U15033 (N_15033,N_14393,N_11251);
xnor U15034 (N_15034,N_11249,N_12781);
and U15035 (N_15035,N_13631,N_12342);
or U15036 (N_15036,N_14069,N_12325);
and U15037 (N_15037,N_11580,N_12002);
nand U15038 (N_15038,N_11441,N_13211);
nand U15039 (N_15039,N_13833,N_13780);
nor U15040 (N_15040,N_14810,N_12202);
and U15041 (N_15041,N_14546,N_11934);
nand U15042 (N_15042,N_10359,N_11330);
nand U15043 (N_15043,N_10638,N_14608);
or U15044 (N_15044,N_14566,N_13931);
nor U15045 (N_15045,N_13567,N_12193);
or U15046 (N_15046,N_13718,N_11502);
nand U15047 (N_15047,N_12844,N_12017);
nor U15048 (N_15048,N_12030,N_11630);
xnor U15049 (N_15049,N_12967,N_11228);
nand U15050 (N_15050,N_12726,N_11421);
nand U15051 (N_15051,N_14136,N_13483);
nand U15052 (N_15052,N_11811,N_12270);
nand U15053 (N_15053,N_14953,N_14585);
nand U15054 (N_15054,N_13760,N_13727);
nor U15055 (N_15055,N_10273,N_13537);
xor U15056 (N_15056,N_11747,N_10755);
nand U15057 (N_15057,N_10015,N_12783);
nor U15058 (N_15058,N_11923,N_10828);
nand U15059 (N_15059,N_12942,N_13520);
xor U15060 (N_15060,N_12836,N_13160);
nor U15061 (N_15061,N_13800,N_13802);
nand U15062 (N_15062,N_12889,N_14827);
or U15063 (N_15063,N_13393,N_11037);
or U15064 (N_15064,N_14223,N_13268);
and U15065 (N_15065,N_13655,N_12935);
or U15066 (N_15066,N_11842,N_13378);
nand U15067 (N_15067,N_12898,N_13291);
xnor U15068 (N_15068,N_12331,N_11087);
nand U15069 (N_15069,N_11234,N_14820);
xor U15070 (N_15070,N_10110,N_10004);
xor U15071 (N_15071,N_14441,N_14869);
nand U15072 (N_15072,N_11907,N_11645);
and U15073 (N_15073,N_10006,N_10929);
or U15074 (N_15074,N_14812,N_14486);
nor U15075 (N_15075,N_12178,N_10132);
nand U15076 (N_15076,N_14843,N_11759);
xor U15077 (N_15077,N_14061,N_12300);
nand U15078 (N_15078,N_13016,N_13048);
nor U15079 (N_15079,N_11791,N_10102);
or U15080 (N_15080,N_12038,N_11932);
nor U15081 (N_15081,N_13105,N_13256);
and U15082 (N_15082,N_12493,N_10028);
nor U15083 (N_15083,N_14543,N_11702);
and U15084 (N_15084,N_11287,N_13353);
nand U15085 (N_15085,N_11601,N_13799);
or U15086 (N_15086,N_13429,N_11629);
or U15087 (N_15087,N_11976,N_13887);
nor U15088 (N_15088,N_13757,N_11690);
or U15089 (N_15089,N_13039,N_12091);
or U15090 (N_15090,N_14016,N_11940);
xor U15091 (N_15091,N_13910,N_12174);
xnor U15092 (N_15092,N_14348,N_13262);
or U15093 (N_15093,N_10649,N_11264);
nand U15094 (N_15094,N_11962,N_11399);
xor U15095 (N_15095,N_10375,N_11205);
and U15096 (N_15096,N_12360,N_12434);
nand U15097 (N_15097,N_14251,N_14421);
xnor U15098 (N_15098,N_13509,N_14078);
xnor U15099 (N_15099,N_11429,N_10148);
or U15100 (N_15100,N_12686,N_14817);
nand U15101 (N_15101,N_14889,N_14844);
xnor U15102 (N_15102,N_12226,N_13731);
xor U15103 (N_15103,N_14095,N_13187);
nand U15104 (N_15104,N_10945,N_14615);
or U15105 (N_15105,N_11807,N_12636);
nand U15106 (N_15106,N_12142,N_14627);
nand U15107 (N_15107,N_10352,N_11154);
or U15108 (N_15108,N_14811,N_12590);
xnor U15109 (N_15109,N_11256,N_12779);
nor U15110 (N_15110,N_14231,N_12734);
nor U15111 (N_15111,N_13664,N_13492);
nor U15112 (N_15112,N_12536,N_12409);
nor U15113 (N_15113,N_14775,N_14765);
nand U15114 (N_15114,N_13025,N_13672);
or U15115 (N_15115,N_13452,N_11563);
nor U15116 (N_15116,N_11127,N_14771);
nand U15117 (N_15117,N_10286,N_10205);
and U15118 (N_15118,N_11863,N_14093);
nand U15119 (N_15119,N_11175,N_14279);
nand U15120 (N_15120,N_14891,N_10407);
xnor U15121 (N_15121,N_11297,N_10770);
nor U15122 (N_15122,N_13488,N_13365);
or U15123 (N_15123,N_12388,N_10486);
or U15124 (N_15124,N_11944,N_14792);
nor U15125 (N_15125,N_11440,N_14362);
xor U15126 (N_15126,N_10926,N_11659);
nor U15127 (N_15127,N_13148,N_12111);
or U15128 (N_15128,N_13647,N_12698);
nor U15129 (N_15129,N_12778,N_13611);
xnor U15130 (N_15130,N_12653,N_11606);
and U15131 (N_15131,N_14667,N_10960);
nand U15132 (N_15132,N_14145,N_11374);
xor U15133 (N_15133,N_14268,N_14902);
xnor U15134 (N_15134,N_12981,N_14135);
and U15135 (N_15135,N_10117,N_13696);
nand U15136 (N_15136,N_11681,N_14311);
nor U15137 (N_15137,N_10878,N_14939);
xnor U15138 (N_15138,N_14727,N_14328);
and U15139 (N_15139,N_12658,N_10833);
and U15140 (N_15140,N_12158,N_12065);
nand U15141 (N_15141,N_13563,N_13546);
nand U15142 (N_15142,N_10194,N_12064);
xnor U15143 (N_15143,N_11617,N_12309);
and U15144 (N_15144,N_10387,N_12659);
xor U15145 (N_15145,N_12947,N_12149);
nand U15146 (N_15146,N_11847,N_14371);
and U15147 (N_15147,N_14090,N_10955);
nor U15148 (N_15148,N_10776,N_14720);
or U15149 (N_15149,N_10645,N_14332);
nor U15150 (N_15150,N_12170,N_12556);
nor U15151 (N_15151,N_13164,N_12943);
nor U15152 (N_15152,N_13857,N_12864);
xnor U15153 (N_15153,N_10094,N_10618);
nand U15154 (N_15154,N_10503,N_13572);
nor U15155 (N_15155,N_12444,N_10760);
nand U15156 (N_15156,N_14446,N_14665);
and U15157 (N_15157,N_10850,N_12912);
nand U15158 (N_15158,N_12752,N_13624);
nor U15159 (N_15159,N_14507,N_11953);
or U15160 (N_15160,N_10839,N_10548);
nor U15161 (N_15161,N_11883,N_11189);
or U15162 (N_15162,N_13769,N_14555);
or U15163 (N_15163,N_14607,N_12794);
or U15164 (N_15164,N_10731,N_10622);
or U15165 (N_15165,N_10272,N_14644);
nand U15166 (N_15166,N_14540,N_11114);
nand U15167 (N_15167,N_13671,N_12440);
xnor U15168 (N_15168,N_12394,N_13366);
and U15169 (N_15169,N_14037,N_14287);
or U15170 (N_15170,N_10353,N_10520);
and U15171 (N_15171,N_14935,N_13103);
nor U15172 (N_15172,N_14228,N_13607);
xnor U15173 (N_15173,N_10677,N_12265);
and U15174 (N_15174,N_14267,N_11488);
xnor U15175 (N_15175,N_10086,N_14519);
nor U15176 (N_15176,N_14304,N_10975);
nand U15177 (N_15177,N_10651,N_13374);
xor U15178 (N_15178,N_11292,N_12060);
nand U15179 (N_15179,N_14830,N_14545);
and U15180 (N_15180,N_10999,N_14339);
and U15181 (N_15181,N_13410,N_11147);
nor U15182 (N_15182,N_13225,N_11608);
or U15183 (N_15183,N_10901,N_12683);
or U15184 (N_15184,N_10320,N_14338);
nand U15185 (N_15185,N_13561,N_12731);
nor U15186 (N_15186,N_13243,N_11711);
and U15187 (N_15187,N_11151,N_14386);
and U15188 (N_15188,N_13240,N_14297);
xnor U15189 (N_15189,N_11047,N_10652);
nor U15190 (N_15190,N_14885,N_10749);
and U15191 (N_15191,N_12240,N_10123);
and U15192 (N_15192,N_10414,N_12763);
xor U15193 (N_15193,N_13007,N_10594);
nor U15194 (N_15194,N_12283,N_12453);
xnor U15195 (N_15195,N_11816,N_13170);
and U15196 (N_15196,N_12983,N_11253);
nor U15197 (N_15197,N_10299,N_12454);
and U15198 (N_15198,N_14334,N_13344);
nor U15199 (N_15199,N_14213,N_14407);
or U15200 (N_15200,N_11722,N_10052);
and U15201 (N_15201,N_14686,N_11473);
xor U15202 (N_15202,N_11689,N_11491);
nor U15203 (N_15203,N_11215,N_11223);
and U15204 (N_15204,N_14350,N_11221);
nand U15205 (N_15205,N_12628,N_11103);
xor U15206 (N_15206,N_12774,N_13436);
nor U15207 (N_15207,N_14207,N_14342);
nand U15208 (N_15208,N_10175,N_14696);
or U15209 (N_15209,N_14498,N_12470);
and U15210 (N_15210,N_14631,N_14951);
nand U15211 (N_15211,N_10722,N_11217);
xor U15212 (N_15212,N_14225,N_13348);
nand U15213 (N_15213,N_14680,N_11941);
xnor U15214 (N_15214,N_11112,N_13486);
or U15215 (N_15215,N_14955,N_13111);
and U15216 (N_15216,N_12400,N_10680);
xor U15217 (N_15217,N_10268,N_13400);
xnor U15218 (N_15218,N_13144,N_10979);
nand U15219 (N_15219,N_14624,N_12319);
nand U15220 (N_15220,N_11583,N_14013);
nand U15221 (N_15221,N_10806,N_11823);
nand U15222 (N_15222,N_14734,N_13040);
nand U15223 (N_15223,N_13545,N_11386);
xor U15224 (N_15224,N_11731,N_12259);
or U15225 (N_15225,N_10987,N_14903);
and U15226 (N_15226,N_10466,N_10312);
nand U15227 (N_15227,N_13856,N_13207);
xor U15228 (N_15228,N_10025,N_11542);
nor U15229 (N_15229,N_13123,N_11872);
xor U15230 (N_15230,N_12141,N_14060);
and U15231 (N_15231,N_11093,N_13828);
nor U15232 (N_15232,N_11202,N_13334);
nor U15233 (N_15233,N_10203,N_12974);
nor U15234 (N_15234,N_10907,N_13450);
nand U15235 (N_15235,N_11260,N_11159);
or U15236 (N_15236,N_13035,N_13868);
nor U15237 (N_15237,N_13066,N_14871);
xor U15238 (N_15238,N_14124,N_12369);
xor U15239 (N_15239,N_13734,N_13294);
nand U15240 (N_15240,N_14161,N_14751);
or U15241 (N_15241,N_14881,N_12784);
xor U15242 (N_15242,N_12081,N_11050);
xnor U15243 (N_15243,N_12274,N_12068);
nor U15244 (N_15244,N_14893,N_11758);
nor U15245 (N_15245,N_12292,N_14581);
xnor U15246 (N_15246,N_13496,N_13119);
and U15247 (N_15247,N_12431,N_13568);
or U15248 (N_15248,N_13009,N_10475);
or U15249 (N_15249,N_13635,N_13430);
or U15250 (N_15250,N_14957,N_10662);
nand U15251 (N_15251,N_12245,N_13308);
nand U15252 (N_15252,N_13468,N_13335);
and U15253 (N_15253,N_11334,N_10947);
nor U15254 (N_15254,N_13658,N_12813);
nand U15255 (N_15255,N_11232,N_12147);
xnor U15256 (N_15256,N_13790,N_14529);
nor U15257 (N_15257,N_14094,N_10916);
xor U15258 (N_15258,N_14243,N_14969);
xor U15259 (N_15259,N_12834,N_13487);
nand U15260 (N_15260,N_10444,N_13596);
or U15261 (N_15261,N_14741,N_12346);
or U15262 (N_15262,N_12402,N_14112);
and U15263 (N_15263,N_10379,N_13075);
nor U15264 (N_15264,N_10984,N_14198);
or U15265 (N_15265,N_13191,N_11476);
nor U15266 (N_15266,N_13118,N_14544);
and U15267 (N_15267,N_11226,N_14099);
and U15268 (N_15268,N_12381,N_14829);
or U15269 (N_15269,N_10697,N_12507);
xnor U15270 (N_15270,N_10306,N_14925);
nand U15271 (N_15271,N_11383,N_10780);
nor U15272 (N_15272,N_10950,N_12796);
nor U15273 (N_15273,N_13986,N_10213);
and U15274 (N_15274,N_11055,N_11431);
and U15275 (N_15275,N_11769,N_11277);
and U15276 (N_15276,N_12273,N_11924);
nor U15277 (N_15277,N_11977,N_11528);
and U15278 (N_15278,N_14977,N_10187);
xnor U15279 (N_15279,N_11867,N_14577);
nand U15280 (N_15280,N_12609,N_13088);
nor U15281 (N_15281,N_12839,N_13491);
or U15282 (N_15282,N_10706,N_11169);
or U15283 (N_15283,N_12955,N_12106);
nor U15284 (N_15284,N_13085,N_12820);
or U15285 (N_15285,N_13775,N_12786);
or U15286 (N_15286,N_12993,N_14025);
or U15287 (N_15287,N_14598,N_11633);
and U15288 (N_15288,N_13888,N_11460);
and U15289 (N_15289,N_10589,N_14987);
or U15290 (N_15290,N_11620,N_12451);
and U15291 (N_15291,N_12392,N_11650);
or U15292 (N_15292,N_12128,N_14333);
and U15293 (N_15293,N_12627,N_13714);
or U15294 (N_15294,N_13894,N_14516);
nor U15295 (N_15295,N_10801,N_10817);
nand U15296 (N_15296,N_14066,N_13804);
xor U15297 (N_15297,N_14453,N_10497);
or U15298 (N_15298,N_11339,N_10479);
and U15299 (N_15299,N_12539,N_10150);
xnor U15300 (N_15300,N_12735,N_10914);
nor U15301 (N_15301,N_10073,N_13590);
and U15302 (N_15302,N_13095,N_11323);
and U15303 (N_15303,N_11720,N_14147);
nand U15304 (N_15304,N_14578,N_11566);
nor U15305 (N_15305,N_14678,N_14439);
and U15306 (N_15306,N_13772,N_11149);
xnor U15307 (N_15307,N_13379,N_12662);
nand U15308 (N_15308,N_13555,N_12020);
xor U15309 (N_15309,N_11225,N_10454);
nor U15310 (N_15310,N_13606,N_14722);
nor U15311 (N_15311,N_13598,N_11598);
or U15312 (N_15312,N_13628,N_11523);
xor U15313 (N_15313,N_11879,N_12681);
and U15314 (N_15314,N_11182,N_11641);
nand U15315 (N_15315,N_10346,N_12625);
and U15316 (N_15316,N_12586,N_13064);
nor U15317 (N_15317,N_12574,N_11117);
and U15318 (N_15318,N_11581,N_11445);
xnor U15319 (N_15319,N_14058,N_13154);
and U15320 (N_15320,N_11257,N_14814);
nor U15321 (N_15321,N_10282,N_12256);
or U15322 (N_15322,N_11336,N_14675);
xor U15323 (N_15323,N_14752,N_14779);
and U15324 (N_15324,N_11826,N_11265);
nand U15325 (N_15325,N_10679,N_13390);
nor U15326 (N_15326,N_14520,N_12320);
nor U15327 (N_15327,N_12757,N_12503);
or U15328 (N_15328,N_11195,N_14033);
nand U15329 (N_15329,N_12472,N_10787);
xor U15330 (N_15330,N_12776,N_14401);
xnor U15331 (N_15331,N_12385,N_10010);
or U15332 (N_15332,N_13416,N_13425);
nor U15333 (N_15333,N_11560,N_11083);
xnor U15334 (N_15334,N_10014,N_10794);
nor U15335 (N_15335,N_12411,N_14419);
nand U15336 (N_15336,N_14366,N_11596);
xor U15337 (N_15337,N_10932,N_12442);
xnor U15338 (N_15338,N_13630,N_11344);
nand U15339 (N_15339,N_13852,N_14254);
or U15340 (N_15340,N_14588,N_14126);
nor U15341 (N_15341,N_12016,N_12297);
nor U15342 (N_15342,N_10072,N_13543);
nor U15343 (N_15343,N_10683,N_12284);
and U15344 (N_15344,N_14657,N_13472);
or U15345 (N_15345,N_12554,N_11318);
nand U15346 (N_15346,N_13969,N_10020);
and U15347 (N_15347,N_14372,N_13923);
xor U15348 (N_15348,N_11875,N_11110);
nor U15349 (N_15349,N_14477,N_11651);
nor U15350 (N_15350,N_11539,N_13107);
nand U15351 (N_15351,N_11700,N_11041);
nand U15352 (N_15352,N_10954,N_10767);
nand U15353 (N_15353,N_13426,N_14772);
xor U15354 (N_15354,N_13172,N_12428);
and U15355 (N_15355,N_13203,N_13900);
nand U15356 (N_15356,N_11059,N_12349);
xor U15357 (N_15357,N_12498,N_13666);
or U15358 (N_15358,N_11136,N_13873);
xnor U15359 (N_15359,N_13169,N_12759);
nor U15360 (N_15360,N_13909,N_12116);
nand U15361 (N_15361,N_10511,N_10873);
nand U15362 (N_15362,N_12918,N_14807);
or U15363 (N_15363,N_12295,N_14580);
xor U15364 (N_15364,N_12758,N_13947);
nand U15365 (N_15365,N_12333,N_11027);
nand U15366 (N_15366,N_14137,N_11889);
and U15367 (N_15367,N_11124,N_13012);
nand U15368 (N_15368,N_13539,N_12560);
nand U15369 (N_15369,N_11394,N_11004);
nor U15370 (N_15370,N_10935,N_10169);
and U15371 (N_15371,N_10058,N_12315);
xor U15372 (N_15372,N_10388,N_10758);
nor U15373 (N_15373,N_14703,N_10993);
and U15374 (N_15374,N_11247,N_12638);
and U15375 (N_15375,N_14015,N_10019);
and U15376 (N_15376,N_12549,N_10812);
or U15377 (N_15377,N_10131,N_12415);
nand U15378 (N_15378,N_12694,N_14782);
or U15379 (N_15379,N_11834,N_11852);
xnor U15380 (N_15380,N_14156,N_10921);
nand U15381 (N_15381,N_14685,N_13327);
and U15382 (N_15382,N_10524,N_12115);
nor U15383 (N_15383,N_12233,N_14799);
nor U15384 (N_15384,N_10537,N_14396);
nor U15385 (N_15385,N_11130,N_13594);
nor U15386 (N_15386,N_11506,N_10112);
or U15387 (N_15387,N_12216,N_14291);
or U15388 (N_15388,N_10666,N_13319);
or U15389 (N_15389,N_13358,N_13116);
or U15390 (N_15390,N_12952,N_14062);
or U15391 (N_15391,N_13604,N_10887);
and U15392 (N_15392,N_11998,N_12610);
nand U15393 (N_15393,N_11058,N_14172);
nor U15394 (N_15394,N_11453,N_13973);
or U15395 (N_15395,N_14408,N_11557);
nor U15396 (N_15396,N_11554,N_14633);
or U15397 (N_15397,N_14563,N_13741);
nor U15398 (N_15398,N_13381,N_14011);
nand U15399 (N_15399,N_13254,N_10120);
and U15400 (N_15400,N_10724,N_10055);
xnor U15401 (N_15401,N_13299,N_12062);
xnor U15402 (N_15402,N_14226,N_12340);
nor U15403 (N_15403,N_10151,N_12887);
or U15404 (N_15404,N_11125,N_11485);
xnor U15405 (N_15405,N_12288,N_13783);
nand U15406 (N_15406,N_12249,N_12537);
and U15407 (N_15407,N_13503,N_13401);
nor U15408 (N_15408,N_11403,N_12018);
xnor U15409 (N_15409,N_13128,N_12232);
and U15410 (N_15410,N_10326,N_13467);
or U15411 (N_15411,N_12148,N_14629);
nor U15412 (N_15412,N_12738,N_14125);
and U15413 (N_15413,N_12087,N_12634);
nor U15414 (N_15414,N_11870,N_14077);
or U15415 (N_15415,N_13943,N_13456);
and U15416 (N_15416,N_10751,N_12410);
nor U15417 (N_15417,N_13479,N_14845);
or U15418 (N_15418,N_13558,N_10753);
and U15419 (N_15419,N_11229,N_12092);
or U15420 (N_15420,N_14642,N_12122);
nand U15421 (N_15421,N_14316,N_13738);
or U15422 (N_15422,N_13370,N_14709);
xnor U15423 (N_15423,N_12531,N_10658);
xnor U15424 (N_15424,N_11712,N_11196);
xnor U15425 (N_15425,N_14052,N_12407);
and U15426 (N_15426,N_13139,N_13071);
nand U15427 (N_15427,N_12403,N_14433);
nand U15428 (N_15428,N_14239,N_14940);
xor U15429 (N_15429,N_13082,N_13722);
xor U15430 (N_15430,N_10218,N_13073);
xnor U15431 (N_15431,N_11948,N_12978);
nor U15432 (N_15432,N_12773,N_12593);
and U15433 (N_15433,N_13253,N_10202);
and U15434 (N_15434,N_13776,N_14199);
nand U15435 (N_15435,N_12576,N_12963);
or U15436 (N_15436,N_13615,N_11204);
nand U15437 (N_15437,N_13131,N_14791);
xor U15438 (N_15438,N_12721,N_13417);
xor U15439 (N_15439,N_12562,N_12931);
xor U15440 (N_15440,N_11377,N_13580);
nor U15441 (N_15441,N_11814,N_12050);
nand U15442 (N_15442,N_12579,N_12742);
and U15443 (N_15443,N_12640,N_11496);
nor U15444 (N_15444,N_10757,N_11568);
or U15445 (N_15445,N_11550,N_11589);
nand U15446 (N_15446,N_10371,N_14708);
nand U15447 (N_15447,N_12221,N_10583);
xnor U15448 (N_15448,N_11558,N_10243);
xor U15449 (N_15449,N_14390,N_11745);
or U15450 (N_15450,N_11882,N_11611);
xor U15451 (N_15451,N_13142,N_10968);
and U15452 (N_15452,N_13711,N_10124);
nor U15453 (N_15453,N_14170,N_11910);
xnor U15454 (N_15454,N_12005,N_10456);
or U15455 (N_15455,N_13141,N_10316);
or U15456 (N_15456,N_14035,N_10347);
and U15457 (N_15457,N_10976,N_13493);
nor U15458 (N_15458,N_12569,N_13215);
nor U15459 (N_15459,N_14978,N_10489);
and U15460 (N_15460,N_11656,N_10095);
or U15461 (N_15461,N_10703,N_12210);
nor U15462 (N_15462,N_11417,N_14313);
nand U15463 (N_15463,N_10140,N_13091);
nor U15464 (N_15464,N_14510,N_12334);
nor U15465 (N_15465,N_12605,N_14144);
nand U15466 (N_15466,N_11439,N_10641);
xor U15467 (N_15467,N_14394,N_12448);
xor U15468 (N_15468,N_14534,N_11987);
xnor U15469 (N_15469,N_10255,N_14963);
xor U15470 (N_15470,N_13538,N_12207);
nor U15471 (N_15471,N_10366,N_13423);
or U15472 (N_15472,N_12526,N_11508);
xnor U15473 (N_15473,N_11663,N_14204);
and U15474 (N_15474,N_13174,N_13395);
nand U15475 (N_15475,N_10217,N_12473);
and U15476 (N_15476,N_10823,N_10191);
or U15477 (N_15477,N_11753,N_11040);
or U15478 (N_15478,N_10464,N_13886);
and U15479 (N_15479,N_13278,N_10313);
and U15480 (N_15480,N_12485,N_10170);
or U15481 (N_15481,N_11201,N_11770);
nand U15482 (N_15482,N_12809,N_11744);
nor U15483 (N_15483,N_13662,N_10474);
xnor U15484 (N_15484,N_13002,N_10233);
or U15485 (N_15485,N_13277,N_14105);
and U15486 (N_15486,N_13847,N_13026);
nand U15487 (N_15487,N_14719,N_14743);
xor U15488 (N_15488,N_11132,N_12479);
or U15489 (N_15489,N_14479,N_10844);
or U15490 (N_15490,N_13500,N_10593);
or U15491 (N_15491,N_13595,N_10813);
and U15492 (N_15492,N_13901,N_13968);
and U15493 (N_15493,N_10991,N_11760);
and U15494 (N_15494,N_13036,N_13418);
and U15495 (N_15495,N_14616,N_13816);
nor U15496 (N_15496,N_11224,N_13385);
and U15497 (N_15497,N_10000,N_12460);
xnor U15498 (N_15498,N_14068,N_10398);
xnor U15499 (N_15499,N_10851,N_11121);
and U15500 (N_15500,N_12644,N_13382);
nor U15501 (N_15501,N_10078,N_13420);
or U15502 (N_15502,N_10458,N_14377);
nand U15503 (N_15503,N_14494,N_11212);
or U15504 (N_15504,N_11274,N_12868);
xor U15505 (N_15505,N_12775,N_11974);
xor U15506 (N_15506,N_10676,N_12849);
or U15507 (N_15507,N_13213,N_10113);
nor U15508 (N_15508,N_12769,N_10937);
nand U15509 (N_15509,N_13867,N_10973);
and U15510 (N_15510,N_11701,N_13183);
and U15511 (N_15511,N_11694,N_10635);
nand U15512 (N_15512,N_13740,N_11348);
or U15513 (N_15513,N_12728,N_13667);
xnor U15514 (N_15514,N_11773,N_11380);
nor U15515 (N_15515,N_12672,N_12746);
or U15516 (N_15516,N_13232,N_10704);
nor U15517 (N_15517,N_14549,N_14224);
or U15518 (N_15518,N_13175,N_11997);
nor U15519 (N_15519,N_14937,N_12246);
or U15520 (N_15520,N_14659,N_11016);
and U15521 (N_15521,N_10111,N_10013);
and U15522 (N_15522,N_14527,N_10892);
xor U15523 (N_15523,N_14950,N_14662);
or U15524 (N_15524,N_12269,N_10063);
nand U15525 (N_15525,N_13527,N_13041);
or U15526 (N_15526,N_11137,N_13899);
nor U15527 (N_15527,N_12900,N_12919);
xor U15528 (N_15528,N_13678,N_13245);
nor U15529 (N_15529,N_11404,N_13835);
nand U15530 (N_15530,N_11599,N_10167);
or U15531 (N_15531,N_12570,N_13526);
nor U15532 (N_15532,N_14054,N_12906);
xnor U15533 (N_15533,N_11762,N_13368);
and U15534 (N_15534,N_14299,N_10792);
and U15535 (N_15535,N_14626,N_14295);
and U15536 (N_15536,N_10895,N_11119);
or U15537 (N_15537,N_14018,N_10532);
nor U15538 (N_15538,N_11461,N_14801);
or U15539 (N_15539,N_10295,N_13958);
or U15540 (N_15540,N_10036,N_14508);
nor U15541 (N_15541,N_11302,N_12152);
nand U15542 (N_15542,N_11077,N_10105);
or U15543 (N_15543,N_10488,N_11714);
or U15544 (N_15544,N_11122,N_13309);
nor U15545 (N_15545,N_11774,N_13336);
xnor U15546 (N_15546,N_12523,N_13811);
nor U15547 (N_15547,N_11134,N_11310);
and U15548 (N_15548,N_13540,N_13946);
and U15549 (N_15549,N_11288,N_13771);
xor U15550 (N_15550,N_11315,N_13011);
or U15551 (N_15551,N_14431,N_13865);
or U15552 (N_15552,N_11727,N_13434);
and U15553 (N_15553,N_13570,N_14864);
nand U15554 (N_15554,N_12097,N_13898);
or U15555 (N_15555,N_13853,N_14215);
or U15556 (N_15556,N_13442,N_10143);
or U15557 (N_15557,N_12012,N_14067);
and U15558 (N_15558,N_13349,N_13480);
and U15559 (N_15559,N_14100,N_12612);
nand U15560 (N_15560,N_12059,N_12165);
and U15561 (N_15561,N_12733,N_14012);
and U15562 (N_15562,N_12484,N_12489);
nor U15563 (N_15563,N_11899,N_10556);
nor U15564 (N_15564,N_11734,N_12399);
or U15565 (N_15565,N_14748,N_12700);
nand U15566 (N_15566,N_10875,N_12604);
and U15567 (N_15567,N_12622,N_13777);
xnor U15568 (N_15568,N_10994,N_14182);
nor U15569 (N_15569,N_14276,N_14117);
nor U15570 (N_15570,N_12575,N_12267);
or U15571 (N_15571,N_12513,N_12716);
and U15572 (N_15572,N_14497,N_13102);
nand U15573 (N_15573,N_10485,N_14245);
or U15574 (N_15574,N_10917,N_11886);
nand U15575 (N_15575,N_11674,N_10436);
xor U15576 (N_15576,N_14818,N_14021);
nand U15577 (N_15577,N_13206,N_11634);
xor U15578 (N_15578,N_14973,N_11422);
nor U15579 (N_15579,N_11002,N_10746);
and U15580 (N_15580,N_12764,N_10739);
or U15581 (N_15581,N_13341,N_10374);
and U15582 (N_15582,N_12129,N_13072);
xor U15583 (N_15583,N_10495,N_11325);
nor U15584 (N_15584,N_10848,N_14038);
or U15585 (N_15585,N_11824,N_14777);
or U15586 (N_15586,N_12862,N_10734);
xor U15587 (N_15587,N_10995,N_12907);
nor U15588 (N_15588,N_13557,N_14548);
and U15589 (N_15589,N_12635,N_14106);
or U15590 (N_15590,N_11305,N_11725);
nor U15591 (N_15591,N_13997,N_13469);
nand U15592 (N_15592,N_11777,N_11167);
xnor U15593 (N_15593,N_13838,N_12413);
and U15594 (N_15594,N_10546,N_14417);
nor U15595 (N_15595,N_12200,N_13525);
nor U15596 (N_15596,N_13399,N_10165);
xor U15597 (N_15597,N_14046,N_11618);
or U15598 (N_15598,N_11458,N_13930);
nand U15599 (N_15599,N_12387,N_14848);
nand U15600 (N_15600,N_10669,N_13252);
nand U15601 (N_15601,N_10236,N_11005);
or U15602 (N_15602,N_14261,N_13952);
or U15603 (N_15603,N_10235,N_11984);
or U15604 (N_15604,N_10082,N_10412);
xnor U15605 (N_15605,N_12368,N_11682);
and U15606 (N_15606,N_14838,N_11779);
nand U15607 (N_15607,N_13286,N_11230);
or U15608 (N_15608,N_10118,N_14044);
xor U15609 (N_15609,N_12171,N_14668);
and U15610 (N_15610,N_12217,N_11423);
nand U15611 (N_15611,N_12094,N_12028);
or U15612 (N_15612,N_11942,N_13851);
or U15613 (N_15613,N_12951,N_14788);
or U15614 (N_15614,N_12755,N_13196);
nand U15615 (N_15615,N_11893,N_13941);
nand U15616 (N_15616,N_10031,N_10804);
or U15617 (N_15617,N_14331,N_10431);
and U15618 (N_15618,N_11014,N_14173);
and U15619 (N_15619,N_12379,N_11971);
and U15620 (N_15620,N_10279,N_12751);
or U15621 (N_15621,N_12780,N_12098);
xor U15622 (N_15622,N_14842,N_12139);
nand U15623 (N_15623,N_10933,N_11415);
xnor U15624 (N_15624,N_11820,N_11751);
nand U15625 (N_15625,N_11475,N_13179);
nor U15626 (N_15626,N_14584,N_12916);
nor U15627 (N_15627,N_13610,N_14841);
and U15628 (N_15628,N_13951,N_13003);
nor U15629 (N_15629,N_10309,N_11029);
xor U15630 (N_15630,N_13143,N_12666);
nand U15631 (N_15631,N_10447,N_13427);
nor U15632 (N_15632,N_14070,N_13751);
xor U15633 (N_15633,N_11054,N_10700);
xnor U15634 (N_15634,N_11975,N_13640);
xnor U15635 (N_15635,N_14769,N_11053);
or U15636 (N_15636,N_10231,N_14958);
xnor U15637 (N_15637,N_10463,N_13643);
and U15638 (N_15638,N_13097,N_11294);
or U15639 (N_15639,N_14906,N_13398);
or U15640 (N_15640,N_11790,N_11089);
xor U15641 (N_15641,N_11032,N_14491);
or U15642 (N_15642,N_13431,N_11430);
and U15643 (N_15643,N_14606,N_11275);
nor U15644 (N_15644,N_11063,N_11595);
xnor U15645 (N_15645,N_10329,N_12328);
xnor U15646 (N_15646,N_10693,N_10501);
or U15647 (N_15647,N_11812,N_13814);
and U15648 (N_15648,N_13217,N_11843);
and U15649 (N_15649,N_13386,N_12244);
nand U15650 (N_15650,N_14525,N_14427);
and U15651 (N_15651,N_12515,N_12691);
nand U15652 (N_15652,N_10835,N_10939);
xor U15653 (N_15653,N_13077,N_11360);
and U15654 (N_15654,N_11705,N_10001);
nor U15655 (N_15655,N_11237,N_11100);
xor U15656 (N_15656,N_12633,N_13755);
nor U15657 (N_15657,N_11990,N_11704);
xor U15658 (N_15658,N_13942,N_13490);
nand U15659 (N_15659,N_12312,N_12581);
or U15660 (N_15660,N_10530,N_13933);
xor U15661 (N_15661,N_13831,N_11443);
or U15662 (N_15662,N_14728,N_10983);
and U15663 (N_15663,N_10837,N_12159);
and U15664 (N_15664,N_13698,N_12182);
xor U15665 (N_15665,N_12715,N_12354);
xor U15666 (N_15666,N_12228,N_14822);
nor U15667 (N_15667,N_12031,N_14613);
nor U15668 (N_15668,N_10971,N_14042);
or U15669 (N_15669,N_11979,N_14552);
nand U15670 (N_15670,N_14846,N_12982);
and U15671 (N_15671,N_13818,N_14914);
nand U15672 (N_15672,N_10049,N_10109);
nor U15673 (N_15673,N_14159,N_12971);
and U15674 (N_15674,N_12261,N_10610);
and U15675 (N_15675,N_14379,N_11181);
nand U15676 (N_15676,N_12941,N_11081);
and U15677 (N_15677,N_11825,N_13383);
or U15678 (N_15678,N_12926,N_13145);
xnor U15679 (N_15679,N_10864,N_10876);
and U15680 (N_15680,N_10323,N_14392);
and U15681 (N_15681,N_12777,N_12287);
nor U15682 (N_15682,N_13415,N_14513);
or U15683 (N_15683,N_10372,N_14264);
or U15684 (N_15684,N_14660,N_11524);
xnor U15685 (N_15685,N_14773,N_13193);
xor U15686 (N_15686,N_12817,N_11177);
nand U15687 (N_15687,N_10208,N_14423);
and U15688 (N_15688,N_12254,N_10145);
nor U15689 (N_15689,N_13984,N_13140);
xnor U15690 (N_15690,N_14171,N_10465);
nor U15691 (N_15691,N_12917,N_14887);
nand U15692 (N_15692,N_10507,N_14302);
and U15693 (N_15693,N_12641,N_11805);
and U15694 (N_15694,N_12441,N_12865);
xor U15695 (N_15695,N_10059,N_10331);
nand U15696 (N_15696,N_10376,N_12891);
nand U15697 (N_15697,N_12760,N_13029);
or U15698 (N_15698,N_13817,N_11635);
and U15699 (N_15699,N_11208,N_14165);
xnor U15700 (N_15700,N_10996,N_12490);
xor U15701 (N_15701,N_14189,N_14564);
or U15702 (N_15702,N_12421,N_14652);
and U15703 (N_15703,N_11308,N_13651);
xor U15704 (N_15704,N_10108,N_12447);
xnor U15705 (N_15705,N_12127,N_13634);
nand U15706 (N_15706,N_14092,N_13993);
nand U15707 (N_15707,N_14493,N_12191);
or U15708 (N_15708,N_12508,N_11389);
or U15709 (N_15709,N_12973,N_14713);
nand U15710 (N_15710,N_11536,N_12799);
nor U15711 (N_15711,N_10433,N_10928);
and U15712 (N_15712,N_12239,N_11233);
xnor U15713 (N_15713,N_14118,N_13550);
nor U15714 (N_15714,N_14006,N_13633);
and U15715 (N_15715,N_10654,N_12690);
nand U15716 (N_15716,N_13275,N_12876);
nand U15717 (N_15717,N_11838,N_14457);
nand U15718 (N_15718,N_11152,N_13194);
or U15719 (N_15719,N_10012,N_12550);
or U15720 (N_15720,N_12036,N_14847);
nand U15721 (N_15721,N_14266,N_10847);
or U15722 (N_15722,N_11433,N_11660);
nor U15723 (N_15723,N_11555,N_13209);
xor U15724 (N_15724,N_11118,N_13670);
nand U15725 (N_15725,N_12276,N_14387);
nor U15726 (N_15726,N_11576,N_10425);
or U15727 (N_15727,N_11388,N_14892);
nand U15728 (N_15728,N_12538,N_12859);
xnor U15729 (N_15729,N_14535,N_12992);
nand U15730 (N_15730,N_14942,N_10855);
or U15731 (N_15731,N_12166,N_13877);
nor U15732 (N_15732,N_11500,N_14323);
nor U15733 (N_15733,N_12826,N_12305);
nor U15734 (N_15734,N_12822,N_13284);
nand U15735 (N_15735,N_14908,N_13820);
nand U15736 (N_15736,N_12882,N_11462);
nand U15737 (N_15737,N_13907,N_12603);
nor U15738 (N_15738,N_14900,N_11094);
and U15739 (N_15739,N_10732,N_10889);
or U15740 (N_15740,N_14991,N_11026);
or U15741 (N_15741,N_12177,N_10317);
nor U15742 (N_15742,N_13612,N_14770);
xnor U15743 (N_15743,N_11090,N_10384);
xnor U15744 (N_15744,N_11076,N_11730);
and U15745 (N_15745,N_12435,N_10843);
xnor U15746 (N_15746,N_11395,N_10091);
and U15747 (N_15747,N_14998,N_14180);
nor U15748 (N_15748,N_13057,N_10280);
nand U15749 (N_15749,N_14840,N_14487);
xnor U15750 (N_15750,N_11003,N_14233);
or U15751 (N_15751,N_12383,N_12511);
or U15752 (N_15752,N_13298,N_10419);
or U15753 (N_15753,N_13642,N_12035);
xor U15754 (N_15754,N_13134,N_14461);
and U15755 (N_15755,N_14113,N_12222);
xnor U15756 (N_15756,N_10561,N_13915);
and U15757 (N_15757,N_13402,N_10591);
or U15758 (N_15758,N_13623,N_12125);
and U15759 (N_15759,N_11411,N_13602);
and U15760 (N_15760,N_10064,N_11548);
or U15761 (N_15761,N_13101,N_12494);
xor U15762 (N_15762,N_14835,N_14674);
xor U15763 (N_15763,N_10502,N_12850);
or U15764 (N_15764,N_12121,N_10784);
xor U15765 (N_15765,N_10098,N_13043);
and U15766 (N_15766,N_11409,N_10023);
or U15767 (N_15767,N_10961,N_12818);
or U15768 (N_15768,N_11290,N_14532);
xor U15769 (N_15769,N_14271,N_13446);
nor U15770 (N_15770,N_13684,N_13473);
or U15771 (N_15771,N_11494,N_11818);
nor U15772 (N_15772,N_10931,N_10789);
or U15773 (N_15773,N_13911,N_10125);
nand U15774 (N_15774,N_13726,N_11952);
and U15775 (N_15775,N_12432,N_13027);
or U15776 (N_15776,N_14539,N_12162);
nand U15777 (N_15777,N_13000,N_13957);
nand U15778 (N_15778,N_12266,N_11600);
nor U15779 (N_15779,N_11418,N_14321);
xnor U15780 (N_15780,N_10585,N_12105);
nor U15781 (N_15781,N_12280,N_11908);
xnor U15782 (N_15782,N_14443,N_14726);
xor U15783 (N_15783,N_11776,N_12466);
xnor U15784 (N_15784,N_10469,N_12401);
xnor U15785 (N_15785,N_10853,N_14915);
and U15786 (N_15786,N_10275,N_10178);
or U15787 (N_15787,N_12022,N_12542);
or U15788 (N_15788,N_13312,N_12190);
or U15789 (N_15789,N_11345,N_11477);
xor U15790 (N_15790,N_13874,N_11578);
and U15791 (N_15791,N_10154,N_14000);
nand U15792 (N_15792,N_10756,N_14882);
nand U15793 (N_15793,N_10476,N_11470);
and U15794 (N_15794,N_14087,N_11570);
xor U15795 (N_15795,N_14677,N_14257);
or U15796 (N_15796,N_12670,N_13972);
nor U15797 (N_15797,N_14194,N_10692);
or U15798 (N_15798,N_12188,N_13222);
xor U15799 (N_15799,N_10083,N_10702);
and U15800 (N_15800,N_11988,N_13347);
or U15801 (N_15801,N_10605,N_10825);
or U15802 (N_15802,N_12307,N_10430);
nand U15803 (N_15803,N_10088,N_11173);
or U15804 (N_15804,N_14877,N_12795);
xnor U15805 (N_15805,N_10333,N_13249);
or U15806 (N_15806,N_14305,N_11531);
or U15807 (N_15807,N_10400,N_12172);
nor U15808 (N_15808,N_11116,N_13301);
and U15809 (N_15809,N_13843,N_13989);
or U15810 (N_15810,N_12598,N_14114);
nor U15811 (N_15811,N_11537,N_12255);
and U15812 (N_15812,N_12645,N_14242);
nand U15813 (N_15813,N_10397,N_10421);
nand U15814 (N_15814,N_10516,N_14970);
and U15815 (N_15815,N_11803,N_10363);
nand U15816 (N_15816,N_11115,N_14993);
or U15817 (N_15817,N_13444,N_12492);
or U15818 (N_15818,N_13728,N_13127);
and U15819 (N_15819,N_13914,N_13862);
or U15820 (N_15820,N_12879,N_12732);
nor U15821 (N_15821,N_11263,N_12377);
xor U15822 (N_15822,N_11780,N_10342);
xor U15823 (N_15823,N_13457,N_10077);
xor U15824 (N_15824,N_11813,N_14965);
and U15825 (N_15825,N_12946,N_10663);
xor U15826 (N_15826,N_14530,N_14047);
nor U15827 (N_15827,N_11028,N_13251);
xnor U15828 (N_15828,N_10087,N_10417);
and U15829 (N_15829,N_14084,N_12160);
nor U15830 (N_15830,N_12717,N_12113);
or U15831 (N_15831,N_14802,N_13971);
nand U15832 (N_15832,N_11698,N_14715);
or U15833 (N_15833,N_13455,N_10810);
and U15834 (N_15834,N_13476,N_13995);
or U15835 (N_15835,N_10214,N_12649);
or U15836 (N_15836,N_10321,N_13044);
xor U15837 (N_15837,N_11193,N_12224);
or U15838 (N_15838,N_14475,N_14651);
or U15839 (N_15839,N_10547,N_14932);
or U15840 (N_15840,N_14797,N_10802);
and U15841 (N_15841,N_10718,N_12707);
or U15842 (N_15842,N_11798,N_11880);
xnor U15843 (N_15843,N_10906,N_13182);
nand U15844 (N_15844,N_10100,N_12391);
xor U15845 (N_15845,N_13660,N_10179);
nand U15846 (N_15846,N_12922,N_10761);
xnor U15847 (N_15847,N_13184,N_10736);
nand U15848 (N_15848,N_10490,N_10365);
or U15849 (N_15849,N_13195,N_11833);
nand U15850 (N_15850,N_11171,N_14628);
nand U15851 (N_15851,N_12578,N_12838);
nand U15852 (N_15852,N_10539,N_10584);
or U15853 (N_15853,N_13202,N_14110);
nand U15854 (N_15854,N_11652,N_10879);
and U15855 (N_15855,N_11018,N_11691);
or U15856 (N_15856,N_13006,N_10778);
nand U15857 (N_15857,N_11587,N_13577);
nor U15858 (N_15858,N_12712,N_13629);
and U15859 (N_15859,N_13210,N_14711);
nor U15860 (N_15860,N_13528,N_10822);
xnor U15861 (N_15861,N_14982,N_11512);
nor U15862 (N_15862,N_11715,N_13345);
and U15863 (N_15863,N_10903,N_14833);
or U15864 (N_15864,N_10199,N_10897);
xor U15865 (N_15865,N_11437,N_13322);
nor U15866 (N_15866,N_13836,N_14634);
xor U15867 (N_15867,N_14910,N_13745);
nand U15868 (N_15868,N_14188,N_13181);
nor U15869 (N_15869,N_14853,N_14059);
nand U15870 (N_15870,N_10311,N_12651);
and U15871 (N_15871,N_13964,N_13547);
xnor U15872 (N_15872,N_11920,N_11795);
nor U15873 (N_15873,N_11398,N_14538);
and U15874 (N_15874,N_14617,N_13793);
or U15875 (N_15875,N_11206,N_12657);
and U15876 (N_15876,N_11513,N_12797);
nand U15877 (N_15877,N_13316,N_14579);
and U15878 (N_15878,N_10925,N_11836);
or U15879 (N_15879,N_13677,N_11414);
nand U15880 (N_15880,N_14438,N_13679);
xor U15881 (N_15881,N_14650,N_13622);
or U15882 (N_15882,N_14464,N_13774);
nand U15883 (N_15883,N_10467,N_13659);
and U15884 (N_15884,N_14346,N_13905);
nor U15885 (N_15885,N_12464,N_12968);
and U15886 (N_15886,N_10158,N_12268);
xor U15887 (N_15887,N_12861,N_11896);
xor U15888 (N_15888,N_14690,N_13566);
nand U15889 (N_15889,N_10318,N_11939);
nand U15890 (N_15890,N_11351,N_12047);
and U15891 (N_15891,N_11111,N_11510);
xor U15892 (N_15892,N_11784,N_12723);
or U15893 (N_15893,N_12564,N_13165);
or U15894 (N_15894,N_12371,N_10011);
nand U15895 (N_15895,N_13511,N_10529);
or U15896 (N_15896,N_13034,N_11420);
nor U15897 (N_15897,N_14619,N_12630);
nor U15898 (N_15898,N_13784,N_12737);
or U15899 (N_15899,N_10182,N_10531);
nand U15900 (N_15900,N_11654,N_14274);
nor U15901 (N_15901,N_11241,N_14216);
and U15902 (N_15902,N_12989,N_13236);
and U15903 (N_15903,N_14088,N_10668);
xnor U15904 (N_15904,N_12123,N_14886);
xor U15905 (N_15905,N_12696,N_14463);
nand U15906 (N_15906,N_11038,N_14129);
and U15907 (N_15907,N_14120,N_11817);
nand U15908 (N_15908,N_14878,N_11393);
or U15909 (N_15909,N_12133,N_11366);
xor U15910 (N_15910,N_11168,N_11096);
or U15911 (N_15911,N_12041,N_10936);
and U15912 (N_15912,N_10341,N_12112);
nand U15913 (N_15913,N_13788,N_12516);
xnor U15914 (N_15914,N_13956,N_14139);
xor U15915 (N_15915,N_14195,N_12013);
nand U15916 (N_15916,N_10160,N_12532);
or U15917 (N_15917,N_12661,N_13013);
nand U15918 (N_15918,N_13342,N_13371);
nand U15919 (N_15919,N_14284,N_12238);
nor U15920 (N_15920,N_14562,N_12821);
or U15921 (N_15921,N_14057,N_10173);
and U15922 (N_15922,N_13153,N_13541);
nand U15923 (N_15923,N_10965,N_13069);
nand U15924 (N_15924,N_10305,N_11543);
and U15925 (N_15925,N_11082,N_13171);
or U15926 (N_15926,N_11703,N_14611);
or U15927 (N_15927,N_14936,N_12743);
and U15928 (N_15928,N_11056,N_13248);
xnor U15929 (N_15929,N_12117,N_13884);
xnor U15930 (N_15930,N_12990,N_13198);
or U15931 (N_15931,N_13564,N_10249);
or U15932 (N_15932,N_12924,N_13405);
and U15933 (N_15933,N_14698,N_14612);
nor U15934 (N_15934,N_12135,N_12830);
xnor U15935 (N_15935,N_12084,N_14614);
xnor U15936 (N_15936,N_10021,N_11677);
or U15937 (N_15937,N_12730,N_14312);
and U15938 (N_15938,N_14808,N_12877);
or U15939 (N_15939,N_14505,N_14868);
xnor U15940 (N_15940,N_12913,N_10428);
and U15941 (N_15941,N_10508,N_11933);
or U15942 (N_15942,N_13988,N_14856);
nand U15943 (N_15943,N_11574,N_10811);
and U15944 (N_15944,N_13311,N_10290);
and U15945 (N_15945,N_10707,N_12524);
nand U15946 (N_15946,N_11713,N_12998);
xor U15947 (N_15947,N_10302,N_10527);
nand U15948 (N_15948,N_10966,N_11179);
or U15949 (N_15949,N_14896,N_12389);
nor U15950 (N_15950,N_12465,N_13185);
or U15951 (N_15951,N_11350,N_14481);
nor U15952 (N_15952,N_10915,N_12972);
nor U15953 (N_15953,N_11917,N_14912);
nor U15954 (N_15954,N_14721,N_10609);
or U15955 (N_15955,N_10192,N_13051);
nand U15956 (N_15956,N_12299,N_10974);
nand U15957 (N_15957,N_10481,N_14451);
or U15958 (N_15958,N_14550,N_13720);
xor U15959 (N_15959,N_10242,N_12520);
or U15960 (N_15960,N_13282,N_13289);
and U15961 (N_15961,N_10368,N_12201);
nand U15962 (N_15962,N_11874,N_14689);
and U15963 (N_15963,N_10521,N_13742);
or U15964 (N_15964,N_10616,N_10568);
or U15965 (N_15965,N_10790,N_11091);
or U15966 (N_15966,N_13789,N_14270);
nand U15967 (N_15967,N_14424,N_12279);
nand U15968 (N_15968,N_10750,N_11128);
and U15969 (N_15969,N_10215,N_10029);
nor U15970 (N_15970,N_10478,N_10034);
nor U15971 (N_15971,N_10060,N_13477);
xor U15972 (N_15972,N_12071,N_14554);
nor U15973 (N_15973,N_13021,N_13008);
and U15974 (N_15974,N_10891,N_10278);
and U15975 (N_15975,N_10473,N_12970);
or U15976 (N_15976,N_11307,N_10390);
and U15977 (N_15977,N_12709,N_11909);
xor U15978 (N_15978,N_11486,N_10606);
nor U15979 (N_15979,N_11678,N_13609);
xnor U15980 (N_15980,N_11490,N_10611);
nor U15981 (N_15981,N_14462,N_11764);
and U15982 (N_15982,N_12236,N_14671);
nand U15983 (N_15983,N_14474,N_12078);
and U15984 (N_15984,N_13979,N_14559);
nand U15985 (N_15985,N_11586,N_12163);
xor U15986 (N_15986,N_10107,N_14349);
nand U15987 (N_15987,N_14414,N_14478);
or U15988 (N_15988,N_14700,N_13639);
and U15989 (N_15989,N_13376,N_10614);
xor U15990 (N_15990,N_13392,N_13721);
xor U15991 (N_15991,N_12608,N_10543);
or U15992 (N_15992,N_10037,N_10558);
nand U15993 (N_15993,N_14500,N_10457);
or U15994 (N_15994,N_12293,N_13648);
xor U15995 (N_15995,N_11381,N_10310);
and U15996 (N_15996,N_10271,N_12803);
xor U15997 (N_15997,N_13809,N_13834);
nor U15998 (N_15998,N_12476,N_10735);
xor U15999 (N_15999,N_10084,N_11174);
and U16000 (N_16000,N_12655,N_10477);
and U16001 (N_16001,N_14975,N_13166);
nand U16002 (N_16002,N_14605,N_14898);
nand U16003 (N_16003,N_11363,N_13499);
or U16004 (N_16004,N_10200,N_12915);
and U16005 (N_16005,N_13974,N_14511);
xor U16006 (N_16006,N_13925,N_14640);
or U16007 (N_16007,N_10902,N_11397);
xnor U16008 (N_16008,N_13146,N_14014);
or U16009 (N_16009,N_10824,N_10207);
and U16010 (N_16010,N_14758,N_13762);
and U16011 (N_16011,N_14318,N_13129);
or U16012 (N_16012,N_12705,N_12406);
nor U16013 (N_16013,N_11765,N_12164);
nand U16014 (N_16014,N_14999,N_11109);
or U16015 (N_16015,N_11749,N_11295);
nor U16016 (N_16016,N_11994,N_10162);
nor U16017 (N_16017,N_11865,N_11186);
xnor U16018 (N_16018,N_10800,N_14027);
or U16019 (N_16019,N_12710,N_10166);
or U16020 (N_16020,N_11250,N_14962);
nand U16021 (N_16021,N_12687,N_11535);
xor U16022 (N_16022,N_12487,N_11876);
xor U16023 (N_16023,N_11748,N_12119);
xnor U16024 (N_16024,N_10090,N_13132);
xnor U16025 (N_16025,N_11419,N_14533);
and U16026 (N_16026,N_12819,N_13305);
nor U16027 (N_16027,N_12345,N_11726);
nor U16028 (N_16028,N_14076,N_14263);
xnor U16029 (N_16029,N_10590,N_10328);
and U16030 (N_16030,N_11162,N_10572);
or U16031 (N_16031,N_10336,N_10450);
or U16032 (N_16032,N_10694,N_11203);
nand U16033 (N_16033,N_13825,N_12547);
nor U16034 (N_16034,N_13204,N_11471);
nor U16035 (N_16035,N_10462,N_14388);
or U16036 (N_16036,N_12429,N_12218);
xnor U16037 (N_16037,N_10894,N_10699);
or U16038 (N_16038,N_12535,N_13149);
or U16039 (N_16039,N_10147,N_13042);
nand U16040 (N_16040,N_10988,N_13530);
xor U16041 (N_16041,N_12220,N_12837);
nand U16042 (N_16042,N_11238,N_12197);
and U16043 (N_16043,N_10541,N_12021);
xor U16044 (N_16044,N_13730,N_10455);
nor U16045 (N_16045,N_11068,N_11626);
nand U16046 (N_16046,N_14941,N_11424);
nand U16047 (N_16047,N_13891,N_12533);
and U16048 (N_16048,N_11986,N_10197);
nand U16049 (N_16049,N_13124,N_11509);
or U16050 (N_16050,N_10634,N_14184);
nand U16051 (N_16051,N_14445,N_14043);
xnor U16052 (N_16052,N_10386,N_14214);
or U16053 (N_16053,N_11480,N_14916);
and U16054 (N_16054,N_12675,N_12703);
or U16055 (N_16055,N_14804,N_11261);
and U16056 (N_16056,N_13724,N_10325);
nand U16057 (N_16057,N_13650,N_13826);
or U16058 (N_16058,N_10373,N_14926);
and U16059 (N_16059,N_10057,N_10446);
nor U16060 (N_16060,N_10958,N_14041);
xnor U16061 (N_16061,N_12607,N_11436);
nor U16062 (N_16062,N_14222,N_11919);
xor U16063 (N_16063,N_13556,N_14237);
or U16064 (N_16064,N_10126,N_13463);
nand U16065 (N_16065,N_12504,N_14310);
nand U16066 (N_16066,N_14750,N_11895);
nor U16067 (N_16067,N_10856,N_10785);
and U16068 (N_16068,N_13737,N_12205);
or U16069 (N_16069,N_12405,N_10096);
nor U16070 (N_16070,N_11283,N_11989);
nand U16071 (N_16071,N_11754,N_13151);
nor U16072 (N_16072,N_11172,N_12996);
nand U16073 (N_16073,N_12702,N_11333);
nor U16074 (N_16074,N_14691,N_10544);
and U16075 (N_16075,N_11092,N_11741);
or U16076 (N_16076,N_13338,N_10266);
and U16077 (N_16077,N_14985,N_12706);
nand U16078 (N_16078,N_11428,N_11868);
and U16079 (N_16079,N_11036,N_14767);
or U16080 (N_16080,N_14413,N_13673);
or U16081 (N_16081,N_13459,N_14335);
and U16082 (N_16082,N_13122,N_11140);
and U16083 (N_16083,N_13350,N_10550);
nand U16084 (N_16084,N_14030,N_10453);
nand U16085 (N_16085,N_10809,N_10868);
and U16086 (N_16086,N_10413,N_13162);
or U16087 (N_16087,N_10858,N_11544);
and U16088 (N_16088,N_12984,N_10862);
xnor U16089 (N_16089,N_13552,N_13384);
or U16090 (N_16090,N_10567,N_13023);
nand U16091 (N_16091,N_11695,N_14260);
or U16092 (N_16092,N_12506,N_11216);
or U16093 (N_16093,N_14319,N_13159);
or U16094 (N_16094,N_13584,N_12885);
nor U16095 (N_16095,N_14315,N_14490);
or U16096 (N_16096,N_12138,N_14625);
nand U16097 (N_16097,N_10959,N_12577);
nor U16098 (N_16098,N_10441,N_10038);
and U16099 (N_16099,N_13542,N_10051);
xnor U16100 (N_16100,N_12741,N_14655);
xnor U16101 (N_16101,N_12910,N_12901);
nand U16102 (N_16102,N_10650,N_12816);
and U16103 (N_16103,N_10636,N_12303);
or U16104 (N_16104,N_13587,N_11160);
xnor U16105 (N_16105,N_13296,N_10137);
nand U16106 (N_16106,N_11602,N_13304);
nor U16107 (N_16107,N_10212,N_11789);
nand U16108 (N_16108,N_13844,N_10405);
xnor U16109 (N_16109,N_14278,N_11286);
or U16110 (N_16110,N_10819,N_11010);
nand U16111 (N_16111,N_10513,N_12828);
nand U16112 (N_16112,N_11218,N_11969);
nor U16113 (N_16113,N_13978,N_13032);
nand U16114 (N_16114,N_11097,N_13419);
xor U16115 (N_16115,N_13690,N_11401);
and U16116 (N_16116,N_10184,N_14669);
xor U16117 (N_16117,N_10181,N_13237);
and U16118 (N_16118,N_14705,N_10340);
nand U16119 (N_16119,N_12080,N_13976);
nand U16120 (N_16120,N_14729,N_12736);
or U16121 (N_16121,N_14567,N_12920);
xnor U16122 (N_16122,N_10239,N_10257);
xor U16123 (N_16123,N_12791,N_13155);
or U16124 (N_16124,N_10670,N_11207);
nand U16125 (N_16125,N_12419,N_14072);
or U16126 (N_16126,N_14308,N_13918);
nor U16127 (N_16127,N_10332,N_11540);
and U16128 (N_16128,N_12477,N_14558);
nand U16129 (N_16129,N_13796,N_11850);
xnor U16130 (N_16130,N_11787,N_12663);
xor U16131 (N_16131,N_12697,N_12278);
nand U16132 (N_16132,N_12914,N_11304);
nand U16133 (N_16133,N_12063,N_13870);
nand U16134 (N_16134,N_13068,N_10952);
nand U16135 (N_16135,N_11291,N_10256);
and U16136 (N_16136,N_10141,N_12615);
nor U16137 (N_16137,N_10733,N_11767);
and U16138 (N_16138,N_14503,N_10253);
and U16139 (N_16139,N_14397,N_11187);
nor U16140 (N_16140,N_13180,N_12815);
nand U16141 (N_16141,N_10512,N_10882);
xnor U16142 (N_16142,N_13765,N_12842);
xor U16143 (N_16143,N_14587,N_12378);
xor U16144 (N_16144,N_10818,N_12438);
and U16145 (N_16145,N_10076,N_10044);
and U16146 (N_16146,N_12469,N_12987);
xnor U16147 (N_16147,N_14193,N_11362);
or U16148 (N_16148,N_12252,N_13513);
xor U16149 (N_16149,N_12618,N_14586);
xor U16150 (N_16150,N_14695,N_13962);
nor U16151 (N_16151,N_14905,N_11648);
xor U16152 (N_16152,N_14537,N_10406);
or U16153 (N_16153,N_11514,N_14575);
or U16154 (N_16154,N_11945,N_13273);
and U16155 (N_16155,N_14190,N_13451);
xnor U16156 (N_16156,N_14602,N_11929);
xnor U16157 (N_16157,N_12977,N_13955);
or U16158 (N_16158,N_12234,N_14492);
and U16159 (N_16159,N_10033,N_10432);
nor U16160 (N_16160,N_12840,N_14980);
and U16161 (N_16161,N_14395,N_14368);
nor U16162 (N_16162,N_10429,N_13234);
xor U16163 (N_16163,N_12680,N_11521);
xor U16164 (N_16164,N_11106,N_13945);
nor U16165 (N_16165,N_12961,N_12637);
and U16166 (N_16166,N_14918,N_14402);
nor U16167 (N_16167,N_11912,N_13433);
and U16168 (N_16168,N_11858,N_10630);
or U16169 (N_16169,N_10709,N_12923);
and U16170 (N_16170,N_10551,N_12770);
xor U16171 (N_16171,N_13412,N_11829);
nor U16172 (N_16172,N_12376,N_14834);
or U16173 (N_16173,N_12856,N_12782);
nor U16174 (N_16174,N_12215,N_11735);
and U16175 (N_16175,N_11866,N_13176);
nor U16176 (N_16176,N_14888,N_12719);
xnor U16177 (N_16177,N_10394,N_10267);
and U16178 (N_16178,N_13020,N_11609);
nand U16179 (N_16179,N_13324,N_11516);
and U16180 (N_16180,N_10493,N_10032);
and U16181 (N_16181,N_12745,N_13932);
and U16182 (N_16182,N_14163,N_12806);
and U16183 (N_16183,N_10338,N_14986);
or U16184 (N_16184,N_11354,N_11271);
and U16185 (N_16185,N_13990,N_10982);
nand U16186 (N_16186,N_12118,N_11000);
nand U16187 (N_16187,N_12086,N_11861);
nor U16188 (N_16188,N_14768,N_14514);
nand U16189 (N_16189,N_11067,N_13871);
xor U16190 (N_16190,N_10343,N_13219);
or U16191 (N_16191,N_12772,N_13317);
nand U16192 (N_16192,N_12074,N_10135);
or U16193 (N_16193,N_10644,N_12184);
and U16194 (N_16194,N_10188,N_10168);
xor U16195 (N_16195,N_13460,N_10101);
nor U16196 (N_16196,N_12899,N_13875);
nor U16197 (N_16197,N_10027,N_12525);
nor U16198 (N_16198,N_12143,N_12253);
nor U16199 (N_16199,N_10719,N_13842);
or U16200 (N_16200,N_11190,N_10714);
and U16201 (N_16201,N_11794,N_10517);
or U16202 (N_16202,N_13578,N_11425);
or U16203 (N_16203,N_11113,N_14485);
or U16204 (N_16204,N_11045,N_12010);
or U16205 (N_16205,N_10355,N_12904);
or U16206 (N_16206,N_10128,N_12072);
nand U16207 (N_16207,N_13573,N_12927);
nand U16208 (N_16208,N_14259,N_11359);
xor U16209 (N_16209,N_11653,N_13786);
or U16210 (N_16210,N_11996,N_13601);
and U16211 (N_16211,N_11696,N_13739);
nor U16212 (N_16212,N_10163,N_14865);
and U16213 (N_16213,N_10905,N_11135);
and U16214 (N_16214,N_12528,N_12322);
xor U16215 (N_16215,N_13795,N_14336);
nand U16216 (N_16216,N_14080,N_13723);
or U16217 (N_16217,N_14426,N_11244);
nor U16218 (N_16218,N_13704,N_10963);
or U16219 (N_16219,N_14687,N_12414);
nor U16220 (N_16220,N_10127,N_10540);
nand U16221 (N_16221,N_11572,N_14604);
nand U16222 (N_16222,N_13773,N_14325);
nand U16223 (N_16223,N_11322,N_13904);
or U16224 (N_16224,N_12452,N_14688);
or U16225 (N_16225,N_10114,N_14249);
and U16226 (N_16226,N_10068,N_14565);
nor U16227 (N_16227,N_14357,N_10685);
nand U16228 (N_16228,N_13961,N_14286);
nand U16229 (N_16229,N_13645,N_11961);
nor U16230 (N_16230,N_14931,N_14785);
nand U16231 (N_16231,N_12347,N_12186);
xnor U16232 (N_16232,N_14152,N_14031);
nor U16233 (N_16233,N_14806,N_13186);
xnor U16234 (N_16234,N_11739,N_13478);
xor U16235 (N_16235,N_11900,N_11101);
and U16236 (N_16236,N_10519,N_10717);
nor U16237 (N_16237,N_10415,N_13307);
or U16238 (N_16238,N_14281,N_10678);
xnor U16239 (N_16239,N_10826,N_13908);
nor U16240 (N_16240,N_13063,N_13703);
xor U16241 (N_16241,N_12175,N_12855);
nand U16242 (N_16242,N_14523,N_12793);
or U16243 (N_16243,N_11503,N_11772);
or U16244 (N_16244,N_14553,N_13438);
xnor U16245 (N_16245,N_12867,N_14656);
xor U16246 (N_16246,N_10725,N_10743);
nor U16247 (N_16247,N_13864,N_12583);
or U16248 (N_16248,N_10845,N_11413);
or U16249 (N_16249,N_12380,N_13295);
or U16250 (N_16250,N_11898,N_14702);
nor U16251 (N_16251,N_10549,N_13756);
or U16252 (N_16252,N_12344,N_10071);
nor U16253 (N_16253,N_11716,N_14272);
nor U16254 (N_16254,N_14026,N_12427);
and U16255 (N_16255,N_10022,N_12761);
nor U16256 (N_16256,N_11408,N_10628);
or U16257 (N_16257,N_11830,N_13080);
and U16258 (N_16258,N_10066,N_12540);
xnor U16259 (N_16259,N_13391,N_13270);
nand U16260 (N_16260,N_13983,N_14130);
nand U16261 (N_16261,N_13519,N_14398);
or U16262 (N_16262,N_10504,N_13321);
or U16263 (N_16263,N_14003,N_10287);
nand U16264 (N_16264,N_12083,N_12792);
nand U16265 (N_16265,N_14440,N_10913);
or U16266 (N_16266,N_11214,N_12949);
or U16267 (N_16267,N_10944,N_10276);
nand U16268 (N_16268,N_12390,N_12829);
nand U16269 (N_16269,N_14007,N_14454);
nor U16270 (N_16270,N_14115,N_13447);
and U16271 (N_16271,N_12704,N_10418);
nor U16272 (N_16272,N_13508,N_14154);
nor U16273 (N_16273,N_14573,N_13247);
xnor U16274 (N_16274,N_10155,N_12257);
nand U16275 (N_16275,N_14449,N_14761);
xor U16276 (N_16276,N_12209,N_10771);
or U16277 (N_16277,N_14850,N_10133);
nor U16278 (N_16278,N_13126,N_10866);
and U16279 (N_16279,N_10580,N_12367);
nor U16280 (N_16280,N_14355,N_14183);
nor U16281 (N_16281,N_11999,N_14167);
and U16282 (N_16282,N_10129,N_12892);
nor U16283 (N_16283,N_11533,N_13880);
nor U16284 (N_16284,N_12321,N_12289);
or U16285 (N_16285,N_13212,N_14557);
and U16286 (N_16286,N_12124,N_11527);
nor U16287 (N_16287,N_11444,N_11197);
nand U16288 (N_16288,N_11559,N_13060);
nor U16289 (N_16289,N_14639,N_11070);
xnor U16290 (N_16290,N_13228,N_11515);
nand U16291 (N_16291,N_13099,N_10997);
or U16292 (N_16292,N_13893,N_14913);
nand U16293 (N_16293,N_11799,N_12296);
or U16294 (N_16294,N_13965,N_13092);
nand U16295 (N_16295,N_12024,N_10382);
xor U16296 (N_16296,N_11227,N_14764);
or U16297 (N_16297,N_10821,N_12009);
xor U16298 (N_16298,N_13657,N_14472);
and U16299 (N_16299,N_14373,N_12936);
or U16300 (N_16300,N_13593,N_13919);
xor U16301 (N_16301,N_11449,N_13589);
or U16302 (N_16302,N_12425,N_11481);
nor U16303 (N_16303,N_14992,N_12088);
xor U16304 (N_16304,N_12613,N_13197);
or U16305 (N_16305,N_11906,N_11844);
and U16306 (N_16306,N_11099,N_12242);
nand U16307 (N_16307,N_14176,N_11231);
xnor U16308 (N_16308,N_11985,N_11466);
xor U16309 (N_16309,N_10596,N_11913);
nand U16310 (N_16310,N_13515,N_12748);
nand U16311 (N_16311,N_13065,N_13883);
nand U16312 (N_16312,N_13627,N_11296);
nor U16313 (N_16313,N_11392,N_13759);
nand U16314 (N_16314,N_11547,N_10046);
nand U16315 (N_16315,N_13585,N_13461);
and U16316 (N_16316,N_11060,N_11792);
and U16317 (N_16317,N_11781,N_14227);
and U16318 (N_16318,N_12517,N_10660);
nor U16319 (N_16319,N_11960,N_13975);
or U16320 (N_16320,N_10602,N_14235);
nor U16321 (N_16321,N_11968,N_11317);
or U16322 (N_16322,N_10254,N_13264);
nor U16323 (N_16323,N_14526,N_10667);
xor U16324 (N_16324,N_11426,N_11655);
nor U16325 (N_16325,N_11788,N_12026);
and U16326 (N_16326,N_10586,N_11802);
xor U16327 (N_16327,N_12587,N_13259);
nor U16328 (N_16328,N_13205,N_14296);
nand U16329 (N_16329,N_11209,N_13135);
and U16330 (N_16330,N_12928,N_14663);
nand U16331 (N_16331,N_11640,N_13653);
nand U16332 (N_16332,N_13991,N_12957);
or U16333 (N_16333,N_12744,N_12339);
xor U16334 (N_16334,N_10748,N_14593);
nor U16335 (N_16335,N_12073,N_11686);
or U16336 (N_16336,N_14778,N_13646);
nor U16337 (N_16337,N_10829,N_12195);
nand U16338 (N_16338,N_14005,N_11356);
nand U16339 (N_16339,N_14049,N_11556);
nand U16340 (N_16340,N_13293,N_11180);
nor U16341 (N_16341,N_12001,N_14509);
nor U16342 (N_16342,N_10927,N_12930);
or U16343 (N_16343,N_13992,N_13715);
nor U16344 (N_16344,N_12559,N_12037);
or U16345 (N_16345,N_13512,N_13397);
xnor U16346 (N_16346,N_14789,N_13680);
xnor U16347 (N_16347,N_11301,N_13421);
nand U16348 (N_16348,N_12467,N_12189);
or U16349 (N_16349,N_10074,N_13708);
xnor U16350 (N_16350,N_14981,N_11022);
and U16351 (N_16351,N_12747,N_11501);
or U16352 (N_16352,N_14024,N_10769);
nor U16353 (N_16353,N_14177,N_14759);
nor U16354 (N_16354,N_11577,N_12801);
nand U16355 (N_16355,N_10535,N_11717);
xor U16356 (N_16356,N_10575,N_12155);
and U16357 (N_16357,N_11925,N_12301);
or U16358 (N_16358,N_14921,N_14051);
nor U16359 (N_16359,N_11391,N_10964);
or U16360 (N_16360,N_12597,N_13813);
xor U16361 (N_16361,N_11564,N_10045);
xor U16362 (N_16362,N_14032,N_14712);
xnor U16363 (N_16363,N_13695,N_11281);
xor U16364 (N_16364,N_11279,N_12958);
xor U16365 (N_16365,N_14399,N_11039);
xor U16366 (N_16366,N_12310,N_14795);
and U16367 (N_16367,N_13343,N_11258);
xor U16368 (N_16368,N_10582,N_11831);
nor U16369 (N_16369,N_10898,N_13190);
and U16370 (N_16370,N_12370,N_11936);
xor U16371 (N_16371,N_13863,N_12251);
or U16372 (N_16372,N_13157,N_13297);
xnor U16373 (N_16373,N_11905,N_14819);
xnor U16374 (N_16374,N_13435,N_14201);
or U16375 (N_16375,N_12695,N_14859);
nor U16376 (N_16376,N_10138,N_14623);
nand U16377 (N_16377,N_12580,N_12976);
and U16378 (N_16378,N_11808,N_14337);
and U16379 (N_16379,N_12243,N_11642);
and U16380 (N_16380,N_11637,N_13700);
or U16381 (N_16381,N_14208,N_12832);
nand U16382 (N_16382,N_12594,N_12685);
or U16383 (N_16383,N_14670,N_11683);
or U16384 (N_16384,N_11079,N_14821);
xnor U16385 (N_16385,N_11857,N_10860);
and U16386 (N_16386,N_11329,N_11378);
and U16387 (N_16387,N_11289,N_12599);
nand U16388 (N_16388,N_14307,N_12688);
nand U16389 (N_16389,N_11043,N_13554);
nor U16390 (N_16390,N_13656,N_13531);
nor U16391 (N_16391,N_11612,N_14256);
and U16392 (N_16392,N_11955,N_13668);
nor U16393 (N_16393,N_11495,N_13290);
and U16394 (N_16394,N_11591,N_11546);
and U16395 (N_16395,N_12883,N_12960);
or U16396 (N_16396,N_13819,N_12055);
xor U16397 (N_16397,N_10189,N_11797);
or U16398 (N_16398,N_10942,N_11676);
nand U16399 (N_16399,N_13408,N_10627);
and U16400 (N_16400,N_10285,N_12896);
and U16401 (N_16401,N_14995,N_10601);
and U16402 (N_16402,N_14645,N_14073);
and U16403 (N_16403,N_14280,N_12313);
nor U16404 (N_16404,N_13010,N_13481);
or U16405 (N_16405,N_10470,N_11474);
nor U16406 (N_16406,N_13049,N_12208);
or U16407 (N_16407,N_13749,N_12673);
nand U16408 (N_16408,N_13691,N_14742);
or U16409 (N_16409,N_11346,N_10204);
nor U16410 (N_16410,N_14450,N_11881);
xnor U16411 (N_16411,N_12846,N_13330);
or U16412 (N_16412,N_12398,N_13693);
and U16413 (N_16413,N_10383,N_12095);
xnor U16414 (N_16414,N_11123,N_13637);
xnor U16415 (N_16415,N_10237,N_12281);
xor U16416 (N_16416,N_13037,N_14381);
nor U16417 (N_16417,N_14269,N_11252);
or U16418 (N_16418,N_10116,N_14360);
or U16419 (N_16419,N_13156,N_11165);
nand U16420 (N_16420,N_12905,N_13766);
xor U16421 (N_16421,N_14738,N_13926);
nand U16422 (N_16422,N_13982,N_10500);
and U16423 (N_16423,N_10980,N_14203);
or U16424 (N_16424,N_10617,N_11517);
or U16425 (N_16425,N_14653,N_12555);
and U16426 (N_16426,N_10499,N_14081);
or U16427 (N_16427,N_13218,N_10258);
nor U16428 (N_16428,N_10570,N_11737);
nor U16429 (N_16429,N_12888,N_12015);
and U16430 (N_16430,N_10361,N_10081);
xnor U16431 (N_16431,N_12043,N_13688);
and U16432 (N_16432,N_12457,N_11627);
nor U16433 (N_16433,N_11657,N_11338);
nor U16434 (N_16434,N_13038,N_12456);
nor U16435 (N_16435,N_14749,N_14437);
xnor U16436 (N_16436,N_13827,N_14960);
nand U16437 (N_16437,N_10924,N_11367);
nand U16438 (N_16438,N_11316,N_13078);
nor U16439 (N_16439,N_10772,N_13050);
nor U16440 (N_16440,N_12749,N_13551);
and U16441 (N_16441,N_10738,N_10815);
xnor U16442 (N_16442,N_12032,N_11950);
xnor U16443 (N_16443,N_11078,N_11525);
nand U16444 (N_16444,N_14468,N_13810);
xor U16445 (N_16445,N_14221,N_11973);
or U16446 (N_16446,N_13807,N_12275);
xor U16447 (N_16447,N_13014,N_13265);
or U16448 (N_16448,N_14899,N_12262);
or U16449 (N_16449,N_14289,N_14482);
xnor U16450 (N_16450,N_10395,N_10206);
nor U16451 (N_16451,N_13710,N_11993);
nor U16452 (N_16452,N_11579,N_13889);
or U16453 (N_16453,N_10797,N_14739);
or U16454 (N_16454,N_14725,N_10344);
nand U16455 (N_16455,N_10335,N_14676);
xnor U16456 (N_16456,N_13719,N_12626);
and U16457 (N_16457,N_14292,N_10841);
or U16458 (N_16458,N_12602,N_10222);
nor U16459 (N_16459,N_12033,N_12374);
or U16460 (N_16460,N_12338,N_13869);
nor U16461 (N_16461,N_10830,N_11903);
xor U16462 (N_16462,N_14019,N_12893);
nor U16463 (N_16463,N_13484,N_14597);
or U16464 (N_16464,N_13387,N_10314);
xnor U16465 (N_16465,N_10888,N_14217);
or U16466 (N_16466,N_13340,N_14796);
and U16467 (N_16467,N_12527,N_13313);
nand U16468 (N_16468,N_14142,N_11832);
xor U16469 (N_16469,N_14370,N_14730);
and U16470 (N_16470,N_12505,N_10911);
and U16471 (N_16471,N_14056,N_10989);
or U16472 (N_16472,N_10260,N_14922);
or U16473 (N_16473,N_10048,N_12386);
nor U16474 (N_16474,N_14706,N_13271);
nand U16475 (N_16475,N_14146,N_11406);
or U16476 (N_16476,N_13927,N_13411);
nor U16477 (N_16477,N_14570,N_12766);
nand U16478 (N_16478,N_13614,N_13676);
xnor U16479 (N_16479,N_12134,N_11049);
or U16480 (N_16480,N_11478,N_12509);
xnor U16481 (N_16481,N_12810,N_13649);
nand U16482 (N_16482,N_14997,N_14460);
nand U16483 (N_16483,N_12285,N_10104);
or U16484 (N_16484,N_11511,N_11884);
nand U16485 (N_16485,N_10893,N_14909);
and U16486 (N_16486,N_13782,N_14428);
and U16487 (N_16487,N_13214,N_14484);
xnor U16488 (N_16488,N_14354,N_12304);
nor U16489 (N_16489,N_13959,N_13824);
xor U16490 (N_16490,N_14694,N_13320);
or U16491 (N_16491,N_12212,N_11211);
or U16492 (N_16492,N_12204,N_12557);
or U16493 (N_16493,N_13079,N_11150);
xnor U16494 (N_16494,N_14071,N_13518);
and U16495 (N_16495,N_12471,N_14824);
xor U16496 (N_16496,N_11255,N_14901);
nor U16497 (N_16497,N_10701,N_12664);
nor U16498 (N_16498,N_14774,N_13808);
nand U16499 (N_16499,N_14641,N_13230);
nor U16500 (N_16500,N_13083,N_13588);
nor U16501 (N_16501,N_12397,N_14762);
or U16502 (N_16502,N_12491,N_10726);
or U16503 (N_16503,N_13924,N_10172);
nand U16504 (N_16504,N_13507,N_11313);
xnor U16505 (N_16505,N_10820,N_10119);
nand U16506 (N_16506,N_14411,N_10391);
nand U16507 (N_16507,N_14367,N_11615);
xor U16508 (N_16508,N_12824,N_13495);
nor U16509 (N_16509,N_10783,N_13158);
or U16510 (N_16510,N_13948,N_10251);
and U16511 (N_16511,N_13189,N_14324);
nand U16512 (N_16512,N_13848,N_10791);
and U16513 (N_16513,N_10566,N_14723);
nor U16514 (N_16514,N_13173,N_13576);
nand U16515 (N_16515,N_14635,N_14430);
nor U16516 (N_16516,N_10923,N_11946);
and U16517 (N_16517,N_13950,N_12468);
and U16518 (N_16518,N_11170,N_12811);
xnor U16519 (N_16519,N_11763,N_12488);
nand U16520 (N_16520,N_10435,N_13440);
nand U16521 (N_16521,N_11670,N_12729);
nand U16522 (N_16522,N_11801,N_10089);
nor U16523 (N_16523,N_14636,N_14205);
or U16524 (N_16524,N_10863,N_10673);
nand U16525 (N_16525,N_11604,N_14162);
and U16526 (N_16526,N_12548,N_14632);
and U16527 (N_16527,N_14376,N_10827);
or U16528 (N_16528,N_13046,N_13548);
or U16529 (N_16529,N_11541,N_11293);
and U16530 (N_16530,N_11341,N_10904);
xnor U16531 (N_16531,N_11298,N_10193);
nand U16532 (N_16532,N_14168,N_12807);
nor U16533 (N_16533,N_10624,N_11740);
or U16534 (N_16534,N_14075,N_12765);
nor U16535 (N_16535,N_10640,N_14420);
nor U16536 (N_16536,N_10632,N_12040);
nand U16537 (N_16537,N_14823,N_14594);
nor U16538 (N_16538,N_11878,N_13255);
xor U16539 (N_16539,N_14322,N_13369);
and U16540 (N_16540,N_12872,N_12595);
or U16541 (N_16541,N_13758,N_13735);
and U16542 (N_16542,N_12650,N_14736);
nor U16543 (N_16543,N_14499,N_10423);
xor U16544 (N_16544,N_14512,N_10626);
and U16545 (N_16545,N_12866,N_13226);
xor U16546 (N_16546,N_10315,N_10788);
or U16547 (N_16547,N_12614,N_10161);
nand U16548 (N_16548,N_12937,N_12753);
nor U16549 (N_16549,N_14123,N_12646);
or U16550 (N_16550,N_11459,N_10522);
and U16551 (N_16551,N_14303,N_11188);
nand U16552 (N_16552,N_11358,N_13323);
nor U16553 (N_16553,N_14116,N_12241);
nand U16554 (N_16554,N_11452,N_12137);
xor U16555 (N_16555,N_12214,N_12496);
xnor U16556 (N_16556,N_11259,N_14556);
nand U16557 (N_16557,N_14849,N_11268);
nor U16558 (N_16558,N_14710,N_13110);
nand U16559 (N_16559,N_14858,N_13269);
nand U16560 (N_16560,N_12326,N_10775);
and U16561 (N_16561,N_11891,N_13471);
and U16562 (N_16562,N_12771,N_13752);
xor U16563 (N_16563,N_10696,N_11918);
nand U16564 (N_16564,N_12768,N_10024);
and U16565 (N_16565,N_12739,N_10487);
nor U16566 (N_16566,N_13292,N_10721);
nor U16567 (N_16567,N_12372,N_10613);
and U16568 (N_16568,N_12708,N_13879);
xor U16569 (N_16569,N_12934,N_12600);
and U16570 (N_16570,N_14158,N_11854);
nor U16571 (N_16571,N_13422,N_11631);
xnor U16572 (N_16572,N_12789,N_13532);
and U16573 (N_16573,N_11161,N_12921);
nand U16574 (N_16574,N_13454,N_13283);
nand U16575 (N_16575,N_11859,N_10705);
xnor U16576 (N_16576,N_10608,N_14944);
nand U16577 (N_16577,N_10356,N_13354);
or U16578 (N_16578,N_13192,N_11349);
nand U16579 (N_16579,N_14920,N_11235);
xnor U16580 (N_16580,N_13015,N_13272);
or U16581 (N_16581,N_14275,N_12110);
nand U16582 (N_16582,N_12365,N_14476);
and U16583 (N_16583,N_11183,N_11311);
nand U16584 (N_16584,N_13019,N_14416);
and U16585 (N_16585,N_11815,N_13768);
xor U16586 (N_16586,N_10545,N_14961);
nor U16587 (N_16587,N_10934,N_14181);
nand U16588 (N_16588,N_13339,N_14359);
or U16589 (N_16589,N_12198,N_12067);
xor U16590 (N_16590,N_10422,N_11723);
nand U16591 (N_16591,N_12948,N_10035);
nand U16592 (N_16592,N_12082,N_12423);
and U16593 (N_16593,N_11352,N_10946);
and U16594 (N_16594,N_14220,N_12568);
nor U16595 (N_16595,N_14976,N_12090);
or U16596 (N_16596,N_14946,N_11742);
nand U16597 (N_16597,N_13326,N_11519);
and U16598 (N_16598,N_14422,N_14298);
or U16599 (N_16599,N_11492,N_10186);
nor U16600 (N_16600,N_14008,N_11688);
and U16601 (N_16601,N_11782,N_13553);
nand U16602 (N_16602,N_13744,N_11593);
xor U16603 (N_16603,N_13928,N_11890);
and U16604 (N_16604,N_11685,N_10533);
or U16605 (N_16605,N_10351,N_10468);
or U16606 (N_16606,N_13223,N_10831);
and U16607 (N_16607,N_14836,N_14109);
nor U16608 (N_16608,N_14127,N_13534);
or U16609 (N_16609,N_14917,N_14202);
xnor U16610 (N_16610,N_11916,N_11991);
nor U16611 (N_16611,N_11133,N_12478);
nor U16612 (N_16612,N_10637,N_13360);
nand U16613 (N_16613,N_13960,N_14218);
xnor U16614 (N_16614,N_10631,N_10263);
or U16615 (N_16615,N_12790,N_11158);
xor U16616 (N_16616,N_14683,N_10247);
xor U16617 (N_16617,N_11575,N_11755);
nor U16618 (N_16618,N_10807,N_11031);
xnor U16619 (N_16619,N_12260,N_14862);
or U16620 (N_16620,N_10146,N_12543);
nand U16621 (N_16621,N_12332,N_14470);
nor U16622 (N_16622,N_13733,N_10871);
nor U16623 (N_16623,N_10615,N_10093);
nor U16624 (N_16624,N_11328,N_10079);
nand U16625 (N_16625,N_14786,N_14258);
nand U16626 (N_16626,N_12179,N_14238);
and U16627 (N_16627,N_14756,N_12999);
xor U16628 (N_16628,N_13712,N_10152);
xor U16629 (N_16629,N_12049,N_12908);
or U16630 (N_16630,N_14825,N_11692);
xor U16631 (N_16631,N_13121,N_10762);
or U16632 (N_16632,N_12327,N_13413);
nor U16633 (N_16633,N_14787,N_11280);
and U16634 (N_16634,N_11184,N_13641);
xnor U16635 (N_16635,N_14766,N_12363);
nand U16636 (N_16636,N_11959,N_14971);
or U16637 (N_16637,N_13571,N_12938);
nand U16638 (N_16638,N_13045,N_11065);
or U16639 (N_16639,N_10492,N_10067);
and U16640 (N_16640,N_12975,N_13859);
nand U16641 (N_16641,N_11721,N_12282);
nor U16642 (N_16642,N_13592,N_13246);
nor U16643 (N_16643,N_13654,N_10292);
nand U16644 (N_16644,N_11718,N_11365);
xnor U16645 (N_16645,N_14681,N_12475);
and U16646 (N_16646,N_11272,N_12962);
xor U16647 (N_16647,N_11254,N_11561);
xor U16648 (N_16648,N_11006,N_12314);
xor U16649 (N_16649,N_14191,N_14085);
or U16650 (N_16650,N_11075,N_13168);
or U16651 (N_16651,N_13944,N_14731);
nand U16652 (N_16652,N_12180,N_11497);
nor U16653 (N_16653,N_14132,N_14693);
nor U16654 (N_16654,N_12248,N_11379);
or U16655 (N_16655,N_12023,N_13120);
nand U16656 (N_16656,N_13084,N_10588);
and U16657 (N_16657,N_10597,N_12007);
and U16658 (N_16658,N_12985,N_14128);
nor U16659 (N_16659,N_13380,N_12362);
nand U16660 (N_16660,N_10744,N_12495);
and U16661 (N_16661,N_10528,N_11809);
xnor U16662 (N_16662,N_11335,N_11966);
or U16663 (N_16663,N_13424,N_12145);
nor U16664 (N_16664,N_11080,N_10176);
and U16665 (N_16665,N_13674,N_10229);
xor U16666 (N_16666,N_10228,N_12986);
and U16667 (N_16667,N_13432,N_14495);
nor U16668 (N_16668,N_10846,N_10842);
and U16669 (N_16669,N_14964,N_10990);
nor U16670 (N_16670,N_12566,N_11015);
nor U16671 (N_16671,N_11964,N_13465);
xor U16672 (N_16672,N_14590,N_11371);
or U16673 (N_16673,N_12812,N_13458);
nand U16674 (N_16674,N_10080,N_10296);
nor U16675 (N_16675,N_12940,N_14560);
nor U16676 (N_16676,N_11340,N_14164);
and U16677 (N_16677,N_10578,N_14448);
and U16678 (N_16678,N_10198,N_11628);
nand U16679 (N_16679,N_13242,N_13235);
nor U16680 (N_16680,N_10909,N_10053);
and U16681 (N_16681,N_10281,N_13967);
nand U16682 (N_16682,N_10209,N_13055);
nand U16683 (N_16683,N_10190,N_11442);
and U16684 (N_16684,N_14938,N_13675);
xnor U16685 (N_16685,N_14684,N_10106);
or U16686 (N_16686,N_10452,N_14200);
xnor U16687 (N_16687,N_10230,N_10564);
nor U16688 (N_16688,N_10525,N_13801);
nand U16689 (N_16689,N_11573,N_13849);
xnor U16690 (N_16690,N_10195,N_11450);
or U16691 (N_16691,N_12499,N_14783);
nor U16692 (N_16692,N_14672,N_14857);
or U16693 (N_16693,N_13895,N_13115);
nor U16694 (N_16694,N_11768,N_10708);
nand U16695 (N_16695,N_12348,N_12450);
or U16696 (N_16696,N_11761,N_14020);
and U16697 (N_16697,N_14861,N_13785);
or U16698 (N_16698,N_14361,N_14247);
nor U16699 (N_16699,N_13104,N_10008);
and U16700 (N_16700,N_10050,N_13866);
xor U16701 (N_16701,N_10227,N_13414);
nand U16702 (N_16702,N_14134,N_13428);
xor U16703 (N_16703,N_12229,N_13878);
xor U16704 (N_16704,N_13409,N_14282);
and U16705 (N_16705,N_12203,N_10377);
nor U16706 (N_16706,N_10297,N_14947);
nor U16707 (N_16707,N_10047,N_12290);
and U16708 (N_16708,N_14083,N_11646);
nand U16709 (N_16709,N_11166,N_10196);
nand U16710 (N_16710,N_14034,N_11614);
xor U16711 (N_16711,N_12000,N_13022);
and U16712 (N_16712,N_11638,N_13364);
and U16713 (N_16713,N_12512,N_10710);
or U16714 (N_16714,N_12359,N_14104);
or U16715 (N_16715,N_13138,N_13560);
or U16716 (N_16716,N_12897,N_11584);
nand U16717 (N_16717,N_13328,N_10773);
and U16718 (N_16718,N_11935,N_13535);
and U16719 (N_16719,N_12103,N_12643);
nand U16720 (N_16720,N_13031,N_11856);
nand U16721 (N_16721,N_10595,N_10224);
or U16722 (N_16722,N_13517,N_12291);
or U16723 (N_16723,N_11410,N_13729);
xor U16724 (N_16724,N_13798,N_12461);
and U16725 (N_16725,N_10523,N_11085);
and U16726 (N_16726,N_10899,N_12693);
and U16727 (N_16727,N_14879,N_11312);
nor U16728 (N_16728,N_12933,N_13669);
nand U16729 (N_16729,N_11030,N_11019);
and U16730 (N_16730,N_10451,N_10402);
and U16731 (N_16731,N_10745,N_14972);
or U16732 (N_16732,N_13779,N_11332);
nand U16733 (N_16733,N_13089,N_13482);
and U16734 (N_16734,N_10642,N_10007);
and U16735 (N_16735,N_11684,N_11483);
nand U16736 (N_16736,N_14244,N_12335);
and U16737 (N_16737,N_14103,N_14536);
and U16738 (N_16738,N_10715,N_14924);
and U16739 (N_16739,N_13453,N_11750);
or U16740 (N_16740,N_13163,N_10367);
xnor U16741 (N_16741,N_14988,N_14949);
nor U16742 (N_16742,N_12682,N_10834);
nand U16743 (N_16743,N_13929,N_10030);
nor U16744 (N_16744,N_11373,N_10354);
or U16745 (N_16745,N_12192,N_12107);
and U16746 (N_16746,N_11538,N_11853);
nor U16747 (N_16747,N_10139,N_11284);
nand U16748 (N_16748,N_11708,N_12571);
xnor U16749 (N_16749,N_12994,N_10872);
or U16750 (N_16750,N_11156,N_11454);
nand U16751 (N_16751,N_10177,N_11592);
xor U16752 (N_16752,N_14506,N_12439);
and U16753 (N_16753,N_12929,N_11793);
or U16754 (N_16754,N_11665,N_10554);
or U16755 (N_16755,N_12286,N_13763);
nand U16756 (N_16756,N_13086,N_11416);
and U16757 (N_16757,N_12932,N_11888);
xnor U16758 (N_16758,N_10854,N_14979);
or U16759 (N_16759,N_12545,N_10607);
and U16760 (N_16760,N_12361,N_13748);
nand U16761 (N_16761,N_12620,N_10043);
and U16762 (N_16762,N_13096,N_14053);
nand U16763 (N_16763,N_14406,N_14211);
nand U16764 (N_16764,N_12689,N_11153);
nor U16765 (N_16765,N_11697,N_12676);
nor U16766 (N_16766,N_11144,N_11446);
xor U16767 (N_16767,N_14210,N_11141);
nand U16768 (N_16768,N_14409,N_11947);
xor U16769 (N_16769,N_12652,N_12787);
or U16770 (N_16770,N_13683,N_13625);
nand U16771 (N_16771,N_12443,N_12014);
xnor U16772 (N_16772,N_13770,N_12647);
or U16773 (N_16773,N_10301,N_13244);
xnor U16774 (N_16774,N_11958,N_14229);
or U16775 (N_16775,N_13717,N_14404);
or U16776 (N_16776,N_13792,N_12714);
nand U16777 (N_16777,N_13231,N_11992);
nor U16778 (N_16778,N_11499,N_12052);
and U16779 (N_16779,N_10682,N_11468);
and U16780 (N_16780,N_10269,N_10814);
xnor U16781 (N_16781,N_12395,N_12802);
or U16782 (N_16782,N_12120,N_10765);
xnor U16783 (N_16783,N_12308,N_11839);
nor U16784 (N_16784,N_14883,N_10157);
nor U16785 (N_16785,N_14501,N_10689);
and U16786 (N_16786,N_14107,N_11142);
nor U16787 (N_16787,N_12591,N_14301);
and U16788 (N_16788,N_12151,N_10727);
nor U16789 (N_16789,N_14442,N_12006);
nand U16790 (N_16790,N_11120,N_10805);
nand U16791 (N_16791,N_13070,N_12298);
nand U16792 (N_16792,N_11669,N_12601);
and U16793 (N_16793,N_12247,N_10234);
xnor U16794 (N_16794,N_10712,N_11405);
and U16795 (N_16795,N_12660,N_14149);
nor U16796 (N_16796,N_14576,N_13117);
and U16797 (N_16797,N_13407,N_13028);
or U16798 (N_16798,N_13523,N_11662);
nor U16799 (N_16799,N_14400,N_13497);
xor U16800 (N_16800,N_13052,N_11484);
nor U16801 (N_16801,N_12109,N_10565);
xnor U16802 (N_16802,N_11752,N_14780);
nor U16803 (N_16803,N_11862,N_11364);
and U16804 (N_16804,N_10445,N_10900);
nand U16805 (N_16805,N_14048,N_14283);
xnor U16806 (N_16806,N_14648,N_13954);
xnor U16807 (N_16807,N_12455,N_13306);
nand U16808 (N_16808,N_13805,N_13406);
nand U16809 (N_16809,N_13582,N_14809);
nand U16810 (N_16810,N_11625,N_11643);
or U16811 (N_16811,N_13200,N_11756);
or U16812 (N_16812,N_12042,N_10136);
xnor U16813 (N_16813,N_12329,N_13692);
nand U16814 (N_16814,N_11616,N_14469);
nand U16815 (N_16815,N_13917,N_14160);
or U16816 (N_16816,N_11623,N_11849);
nand U16817 (N_16817,N_12384,N_13822);
or U16818 (N_16818,N_10438,N_13897);
or U16819 (N_16819,N_10910,N_14805);
or U16820 (N_16820,N_13913,N_14262);
xnor U16821 (N_16821,N_12925,N_12567);
or U16822 (N_16822,N_14265,N_11644);
nand U16823 (N_16823,N_12995,N_13074);
xnor U16824 (N_16824,N_12617,N_13113);
or U16825 (N_16825,N_13761,N_14732);
and U16826 (N_16826,N_10472,N_13689);
nor U16827 (N_16827,N_10557,N_12894);
or U16828 (N_16828,N_11957,N_10223);
nor U16829 (N_16829,N_11337,N_14459);
or U16830 (N_16830,N_10232,N_12114);
and U16831 (N_16831,N_11567,N_13177);
and U16832 (N_16832,N_12541,N_14793);
and U16833 (N_16833,N_10061,N_11368);
xor U16834 (N_16834,N_14839,N_12100);
nor U16835 (N_16835,N_12474,N_13860);
and U16836 (N_16836,N_14798,N_10085);
or U16837 (N_16837,N_11361,N_11044);
and U16838 (N_16838,N_12584,N_12355);
xor U16839 (N_16839,N_13638,N_11326);
xor U16840 (N_16840,N_11222,N_10264);
nor U16841 (N_16841,N_13167,N_14418);
and U16842 (N_16842,N_12227,N_13830);
nor U16843 (N_16843,N_13485,N_11013);
xnor U16844 (N_16844,N_14934,N_10951);
and U16845 (N_16845,N_10308,N_13626);
nand U16846 (N_16846,N_11324,N_10786);
nand U16847 (N_16847,N_14089,N_11504);
and U16848 (N_16848,N_10884,N_10852);
nand U16849 (N_16849,N_10657,N_10420);
xnor U16850 (N_16850,N_14434,N_12631);
and U16851 (N_16851,N_11382,N_13024);
xor U16852 (N_16852,N_10283,N_14232);
nand U16853 (N_16853,N_14911,N_14345);
nand U16854 (N_16854,N_12481,N_10877);
nor U16855 (N_16855,N_10103,N_13603);
nor U16856 (N_16856,N_14568,N_11671);
or U16857 (N_16857,N_10881,N_10350);
nand U16858 (N_16858,N_10164,N_10385);
nor U16859 (N_16859,N_12596,N_14956);
or U16860 (N_16860,N_10574,N_13017);
and U16861 (N_16861,N_11585,N_14747);
and U16862 (N_16862,N_13803,N_11300);
nor U16863 (N_16863,N_11155,N_13716);
and U16864 (N_16864,N_12108,N_10339);
nand U16865 (N_16865,N_11647,N_11487);
or U16866 (N_16866,N_13840,N_14488);
nand U16867 (N_16867,N_12004,N_11736);
and U16868 (N_16868,N_10017,N_13935);
nand U16869 (N_16869,N_11084,N_14352);
or U16870 (N_16870,N_12069,N_11034);
xor U16871 (N_16871,N_12132,N_13697);
xnor U16872 (N_16872,N_11860,N_13618);
nand U16873 (N_16873,N_13620,N_10439);
nor U16874 (N_16874,N_10399,N_12551);
nand U16875 (N_16875,N_10334,N_12183);
or U16876 (N_16876,N_13062,N_11191);
nor U16877 (N_16877,N_13619,N_13936);
or U16878 (N_16878,N_14502,N_11636);
nand U16879 (N_16879,N_12853,N_14378);
xnor U16880 (N_16880,N_13375,N_13464);
nand U16881 (N_16881,N_12219,N_13701);
nor U16882 (N_16882,N_12648,N_13994);
and U16883 (N_16883,N_10491,N_14647);
nand U16884 (N_16884,N_12027,N_10681);
nand U16885 (N_16885,N_13949,N_10483);
nor U16886 (N_16886,N_12422,N_13806);
nor U16887 (N_16887,N_13882,N_13220);
nor U16888 (N_16888,N_11639,N_14561);
or U16889 (N_16889,N_12264,N_12057);
nor U16890 (N_16890,N_11009,N_11370);
xnor U16891 (N_16891,N_13152,N_10042);
or U16892 (N_16892,N_10459,N_14456);
xor U16893 (N_16893,N_12449,N_14679);
nand U16894 (N_16894,N_10225,N_12213);
xor U16895 (N_16895,N_10832,N_14186);
or U16896 (N_16896,N_13314,N_14863);
nand U16897 (N_16897,N_10156,N_13258);
and U16898 (N_16898,N_11956,N_12199);
and U16899 (N_16899,N_14919,N_14317);
and U16900 (N_16900,N_14894,N_11821);
or U16901 (N_16901,N_13544,N_10559);
or U16902 (N_16902,N_13005,N_12433);
nor U16903 (N_16903,N_10291,N_13533);
xnor U16904 (N_16904,N_12075,N_14875);
xnor U16905 (N_16905,N_11435,N_11457);
nand U16906 (N_16906,N_10861,N_13981);
and U16907 (N_16907,N_13466,N_13367);
and U16908 (N_16908,N_14754,N_12230);
and U16909 (N_16909,N_10981,N_14385);
nor U16910 (N_16910,N_12553,N_14447);
nor U16911 (N_16911,N_14028,N_13056);
xnor U16912 (N_16912,N_13498,N_11520);
nor U16913 (N_16913,N_13403,N_13916);
nand U16914 (N_16914,N_10534,N_10711);
nor U16915 (N_16915,N_10337,N_11846);
nor U16916 (N_16916,N_12667,N_14974);
nor U16917 (N_16917,N_11402,N_13661);
xor U16918 (N_16918,N_14895,N_10560);
xnor U16919 (N_16919,N_13562,N_10219);
nand U16920 (N_16920,N_11963,N_11530);
xor U16921 (N_16921,N_13359,N_10953);
xor U16922 (N_16922,N_14036,N_10690);
nand U16923 (N_16923,N_11983,N_14040);
nor U16924 (N_16924,N_13389,N_14760);
nor U16925 (N_16925,N_12408,N_13912);
xor U16926 (N_16926,N_11001,N_13448);
xnor U16927 (N_16927,N_10389,N_11025);
xnor U16928 (N_16928,N_12945,N_13285);
and U16929 (N_16929,N_14666,N_14595);
xnor U16930 (N_16930,N_14904,N_12044);
nor U16931 (N_16931,N_11353,N_10838);
nand U16932 (N_16932,N_11810,N_10986);
xnor U16933 (N_16933,N_11667,N_13356);
or U16934 (N_16934,N_11267,N_10259);
nor U16935 (N_16935,N_14551,N_13109);
xor U16936 (N_16936,N_12323,N_14781);
nor U16937 (N_16937,N_11597,N_10265);
and U16938 (N_16938,N_11902,N_12046);
nand U16939 (N_16939,N_11246,N_10277);
nand U16940 (N_16940,N_13357,N_14196);
or U16941 (N_16941,N_12154,N_13764);
and U16942 (N_16942,N_14294,N_11327);
nand U16943 (N_16943,N_13890,N_11851);
nor U16944 (N_16944,N_13388,N_12418);
and U16945 (N_16945,N_12713,N_14343);
xnor U16946 (N_16946,N_12814,N_12588);
nor U16947 (N_16947,N_13707,N_13208);
nor U16948 (N_16948,N_12858,N_10729);
nor U16949 (N_16949,N_14023,N_13263);
and U16950 (N_16950,N_12890,N_10426);
xor U16951 (N_16951,N_12767,N_14994);
nor U16952 (N_16952,N_14574,N_10970);
and U16953 (N_16953,N_11827,N_10849);
nor U16954 (N_16954,N_13861,N_10675);
or U16955 (N_16955,N_12302,N_12358);
xnor U16956 (N_16956,N_12311,N_10180);
nand U16957 (N_16957,N_12552,N_13133);
xnor U16958 (N_16958,N_11529,N_13404);
and U16959 (N_16959,N_13709,N_12101);
nor U16960 (N_16960,N_14637,N_12104);
xor U16961 (N_16961,N_11064,N_10378);
or U16962 (N_16962,N_14496,N_11892);
xnor U16963 (N_16963,N_14185,N_12483);
or U16964 (N_16964,N_11095,N_12272);
xor U16965 (N_16965,N_14622,N_10620);
and U16966 (N_16966,N_14212,N_13394);
nor U16967 (N_16967,N_11086,N_12051);
nand U16968 (N_16968,N_10056,N_13439);
and U16969 (N_16969,N_14854,N_14620);
and U16970 (N_16970,N_12250,N_11331);
nor U16971 (N_16971,N_14375,N_13706);
or U16972 (N_16972,N_10967,N_14610);
and U16973 (N_16973,N_13652,N_10185);
nor U16974 (N_16974,N_10941,N_13332);
nor U16975 (N_16975,N_10962,N_13791);
or U16976 (N_16976,N_12964,N_12903);
or U16977 (N_16977,N_12558,N_10411);
nand U16978 (N_16978,N_13686,N_14273);
and U16979 (N_16979,N_12860,N_10943);
xor U16980 (N_16980,N_14989,N_12563);
or U16981 (N_16981,N_13787,N_10612);
xor U16982 (N_16982,N_11200,N_12514);
nor U16983 (N_16983,N_12277,N_13581);
nand U16984 (N_16984,N_10142,N_12835);
or U16985 (N_16985,N_12393,N_11024);
or U16986 (N_16986,N_11943,N_11033);
xor U16987 (N_16987,N_14717,N_12911);
xor U16988 (N_16988,N_13922,N_12678);
xnor U16989 (N_16989,N_13599,N_10779);
and U16990 (N_16990,N_13137,N_10097);
and U16991 (N_16991,N_11552,N_12669);
nor U16992 (N_16992,N_10121,N_11911);
and U16993 (N_16993,N_12341,N_12629);
xor U16994 (N_16994,N_12318,N_14330);
or U16995 (N_16995,N_11069,N_14329);
xor U16996 (N_16996,N_14952,N_12665);
and U16997 (N_16997,N_10948,N_14174);
nand U16998 (N_16998,N_11306,N_14148);
xnor U16999 (N_16999,N_14930,N_13333);
nor U17000 (N_17000,N_13047,N_14569);
and U17001 (N_17001,N_10896,N_10294);
nor U17002 (N_17002,N_12501,N_13781);
xnor U17003 (N_17003,N_13797,N_11978);
nor U17004 (N_17004,N_14813,N_14384);
nor U17005 (N_17005,N_10648,N_14733);
nand U17006 (N_17006,N_12039,N_13261);
nor U17007 (N_17007,N_14601,N_11982);
or U17008 (N_17008,N_12902,N_10381);
nor U17009 (N_17009,N_12546,N_13346);
or U17010 (N_17010,N_13233,N_12831);
nand U17011 (N_17011,N_10396,N_10633);
or U17012 (N_17012,N_11800,N_10723);
or U17013 (N_17013,N_11012,N_10793);
or U17014 (N_17014,N_10716,N_13767);
and U17015 (N_17015,N_12306,N_14344);
xnor U17016 (N_17016,N_12352,N_13812);
or U17017 (N_17017,N_11412,N_11551);
xor U17018 (N_17018,N_12079,N_11273);
xnor U17019 (N_17019,N_14515,N_11545);
xnor U17020 (N_17020,N_10918,N_13361);
and U17021 (N_17021,N_13892,N_14661);
xor U17022 (N_17022,N_14763,N_10494);
and U17023 (N_17023,N_11400,N_13632);
nor U17024 (N_17024,N_10440,N_12668);
and U17025 (N_17025,N_12356,N_12997);
or U17026 (N_17026,N_11482,N_11309);
or U17027 (N_17027,N_13004,N_11565);
nor U17028 (N_17028,N_12979,N_14455);
nor U17029 (N_17029,N_12025,N_14101);
xnor U17030 (N_17030,N_10238,N_10720);
and U17031 (N_17031,N_12881,N_11248);
nor U17032 (N_17032,N_11213,N_11219);
xnor U17033 (N_17033,N_11897,N_11621);
or U17034 (N_17034,N_11199,N_12854);
nor U17035 (N_17035,N_11938,N_11693);
or U17036 (N_17036,N_14630,N_12724);
nor U17037 (N_17037,N_12337,N_11008);
xnor U17038 (N_17038,N_13114,N_10357);
nor U17039 (N_17039,N_10289,N_13885);
or U17040 (N_17040,N_13489,N_13736);
nand U17041 (N_17041,N_11828,N_14504);
nor U17042 (N_17042,N_10865,N_12534);
xnor U17043 (N_17043,N_11432,N_11965);
and U17044 (N_17044,N_13934,N_13996);
xnor U17045 (N_17045,N_12181,N_12953);
nor U17046 (N_17046,N_11894,N_12679);
or U17047 (N_17047,N_12582,N_12093);
and U17048 (N_17048,N_14458,N_12671);
and U17049 (N_17049,N_12585,N_10653);
and U17050 (N_17050,N_14473,N_14699);
nand U17051 (N_17051,N_13227,N_11376);
nand U17052 (N_17052,N_14039,N_13462);
and U17053 (N_17053,N_12880,N_10886);
and U17054 (N_17054,N_13841,N_14716);
or U17055 (N_17055,N_13682,N_11176);
nand U17056 (N_17056,N_14004,N_11194);
xnor U17057 (N_17057,N_11343,N_11148);
or U17058 (N_17058,N_13617,N_11357);
nor U17059 (N_17059,N_13687,N_13832);
xnor U17060 (N_17060,N_13881,N_11775);
xnor U17061 (N_17061,N_11666,N_10656);
or U17062 (N_17062,N_13018,N_12845);
or U17063 (N_17063,N_13090,N_10248);
and U17064 (N_17064,N_14230,N_14872);
xnor U17065 (N_17065,N_14643,N_10665);
nand U17066 (N_17066,N_14943,N_12518);
nand U17067 (N_17067,N_14436,N_12788);
or U17068 (N_17068,N_14197,N_14063);
nor U17069 (N_17069,N_11949,N_12056);
nand U17070 (N_17070,N_10912,N_11532);
or U17071 (N_17071,N_14252,N_11549);
nor U17072 (N_17072,N_12522,N_10920);
xor U17073 (N_17073,N_12684,N_11163);
nand U17074 (N_17074,N_11877,N_11104);
and U17075 (N_17075,N_10840,N_14757);
nand U17076 (N_17076,N_11873,N_13702);
nand U17077 (N_17077,N_13854,N_14592);
and U17078 (N_17078,N_14157,N_14603);
nand U17079 (N_17079,N_14001,N_13953);
nand U17080 (N_17080,N_10130,N_12019);
nor U17081 (N_17081,N_12066,N_14178);
and U17082 (N_17082,N_10576,N_12294);
or U17083 (N_17083,N_10808,N_12497);
nor U17084 (N_17084,N_14022,N_14654);
and U17085 (N_17085,N_12211,N_13579);
and U17086 (N_17086,N_11869,N_14517);
xnor U17087 (N_17087,N_12624,N_13906);
nor U17088 (N_17088,N_10972,N_12592);
nand U17089 (N_17089,N_10220,N_14954);
and U17090 (N_17090,N_12463,N_13903);
and U17091 (N_17091,N_10240,N_12785);
nand U17092 (N_17092,N_12396,N_11243);
xnor U17093 (N_17093,N_10526,N_10062);
and U17094 (N_17094,N_13966,N_14151);
or U17095 (N_17095,N_12589,N_10330);
and U17096 (N_17096,N_14380,N_14815);
or U17097 (N_17097,N_10009,N_12156);
or U17098 (N_17098,N_12144,N_10303);
xor U17099 (N_17099,N_11928,N_11146);
nor U17100 (N_17100,N_12606,N_11498);
or U17101 (N_17101,N_11914,N_13276);
nor U17102 (N_17102,N_13250,N_11951);
nor U17103 (N_17103,N_10754,N_12350);
or U17104 (N_17104,N_10410,N_11011);
or U17105 (N_17105,N_13067,N_14326);
and U17106 (N_17106,N_13279,N_12991);
xnor U17107 (N_17107,N_12502,N_14714);
nor U17108 (N_17108,N_13753,N_13850);
or U17109 (N_17109,N_13977,N_14415);
xnor U17110 (N_17110,N_12573,N_12070);
nor U17111 (N_17111,N_13855,N_14860);
and U17112 (N_17112,N_10284,N_10252);
or U17113 (N_17113,N_11967,N_10796);
and U17114 (N_17114,N_12873,N_11463);
and U17115 (N_17115,N_10514,N_12437);
and U17116 (N_17116,N_10245,N_11464);
xnor U17117 (N_17117,N_10816,N_14471);
and U17118 (N_17118,N_13061,N_13663);
nand U17119 (N_17119,N_11926,N_11282);
and U17120 (N_17120,N_12718,N_13837);
nor U17121 (N_17121,N_14646,N_11020);
nand U17122 (N_17122,N_12825,N_11840);
xor U17123 (N_17123,N_12843,N_14138);
nor U17124 (N_17124,N_11321,N_13823);
or U17125 (N_17125,N_14837,N_14701);
xor U17126 (N_17126,N_11588,N_11901);
or U17127 (N_17127,N_14870,N_12136);
nor U17128 (N_17128,N_10210,N_12692);
nor U17129 (N_17129,N_11434,N_12263);
or U17130 (N_17130,N_13470,N_14175);
xor U17131 (N_17131,N_10496,N_13112);
and U17132 (N_17132,N_13318,N_12008);
or U17133 (N_17133,N_11526,N_10647);
nand U17134 (N_17134,N_11240,N_11766);
nand U17135 (N_17135,N_13355,N_14582);
nor U17136 (N_17136,N_12954,N_12800);
nor U17137 (N_17137,N_13872,N_10065);
xnor U17138 (N_17138,N_13274,N_13445);
nand U17139 (N_17139,N_12956,N_11699);
nor U17140 (N_17140,N_12187,N_14079);
and U17141 (N_17141,N_14465,N_14968);
xnor U17142 (N_17142,N_10041,N_11848);
or U17143 (N_17143,N_12462,N_11407);
nand U17144 (N_17144,N_13506,N_10661);
or U17145 (N_17145,N_13087,N_14219);
nand U17146 (N_17146,N_12720,N_13241);
xnor U17147 (N_17147,N_13597,N_13094);
and U17148 (N_17148,N_11355,N_13281);
and U17149 (N_17149,N_12966,N_12424);
or U17150 (N_17150,N_14658,N_14320);
xnor U17151 (N_17151,N_12168,N_10600);
and U17152 (N_17152,N_10300,N_12565);
or U17153 (N_17153,N_11675,N_11427);
nand U17154 (N_17154,N_10747,N_11622);
nor U17155 (N_17155,N_14816,N_13238);
nor U17156 (N_17156,N_11687,N_14967);
and U17157 (N_17157,N_14143,N_14866);
or U17158 (N_17158,N_13474,N_10364);
or U17159 (N_17159,N_10874,N_10664);
xnor U17160 (N_17160,N_12529,N_14356);
nand U17161 (N_17161,N_10408,N_10672);
and U17162 (N_17162,N_12674,N_13858);
and U17163 (N_17163,N_14091,N_12126);
xor U17164 (N_17164,N_12827,N_13750);
nor U17165 (N_17165,N_12416,N_14119);
or U17166 (N_17166,N_14314,N_11456);
nand U17167 (N_17167,N_14155,N_14873);
and U17168 (N_17168,N_12089,N_13058);
and U17169 (N_17169,N_13372,N_13331);
nor U17170 (N_17170,N_11980,N_10122);
xor U17171 (N_17171,N_12677,N_10246);
or U17172 (N_17172,N_10324,N_10401);
and U17173 (N_17173,N_10782,N_14002);
nand U17174 (N_17174,N_14206,N_14744);
and U17175 (N_17175,N_12011,N_13505);
nor U17176 (N_17176,N_12420,N_11710);
and U17177 (N_17177,N_10498,N_12959);
nor U17178 (N_17178,N_13310,N_12196);
and U17179 (N_17179,N_11098,N_10510);
nor U17180 (N_17180,N_10039,N_14746);
nand U17181 (N_17181,N_10216,N_10261);
nand U17182 (N_17182,N_14369,N_10542);
or U17183 (N_17183,N_11074,N_14800);
nor U17184 (N_17184,N_10437,N_13178);
nor U17185 (N_17185,N_11007,N_12085);
or U17186 (N_17186,N_11185,N_13266);
nor U17187 (N_17187,N_10985,N_13613);
nand U17188 (N_17188,N_11661,N_14737);
xor U17189 (N_17189,N_14444,N_10327);
nor U17190 (N_17190,N_10867,N_11072);
nor U17191 (N_17191,N_14309,N_10538);
nor U17192 (N_17192,N_11472,N_14707);
xor U17193 (N_17193,N_13521,N_10795);
or U17194 (N_17194,N_14776,N_10587);
or U17195 (N_17195,N_11108,N_10713);
xor U17196 (N_17196,N_12426,N_11465);
nor U17197 (N_17197,N_10304,N_10643);
nand U17198 (N_17198,N_14928,N_12621);
or U17199 (N_17199,N_14745,N_10393);
nor U17200 (N_17200,N_11785,N_11668);
or U17201 (N_17201,N_10569,N_10409);
xor U17202 (N_17202,N_12176,N_14098);
nand U17203 (N_17203,N_12404,N_11507);
or U17204 (N_17204,N_13524,N_13325);
xnor U17205 (N_17205,N_13921,N_12482);
xor U17206 (N_17206,N_12833,N_10604);
xnor U17207 (N_17207,N_12003,N_10293);
xor U17208 (N_17208,N_11887,N_14288);
or U17209 (N_17209,N_12185,N_10134);
nor U17210 (N_17210,N_14055,N_13136);
nor U17211 (N_17211,N_13608,N_12430);
nor U17212 (N_17212,N_13260,N_14248);
and U17213 (N_17213,N_10629,N_12417);
xor U17214 (N_17214,N_10362,N_11369);
or U17215 (N_17215,N_13501,N_14572);
or U17216 (N_17216,N_14638,N_11270);
or U17217 (N_17217,N_13600,N_12642);
nor U17218 (N_17218,N_11057,N_14050);
xor U17219 (N_17219,N_13093,N_10623);
or U17220 (N_17220,N_14984,N_11048);
and U17221 (N_17221,N_10070,N_14983);
xnor U17222 (N_17222,N_12874,N_11157);
xor U17223 (N_17223,N_10969,N_12754);
or U17224 (N_17224,N_10509,N_13876);
and U17225 (N_17225,N_14784,N_13621);
xnor U17226 (N_17226,N_13980,N_14948);
and U17227 (N_17227,N_14521,N_13514);
nand U17228 (N_17228,N_13938,N_14432);
nor U17229 (N_17229,N_14600,N_11239);
and U17230 (N_17230,N_12317,N_13443);
and U17231 (N_17231,N_11469,N_12530);
nand U17232 (N_17232,N_13130,N_12480);
nor U17233 (N_17233,N_12446,N_13845);
and U17234 (N_17234,N_12805,N_11390);
and U17235 (N_17235,N_11303,N_13699);
nor U17236 (N_17236,N_11266,N_10885);
nor U17237 (N_17237,N_14140,N_10174);
or U17238 (N_17238,N_14435,N_14064);
and U17239 (N_17239,N_14383,N_12521);
or U17240 (N_17240,N_14927,N_11107);
nor U17241 (N_17241,N_12616,N_10434);
or U17242 (N_17242,N_11375,N_10798);
xnor U17243 (N_17243,N_11236,N_12727);
and U17244 (N_17244,N_12870,N_11319);
and U17245 (N_17245,N_11143,N_12353);
or U17246 (N_17246,N_13896,N_14150);
nor U17247 (N_17247,N_12699,N_13494);
and U17248 (N_17248,N_11603,N_13449);
or U17249 (N_17249,N_11728,N_14086);
nor U17250 (N_17250,N_14374,N_14599);
xor U17251 (N_17251,N_13559,N_10515);
and U17252 (N_17252,N_10698,N_11706);
or U17253 (N_17253,N_13694,N_13937);
or U17254 (N_17254,N_13161,N_11981);
nand U17255 (N_17255,N_10759,N_11937);
and U17256 (N_17256,N_10998,N_12851);
nand U17257 (N_17257,N_14724,N_12798);
nor U17258 (N_17258,N_11220,N_10555);
nand U17259 (N_17259,N_14790,N_10026);
xor U17260 (N_17260,N_12500,N_13106);
nand U17261 (N_17261,N_12343,N_14363);
nand U17262 (N_17262,N_13224,N_10571);
nand U17263 (N_17263,N_13636,N_13221);
or U17264 (N_17264,N_11385,N_14133);
nor U17265 (N_17265,N_11931,N_10443);
or U17266 (N_17266,N_14826,N_14403);
or U17267 (N_17267,N_14425,N_11746);
or U17268 (N_17268,N_13287,N_11724);
or U17269 (N_17269,N_11738,N_14010);
and U17270 (N_17270,N_10482,N_10603);
or U17271 (N_17271,N_12519,N_14489);
nand U17272 (N_17272,N_13475,N_14096);
or U17273 (N_17273,N_13565,N_11733);
nor U17274 (N_17274,N_14621,N_12436);
xor U17275 (N_17275,N_13829,N_10153);
xor U17276 (N_17276,N_12886,N_12510);
nor U17277 (N_17277,N_14740,N_11518);
or U17278 (N_17278,N_10480,N_14933);
xnor U17279 (N_17279,N_12316,N_12965);
or U17280 (N_17280,N_11845,N_10764);
xor U17281 (N_17281,N_11129,N_13337);
and U17282 (N_17282,N_14391,N_13574);
nor U17283 (N_17283,N_10054,N_10424);
xnor U17284 (N_17284,N_11673,N_10870);
xnor U17285 (N_17285,N_10322,N_10659);
nor U17286 (N_17286,N_14131,N_13216);
nand U17287 (N_17287,N_12884,N_11262);
or U17288 (N_17288,N_12169,N_12654);
nor U17289 (N_17289,N_11479,N_11276);
or U17290 (N_17290,N_14340,N_13987);
and U17291 (N_17291,N_10908,N_11954);
nand U17292 (N_17292,N_12194,N_10298);
and U17293 (N_17293,N_14347,N_14692);
nor U17294 (N_17294,N_10403,N_10348);
and U17295 (N_17295,N_10674,N_11904);
or U17296 (N_17296,N_10506,N_10201);
nor U17297 (N_17297,N_11930,N_13315);
xor U17298 (N_17298,N_10781,N_10370);
and U17299 (N_17299,N_13536,N_12029);
nor U17300 (N_17300,N_11447,N_12077);
xor U17301 (N_17301,N_14141,N_12852);
nor U17302 (N_17302,N_12231,N_10577);
xor U17303 (N_17303,N_14618,N_11885);
or U17304 (N_17304,N_11396,N_12258);
nand U17305 (N_17305,N_11052,N_14065);
and U17306 (N_17306,N_14803,N_14541);
and U17307 (N_17307,N_10262,N_10345);
nor U17308 (N_17308,N_10416,N_11921);
nand U17309 (N_17309,N_12939,N_12804);
xnor U17310 (N_17310,N_14327,N_10752);
xnor U17311 (N_17311,N_13549,N_11387);
or U17312 (N_17312,N_14649,N_10144);
xor U17313 (N_17313,N_10763,N_10183);
xnor U17314 (N_17314,N_12632,N_12225);
or U17315 (N_17315,N_14735,N_11553);
nand U17316 (N_17316,N_12237,N_10919);
xnor U17317 (N_17317,N_10730,N_14990);
nand U17318 (N_17318,N_14102,N_12623);
or U17319 (N_17319,N_13147,N_11342);
nand U17320 (N_17320,N_11605,N_14528);
xnor U17321 (N_17321,N_11927,N_11023);
nor U17322 (N_17322,N_13529,N_14111);
nand U17323 (N_17323,N_14832,N_12445);
nor U17324 (N_17324,N_11299,N_14755);
xnor U17325 (N_17325,N_11719,N_10115);
nor U17326 (N_17326,N_14874,N_10518);
and U17327 (N_17327,N_10869,N_10442);
xor U17328 (N_17328,N_10619,N_10460);
xor U17329 (N_17329,N_13257,N_12131);
nor U17330 (N_17330,N_14673,N_10319);
or U17331 (N_17331,N_14452,N_10691);
or U17332 (N_17332,N_13504,N_10171);
or U17333 (N_17333,N_13846,N_11145);
and U17334 (N_17334,N_11131,N_10226);
nor U17335 (N_17335,N_12871,N_13267);
and U17336 (N_17336,N_11632,N_10211);
nor U17337 (N_17337,N_14166,N_10221);
or U17338 (N_17338,N_13725,N_14341);
and U17339 (N_17339,N_13351,N_13188);
nor U17340 (N_17340,N_10159,N_11021);
or U17341 (N_17341,N_10581,N_14209);
nor U17342 (N_17342,N_12053,N_12223);
nor U17343 (N_17343,N_10449,N_12235);
or U17344 (N_17344,N_10621,N_13939);
nand U17345 (N_17345,N_11066,N_10940);
or U17346 (N_17346,N_10803,N_12058);
nand U17347 (N_17347,N_11035,N_13352);
xor U17348 (N_17348,N_10686,N_14074);
nand U17349 (N_17349,N_14852,N_13229);
or U17350 (N_17350,N_11819,N_12045);
nand U17351 (N_17351,N_11970,N_10655);
nor U17352 (N_17352,N_14250,N_11017);
xnor U17353 (N_17353,N_14609,N_14831);
and U17354 (N_17354,N_11709,N_14122);
or U17355 (N_17355,N_14524,N_12944);
xnor U17356 (N_17356,N_13665,N_12130);
nand U17357 (N_17357,N_14966,N_13076);
or U17358 (N_17358,N_12857,N_10978);
xor U17359 (N_17359,N_10360,N_14531);
and U17360 (N_17360,N_12054,N_12357);
nor U17361 (N_17361,N_10380,N_14351);
and U17362 (N_17362,N_11320,N_11658);
xnor U17363 (N_17363,N_12330,N_10857);
nor U17364 (N_17364,N_11582,N_11796);
nand U17365 (N_17365,N_12740,N_12206);
nor U17366 (N_17366,N_14353,N_13053);
and U17367 (N_17367,N_11864,N_14467);
nand U17368 (N_17368,N_12486,N_11102);
and U17369 (N_17369,N_10069,N_12061);
or U17370 (N_17370,N_10938,N_14300);
nand U17371 (N_17371,N_11679,N_14996);
and U17372 (N_17372,N_12412,N_10639);
xor U17373 (N_17373,N_13108,N_11786);
nor U17374 (N_17374,N_12375,N_11619);
nand U17375 (N_17375,N_14290,N_10737);
or U17376 (N_17376,N_14855,N_11138);
or U17377 (N_17377,N_14907,N_13920);
and U17378 (N_17378,N_14255,N_11051);
or U17379 (N_17379,N_14187,N_13201);
nand U17380 (N_17380,N_10505,N_14959);
nand U17381 (N_17381,N_10836,N_12544);
xor U17382 (N_17382,N_10002,N_14664);
nand U17383 (N_17383,N_11534,N_11505);
nand U17384 (N_17384,N_10598,N_13059);
and U17385 (N_17385,N_13199,N_10270);
nand U17386 (N_17386,N_10092,N_10777);
xnor U17387 (N_17387,N_10562,N_10728);
or U17388 (N_17388,N_14429,N_12336);
xnor U17389 (N_17389,N_12271,N_12173);
xnor U17390 (N_17390,N_11164,N_10016);
or U17391 (N_17391,N_11088,N_11192);
and U17392 (N_17392,N_10774,N_11571);
nor U17393 (N_17393,N_13441,N_13001);
nor U17394 (N_17394,N_13583,N_12950);
nand U17395 (N_17395,N_13815,N_10404);
nand U17396 (N_17396,N_11384,N_14480);
xor U17397 (N_17397,N_14589,N_10349);
xor U17398 (N_17398,N_10244,N_11837);
xor U17399 (N_17399,N_12847,N_13732);
or U17400 (N_17400,N_13396,N_14192);
or U17401 (N_17401,N_13970,N_14571);
nand U17402 (N_17402,N_11372,N_11783);
nor U17403 (N_17403,N_10695,N_11489);
and U17404 (N_17404,N_14240,N_10687);
or U17405 (N_17405,N_13794,N_11672);
nand U17406 (N_17406,N_11448,N_13743);
or U17407 (N_17407,N_13100,N_12895);
and U17408 (N_17408,N_13705,N_10018);
and U17409 (N_17409,N_10930,N_10579);
and U17410 (N_17410,N_13150,N_12382);
and U17411 (N_17411,N_11105,N_11835);
and U17412 (N_17412,N_10471,N_12458);
and U17413 (N_17413,N_11871,N_12146);
and U17414 (N_17414,N_12140,N_10358);
and U17415 (N_17415,N_14029,N_13985);
nand U17416 (N_17416,N_13681,N_12096);
xor U17417 (N_17417,N_14542,N_11778);
nand U17418 (N_17418,N_12351,N_14884);
xor U17419 (N_17419,N_13239,N_13616);
or U17420 (N_17420,N_12619,N_10448);
nor U17421 (N_17421,N_11285,N_14365);
or U17422 (N_17422,N_11073,N_10484);
nor U17423 (N_17423,N_12909,N_14828);
nand U17424 (N_17424,N_12161,N_13575);
nand U17425 (N_17425,N_10274,N_12711);
and U17426 (N_17426,N_14794,N_13033);
or U17427 (N_17427,N_11438,N_14596);
or U17428 (N_17428,N_12823,N_10922);
and U17429 (N_17429,N_12102,N_10688);
nand U17430 (N_17430,N_10461,N_11624);
or U17431 (N_17431,N_13377,N_13963);
xnor U17432 (N_17432,N_11590,N_12034);
nor U17433 (N_17433,N_10883,N_14412);
or U17434 (N_17434,N_10740,N_11915);
xnor U17435 (N_17435,N_13437,N_14108);
or U17436 (N_17436,N_10625,N_11269);
or U17437 (N_17437,N_11995,N_10250);
nand U17438 (N_17438,N_11771,N_14097);
nand U17439 (N_17439,N_11732,N_12656);
and U17440 (N_17440,N_12980,N_11347);
and U17441 (N_17441,N_13098,N_11729);
nand U17442 (N_17442,N_14241,N_11245);
nand U17443 (N_17443,N_10859,N_14253);
nand U17444 (N_17444,N_13502,N_10741);
xor U17445 (N_17445,N_12157,N_14704);
nor U17446 (N_17446,N_12153,N_12373);
and U17447 (N_17447,N_13998,N_12875);
and U17448 (N_17448,N_10427,N_14389);
nor U17449 (N_17449,N_12364,N_11522);
xnor U17450 (N_17450,N_10149,N_12808);
or U17451 (N_17451,N_11178,N_14851);
and U17452 (N_17452,N_11314,N_10977);
nor U17453 (N_17453,N_14583,N_11493);
xor U17454 (N_17454,N_13586,N_13510);
nand U17455 (N_17455,N_10992,N_12366);
nand U17456 (N_17456,N_11841,N_12076);
or U17457 (N_17457,N_13902,N_14929);
and U17458 (N_17458,N_10957,N_13363);
nand U17459 (N_17459,N_11126,N_12701);
or U17460 (N_17460,N_13839,N_10956);
nand U17461 (N_17461,N_14410,N_10552);
nand U17462 (N_17462,N_10392,N_13300);
nor U17463 (N_17463,N_11451,N_10075);
and U17464 (N_17464,N_10646,N_14867);
and U17465 (N_17465,N_10040,N_13713);
and U17466 (N_17466,N_13754,N_14547);
or U17467 (N_17467,N_12048,N_13280);
xnor U17468 (N_17468,N_12324,N_13125);
xor U17469 (N_17469,N_12762,N_10890);
and U17470 (N_17470,N_10536,N_14234);
nor U17471 (N_17471,N_11071,N_12863);
nor U17472 (N_17472,N_13747,N_13302);
nand U17473 (N_17473,N_11610,N_14897);
nand U17474 (N_17474,N_10768,N_14277);
nor U17475 (N_17475,N_14718,N_10288);
xnor U17476 (N_17476,N_10099,N_11455);
nor U17477 (N_17477,N_14382,N_12969);
or U17478 (N_17478,N_14697,N_14518);
nand U17479 (N_17479,N_14293,N_10671);
or U17480 (N_17480,N_10766,N_10241);
nor U17481 (N_17481,N_11743,N_11278);
nor U17482 (N_17482,N_11210,N_11822);
or U17483 (N_17483,N_11804,N_12459);
xor U17484 (N_17484,N_12725,N_11467);
or U17485 (N_17485,N_13030,N_11139);
xnor U17486 (N_17486,N_11649,N_14466);
and U17487 (N_17487,N_11062,N_11680);
and U17488 (N_17488,N_10949,N_14753);
and U17489 (N_17489,N_11613,N_14153);
or U17490 (N_17490,N_13329,N_12639);
and U17491 (N_17491,N_11757,N_14876);
nand U17492 (N_17492,N_14236,N_10573);
nor U17493 (N_17493,N_14522,N_12878);
xor U17494 (N_17494,N_13591,N_12750);
nand U17495 (N_17495,N_11562,N_14045);
or U17496 (N_17496,N_10799,N_14364);
xnor U17497 (N_17497,N_14121,N_10880);
nor U17498 (N_17498,N_14358,N_12988);
or U17499 (N_17499,N_14179,N_10592);
xnor U17500 (N_17500,N_11967,N_11003);
xnor U17501 (N_17501,N_10246,N_14837);
and U17502 (N_17502,N_13337,N_10121);
nor U17503 (N_17503,N_13290,N_12654);
nand U17504 (N_17504,N_13170,N_11518);
xor U17505 (N_17505,N_10761,N_12226);
and U17506 (N_17506,N_14424,N_14453);
or U17507 (N_17507,N_12572,N_14868);
or U17508 (N_17508,N_13940,N_11416);
or U17509 (N_17509,N_14842,N_12564);
and U17510 (N_17510,N_14344,N_13793);
xor U17511 (N_17511,N_12767,N_12283);
nand U17512 (N_17512,N_11078,N_10520);
xor U17513 (N_17513,N_11755,N_14242);
xor U17514 (N_17514,N_10220,N_11179);
nor U17515 (N_17515,N_13519,N_12839);
xnor U17516 (N_17516,N_14284,N_10275);
nand U17517 (N_17517,N_12531,N_10872);
nand U17518 (N_17518,N_11864,N_11556);
or U17519 (N_17519,N_13062,N_10691);
or U17520 (N_17520,N_11157,N_10992);
xnor U17521 (N_17521,N_13552,N_13313);
xnor U17522 (N_17522,N_11509,N_14242);
nand U17523 (N_17523,N_12590,N_14779);
nor U17524 (N_17524,N_10231,N_10100);
and U17525 (N_17525,N_14833,N_13212);
nor U17526 (N_17526,N_14052,N_10092);
nor U17527 (N_17527,N_13844,N_14791);
nor U17528 (N_17528,N_14111,N_10060);
nor U17529 (N_17529,N_10908,N_12697);
nor U17530 (N_17530,N_10704,N_12671);
nand U17531 (N_17531,N_10995,N_14648);
xnor U17532 (N_17532,N_14929,N_14992);
xnor U17533 (N_17533,N_10834,N_10692);
nand U17534 (N_17534,N_10743,N_12894);
and U17535 (N_17535,N_10832,N_14526);
nand U17536 (N_17536,N_12293,N_11721);
and U17537 (N_17537,N_13004,N_14332);
xnor U17538 (N_17538,N_10013,N_13987);
xnor U17539 (N_17539,N_11419,N_11443);
nor U17540 (N_17540,N_13569,N_10900);
nor U17541 (N_17541,N_10818,N_11790);
or U17542 (N_17542,N_13525,N_13860);
or U17543 (N_17543,N_14655,N_11158);
nand U17544 (N_17544,N_14403,N_10734);
nor U17545 (N_17545,N_10398,N_10754);
nand U17546 (N_17546,N_11420,N_12643);
and U17547 (N_17547,N_14071,N_14232);
xor U17548 (N_17548,N_10880,N_13379);
nand U17549 (N_17549,N_10221,N_14876);
nor U17550 (N_17550,N_14340,N_10969);
xor U17551 (N_17551,N_14267,N_10840);
or U17552 (N_17552,N_13884,N_12665);
xnor U17553 (N_17553,N_13556,N_14217);
nand U17554 (N_17554,N_14465,N_14514);
xnor U17555 (N_17555,N_11987,N_12017);
xor U17556 (N_17556,N_13474,N_13787);
xnor U17557 (N_17557,N_10762,N_10246);
and U17558 (N_17558,N_12996,N_13898);
and U17559 (N_17559,N_11106,N_13808);
xnor U17560 (N_17560,N_10845,N_13666);
and U17561 (N_17561,N_12745,N_10031);
xor U17562 (N_17562,N_10178,N_13501);
nor U17563 (N_17563,N_12577,N_11657);
and U17564 (N_17564,N_10057,N_14836);
nor U17565 (N_17565,N_13175,N_13135);
nor U17566 (N_17566,N_11671,N_12624);
or U17567 (N_17567,N_13132,N_10111);
or U17568 (N_17568,N_14750,N_14244);
xnor U17569 (N_17569,N_14302,N_14761);
xnor U17570 (N_17570,N_10194,N_11146);
and U17571 (N_17571,N_11277,N_14417);
or U17572 (N_17572,N_13273,N_14795);
xor U17573 (N_17573,N_11315,N_13734);
or U17574 (N_17574,N_14775,N_11147);
or U17575 (N_17575,N_10449,N_11559);
nor U17576 (N_17576,N_12165,N_11900);
nand U17577 (N_17577,N_12297,N_14233);
xnor U17578 (N_17578,N_12276,N_12436);
and U17579 (N_17579,N_14466,N_10108);
nor U17580 (N_17580,N_10695,N_11769);
and U17581 (N_17581,N_14776,N_13385);
nand U17582 (N_17582,N_14055,N_13690);
and U17583 (N_17583,N_12603,N_11085);
nand U17584 (N_17584,N_14196,N_12309);
or U17585 (N_17585,N_11377,N_14118);
xnor U17586 (N_17586,N_14245,N_12475);
or U17587 (N_17587,N_10566,N_14810);
or U17588 (N_17588,N_10036,N_10678);
nor U17589 (N_17589,N_10494,N_14233);
and U17590 (N_17590,N_10834,N_11113);
and U17591 (N_17591,N_12035,N_11215);
and U17592 (N_17592,N_12530,N_13638);
xor U17593 (N_17593,N_13143,N_11500);
nor U17594 (N_17594,N_13907,N_11195);
and U17595 (N_17595,N_12080,N_13992);
and U17596 (N_17596,N_11975,N_14045);
nand U17597 (N_17597,N_10893,N_12457);
xor U17598 (N_17598,N_14949,N_13719);
xnor U17599 (N_17599,N_10071,N_11906);
and U17600 (N_17600,N_12453,N_11647);
and U17601 (N_17601,N_14395,N_14312);
xnor U17602 (N_17602,N_12955,N_14851);
or U17603 (N_17603,N_13193,N_13196);
or U17604 (N_17604,N_13977,N_10347);
nor U17605 (N_17605,N_13197,N_11850);
nor U17606 (N_17606,N_12208,N_13115);
nand U17607 (N_17607,N_12922,N_12764);
nor U17608 (N_17608,N_12450,N_10486);
nand U17609 (N_17609,N_12362,N_10252);
or U17610 (N_17610,N_13342,N_14892);
xor U17611 (N_17611,N_12582,N_10601);
nor U17612 (N_17612,N_14717,N_11707);
nor U17613 (N_17613,N_10334,N_10092);
nor U17614 (N_17614,N_13684,N_14892);
and U17615 (N_17615,N_12439,N_13490);
nand U17616 (N_17616,N_11364,N_10072);
xnor U17617 (N_17617,N_14522,N_13477);
nor U17618 (N_17618,N_14564,N_10931);
xnor U17619 (N_17619,N_14107,N_14937);
and U17620 (N_17620,N_12366,N_10505);
or U17621 (N_17621,N_13560,N_14744);
nand U17622 (N_17622,N_10120,N_14060);
xor U17623 (N_17623,N_12742,N_11746);
or U17624 (N_17624,N_13271,N_12676);
nand U17625 (N_17625,N_10748,N_11080);
and U17626 (N_17626,N_10645,N_13029);
nor U17627 (N_17627,N_10577,N_14477);
xnor U17628 (N_17628,N_13063,N_14468);
xor U17629 (N_17629,N_11496,N_14112);
and U17630 (N_17630,N_13281,N_13075);
nand U17631 (N_17631,N_11948,N_10617);
xor U17632 (N_17632,N_10208,N_12006);
and U17633 (N_17633,N_12782,N_11158);
nor U17634 (N_17634,N_13449,N_10144);
xor U17635 (N_17635,N_14729,N_13592);
or U17636 (N_17636,N_11659,N_11061);
or U17637 (N_17637,N_10154,N_12495);
xnor U17638 (N_17638,N_12631,N_11420);
nor U17639 (N_17639,N_12859,N_12885);
or U17640 (N_17640,N_13812,N_12711);
and U17641 (N_17641,N_13743,N_10020);
or U17642 (N_17642,N_10171,N_10302);
xnor U17643 (N_17643,N_14101,N_12233);
xor U17644 (N_17644,N_13020,N_11016);
nand U17645 (N_17645,N_13772,N_10929);
nor U17646 (N_17646,N_11966,N_10938);
nand U17647 (N_17647,N_14456,N_10545);
and U17648 (N_17648,N_14685,N_13788);
nand U17649 (N_17649,N_14960,N_11976);
and U17650 (N_17650,N_14570,N_13319);
nand U17651 (N_17651,N_12924,N_10909);
nor U17652 (N_17652,N_14522,N_10170);
nor U17653 (N_17653,N_12857,N_12027);
nor U17654 (N_17654,N_10967,N_13454);
nor U17655 (N_17655,N_11313,N_12296);
or U17656 (N_17656,N_14174,N_11044);
and U17657 (N_17657,N_10523,N_10725);
xor U17658 (N_17658,N_11688,N_12203);
and U17659 (N_17659,N_12433,N_11671);
nand U17660 (N_17660,N_12603,N_13504);
or U17661 (N_17661,N_13983,N_14378);
xnor U17662 (N_17662,N_14974,N_13156);
or U17663 (N_17663,N_12994,N_13121);
nand U17664 (N_17664,N_13051,N_13675);
nor U17665 (N_17665,N_14671,N_13669);
xor U17666 (N_17666,N_11387,N_11989);
nand U17667 (N_17667,N_13425,N_11388);
xnor U17668 (N_17668,N_12822,N_14328);
and U17669 (N_17669,N_14268,N_11690);
nor U17670 (N_17670,N_14879,N_13737);
nand U17671 (N_17671,N_12270,N_10301);
xnor U17672 (N_17672,N_11552,N_14379);
nand U17673 (N_17673,N_12639,N_11106);
or U17674 (N_17674,N_13092,N_12325);
xor U17675 (N_17675,N_11559,N_14012);
nor U17676 (N_17676,N_13584,N_13198);
nand U17677 (N_17677,N_10099,N_10248);
nor U17678 (N_17678,N_10043,N_13060);
nor U17679 (N_17679,N_10345,N_12846);
or U17680 (N_17680,N_14461,N_13786);
nand U17681 (N_17681,N_14234,N_11262);
xor U17682 (N_17682,N_12859,N_11316);
and U17683 (N_17683,N_12523,N_14853);
nor U17684 (N_17684,N_13097,N_13056);
nand U17685 (N_17685,N_13548,N_11058);
xnor U17686 (N_17686,N_13184,N_14693);
or U17687 (N_17687,N_13979,N_10330);
or U17688 (N_17688,N_10858,N_14423);
and U17689 (N_17689,N_12794,N_11711);
xnor U17690 (N_17690,N_10134,N_10880);
xor U17691 (N_17691,N_10089,N_12308);
nand U17692 (N_17692,N_10210,N_12499);
and U17693 (N_17693,N_11376,N_12649);
xor U17694 (N_17694,N_12703,N_10064);
or U17695 (N_17695,N_13512,N_14434);
and U17696 (N_17696,N_12714,N_12934);
xor U17697 (N_17697,N_12177,N_11968);
nand U17698 (N_17698,N_10365,N_12141);
xnor U17699 (N_17699,N_14896,N_14510);
nand U17700 (N_17700,N_14774,N_12592);
and U17701 (N_17701,N_13028,N_13092);
xor U17702 (N_17702,N_10451,N_13792);
nor U17703 (N_17703,N_10599,N_12248);
and U17704 (N_17704,N_10507,N_13754);
nand U17705 (N_17705,N_13896,N_14026);
nor U17706 (N_17706,N_10581,N_12860);
xor U17707 (N_17707,N_11469,N_10099);
xnor U17708 (N_17708,N_14171,N_10025);
nor U17709 (N_17709,N_13388,N_13353);
nand U17710 (N_17710,N_11393,N_12715);
xor U17711 (N_17711,N_14056,N_13666);
nor U17712 (N_17712,N_10207,N_10718);
nand U17713 (N_17713,N_14734,N_11838);
nor U17714 (N_17714,N_11267,N_14064);
nor U17715 (N_17715,N_12786,N_10350);
xnor U17716 (N_17716,N_11475,N_12035);
xor U17717 (N_17717,N_10875,N_13914);
or U17718 (N_17718,N_12286,N_14310);
xor U17719 (N_17719,N_11116,N_12553);
nor U17720 (N_17720,N_13637,N_10242);
and U17721 (N_17721,N_13653,N_12890);
and U17722 (N_17722,N_13474,N_14587);
xor U17723 (N_17723,N_11256,N_13684);
xnor U17724 (N_17724,N_13110,N_13753);
or U17725 (N_17725,N_14919,N_12542);
and U17726 (N_17726,N_13623,N_13686);
nand U17727 (N_17727,N_10748,N_10126);
nand U17728 (N_17728,N_12614,N_11364);
nand U17729 (N_17729,N_10582,N_14954);
xnor U17730 (N_17730,N_14332,N_11219);
xnor U17731 (N_17731,N_11778,N_10226);
xor U17732 (N_17732,N_13008,N_14829);
nand U17733 (N_17733,N_10169,N_10859);
or U17734 (N_17734,N_11327,N_11592);
or U17735 (N_17735,N_11204,N_13820);
and U17736 (N_17736,N_10749,N_10844);
or U17737 (N_17737,N_14130,N_14467);
or U17738 (N_17738,N_13725,N_13949);
nand U17739 (N_17739,N_11590,N_10462);
and U17740 (N_17740,N_10843,N_13509);
or U17741 (N_17741,N_10819,N_11392);
nand U17742 (N_17742,N_10813,N_14914);
nand U17743 (N_17743,N_13557,N_14770);
nor U17744 (N_17744,N_11169,N_14640);
and U17745 (N_17745,N_13383,N_11842);
nor U17746 (N_17746,N_10989,N_12974);
or U17747 (N_17747,N_13681,N_11589);
and U17748 (N_17748,N_13030,N_13711);
or U17749 (N_17749,N_12263,N_10488);
and U17750 (N_17750,N_10699,N_13502);
or U17751 (N_17751,N_13568,N_11949);
xor U17752 (N_17752,N_13094,N_14380);
or U17753 (N_17753,N_14667,N_14999);
and U17754 (N_17754,N_14010,N_10854);
nor U17755 (N_17755,N_13298,N_10050);
nand U17756 (N_17756,N_12846,N_13732);
nand U17757 (N_17757,N_13165,N_10887);
and U17758 (N_17758,N_12297,N_14062);
nor U17759 (N_17759,N_11743,N_12463);
nand U17760 (N_17760,N_10151,N_14960);
and U17761 (N_17761,N_13437,N_13155);
nand U17762 (N_17762,N_12294,N_10896);
xnor U17763 (N_17763,N_13949,N_12146);
xor U17764 (N_17764,N_12447,N_12446);
xor U17765 (N_17765,N_11515,N_11493);
or U17766 (N_17766,N_12134,N_13340);
xnor U17767 (N_17767,N_12649,N_14941);
nand U17768 (N_17768,N_10339,N_12372);
or U17769 (N_17769,N_12939,N_11248);
xnor U17770 (N_17770,N_10929,N_12193);
nand U17771 (N_17771,N_11535,N_11690);
xor U17772 (N_17772,N_14817,N_13776);
xor U17773 (N_17773,N_11107,N_10105);
or U17774 (N_17774,N_12288,N_12384);
or U17775 (N_17775,N_12190,N_12810);
xor U17776 (N_17776,N_14195,N_12572);
nor U17777 (N_17777,N_12406,N_13774);
xor U17778 (N_17778,N_14976,N_10936);
xnor U17779 (N_17779,N_11759,N_12028);
or U17780 (N_17780,N_14203,N_13041);
xnor U17781 (N_17781,N_11499,N_14545);
nand U17782 (N_17782,N_11786,N_14313);
nor U17783 (N_17783,N_10382,N_12372);
and U17784 (N_17784,N_11473,N_14807);
nor U17785 (N_17785,N_10354,N_14395);
or U17786 (N_17786,N_12981,N_13420);
xnor U17787 (N_17787,N_12148,N_12161);
or U17788 (N_17788,N_11549,N_14081);
nor U17789 (N_17789,N_12512,N_13239);
xnor U17790 (N_17790,N_13581,N_14954);
nor U17791 (N_17791,N_10946,N_10871);
nand U17792 (N_17792,N_14511,N_11948);
or U17793 (N_17793,N_14806,N_13851);
nor U17794 (N_17794,N_14752,N_10922);
or U17795 (N_17795,N_14268,N_10519);
xnor U17796 (N_17796,N_10207,N_12437);
nor U17797 (N_17797,N_13674,N_12030);
and U17798 (N_17798,N_12512,N_14016);
nand U17799 (N_17799,N_13619,N_10522);
nor U17800 (N_17800,N_10105,N_10708);
nand U17801 (N_17801,N_11500,N_14858);
nor U17802 (N_17802,N_14185,N_13091);
nand U17803 (N_17803,N_11826,N_13486);
xor U17804 (N_17804,N_13848,N_14392);
nor U17805 (N_17805,N_14112,N_10827);
and U17806 (N_17806,N_13835,N_11410);
and U17807 (N_17807,N_10491,N_10441);
xor U17808 (N_17808,N_12144,N_12786);
and U17809 (N_17809,N_12453,N_13160);
or U17810 (N_17810,N_14403,N_10724);
xnor U17811 (N_17811,N_14689,N_12474);
xnor U17812 (N_17812,N_10924,N_12993);
or U17813 (N_17813,N_14675,N_12059);
nor U17814 (N_17814,N_12846,N_10771);
and U17815 (N_17815,N_13060,N_14035);
nand U17816 (N_17816,N_12412,N_14469);
and U17817 (N_17817,N_10415,N_13578);
nand U17818 (N_17818,N_10485,N_11377);
or U17819 (N_17819,N_11231,N_12061);
and U17820 (N_17820,N_11906,N_14241);
nor U17821 (N_17821,N_12695,N_10837);
and U17822 (N_17822,N_10113,N_12716);
or U17823 (N_17823,N_11477,N_12458);
and U17824 (N_17824,N_12368,N_13287);
nand U17825 (N_17825,N_11018,N_12632);
xor U17826 (N_17826,N_13183,N_14949);
or U17827 (N_17827,N_12057,N_12203);
or U17828 (N_17828,N_13362,N_11691);
nor U17829 (N_17829,N_13944,N_11756);
xor U17830 (N_17830,N_10063,N_14924);
and U17831 (N_17831,N_12233,N_12255);
or U17832 (N_17832,N_14607,N_11087);
or U17833 (N_17833,N_10204,N_14197);
or U17834 (N_17834,N_13394,N_14330);
xor U17835 (N_17835,N_11384,N_13857);
nand U17836 (N_17836,N_10025,N_11861);
and U17837 (N_17837,N_11435,N_14265);
and U17838 (N_17838,N_11799,N_11632);
xor U17839 (N_17839,N_14197,N_13061);
nand U17840 (N_17840,N_11193,N_12318);
nand U17841 (N_17841,N_14535,N_14356);
xnor U17842 (N_17842,N_10791,N_11674);
nand U17843 (N_17843,N_10924,N_11873);
nor U17844 (N_17844,N_14875,N_10583);
or U17845 (N_17845,N_11029,N_14542);
or U17846 (N_17846,N_13173,N_10900);
nand U17847 (N_17847,N_12038,N_12893);
xnor U17848 (N_17848,N_11641,N_10659);
and U17849 (N_17849,N_12458,N_12721);
or U17850 (N_17850,N_10888,N_11014);
or U17851 (N_17851,N_13922,N_14275);
xnor U17852 (N_17852,N_14487,N_11466);
xnor U17853 (N_17853,N_10742,N_12943);
or U17854 (N_17854,N_10204,N_11673);
and U17855 (N_17855,N_12678,N_12426);
nand U17856 (N_17856,N_10847,N_12332);
or U17857 (N_17857,N_13696,N_12163);
xor U17858 (N_17858,N_11493,N_14848);
nor U17859 (N_17859,N_13417,N_11335);
nor U17860 (N_17860,N_14347,N_11087);
nor U17861 (N_17861,N_10298,N_14290);
nand U17862 (N_17862,N_11597,N_11575);
nor U17863 (N_17863,N_14109,N_11572);
and U17864 (N_17864,N_10542,N_11835);
or U17865 (N_17865,N_11677,N_11544);
xnor U17866 (N_17866,N_11349,N_14287);
xor U17867 (N_17867,N_13209,N_14641);
nand U17868 (N_17868,N_13360,N_12497);
or U17869 (N_17869,N_10259,N_10200);
nand U17870 (N_17870,N_14098,N_13354);
or U17871 (N_17871,N_13999,N_13215);
and U17872 (N_17872,N_10998,N_13785);
and U17873 (N_17873,N_14001,N_11843);
and U17874 (N_17874,N_11135,N_10689);
nor U17875 (N_17875,N_14211,N_11638);
nand U17876 (N_17876,N_10081,N_10412);
nand U17877 (N_17877,N_13375,N_10517);
or U17878 (N_17878,N_11691,N_13025);
nor U17879 (N_17879,N_13385,N_11038);
nor U17880 (N_17880,N_13047,N_12977);
and U17881 (N_17881,N_11591,N_14867);
nand U17882 (N_17882,N_14322,N_10691);
nand U17883 (N_17883,N_14531,N_14162);
or U17884 (N_17884,N_11659,N_10575);
or U17885 (N_17885,N_14842,N_10207);
xor U17886 (N_17886,N_14321,N_10762);
nand U17887 (N_17887,N_13658,N_11140);
nand U17888 (N_17888,N_13628,N_11184);
nand U17889 (N_17889,N_14093,N_10438);
xor U17890 (N_17890,N_10456,N_11263);
xor U17891 (N_17891,N_11878,N_14875);
or U17892 (N_17892,N_11524,N_11828);
xor U17893 (N_17893,N_11830,N_14500);
xnor U17894 (N_17894,N_11303,N_11984);
nor U17895 (N_17895,N_13490,N_14736);
and U17896 (N_17896,N_12276,N_13406);
or U17897 (N_17897,N_11752,N_12647);
or U17898 (N_17898,N_10840,N_11580);
nand U17899 (N_17899,N_13298,N_13111);
nand U17900 (N_17900,N_10259,N_14002);
xor U17901 (N_17901,N_11300,N_11930);
or U17902 (N_17902,N_12276,N_10545);
and U17903 (N_17903,N_11899,N_12860);
nor U17904 (N_17904,N_14948,N_11727);
or U17905 (N_17905,N_11096,N_12563);
nor U17906 (N_17906,N_12949,N_10703);
nor U17907 (N_17907,N_13590,N_11881);
or U17908 (N_17908,N_11404,N_12055);
nor U17909 (N_17909,N_13510,N_12679);
and U17910 (N_17910,N_11795,N_11005);
and U17911 (N_17911,N_10810,N_13551);
and U17912 (N_17912,N_13683,N_13167);
and U17913 (N_17913,N_13689,N_10320);
nand U17914 (N_17914,N_12741,N_11576);
nor U17915 (N_17915,N_12901,N_13939);
xnor U17916 (N_17916,N_12865,N_12835);
or U17917 (N_17917,N_11330,N_14900);
or U17918 (N_17918,N_10297,N_13010);
nand U17919 (N_17919,N_11748,N_13669);
xor U17920 (N_17920,N_14524,N_13836);
nor U17921 (N_17921,N_10125,N_12232);
or U17922 (N_17922,N_10662,N_10094);
nand U17923 (N_17923,N_13674,N_10536);
and U17924 (N_17924,N_10562,N_10743);
or U17925 (N_17925,N_13436,N_11550);
nand U17926 (N_17926,N_14614,N_12114);
nand U17927 (N_17927,N_12768,N_12242);
nand U17928 (N_17928,N_13729,N_13571);
or U17929 (N_17929,N_12465,N_13191);
or U17930 (N_17930,N_12711,N_13292);
nor U17931 (N_17931,N_14540,N_11721);
or U17932 (N_17932,N_14545,N_10973);
nor U17933 (N_17933,N_12157,N_12331);
or U17934 (N_17934,N_13020,N_14135);
and U17935 (N_17935,N_11187,N_11100);
xor U17936 (N_17936,N_10790,N_10306);
xor U17937 (N_17937,N_11868,N_11117);
xnor U17938 (N_17938,N_13924,N_12649);
nand U17939 (N_17939,N_12960,N_11073);
nor U17940 (N_17940,N_10684,N_14517);
nor U17941 (N_17941,N_14497,N_10214);
nand U17942 (N_17942,N_12806,N_14416);
and U17943 (N_17943,N_10825,N_10849);
nor U17944 (N_17944,N_14756,N_10161);
xor U17945 (N_17945,N_11461,N_12131);
nor U17946 (N_17946,N_11958,N_11957);
xnor U17947 (N_17947,N_14575,N_12767);
nand U17948 (N_17948,N_11259,N_13819);
xnor U17949 (N_17949,N_14302,N_12640);
or U17950 (N_17950,N_10430,N_10406);
nor U17951 (N_17951,N_12000,N_11344);
or U17952 (N_17952,N_14533,N_12999);
xnor U17953 (N_17953,N_11608,N_13290);
nand U17954 (N_17954,N_13566,N_12890);
nand U17955 (N_17955,N_13337,N_13022);
nand U17956 (N_17956,N_10423,N_14237);
xor U17957 (N_17957,N_13768,N_12462);
xnor U17958 (N_17958,N_13476,N_12692);
nand U17959 (N_17959,N_10969,N_12926);
or U17960 (N_17960,N_13736,N_13660);
nor U17961 (N_17961,N_11085,N_14760);
nor U17962 (N_17962,N_12523,N_13590);
or U17963 (N_17963,N_13344,N_14279);
nor U17964 (N_17964,N_12216,N_12415);
and U17965 (N_17965,N_10582,N_11407);
and U17966 (N_17966,N_14216,N_14778);
nor U17967 (N_17967,N_14967,N_13540);
nor U17968 (N_17968,N_13605,N_11118);
or U17969 (N_17969,N_12301,N_13779);
nand U17970 (N_17970,N_14760,N_12675);
nand U17971 (N_17971,N_13465,N_14550);
nor U17972 (N_17972,N_14779,N_11334);
or U17973 (N_17973,N_12190,N_13968);
xor U17974 (N_17974,N_11436,N_10181);
and U17975 (N_17975,N_11037,N_10025);
and U17976 (N_17976,N_14389,N_14587);
nor U17977 (N_17977,N_11699,N_12383);
nor U17978 (N_17978,N_12535,N_11350);
or U17979 (N_17979,N_10163,N_10065);
nor U17980 (N_17980,N_10485,N_14833);
nand U17981 (N_17981,N_12727,N_12234);
nor U17982 (N_17982,N_11581,N_14638);
nand U17983 (N_17983,N_13924,N_12916);
nor U17984 (N_17984,N_10167,N_14164);
nor U17985 (N_17985,N_13767,N_11848);
or U17986 (N_17986,N_10252,N_14439);
nor U17987 (N_17987,N_14231,N_10524);
or U17988 (N_17988,N_10886,N_13766);
nand U17989 (N_17989,N_13524,N_12002);
nor U17990 (N_17990,N_12480,N_12355);
nand U17991 (N_17991,N_11123,N_10514);
xnor U17992 (N_17992,N_13672,N_14397);
nor U17993 (N_17993,N_13036,N_12532);
nand U17994 (N_17994,N_10074,N_13900);
xnor U17995 (N_17995,N_13815,N_14659);
xor U17996 (N_17996,N_13385,N_14775);
nand U17997 (N_17997,N_10898,N_13629);
xor U17998 (N_17998,N_11221,N_13127);
xor U17999 (N_17999,N_14105,N_14447);
nor U18000 (N_18000,N_10709,N_10229);
xor U18001 (N_18001,N_14650,N_11846);
nor U18002 (N_18002,N_12062,N_12531);
or U18003 (N_18003,N_10087,N_13339);
and U18004 (N_18004,N_11427,N_11837);
and U18005 (N_18005,N_11949,N_12342);
and U18006 (N_18006,N_12441,N_13912);
nor U18007 (N_18007,N_11210,N_13397);
nand U18008 (N_18008,N_11308,N_11437);
nand U18009 (N_18009,N_14276,N_11298);
nand U18010 (N_18010,N_11788,N_14726);
or U18011 (N_18011,N_14619,N_11878);
nand U18012 (N_18012,N_11527,N_13928);
nand U18013 (N_18013,N_13650,N_14038);
nand U18014 (N_18014,N_12584,N_11922);
nand U18015 (N_18015,N_10437,N_13345);
xor U18016 (N_18016,N_14956,N_12465);
or U18017 (N_18017,N_14428,N_14333);
xor U18018 (N_18018,N_10292,N_13192);
and U18019 (N_18019,N_14734,N_11085);
and U18020 (N_18020,N_13247,N_14576);
nand U18021 (N_18021,N_12125,N_13476);
or U18022 (N_18022,N_12512,N_12060);
or U18023 (N_18023,N_12263,N_12664);
and U18024 (N_18024,N_13566,N_14125);
nor U18025 (N_18025,N_13483,N_13772);
or U18026 (N_18026,N_11309,N_12831);
nor U18027 (N_18027,N_10329,N_12493);
nor U18028 (N_18028,N_14744,N_10574);
xnor U18029 (N_18029,N_12502,N_10452);
and U18030 (N_18030,N_10451,N_10280);
nand U18031 (N_18031,N_10838,N_14852);
xnor U18032 (N_18032,N_14249,N_13988);
xor U18033 (N_18033,N_13566,N_11724);
nand U18034 (N_18034,N_12911,N_14366);
nand U18035 (N_18035,N_14285,N_13452);
or U18036 (N_18036,N_11964,N_10752);
nand U18037 (N_18037,N_13243,N_13676);
nor U18038 (N_18038,N_12755,N_10744);
nand U18039 (N_18039,N_10523,N_10943);
nand U18040 (N_18040,N_12904,N_11047);
nand U18041 (N_18041,N_13804,N_14965);
and U18042 (N_18042,N_11188,N_10702);
nor U18043 (N_18043,N_12879,N_13927);
nor U18044 (N_18044,N_11625,N_14654);
or U18045 (N_18045,N_13139,N_12364);
and U18046 (N_18046,N_11608,N_11945);
or U18047 (N_18047,N_12666,N_14380);
nor U18048 (N_18048,N_12339,N_12243);
and U18049 (N_18049,N_13774,N_14408);
nand U18050 (N_18050,N_10359,N_13163);
nor U18051 (N_18051,N_10233,N_14800);
xor U18052 (N_18052,N_13096,N_13720);
xnor U18053 (N_18053,N_14715,N_11206);
xor U18054 (N_18054,N_10704,N_11155);
xnor U18055 (N_18055,N_12836,N_12813);
and U18056 (N_18056,N_11222,N_12345);
xnor U18057 (N_18057,N_11425,N_14080);
and U18058 (N_18058,N_14090,N_14491);
xnor U18059 (N_18059,N_12593,N_14865);
or U18060 (N_18060,N_12327,N_11324);
xor U18061 (N_18061,N_12587,N_14509);
or U18062 (N_18062,N_11637,N_11072);
and U18063 (N_18063,N_10187,N_12062);
nand U18064 (N_18064,N_13386,N_13498);
nand U18065 (N_18065,N_12177,N_14612);
or U18066 (N_18066,N_11528,N_10662);
nor U18067 (N_18067,N_10575,N_11323);
nand U18068 (N_18068,N_14171,N_14101);
and U18069 (N_18069,N_14515,N_12683);
nor U18070 (N_18070,N_12059,N_14194);
nand U18071 (N_18071,N_12516,N_12039);
nand U18072 (N_18072,N_12945,N_12078);
or U18073 (N_18073,N_14429,N_13704);
nor U18074 (N_18074,N_13048,N_14212);
nor U18075 (N_18075,N_11156,N_10575);
or U18076 (N_18076,N_11473,N_10217);
or U18077 (N_18077,N_14428,N_13511);
xnor U18078 (N_18078,N_12458,N_12784);
nor U18079 (N_18079,N_10515,N_14345);
nand U18080 (N_18080,N_13628,N_13659);
nor U18081 (N_18081,N_14270,N_12603);
xor U18082 (N_18082,N_13024,N_13820);
nand U18083 (N_18083,N_10329,N_11430);
or U18084 (N_18084,N_14104,N_11122);
and U18085 (N_18085,N_14845,N_10495);
or U18086 (N_18086,N_10782,N_13473);
nand U18087 (N_18087,N_13706,N_12779);
nand U18088 (N_18088,N_11853,N_13560);
or U18089 (N_18089,N_13703,N_13654);
or U18090 (N_18090,N_10747,N_10630);
nor U18091 (N_18091,N_14165,N_14532);
nor U18092 (N_18092,N_10330,N_13860);
and U18093 (N_18093,N_12789,N_11453);
xnor U18094 (N_18094,N_10234,N_14685);
xor U18095 (N_18095,N_11318,N_12693);
nand U18096 (N_18096,N_10017,N_12827);
and U18097 (N_18097,N_11922,N_11331);
or U18098 (N_18098,N_14117,N_11659);
nor U18099 (N_18099,N_13445,N_12723);
nor U18100 (N_18100,N_11715,N_10166);
xor U18101 (N_18101,N_12353,N_10444);
nor U18102 (N_18102,N_10226,N_11296);
xnor U18103 (N_18103,N_11491,N_11040);
nor U18104 (N_18104,N_14728,N_11668);
nor U18105 (N_18105,N_13985,N_10224);
xor U18106 (N_18106,N_12491,N_12898);
or U18107 (N_18107,N_13342,N_10095);
or U18108 (N_18108,N_14206,N_10788);
or U18109 (N_18109,N_13861,N_11272);
nor U18110 (N_18110,N_13545,N_13350);
nor U18111 (N_18111,N_11934,N_11398);
nand U18112 (N_18112,N_10796,N_11261);
and U18113 (N_18113,N_12477,N_11576);
nand U18114 (N_18114,N_10962,N_11963);
or U18115 (N_18115,N_10957,N_14793);
nor U18116 (N_18116,N_10243,N_14034);
nand U18117 (N_18117,N_12250,N_12738);
or U18118 (N_18118,N_12510,N_10678);
xnor U18119 (N_18119,N_13222,N_11961);
nor U18120 (N_18120,N_12409,N_13982);
xnor U18121 (N_18121,N_13657,N_12489);
nand U18122 (N_18122,N_13236,N_10645);
xnor U18123 (N_18123,N_12644,N_11741);
nor U18124 (N_18124,N_12397,N_13813);
or U18125 (N_18125,N_14975,N_12457);
nand U18126 (N_18126,N_10278,N_13291);
nor U18127 (N_18127,N_12463,N_13029);
nor U18128 (N_18128,N_11803,N_14067);
nor U18129 (N_18129,N_10062,N_13442);
nand U18130 (N_18130,N_14183,N_13860);
xor U18131 (N_18131,N_12028,N_13011);
nor U18132 (N_18132,N_12560,N_14352);
xnor U18133 (N_18133,N_13140,N_11062);
xor U18134 (N_18134,N_12729,N_14032);
nand U18135 (N_18135,N_11290,N_11208);
or U18136 (N_18136,N_10034,N_13462);
xor U18137 (N_18137,N_13725,N_10713);
xor U18138 (N_18138,N_14062,N_13026);
xnor U18139 (N_18139,N_11833,N_12857);
or U18140 (N_18140,N_12520,N_10859);
nand U18141 (N_18141,N_10780,N_11267);
or U18142 (N_18142,N_14413,N_12508);
or U18143 (N_18143,N_10355,N_11131);
or U18144 (N_18144,N_14718,N_11811);
and U18145 (N_18145,N_12843,N_11778);
nor U18146 (N_18146,N_11747,N_11276);
nor U18147 (N_18147,N_14326,N_14341);
nand U18148 (N_18148,N_10074,N_11206);
nor U18149 (N_18149,N_12440,N_13081);
xnor U18150 (N_18150,N_11549,N_13574);
xor U18151 (N_18151,N_12401,N_14275);
and U18152 (N_18152,N_12229,N_12849);
xnor U18153 (N_18153,N_13275,N_13353);
xor U18154 (N_18154,N_11447,N_14091);
or U18155 (N_18155,N_12559,N_12139);
xor U18156 (N_18156,N_11308,N_10458);
or U18157 (N_18157,N_11865,N_13986);
or U18158 (N_18158,N_10758,N_13261);
xnor U18159 (N_18159,N_13632,N_14273);
nand U18160 (N_18160,N_13692,N_12554);
nor U18161 (N_18161,N_11899,N_13583);
and U18162 (N_18162,N_14434,N_11870);
or U18163 (N_18163,N_13392,N_14563);
nor U18164 (N_18164,N_14661,N_12125);
nor U18165 (N_18165,N_13727,N_13047);
xnor U18166 (N_18166,N_10895,N_12409);
nand U18167 (N_18167,N_10999,N_12753);
or U18168 (N_18168,N_11442,N_10807);
or U18169 (N_18169,N_10644,N_12007);
and U18170 (N_18170,N_10784,N_13677);
or U18171 (N_18171,N_10220,N_12752);
or U18172 (N_18172,N_12770,N_14230);
and U18173 (N_18173,N_11523,N_11533);
nand U18174 (N_18174,N_11163,N_13775);
or U18175 (N_18175,N_11050,N_11002);
xor U18176 (N_18176,N_14158,N_14558);
nor U18177 (N_18177,N_14257,N_14058);
xor U18178 (N_18178,N_13534,N_13928);
and U18179 (N_18179,N_12303,N_12700);
or U18180 (N_18180,N_14861,N_11995);
xnor U18181 (N_18181,N_10131,N_14296);
nor U18182 (N_18182,N_10379,N_11018);
nand U18183 (N_18183,N_14599,N_11947);
nand U18184 (N_18184,N_10625,N_13903);
and U18185 (N_18185,N_13791,N_13191);
or U18186 (N_18186,N_13734,N_13922);
and U18187 (N_18187,N_12874,N_12024);
and U18188 (N_18188,N_11693,N_12189);
or U18189 (N_18189,N_11956,N_10885);
nand U18190 (N_18190,N_10251,N_10861);
nor U18191 (N_18191,N_10232,N_13402);
nand U18192 (N_18192,N_10059,N_13064);
or U18193 (N_18193,N_11299,N_11264);
xnor U18194 (N_18194,N_11748,N_14468);
xor U18195 (N_18195,N_11172,N_10771);
xor U18196 (N_18196,N_13771,N_14109);
nand U18197 (N_18197,N_13274,N_12096);
xor U18198 (N_18198,N_10765,N_10101);
xnor U18199 (N_18199,N_12076,N_12345);
nor U18200 (N_18200,N_10699,N_12996);
nor U18201 (N_18201,N_11451,N_13030);
nor U18202 (N_18202,N_12731,N_10465);
nand U18203 (N_18203,N_10781,N_12780);
and U18204 (N_18204,N_12561,N_14293);
nand U18205 (N_18205,N_13910,N_10352);
nor U18206 (N_18206,N_10159,N_11576);
nand U18207 (N_18207,N_14039,N_12523);
and U18208 (N_18208,N_10154,N_14124);
nor U18209 (N_18209,N_11925,N_14571);
nand U18210 (N_18210,N_12428,N_10250);
nand U18211 (N_18211,N_14104,N_11840);
and U18212 (N_18212,N_12368,N_12939);
or U18213 (N_18213,N_14268,N_12641);
and U18214 (N_18214,N_11891,N_13841);
nor U18215 (N_18215,N_11355,N_11357);
or U18216 (N_18216,N_11887,N_11575);
nand U18217 (N_18217,N_14357,N_13318);
xor U18218 (N_18218,N_14919,N_14368);
or U18219 (N_18219,N_11032,N_13061);
xnor U18220 (N_18220,N_13158,N_12836);
or U18221 (N_18221,N_12167,N_12992);
nand U18222 (N_18222,N_12501,N_14542);
nor U18223 (N_18223,N_11497,N_12553);
xnor U18224 (N_18224,N_11410,N_11054);
and U18225 (N_18225,N_13534,N_11836);
and U18226 (N_18226,N_11076,N_14802);
or U18227 (N_18227,N_14432,N_14192);
nand U18228 (N_18228,N_13639,N_10764);
and U18229 (N_18229,N_11903,N_10005);
and U18230 (N_18230,N_12991,N_11431);
and U18231 (N_18231,N_12039,N_10082);
nor U18232 (N_18232,N_11465,N_11017);
or U18233 (N_18233,N_11130,N_13179);
xor U18234 (N_18234,N_13563,N_14043);
xnor U18235 (N_18235,N_12370,N_14821);
and U18236 (N_18236,N_13731,N_10151);
nor U18237 (N_18237,N_10598,N_14635);
and U18238 (N_18238,N_10574,N_14334);
xor U18239 (N_18239,N_14903,N_11335);
xor U18240 (N_18240,N_11115,N_11196);
or U18241 (N_18241,N_11928,N_12559);
or U18242 (N_18242,N_10256,N_10015);
or U18243 (N_18243,N_14688,N_11693);
nor U18244 (N_18244,N_11029,N_10981);
nor U18245 (N_18245,N_14752,N_14595);
or U18246 (N_18246,N_14974,N_11873);
nor U18247 (N_18247,N_10476,N_10724);
or U18248 (N_18248,N_11377,N_13876);
xnor U18249 (N_18249,N_12920,N_14101);
xnor U18250 (N_18250,N_11685,N_12589);
nor U18251 (N_18251,N_12415,N_14861);
xor U18252 (N_18252,N_13392,N_12934);
nor U18253 (N_18253,N_13820,N_11698);
nor U18254 (N_18254,N_14719,N_13112);
xor U18255 (N_18255,N_12306,N_13162);
xor U18256 (N_18256,N_11877,N_11860);
xor U18257 (N_18257,N_12154,N_14517);
and U18258 (N_18258,N_14000,N_13387);
and U18259 (N_18259,N_13890,N_13937);
xnor U18260 (N_18260,N_13113,N_14898);
nand U18261 (N_18261,N_12853,N_13514);
xor U18262 (N_18262,N_13359,N_12265);
and U18263 (N_18263,N_14048,N_11097);
xor U18264 (N_18264,N_14554,N_13211);
nand U18265 (N_18265,N_11914,N_11414);
nand U18266 (N_18266,N_12137,N_12378);
or U18267 (N_18267,N_12480,N_10228);
nand U18268 (N_18268,N_11049,N_12642);
xor U18269 (N_18269,N_10199,N_13408);
or U18270 (N_18270,N_13280,N_10822);
nand U18271 (N_18271,N_13048,N_14796);
or U18272 (N_18272,N_14423,N_12272);
or U18273 (N_18273,N_14013,N_10036);
xnor U18274 (N_18274,N_11126,N_10982);
or U18275 (N_18275,N_14806,N_10522);
and U18276 (N_18276,N_12040,N_11396);
nand U18277 (N_18277,N_14886,N_11330);
or U18278 (N_18278,N_10817,N_11898);
nor U18279 (N_18279,N_11062,N_13446);
or U18280 (N_18280,N_13598,N_13413);
nor U18281 (N_18281,N_14027,N_11362);
nor U18282 (N_18282,N_10306,N_12854);
nand U18283 (N_18283,N_12325,N_13485);
nor U18284 (N_18284,N_12894,N_10420);
nand U18285 (N_18285,N_13340,N_13862);
and U18286 (N_18286,N_14136,N_10140);
xnor U18287 (N_18287,N_11230,N_14066);
nand U18288 (N_18288,N_13641,N_11752);
nand U18289 (N_18289,N_13780,N_14306);
nor U18290 (N_18290,N_10153,N_11650);
nor U18291 (N_18291,N_13788,N_11325);
or U18292 (N_18292,N_13833,N_14667);
xnor U18293 (N_18293,N_11429,N_13010);
or U18294 (N_18294,N_13803,N_14883);
nand U18295 (N_18295,N_14549,N_10599);
xnor U18296 (N_18296,N_12513,N_14325);
and U18297 (N_18297,N_11209,N_12115);
xor U18298 (N_18298,N_11662,N_14897);
nor U18299 (N_18299,N_11387,N_11034);
xnor U18300 (N_18300,N_12327,N_14337);
nand U18301 (N_18301,N_13742,N_13892);
and U18302 (N_18302,N_11648,N_10399);
xnor U18303 (N_18303,N_14054,N_13931);
xor U18304 (N_18304,N_12904,N_12754);
nand U18305 (N_18305,N_13034,N_13252);
and U18306 (N_18306,N_12306,N_12500);
and U18307 (N_18307,N_11557,N_12878);
nand U18308 (N_18308,N_13411,N_12780);
nor U18309 (N_18309,N_11271,N_14458);
nor U18310 (N_18310,N_12272,N_11274);
and U18311 (N_18311,N_13006,N_10926);
xor U18312 (N_18312,N_12090,N_10844);
xnor U18313 (N_18313,N_10722,N_13044);
or U18314 (N_18314,N_14186,N_12608);
nand U18315 (N_18315,N_10947,N_14365);
nor U18316 (N_18316,N_14263,N_11262);
nand U18317 (N_18317,N_12161,N_10801);
nor U18318 (N_18318,N_11611,N_14639);
and U18319 (N_18319,N_10550,N_14772);
xnor U18320 (N_18320,N_12648,N_10632);
xor U18321 (N_18321,N_12203,N_11801);
nor U18322 (N_18322,N_13602,N_12116);
nor U18323 (N_18323,N_14139,N_11860);
or U18324 (N_18324,N_14563,N_10525);
and U18325 (N_18325,N_14962,N_13131);
or U18326 (N_18326,N_13079,N_12001);
and U18327 (N_18327,N_11347,N_10779);
nand U18328 (N_18328,N_13035,N_11913);
xor U18329 (N_18329,N_13973,N_10461);
nand U18330 (N_18330,N_13813,N_11949);
and U18331 (N_18331,N_11522,N_14958);
nand U18332 (N_18332,N_10047,N_11687);
and U18333 (N_18333,N_11739,N_14229);
or U18334 (N_18334,N_13239,N_11710);
nor U18335 (N_18335,N_10779,N_13147);
and U18336 (N_18336,N_10517,N_13956);
or U18337 (N_18337,N_12446,N_14997);
nor U18338 (N_18338,N_14226,N_11291);
nand U18339 (N_18339,N_10490,N_11417);
and U18340 (N_18340,N_11856,N_10862);
nand U18341 (N_18341,N_13309,N_13966);
and U18342 (N_18342,N_12122,N_13119);
nor U18343 (N_18343,N_14624,N_12899);
nor U18344 (N_18344,N_13485,N_10475);
nand U18345 (N_18345,N_11632,N_10840);
and U18346 (N_18346,N_14777,N_10453);
xnor U18347 (N_18347,N_10805,N_14180);
nor U18348 (N_18348,N_10607,N_10660);
nand U18349 (N_18349,N_11823,N_14297);
or U18350 (N_18350,N_10015,N_13446);
nand U18351 (N_18351,N_14298,N_13691);
nor U18352 (N_18352,N_11823,N_11393);
nor U18353 (N_18353,N_11120,N_13790);
nor U18354 (N_18354,N_13514,N_10847);
nor U18355 (N_18355,N_10352,N_14044);
or U18356 (N_18356,N_11273,N_12387);
and U18357 (N_18357,N_14727,N_11433);
or U18358 (N_18358,N_12652,N_12438);
nand U18359 (N_18359,N_13801,N_11073);
and U18360 (N_18360,N_12815,N_10103);
or U18361 (N_18361,N_11730,N_11329);
nand U18362 (N_18362,N_12264,N_14482);
xor U18363 (N_18363,N_14691,N_12489);
or U18364 (N_18364,N_12460,N_10738);
or U18365 (N_18365,N_12098,N_14909);
and U18366 (N_18366,N_14116,N_14888);
nand U18367 (N_18367,N_11758,N_11122);
xnor U18368 (N_18368,N_11176,N_11440);
or U18369 (N_18369,N_14792,N_11074);
xnor U18370 (N_18370,N_14466,N_14747);
and U18371 (N_18371,N_13236,N_14696);
nand U18372 (N_18372,N_10703,N_11146);
and U18373 (N_18373,N_14403,N_13556);
xor U18374 (N_18374,N_12809,N_11424);
xor U18375 (N_18375,N_14989,N_10710);
nand U18376 (N_18376,N_10110,N_12999);
and U18377 (N_18377,N_10602,N_14867);
and U18378 (N_18378,N_12146,N_14322);
and U18379 (N_18379,N_11755,N_11392);
nand U18380 (N_18380,N_10298,N_13055);
or U18381 (N_18381,N_11754,N_12970);
and U18382 (N_18382,N_10317,N_12436);
xnor U18383 (N_18383,N_14081,N_14292);
xor U18384 (N_18384,N_10784,N_10440);
nor U18385 (N_18385,N_13689,N_10846);
and U18386 (N_18386,N_12441,N_12963);
xor U18387 (N_18387,N_13523,N_12073);
nand U18388 (N_18388,N_14133,N_13509);
nand U18389 (N_18389,N_12231,N_12279);
xor U18390 (N_18390,N_11181,N_11182);
and U18391 (N_18391,N_12817,N_10286);
nand U18392 (N_18392,N_13600,N_11909);
or U18393 (N_18393,N_14186,N_11227);
nand U18394 (N_18394,N_14440,N_13458);
nor U18395 (N_18395,N_13300,N_11077);
and U18396 (N_18396,N_11886,N_13014);
xnor U18397 (N_18397,N_13366,N_11982);
nor U18398 (N_18398,N_14168,N_14216);
nand U18399 (N_18399,N_10366,N_11639);
xnor U18400 (N_18400,N_12574,N_13728);
or U18401 (N_18401,N_10479,N_11930);
or U18402 (N_18402,N_14614,N_12908);
nor U18403 (N_18403,N_11937,N_11560);
nand U18404 (N_18404,N_14680,N_10394);
and U18405 (N_18405,N_13505,N_11896);
or U18406 (N_18406,N_11273,N_14606);
or U18407 (N_18407,N_10196,N_14551);
and U18408 (N_18408,N_10765,N_14298);
or U18409 (N_18409,N_10764,N_14061);
and U18410 (N_18410,N_11700,N_10461);
or U18411 (N_18411,N_11067,N_10130);
and U18412 (N_18412,N_11396,N_10259);
nor U18413 (N_18413,N_14331,N_14839);
nand U18414 (N_18414,N_14579,N_10608);
nand U18415 (N_18415,N_11547,N_12097);
and U18416 (N_18416,N_11191,N_11803);
xnor U18417 (N_18417,N_13432,N_11791);
nand U18418 (N_18418,N_11988,N_10385);
xnor U18419 (N_18419,N_14919,N_13202);
xor U18420 (N_18420,N_10077,N_12532);
or U18421 (N_18421,N_10022,N_14291);
nor U18422 (N_18422,N_14435,N_13870);
xnor U18423 (N_18423,N_10561,N_12416);
nand U18424 (N_18424,N_14160,N_13892);
or U18425 (N_18425,N_11750,N_11565);
xor U18426 (N_18426,N_10722,N_11770);
nor U18427 (N_18427,N_11764,N_11078);
xor U18428 (N_18428,N_11438,N_10483);
xnor U18429 (N_18429,N_12469,N_12718);
xor U18430 (N_18430,N_13763,N_11607);
nor U18431 (N_18431,N_12975,N_13507);
nor U18432 (N_18432,N_11809,N_13297);
or U18433 (N_18433,N_12691,N_10863);
or U18434 (N_18434,N_11396,N_13228);
nor U18435 (N_18435,N_14367,N_11112);
or U18436 (N_18436,N_10462,N_13016);
and U18437 (N_18437,N_14932,N_11739);
or U18438 (N_18438,N_14061,N_12565);
or U18439 (N_18439,N_12693,N_13692);
or U18440 (N_18440,N_13011,N_10740);
nand U18441 (N_18441,N_10813,N_12504);
or U18442 (N_18442,N_10229,N_11709);
and U18443 (N_18443,N_13213,N_13999);
xor U18444 (N_18444,N_13077,N_12923);
nor U18445 (N_18445,N_13897,N_12702);
nor U18446 (N_18446,N_11993,N_12036);
nand U18447 (N_18447,N_10149,N_14610);
nand U18448 (N_18448,N_12743,N_11065);
nor U18449 (N_18449,N_14186,N_13146);
and U18450 (N_18450,N_11268,N_14312);
and U18451 (N_18451,N_10313,N_13672);
nand U18452 (N_18452,N_14996,N_12857);
nor U18453 (N_18453,N_10275,N_10709);
xnor U18454 (N_18454,N_13170,N_11541);
and U18455 (N_18455,N_13560,N_14503);
xnor U18456 (N_18456,N_10912,N_10142);
or U18457 (N_18457,N_10674,N_14186);
nor U18458 (N_18458,N_13448,N_14511);
nand U18459 (N_18459,N_11790,N_14640);
xor U18460 (N_18460,N_11501,N_14938);
xor U18461 (N_18461,N_12954,N_10366);
xor U18462 (N_18462,N_13177,N_14568);
and U18463 (N_18463,N_11633,N_11552);
nor U18464 (N_18464,N_10822,N_10061);
or U18465 (N_18465,N_10763,N_11914);
nand U18466 (N_18466,N_14754,N_12498);
xnor U18467 (N_18467,N_14725,N_11563);
and U18468 (N_18468,N_12858,N_10915);
xor U18469 (N_18469,N_10850,N_12653);
and U18470 (N_18470,N_14050,N_10905);
xor U18471 (N_18471,N_14613,N_12679);
or U18472 (N_18472,N_13664,N_10407);
or U18473 (N_18473,N_14997,N_14117);
xnor U18474 (N_18474,N_13278,N_14212);
xor U18475 (N_18475,N_10055,N_10971);
or U18476 (N_18476,N_13903,N_12287);
nand U18477 (N_18477,N_13766,N_10949);
and U18478 (N_18478,N_13496,N_10958);
xor U18479 (N_18479,N_10410,N_13631);
nand U18480 (N_18480,N_14620,N_12482);
nor U18481 (N_18481,N_13421,N_13717);
nor U18482 (N_18482,N_13376,N_11558);
and U18483 (N_18483,N_13471,N_11362);
xnor U18484 (N_18484,N_13892,N_13088);
or U18485 (N_18485,N_11109,N_13759);
and U18486 (N_18486,N_14596,N_12062);
nand U18487 (N_18487,N_12637,N_10807);
and U18488 (N_18488,N_11289,N_14530);
or U18489 (N_18489,N_14751,N_14508);
xnor U18490 (N_18490,N_13044,N_11035);
or U18491 (N_18491,N_11424,N_11923);
xor U18492 (N_18492,N_13309,N_14875);
and U18493 (N_18493,N_13038,N_11431);
nand U18494 (N_18494,N_14792,N_14944);
xor U18495 (N_18495,N_10251,N_11254);
xor U18496 (N_18496,N_13693,N_13385);
xnor U18497 (N_18497,N_14173,N_11551);
or U18498 (N_18498,N_12223,N_13543);
and U18499 (N_18499,N_10285,N_14363);
and U18500 (N_18500,N_13039,N_14663);
nand U18501 (N_18501,N_10119,N_10061);
xnor U18502 (N_18502,N_14722,N_10726);
nand U18503 (N_18503,N_14615,N_12204);
and U18504 (N_18504,N_14069,N_10495);
nor U18505 (N_18505,N_11376,N_13014);
and U18506 (N_18506,N_14455,N_13771);
and U18507 (N_18507,N_10532,N_14044);
and U18508 (N_18508,N_14101,N_10452);
nand U18509 (N_18509,N_12639,N_10508);
xor U18510 (N_18510,N_12995,N_10155);
xor U18511 (N_18511,N_11188,N_11750);
nor U18512 (N_18512,N_10827,N_12357);
xnor U18513 (N_18513,N_13714,N_14002);
nor U18514 (N_18514,N_10013,N_10586);
nor U18515 (N_18515,N_11274,N_13598);
nor U18516 (N_18516,N_13381,N_10637);
nor U18517 (N_18517,N_10150,N_10729);
or U18518 (N_18518,N_14453,N_10042);
nor U18519 (N_18519,N_10168,N_13605);
nor U18520 (N_18520,N_13946,N_13397);
nor U18521 (N_18521,N_14781,N_10208);
nand U18522 (N_18522,N_12711,N_10001);
or U18523 (N_18523,N_10007,N_11144);
nand U18524 (N_18524,N_14303,N_11171);
nand U18525 (N_18525,N_11523,N_12712);
or U18526 (N_18526,N_13147,N_13839);
nand U18527 (N_18527,N_10562,N_14206);
or U18528 (N_18528,N_10732,N_12929);
nor U18529 (N_18529,N_13703,N_13219);
nor U18530 (N_18530,N_12256,N_14618);
nand U18531 (N_18531,N_11238,N_11969);
nor U18532 (N_18532,N_14558,N_14728);
nand U18533 (N_18533,N_12368,N_12033);
nor U18534 (N_18534,N_12579,N_14140);
xnor U18535 (N_18535,N_14162,N_12356);
xor U18536 (N_18536,N_11820,N_10456);
nor U18537 (N_18537,N_11093,N_13018);
and U18538 (N_18538,N_11015,N_12158);
nand U18539 (N_18539,N_13191,N_14534);
xnor U18540 (N_18540,N_10918,N_14218);
and U18541 (N_18541,N_14404,N_10087);
nor U18542 (N_18542,N_11344,N_11989);
and U18543 (N_18543,N_11870,N_13891);
nor U18544 (N_18544,N_11002,N_12370);
or U18545 (N_18545,N_10950,N_11460);
xnor U18546 (N_18546,N_10094,N_10289);
or U18547 (N_18547,N_13872,N_10592);
and U18548 (N_18548,N_14887,N_12045);
or U18549 (N_18549,N_14209,N_12027);
nor U18550 (N_18550,N_12254,N_10535);
nand U18551 (N_18551,N_14169,N_14805);
and U18552 (N_18552,N_13704,N_11593);
nand U18553 (N_18553,N_11667,N_13816);
nand U18554 (N_18554,N_14447,N_11279);
nand U18555 (N_18555,N_10600,N_10423);
xor U18556 (N_18556,N_14975,N_14454);
or U18557 (N_18557,N_11071,N_13773);
and U18558 (N_18558,N_11576,N_12854);
or U18559 (N_18559,N_13249,N_13710);
nor U18560 (N_18560,N_12236,N_11301);
or U18561 (N_18561,N_12366,N_10425);
and U18562 (N_18562,N_13104,N_10960);
xnor U18563 (N_18563,N_10215,N_11729);
xnor U18564 (N_18564,N_10142,N_13121);
nand U18565 (N_18565,N_14066,N_10328);
and U18566 (N_18566,N_10850,N_11732);
and U18567 (N_18567,N_13557,N_13177);
xor U18568 (N_18568,N_10930,N_11166);
and U18569 (N_18569,N_13658,N_14656);
xnor U18570 (N_18570,N_13127,N_13646);
nor U18571 (N_18571,N_13218,N_14573);
and U18572 (N_18572,N_11912,N_11251);
and U18573 (N_18573,N_13847,N_14829);
and U18574 (N_18574,N_12878,N_14607);
or U18575 (N_18575,N_11668,N_13267);
nand U18576 (N_18576,N_11649,N_11102);
nor U18577 (N_18577,N_10151,N_10436);
xnor U18578 (N_18578,N_10964,N_14940);
xor U18579 (N_18579,N_13601,N_10137);
nor U18580 (N_18580,N_13434,N_14841);
or U18581 (N_18581,N_14962,N_11938);
xor U18582 (N_18582,N_10608,N_12260);
nor U18583 (N_18583,N_13380,N_10709);
or U18584 (N_18584,N_13772,N_10845);
xor U18585 (N_18585,N_13039,N_12683);
nor U18586 (N_18586,N_13900,N_12239);
nand U18587 (N_18587,N_11187,N_11522);
xnor U18588 (N_18588,N_10377,N_12593);
nor U18589 (N_18589,N_11147,N_12163);
xor U18590 (N_18590,N_11580,N_11164);
nand U18591 (N_18591,N_13794,N_11604);
or U18592 (N_18592,N_14329,N_13903);
xnor U18593 (N_18593,N_11265,N_12079);
or U18594 (N_18594,N_11942,N_10967);
nor U18595 (N_18595,N_11197,N_12513);
nand U18596 (N_18596,N_13587,N_12561);
nand U18597 (N_18597,N_10336,N_12580);
nand U18598 (N_18598,N_12056,N_12160);
and U18599 (N_18599,N_11541,N_11246);
xnor U18600 (N_18600,N_13061,N_10141);
xor U18601 (N_18601,N_13216,N_10898);
xnor U18602 (N_18602,N_12151,N_14611);
nor U18603 (N_18603,N_13388,N_12394);
xor U18604 (N_18604,N_11680,N_11960);
nand U18605 (N_18605,N_10047,N_12976);
and U18606 (N_18606,N_10057,N_11983);
nand U18607 (N_18607,N_12393,N_13045);
nand U18608 (N_18608,N_11782,N_12494);
nand U18609 (N_18609,N_13695,N_13491);
xor U18610 (N_18610,N_11780,N_14247);
nand U18611 (N_18611,N_12691,N_12682);
xnor U18612 (N_18612,N_10845,N_11561);
or U18613 (N_18613,N_10228,N_12743);
nand U18614 (N_18614,N_14186,N_13099);
and U18615 (N_18615,N_10122,N_14400);
or U18616 (N_18616,N_12544,N_12900);
nor U18617 (N_18617,N_11930,N_14833);
or U18618 (N_18618,N_14758,N_12191);
nand U18619 (N_18619,N_13653,N_12803);
nor U18620 (N_18620,N_14971,N_10775);
or U18621 (N_18621,N_14163,N_11708);
or U18622 (N_18622,N_10498,N_11243);
or U18623 (N_18623,N_13176,N_13424);
nand U18624 (N_18624,N_13910,N_11749);
nand U18625 (N_18625,N_10681,N_14033);
and U18626 (N_18626,N_14782,N_11598);
or U18627 (N_18627,N_12176,N_11781);
or U18628 (N_18628,N_14681,N_11260);
or U18629 (N_18629,N_11798,N_12833);
or U18630 (N_18630,N_10751,N_11531);
and U18631 (N_18631,N_13312,N_14381);
xnor U18632 (N_18632,N_10827,N_12648);
and U18633 (N_18633,N_10462,N_11810);
nor U18634 (N_18634,N_12670,N_14749);
xnor U18635 (N_18635,N_12949,N_13792);
or U18636 (N_18636,N_11815,N_10029);
nand U18637 (N_18637,N_14708,N_12024);
xor U18638 (N_18638,N_11925,N_10649);
nor U18639 (N_18639,N_13951,N_14928);
or U18640 (N_18640,N_12801,N_11248);
or U18641 (N_18641,N_14953,N_12554);
xnor U18642 (N_18642,N_13212,N_10732);
or U18643 (N_18643,N_11829,N_10299);
or U18644 (N_18644,N_14343,N_12642);
xor U18645 (N_18645,N_10975,N_10478);
and U18646 (N_18646,N_13264,N_11341);
xor U18647 (N_18647,N_13972,N_13611);
nor U18648 (N_18648,N_12756,N_11514);
nor U18649 (N_18649,N_11640,N_12123);
nand U18650 (N_18650,N_14767,N_13463);
nor U18651 (N_18651,N_14994,N_13335);
nor U18652 (N_18652,N_13577,N_12218);
nor U18653 (N_18653,N_12272,N_10800);
nand U18654 (N_18654,N_10778,N_10797);
or U18655 (N_18655,N_14358,N_11296);
and U18656 (N_18656,N_11806,N_12143);
xor U18657 (N_18657,N_12823,N_14881);
nor U18658 (N_18658,N_12182,N_12125);
or U18659 (N_18659,N_13575,N_10767);
or U18660 (N_18660,N_10587,N_12497);
or U18661 (N_18661,N_11456,N_13992);
and U18662 (N_18662,N_12828,N_11077);
and U18663 (N_18663,N_13167,N_10167);
nand U18664 (N_18664,N_10021,N_12233);
nand U18665 (N_18665,N_12419,N_10259);
and U18666 (N_18666,N_10685,N_14938);
nand U18667 (N_18667,N_13103,N_12389);
nor U18668 (N_18668,N_10010,N_14705);
nand U18669 (N_18669,N_13198,N_10149);
nor U18670 (N_18670,N_11212,N_14154);
and U18671 (N_18671,N_12511,N_10208);
nor U18672 (N_18672,N_10381,N_10239);
nor U18673 (N_18673,N_10353,N_12711);
or U18674 (N_18674,N_14282,N_14185);
and U18675 (N_18675,N_10085,N_10106);
nor U18676 (N_18676,N_13919,N_10106);
and U18677 (N_18677,N_14619,N_11644);
xnor U18678 (N_18678,N_14889,N_10507);
nor U18679 (N_18679,N_14975,N_12258);
and U18680 (N_18680,N_10955,N_13296);
nand U18681 (N_18681,N_10092,N_12000);
xnor U18682 (N_18682,N_12826,N_14260);
or U18683 (N_18683,N_14306,N_13587);
xor U18684 (N_18684,N_13890,N_11075);
and U18685 (N_18685,N_14238,N_13281);
nor U18686 (N_18686,N_14121,N_11669);
nand U18687 (N_18687,N_11062,N_13184);
nand U18688 (N_18688,N_14211,N_14367);
nor U18689 (N_18689,N_11639,N_10738);
or U18690 (N_18690,N_13915,N_10522);
xor U18691 (N_18691,N_14474,N_10062);
or U18692 (N_18692,N_10859,N_11821);
nor U18693 (N_18693,N_10923,N_14121);
xor U18694 (N_18694,N_12595,N_12374);
xnor U18695 (N_18695,N_13960,N_10745);
and U18696 (N_18696,N_12511,N_11096);
nor U18697 (N_18697,N_13508,N_12608);
xnor U18698 (N_18698,N_12268,N_14945);
or U18699 (N_18699,N_12534,N_11634);
nand U18700 (N_18700,N_12301,N_12372);
xor U18701 (N_18701,N_13549,N_13020);
nor U18702 (N_18702,N_10652,N_11035);
nand U18703 (N_18703,N_12474,N_10296);
xnor U18704 (N_18704,N_12297,N_10463);
or U18705 (N_18705,N_10784,N_14785);
nor U18706 (N_18706,N_14987,N_11145);
nand U18707 (N_18707,N_13664,N_10984);
xnor U18708 (N_18708,N_13534,N_14155);
or U18709 (N_18709,N_10252,N_10194);
and U18710 (N_18710,N_13056,N_12833);
nor U18711 (N_18711,N_11886,N_10613);
xor U18712 (N_18712,N_11827,N_14725);
nand U18713 (N_18713,N_13377,N_10569);
nand U18714 (N_18714,N_11988,N_14400);
nor U18715 (N_18715,N_10015,N_13070);
and U18716 (N_18716,N_11228,N_13676);
and U18717 (N_18717,N_13483,N_10502);
and U18718 (N_18718,N_12489,N_11008);
and U18719 (N_18719,N_10099,N_13032);
and U18720 (N_18720,N_11771,N_12701);
xnor U18721 (N_18721,N_10197,N_11574);
and U18722 (N_18722,N_11200,N_12590);
nand U18723 (N_18723,N_13727,N_13238);
nand U18724 (N_18724,N_12913,N_10344);
nand U18725 (N_18725,N_14141,N_10041);
nor U18726 (N_18726,N_13204,N_10662);
nand U18727 (N_18727,N_14124,N_14133);
nor U18728 (N_18728,N_12380,N_10722);
nand U18729 (N_18729,N_10755,N_14453);
nand U18730 (N_18730,N_10990,N_11645);
nor U18731 (N_18731,N_10407,N_13048);
or U18732 (N_18732,N_14230,N_10791);
nor U18733 (N_18733,N_13079,N_13448);
nand U18734 (N_18734,N_13599,N_11653);
xor U18735 (N_18735,N_13883,N_13081);
and U18736 (N_18736,N_12141,N_10855);
or U18737 (N_18737,N_12978,N_11954);
xnor U18738 (N_18738,N_14304,N_10284);
and U18739 (N_18739,N_10455,N_14481);
and U18740 (N_18740,N_12478,N_10981);
and U18741 (N_18741,N_14587,N_14937);
and U18742 (N_18742,N_12117,N_14918);
or U18743 (N_18743,N_14279,N_10808);
nand U18744 (N_18744,N_12568,N_12384);
nand U18745 (N_18745,N_12256,N_14373);
and U18746 (N_18746,N_11205,N_12066);
and U18747 (N_18747,N_11707,N_11873);
xnor U18748 (N_18748,N_12015,N_13053);
and U18749 (N_18749,N_11265,N_12780);
nor U18750 (N_18750,N_12609,N_11901);
xor U18751 (N_18751,N_10254,N_10550);
and U18752 (N_18752,N_13228,N_12802);
and U18753 (N_18753,N_10841,N_13584);
xnor U18754 (N_18754,N_13909,N_10150);
or U18755 (N_18755,N_14502,N_12341);
nand U18756 (N_18756,N_13668,N_12850);
nand U18757 (N_18757,N_10675,N_12654);
xnor U18758 (N_18758,N_14555,N_10911);
nand U18759 (N_18759,N_12359,N_13562);
and U18760 (N_18760,N_10635,N_10262);
nor U18761 (N_18761,N_10754,N_10211);
nor U18762 (N_18762,N_13693,N_14397);
and U18763 (N_18763,N_14795,N_10780);
or U18764 (N_18764,N_13930,N_10431);
nor U18765 (N_18765,N_14917,N_14767);
and U18766 (N_18766,N_13696,N_10531);
nand U18767 (N_18767,N_14012,N_14409);
or U18768 (N_18768,N_14119,N_13252);
and U18769 (N_18769,N_13807,N_13018);
nor U18770 (N_18770,N_11093,N_14041);
nand U18771 (N_18771,N_10914,N_10858);
or U18772 (N_18772,N_14774,N_12182);
xor U18773 (N_18773,N_12826,N_10092);
nand U18774 (N_18774,N_10503,N_12650);
nor U18775 (N_18775,N_10829,N_13789);
nor U18776 (N_18776,N_10646,N_10278);
nor U18777 (N_18777,N_10699,N_10849);
and U18778 (N_18778,N_12654,N_12689);
and U18779 (N_18779,N_14132,N_13580);
xor U18780 (N_18780,N_12656,N_10536);
or U18781 (N_18781,N_13228,N_14456);
nand U18782 (N_18782,N_13043,N_10358);
or U18783 (N_18783,N_14049,N_13324);
or U18784 (N_18784,N_13456,N_14039);
nand U18785 (N_18785,N_11511,N_14895);
and U18786 (N_18786,N_13571,N_12400);
and U18787 (N_18787,N_14272,N_10913);
nand U18788 (N_18788,N_14300,N_13689);
nand U18789 (N_18789,N_11911,N_14929);
nand U18790 (N_18790,N_12921,N_12838);
and U18791 (N_18791,N_14882,N_12808);
nor U18792 (N_18792,N_14533,N_14065);
and U18793 (N_18793,N_12227,N_12094);
nor U18794 (N_18794,N_12673,N_11607);
or U18795 (N_18795,N_10724,N_10310);
nand U18796 (N_18796,N_13588,N_12624);
nor U18797 (N_18797,N_13521,N_11045);
or U18798 (N_18798,N_13352,N_11576);
nand U18799 (N_18799,N_10446,N_11190);
xor U18800 (N_18800,N_10390,N_12006);
nor U18801 (N_18801,N_12729,N_14020);
xor U18802 (N_18802,N_12098,N_10049);
or U18803 (N_18803,N_10129,N_11977);
nor U18804 (N_18804,N_13145,N_12621);
nand U18805 (N_18805,N_13088,N_14968);
nor U18806 (N_18806,N_12240,N_14420);
or U18807 (N_18807,N_13907,N_12661);
xnor U18808 (N_18808,N_13611,N_10782);
xnor U18809 (N_18809,N_12452,N_14543);
or U18810 (N_18810,N_12763,N_14518);
and U18811 (N_18811,N_13903,N_10716);
or U18812 (N_18812,N_11591,N_10829);
nor U18813 (N_18813,N_14109,N_12823);
nand U18814 (N_18814,N_12685,N_11609);
nand U18815 (N_18815,N_11970,N_12365);
or U18816 (N_18816,N_12135,N_13031);
xnor U18817 (N_18817,N_12881,N_14666);
or U18818 (N_18818,N_12573,N_12693);
nand U18819 (N_18819,N_12049,N_14393);
nor U18820 (N_18820,N_13115,N_14909);
and U18821 (N_18821,N_14025,N_10334);
nor U18822 (N_18822,N_13572,N_11816);
nand U18823 (N_18823,N_13550,N_12090);
nor U18824 (N_18824,N_12017,N_14365);
nand U18825 (N_18825,N_13096,N_13741);
nor U18826 (N_18826,N_13576,N_13591);
nor U18827 (N_18827,N_13758,N_13752);
xor U18828 (N_18828,N_10367,N_12923);
nand U18829 (N_18829,N_10830,N_11875);
or U18830 (N_18830,N_12736,N_12255);
nor U18831 (N_18831,N_14256,N_12642);
xor U18832 (N_18832,N_12217,N_10373);
xnor U18833 (N_18833,N_14419,N_10844);
and U18834 (N_18834,N_12274,N_13762);
or U18835 (N_18835,N_11512,N_11488);
or U18836 (N_18836,N_12911,N_12411);
xnor U18837 (N_18837,N_10436,N_12721);
and U18838 (N_18838,N_11771,N_13870);
nand U18839 (N_18839,N_13182,N_11178);
and U18840 (N_18840,N_13673,N_10461);
and U18841 (N_18841,N_12149,N_14557);
nor U18842 (N_18842,N_13142,N_13360);
nand U18843 (N_18843,N_12110,N_14369);
and U18844 (N_18844,N_11176,N_10267);
or U18845 (N_18845,N_12291,N_10022);
xor U18846 (N_18846,N_13374,N_11074);
or U18847 (N_18847,N_11412,N_11955);
and U18848 (N_18848,N_11563,N_11815);
nand U18849 (N_18849,N_10225,N_11674);
nand U18850 (N_18850,N_14145,N_11332);
xor U18851 (N_18851,N_12038,N_13373);
nand U18852 (N_18852,N_12152,N_13685);
and U18853 (N_18853,N_10024,N_13912);
xnor U18854 (N_18854,N_12692,N_13290);
nor U18855 (N_18855,N_13730,N_12541);
or U18856 (N_18856,N_14988,N_10303);
xor U18857 (N_18857,N_10323,N_11498);
nand U18858 (N_18858,N_11677,N_11577);
and U18859 (N_18859,N_12650,N_13362);
or U18860 (N_18860,N_12227,N_11115);
xor U18861 (N_18861,N_12091,N_13346);
nor U18862 (N_18862,N_12103,N_12609);
nand U18863 (N_18863,N_12568,N_11082);
and U18864 (N_18864,N_13018,N_12841);
and U18865 (N_18865,N_13681,N_12027);
and U18866 (N_18866,N_13043,N_14012);
or U18867 (N_18867,N_11587,N_14874);
xnor U18868 (N_18868,N_12771,N_12390);
nand U18869 (N_18869,N_11713,N_12525);
nor U18870 (N_18870,N_13390,N_14209);
nand U18871 (N_18871,N_10908,N_11898);
nor U18872 (N_18872,N_14073,N_10381);
xor U18873 (N_18873,N_12794,N_12744);
or U18874 (N_18874,N_10272,N_10183);
xor U18875 (N_18875,N_12874,N_10809);
xnor U18876 (N_18876,N_11407,N_12813);
and U18877 (N_18877,N_13940,N_12989);
nand U18878 (N_18878,N_12255,N_11852);
or U18879 (N_18879,N_13686,N_14243);
nor U18880 (N_18880,N_12951,N_10340);
nor U18881 (N_18881,N_10884,N_10209);
nor U18882 (N_18882,N_13325,N_14450);
xnor U18883 (N_18883,N_13043,N_13651);
nand U18884 (N_18884,N_11487,N_11225);
and U18885 (N_18885,N_12425,N_13180);
xor U18886 (N_18886,N_13413,N_12223);
and U18887 (N_18887,N_13392,N_14113);
and U18888 (N_18888,N_10273,N_10286);
and U18889 (N_18889,N_10766,N_11726);
or U18890 (N_18890,N_11062,N_10137);
and U18891 (N_18891,N_14119,N_11971);
xor U18892 (N_18892,N_10582,N_10881);
nor U18893 (N_18893,N_10652,N_14980);
and U18894 (N_18894,N_10606,N_12518);
or U18895 (N_18895,N_13151,N_10002);
nor U18896 (N_18896,N_12748,N_12827);
and U18897 (N_18897,N_11609,N_13220);
nand U18898 (N_18898,N_12402,N_13661);
and U18899 (N_18899,N_13938,N_12257);
and U18900 (N_18900,N_10707,N_13336);
nor U18901 (N_18901,N_10218,N_13803);
xor U18902 (N_18902,N_12630,N_10177);
xnor U18903 (N_18903,N_10705,N_13068);
xor U18904 (N_18904,N_12596,N_10616);
and U18905 (N_18905,N_13306,N_10950);
nand U18906 (N_18906,N_10367,N_13534);
and U18907 (N_18907,N_10144,N_11311);
or U18908 (N_18908,N_13082,N_12899);
nor U18909 (N_18909,N_13017,N_13073);
xnor U18910 (N_18910,N_12209,N_13164);
and U18911 (N_18911,N_14692,N_11715);
or U18912 (N_18912,N_12759,N_13107);
and U18913 (N_18913,N_12481,N_10685);
nor U18914 (N_18914,N_13505,N_12666);
nand U18915 (N_18915,N_10574,N_14453);
nand U18916 (N_18916,N_11003,N_11464);
and U18917 (N_18917,N_10675,N_14087);
nand U18918 (N_18918,N_12724,N_10308);
or U18919 (N_18919,N_13670,N_13271);
xnor U18920 (N_18920,N_14999,N_12386);
and U18921 (N_18921,N_10541,N_14566);
or U18922 (N_18922,N_12941,N_13772);
and U18923 (N_18923,N_14065,N_10048);
xnor U18924 (N_18924,N_10899,N_10323);
nor U18925 (N_18925,N_10425,N_10695);
nand U18926 (N_18926,N_10035,N_12712);
or U18927 (N_18927,N_14737,N_10123);
and U18928 (N_18928,N_11555,N_14101);
xnor U18929 (N_18929,N_11996,N_12880);
and U18930 (N_18930,N_13172,N_12218);
nand U18931 (N_18931,N_10672,N_11874);
nor U18932 (N_18932,N_13012,N_11059);
or U18933 (N_18933,N_10089,N_13057);
nand U18934 (N_18934,N_14975,N_14838);
nor U18935 (N_18935,N_13223,N_11636);
nand U18936 (N_18936,N_11749,N_11776);
nor U18937 (N_18937,N_14836,N_14670);
xnor U18938 (N_18938,N_10134,N_10903);
xor U18939 (N_18939,N_12925,N_14037);
nor U18940 (N_18940,N_12878,N_13567);
xor U18941 (N_18941,N_11950,N_12153);
nor U18942 (N_18942,N_14003,N_13983);
or U18943 (N_18943,N_11746,N_14631);
or U18944 (N_18944,N_12223,N_11088);
nand U18945 (N_18945,N_14114,N_10078);
nor U18946 (N_18946,N_13532,N_12908);
nor U18947 (N_18947,N_12310,N_12565);
nor U18948 (N_18948,N_12167,N_12271);
xor U18949 (N_18949,N_13650,N_10568);
or U18950 (N_18950,N_12555,N_13175);
xor U18951 (N_18951,N_14488,N_14228);
nor U18952 (N_18952,N_11113,N_10309);
and U18953 (N_18953,N_11894,N_10322);
xnor U18954 (N_18954,N_14645,N_14851);
nor U18955 (N_18955,N_12951,N_12048);
nand U18956 (N_18956,N_14077,N_12686);
or U18957 (N_18957,N_10667,N_11935);
and U18958 (N_18958,N_11113,N_12282);
nand U18959 (N_18959,N_14442,N_11831);
xnor U18960 (N_18960,N_13703,N_11758);
nand U18961 (N_18961,N_10845,N_11249);
or U18962 (N_18962,N_10926,N_11325);
xnor U18963 (N_18963,N_14687,N_14598);
nand U18964 (N_18964,N_12161,N_10716);
xnor U18965 (N_18965,N_10450,N_12938);
nor U18966 (N_18966,N_10166,N_13554);
and U18967 (N_18967,N_14465,N_14810);
nand U18968 (N_18968,N_12164,N_10376);
or U18969 (N_18969,N_10069,N_13324);
and U18970 (N_18970,N_12284,N_13176);
or U18971 (N_18971,N_13357,N_14033);
or U18972 (N_18972,N_13266,N_10642);
or U18973 (N_18973,N_14122,N_12420);
xnor U18974 (N_18974,N_11919,N_14756);
nor U18975 (N_18975,N_14485,N_12922);
nand U18976 (N_18976,N_12331,N_13830);
and U18977 (N_18977,N_11914,N_14252);
xor U18978 (N_18978,N_14417,N_10454);
xor U18979 (N_18979,N_10128,N_14536);
xnor U18980 (N_18980,N_12130,N_10445);
xnor U18981 (N_18981,N_11101,N_12771);
and U18982 (N_18982,N_13097,N_10185);
nand U18983 (N_18983,N_10969,N_12764);
or U18984 (N_18984,N_14739,N_14549);
and U18985 (N_18985,N_12709,N_14729);
or U18986 (N_18986,N_12578,N_14885);
and U18987 (N_18987,N_11116,N_10695);
xor U18988 (N_18988,N_13464,N_12514);
and U18989 (N_18989,N_11807,N_14841);
nand U18990 (N_18990,N_11282,N_14107);
nor U18991 (N_18991,N_14108,N_12503);
nor U18992 (N_18992,N_11675,N_13756);
nor U18993 (N_18993,N_12488,N_13205);
nand U18994 (N_18994,N_14064,N_10668);
or U18995 (N_18995,N_12734,N_10233);
or U18996 (N_18996,N_12713,N_11071);
or U18997 (N_18997,N_14963,N_14948);
xor U18998 (N_18998,N_13292,N_12722);
nor U18999 (N_18999,N_13686,N_11198);
nand U19000 (N_19000,N_13262,N_13937);
nand U19001 (N_19001,N_11774,N_11029);
xnor U19002 (N_19002,N_14520,N_12877);
nor U19003 (N_19003,N_12748,N_13415);
nand U19004 (N_19004,N_12083,N_11916);
nand U19005 (N_19005,N_11439,N_11875);
or U19006 (N_19006,N_13870,N_11572);
nor U19007 (N_19007,N_13250,N_13908);
xnor U19008 (N_19008,N_12525,N_12616);
xor U19009 (N_19009,N_13771,N_13576);
or U19010 (N_19010,N_13928,N_10926);
nand U19011 (N_19011,N_11623,N_14022);
nor U19012 (N_19012,N_11438,N_12326);
nor U19013 (N_19013,N_13303,N_11308);
nand U19014 (N_19014,N_10685,N_13006);
nor U19015 (N_19015,N_11714,N_10526);
nor U19016 (N_19016,N_12028,N_12103);
nand U19017 (N_19017,N_14394,N_10941);
nor U19018 (N_19018,N_14060,N_11747);
nor U19019 (N_19019,N_12228,N_14602);
or U19020 (N_19020,N_12636,N_12590);
or U19021 (N_19021,N_14210,N_10824);
nand U19022 (N_19022,N_12561,N_14468);
nor U19023 (N_19023,N_11032,N_11149);
xnor U19024 (N_19024,N_14346,N_14991);
or U19025 (N_19025,N_10246,N_12105);
xor U19026 (N_19026,N_14245,N_12618);
nor U19027 (N_19027,N_13917,N_13111);
nand U19028 (N_19028,N_11709,N_11542);
nor U19029 (N_19029,N_11079,N_13837);
nor U19030 (N_19030,N_10609,N_12903);
or U19031 (N_19031,N_13916,N_10838);
nand U19032 (N_19032,N_13044,N_10422);
nor U19033 (N_19033,N_10500,N_11978);
or U19034 (N_19034,N_11165,N_12173);
xor U19035 (N_19035,N_12317,N_12012);
or U19036 (N_19036,N_13260,N_11303);
xnor U19037 (N_19037,N_10337,N_14497);
nand U19038 (N_19038,N_10982,N_11765);
and U19039 (N_19039,N_13311,N_14187);
xnor U19040 (N_19040,N_14506,N_12441);
or U19041 (N_19041,N_14106,N_10166);
xor U19042 (N_19042,N_10953,N_10360);
and U19043 (N_19043,N_13971,N_10418);
xnor U19044 (N_19044,N_11596,N_13086);
xnor U19045 (N_19045,N_14834,N_11140);
and U19046 (N_19046,N_10808,N_14175);
nor U19047 (N_19047,N_12282,N_11793);
and U19048 (N_19048,N_14573,N_12287);
or U19049 (N_19049,N_11473,N_14026);
nor U19050 (N_19050,N_11529,N_13526);
nand U19051 (N_19051,N_10748,N_12701);
and U19052 (N_19052,N_13934,N_14920);
nand U19053 (N_19053,N_13909,N_13771);
nand U19054 (N_19054,N_13710,N_13434);
or U19055 (N_19055,N_11310,N_11829);
or U19056 (N_19056,N_13505,N_13559);
nor U19057 (N_19057,N_13480,N_11989);
or U19058 (N_19058,N_13651,N_11861);
nor U19059 (N_19059,N_10344,N_13009);
nand U19060 (N_19060,N_13278,N_14407);
and U19061 (N_19061,N_13807,N_14004);
and U19062 (N_19062,N_13390,N_10042);
nand U19063 (N_19063,N_12100,N_10925);
and U19064 (N_19064,N_12803,N_13800);
or U19065 (N_19065,N_12823,N_12521);
nand U19066 (N_19066,N_10456,N_12289);
or U19067 (N_19067,N_12358,N_10301);
or U19068 (N_19068,N_10695,N_10696);
nor U19069 (N_19069,N_12292,N_11247);
or U19070 (N_19070,N_12320,N_12803);
or U19071 (N_19071,N_12811,N_11988);
nand U19072 (N_19072,N_11470,N_10444);
xnor U19073 (N_19073,N_14533,N_12957);
nor U19074 (N_19074,N_11524,N_10141);
or U19075 (N_19075,N_11968,N_10135);
nor U19076 (N_19076,N_14653,N_11797);
or U19077 (N_19077,N_11904,N_14050);
xnor U19078 (N_19078,N_11838,N_10126);
or U19079 (N_19079,N_12830,N_11743);
nand U19080 (N_19080,N_12937,N_12961);
nand U19081 (N_19081,N_10800,N_10403);
nand U19082 (N_19082,N_10392,N_11804);
nor U19083 (N_19083,N_14798,N_13158);
and U19084 (N_19084,N_11796,N_11329);
nor U19085 (N_19085,N_13630,N_13373);
xnor U19086 (N_19086,N_14853,N_11119);
and U19087 (N_19087,N_10291,N_14370);
or U19088 (N_19088,N_10530,N_10548);
and U19089 (N_19089,N_11960,N_14532);
xnor U19090 (N_19090,N_10111,N_14291);
nand U19091 (N_19091,N_13816,N_14613);
nand U19092 (N_19092,N_11644,N_14056);
xor U19093 (N_19093,N_12963,N_10093);
or U19094 (N_19094,N_10383,N_11003);
nand U19095 (N_19095,N_14008,N_14104);
and U19096 (N_19096,N_13456,N_10181);
or U19097 (N_19097,N_14722,N_12397);
nor U19098 (N_19098,N_11018,N_12064);
and U19099 (N_19099,N_14863,N_12659);
xor U19100 (N_19100,N_11602,N_10919);
nand U19101 (N_19101,N_12921,N_12320);
nor U19102 (N_19102,N_14294,N_14932);
nor U19103 (N_19103,N_10151,N_10237);
or U19104 (N_19104,N_11509,N_12976);
xor U19105 (N_19105,N_12522,N_10341);
or U19106 (N_19106,N_14571,N_11897);
nand U19107 (N_19107,N_14854,N_12057);
and U19108 (N_19108,N_10457,N_11323);
or U19109 (N_19109,N_12620,N_13582);
xnor U19110 (N_19110,N_11747,N_13206);
or U19111 (N_19111,N_11516,N_13174);
and U19112 (N_19112,N_13769,N_13811);
and U19113 (N_19113,N_13760,N_13838);
nor U19114 (N_19114,N_11967,N_11118);
nand U19115 (N_19115,N_11273,N_12405);
nand U19116 (N_19116,N_13055,N_10104);
nor U19117 (N_19117,N_11789,N_14673);
xor U19118 (N_19118,N_10552,N_11594);
nor U19119 (N_19119,N_11598,N_13812);
nand U19120 (N_19120,N_11249,N_14371);
nand U19121 (N_19121,N_12966,N_14684);
and U19122 (N_19122,N_14285,N_12508);
and U19123 (N_19123,N_12826,N_14656);
nand U19124 (N_19124,N_13713,N_14413);
or U19125 (N_19125,N_13307,N_10046);
and U19126 (N_19126,N_10239,N_13453);
or U19127 (N_19127,N_12274,N_10274);
xor U19128 (N_19128,N_12674,N_11767);
nor U19129 (N_19129,N_14540,N_14877);
xnor U19130 (N_19130,N_14391,N_14871);
nor U19131 (N_19131,N_11277,N_12235);
nor U19132 (N_19132,N_10147,N_13671);
nor U19133 (N_19133,N_13760,N_14871);
nor U19134 (N_19134,N_12950,N_13317);
xor U19135 (N_19135,N_13742,N_14611);
xor U19136 (N_19136,N_13788,N_13262);
nor U19137 (N_19137,N_13073,N_12400);
and U19138 (N_19138,N_12096,N_13419);
nor U19139 (N_19139,N_13204,N_11830);
nor U19140 (N_19140,N_10614,N_14632);
and U19141 (N_19141,N_10314,N_10433);
nor U19142 (N_19142,N_10408,N_11247);
xor U19143 (N_19143,N_11923,N_14708);
or U19144 (N_19144,N_14701,N_10688);
or U19145 (N_19145,N_13846,N_13478);
nand U19146 (N_19146,N_14522,N_14021);
and U19147 (N_19147,N_13772,N_13065);
or U19148 (N_19148,N_10348,N_10182);
nand U19149 (N_19149,N_14372,N_11648);
xnor U19150 (N_19150,N_10040,N_13207);
and U19151 (N_19151,N_10932,N_10819);
xor U19152 (N_19152,N_12649,N_12544);
nor U19153 (N_19153,N_12429,N_12816);
nand U19154 (N_19154,N_13733,N_11205);
xor U19155 (N_19155,N_13725,N_11399);
or U19156 (N_19156,N_10695,N_14767);
xnor U19157 (N_19157,N_14844,N_12824);
xor U19158 (N_19158,N_11244,N_13731);
and U19159 (N_19159,N_13759,N_11956);
nand U19160 (N_19160,N_11545,N_10182);
xnor U19161 (N_19161,N_10010,N_12817);
nor U19162 (N_19162,N_13891,N_14357);
nor U19163 (N_19163,N_10940,N_14070);
or U19164 (N_19164,N_12144,N_12693);
or U19165 (N_19165,N_11779,N_13400);
and U19166 (N_19166,N_10052,N_13181);
nand U19167 (N_19167,N_11598,N_10386);
and U19168 (N_19168,N_11670,N_14088);
nand U19169 (N_19169,N_13017,N_14363);
xor U19170 (N_19170,N_11494,N_11039);
nor U19171 (N_19171,N_13209,N_14597);
or U19172 (N_19172,N_13447,N_14901);
and U19173 (N_19173,N_14499,N_14813);
xor U19174 (N_19174,N_13066,N_13394);
nand U19175 (N_19175,N_12759,N_14186);
and U19176 (N_19176,N_11078,N_14007);
xnor U19177 (N_19177,N_10744,N_14575);
nand U19178 (N_19178,N_11572,N_12562);
nand U19179 (N_19179,N_10447,N_12652);
or U19180 (N_19180,N_11579,N_12019);
or U19181 (N_19181,N_11548,N_13583);
and U19182 (N_19182,N_12696,N_14390);
nand U19183 (N_19183,N_14590,N_14684);
nand U19184 (N_19184,N_11465,N_13628);
and U19185 (N_19185,N_10910,N_14931);
or U19186 (N_19186,N_10506,N_12770);
or U19187 (N_19187,N_14542,N_13745);
and U19188 (N_19188,N_10345,N_11463);
nor U19189 (N_19189,N_14417,N_13800);
nand U19190 (N_19190,N_10960,N_10812);
xnor U19191 (N_19191,N_11059,N_12546);
or U19192 (N_19192,N_14595,N_13601);
nor U19193 (N_19193,N_11335,N_10275);
or U19194 (N_19194,N_12599,N_11011);
xnor U19195 (N_19195,N_14210,N_11808);
and U19196 (N_19196,N_11892,N_11835);
or U19197 (N_19197,N_13304,N_14890);
or U19198 (N_19198,N_14428,N_10326);
nor U19199 (N_19199,N_11264,N_12591);
xnor U19200 (N_19200,N_12813,N_12584);
nand U19201 (N_19201,N_14068,N_11213);
xnor U19202 (N_19202,N_12426,N_10834);
nand U19203 (N_19203,N_12156,N_14410);
nand U19204 (N_19204,N_11629,N_11420);
and U19205 (N_19205,N_10998,N_12038);
nor U19206 (N_19206,N_12262,N_13706);
nor U19207 (N_19207,N_11493,N_12373);
nor U19208 (N_19208,N_10069,N_14649);
or U19209 (N_19209,N_14879,N_10372);
nand U19210 (N_19210,N_13358,N_10586);
nor U19211 (N_19211,N_13219,N_12428);
nand U19212 (N_19212,N_13626,N_12802);
nand U19213 (N_19213,N_13365,N_13248);
nand U19214 (N_19214,N_10414,N_12503);
and U19215 (N_19215,N_14639,N_13892);
or U19216 (N_19216,N_13541,N_12184);
or U19217 (N_19217,N_13421,N_11440);
nor U19218 (N_19218,N_13675,N_13824);
or U19219 (N_19219,N_12136,N_12308);
nor U19220 (N_19220,N_13936,N_12649);
nand U19221 (N_19221,N_14723,N_14677);
and U19222 (N_19222,N_11684,N_14738);
or U19223 (N_19223,N_13524,N_12991);
and U19224 (N_19224,N_12400,N_12719);
nand U19225 (N_19225,N_11356,N_11019);
or U19226 (N_19226,N_14821,N_12100);
or U19227 (N_19227,N_11070,N_13155);
nand U19228 (N_19228,N_10733,N_12763);
xnor U19229 (N_19229,N_12986,N_13569);
nor U19230 (N_19230,N_14455,N_13694);
or U19231 (N_19231,N_14894,N_13342);
and U19232 (N_19232,N_11436,N_10973);
xnor U19233 (N_19233,N_14840,N_14994);
nor U19234 (N_19234,N_12857,N_11864);
nand U19235 (N_19235,N_13467,N_11878);
xnor U19236 (N_19236,N_10204,N_13522);
nor U19237 (N_19237,N_12868,N_11829);
or U19238 (N_19238,N_12971,N_10728);
nand U19239 (N_19239,N_12064,N_12285);
nor U19240 (N_19240,N_13482,N_12566);
and U19241 (N_19241,N_13366,N_14026);
nor U19242 (N_19242,N_11095,N_11535);
nand U19243 (N_19243,N_13606,N_11152);
and U19244 (N_19244,N_13153,N_10991);
xor U19245 (N_19245,N_13908,N_10397);
or U19246 (N_19246,N_14168,N_13656);
xnor U19247 (N_19247,N_13709,N_13806);
nand U19248 (N_19248,N_10482,N_10897);
nor U19249 (N_19249,N_14832,N_14983);
or U19250 (N_19250,N_10147,N_13875);
and U19251 (N_19251,N_14819,N_14784);
nand U19252 (N_19252,N_13256,N_11460);
xor U19253 (N_19253,N_10290,N_12447);
xnor U19254 (N_19254,N_14536,N_11451);
and U19255 (N_19255,N_10675,N_10354);
and U19256 (N_19256,N_13576,N_11875);
nor U19257 (N_19257,N_12587,N_12990);
or U19258 (N_19258,N_14915,N_14682);
or U19259 (N_19259,N_10202,N_11412);
or U19260 (N_19260,N_12811,N_13457);
xnor U19261 (N_19261,N_12612,N_10317);
nor U19262 (N_19262,N_12372,N_13394);
or U19263 (N_19263,N_12959,N_14877);
xnor U19264 (N_19264,N_10057,N_11475);
or U19265 (N_19265,N_11526,N_10785);
and U19266 (N_19266,N_14265,N_10525);
nand U19267 (N_19267,N_12992,N_10874);
nand U19268 (N_19268,N_13390,N_13058);
and U19269 (N_19269,N_12309,N_14502);
nand U19270 (N_19270,N_12806,N_11230);
or U19271 (N_19271,N_13194,N_10133);
nor U19272 (N_19272,N_11085,N_14471);
nand U19273 (N_19273,N_10931,N_11739);
nand U19274 (N_19274,N_13144,N_14248);
nor U19275 (N_19275,N_10755,N_14081);
or U19276 (N_19276,N_11015,N_14574);
nor U19277 (N_19277,N_14407,N_11285);
nand U19278 (N_19278,N_13624,N_11141);
or U19279 (N_19279,N_10085,N_14359);
nand U19280 (N_19280,N_13742,N_11993);
or U19281 (N_19281,N_12696,N_11560);
or U19282 (N_19282,N_14465,N_12560);
nand U19283 (N_19283,N_14992,N_13830);
nand U19284 (N_19284,N_10260,N_12495);
nand U19285 (N_19285,N_14214,N_13450);
and U19286 (N_19286,N_10132,N_14655);
nor U19287 (N_19287,N_12702,N_14644);
nor U19288 (N_19288,N_12187,N_14623);
nor U19289 (N_19289,N_14766,N_10142);
nor U19290 (N_19290,N_11694,N_10674);
or U19291 (N_19291,N_10829,N_12070);
or U19292 (N_19292,N_11178,N_13284);
nor U19293 (N_19293,N_13719,N_12191);
nor U19294 (N_19294,N_12542,N_13582);
and U19295 (N_19295,N_10478,N_13838);
nand U19296 (N_19296,N_10302,N_14541);
or U19297 (N_19297,N_13286,N_11307);
or U19298 (N_19298,N_10609,N_11056);
xor U19299 (N_19299,N_11562,N_13954);
xor U19300 (N_19300,N_12809,N_11751);
xnor U19301 (N_19301,N_13239,N_10643);
xnor U19302 (N_19302,N_11708,N_14577);
nand U19303 (N_19303,N_10472,N_10207);
nor U19304 (N_19304,N_10650,N_14596);
and U19305 (N_19305,N_13889,N_12908);
nor U19306 (N_19306,N_10231,N_13840);
nand U19307 (N_19307,N_12382,N_13251);
nor U19308 (N_19308,N_13273,N_10083);
or U19309 (N_19309,N_14299,N_14998);
xor U19310 (N_19310,N_10357,N_12008);
nor U19311 (N_19311,N_11491,N_13099);
xnor U19312 (N_19312,N_12265,N_10509);
nand U19313 (N_19313,N_11919,N_14029);
nor U19314 (N_19314,N_10295,N_12841);
or U19315 (N_19315,N_12726,N_13274);
or U19316 (N_19316,N_10903,N_10207);
or U19317 (N_19317,N_11364,N_14620);
nand U19318 (N_19318,N_14097,N_11218);
nand U19319 (N_19319,N_14926,N_14742);
and U19320 (N_19320,N_11359,N_14276);
nor U19321 (N_19321,N_11146,N_14715);
and U19322 (N_19322,N_11036,N_11581);
nand U19323 (N_19323,N_12422,N_12541);
and U19324 (N_19324,N_11146,N_12908);
or U19325 (N_19325,N_12392,N_11146);
xor U19326 (N_19326,N_10985,N_12850);
xnor U19327 (N_19327,N_14366,N_10413);
nand U19328 (N_19328,N_12487,N_11677);
and U19329 (N_19329,N_13093,N_11002);
xnor U19330 (N_19330,N_13712,N_12385);
and U19331 (N_19331,N_10136,N_14481);
nor U19332 (N_19332,N_12964,N_11039);
and U19333 (N_19333,N_11779,N_14361);
nand U19334 (N_19334,N_13034,N_11142);
nand U19335 (N_19335,N_13447,N_11277);
nor U19336 (N_19336,N_11606,N_14706);
or U19337 (N_19337,N_12544,N_13876);
nor U19338 (N_19338,N_12401,N_12932);
xnor U19339 (N_19339,N_13162,N_10386);
nor U19340 (N_19340,N_10579,N_11340);
xor U19341 (N_19341,N_14175,N_10847);
xnor U19342 (N_19342,N_14808,N_14585);
or U19343 (N_19343,N_13789,N_11183);
xor U19344 (N_19344,N_13858,N_13976);
xnor U19345 (N_19345,N_14080,N_11892);
and U19346 (N_19346,N_11010,N_10168);
and U19347 (N_19347,N_12131,N_13487);
nor U19348 (N_19348,N_12310,N_13420);
nor U19349 (N_19349,N_11436,N_14658);
or U19350 (N_19350,N_13946,N_12253);
and U19351 (N_19351,N_10661,N_14848);
or U19352 (N_19352,N_13796,N_11800);
nor U19353 (N_19353,N_13877,N_14036);
xnor U19354 (N_19354,N_13256,N_10849);
nand U19355 (N_19355,N_10992,N_10401);
nor U19356 (N_19356,N_12677,N_12859);
and U19357 (N_19357,N_11861,N_13563);
nor U19358 (N_19358,N_13391,N_11426);
or U19359 (N_19359,N_13576,N_14183);
nor U19360 (N_19360,N_14646,N_14685);
xnor U19361 (N_19361,N_14581,N_14265);
nand U19362 (N_19362,N_13926,N_10647);
nor U19363 (N_19363,N_12444,N_12184);
or U19364 (N_19364,N_13491,N_13542);
nand U19365 (N_19365,N_14811,N_10312);
nor U19366 (N_19366,N_10475,N_13717);
xnor U19367 (N_19367,N_11010,N_13438);
nand U19368 (N_19368,N_10402,N_12900);
nor U19369 (N_19369,N_12582,N_10135);
and U19370 (N_19370,N_10556,N_11203);
and U19371 (N_19371,N_14776,N_12503);
and U19372 (N_19372,N_10533,N_14252);
nor U19373 (N_19373,N_13137,N_10790);
and U19374 (N_19374,N_12150,N_13927);
xnor U19375 (N_19375,N_13951,N_11331);
xnor U19376 (N_19376,N_13314,N_12485);
xor U19377 (N_19377,N_10776,N_14001);
and U19378 (N_19378,N_10955,N_11442);
nand U19379 (N_19379,N_10778,N_13820);
and U19380 (N_19380,N_14662,N_12565);
and U19381 (N_19381,N_14521,N_10209);
nand U19382 (N_19382,N_11771,N_13244);
nand U19383 (N_19383,N_14494,N_13479);
nand U19384 (N_19384,N_13387,N_11786);
and U19385 (N_19385,N_11854,N_13484);
or U19386 (N_19386,N_13889,N_12836);
nor U19387 (N_19387,N_12276,N_10128);
or U19388 (N_19388,N_14617,N_12841);
or U19389 (N_19389,N_12533,N_14934);
xor U19390 (N_19390,N_11796,N_11080);
and U19391 (N_19391,N_14461,N_10950);
xor U19392 (N_19392,N_13311,N_13853);
nand U19393 (N_19393,N_11057,N_14404);
or U19394 (N_19394,N_11669,N_10701);
and U19395 (N_19395,N_11382,N_13391);
xor U19396 (N_19396,N_12115,N_12765);
nor U19397 (N_19397,N_14275,N_10576);
nand U19398 (N_19398,N_13746,N_13041);
nand U19399 (N_19399,N_12600,N_11021);
xor U19400 (N_19400,N_14704,N_13201);
and U19401 (N_19401,N_13379,N_12331);
or U19402 (N_19402,N_10712,N_14714);
or U19403 (N_19403,N_14518,N_12846);
xnor U19404 (N_19404,N_12038,N_12813);
or U19405 (N_19405,N_13914,N_14911);
nand U19406 (N_19406,N_13917,N_10165);
xor U19407 (N_19407,N_13943,N_13893);
nand U19408 (N_19408,N_13565,N_14106);
or U19409 (N_19409,N_11574,N_11707);
xnor U19410 (N_19410,N_13410,N_10027);
nor U19411 (N_19411,N_14312,N_11452);
xnor U19412 (N_19412,N_12539,N_12300);
nor U19413 (N_19413,N_14533,N_10948);
nor U19414 (N_19414,N_10913,N_12109);
and U19415 (N_19415,N_12490,N_14755);
and U19416 (N_19416,N_11983,N_10314);
or U19417 (N_19417,N_13852,N_10428);
nand U19418 (N_19418,N_11199,N_11734);
and U19419 (N_19419,N_12320,N_14249);
or U19420 (N_19420,N_11350,N_12982);
and U19421 (N_19421,N_14116,N_13153);
and U19422 (N_19422,N_10367,N_12547);
xor U19423 (N_19423,N_10764,N_13668);
xnor U19424 (N_19424,N_11349,N_10696);
and U19425 (N_19425,N_10908,N_12021);
or U19426 (N_19426,N_14287,N_13504);
xnor U19427 (N_19427,N_12846,N_11782);
nor U19428 (N_19428,N_13398,N_14189);
and U19429 (N_19429,N_10510,N_10689);
and U19430 (N_19430,N_12720,N_11522);
nor U19431 (N_19431,N_11356,N_11046);
nand U19432 (N_19432,N_11027,N_10905);
nor U19433 (N_19433,N_12413,N_14942);
nor U19434 (N_19434,N_10684,N_12517);
nor U19435 (N_19435,N_13692,N_12840);
xor U19436 (N_19436,N_13346,N_13986);
nand U19437 (N_19437,N_11832,N_12627);
nor U19438 (N_19438,N_14565,N_10401);
and U19439 (N_19439,N_13673,N_14110);
nand U19440 (N_19440,N_14112,N_10238);
and U19441 (N_19441,N_13730,N_12485);
nand U19442 (N_19442,N_12764,N_14471);
and U19443 (N_19443,N_10857,N_11905);
or U19444 (N_19444,N_11415,N_10051);
nor U19445 (N_19445,N_12591,N_12079);
or U19446 (N_19446,N_12877,N_10343);
and U19447 (N_19447,N_13730,N_12046);
nand U19448 (N_19448,N_12092,N_10277);
or U19449 (N_19449,N_13707,N_14804);
nand U19450 (N_19450,N_10408,N_14932);
nand U19451 (N_19451,N_13212,N_14143);
xor U19452 (N_19452,N_12361,N_11564);
and U19453 (N_19453,N_14886,N_12263);
nor U19454 (N_19454,N_14170,N_10468);
and U19455 (N_19455,N_13656,N_14350);
and U19456 (N_19456,N_11786,N_14487);
or U19457 (N_19457,N_11164,N_11628);
xor U19458 (N_19458,N_13980,N_14724);
nor U19459 (N_19459,N_11032,N_12773);
nand U19460 (N_19460,N_12657,N_10809);
and U19461 (N_19461,N_13260,N_14835);
xnor U19462 (N_19462,N_10843,N_10009);
xor U19463 (N_19463,N_12866,N_12307);
or U19464 (N_19464,N_12295,N_12165);
xnor U19465 (N_19465,N_12767,N_14596);
nand U19466 (N_19466,N_12090,N_12441);
or U19467 (N_19467,N_10290,N_10559);
nand U19468 (N_19468,N_13491,N_13363);
and U19469 (N_19469,N_13404,N_14061);
nand U19470 (N_19470,N_13836,N_13586);
and U19471 (N_19471,N_10889,N_14203);
and U19472 (N_19472,N_12442,N_13650);
and U19473 (N_19473,N_14344,N_10375);
nor U19474 (N_19474,N_12038,N_14544);
nor U19475 (N_19475,N_13035,N_10182);
nor U19476 (N_19476,N_11340,N_13974);
xnor U19477 (N_19477,N_11848,N_11752);
xor U19478 (N_19478,N_14289,N_13793);
nand U19479 (N_19479,N_12718,N_11072);
nor U19480 (N_19480,N_10337,N_10054);
nor U19481 (N_19481,N_13469,N_13863);
nor U19482 (N_19482,N_10166,N_10880);
nor U19483 (N_19483,N_10302,N_10666);
nor U19484 (N_19484,N_11377,N_10116);
nor U19485 (N_19485,N_14611,N_10308);
xor U19486 (N_19486,N_10281,N_12799);
nor U19487 (N_19487,N_14592,N_11114);
and U19488 (N_19488,N_11377,N_11931);
or U19489 (N_19489,N_14715,N_11661);
nor U19490 (N_19490,N_14035,N_14727);
and U19491 (N_19491,N_11412,N_12256);
nand U19492 (N_19492,N_14890,N_12944);
or U19493 (N_19493,N_13551,N_13570);
nand U19494 (N_19494,N_10371,N_11393);
or U19495 (N_19495,N_11055,N_12492);
xnor U19496 (N_19496,N_10728,N_13467);
nand U19497 (N_19497,N_13291,N_11872);
xor U19498 (N_19498,N_10462,N_10340);
nor U19499 (N_19499,N_13878,N_13225);
xnor U19500 (N_19500,N_10933,N_13521);
nor U19501 (N_19501,N_10474,N_10771);
xnor U19502 (N_19502,N_13013,N_14999);
xor U19503 (N_19503,N_11993,N_12759);
and U19504 (N_19504,N_13073,N_12798);
and U19505 (N_19505,N_14521,N_13101);
nand U19506 (N_19506,N_11543,N_12477);
or U19507 (N_19507,N_10733,N_11493);
or U19508 (N_19508,N_11193,N_13747);
and U19509 (N_19509,N_13909,N_11702);
nand U19510 (N_19510,N_11716,N_13030);
xor U19511 (N_19511,N_11766,N_10677);
nor U19512 (N_19512,N_14987,N_11330);
nand U19513 (N_19513,N_14329,N_14056);
and U19514 (N_19514,N_13569,N_13297);
or U19515 (N_19515,N_14383,N_14431);
or U19516 (N_19516,N_10908,N_12258);
nor U19517 (N_19517,N_11435,N_14961);
nand U19518 (N_19518,N_11824,N_10412);
and U19519 (N_19519,N_11256,N_10846);
or U19520 (N_19520,N_11632,N_10556);
xnor U19521 (N_19521,N_13153,N_11700);
and U19522 (N_19522,N_14431,N_10357);
xor U19523 (N_19523,N_13495,N_14130);
and U19524 (N_19524,N_11178,N_11611);
or U19525 (N_19525,N_14606,N_12908);
nand U19526 (N_19526,N_14815,N_11149);
nand U19527 (N_19527,N_10141,N_12777);
xnor U19528 (N_19528,N_12544,N_11021);
nand U19529 (N_19529,N_10913,N_13091);
nand U19530 (N_19530,N_11390,N_11580);
nor U19531 (N_19531,N_12573,N_12814);
and U19532 (N_19532,N_11366,N_13365);
and U19533 (N_19533,N_12439,N_13946);
and U19534 (N_19534,N_12457,N_13410);
or U19535 (N_19535,N_12941,N_13927);
xnor U19536 (N_19536,N_13690,N_11742);
nor U19537 (N_19537,N_11814,N_12985);
nand U19538 (N_19538,N_12056,N_11354);
nand U19539 (N_19539,N_10990,N_11539);
xor U19540 (N_19540,N_14380,N_11287);
xnor U19541 (N_19541,N_10014,N_11643);
nand U19542 (N_19542,N_14612,N_10983);
or U19543 (N_19543,N_14402,N_14299);
or U19544 (N_19544,N_13269,N_11363);
or U19545 (N_19545,N_13914,N_14219);
xnor U19546 (N_19546,N_10996,N_14227);
and U19547 (N_19547,N_11818,N_10236);
nor U19548 (N_19548,N_11551,N_13514);
nor U19549 (N_19549,N_10202,N_12169);
or U19550 (N_19550,N_13908,N_14685);
nand U19551 (N_19551,N_11708,N_14369);
and U19552 (N_19552,N_11793,N_13176);
or U19553 (N_19553,N_13871,N_12844);
nand U19554 (N_19554,N_13426,N_12280);
and U19555 (N_19555,N_13093,N_10657);
nor U19556 (N_19556,N_10949,N_10858);
xor U19557 (N_19557,N_14434,N_11244);
nand U19558 (N_19558,N_13608,N_13529);
and U19559 (N_19559,N_11592,N_10377);
nand U19560 (N_19560,N_11021,N_14834);
nand U19561 (N_19561,N_10147,N_14498);
nand U19562 (N_19562,N_10299,N_10932);
or U19563 (N_19563,N_14001,N_12887);
and U19564 (N_19564,N_13972,N_12963);
and U19565 (N_19565,N_11807,N_14468);
or U19566 (N_19566,N_11126,N_14131);
nand U19567 (N_19567,N_10406,N_13268);
nor U19568 (N_19568,N_11312,N_14402);
xnor U19569 (N_19569,N_11599,N_14283);
nor U19570 (N_19570,N_11834,N_10525);
or U19571 (N_19571,N_13018,N_10711);
xor U19572 (N_19572,N_12870,N_12943);
nand U19573 (N_19573,N_13658,N_12318);
or U19574 (N_19574,N_11304,N_13941);
and U19575 (N_19575,N_10633,N_14241);
and U19576 (N_19576,N_14547,N_13511);
xnor U19577 (N_19577,N_13292,N_14251);
xor U19578 (N_19578,N_12002,N_11417);
xnor U19579 (N_19579,N_14565,N_10932);
or U19580 (N_19580,N_10089,N_11486);
nor U19581 (N_19581,N_12937,N_13756);
and U19582 (N_19582,N_12032,N_12533);
nand U19583 (N_19583,N_10448,N_10197);
nand U19584 (N_19584,N_14310,N_14663);
xnor U19585 (N_19585,N_14912,N_14972);
or U19586 (N_19586,N_13699,N_11508);
nand U19587 (N_19587,N_13108,N_13484);
and U19588 (N_19588,N_13172,N_14264);
nor U19589 (N_19589,N_12789,N_10928);
nand U19590 (N_19590,N_12773,N_12659);
or U19591 (N_19591,N_11124,N_10319);
nand U19592 (N_19592,N_10940,N_13088);
nor U19593 (N_19593,N_14761,N_14525);
and U19594 (N_19594,N_14254,N_11928);
nand U19595 (N_19595,N_11359,N_13832);
xor U19596 (N_19596,N_13318,N_12637);
and U19597 (N_19597,N_14017,N_13990);
or U19598 (N_19598,N_10915,N_14778);
and U19599 (N_19599,N_10359,N_10635);
or U19600 (N_19600,N_10388,N_11342);
nor U19601 (N_19601,N_11536,N_12631);
nor U19602 (N_19602,N_10882,N_14669);
nor U19603 (N_19603,N_13242,N_12783);
xor U19604 (N_19604,N_12735,N_13230);
and U19605 (N_19605,N_14978,N_13978);
xnor U19606 (N_19606,N_14791,N_10484);
nor U19607 (N_19607,N_14845,N_14729);
nor U19608 (N_19608,N_11035,N_13783);
xnor U19609 (N_19609,N_13441,N_10841);
xnor U19610 (N_19610,N_10503,N_13343);
xnor U19611 (N_19611,N_12300,N_13768);
and U19612 (N_19612,N_10097,N_12207);
or U19613 (N_19613,N_13505,N_14053);
nand U19614 (N_19614,N_10004,N_10668);
nand U19615 (N_19615,N_10172,N_12777);
nor U19616 (N_19616,N_11335,N_12470);
nor U19617 (N_19617,N_10840,N_10565);
or U19618 (N_19618,N_10610,N_11302);
nor U19619 (N_19619,N_14332,N_12280);
xor U19620 (N_19620,N_10221,N_13560);
or U19621 (N_19621,N_12529,N_12815);
xnor U19622 (N_19622,N_13119,N_11097);
or U19623 (N_19623,N_12729,N_12191);
nor U19624 (N_19624,N_13015,N_13553);
nand U19625 (N_19625,N_13744,N_13333);
nor U19626 (N_19626,N_14677,N_14150);
and U19627 (N_19627,N_10722,N_14344);
nor U19628 (N_19628,N_12222,N_10518);
xor U19629 (N_19629,N_12848,N_10412);
nor U19630 (N_19630,N_12154,N_10589);
nand U19631 (N_19631,N_13060,N_12808);
and U19632 (N_19632,N_11802,N_14352);
xor U19633 (N_19633,N_10288,N_12500);
nand U19634 (N_19634,N_10130,N_10393);
nor U19635 (N_19635,N_12204,N_11366);
or U19636 (N_19636,N_12778,N_11063);
xor U19637 (N_19637,N_12758,N_13802);
nand U19638 (N_19638,N_14662,N_11344);
nand U19639 (N_19639,N_12416,N_10087);
nor U19640 (N_19640,N_12690,N_14839);
or U19641 (N_19641,N_12545,N_12806);
xor U19642 (N_19642,N_13921,N_14523);
nor U19643 (N_19643,N_13226,N_12916);
nand U19644 (N_19644,N_13270,N_14729);
nand U19645 (N_19645,N_13298,N_13796);
xnor U19646 (N_19646,N_13327,N_10531);
nand U19647 (N_19647,N_10757,N_13883);
or U19648 (N_19648,N_14417,N_10781);
and U19649 (N_19649,N_11065,N_14274);
or U19650 (N_19650,N_12214,N_14692);
nor U19651 (N_19651,N_14489,N_12573);
nand U19652 (N_19652,N_12729,N_10685);
nand U19653 (N_19653,N_14525,N_13150);
nand U19654 (N_19654,N_10293,N_14583);
nand U19655 (N_19655,N_13812,N_14745);
and U19656 (N_19656,N_10423,N_14517);
nor U19657 (N_19657,N_12226,N_12102);
or U19658 (N_19658,N_11028,N_13873);
or U19659 (N_19659,N_11316,N_14583);
nor U19660 (N_19660,N_13966,N_14716);
nor U19661 (N_19661,N_12393,N_12226);
or U19662 (N_19662,N_11721,N_10942);
and U19663 (N_19663,N_14571,N_11327);
xnor U19664 (N_19664,N_13597,N_13008);
or U19665 (N_19665,N_13378,N_11880);
nand U19666 (N_19666,N_10068,N_14250);
and U19667 (N_19667,N_10812,N_11754);
or U19668 (N_19668,N_12566,N_10410);
nor U19669 (N_19669,N_11351,N_13478);
and U19670 (N_19670,N_10617,N_11349);
and U19671 (N_19671,N_11350,N_10437);
or U19672 (N_19672,N_11727,N_13989);
nand U19673 (N_19673,N_12069,N_13355);
nand U19674 (N_19674,N_13289,N_14659);
nand U19675 (N_19675,N_10543,N_11140);
xor U19676 (N_19676,N_12407,N_12748);
and U19677 (N_19677,N_11986,N_11848);
nand U19678 (N_19678,N_12773,N_11415);
and U19679 (N_19679,N_12823,N_11414);
nor U19680 (N_19680,N_14395,N_11428);
and U19681 (N_19681,N_10520,N_13784);
and U19682 (N_19682,N_10489,N_14703);
xor U19683 (N_19683,N_12247,N_10586);
nand U19684 (N_19684,N_13332,N_14149);
and U19685 (N_19685,N_11799,N_14032);
xnor U19686 (N_19686,N_14369,N_11712);
nand U19687 (N_19687,N_11317,N_10001);
or U19688 (N_19688,N_12263,N_14385);
or U19689 (N_19689,N_10138,N_11860);
and U19690 (N_19690,N_10184,N_10572);
nor U19691 (N_19691,N_14601,N_14856);
nand U19692 (N_19692,N_13218,N_12515);
nor U19693 (N_19693,N_12205,N_11889);
nor U19694 (N_19694,N_14644,N_14932);
xor U19695 (N_19695,N_14090,N_11699);
nand U19696 (N_19696,N_13898,N_13446);
and U19697 (N_19697,N_14029,N_11499);
or U19698 (N_19698,N_12052,N_14070);
nand U19699 (N_19699,N_13727,N_14790);
nor U19700 (N_19700,N_13741,N_13583);
or U19701 (N_19701,N_13298,N_13688);
xnor U19702 (N_19702,N_12976,N_13234);
xnor U19703 (N_19703,N_13819,N_11396);
and U19704 (N_19704,N_13616,N_13050);
nand U19705 (N_19705,N_11327,N_12082);
nand U19706 (N_19706,N_13677,N_10535);
nand U19707 (N_19707,N_12568,N_13631);
and U19708 (N_19708,N_12553,N_14413);
xor U19709 (N_19709,N_11886,N_12782);
nand U19710 (N_19710,N_12310,N_13925);
and U19711 (N_19711,N_11879,N_10023);
nor U19712 (N_19712,N_10830,N_13585);
and U19713 (N_19713,N_10997,N_12425);
and U19714 (N_19714,N_14448,N_10873);
or U19715 (N_19715,N_14596,N_13746);
nor U19716 (N_19716,N_11525,N_11963);
or U19717 (N_19717,N_13574,N_11586);
nand U19718 (N_19718,N_11197,N_12870);
nor U19719 (N_19719,N_11391,N_10130);
nand U19720 (N_19720,N_10274,N_12355);
nor U19721 (N_19721,N_10737,N_10588);
xor U19722 (N_19722,N_11906,N_13814);
nand U19723 (N_19723,N_14144,N_12021);
nand U19724 (N_19724,N_10802,N_14919);
or U19725 (N_19725,N_13601,N_12006);
or U19726 (N_19726,N_13970,N_14228);
and U19727 (N_19727,N_12058,N_10149);
and U19728 (N_19728,N_10350,N_14202);
and U19729 (N_19729,N_12032,N_14020);
nand U19730 (N_19730,N_13522,N_11175);
nor U19731 (N_19731,N_12053,N_13112);
nand U19732 (N_19732,N_12885,N_12704);
and U19733 (N_19733,N_11794,N_14104);
and U19734 (N_19734,N_14688,N_11784);
and U19735 (N_19735,N_11453,N_13044);
and U19736 (N_19736,N_12748,N_14184);
or U19737 (N_19737,N_10162,N_14721);
nor U19738 (N_19738,N_12398,N_12470);
xor U19739 (N_19739,N_14847,N_12353);
nor U19740 (N_19740,N_12890,N_14929);
and U19741 (N_19741,N_10131,N_14163);
or U19742 (N_19742,N_12218,N_14651);
nand U19743 (N_19743,N_11086,N_13584);
and U19744 (N_19744,N_13959,N_11569);
nand U19745 (N_19745,N_10730,N_13344);
nor U19746 (N_19746,N_12381,N_12300);
and U19747 (N_19747,N_11279,N_13708);
nor U19748 (N_19748,N_10836,N_13868);
or U19749 (N_19749,N_10380,N_11096);
nand U19750 (N_19750,N_13784,N_10759);
nor U19751 (N_19751,N_11514,N_12515);
nor U19752 (N_19752,N_13806,N_11917);
nand U19753 (N_19753,N_13102,N_11820);
nor U19754 (N_19754,N_13554,N_13762);
nor U19755 (N_19755,N_14682,N_10308);
nor U19756 (N_19756,N_13636,N_11309);
nor U19757 (N_19757,N_13450,N_13414);
xor U19758 (N_19758,N_12002,N_12568);
xor U19759 (N_19759,N_10057,N_12100);
nor U19760 (N_19760,N_11862,N_13012);
xnor U19761 (N_19761,N_10621,N_12339);
xor U19762 (N_19762,N_14264,N_10198);
or U19763 (N_19763,N_13156,N_14696);
or U19764 (N_19764,N_11628,N_11943);
and U19765 (N_19765,N_10475,N_11435);
or U19766 (N_19766,N_13183,N_10853);
nor U19767 (N_19767,N_11696,N_12759);
and U19768 (N_19768,N_11309,N_12522);
xnor U19769 (N_19769,N_12793,N_14536);
or U19770 (N_19770,N_13621,N_11075);
nor U19771 (N_19771,N_10525,N_13287);
nand U19772 (N_19772,N_11527,N_10129);
or U19773 (N_19773,N_13579,N_12596);
and U19774 (N_19774,N_14703,N_13170);
nand U19775 (N_19775,N_11794,N_10464);
and U19776 (N_19776,N_13718,N_14034);
xnor U19777 (N_19777,N_13811,N_12893);
xnor U19778 (N_19778,N_13538,N_10765);
xnor U19779 (N_19779,N_14977,N_14672);
and U19780 (N_19780,N_13043,N_12186);
xnor U19781 (N_19781,N_13962,N_12307);
nor U19782 (N_19782,N_10477,N_12425);
and U19783 (N_19783,N_14001,N_14800);
xor U19784 (N_19784,N_10807,N_14793);
or U19785 (N_19785,N_13271,N_10424);
nand U19786 (N_19786,N_11375,N_12453);
xnor U19787 (N_19787,N_12768,N_11216);
xnor U19788 (N_19788,N_14720,N_14820);
nor U19789 (N_19789,N_14372,N_13632);
nor U19790 (N_19790,N_11258,N_14835);
nand U19791 (N_19791,N_13179,N_14725);
and U19792 (N_19792,N_12706,N_10139);
nand U19793 (N_19793,N_12044,N_14891);
nand U19794 (N_19794,N_12350,N_10314);
or U19795 (N_19795,N_12155,N_10641);
and U19796 (N_19796,N_14256,N_14603);
or U19797 (N_19797,N_14043,N_14073);
nand U19798 (N_19798,N_14656,N_10539);
nor U19799 (N_19799,N_11925,N_13816);
xor U19800 (N_19800,N_10023,N_13507);
and U19801 (N_19801,N_12788,N_11142);
or U19802 (N_19802,N_11237,N_12779);
or U19803 (N_19803,N_13259,N_12171);
nor U19804 (N_19804,N_14787,N_11872);
and U19805 (N_19805,N_12891,N_13226);
nand U19806 (N_19806,N_14037,N_13701);
and U19807 (N_19807,N_10119,N_14785);
and U19808 (N_19808,N_11720,N_12095);
or U19809 (N_19809,N_14616,N_13839);
or U19810 (N_19810,N_11494,N_10876);
nand U19811 (N_19811,N_11818,N_12747);
nor U19812 (N_19812,N_10579,N_13740);
xor U19813 (N_19813,N_11354,N_14600);
or U19814 (N_19814,N_10401,N_14395);
and U19815 (N_19815,N_11302,N_10001);
nand U19816 (N_19816,N_12070,N_11066);
xor U19817 (N_19817,N_13345,N_14011);
and U19818 (N_19818,N_11921,N_12234);
xnor U19819 (N_19819,N_10953,N_11924);
nand U19820 (N_19820,N_11922,N_11296);
nor U19821 (N_19821,N_13945,N_10544);
or U19822 (N_19822,N_13687,N_10392);
and U19823 (N_19823,N_10345,N_13721);
xnor U19824 (N_19824,N_11565,N_11266);
and U19825 (N_19825,N_10889,N_14886);
xnor U19826 (N_19826,N_11786,N_11501);
nor U19827 (N_19827,N_12361,N_11441);
nand U19828 (N_19828,N_14536,N_11722);
xor U19829 (N_19829,N_11722,N_10086);
nor U19830 (N_19830,N_10391,N_13424);
and U19831 (N_19831,N_14671,N_10079);
or U19832 (N_19832,N_11526,N_13784);
nor U19833 (N_19833,N_11015,N_11442);
or U19834 (N_19834,N_11771,N_10542);
nor U19835 (N_19835,N_10540,N_11018);
nor U19836 (N_19836,N_14040,N_11393);
and U19837 (N_19837,N_10884,N_13398);
and U19838 (N_19838,N_13618,N_14415);
nor U19839 (N_19839,N_12974,N_14106);
or U19840 (N_19840,N_13948,N_12192);
nand U19841 (N_19841,N_12307,N_10321);
xor U19842 (N_19842,N_10199,N_13931);
xor U19843 (N_19843,N_13135,N_12046);
or U19844 (N_19844,N_14454,N_11174);
xor U19845 (N_19845,N_12813,N_10931);
nand U19846 (N_19846,N_13529,N_10084);
nor U19847 (N_19847,N_14077,N_10770);
nor U19848 (N_19848,N_10204,N_10793);
or U19849 (N_19849,N_10105,N_10324);
nand U19850 (N_19850,N_12171,N_10283);
or U19851 (N_19851,N_14029,N_11103);
nand U19852 (N_19852,N_10679,N_12984);
or U19853 (N_19853,N_11450,N_11981);
nor U19854 (N_19854,N_12207,N_12157);
xor U19855 (N_19855,N_14724,N_11727);
or U19856 (N_19856,N_14053,N_10241);
nor U19857 (N_19857,N_11801,N_14922);
nor U19858 (N_19858,N_10850,N_14930);
nand U19859 (N_19859,N_12835,N_13390);
nor U19860 (N_19860,N_13159,N_14732);
or U19861 (N_19861,N_11343,N_10488);
nand U19862 (N_19862,N_13361,N_14656);
xnor U19863 (N_19863,N_13737,N_12002);
xnor U19864 (N_19864,N_14277,N_10419);
xnor U19865 (N_19865,N_13390,N_14284);
or U19866 (N_19866,N_13969,N_12874);
and U19867 (N_19867,N_12163,N_12603);
nand U19868 (N_19868,N_10722,N_13144);
and U19869 (N_19869,N_11343,N_10494);
xnor U19870 (N_19870,N_13667,N_13683);
and U19871 (N_19871,N_14331,N_12943);
xor U19872 (N_19872,N_11789,N_12812);
nand U19873 (N_19873,N_12697,N_12792);
and U19874 (N_19874,N_11139,N_12263);
or U19875 (N_19875,N_11657,N_10883);
xnor U19876 (N_19876,N_14857,N_12267);
nor U19877 (N_19877,N_14034,N_11973);
or U19878 (N_19878,N_14645,N_13905);
xnor U19879 (N_19879,N_12865,N_12303);
nor U19880 (N_19880,N_14680,N_12078);
nor U19881 (N_19881,N_13026,N_11288);
xnor U19882 (N_19882,N_10748,N_10474);
and U19883 (N_19883,N_11029,N_12783);
nor U19884 (N_19884,N_10227,N_11613);
or U19885 (N_19885,N_12385,N_10777);
nand U19886 (N_19886,N_12249,N_14683);
and U19887 (N_19887,N_14872,N_14791);
nand U19888 (N_19888,N_12620,N_11669);
or U19889 (N_19889,N_10283,N_14959);
xor U19890 (N_19890,N_14101,N_12615);
and U19891 (N_19891,N_10550,N_12295);
or U19892 (N_19892,N_10644,N_10204);
nor U19893 (N_19893,N_14285,N_11759);
nor U19894 (N_19894,N_12278,N_11632);
or U19895 (N_19895,N_14840,N_14303);
nand U19896 (N_19896,N_14798,N_10484);
and U19897 (N_19897,N_14305,N_14845);
nand U19898 (N_19898,N_14936,N_11145);
nor U19899 (N_19899,N_12128,N_14172);
or U19900 (N_19900,N_12120,N_14772);
nand U19901 (N_19901,N_10782,N_11660);
and U19902 (N_19902,N_12655,N_14041);
and U19903 (N_19903,N_13890,N_10203);
xor U19904 (N_19904,N_14319,N_13150);
and U19905 (N_19905,N_13694,N_13558);
xnor U19906 (N_19906,N_14652,N_14219);
and U19907 (N_19907,N_10856,N_11758);
nor U19908 (N_19908,N_13591,N_13239);
nor U19909 (N_19909,N_12569,N_13045);
xor U19910 (N_19910,N_12836,N_14533);
or U19911 (N_19911,N_10245,N_13608);
or U19912 (N_19912,N_12222,N_13289);
xor U19913 (N_19913,N_12540,N_11084);
nor U19914 (N_19914,N_11028,N_13384);
nor U19915 (N_19915,N_12748,N_13911);
or U19916 (N_19916,N_13798,N_14441);
nand U19917 (N_19917,N_10404,N_13136);
or U19918 (N_19918,N_10055,N_14902);
or U19919 (N_19919,N_14484,N_12442);
nor U19920 (N_19920,N_12146,N_11251);
nand U19921 (N_19921,N_11773,N_14885);
and U19922 (N_19922,N_13249,N_13514);
nand U19923 (N_19923,N_13875,N_10768);
or U19924 (N_19924,N_12880,N_12506);
and U19925 (N_19925,N_14701,N_14680);
and U19926 (N_19926,N_13634,N_12864);
nand U19927 (N_19927,N_14060,N_11667);
xor U19928 (N_19928,N_14963,N_11903);
nor U19929 (N_19929,N_12366,N_11553);
nand U19930 (N_19930,N_10238,N_12797);
nor U19931 (N_19931,N_11269,N_11735);
nand U19932 (N_19932,N_14271,N_11371);
or U19933 (N_19933,N_13238,N_10783);
xor U19934 (N_19934,N_13412,N_11974);
nand U19935 (N_19935,N_11018,N_13918);
nand U19936 (N_19936,N_10214,N_14831);
or U19937 (N_19937,N_11557,N_13060);
xor U19938 (N_19938,N_14377,N_13271);
xor U19939 (N_19939,N_11508,N_10264);
and U19940 (N_19940,N_14079,N_10764);
or U19941 (N_19941,N_13364,N_13330);
nand U19942 (N_19942,N_14124,N_13899);
and U19943 (N_19943,N_12508,N_11165);
and U19944 (N_19944,N_12487,N_12628);
and U19945 (N_19945,N_12357,N_12094);
nand U19946 (N_19946,N_10550,N_12743);
and U19947 (N_19947,N_12580,N_13709);
or U19948 (N_19948,N_11459,N_14066);
and U19949 (N_19949,N_14715,N_12106);
or U19950 (N_19950,N_14224,N_11473);
xnor U19951 (N_19951,N_14047,N_14322);
xnor U19952 (N_19952,N_14488,N_11017);
or U19953 (N_19953,N_14987,N_12054);
nand U19954 (N_19954,N_12509,N_12885);
nand U19955 (N_19955,N_12786,N_10755);
nor U19956 (N_19956,N_11024,N_12012);
nor U19957 (N_19957,N_10461,N_11013);
and U19958 (N_19958,N_13983,N_13114);
and U19959 (N_19959,N_10602,N_13943);
nand U19960 (N_19960,N_11349,N_13170);
xor U19961 (N_19961,N_13949,N_13587);
and U19962 (N_19962,N_13500,N_14123);
nand U19963 (N_19963,N_10066,N_11243);
nand U19964 (N_19964,N_11729,N_10279);
nand U19965 (N_19965,N_10704,N_12902);
xnor U19966 (N_19966,N_10503,N_13538);
xor U19967 (N_19967,N_12996,N_12938);
nor U19968 (N_19968,N_11795,N_10807);
and U19969 (N_19969,N_13292,N_11644);
and U19970 (N_19970,N_14901,N_13862);
nor U19971 (N_19971,N_13253,N_11174);
or U19972 (N_19972,N_13836,N_10830);
and U19973 (N_19973,N_13873,N_10201);
nor U19974 (N_19974,N_11675,N_10065);
or U19975 (N_19975,N_12855,N_10996);
nor U19976 (N_19976,N_11125,N_12029);
nand U19977 (N_19977,N_12481,N_11681);
or U19978 (N_19978,N_10893,N_13993);
nand U19979 (N_19979,N_10717,N_10249);
nor U19980 (N_19980,N_10750,N_10150);
xor U19981 (N_19981,N_14333,N_14059);
nor U19982 (N_19982,N_14754,N_11204);
nor U19983 (N_19983,N_10507,N_13405);
and U19984 (N_19984,N_13714,N_14372);
and U19985 (N_19985,N_12034,N_10705);
nand U19986 (N_19986,N_13121,N_12631);
nor U19987 (N_19987,N_12505,N_10393);
and U19988 (N_19988,N_10785,N_14351);
nand U19989 (N_19989,N_10415,N_12635);
and U19990 (N_19990,N_13546,N_10687);
or U19991 (N_19991,N_10189,N_10267);
and U19992 (N_19992,N_11596,N_11113);
or U19993 (N_19993,N_12374,N_12773);
nor U19994 (N_19994,N_10866,N_10539);
or U19995 (N_19995,N_14498,N_13121);
or U19996 (N_19996,N_12511,N_13448);
nor U19997 (N_19997,N_14175,N_11278);
nor U19998 (N_19998,N_10568,N_10907);
or U19999 (N_19999,N_12165,N_14236);
nor U20000 (N_20000,N_19428,N_19722);
nor U20001 (N_20001,N_17468,N_15027);
and U20002 (N_20002,N_19088,N_18272);
nor U20003 (N_20003,N_19574,N_18828);
and U20004 (N_20004,N_19946,N_19342);
nor U20005 (N_20005,N_19228,N_15322);
xor U20006 (N_20006,N_15776,N_15760);
nand U20007 (N_20007,N_19886,N_15733);
and U20008 (N_20008,N_19346,N_15608);
xor U20009 (N_20009,N_15338,N_15844);
and U20010 (N_20010,N_17899,N_19027);
nand U20011 (N_20011,N_15549,N_18624);
nand U20012 (N_20012,N_18056,N_16787);
nand U20013 (N_20013,N_18012,N_15892);
and U20014 (N_20014,N_16043,N_18436);
xor U20015 (N_20015,N_17135,N_18871);
nor U20016 (N_20016,N_16335,N_17259);
xor U20017 (N_20017,N_18152,N_17124);
nand U20018 (N_20018,N_15618,N_16398);
nand U20019 (N_20019,N_15901,N_17798);
nor U20020 (N_20020,N_15152,N_17353);
xor U20021 (N_20021,N_18791,N_17216);
nand U20022 (N_20022,N_18475,N_16637);
nor U20023 (N_20023,N_19581,N_15367);
or U20024 (N_20024,N_16524,N_18002);
nor U20025 (N_20025,N_17619,N_15454);
nand U20026 (N_20026,N_16230,N_15688);
or U20027 (N_20027,N_15574,N_15645);
or U20028 (N_20028,N_16924,N_19188);
xnor U20029 (N_20029,N_17527,N_17816);
and U20030 (N_20030,N_18036,N_19204);
nor U20031 (N_20031,N_18688,N_18532);
or U20032 (N_20032,N_19130,N_17033);
or U20033 (N_20033,N_16520,N_19795);
xnor U20034 (N_20034,N_17334,N_18627);
xor U20035 (N_20035,N_17976,N_15221);
nand U20036 (N_20036,N_16134,N_18288);
nor U20037 (N_20037,N_18111,N_17207);
nand U20038 (N_20038,N_18852,N_15088);
nor U20039 (N_20039,N_19250,N_16047);
and U20040 (N_20040,N_19236,N_19736);
nor U20041 (N_20041,N_18394,N_18356);
xor U20042 (N_20042,N_18809,N_19281);
xnor U20043 (N_20043,N_18812,N_18737);
and U20044 (N_20044,N_19080,N_17595);
and U20045 (N_20045,N_16965,N_19288);
or U20046 (N_20046,N_18529,N_17993);
xor U20047 (N_20047,N_16336,N_18541);
nand U20048 (N_20048,N_16364,N_15311);
nor U20049 (N_20049,N_17673,N_16585);
xnor U20050 (N_20050,N_16625,N_19006);
nor U20051 (N_20051,N_18962,N_17845);
nor U20052 (N_20052,N_19920,N_18198);
or U20053 (N_20053,N_16807,N_17854);
and U20054 (N_20054,N_15658,N_18298);
xor U20055 (N_20055,N_16857,N_16062);
xor U20056 (N_20056,N_18146,N_15796);
nor U20057 (N_20057,N_18526,N_16796);
nand U20058 (N_20058,N_15328,N_16988);
nor U20059 (N_20059,N_18017,N_16837);
nand U20060 (N_20060,N_17743,N_15672);
or U20061 (N_20061,N_16792,N_19845);
nor U20062 (N_20062,N_19796,N_15607);
and U20063 (N_20063,N_15537,N_15290);
xnor U20064 (N_20064,N_19153,N_19049);
xnor U20065 (N_20065,N_15067,N_15742);
or U20066 (N_20066,N_17592,N_16859);
xnor U20067 (N_20067,N_16953,N_19679);
xnor U20068 (N_20068,N_18981,N_17591);
or U20069 (N_20069,N_19460,N_16028);
nor U20070 (N_20070,N_18866,N_16962);
nand U20071 (N_20071,N_17907,N_19077);
nand U20072 (N_20072,N_16041,N_15186);
or U20073 (N_20073,N_19136,N_15546);
and U20074 (N_20074,N_18634,N_17515);
xor U20075 (N_20075,N_18292,N_16082);
and U20076 (N_20076,N_15223,N_17451);
and U20077 (N_20077,N_19430,N_18456);
nand U20078 (N_20078,N_16921,N_16730);
xor U20079 (N_20079,N_19494,N_15061);
xor U20080 (N_20080,N_18788,N_18760);
and U20081 (N_20081,N_15967,N_17972);
nand U20082 (N_20082,N_18531,N_18948);
or U20083 (N_20083,N_18903,N_15771);
xnor U20084 (N_20084,N_17099,N_18655);
and U20085 (N_20085,N_18051,N_15205);
and U20086 (N_20086,N_16052,N_15199);
xnor U20087 (N_20087,N_19249,N_16534);
xnor U20088 (N_20088,N_18187,N_17089);
or U20089 (N_20089,N_17088,N_18346);
xor U20090 (N_20090,N_16665,N_19023);
or U20091 (N_20091,N_18675,N_18970);
or U20092 (N_20092,N_17540,N_17837);
nand U20093 (N_20093,N_17891,N_15578);
nand U20094 (N_20094,N_19200,N_16133);
nand U20095 (N_20095,N_19354,N_16964);
nor U20096 (N_20096,N_16367,N_19894);
nand U20097 (N_20097,N_17681,N_16247);
or U20098 (N_20098,N_17262,N_19776);
nor U20099 (N_20099,N_16113,N_18899);
xor U20100 (N_20100,N_19386,N_17424);
xor U20101 (N_20101,N_16250,N_17118);
and U20102 (N_20102,N_17544,N_16155);
nand U20103 (N_20103,N_15123,N_16543);
or U20104 (N_20104,N_16803,N_16118);
or U20105 (N_20105,N_17714,N_16768);
nor U20106 (N_20106,N_17422,N_15845);
and U20107 (N_20107,N_17943,N_15218);
nor U20108 (N_20108,N_18207,N_19631);
nor U20109 (N_20109,N_18229,N_17096);
nor U20110 (N_20110,N_15837,N_18328);
and U20111 (N_20111,N_19507,N_19579);
nand U20112 (N_20112,N_19693,N_18433);
and U20113 (N_20113,N_15450,N_17774);
or U20114 (N_20114,N_19757,N_19569);
xor U20115 (N_20115,N_18022,N_19968);
or U20116 (N_20116,N_18885,N_15079);
and U20117 (N_20117,N_18195,N_16242);
and U20118 (N_20118,N_19559,N_18727);
xor U20119 (N_20119,N_18883,N_16575);
nand U20120 (N_20120,N_16437,N_19211);
nor U20121 (N_20121,N_18633,N_19554);
nor U20122 (N_20122,N_18900,N_17065);
or U20123 (N_20123,N_16183,N_18957);
xnor U20124 (N_20124,N_17287,N_19930);
nand U20125 (N_20125,N_15793,N_19252);
or U20126 (N_20126,N_17375,N_19667);
xor U20127 (N_20127,N_15619,N_18635);
and U20128 (N_20128,N_19974,N_17805);
nor U20129 (N_20129,N_18336,N_16209);
nand U20130 (N_20130,N_16349,N_18877);
nand U20131 (N_20131,N_17370,N_19867);
nor U20132 (N_20132,N_15911,N_15504);
and U20133 (N_20133,N_16533,N_15728);
xor U20134 (N_20134,N_17178,N_18088);
xor U20135 (N_20135,N_17426,N_19329);
and U20136 (N_20136,N_16614,N_19912);
or U20137 (N_20137,N_18845,N_19786);
nor U20138 (N_20138,N_15518,N_18466);
nor U20139 (N_20139,N_18372,N_17935);
xnor U20140 (N_20140,N_15600,N_18654);
or U20141 (N_20141,N_19371,N_18452);
and U20142 (N_20142,N_19962,N_19126);
or U20143 (N_20143,N_16726,N_15001);
or U20144 (N_20144,N_15550,N_16698);
nand U20145 (N_20145,N_15075,N_17877);
nor U20146 (N_20146,N_17824,N_17603);
nor U20147 (N_20147,N_17889,N_15990);
nor U20148 (N_20148,N_16817,N_15082);
nor U20149 (N_20149,N_15120,N_16111);
nand U20150 (N_20150,N_16345,N_18125);
nor U20151 (N_20151,N_17499,N_17423);
or U20152 (N_20152,N_16695,N_19135);
or U20153 (N_20153,N_17026,N_15099);
nand U20154 (N_20154,N_17647,N_17825);
nand U20155 (N_20155,N_17330,N_17699);
or U20156 (N_20156,N_15192,N_15856);
xnor U20157 (N_20157,N_15236,N_19885);
nor U20158 (N_20158,N_16539,N_19519);
and U20159 (N_20159,N_15973,N_15206);
and U20160 (N_20160,N_16213,N_15446);
nand U20161 (N_20161,N_15468,N_16805);
or U20162 (N_20162,N_17038,N_15375);
xnor U20163 (N_20163,N_15102,N_15269);
or U20164 (N_20164,N_17839,N_18869);
or U20165 (N_20165,N_17497,N_16691);
nand U20166 (N_20166,N_17585,N_16499);
nor U20167 (N_20167,N_16622,N_19546);
and U20168 (N_20168,N_17432,N_16329);
nand U20169 (N_20169,N_19378,N_19239);
or U20170 (N_20170,N_16794,N_17460);
xnor U20171 (N_20171,N_15568,N_17878);
and U20172 (N_20172,N_16968,N_18909);
nand U20173 (N_20173,N_19840,N_19452);
nand U20174 (N_20174,N_17183,N_16724);
and U20175 (N_20175,N_19585,N_17611);
nor U20176 (N_20176,N_19924,N_19043);
nor U20177 (N_20177,N_18060,N_16684);
or U20178 (N_20178,N_17550,N_18431);
nand U20179 (N_20179,N_15731,N_16451);
and U20180 (N_20180,N_19688,N_19549);
xor U20181 (N_20181,N_17730,N_16806);
and U20182 (N_20182,N_19122,N_16468);
or U20183 (N_20183,N_17163,N_17503);
xnor U20184 (N_20184,N_15430,N_17498);
nand U20185 (N_20185,N_16220,N_17618);
nand U20186 (N_20186,N_15178,N_18488);
nor U20187 (N_20187,N_18177,N_18956);
or U20188 (N_20188,N_16982,N_16136);
nand U20189 (N_20189,N_19727,N_15409);
and U20190 (N_20190,N_15467,N_18745);
or U20191 (N_20191,N_18273,N_15745);
nor U20192 (N_20192,N_15381,N_19531);
nand U20193 (N_20193,N_17741,N_15126);
nand U20194 (N_20194,N_16606,N_18813);
nand U20195 (N_20195,N_15165,N_19480);
xor U20196 (N_20196,N_19651,N_15867);
nand U20197 (N_20197,N_17322,N_17105);
or U20198 (N_20198,N_19540,N_19595);
nor U20199 (N_20199,N_15840,N_19301);
xnor U20200 (N_20200,N_16702,N_19289);
and U20201 (N_20201,N_19109,N_15809);
or U20202 (N_20202,N_15954,N_15599);
xor U20203 (N_20203,N_18639,N_18427);
nor U20204 (N_20204,N_17631,N_16010);
nor U20205 (N_20205,N_15458,N_18483);
nand U20206 (N_20206,N_17159,N_16605);
and U20207 (N_20207,N_15853,N_18241);
xor U20208 (N_20208,N_15457,N_19223);
nor U20209 (N_20209,N_19745,N_19768);
xor U20210 (N_20210,N_17395,N_17505);
nor U20211 (N_20211,N_17523,N_17855);
or U20212 (N_20212,N_17478,N_19317);
nand U20213 (N_20213,N_15652,N_16458);
and U20214 (N_20214,N_17997,N_15233);
nor U20215 (N_20215,N_17371,N_18110);
and U20216 (N_20216,N_16497,N_15893);
nand U20217 (N_20217,N_15969,N_17329);
or U20218 (N_20218,N_19983,N_17867);
or U20219 (N_20219,N_19599,N_17806);
xnor U20220 (N_20220,N_15267,N_19202);
and U20221 (N_20221,N_18700,N_19992);
or U20222 (N_20222,N_17193,N_19299);
or U20223 (N_20223,N_19509,N_16054);
nand U20224 (N_20224,N_15749,N_18902);
xor U20225 (N_20225,N_19809,N_15052);
nand U20226 (N_20226,N_19053,N_15250);
or U20227 (N_20227,N_17320,N_17394);
or U20228 (N_20228,N_18611,N_19298);
and U20229 (N_20229,N_15654,N_19799);
nand U20230 (N_20230,N_15820,N_15665);
and U20231 (N_20231,N_17533,N_18095);
xnor U20232 (N_20232,N_18335,N_18106);
nor U20233 (N_20233,N_15810,N_17823);
and U20234 (N_20234,N_18920,N_15396);
nor U20235 (N_20235,N_15303,N_17166);
nand U20236 (N_20236,N_17056,N_15506);
and U20237 (N_20237,N_16419,N_17693);
xor U20238 (N_20238,N_16288,N_15648);
nor U20239 (N_20239,N_18143,N_15740);
nand U20240 (N_20240,N_19037,N_16132);
and U20241 (N_20241,N_18257,N_16971);
or U20242 (N_20242,N_15297,N_19062);
xnor U20243 (N_20243,N_18856,N_19705);
or U20244 (N_20244,N_17581,N_17017);
nor U20245 (N_20245,N_17474,N_16512);
and U20246 (N_20246,N_18600,N_17787);
nand U20247 (N_20247,N_15646,N_15923);
and U20248 (N_20248,N_19785,N_16408);
and U20249 (N_20249,N_16391,N_16005);
nor U20250 (N_20250,N_19898,N_19957);
nor U20251 (N_20251,N_15565,N_18862);
nand U20252 (N_20252,N_15933,N_16931);
xnor U20253 (N_20253,N_18572,N_15542);
and U20254 (N_20254,N_16973,N_17010);
and U20255 (N_20255,N_19133,N_18952);
nor U20256 (N_20256,N_17793,N_18720);
nand U20257 (N_20257,N_15916,N_16620);
nor U20258 (N_20258,N_18113,N_19143);
xnor U20259 (N_20259,N_16358,N_19831);
nand U20260 (N_20260,N_15175,N_17187);
xor U20261 (N_20261,N_16018,N_17189);
nor U20262 (N_20262,N_19721,N_17727);
nor U20263 (N_20263,N_19230,N_18797);
and U20264 (N_20264,N_17378,N_18690);
and U20265 (N_20265,N_19580,N_16293);
nor U20266 (N_20266,N_16441,N_17936);
and U20267 (N_20267,N_17555,N_17362);
or U20268 (N_20268,N_15639,N_18398);
nand U20269 (N_20269,N_17804,N_17399);
or U20270 (N_20270,N_19773,N_17345);
xor U20271 (N_20271,N_15805,N_17041);
nor U20272 (N_20272,N_15530,N_19150);
nand U20273 (N_20273,N_18965,N_19673);
xnor U20274 (N_20274,N_18592,N_17062);
and U20275 (N_20275,N_18940,N_17649);
nand U20276 (N_20276,N_15072,N_15818);
nand U20277 (N_20277,N_15266,N_19610);
and U20278 (N_20278,N_15156,N_15469);
nand U20279 (N_20279,N_18971,N_15693);
or U20280 (N_20280,N_19873,N_19843);
xor U20281 (N_20281,N_16906,N_15314);
and U20282 (N_20282,N_17779,N_19600);
or U20283 (N_20283,N_15699,N_18988);
nand U20284 (N_20284,N_17130,N_18549);
or U20285 (N_20285,N_19694,N_18694);
xnor U20286 (N_20286,N_15014,N_15750);
or U20287 (N_20287,N_18937,N_18975);
and U20288 (N_20288,N_18689,N_15927);
nor U20289 (N_20289,N_15276,N_17875);
nand U20290 (N_20290,N_16330,N_17098);
or U20291 (N_20291,N_19454,N_15891);
nand U20292 (N_20292,N_17682,N_19921);
xnor U20293 (N_20293,N_18656,N_18983);
and U20294 (N_20294,N_19641,N_16501);
and U20295 (N_20295,N_17713,N_17167);
or U20296 (N_20296,N_15062,N_16646);
xnor U20297 (N_20297,N_17171,N_19351);
and U20298 (N_20298,N_16619,N_15497);
xnor U20299 (N_20299,N_19309,N_19189);
nor U20300 (N_20300,N_19167,N_15637);
and U20301 (N_20301,N_16845,N_15134);
nand U20302 (N_20302,N_18776,N_19429);
and U20303 (N_20303,N_18015,N_17408);
nor U20304 (N_20304,N_15517,N_16117);
xor U20305 (N_20305,N_15798,N_17236);
xnor U20306 (N_20306,N_19238,N_17176);
nand U20307 (N_20307,N_15945,N_16483);
nand U20308 (N_20308,N_19565,N_18625);
nand U20309 (N_20309,N_17464,N_15885);
nor U20310 (N_20310,N_18384,N_16003);
xor U20311 (N_20311,N_18616,N_17517);
nand U20312 (N_20312,N_16643,N_19560);
nor U20313 (N_20313,N_18217,N_19008);
or U20314 (N_20314,N_18942,N_15115);
nand U20315 (N_20315,N_17536,N_19817);
nand U20316 (N_20316,N_18594,N_15025);
or U20317 (N_20317,N_19304,N_16092);
nor U20318 (N_20318,N_16399,N_17414);
or U20319 (N_20319,N_17608,N_15439);
and U20320 (N_20320,N_18360,N_19159);
nor U20321 (N_20321,N_18395,N_17597);
and U20322 (N_20322,N_18705,N_17077);
nor U20323 (N_20323,N_18619,N_17994);
xnor U20324 (N_20324,N_18787,N_19089);
xnor U20325 (N_20325,N_17104,N_15044);
nand U20326 (N_20326,N_17092,N_17147);
xor U20327 (N_20327,N_18057,N_19407);
or U20328 (N_20328,N_19515,N_16566);
nand U20329 (N_20329,N_17679,N_16356);
nand U20330 (N_20330,N_15757,N_15685);
or U20331 (N_20331,N_16257,N_16269);
xnor U20332 (N_20332,N_15295,N_16189);
nor U20333 (N_20333,N_16940,N_18240);
or U20334 (N_20334,N_16311,N_19608);
nand U20335 (N_20335,N_17838,N_15159);
and U20336 (N_20336,N_15959,N_17304);
or U20337 (N_20337,N_18204,N_16781);
nand U20338 (N_20338,N_15936,N_19657);
nor U20339 (N_20339,N_16736,N_15752);
and U20340 (N_20340,N_15071,N_17925);
nor U20341 (N_20341,N_17296,N_18978);
nor U20342 (N_20342,N_18556,N_15437);
xnor U20343 (N_20343,N_19634,N_15717);
xnor U20344 (N_20344,N_17924,N_15584);
or U20345 (N_20345,N_19320,N_18873);
and U20346 (N_20346,N_19165,N_15009);
or U20347 (N_20347,N_15922,N_15739);
nand U20348 (N_20348,N_19087,N_17857);
and U20349 (N_20349,N_15065,N_17518);
nand U20350 (N_20350,N_15859,N_15874);
nand U20351 (N_20351,N_15358,N_18476);
nor U20352 (N_20352,N_19573,N_15794);
or U20353 (N_20353,N_18922,N_19423);
or U20354 (N_20354,N_18440,N_16418);
nand U20355 (N_20355,N_18622,N_15698);
nand U20356 (N_20356,N_15906,N_15208);
or U20357 (N_20357,N_17613,N_15664);
or U20358 (N_20358,N_19233,N_17847);
nor U20359 (N_20359,N_17734,N_19503);
nor U20360 (N_20360,N_18679,N_19710);
xnor U20361 (N_20361,N_15272,N_19083);
nor U20362 (N_20362,N_19308,N_15692);
and U20363 (N_20363,N_15816,N_18910);
xor U20364 (N_20364,N_19348,N_16528);
or U20365 (N_20365,N_15164,N_19125);
nand U20366 (N_20366,N_18411,N_15133);
nand U20367 (N_20367,N_15012,N_16178);
nand U20368 (N_20368,N_17705,N_19010);
xnor U20369 (N_20369,N_17381,N_18738);
or U20370 (N_20370,N_15668,N_16978);
xnor U20371 (N_20371,N_19652,N_16711);
or U20372 (N_20372,N_18709,N_17722);
nand U20373 (N_20373,N_15228,N_17247);
or U20374 (N_20374,N_17390,N_15800);
and U20375 (N_20375,N_17316,N_18505);
nor U20376 (N_20376,N_15815,N_15320);
nand U20377 (N_20377,N_16650,N_15201);
and U20378 (N_20378,N_15781,N_18716);
nor U20379 (N_20379,N_17846,N_18141);
and U20380 (N_20380,N_15335,N_18001);
nand U20381 (N_20381,N_15103,N_17488);
xor U20382 (N_20382,N_18671,N_15020);
and U20383 (N_20383,N_16179,N_15419);
or U20384 (N_20384,N_15138,N_18210);
and U20385 (N_20385,N_15759,N_16686);
nand U20386 (N_20386,N_17622,N_16211);
nor U20387 (N_20387,N_16375,N_19092);
xor U20388 (N_20388,N_16927,N_18465);
xnor U20389 (N_20389,N_17970,N_17563);
xnor U20390 (N_20390,N_18363,N_16970);
xor U20391 (N_20391,N_15593,N_17690);
nand U20392 (N_20392,N_15538,N_15577);
or U20393 (N_20393,N_15556,N_19905);
or U20394 (N_20394,N_17851,N_18517);
nor U20395 (N_20395,N_16067,N_18365);
nor U20396 (N_20396,N_15579,N_16416);
or U20397 (N_20397,N_18918,N_17756);
and U20398 (N_20398,N_18087,N_15963);
nor U20399 (N_20399,N_17582,N_18853);
or U20400 (N_20400,N_19743,N_17716);
xnor U20401 (N_20401,N_15161,N_16139);
nor U20402 (N_20402,N_15718,N_18994);
nor U20403 (N_20403,N_19616,N_18042);
nor U20404 (N_20404,N_17910,N_17361);
xnor U20405 (N_20405,N_16779,N_19523);
and U20406 (N_20406,N_17580,N_17016);
nand U20407 (N_20407,N_15562,N_16581);
nand U20408 (N_20408,N_15147,N_16945);
nand U20409 (N_20409,N_15225,N_17763);
nand U20410 (N_20410,N_15128,N_19808);
and U20411 (N_20411,N_18596,N_16120);
nor U20412 (N_20412,N_19235,N_19504);
or U20413 (N_20413,N_19622,N_18340);
or U20414 (N_20414,N_16904,N_18601);
xor U20415 (N_20415,N_18354,N_18371);
or U20416 (N_20416,N_19483,N_17045);
nor U20417 (N_20417,N_16180,N_18147);
xnor U20418 (N_20418,N_16503,N_17626);
and U20419 (N_20419,N_16216,N_17433);
or U20420 (N_20420,N_17548,N_18729);
xnor U20421 (N_20421,N_17428,N_18551);
and U20422 (N_20422,N_19478,N_16261);
nand U20423 (N_20423,N_15489,N_19810);
and U20424 (N_20424,N_17977,N_15241);
or U20425 (N_20425,N_18021,N_18339);
and U20426 (N_20426,N_16798,N_18358);
or U20427 (N_20427,N_19267,N_15195);
and U20428 (N_20428,N_15952,N_19815);
xor U20429 (N_20429,N_18628,N_15670);
nor U20430 (N_20430,N_19868,N_16611);
nor U20431 (N_20431,N_19294,N_19942);
xnor U20432 (N_20432,N_15683,N_16853);
and U20433 (N_20433,N_18618,N_18568);
xnor U20434 (N_20434,N_18793,N_16993);
nand U20435 (N_20435,N_17141,N_15522);
or U20436 (N_20436,N_19704,N_15462);
or U20437 (N_20437,N_15732,N_19375);
nand U20438 (N_20438,N_15716,N_18650);
xor U20439 (N_20439,N_18367,N_16746);
nor U20440 (N_20440,N_19081,N_18139);
and U20441 (N_20441,N_18770,N_15063);
or U20442 (N_20442,N_15605,N_17629);
xnor U20443 (N_20443,N_18373,N_16338);
xor U20444 (N_20444,N_17529,N_16011);
nor U20445 (N_20445,N_16061,N_15651);
and U20446 (N_20446,N_15017,N_19266);
nor U20447 (N_20447,N_16019,N_19568);
xor U20448 (N_20448,N_17100,N_15612);
or U20449 (N_20449,N_19388,N_19750);
nand U20450 (N_20450,N_18783,N_15498);
nor U20451 (N_20451,N_16110,N_15934);
or U20452 (N_20452,N_18907,N_17427);
and U20453 (N_20453,N_18421,N_17900);
nand U20454 (N_20454,N_15220,N_16022);
xnor U20455 (N_20455,N_17153,N_17106);
and U20456 (N_20456,N_18115,N_18370);
nand U20457 (N_20457,N_18073,N_15690);
xnor U20458 (N_20458,N_19268,N_18750);
or U20459 (N_20459,N_16164,N_16799);
nand U20460 (N_20460,N_16878,N_16241);
nor U20461 (N_20461,N_19491,N_19970);
xnor U20462 (N_20462,N_16362,N_15780);
xnor U20463 (N_20463,N_17393,N_17547);
nand U20464 (N_20464,N_15851,N_18752);
or U20465 (N_20465,N_17560,N_15555);
nand U20466 (N_20466,N_17584,N_17052);
nand U20467 (N_20467,N_15171,N_15399);
and U20468 (N_20468,N_15894,N_18463);
xnor U20469 (N_20469,N_19005,N_19174);
nor U20470 (N_20470,N_18610,N_19687);
xnor U20471 (N_20471,N_16559,N_17029);
nor U20472 (N_20472,N_19038,N_16071);
or U20473 (N_20473,N_15558,N_15408);
nand U20474 (N_20474,N_15289,N_18322);
nor U20475 (N_20475,N_19814,N_18070);
nand U20476 (N_20476,N_15452,N_15197);
and U20477 (N_20477,N_18097,N_16480);
nand U20478 (N_20478,N_17121,N_18382);
xor U20479 (N_20479,N_16849,N_17444);
nand U20480 (N_20480,N_16640,N_17530);
nand U20481 (N_20481,N_19698,N_16759);
nand U20482 (N_20482,N_17559,N_17343);
nor U20483 (N_20483,N_19564,N_19042);
nor U20484 (N_20484,N_16772,N_17439);
and U20485 (N_20485,N_19668,N_19115);
xor U20486 (N_20486,N_19696,N_19613);
nor U20487 (N_20487,N_16481,N_17279);
xnor U20488 (N_20488,N_18362,N_16225);
and U20489 (N_20489,N_17278,N_19833);
and U20490 (N_20490,N_19940,N_15621);
nand U20491 (N_20491,N_16170,N_17678);
and U20492 (N_20492,N_18698,N_19561);
and U20493 (N_20493,N_16332,N_16603);
nand U20494 (N_20494,N_18886,N_18528);
xnor U20495 (N_20495,N_16763,N_19457);
or U20496 (N_20496,N_19258,N_18170);
xnor U20497 (N_20497,N_15630,N_15459);
and U20498 (N_20498,N_15814,N_18581);
nand U20499 (N_20499,N_15056,N_19665);
or U20500 (N_20500,N_18482,N_18123);
xor U20501 (N_20501,N_17357,N_16827);
nand U20502 (N_20502,N_15416,N_19160);
xor U20503 (N_20503,N_15136,N_15019);
xnor U20504 (N_20504,N_17271,N_17813);
xnor U20505 (N_20505,N_18416,N_19307);
and U20506 (N_20506,N_16195,N_18464);
nand U20507 (N_20507,N_16749,N_17605);
or U20508 (N_20508,N_17586,N_16960);
xor U20509 (N_20509,N_16299,N_19431);
or U20510 (N_20510,N_16440,N_18567);
xnor U20511 (N_20511,N_18318,N_17656);
and U20512 (N_20512,N_16688,N_15015);
xnor U20513 (N_20513,N_17235,N_18485);
xnor U20514 (N_20514,N_15334,N_17440);
xor U20515 (N_20515,N_19416,N_19325);
or U20516 (N_20516,N_16991,N_16513);
or U20517 (N_20517,N_17028,N_17190);
nor U20518 (N_20518,N_17257,N_16900);
or U20519 (N_20519,N_18539,N_19413);
and U20520 (N_20520,N_18406,N_15992);
or U20521 (N_20521,N_18238,N_17403);
xnor U20522 (N_20522,N_15962,N_16996);
nor U20523 (N_20523,N_18102,N_16893);
nand U20524 (N_20524,N_19517,N_19112);
xnor U20525 (N_20525,N_16564,N_15214);
nand U20526 (N_20526,N_18030,N_18764);
nor U20527 (N_20527,N_18179,N_15047);
nand U20528 (N_20528,N_18267,N_17797);
xnor U20529 (N_20529,N_18048,N_19097);
nand U20530 (N_20530,N_18453,N_16571);
xnor U20531 (N_20531,N_18389,N_17286);
nor U20532 (N_20532,N_19365,N_15787);
and U20533 (N_20533,N_17177,N_19444);
and U20534 (N_20534,N_18708,N_15950);
nand U20535 (N_20535,N_16368,N_16436);
xor U20536 (N_20536,N_15634,N_15778);
and U20537 (N_20537,N_17298,N_18457);
or U20538 (N_20538,N_19374,N_15753);
xnor U20539 (N_20539,N_19749,N_16281);
xnor U20540 (N_20540,N_15093,N_19532);
xnor U20541 (N_20541,N_19954,N_15912);
and U20542 (N_20542,N_16633,N_17612);
nand U20543 (N_20543,N_19347,N_18941);
nor U20544 (N_20544,N_18347,N_18053);
nor U20545 (N_20545,N_17027,N_18327);
xor U20546 (N_20546,N_15521,N_16291);
xor U20547 (N_20547,N_19229,N_18979);
xor U20548 (N_20548,N_17379,N_17643);
nor U20549 (N_20549,N_15144,N_16850);
xnor U20550 (N_20550,N_18038,N_16314);
or U20551 (N_20551,N_17342,N_15590);
nor U20552 (N_20552,N_16556,N_16720);
nor U20553 (N_20553,N_16239,N_19035);
nor U20554 (N_20554,N_15281,N_19708);
xor U20555 (N_20555,N_15304,N_15109);
and U20556 (N_20556,N_16678,N_19368);
xnor U20557 (N_20557,N_17745,N_16057);
xnor U20558 (N_20558,N_15362,N_19287);
nor U20559 (N_20559,N_19516,N_19078);
or U20560 (N_20560,N_15013,N_15935);
or U20561 (N_20561,N_16487,N_15280);
nor U20562 (N_20562,N_16306,N_15400);
nor U20563 (N_20563,N_16263,N_16636);
nor U20564 (N_20564,N_19448,N_18281);
or U20565 (N_20565,N_17049,N_16033);
nand U20566 (N_20566,N_19664,N_17694);
xnor U20567 (N_20567,N_19313,N_18535);
xnor U20568 (N_20568,N_18746,N_15278);
or U20569 (N_20569,N_15149,N_19296);
and U20570 (N_20570,N_15655,N_17064);
nand U20571 (N_20571,N_18613,N_16545);
nor U20572 (N_20572,N_18707,N_17463);
and U20573 (N_20573,N_15587,N_18995);
and U20574 (N_20574,N_18666,N_18864);
or U20575 (N_20575,N_19996,N_15264);
nor U20576 (N_20576,N_19086,N_18673);
nor U20577 (N_20577,N_15914,N_17142);
and U20578 (N_20578,N_16936,N_16762);
nor U20579 (N_20579,N_17009,N_15724);
xnor U20580 (N_20580,N_19877,N_19290);
or U20581 (N_20581,N_19987,N_19123);
nor U20582 (N_20582,N_17646,N_18124);
and U20583 (N_20583,N_17766,N_18930);
or U20584 (N_20584,N_18129,N_18448);
nor U20585 (N_20585,N_16128,N_19052);
or U20586 (N_20586,N_18277,N_17084);
nor U20587 (N_20587,N_18833,N_19807);
nand U20588 (N_20588,N_15957,N_18566);
and U20589 (N_20589,N_17496,N_19870);
nor U20590 (N_20590,N_16433,N_19206);
xnor U20591 (N_20591,N_18282,N_18848);
or U20592 (N_20592,N_16030,N_17228);
or U20593 (N_20593,N_19658,N_19906);
nor U20594 (N_20594,N_18154,N_16403);
and U20595 (N_20595,N_18766,N_16708);
or U20596 (N_20596,N_16689,N_17868);
and U20597 (N_20597,N_16185,N_18626);
and U20598 (N_20598,N_17175,N_16448);
or U20599 (N_20599,N_16434,N_17397);
nand U20600 (N_20600,N_19606,N_17447);
nand U20601 (N_20601,N_16007,N_17969);
nor U20602 (N_20602,N_16072,N_17149);
or U20603 (N_20603,N_17134,N_19098);
xnor U20604 (N_20604,N_15096,N_15783);
and U20605 (N_20605,N_16182,N_17144);
nand U20606 (N_20606,N_19542,N_15972);
xnor U20607 (N_20607,N_17288,N_18511);
xor U20608 (N_20608,N_19901,N_18917);
and U20609 (N_20609,N_15527,N_18801);
xor U20610 (N_20610,N_18332,N_17072);
or U20611 (N_20611,N_19591,N_16304);
nor U20612 (N_20612,N_15417,N_17005);
and U20613 (N_20613,N_15150,N_15821);
nor U20614 (N_20614,N_15513,N_16656);
xnor U20615 (N_20615,N_18035,N_19302);
nand U20616 (N_20616,N_19237,N_16114);
or U20617 (N_20617,N_17306,N_15434);
or U20618 (N_20618,N_19701,N_15106);
and U20619 (N_20619,N_19754,N_19274);
nand U20620 (N_20620,N_15879,N_16363);
nor U20621 (N_20621,N_17905,N_19811);
nand U20622 (N_20622,N_17942,N_18311);
and U20623 (N_20623,N_19955,N_15647);
and U20624 (N_20624,N_19923,N_15650);
nand U20625 (N_20625,N_19007,N_19158);
and U20626 (N_20626,N_17531,N_17948);
nor U20627 (N_20627,N_17410,N_16407);
nor U20628 (N_20628,N_15325,N_18285);
nor U20629 (N_20629,N_17264,N_17184);
xor U20630 (N_20630,N_16775,N_16267);
xnor U20631 (N_20631,N_16040,N_16121);
nor U20632 (N_20632,N_15209,N_15180);
nor U20633 (N_20633,N_17616,N_19312);
xnor U20634 (N_20634,N_19994,N_17865);
nor U20635 (N_20635,N_17717,N_18052);
nor U20636 (N_20636,N_15726,N_18830);
nand U20637 (N_20637,N_18875,N_17040);
and U20638 (N_20638,N_15673,N_17415);
and U20639 (N_20639,N_16421,N_18101);
nor U20640 (N_20640,N_18713,N_18762);
xor U20641 (N_20641,N_17660,N_19897);
xor U20642 (N_20642,N_16942,N_15838);
nor U20643 (N_20643,N_19964,N_19530);
nor U20644 (N_20644,N_16560,N_17051);
nand U20645 (N_20645,N_16694,N_16422);
nand U20646 (N_20646,N_18725,N_15691);
nand U20647 (N_20647,N_17061,N_18061);
and U20648 (N_20648,N_16204,N_16541);
nor U20649 (N_20649,N_15674,N_17686);
nand U20650 (N_20650,N_15386,N_16105);
and U20651 (N_20651,N_15788,N_16747);
xnor U20652 (N_20652,N_18696,N_19640);
or U20653 (N_20653,N_19672,N_15438);
and U20654 (N_20654,N_19555,N_18401);
xnor U20655 (N_20655,N_15847,N_15900);
and U20656 (N_20656,N_15305,N_17985);
xor U20657 (N_20657,N_19095,N_16540);
or U20658 (N_20658,N_17110,N_19760);
nand U20659 (N_20659,N_17358,N_18006);
or U20660 (N_20660,N_19711,N_16526);
nor U20661 (N_20661,N_18489,N_16006);
or U20662 (N_20662,N_16176,N_18295);
nand U20663 (N_20663,N_19772,N_19830);
and U20664 (N_20664,N_15054,N_15575);
nand U20665 (N_20665,N_17290,N_19419);
or U20666 (N_20666,N_17802,N_17363);
or U20667 (N_20667,N_15586,N_15222);
nand U20668 (N_20668,N_16352,N_17060);
nor U20669 (N_20669,N_15842,N_19340);
nand U20670 (N_20670,N_19735,N_19685);
nand U20671 (N_20671,N_19813,N_16467);
nor U20672 (N_20672,N_15007,N_19660);
nor U20673 (N_20673,N_16938,N_15877);
xor U20674 (N_20674,N_19680,N_16612);
xor U20675 (N_20675,N_16090,N_17349);
or U20676 (N_20676,N_18739,N_18443);
or U20677 (N_20677,N_17311,N_15257);
xnor U20678 (N_20678,N_17615,N_19225);
nor U20679 (N_20679,N_18243,N_17908);
and U20680 (N_20680,N_16286,N_17753);
and U20681 (N_20681,N_16860,N_15979);
nand U20682 (N_20682,N_18148,N_17589);
nand U20683 (N_20683,N_18268,N_16552);
and U20684 (N_20684,N_17648,N_19068);
nand U20685 (N_20685,N_18319,N_16361);
nor U20686 (N_20686,N_19659,N_16202);
and U20687 (N_20687,N_16889,N_15508);
nand U20688 (N_20688,N_17075,N_15385);
xor U20689 (N_20689,N_16627,N_15095);
xor U20690 (N_20690,N_19057,N_18823);
nor U20691 (N_20691,N_18265,N_19376);
nand U20692 (N_20692,N_17103,N_17457);
or U20693 (N_20693,N_19142,N_16593);
nand U20694 (N_20694,N_17243,N_18424);
xor U20695 (N_20695,N_15775,N_18495);
and U20696 (N_20696,N_19253,N_15925);
nand U20697 (N_20697,N_16669,N_15540);
xor U20698 (N_20698,N_17990,N_18203);
and U20699 (N_20699,N_17607,N_15779);
nand U20700 (N_20700,N_16967,N_19403);
or U20701 (N_20701,N_19733,N_16855);
and U20702 (N_20702,N_16077,N_16641);
or U20703 (N_20703,N_18076,N_16657);
or U20704 (N_20704,N_15929,N_16891);
nand U20705 (N_20705,N_17627,N_16268);
xor U20706 (N_20706,N_17736,N_19154);
or U20707 (N_20707,N_19139,N_16981);
xor U20708 (N_20708,N_15460,N_17011);
or U20709 (N_20709,N_15529,N_17632);
nor U20710 (N_20710,N_15287,N_18747);
nand U20711 (N_20711,N_15226,N_19019);
nand U20712 (N_20712,N_19015,N_18304);
or U20713 (N_20713,N_19654,N_15616);
or U20714 (N_20714,N_17881,N_16735);
xnor U20715 (N_20715,N_19740,N_19327);
nor U20716 (N_20716,N_18135,N_15870);
or U20717 (N_20717,N_18196,N_17401);
and U20718 (N_20718,N_15475,N_17158);
xnor U20719 (N_20719,N_16535,N_18742);
nor U20720 (N_20720,N_16277,N_17789);
xnor U20721 (N_20721,N_19127,N_19943);
nand U20722 (N_20722,N_15137,N_17081);
xor U20723 (N_20723,N_15899,N_17200);
nand U20724 (N_20724,N_18985,N_18664);
xor U20725 (N_20725,N_18287,N_17663);
nor U20726 (N_20726,N_18976,N_18506);
and U20727 (N_20727,N_15121,N_15414);
xor U20728 (N_20728,N_15709,N_17834);
and U20729 (N_20729,N_16466,N_18116);
and U20730 (N_20730,N_15488,N_15286);
nand U20731 (N_20731,N_15811,N_16187);
or U20732 (N_20732,N_15617,N_19512);
xor U20733 (N_20733,N_19196,N_19969);
nand U20734 (N_20734,N_16334,N_18771);
and U20735 (N_20735,N_18769,N_19825);
nand U20736 (N_20736,N_16677,N_18993);
nor U20737 (N_20737,N_15589,N_19278);
or U20738 (N_20738,N_18807,N_19662);
nand U20739 (N_20739,N_18227,N_18997);
nand U20740 (N_20740,N_18608,N_18923);
nor U20741 (N_20741,N_18353,N_17764);
and U20742 (N_20742,N_18894,N_17242);
nand U20743 (N_20743,N_15083,N_16380);
and U20744 (N_20744,N_19900,N_15263);
xnor U20745 (N_20745,N_15653,N_16290);
or U20746 (N_20746,N_18283,N_16075);
and U20747 (N_20747,N_15991,N_16476);
and U20748 (N_20748,N_16206,N_19214);
or U20749 (N_20749,N_15582,N_18540);
nand U20750 (N_20750,N_17528,N_15424);
or U20751 (N_20751,N_19739,N_17919);
nor U20752 (N_20752,N_16870,N_15614);
xnor U20753 (N_20753,N_16770,N_18534);
nor U20754 (N_20754,N_18623,N_19149);
nor U20755 (N_20755,N_19106,N_15456);
or U20756 (N_20756,N_19138,N_17941);
nand U20757 (N_20757,N_16346,N_15965);
nand U20758 (N_20758,N_17903,N_16138);
xnor U20759 (N_20759,N_15184,N_15094);
or U20760 (N_20760,N_19783,N_18004);
and U20761 (N_20761,N_17256,N_16760);
or U20762 (N_20762,N_17691,N_17265);
xnor U20763 (N_20763,N_16687,N_19396);
xnor U20764 (N_20764,N_19936,N_18521);
nand U20765 (N_20765,N_16764,N_15135);
nand U20766 (N_20766,N_15169,N_17076);
or U20767 (N_20767,N_18558,N_18838);
nor U20768 (N_20768,N_16531,N_15832);
xnor U20769 (N_20769,N_16562,N_15229);
or U20770 (N_20770,N_16078,N_19851);
xnor U20771 (N_20771,N_17442,N_19986);
or U20772 (N_20772,N_19061,N_16892);
nand U20773 (N_20773,N_16372,N_15157);
and U20774 (N_20774,N_16366,N_16621);
nand U20775 (N_20775,N_19372,N_19681);
nand U20776 (N_20776,N_19193,N_15544);
nor U20777 (N_20777,N_15887,N_17949);
nand U20778 (N_20778,N_16094,N_19040);
or U20779 (N_20779,N_16478,N_16800);
and U20780 (N_20780,N_19932,N_16653);
nand U20781 (N_20781,N_19789,N_18086);
nor U20782 (N_20782,N_18091,N_19114);
or U20783 (N_20783,N_16410,N_18313);
and U20784 (N_20784,N_16661,N_15904);
nor U20785 (N_20785,N_19026,N_17651);
nor U20786 (N_20786,N_18763,N_15702);
xnor U20787 (N_20787,N_18260,N_18250);
nor U20788 (N_20788,N_18080,N_18399);
xor U20789 (N_20789,N_19198,N_19611);
and U20790 (N_20790,N_16925,N_19666);
nor U20791 (N_20791,N_15622,N_15737);
and U20792 (N_20792,N_17765,N_16660);
and U20793 (N_20793,N_17653,N_17448);
xor U20794 (N_20794,N_15871,N_16432);
nor U20795 (N_20795,N_16992,N_15190);
or U20796 (N_20796,N_15039,N_17923);
nor U20797 (N_20797,N_19456,N_16879);
xor U20798 (N_20798,N_16789,N_17095);
nor U20799 (N_20799,N_18344,N_18114);
or U20800 (N_20800,N_15628,N_18645);
nand U20801 (N_20801,N_17091,N_15846);
nor U20802 (N_20802,N_19966,N_17578);
nor U20803 (N_20803,N_16734,N_18142);
and U20804 (N_20804,N_18921,N_19838);
nor U20805 (N_20805,N_18522,N_19856);
nor U20806 (N_20806,N_17721,N_15084);
or U20807 (N_20807,N_19475,N_17145);
nor U20808 (N_20808,N_18315,N_16858);
nor U20809 (N_20809,N_17126,N_19116);
nand U20810 (N_20810,N_18157,N_19853);
or U20811 (N_20811,N_19254,N_18632);
xnor U20812 (N_20812,N_15857,N_16567);
nand U20813 (N_20813,N_15499,N_16565);
xnor U20814 (N_20814,N_17710,N_19036);
xnor U20815 (N_20815,N_15949,N_17782);
xnor U20816 (N_20816,N_16511,N_16192);
or U20817 (N_20817,N_19319,N_15795);
or U20818 (N_20818,N_18736,N_15998);
xnor U20819 (N_20819,N_17636,N_16966);
and U20820 (N_20820,N_18180,N_16167);
xnor U20821 (N_20821,N_17759,N_17570);
nand U20822 (N_20822,N_15640,N_18523);
and U20823 (N_20823,N_18741,N_16521);
or U20824 (N_20824,N_16809,N_16802);
or U20825 (N_20825,N_19904,N_17493);
or U20826 (N_20826,N_16907,N_19828);
and U20827 (N_20827,N_16152,N_15875);
nand U20828 (N_20828,N_18312,N_18802);
or U20829 (N_20829,N_15493,N_18418);
or U20830 (N_20830,N_17347,N_18150);
nor U20831 (N_20831,N_18636,N_15872);
or U20832 (N_20832,N_18252,N_17999);
nand U20833 (N_20833,N_17481,N_17770);
and U20834 (N_20834,N_16727,N_19880);
and U20835 (N_20835,N_18710,N_16574);
or U20836 (N_20836,N_15581,N_19292);
nor U20837 (N_20837,N_16184,N_18303);
nand U20838 (N_20838,N_19462,N_15040);
xor U20839 (N_20839,N_19578,N_18513);
nor U20840 (N_20840,N_15132,N_16454);
and U20841 (N_20841,N_18133,N_17355);
and U20842 (N_20842,N_19496,N_19793);
and U20843 (N_20843,N_15802,N_17482);
xnor U20844 (N_20844,N_15543,N_15026);
or U20845 (N_20845,N_19181,N_19212);
xnor U20846 (N_20846,N_18704,N_19247);
nand U20847 (N_20847,N_18063,N_18602);
or U20848 (N_20848,N_19505,N_16379);
and U20849 (N_20849,N_15876,N_19251);
or U20850 (N_20850,N_19860,N_18462);
or U20851 (N_20851,N_16710,N_19315);
nor U20852 (N_20852,N_18477,N_15238);
nand U20853 (N_20853,N_19050,N_19945);
xnor U20854 (N_20854,N_16712,N_15836);
xor U20855 (N_20855,N_18171,N_17404);
nor U20856 (N_20856,N_18959,N_15501);
or U20857 (N_20857,N_19863,N_19669);
nand U20858 (N_20858,N_19547,N_16791);
nand U20859 (N_20859,N_18646,N_17513);
nand U20860 (N_20860,N_15421,N_16623);
nor U20861 (N_20861,N_18653,N_19144);
and U20862 (N_20862,N_16357,N_15181);
and U20863 (N_20863,N_18712,N_17723);
nor U20864 (N_20864,N_16226,N_17866);
and U20865 (N_20865,N_18638,N_16638);
and U20866 (N_20866,N_19963,N_17254);
and U20867 (N_20867,N_18805,N_19802);
xor U20868 (N_20868,N_18175,N_16652);
or U20869 (N_20869,N_16127,N_18291);
and U20870 (N_20870,N_17982,N_15345);
xor U20871 (N_20871,N_18297,N_19949);
and U20872 (N_20872,N_17365,N_15042);
or U20873 (N_20873,N_17302,N_18547);
and U20874 (N_20874,N_16234,N_19137);
nand U20875 (N_20875,N_19907,N_18850);
nand U20876 (N_20876,N_15641,N_15947);
nand U20877 (N_20877,N_16584,N_17225);
xnor U20878 (N_20878,N_16320,N_15704);
xnor U20879 (N_20879,N_16507,N_19761);
nand U20880 (N_20880,N_17082,N_19629);
and U20881 (N_20881,N_18455,N_16074);
or U20882 (N_20882,N_15119,N_18786);
or U20883 (N_20883,N_15074,N_19164);
xor U20884 (N_20884,N_18158,N_16949);
xor U20885 (N_20885,N_16310,N_17561);
or U20886 (N_20886,N_18374,N_15114);
or U20887 (N_20887,N_16001,N_15033);
nand U20888 (N_20888,N_18614,N_16926);
or U20889 (N_20889,N_17312,N_17769);
and U20890 (N_20890,N_17738,N_15791);
nand U20891 (N_20891,N_15183,N_19605);
nor U20892 (N_20892,N_17275,N_19210);
and U20893 (N_20893,N_18220,N_17419);
nand U20894 (N_20894,N_18491,N_16489);
xnor U20895 (N_20895,N_17835,N_16137);
xor U20896 (N_20896,N_19163,N_18206);
nand U20897 (N_20897,N_15903,N_15293);
nor U20898 (N_20898,N_17114,N_16999);
or U20899 (N_20899,N_17226,N_19948);
or U20900 (N_20900,N_17458,N_16271);
xor U20901 (N_20901,N_17703,N_16065);
or U20902 (N_20902,N_15557,N_17596);
nor U20903 (N_20903,N_19343,N_17150);
or U20904 (N_20904,N_17151,N_16331);
nand U20905 (N_20905,N_18183,N_19746);
and U20906 (N_20906,N_19121,N_18554);
and U20907 (N_20907,N_17086,N_19141);
nand U20908 (N_20908,N_17181,N_19260);
nand U20909 (N_20909,N_18914,N_16103);
and U20910 (N_20910,N_19499,N_17161);
nor U20911 (N_20911,N_19393,N_18486);
and U20912 (N_20912,N_19684,N_15361);
nor U20913 (N_20913,N_19209,N_16663);
nand U20914 (N_20914,N_17811,N_17841);
xnor U20915 (N_20915,N_18033,N_16758);
or U20916 (N_20916,N_17360,N_17160);
and U20917 (N_20917,N_19543,N_16670);
nand U20918 (N_20918,N_18938,N_18155);
xor U20919 (N_20919,N_17957,N_19682);
or U20920 (N_20920,N_19525,N_18681);
or U20921 (N_20921,N_19310,N_19146);
xnor U20922 (N_20922,N_19764,N_19119);
nor U20923 (N_20923,N_19492,N_17974);
nor U20924 (N_20924,N_16527,N_16344);
xor U20925 (N_20925,N_18254,N_19065);
and U20926 (N_20926,N_17387,N_19168);
nor U20927 (N_20927,N_16285,N_17920);
xnor U20928 (N_20928,N_18893,N_17172);
xnor U20929 (N_20929,N_18951,N_15080);
xor U20930 (N_20930,N_15251,N_16905);
and U20931 (N_20931,N_18144,N_15392);
or U20932 (N_20932,N_16051,N_18831);
or U20933 (N_20933,N_17964,N_16093);
nand U20934 (N_20934,N_18223,N_19584);
xor U20935 (N_20935,N_18683,N_15486);
xnor U20936 (N_20936,N_18333,N_16235);
nor U20937 (N_20937,N_18789,N_18835);
nand U20938 (N_20938,N_19379,N_18961);
and U20939 (N_20939,N_19455,N_18377);
xor U20940 (N_20940,N_15917,N_17666);
or U20941 (N_20941,N_19072,N_17354);
xor U20942 (N_20942,N_19079,N_19391);
xor U20943 (N_20943,N_19243,N_15881);
or U20944 (N_20944,N_17485,N_17332);
nor U20945 (N_20945,N_17670,N_19902);
and U20946 (N_20946,N_19366,N_16032);
or U20947 (N_20947,N_17437,N_15436);
nor U20948 (N_20948,N_15154,N_19445);
or U20949 (N_20949,N_18691,N_15748);
nor U20950 (N_20950,N_19777,N_17420);
or U20951 (N_20951,N_16899,N_18928);
xnor U20952 (N_20952,N_19345,N_15262);
and U20953 (N_20953,N_16080,N_17880);
xor U20954 (N_20954,N_18334,N_17707);
xnor U20955 (N_20955,N_15346,N_17034);
and U20956 (N_20956,N_18216,N_15528);
or U20957 (N_20957,N_19273,N_19642);
or U20958 (N_20958,N_17809,N_18982);
nand U20959 (N_20959,N_16510,N_18659);
nand U20960 (N_20960,N_16530,N_19589);
nor U20961 (N_20961,N_15127,N_19284);
or U20962 (N_20962,N_16153,N_18992);
or U20963 (N_20963,N_15719,N_17775);
and U20964 (N_20964,N_18587,N_15333);
xor U20965 (N_20965,N_19816,N_19527);
nand U20966 (N_20966,N_18967,N_18744);
and U20967 (N_20967,N_18640,N_19175);
xor U20968 (N_20968,N_16795,N_16917);
nor U20969 (N_20969,N_15016,N_19759);
nor U20970 (N_20970,N_16977,N_19326);
and U20971 (N_20971,N_18369,N_15675);
nand U20972 (N_20972,N_19330,N_19592);
xnor U20973 (N_20973,N_19013,N_15735);
xor U20974 (N_20974,N_15426,N_17628);
nand U20975 (N_20975,N_16319,N_16843);
nor U20976 (N_20976,N_17992,N_18731);
and U20977 (N_20977,N_18620,N_18897);
nand U20978 (N_20978,N_18425,N_17066);
nand U20979 (N_20979,N_16748,N_16307);
xnor U20980 (N_20980,N_16274,N_17014);
nor U20981 (N_20981,N_18163,N_16783);
nand U20982 (N_20982,N_18205,N_19882);
nor U20983 (N_20983,N_15829,N_18084);
or U20984 (N_20984,N_16219,N_18944);
nor U20985 (N_20985,N_17692,N_16143);
or U20986 (N_20986,N_17577,N_19381);
nand U20987 (N_20987,N_19255,N_17952);
and U20988 (N_20988,N_17108,N_19357);
nand U20989 (N_20989,N_17885,N_17593);
nand U20990 (N_20990,N_15196,N_18027);
nand U20991 (N_20991,N_16819,N_15626);
and U20992 (N_20992,N_17018,N_18884);
nor U20993 (N_20993,N_16649,N_18194);
xnor U20994 (N_20994,N_19751,N_16975);
or U20995 (N_20995,N_16756,N_17971);
xnor U20996 (N_20996,N_15721,N_15188);
xnor U20997 (N_20997,N_16600,N_18007);
nor U20998 (N_20998,N_17894,N_18836);
nand U20999 (N_20999,N_15705,N_19032);
nor U21000 (N_21000,N_19707,N_15261);
nor U21001 (N_21001,N_18735,N_18323);
and U21002 (N_21002,N_18732,N_16824);
or U21003 (N_21003,N_19264,N_18164);
nor U21004 (N_21004,N_15355,N_15573);
nand U21005 (N_21005,N_18099,N_19720);
xnor U21006 (N_21006,N_19717,N_19596);
xor U21007 (N_21007,N_18385,N_19199);
xnor U21008 (N_21008,N_16413,N_19820);
and U21009 (N_21009,N_16201,N_18728);
or U21010 (N_21010,N_19959,N_18055);
or U21011 (N_21011,N_16369,N_18768);
or U21012 (N_21012,N_16386,N_15785);
nand U21013 (N_21013,N_19389,N_17069);
xnor U21014 (N_21014,N_19369,N_16866);
xnor U21015 (N_21015,N_16707,N_18409);
xnor U21016 (N_21016,N_18964,N_18784);
or U21017 (N_21017,N_19421,N_19822);
and U21018 (N_21018,N_16070,N_17085);
or U21019 (N_21019,N_19985,N_18379);
nand U21020 (N_21020,N_18230,N_16961);
or U21021 (N_21021,N_19878,N_19805);
nand U21022 (N_21022,N_17760,N_17206);
xnor U21023 (N_21023,N_16516,N_19545);
or U21024 (N_21024,N_17308,N_16197);
or U21025 (N_21025,N_15895,N_15754);
nand U21026 (N_21026,N_17859,N_18779);
xnor U21027 (N_21027,N_19021,N_16404);
nand U21028 (N_21028,N_19978,N_16328);
nor U21029 (N_21029,N_16161,N_17315);
xor U21030 (N_21030,N_16060,N_17819);
and U21031 (N_21031,N_18445,N_17571);
or U21032 (N_21032,N_16181,N_19058);
xnor U21033 (N_21033,N_18849,N_15596);
nand U21034 (N_21034,N_18740,N_16928);
or U21035 (N_21035,N_16505,N_15994);
and U21036 (N_21036,N_18244,N_18847);
nor U21037 (N_21037,N_19744,N_17473);
xor U21038 (N_21038,N_15858,N_15193);
and U21039 (N_21039,N_17333,N_18130);
nand U21040 (N_21040,N_19501,N_15216);
nand U21041 (N_21041,N_16769,N_16632);
or U21042 (N_21042,N_18224,N_18320);
and U21043 (N_21043,N_17131,N_15246);
nor U21044 (N_21044,N_16125,N_16035);
xnor U21045 (N_21045,N_19412,N_19222);
xnor U21046 (N_21046,N_17917,N_15708);
xor U21047 (N_21047,N_16538,N_18935);
or U21048 (N_21048,N_15720,N_16000);
nor U21049 (N_21049,N_18094,N_18019);
xnor U21050 (N_21050,N_17258,N_19826);
nor U21051 (N_21051,N_19500,N_15466);
nor U21052 (N_21052,N_19769,N_16589);
nand U21053 (N_21053,N_17491,N_16166);
or U21054 (N_21054,N_16425,N_18469);
nor U21055 (N_21055,N_18757,N_15274);
nor U21056 (N_21056,N_15703,N_15603);
nand U21057 (N_21057,N_18496,N_16190);
nand U21058 (N_21058,N_16099,N_18381);
or U21059 (N_21059,N_15715,N_15046);
xor U21060 (N_21060,N_19208,N_15429);
nor U21061 (N_21061,N_19827,N_15841);
nand U21062 (N_21062,N_16923,N_17882);
and U21063 (N_21063,N_18258,N_18444);
nor U21064 (N_21064,N_19781,N_16751);
or U21065 (N_21065,N_18269,N_17402);
nand U21066 (N_21066,N_19590,N_15571);
xor U21067 (N_21067,N_19976,N_19280);
or U21068 (N_21068,N_17762,N_16159);
nand U21069 (N_21069,N_16147,N_15234);
or U21070 (N_21070,N_18773,N_15227);
nor U21071 (N_21071,N_19876,N_19166);
and U21072 (N_21072,N_15435,N_18913);
or U21073 (N_21073,N_15638,N_18637);
nor U21074 (N_21074,N_19619,N_15494);
and U21075 (N_21075,N_17139,N_17090);
xor U21076 (N_21076,N_19474,N_18074);
and U21077 (N_21077,N_17301,N_16815);
or U21078 (N_21078,N_17455,N_15500);
nor U21079 (N_21079,N_19467,N_16693);
xor U21080 (N_21080,N_15679,N_17573);
xor U21081 (N_21081,N_15968,N_19470);
or U21082 (N_21082,N_19770,N_18062);
nand U21083 (N_21083,N_18839,N_19399);
and U21084 (N_21084,N_18054,N_19965);
and U21085 (N_21085,N_19030,N_18066);
and U21086 (N_21086,N_17871,N_19242);
and U21087 (N_21087,N_15747,N_17940);
nor U21088 (N_21088,N_15202,N_15919);
nand U21089 (N_21089,N_16525,N_16655);
nor U21090 (N_21090,N_18550,N_19550);
nand U21091 (N_21091,N_15427,N_17093);
nand U21092 (N_21092,N_15339,N_16427);
or U21093 (N_21093,N_18350,N_19849);
and U21094 (N_21094,N_16084,N_15694);
nand U21095 (N_21095,N_18293,N_19747);
or U21096 (N_21096,N_16985,N_15087);
or U21097 (N_21097,N_19076,N_16264);
and U21098 (N_21098,N_17043,N_18134);
xor U21099 (N_21099,N_19692,N_19203);
xnor U21100 (N_21100,N_15681,N_18451);
xnor U21101 (N_21101,N_19528,N_17955);
xor U21102 (N_21102,N_16814,N_17170);
and U21103 (N_21103,N_17116,N_16430);
or U21104 (N_21104,N_15200,N_16131);
xor U21105 (N_21105,N_19756,N_18912);
and U21106 (N_21106,N_16553,N_16983);
nand U21107 (N_21107,N_15491,N_19521);
nand U21108 (N_21108,N_17844,N_16716);
and U21109 (N_21109,N_16778,N_17109);
xnor U21110 (N_21110,N_15863,N_16106);
or U21111 (N_21111,N_17958,N_19630);
or U21112 (N_21112,N_18122,N_17138);
xnor U21113 (N_21113,N_19031,N_18136);
or U21114 (N_21114,N_19858,N_19835);
or U21115 (N_21115,N_15824,N_19406);
or U21116 (N_21116,N_16292,N_18430);
or U21117 (N_21117,N_16939,N_15822);
and U21118 (N_21118,N_15482,N_15076);
xor U21119 (N_21119,N_15695,N_19321);
nand U21120 (N_21120,N_17500,N_16937);
or U21121 (N_21121,N_16305,N_19349);
or U21122 (N_21122,N_17125,N_16549);
nor U21123 (N_21123,N_17219,N_17046);
xor U21124 (N_21124,N_15743,N_15955);
nand U21125 (N_21125,N_16995,N_18590);
and U21126 (N_21126,N_17374,N_15812);
and U21127 (N_21127,N_15418,N_16351);
nand U21128 (N_21128,N_18684,N_15428);
and U21129 (N_21129,N_15902,N_18166);
nor U21130 (N_21130,N_15831,N_18840);
or U21131 (N_21131,N_17677,N_19100);
and U21132 (N_21132,N_18598,N_15376);
or U21133 (N_21133,N_17557,N_17983);
and U21134 (N_21134,N_18162,N_17266);
and U21135 (N_21135,N_17299,N_19039);
or U21136 (N_21136,N_17567,N_19766);
nand U21137 (N_21137,N_18064,N_16096);
or U21138 (N_21138,N_16104,N_16371);
nor U21139 (N_21139,N_18612,N_17998);
nand U21140 (N_21140,N_19184,N_18916);
or U21141 (N_21141,N_18767,N_19656);
nor U21142 (N_21142,N_16484,N_16576);
xor U21143 (N_21143,N_19218,N_17328);
and U21144 (N_21144,N_17245,N_19498);
or U21145 (N_21145,N_18508,N_19874);
nand U21146 (N_21146,N_16522,N_19051);
nor U21147 (N_21147,N_15070,N_19140);
nand U21148 (N_21148,N_17155,N_16682);
nor U21149 (N_21149,N_19741,N_17023);
or U21150 (N_21150,N_15342,N_18018);
xnor U21151 (N_21151,N_18719,N_19635);
and U21152 (N_21152,N_15130,N_16618);
or U21153 (N_21153,N_19529,N_16374);
nand U21154 (N_21154,N_15946,N_16021);
xnor U21155 (N_21155,N_19476,N_15299);
or U21156 (N_21156,N_17364,N_19048);
or U21157 (N_21157,N_17886,N_17490);
xor U21158 (N_21158,N_15930,N_17640);
nand U21159 (N_21159,N_17869,N_19628);
nor U21160 (N_21160,N_17671,N_15113);
nor U21161 (N_21161,N_15243,N_15153);
and U21162 (N_21162,N_18803,N_17020);
and U21163 (N_21163,N_17438,N_18096);
and U21164 (N_21164,N_18156,N_17568);
xor U21165 (N_21165,N_15738,N_19626);
xnor U21166 (N_21166,N_17169,N_19263);
nand U21167 (N_21167,N_15852,N_15727);
xor U21168 (N_21168,N_15336,N_15890);
nand U21169 (N_21169,N_16851,N_17385);
nand U21170 (N_21170,N_15828,N_18208);
and U21171 (N_21171,N_18209,N_15907);
nor U21172 (N_21172,N_18661,N_16321);
nand U21173 (N_21173,N_18509,N_17931);
nor U21174 (N_21174,N_15797,N_18987);
nand U21175 (N_21175,N_15585,N_15380);
nor U21176 (N_21176,N_15684,N_16169);
or U21177 (N_21177,N_16626,N_18868);
and U21178 (N_21178,N_18121,N_18676);
xnor U21179 (N_21179,N_18561,N_15613);
nand U21180 (N_21180,N_19103,N_19458);
nor U21181 (N_21181,N_18234,N_18414);
or U21182 (N_21182,N_17044,N_17366);
xnor U21183 (N_21183,N_17635,N_15363);
or U21184 (N_21184,N_17122,N_18494);
nor U21185 (N_21185,N_16546,N_18652);
or U21186 (N_21186,N_17872,N_18794);
nor U21187 (N_21187,N_16692,N_19881);
or U21188 (N_21188,N_18861,N_16517);
nor U21189 (N_21189,N_18621,N_19804);
nor U21190 (N_21190,N_18533,N_17006);
nor U21191 (N_21191,N_17384,N_18450);
xnor U21192 (N_21192,N_17339,N_18966);
xnor U21193 (N_21193,N_16300,N_16029);
and U21194 (N_21194,N_19054,N_19303);
nor U21195 (N_21195,N_17556,N_19487);
xnor U21196 (N_21196,N_16272,N_15259);
and U21197 (N_21197,N_16717,N_18846);
nor U21198 (N_21198,N_16958,N_19587);
nand U21199 (N_21199,N_16723,N_16223);
and U21200 (N_21200,N_18895,N_15763);
and U21201 (N_21201,N_17739,N_17606);
or U21202 (N_21202,N_18410,N_18256);
or U21203 (N_21203,N_18953,N_19495);
or U21204 (N_21204,N_16038,N_17291);
and U21205 (N_21205,N_16188,N_19683);
and U21206 (N_21206,N_18504,N_15559);
xor U21207 (N_21207,N_17870,N_16055);
and U21208 (N_21208,N_16634,N_17282);
or U21209 (N_21209,N_18772,N_15511);
nor U21210 (N_21210,N_15888,N_17048);
xnor U21211 (N_21211,N_18841,N_19033);
nand U21212 (N_21212,N_15883,N_19227);
and U21213 (N_21213,N_17261,N_19439);
xnor U21214 (N_21214,N_19951,N_17624);
nand U21215 (N_21215,N_15477,N_18083);
nand U21216 (N_21216,N_17025,N_15049);
xnor U21217 (N_21217,N_19661,N_19221);
nor U21218 (N_21218,N_19650,N_17204);
xor U21219 (N_21219,N_19973,N_17810);
xor U21220 (N_21220,N_17777,N_17980);
and U21221 (N_21221,N_17479,N_15447);
and U21222 (N_21222,N_16644,N_17508);
xnor U21223 (N_21223,N_18271,N_15971);
and U21224 (N_21224,N_16494,N_16950);
or U21225 (N_21225,N_16412,N_16659);
or U21226 (N_21226,N_15442,N_18947);
xor U21227 (N_21227,N_17572,N_16908);
xnor U21228 (N_21228,N_17667,N_15644);
xnor U21229 (N_21229,N_17833,N_18889);
nor U21230 (N_21230,N_19908,N_17944);
xor U21231 (N_21231,N_18514,N_17132);
or U21232 (N_21232,N_15224,N_15766);
or U21233 (N_21233,N_19339,N_17185);
or U21234 (N_21234,N_18404,N_16662);
or U21235 (N_21235,N_16081,N_15860);
nor U21236 (N_21236,N_17180,N_19771);
and U21237 (N_21237,N_19440,N_15696);
nor U21238 (N_21238,N_16378,N_18582);
nand U21239 (N_21239,N_16766,N_19919);
nand U21240 (N_21240,N_16586,N_19824);
xor U21241 (N_21241,N_17702,N_18393);
and U21242 (N_21242,N_15503,N_16423);
nand U21243 (N_21243,N_19649,N_15803);
and U21244 (N_21244,N_15985,N_17188);
nor U21245 (N_21245,N_18357,N_19129);
or U21246 (N_21246,N_15387,N_18289);
xor U21247 (N_21247,N_19653,N_18169);
and U21248 (N_21248,N_18780,N_19742);
and U21249 (N_21249,N_16014,N_15366);
or U21250 (N_21250,N_16676,N_17898);
nand U21251 (N_21251,N_17094,N_19479);
and U21252 (N_21252,N_19425,N_17758);
nand U21253 (N_21253,N_17398,N_16554);
or U21254 (N_21254,N_17337,N_17514);
nand U21255 (N_21255,N_15977,N_18898);
nand U21256 (N_21256,N_16667,N_16920);
and U21257 (N_21257,N_19075,N_15882);
xor U21258 (N_21258,N_16083,N_16550);
xor U21259 (N_21259,N_15920,N_15666);
nor U21260 (N_21260,N_16882,N_16887);
nor U21261 (N_21261,N_17558,N_17786);
nand U21262 (N_21262,N_18854,N_15913);
nor U21263 (N_21263,N_15245,N_15623);
nand U21264 (N_21264,N_19411,N_15898);
xnor U21265 (N_21265,N_17754,N_18722);
or U21266 (N_21266,N_19245,N_18218);
and U21267 (N_21267,N_17991,N_16395);
nand U21268 (N_21268,N_17800,N_16173);
nand U21269 (N_21269,N_17059,N_16465);
and U21270 (N_21270,N_17732,N_15323);
nor U21271 (N_21271,N_18185,N_17507);
nor U21272 (N_21272,N_17047,N_18191);
xnor U21273 (N_21273,N_17227,N_18296);
nor U21274 (N_21274,N_18392,N_19854);
xor U21275 (N_21275,N_16861,N_16449);
xnor U21276 (N_21276,N_16322,N_18024);
and U21277 (N_21277,N_19848,N_16027);
and U21278 (N_21278,N_19618,N_17913);
and U21279 (N_21279,N_17292,N_15897);
or U21280 (N_21280,N_16897,N_16470);
nor U21281 (N_21281,N_16063,N_19451);
and U21282 (N_21282,N_18996,N_17434);
nor U21283 (N_21283,N_15918,N_18588);
nor U21284 (N_21284,N_16266,N_19427);
or U21285 (N_21285,N_16598,N_16337);
xnor U21286 (N_21286,N_19913,N_16862);
xnor U21287 (N_21287,N_18025,N_16718);
nand U21288 (N_21288,N_18977,N_17749);
and U21289 (N_21289,N_18668,N_17087);
and U21290 (N_21290,N_17211,N_16706);
nor U21291 (N_21291,N_15051,N_16126);
xor U21292 (N_21292,N_17953,N_19995);
nand U21293 (N_21293,N_17238,N_18663);
xor U21294 (N_21294,N_19832,N_16722);
or U21295 (N_21295,N_17154,N_19246);
nand U21296 (N_21296,N_16733,N_16597);
and U21297 (N_21297,N_18247,N_17459);
and U21298 (N_21298,N_17664,N_15410);
xnor U21299 (N_21299,N_18215,N_16085);
xnor U21300 (N_21300,N_19645,N_19132);
or U21301 (N_21301,N_15986,N_17767);
xnor U21302 (N_21302,N_19609,N_15004);
and U21303 (N_21303,N_16854,N_17416);
nand U21304 (N_21304,N_16569,N_18082);
xor U21305 (N_21305,N_15632,N_18911);
and U21306 (N_21306,N_15177,N_19311);
or U21307 (N_21307,N_16324,N_16193);
nand U21308 (N_21308,N_18630,N_17281);
xor U21309 (N_21309,N_19056,N_19938);
xnor U21310 (N_21310,N_17314,N_18168);
nor U21311 (N_21311,N_18105,N_19306);
and U21312 (N_21312,N_18827,N_17937);
nor U21313 (N_21313,N_19067,N_18078);
and U21314 (N_21314,N_16233,N_19071);
xor U21315 (N_21315,N_15038,N_18545);
nand U21316 (N_21316,N_18518,N_15404);
nand U21317 (N_21317,N_16461,N_19522);
nand U21318 (N_21318,N_17506,N_15035);
and U21319 (N_21319,N_17807,N_18046);
xnor U21320 (N_21320,N_19156,N_15356);
nor U21321 (N_21321,N_18660,N_15595);
nand U21322 (N_21322,N_17554,N_18778);
and U21323 (N_21323,N_17350,N_17785);
or U21324 (N_21324,N_15604,N_19446);
nand U21325 (N_21325,N_17074,N_18316);
xnor U21326 (N_21326,N_15931,N_15248);
nor U21327 (N_21327,N_15377,N_18718);
xnor U21328 (N_21328,N_17436,N_15307);
or U21329 (N_21329,N_16834,N_16745);
and U21330 (N_21330,N_19910,N_15002);
or U21331 (N_21331,N_17409,N_17752);
and U21332 (N_21332,N_15510,N_16002);
or U21333 (N_21333,N_19433,N_17267);
nor U21334 (N_21334,N_18039,N_18388);
xor U21335 (N_21335,N_17956,N_16479);
or U21336 (N_21336,N_17240,N_17405);
nand U21337 (N_21337,N_15060,N_15509);
xor U21338 (N_21338,N_19879,N_15905);
xnor U21339 (N_21339,N_17532,N_16871);
and U21340 (N_21340,N_18026,N_18880);
and U21341 (N_21341,N_16829,N_17639);
xor U21342 (N_21342,N_15441,N_18527);
and U21343 (N_21343,N_17614,N_19864);
and U21344 (N_21344,N_19544,N_17477);
xor U21345 (N_21345,N_19925,N_18331);
nand U21346 (N_21346,N_17856,N_16895);
and U21347 (N_21347,N_18896,N_18306);
or U21348 (N_21348,N_18458,N_16901);
nor U21349 (N_21349,N_15723,N_15384);
xnor U21350 (N_21350,N_19834,N_19597);
xor U21351 (N_21351,N_18701,N_19275);
xnor U21352 (N_21352,N_18190,N_18826);
xnor U21353 (N_21353,N_19961,N_15707);
or U21354 (N_21354,N_15282,N_19603);
xnor U21355 (N_21355,N_19778,N_18824);
nor U21356 (N_21356,N_16666,N_18881);
and U21357 (N_21357,N_18605,N_18437);
xor U21358 (N_21358,N_19939,N_16097);
nand U21359 (N_21359,N_16801,N_18309);
nand U21360 (N_21360,N_18184,N_19148);
xor U21361 (N_21361,N_15948,N_19779);
and U21362 (N_21362,N_19145,N_16868);
xor U21363 (N_21363,N_16275,N_16588);
nor U21364 (N_21364,N_19857,N_16788);
or U21365 (N_21365,N_16509,N_19020);
or U21366 (N_21366,N_18774,N_16390);
xnor U21367 (N_21367,N_18117,N_15978);
xor U21368 (N_21368,N_19262,N_16409);
or U21369 (N_21369,N_15313,N_17781);
nand U21370 (N_21370,N_17934,N_15162);
xnor U21371 (N_21371,N_19842,N_18266);
and U21372 (N_21372,N_18072,N_15053);
or U21373 (N_21373,N_18290,N_15909);
nor U21374 (N_21374,N_19000,N_16629);
xor U21375 (N_21375,N_19248,N_18202);
and U21376 (N_21376,N_18197,N_16786);
nor U21377 (N_21377,N_19011,N_19493);
nor U21378 (N_21378,N_17883,N_19627);
nor U21379 (N_21379,N_15078,N_18759);
nand U21380 (N_21380,N_19437,N_19734);
xor U21381 (N_21381,N_15611,N_16194);
nor U21382 (N_21382,N_15868,N_18984);
and U21383 (N_21383,N_19991,N_16203);
xnor U21384 (N_21384,N_16119,N_17522);
nand U21385 (N_21385,N_19490,N_16986);
or U21386 (N_21386,N_15807,N_16287);
nand U21387 (N_21387,N_19231,N_19884);
xor U21388 (N_21388,N_19892,N_17912);
nor U21389 (N_21389,N_18413,N_16725);
nand U21390 (N_21390,N_16561,N_16360);
nor U21391 (N_21391,N_16890,N_18188);
nand U21392 (N_21392,N_19915,N_15471);
xor U21393 (N_21393,N_18573,N_15443);
nor U21394 (N_21394,N_17297,N_15444);
and U21395 (N_21395,N_17336,N_19899);
xnor U21396 (N_21396,N_17191,N_18775);
xnor U21397 (N_21397,N_17950,N_17922);
nor U21398 (N_21398,N_17720,N_16731);
nand U21399 (N_21399,N_18544,N_18519);
nor U21400 (N_21400,N_18029,N_16767);
nand U21401 (N_21401,N_19602,N_17268);
and U21402 (N_21402,N_19941,N_15854);
or U21403 (N_21403,N_17471,N_16008);
nand U21404 (N_21404,N_19792,N_16259);
and U21405 (N_21405,N_19604,N_15566);
or U21406 (N_21406,N_19070,N_19612);
or U21407 (N_21407,N_17987,N_17143);
nand U21408 (N_21408,N_19689,N_17884);
xnor U21409 (N_21409,N_16934,N_16428);
nand U21410 (N_21410,N_16447,N_16491);
nand U21411 (N_21411,N_18081,N_15098);
nor U21412 (N_21412,N_19972,N_19328);
and U21413 (N_21413,N_17657,N_19316);
nand U21414 (N_21414,N_19526,N_17598);
and U21415 (N_21415,N_15656,N_18946);
xor U21416 (N_21416,N_19282,N_19353);
xor U21417 (N_21417,N_18968,N_17960);
nand U21418 (N_21418,N_15018,N_16381);
nor U21419 (N_21419,N_15932,N_18232);
xor U21420 (N_21420,N_15232,N_19775);
and U21421 (N_21421,N_15580,N_16737);
or U21422 (N_21422,N_16696,N_19224);
nand U21423 (N_21423,N_17828,N_18730);
nand U21424 (N_21424,N_17609,N_16248);
and U21425 (N_21425,N_16628,N_18585);
or U21426 (N_21426,N_16073,N_15649);
nor U21427 (N_21427,N_18924,N_18843);
and U21428 (N_21428,N_16243,N_18890);
nor U21429 (N_21429,N_16420,N_18010);
xor U21430 (N_21430,N_16050,N_17220);
nor U21431 (N_21431,N_18023,N_17927);
nor U21432 (N_21432,N_19539,N_16742);
xor U21433 (N_21433,N_17791,N_18351);
and U21434 (N_21434,N_17848,N_16607);
xnor U21435 (N_21435,N_15167,N_19566);
nor U21436 (N_21436,N_16592,N_16198);
nor U21437 (N_21437,N_17015,N_16207);
or U21438 (N_21438,N_15615,N_17246);
nor U21439 (N_21439,N_16482,N_19510);
nor U21440 (N_21440,N_16012,N_18492);
and U21441 (N_21441,N_17063,N_16100);
or U21442 (N_21442,N_15407,N_19464);
nor U21443 (N_21443,N_19709,N_18225);
xnor U21444 (N_21444,N_16426,N_17249);
nand U21445 (N_21445,N_17929,N_17199);
xor U21446 (N_21446,N_18754,N_16214);
nand U21447 (N_21447,N_16122,N_19134);
xnor U21448 (N_21448,N_17729,N_18501);
nand U21449 (N_21449,N_17146,N_17179);
nor U21450 (N_21450,N_19639,N_19695);
and U21451 (N_21451,N_15591,N_17509);
nand U21452 (N_21452,N_15158,N_16376);
or U21453 (N_21453,N_15249,N_18429);
nor U21454 (N_21454,N_17260,N_17695);
nand U21455 (N_21455,N_16675,N_19402);
nand U21456 (N_21456,N_17441,N_16135);
nor U21457 (N_21457,N_15507,N_18441);
or U21458 (N_21458,N_17587,N_16400);
and U21459 (N_21459,N_18286,N_15340);
nand U21460 (N_21460,N_19790,N_16608);
xnor U21461 (N_21461,N_19934,N_19719);
nand U21462 (N_21462,N_15240,N_17830);
and U21463 (N_21463,N_15331,N_17771);
nand U21464 (N_21464,N_15682,N_19865);
nor U21465 (N_21465,N_19952,N_15101);
or U21466 (N_21466,N_19105,N_18945);
nor U21467 (N_21467,N_15237,N_16714);
nor U21468 (N_21468,N_18500,N_17803);
and U21469 (N_21469,N_16797,N_18530);
or U21470 (N_21470,N_17502,N_19270);
xnor U21471 (N_21471,N_16265,N_19723);
xor U21472 (N_21472,N_16270,N_17620);
xnor U21473 (N_21473,N_19725,N_19405);
xor U21474 (N_21474,N_16874,N_15324);
xor U21475 (N_21475,N_19601,N_16568);
nand U21476 (N_21476,N_16599,N_17461);
and U21477 (N_21477,N_18597,N_18325);
xnor U21478 (N_21478,N_16715,N_18576);
xnor U21479 (N_21479,N_15479,N_19385);
xor U21480 (N_21480,N_18785,N_18546);
xor U21481 (N_21481,N_15423,N_15354);
or U21482 (N_21482,N_18543,N_16864);
nand U21483 (N_21483,N_15374,N_15308);
nor U21484 (N_21484,N_17263,N_15382);
xnor U21485 (N_21485,N_18127,N_17037);
nor U21486 (N_21486,N_18391,N_16088);
or U21487 (N_21487,N_15285,N_15896);
nand U21488 (N_21488,N_16645,N_16979);
or U21489 (N_21489,N_18235,N_17849);
or U21490 (N_21490,N_15100,N_15642);
nor U21491 (N_21491,N_17321,N_18043);
nand U21492 (N_21492,N_17599,N_19691);
xnor U21493 (N_21493,N_19009,N_19536);
and U21494 (N_21494,N_17208,N_18678);
nor U21495 (N_21495,N_17890,N_19217);
nor U21496 (N_21496,N_18417,N_17579);
nor U21497 (N_21497,N_19621,N_18192);
xnor U21498 (N_21498,N_18524,N_18454);
or U21499 (N_21499,N_16315,N_16396);
nand U21500 (N_21500,N_18089,N_17901);
nor U21501 (N_21501,N_19069,N_18402);
or U21502 (N_21502,N_17487,N_19063);
xnor U21503 (N_21503,N_17784,N_15886);
xor U21504 (N_21504,N_16867,N_17373);
and U21505 (N_21505,N_18261,N_19120);
xor U21506 (N_21506,N_16782,N_18499);
or U21507 (N_21507,N_18400,N_15321);
and U21508 (N_21508,N_18711,N_15956);
or U21509 (N_21509,N_19918,N_19004);
or U21510 (N_21510,N_15714,N_15741);
and U21511 (N_21511,N_16472,N_15461);
nand U21512 (N_21512,N_16474,N_17700);
nor U21513 (N_21513,N_15826,N_19625);
xnor U21514 (N_21514,N_17406,N_19481);
or U21515 (N_21515,N_19859,N_15316);
and U21516 (N_21516,N_18330,N_18419);
nand U21517 (N_21517,N_17685,N_16852);
nor U21518 (N_21518,N_19387,N_16236);
and U21519 (N_21519,N_19335,N_18901);
nand U21520 (N_21520,N_15970,N_15268);
nor U21521 (N_21521,N_19617,N_15312);
and U21522 (N_21522,N_19514,N_17534);
xnor U21523 (N_21523,N_16750,N_18126);
nor U21524 (N_21524,N_15773,N_17407);
nand U21525 (N_21525,N_16102,N_16912);
or U21526 (N_21526,N_17661,N_17897);
or U21527 (N_21527,N_17718,N_18131);
xnor U21528 (N_21528,N_19914,N_15023);
nor U21529 (N_21529,N_17696,N_18397);
or U21530 (N_21530,N_19219,N_19216);
nor U21531 (N_21531,N_18651,N_18103);
or U21532 (N_21532,N_19014,N_16615);
xor U21533 (N_21533,N_17067,N_19508);
xnor U21534 (N_21534,N_19895,N_19588);
nand U21535 (N_21535,N_16141,N_15310);
and U21536 (N_21536,N_18687,N_15403);
and U21537 (N_21537,N_16196,N_18037);
and U21538 (N_21538,N_19074,N_17689);
and U21539 (N_21539,N_16485,N_19728);
nor U21540 (N_21540,N_17706,N_16255);
and U21541 (N_21541,N_15415,N_15064);
nand U21542 (N_21542,N_18159,N_15189);
xor U21543 (N_21543,N_16312,N_18449);
nand U21544 (N_21544,N_17988,N_15378);
or U21545 (N_21545,N_17232,N_19461);
or U21546 (N_21546,N_17895,N_16743);
xor U21547 (N_21547,N_19117,N_17542);
or U21548 (N_21548,N_17826,N_19675);
nand U21549 (N_21549,N_15091,N_19367);
nor U21550 (N_21550,N_15097,N_16683);
or U21551 (N_21551,N_18724,N_16068);
and U21552 (N_21552,N_16739,N_19060);
xor U21553 (N_21553,N_19410,N_16151);
nand U21554 (N_21554,N_19513,N_17916);
nand U21555 (N_21555,N_15483,N_18075);
nor U21556 (N_21556,N_19269,N_19382);
and U21557 (N_21557,N_17621,N_19690);
nand U21558 (N_21558,N_17701,N_15373);
xor U21559 (N_21559,N_17551,N_18963);
xnor U21560 (N_21560,N_19297,N_15364);
xor U21561 (N_21561,N_15627,N_19194);
nand U21562 (N_21562,N_17659,N_15636);
xor U21563 (N_21563,N_19426,N_17966);
xor U21564 (N_21564,N_19575,N_19502);
and U21565 (N_21565,N_18756,N_17352);
and U21566 (N_21566,N_18201,N_18662);
and U21567 (N_21567,N_18478,N_15873);
nand U21568 (N_21568,N_16302,N_17136);
xnor U21569 (N_21569,N_19998,N_17209);
and U21570 (N_21570,N_19488,N_17757);
nand U21571 (N_21571,N_16914,N_16435);
nor U21572 (N_21572,N_17115,N_18407);
or U21573 (N_21573,N_16394,N_19291);
xor U21574 (N_21574,N_17241,N_17470);
nor U21575 (N_21575,N_16066,N_16348);
or U21576 (N_21576,N_16023,N_15111);
nand U21577 (N_21577,N_18820,N_15569);
or U21578 (N_21578,N_16826,N_18796);
xor U21579 (N_21579,N_18939,N_17053);
or U21580 (N_21580,N_17926,N_16873);
nor U21581 (N_21581,N_18426,N_16555);
nor U21582 (N_21582,N_17668,N_16205);
and U21583 (N_21583,N_15817,N_16508);
nor U21584 (N_21584,N_15041,N_15005);
and U21585 (N_21585,N_15317,N_19767);
nand U21586 (N_21586,N_19295,N_19404);
xnor U21587 (N_21587,N_18512,N_19179);
and U21588 (N_21588,N_17637,N_19417);
xor U21589 (N_21589,N_16744,N_19397);
nand U21590 (N_21590,N_15211,N_15849);
nor U21591 (N_21591,N_19082,N_19186);
xor U21592 (N_21592,N_17965,N_16488);
nand U21593 (N_21593,N_15552,N_18643);
and U21594 (N_21594,N_16793,N_15309);
and U21595 (N_21595,N_19418,N_15476);
or U21596 (N_21596,N_18810,N_15541);
nor U21597 (N_21597,N_15713,N_15594);
xor U21598 (N_21598,N_15547,N_17697);
and U21599 (N_21599,N_15601,N_18617);
or U21600 (N_21600,N_19765,N_15204);
and U21601 (N_21601,N_19888,N_19177);
xnor U21602 (N_21602,N_16833,N_16429);
or U21603 (N_21603,N_17486,N_15678);
and U21604 (N_21604,N_18299,N_15523);
nor U21605 (N_21605,N_17202,N_15160);
nor U21606 (N_21606,N_15774,N_16199);
nand U21607 (N_21607,N_16804,N_15539);
xnor U21608 (N_21608,N_18631,N_16785);
nand U21609 (N_21609,N_18904,N_15217);
xnor U21610 (N_21610,N_18349,N_17449);
or U21611 (N_21611,N_18934,N_17827);
nand U21612 (N_21612,N_19151,N_19801);
xor U21613 (N_21613,N_17740,N_16956);
or U21614 (N_21614,N_16699,N_16954);
nor U21615 (N_21615,N_19869,N_15532);
or U21616 (N_21616,N_19633,N_15974);
nand U21617 (N_21617,N_18058,N_15116);
xor U21618 (N_21618,N_17001,N_18008);
or U21619 (N_21619,N_16654,N_15170);
and U21620 (N_21620,N_15819,N_19655);
nor U21621 (N_21621,N_19678,N_17553);
xor U21622 (N_21622,N_17525,N_18927);
xor U21623 (N_21623,N_18586,N_18950);
xor U21624 (N_21624,N_16536,N_17475);
nor U21625 (N_21625,N_15173,N_15371);
or U21626 (N_21626,N_16036,N_17687);
and U21627 (N_21627,N_19025,N_18471);
nand U21628 (N_21628,N_18991,N_15490);
xor U21629 (N_21629,N_15104,N_16780);
nand U21630 (N_21630,N_18013,N_15043);
nor U21631 (N_21631,N_17623,N_19359);
and U21632 (N_21632,N_19598,N_15085);
and U21633 (N_21633,N_17221,N_15786);
xnor U21634 (N_21634,N_15746,N_17244);
and U21635 (N_21635,N_15944,N_18329);
or U21636 (N_21636,N_15764,N_19265);
and U21637 (N_21637,N_19128,N_15291);
nand U21638 (N_21638,N_19336,N_19903);
and U21639 (N_21639,N_15270,N_15393);
or U21640 (N_21640,N_15689,N_18537);
and U21641 (N_21641,N_17210,N_19283);
or U21642 (N_21642,N_18326,N_15370);
nand U21643 (N_21643,N_19034,N_18955);
nand U21644 (N_21644,N_19738,N_16280);
or U21645 (N_21645,N_17864,N_18606);
xnor U21646 (N_21646,N_15667,N_16108);
nand U21647 (N_21647,N_19334,N_19850);
nor U21648 (N_21648,N_17284,N_19732);
nand U21649 (N_21649,N_16732,N_18497);
nand U21650 (N_21650,N_15298,N_15059);
nor U21651 (N_21651,N_18028,N_18958);
and U21652 (N_21652,N_18905,N_15502);
xnor U21653 (N_21653,N_18226,N_16685);
xnor U21654 (N_21654,N_16355,N_17196);
nand U21655 (N_21655,N_17164,N_18140);
nand U21656 (N_21656,N_18310,N_16532);
or U21657 (N_21657,N_19215,N_18892);
nand U21658 (N_21658,N_16671,N_18153);
nand U21659 (N_21659,N_19715,N_16902);
and U21660 (N_21660,N_19314,N_19271);
or U21661 (N_21661,N_19486,N_19537);
nor U21662 (N_21662,N_17654,N_16713);
nand U21663 (N_21663,N_18222,N_17674);
and U21664 (N_21664,N_15660,N_19172);
nor U21665 (N_21665,N_15273,N_19213);
nor U21666 (N_21666,N_16475,N_17230);
nor U21667 (N_21667,N_19155,N_17386);
nand U21668 (N_21668,N_19377,N_19279);
or U21669 (N_21669,N_15394,N_19997);
xnor U21670 (N_21670,N_15176,N_17102);
or U21671 (N_21671,N_17000,N_17780);
nand U21672 (N_21672,N_15432,N_15669);
nand U21673 (N_21673,N_15710,N_17222);
and U21674 (N_21674,N_19293,N_15964);
xor U21675 (N_21675,N_17887,N_18470);
nand U21676 (N_21676,N_15352,N_18003);
nand U21677 (N_21677,N_16172,N_19124);
xnor U21678 (N_21678,N_16579,N_18014);
nor U21679 (N_21679,N_16492,N_16262);
and U21680 (N_21680,N_17310,N_17327);
xor U21681 (N_21681,N_16168,N_16087);
xor U21682 (N_21682,N_15700,N_18251);
xnor U21683 (N_21683,N_18422,N_19107);
and U21684 (N_21684,N_17574,N_17704);
and U21685 (N_21685,N_16929,N_18302);
xor U21686 (N_21686,N_17480,N_19643);
and U21687 (N_21687,N_15090,N_15000);
xor U21688 (N_21688,N_17698,N_16238);
nand U21689 (N_21689,N_17947,N_18211);
nor U21690 (N_21690,N_15687,N_17012);
or U21691 (N_21691,N_17630,N_15534);
xnor U21692 (N_21692,N_16370,N_17213);
or U21693 (N_21693,N_15958,N_18090);
and U21694 (N_21694,N_16039,N_17858);
nor U21695 (N_21695,N_16240,N_15659);
nand U21696 (N_21696,N_19755,N_18932);
nand U21697 (N_21697,N_18714,N_16016);
and U21698 (N_21698,N_16808,N_19798);
nand U21699 (N_21699,N_19887,N_18248);
or U21700 (N_21700,N_17346,N_19497);
or U21701 (N_21701,N_17073,N_16865);
or U21702 (N_21702,N_15279,N_16617);
nor U21703 (N_21703,N_15343,N_16943);
or U21704 (N_21704,N_16915,N_15172);
nor U21705 (N_21705,N_18420,N_15827);
nand U21706 (N_21706,N_16911,N_19059);
xnor U21707 (N_21707,N_19463,N_19473);
nor U21708 (N_21708,N_16880,N_15353);
nor U21709 (N_21709,N_15789,N_18751);
and U21710 (N_21710,N_17388,N_17003);
nor U21711 (N_21711,N_15839,N_18702);
or U21712 (N_21712,N_19558,N_18642);
nand U21713 (N_21713,N_18560,N_18390);
xnor U21714 (N_21714,N_18119,N_18387);
or U21715 (N_21715,N_15790,N_16444);
and U21716 (N_21716,N_17465,N_19718);
nand U21717 (N_21717,N_17921,N_19636);
or U21718 (N_21718,N_17852,N_19370);
nor U21719 (N_21719,N_17030,N_19073);
and U21720 (N_21720,N_15142,N_18887);
xnor U21721 (N_21721,N_19465,N_19469);
and U21722 (N_21722,N_17035,N_17452);
or U21723 (N_21723,N_16719,N_15830);
nor U21724 (N_21724,N_19960,N_16583);
or U21725 (N_21725,N_17057,N_16504);
xnor U21726 (N_21726,N_15850,N_16154);
and U21727 (N_21727,N_16453,N_19045);
nor U21728 (N_21728,N_19447,N_15553);
nand U21729 (N_21729,N_17294,N_18667);
nor U21730 (N_21730,N_18717,N_19197);
nor U21731 (N_21731,N_16998,N_18834);
and U21732 (N_21732,N_19420,N_15987);
nand U21733 (N_21733,N_15351,N_19046);
or U21734 (N_21734,N_18998,N_19847);
and U21735 (N_21735,N_17192,N_16442);
nor U21736 (N_21736,N_18800,N_18355);
and U21737 (N_21737,N_19272,N_17253);
nand U21738 (N_21738,N_18490,N_16841);
xor U21739 (N_21739,N_19981,N_16668);
and U21740 (N_21740,N_15010,N_18734);
nor U21741 (N_21741,N_17250,N_15554);
nor U21742 (N_21742,N_16260,N_16957);
and U21743 (N_21743,N_18669,N_16703);
and U21744 (N_21744,N_17915,N_19556);
xor U21745 (N_21745,N_19361,N_19096);
nor U21746 (N_21746,N_18093,N_18589);
or U21747 (N_21747,N_19823,N_17218);
or U21748 (N_21748,N_16024,N_15166);
xnor U21749 (N_21749,N_17472,N_19191);
and U21750 (N_21750,N_19928,N_18460);
xnor U21751 (N_21751,N_18236,N_16757);
nand U21752 (N_21752,N_17549,N_17821);
or U21753 (N_21753,N_19794,N_19344);
and U21754 (N_21754,N_18077,N_15470);
nor U21755 (N_21755,N_19883,N_18107);
xor U21756 (N_21756,N_19839,N_15081);
nor U21757 (N_21757,N_17120,N_16115);
or U21758 (N_21758,N_16839,N_15676);
and U21759 (N_21759,N_15564,N_18245);
xor U21760 (N_21760,N_16495,N_17083);
and U21761 (N_21761,N_19205,N_18439);
nor U21762 (N_21762,N_16591,N_15148);
and U21763 (N_21763,N_18345,N_17526);
or U21764 (N_21764,N_19471,N_16388);
xnor U21765 (N_21765,N_19201,N_16144);
nor U21766 (N_21766,N_16439,N_16464);
nor U21767 (N_21767,N_19064,N_18151);
xnor U21768 (N_21768,N_15941,N_16680);
and U21769 (N_21769,N_16031,N_17233);
nand U21770 (N_21770,N_17676,N_17317);
or U21771 (N_21771,N_19929,N_16296);
nor U21772 (N_21772,N_17307,N_18564);
xnor U21773 (N_21773,N_16471,N_16116);
or U21774 (N_21774,N_16518,N_19300);
nand U21775 (N_21775,N_17794,N_18867);
xnor U21776 (N_21776,N_17933,N_16231);
or U21777 (N_21777,N_17205,N_19232);
and U21778 (N_21778,N_15792,N_15401);
and U21779 (N_21779,N_19520,N_15006);
xnor U21780 (N_21780,N_15073,N_17521);
nor U21781 (N_21781,N_17602,N_19012);
nand U21782 (N_21782,N_18213,N_15915);
nor U21783 (N_21783,N_17429,N_17801);
nand U21784 (N_21784,N_16459,N_16647);
nor U21785 (N_21785,N_17129,N_18548);
or U21786 (N_21786,N_19999,N_18481);
or U21787 (N_21787,N_19975,N_18317);
or U21788 (N_21788,N_18434,N_18034);
nor U21789 (N_21789,N_17198,N_18321);
nor U21790 (N_21790,N_15548,N_18870);
nand U21791 (N_21791,N_16316,N_18120);
or U21792 (N_21792,N_16771,N_18723);
nor U21793 (N_21793,N_15163,N_19390);
xor U21794 (N_21794,N_17962,N_18811);
nor U21795 (N_21795,N_18338,N_15525);
nor U21796 (N_21796,N_17861,N_16974);
and U21797 (N_21797,N_15560,N_15315);
nor U21798 (N_21798,N_18173,N_16578);
and U21799 (N_21799,N_16365,N_17467);
or U21800 (N_21800,N_17466,N_15412);
or U21801 (N_21801,N_16894,N_16308);
and U21802 (N_21802,N_15862,N_16624);
xnor U21803 (N_21803,N_17959,N_16700);
nand U21804 (N_21804,N_19257,N_18686);
and U21805 (N_21805,N_19967,N_17512);
nand U21806 (N_21806,N_16997,N_15213);
and U21807 (N_21807,N_18936,N_17535);
xor U21808 (N_21808,N_16150,N_19241);
nand U21809 (N_21809,N_15110,N_19384);
or U21810 (N_21810,N_19577,N_17313);
nor U21811 (N_21811,N_19931,N_17724);
or U21812 (N_21812,N_15671,N_17932);
xnor U21813 (N_21813,N_17815,N_17954);
or U21814 (N_21814,N_19944,N_19716);
xor U21815 (N_21815,N_16157,N_18049);
and U21816 (N_21816,N_16017,N_15397);
xnor U21817 (N_21817,N_16822,N_15520);
nor U21818 (N_21818,N_17248,N_18851);
nor U21819 (N_21819,N_16577,N_16284);
and U21820 (N_21820,N_15770,N_18816);
and U21821 (N_21821,N_15445,N_19484);
or U21822 (N_21822,N_18943,N_15975);
xnor U21823 (N_21823,N_17435,N_16142);
xnor U21824 (N_21824,N_19187,N_19911);
or U21825 (N_21825,N_19318,N_15140);
nand U21826 (N_21826,N_19084,N_16679);
nor U21827 (N_21827,N_17071,N_16246);
xor U21828 (N_21828,N_16729,N_19582);
xor U21829 (N_21829,N_18108,N_19871);
and U21830 (N_21830,N_17888,N_18294);
and U21831 (N_21831,N_15359,N_18242);
xor U21832 (N_21832,N_15003,N_15185);
nand U21833 (N_21833,N_19947,N_16384);
nand U21834 (N_21834,N_19442,N_18974);
or U21835 (N_21835,N_15485,N_18593);
and U21836 (N_21836,N_17812,N_16350);
or U21837 (N_21837,N_19614,N_17356);
or U21838 (N_21838,N_17107,N_17123);
nor U21839 (N_21839,N_18648,N_18128);
xor U21840 (N_21840,N_18280,N_17633);
and U21841 (N_21841,N_18542,N_17746);
and U21842 (N_21842,N_17879,N_15938);
nor U21843 (N_21843,N_17504,N_16325);
xnor U21844 (N_21844,N_16697,N_17683);
or U21845 (N_21845,N_17995,N_17684);
xnor U21846 (N_21846,N_16631,N_15045);
xnor U21847 (N_21847,N_17392,N_15495);
nand U21848 (N_21848,N_17068,N_15570);
nand U21849 (N_21849,N_18933,N_16994);
and U21850 (N_21850,N_18753,N_17019);
nand U21851 (N_21851,N_19677,N_17377);
xor U21852 (N_21852,N_18575,N_16228);
or U21853 (N_21853,N_17896,N_17194);
nor U21854 (N_21854,N_18383,N_15782);
or U21855 (N_21855,N_18559,N_18795);
and U21856 (N_21856,N_17836,N_15583);
nand U21857 (N_21857,N_19324,N_17274);
nand U21858 (N_21858,N_16918,N_16282);
xor U21859 (N_21859,N_19093,N_17070);
or U21860 (N_21860,N_15349,N_18000);
nand U21861 (N_21861,N_15951,N_16523);
xnor U21862 (N_21862,N_17638,N_18047);
xor U21863 (N_21863,N_16548,N_17148);
nor U21864 (N_21864,N_17808,N_16446);
nand U21865 (N_21865,N_16846,N_17318);
or U21866 (N_21866,N_17909,N_15294);
nor U21867 (N_21867,N_18182,N_15563);
and U21868 (N_21868,N_15625,N_16229);
and U21869 (N_21869,N_17483,N_15203);
xor U21870 (N_21870,N_18364,N_16761);
and U21871 (N_21871,N_15319,N_19489);
nand U21872 (N_21872,N_16818,N_16563);
or U21873 (N_21873,N_15736,N_18929);
and U21874 (N_21874,N_17537,N_18908);
or U21875 (N_21875,N_15210,N_15425);
xor U21876 (N_21876,N_19671,N_16515);
nand U21877 (N_21877,N_17335,N_19101);
xnor U21878 (N_21878,N_18859,N_17285);
and U21879 (N_21879,N_16091,N_18980);
and U21880 (N_21880,N_16098,N_17324);
nor U21881 (N_21881,N_16944,N_19571);
nand U21882 (N_21882,N_15921,N_19572);
nor U21883 (N_21883,N_19395,N_19674);
and U21884 (N_21884,N_19409,N_19615);
xnor U21885 (N_21885,N_17520,N_15247);
or U21886 (N_21886,N_16455,N_18178);
nor U21887 (N_21887,N_17814,N_18069);
nand U21888 (N_21888,N_16473,N_16898);
nand U21889 (N_21889,N_17494,N_16848);
and U21890 (N_21890,N_16658,N_19466);
nand U21891 (N_21891,N_18473,N_19424);
or U21892 (N_21892,N_15588,N_16601);
nor U21893 (N_21893,N_19472,N_18879);
and U21894 (N_21894,N_18578,N_15661);
nor U21895 (N_21895,N_18279,N_16237);
nand U21896 (N_21896,N_17850,N_17326);
nand U21897 (N_21897,N_17914,N_16910);
and U21898 (N_21898,N_16790,N_18855);
nor U21899 (N_21899,N_15813,N_15939);
nand U21900 (N_21900,N_15772,N_17772);
xor U21901 (N_21901,N_16107,N_16253);
nand U21902 (N_21902,N_18570,N_18748);
nor U21903 (N_21903,N_15866,N_17501);
nor U21904 (N_21904,N_18005,N_17712);
and U21905 (N_21905,N_18665,N_17004);
nor U21906 (N_21906,N_15472,N_19797);
nor U21907 (N_21907,N_19453,N_18274);
and U21908 (N_21908,N_17728,N_19220);
and U21909 (N_21909,N_16558,N_17601);
and U21910 (N_21910,N_15055,N_16354);
xnor U21911 (N_21911,N_18882,N_15629);
nor U21912 (N_21912,N_15405,N_16674);
nand U21913 (N_21913,N_17873,N_15496);
or U21914 (N_21914,N_19896,N_16948);
or U21915 (N_21915,N_18100,N_17469);
nand U21916 (N_21916,N_17431,N_17840);
nand U21917 (N_21917,N_16514,N_17790);
and U21918 (N_21918,N_16831,N_17945);
nand U21919 (N_21919,N_15631,N_19729);
xor U21920 (N_21920,N_18682,N_16025);
xor U21921 (N_21921,N_16557,N_18368);
and U21922 (N_21922,N_17788,N_15390);
or U21923 (N_21923,N_15848,N_19415);
or U21924 (N_21924,N_18591,N_18607);
nor U21925 (N_21925,N_16888,N_15535);
or U21926 (N_21926,N_15296,N_18603);
xor U21927 (N_21927,N_15347,N_15756);
xnor U21928 (N_21928,N_15997,N_18065);
xnor U21929 (N_21929,N_18857,N_15662);
nor U21930 (N_21930,N_15711,N_16278);
xnor U21931 (N_21931,N_15031,N_19432);
nor U21932 (N_21932,N_19171,N_15701);
and U21933 (N_21933,N_18925,N_15265);
and U21934 (N_21934,N_19548,N_15260);
xor U21935 (N_21935,N_16844,N_19443);
nor U21936 (N_21936,N_18032,N_16616);
xnor U21937 (N_21937,N_18040,N_18863);
nand U21938 (N_21938,N_18677,N_17174);
nor U21939 (N_21939,N_16165,N_16200);
nor U21940 (N_21940,N_19408,N_19477);
nor U21941 (N_21941,N_17610,N_18804);
xor U21942 (N_21942,N_18359,N_16886);
xnor U21943 (N_21943,N_19094,N_16009);
nand U21944 (N_21944,N_16832,N_15953);
or U21945 (N_21945,N_15030,N_15576);
nand U21946 (N_21946,N_18765,N_19841);
xor U21947 (N_21947,N_16089,N_15383);
nor U21948 (N_21948,N_19819,N_19044);
or U21949 (N_21949,N_16547,N_15271);
or U21950 (N_21950,N_16823,N_15058);
nand U21951 (N_21951,N_19104,N_16932);
and U21952 (N_21952,N_19337,N_15048);
nor U21953 (N_21953,N_15231,N_19784);
xor U21954 (N_21954,N_16784,N_16056);
nor U21955 (N_21955,N_18432,N_16594);
xor U21956 (N_21956,N_19332,N_18442);
nand U21957 (N_21957,N_19984,N_16160);
nor U21958 (N_21958,N_18990,N_16212);
xnor U21959 (N_21959,N_17289,N_16342);
and U21960 (N_21960,N_17223,N_16572);
xnor U21961 (N_21961,N_16046,N_19699);
or U21962 (N_21962,N_15105,N_15519);
nor U21963 (N_21963,N_15734,N_18818);
nand U21964 (N_21964,N_18553,N_15996);
and U21965 (N_21965,N_19373,N_17396);
and U21966 (N_21966,N_19195,N_19047);
and U21967 (N_21967,N_15976,N_16602);
xnor U21968 (N_21968,N_16393,N_17973);
nand U21969 (N_21969,N_17672,N_15843);
nand U21970 (N_21970,N_17902,N_19185);
nand U21971 (N_21971,N_18137,N_15531);
xor U21972 (N_21972,N_17036,N_15880);
nor U21973 (N_21973,N_15910,N_16389);
nand U21974 (N_21974,N_18670,N_17725);
xor U21975 (N_21975,N_17832,N_17119);
and U21976 (N_21976,N_18174,N_17214);
and U21977 (N_21977,N_18520,N_16149);
and U21978 (N_21978,N_18085,N_18237);
nand U21979 (N_21979,N_17224,N_16392);
xnor U21980 (N_21980,N_17538,N_15050);
and U21981 (N_21981,N_17280,N_17975);
nand U21982 (N_21982,N_17645,N_18874);
xor U21983 (N_21983,N_19018,N_15369);
nor U21984 (N_21984,N_15643,N_19169);
nand U21985 (N_21985,N_15215,N_18674);
nand U21986 (N_21986,N_17300,N_19787);
nand U21987 (N_21987,N_17152,N_16129);
and U21988 (N_21988,N_15306,N_16881);
nor U21989 (N_21989,N_19993,N_16095);
and U21990 (N_21990,N_16317,N_18447);
or U21991 (N_21991,N_15806,N_18777);
or U21992 (N_21992,N_15762,N_15420);
nor U21993 (N_21993,N_18825,N_17918);
nand U21994 (N_21994,N_18239,N_17303);
and U21995 (N_21995,N_17454,N_16987);
or U21996 (N_21996,N_18405,N_15516);
nand U21997 (N_21997,N_19534,N_16218);
xnor U21998 (N_21998,N_16059,N_16856);
nor U21999 (N_21999,N_17168,N_15198);
or U22000 (N_22000,N_17055,N_19950);
nor U22001 (N_22001,N_18253,N_16877);
or U22002 (N_22002,N_17195,N_16613);
or U22003 (N_22003,N_18132,N_16884);
nand U22004 (N_22004,N_17344,N_18324);
xnor U22005 (N_22005,N_17776,N_15961);
or U22006 (N_22006,N_15029,N_18233);
nor U22007 (N_22007,N_16630,N_18583);
or U22008 (N_22008,N_17137,N_18817);
and U22009 (N_22009,N_19022,N_19400);
and U22010 (N_22010,N_15277,N_15474);
and U22011 (N_22011,N_16519,N_16774);
xnor U22012 (N_22012,N_15112,N_16015);
nand U22013 (N_22013,N_16740,N_16064);
nand U22014 (N_22014,N_18031,N_17726);
xnor U22015 (N_22015,N_18092,N_17928);
or U22016 (N_22016,N_17367,N_16406);
nand U22017 (N_22017,N_15878,N_19111);
and U22018 (N_22018,N_16343,N_19567);
xnor U22019 (N_22019,N_18307,N_15368);
nand U22020 (N_22020,N_15463,N_15024);
nor U22021 (N_22021,N_16835,N_15219);
nor U22022 (N_22022,N_18308,N_17906);
or U22023 (N_22023,N_17842,N_16045);
xnor U22024 (N_22024,N_15995,N_15769);
xor U22025 (N_22025,N_19909,N_18721);
nand U22026 (N_22026,N_19552,N_17382);
or U22027 (N_22027,N_15982,N_18228);
and U22028 (N_22028,N_17380,N_19436);
nor U22029 (N_22029,N_15372,N_16875);
xnor U22030 (N_22030,N_15624,N_19829);
nand U22031 (N_22031,N_15481,N_17711);
or U22032 (N_22032,N_19401,N_18176);
or U22033 (N_22033,N_19414,N_17111);
nand U22034 (N_22034,N_18300,N_19118);
nand U22035 (N_22035,N_18931,N_15940);
nand U22036 (N_22036,N_15411,N_19623);
xor U22037 (N_22037,N_17495,N_17031);
or U22038 (N_22038,N_16053,N_17783);
and U22039 (N_22039,N_15092,N_16963);
nor U22040 (N_22040,N_18525,N_15155);
or U22041 (N_22041,N_18657,N_18011);
or U22042 (N_22042,N_16753,N_18059);
nand U22043 (N_22043,N_17930,N_19180);
or U22044 (N_22044,N_18479,N_18808);
xnor U22045 (N_22045,N_18435,N_17604);
and U22046 (N_22046,N_17680,N_15755);
or U22047 (N_22047,N_16431,N_18264);
nor U22048 (N_22048,N_19341,N_15984);
nand U22049 (N_22049,N_19256,N_18510);
nor U22050 (N_22050,N_18468,N_18858);
nor U22051 (N_22051,N_16215,N_17829);
xor U22052 (N_22052,N_17024,N_17323);
xor U22053 (N_22053,N_16076,N_17421);
nor U22054 (N_22054,N_17255,N_19178);
nor U22055 (N_22055,N_19821,N_15524);
and U22056 (N_22056,N_15327,N_16462);
or U22057 (N_22057,N_18366,N_15988);
xnor U22058 (N_22058,N_15118,N_15635);
xor U22059 (N_22059,N_15765,N_16456);
and U22060 (N_22060,N_18755,N_18467);
nor U22061 (N_22061,N_16876,N_17368);
nand U22062 (N_22062,N_18423,N_18186);
and U22063 (N_22063,N_18263,N_15834);
nand U22064 (N_22064,N_17234,N_18502);
xor U22065 (N_22065,N_15943,N_19434);
and U22066 (N_22066,N_19533,N_18050);
or U22067 (N_22067,N_19110,N_16411);
nor U22068 (N_22068,N_16922,N_18878);
nor U22069 (N_22069,N_18403,N_19438);
nand U22070 (N_22070,N_19676,N_17822);
or U22071 (N_22071,N_19982,N_15292);
nand U22072 (N_22072,N_15706,N_16387);
xor U22073 (N_22073,N_19875,N_16885);
nand U22074 (N_22074,N_18376,N_18703);
and U22075 (N_22075,N_16935,N_16821);
or U22076 (N_22076,N_18906,N_19017);
xor U22077 (N_22077,N_15712,N_16738);
nor U22078 (N_22078,N_19557,N_18815);
xor U22079 (N_22079,N_19855,N_16013);
or U22080 (N_22080,N_19002,N_19686);
or U22081 (N_22081,N_16224,N_19091);
or U22082 (N_22082,N_19173,N_18577);
nor U22083 (N_22083,N_19363,N_16417);
xnor U22084 (N_22084,N_17054,N_17650);
nor U22085 (N_22085,N_17719,N_17456);
nand U22086 (N_22086,N_17688,N_15069);
or U22087 (N_22087,N_15536,N_16227);
xor U22088 (N_22088,N_16020,N_16916);
xnor U22089 (N_22089,N_16340,N_16295);
nand U22090 (N_22090,N_17715,N_17588);
nand U22091 (N_22091,N_16976,N_19748);
or U22092 (N_22092,N_18571,N_18685);
nand U22093 (N_22093,N_17963,N_15107);
nand U22094 (N_22094,N_19726,N_17272);
and U22095 (N_22095,N_18276,N_15337);
nand U22096 (N_22096,N_19240,N_19394);
nand U22097 (N_22097,N_18790,N_19541);
xnor U22098 (N_22098,N_17655,N_15983);
nor U22099 (N_22099,N_17013,N_17989);
nand U22100 (N_22100,N_17340,N_16754);
and U22101 (N_22101,N_18844,N_16896);
and U22102 (N_22102,N_18408,N_15989);
xor U22103 (N_22103,N_18118,N_16026);
xor U22104 (N_22104,N_19003,N_19449);
nand U22105 (N_22105,N_15131,N_19450);
nor U22106 (N_22106,N_15533,N_16930);
nand U22107 (N_22107,N_18396,N_17341);
and U22108 (N_22108,N_18165,N_15657);
nand U22109 (N_22109,N_19953,N_18695);
nor U22110 (N_22110,N_19890,N_17446);
and U22111 (N_22111,N_15329,N_15981);
xor U22112 (N_22112,N_16972,N_15145);
or U22113 (N_22113,N_18221,N_18375);
xor U22114 (N_22114,N_18609,N_17319);
xnor U22115 (N_22115,N_17101,N_16175);
nor U22116 (N_22116,N_16587,N_18726);
nand U22117 (N_22117,N_18219,N_19818);
or U22118 (N_22118,N_16004,N_16989);
and U22119 (N_22119,N_17376,N_15966);
nor U22120 (N_22120,N_19518,N_15480);
nand U22121 (N_22121,N_19806,N_18821);
nand U22122 (N_22122,N_17080,N_17792);
xnor U22123 (N_22123,N_16191,N_15835);
nor U22124 (N_22124,N_17039,N_15034);
or U22125 (N_22125,N_17979,N_17892);
nor U22126 (N_22126,N_18112,N_16776);
nand U22127 (N_22127,N_15823,N_17231);
nor U22128 (N_22128,N_18275,N_19724);
nand U22129 (N_22129,N_18343,N_17817);
and U22130 (N_22130,N_15253,N_16309);
nor U22131 (N_22131,N_19338,N_19152);
xnor U22132 (N_22132,N_17351,N_18580);
nor U22133 (N_22133,N_18380,N_17008);
nor U22134 (N_22134,N_16327,N_16872);
nor U22135 (N_22135,N_15348,N_17669);
or U22136 (N_22136,N_15680,N_18044);
or U22137 (N_22137,N_16401,N_16415);
xor U22138 (N_22138,N_17984,N_16980);
or U22139 (N_22139,N_16909,N_16283);
and U22140 (N_22140,N_18161,N_19576);
and U22141 (N_22141,N_19731,N_17747);
or U22142 (N_22142,N_17007,N_17252);
nor U22143 (N_22143,N_16402,N_15326);
and U22144 (N_22144,N_18989,N_19852);
and U22145 (N_22145,N_15864,N_15389);
and U22146 (N_22146,N_17476,N_15937);
and U22147 (N_22147,N_19927,N_16705);
xor U22148 (N_22148,N_15455,N_17576);
xnor U22149 (N_22149,N_18314,N_18181);
nand U22150 (N_22150,N_18949,N_18109);
or U22151 (N_22151,N_15551,N_19276);
nand U22152 (N_22152,N_18461,N_19989);
or U22153 (N_22153,N_18860,N_17203);
nand U22154 (N_22154,N_19099,N_17634);
nor U22155 (N_22155,N_16672,N_18872);
and U22156 (N_22156,N_17140,N_17417);
xnor U22157 (N_22157,N_16498,N_17519);
or U22158 (N_22158,N_17564,N_15254);
xnor U22159 (N_22159,N_15926,N_15422);
xnor U22160 (N_22160,N_15255,N_19791);
xnor U22161 (N_22161,N_16079,N_15139);
xor U22162 (N_22162,N_19644,N_15021);
nand U22163 (N_22163,N_19956,N_15677);
nand U22164 (N_22164,N_18555,N_16162);
or U22165 (N_22165,N_19511,N_19161);
nor U22166 (N_22166,N_18599,N_15722);
or U22167 (N_22167,N_16298,N_18438);
or U22168 (N_22168,N_19917,N_18743);
and U22169 (N_22169,N_17778,N_16582);
or U22170 (N_22170,N_15207,N_17283);
and U22171 (N_22171,N_18138,N_15230);
nand U22172 (N_22172,N_17675,N_16825);
nand U22173 (N_22173,N_16477,N_19108);
nor U22174 (N_22174,N_19183,N_15808);
nand U22175 (N_22175,N_16208,N_16840);
and U22176 (N_22176,N_17113,N_15993);
nand U22177 (N_22177,N_19207,N_15068);
and U22178 (N_22178,N_15406,N_19713);
nor U22179 (N_22179,N_16450,N_17773);
nand U22180 (N_22180,N_17389,N_19157);
xor U22181 (N_22181,N_19259,N_17309);
or U22182 (N_22182,N_18806,N_19763);
or U22183 (N_22183,N_15360,N_19872);
and U22184 (N_22184,N_19066,N_18680);
and U22185 (N_22185,N_16382,N_15379);
xor U22186 (N_22186,N_19638,N_19029);
xor U22187 (N_22187,N_15256,N_16573);
nand U22188 (N_22188,N_16828,N_16058);
or U22189 (N_22189,N_17761,N_18584);
or U22190 (N_22190,N_16463,N_15751);
or U22191 (N_22191,N_17590,N_17575);
xnor U22192 (N_22192,N_17546,N_19322);
nor U22193 (N_22193,N_19844,N_16836);
and U22194 (N_22194,N_18474,N_19001);
or U22195 (N_22195,N_16919,N_17978);
and U22196 (N_22196,N_19524,N_18563);
or U22197 (N_22197,N_18865,N_15884);
or U22198 (N_22198,N_16486,N_15194);
or U22199 (N_22199,N_17112,N_19085);
or U22200 (N_22200,N_18386,N_15592);
xnor U22201 (N_22201,N_18649,N_16765);
and U22202 (N_22202,N_15433,N_19380);
xnor U22203 (N_22203,N_19570,N_15801);
xor U22204 (N_22204,N_16933,N_16460);
and U22205 (N_22205,N_17173,N_16820);
nand U22206 (N_22206,N_16544,N_19861);
xor U22207 (N_22207,N_19706,N_16502);
or U22208 (N_22208,N_15663,N_17951);
nand U22209 (N_22209,N_18446,N_15182);
xnor U22210 (N_22210,N_17492,N_18270);
xor U22211 (N_22211,N_19176,N_18758);
nand U22212 (N_22212,N_15451,N_17642);
and U22213 (N_22213,N_19812,N_17543);
xnor U22214 (N_22214,N_16373,N_17157);
xor U22215 (N_22215,N_19752,N_17237);
and U22216 (N_22216,N_16595,N_19352);
nor U22217 (N_22217,N_16610,N_18189);
xnor U22218 (N_22218,N_15089,N_18341);
xnor U22219 (N_22219,N_15928,N_16752);
or U22220 (N_22220,N_19889,N_16294);
and U22221 (N_22221,N_15999,N_17539);
xor U22222 (N_22222,N_15413,N_18658);
xor U22223 (N_22223,N_17156,N_15448);
nand U22224 (N_22224,N_15168,N_16537);
nand U22225 (N_22225,N_16146,N_15473);
and U22226 (N_22226,N_19712,N_15865);
nor U22227 (N_22227,N_19846,N_16210);
xor U22228 (N_22228,N_17860,N_15179);
or U22229 (N_22229,N_17425,N_16773);
nand U22230 (N_22230,N_17078,N_17002);
nor U22231 (N_22231,N_18428,N_17058);
nor U22232 (N_22232,N_19364,N_15288);
xor U22233 (N_22233,N_15143,N_15357);
or U22234 (N_22234,N_17239,N_19234);
or U22235 (N_22235,N_19422,N_17562);
xor U22236 (N_22236,N_16609,N_17981);
or U22237 (N_22237,N_16279,N_19594);
xnor U22238 (N_22238,N_18415,N_16496);
nand U22239 (N_22239,N_16217,N_15861);
xnor U22240 (N_22240,N_17748,N_19697);
nor U22241 (N_22241,N_16318,N_16101);
nand U22242 (N_22242,N_16289,N_16109);
nor U22243 (N_22243,N_17862,N_15505);
nand U22244 (N_22244,N_18262,N_17021);
and U22245 (N_22245,N_19916,N_16333);
or U22246 (N_22246,N_16140,N_15146);
xnor U22247 (N_22247,N_19563,N_19663);
or U22248 (N_22248,N_16673,N_16984);
nor U22249 (N_22249,N_19922,N_16249);
xnor U22250 (N_22250,N_15768,N_17511);
xor U22251 (N_22251,N_15908,N_16635);
xor U22252 (N_22252,N_17939,N_18552);
and U22253 (N_22253,N_19670,N_19355);
xnor U22254 (N_22254,N_18352,N_15567);
xnor U22255 (N_22255,N_18829,N_16551);
nor U22256 (N_22256,N_15330,N_16590);
nand U22257 (N_22257,N_18301,N_19646);
or U22258 (N_22258,N_19979,N_17938);
nor U22259 (N_22259,N_18960,N_16969);
xnor U22260 (N_22260,N_15492,N_19028);
nor U22261 (N_22261,N_18487,N_17217);
nand U22262 (N_22262,N_15066,N_18798);
nor U22263 (N_22263,N_16913,N_15767);
nand U22264 (N_22264,N_19971,N_15572);
nand U22265 (N_22265,N_16570,N_15402);
and U22266 (N_22266,N_15725,N_16438);
nand U22267 (N_22267,N_18615,N_18919);
nand U22268 (N_22268,N_18876,N_17127);
and U22269 (N_22269,N_19730,N_19435);
xnor U22270 (N_22270,N_16721,N_16490);
nand U22271 (N_22271,N_19935,N_17489);
or U22272 (N_22272,N_15318,N_17162);
nand U22273 (N_22273,N_19937,N_16158);
nor U22274 (N_22274,N_19782,N_19714);
nor U22275 (N_22275,N_17348,N_17641);
nor U22276 (N_22276,N_17625,N_19762);
and U22277 (N_22277,N_19586,N_18041);
and U22278 (N_22278,N_18412,N_15804);
and U22279 (N_22279,N_16955,N_19362);
or U22280 (N_22280,N_15344,N_15086);
nand U22281 (N_22281,N_17276,N_15388);
or U22282 (N_22282,N_17768,N_16171);
or U22283 (N_22283,N_18604,N_19648);
nor U22284 (N_22284,N_15258,N_16648);
xnor U22285 (N_22285,N_17733,N_15108);
nor U22286 (N_22286,N_17201,N_16728);
nor U22287 (N_22287,N_17853,N_19055);
nor U22288 (N_22288,N_16709,N_15431);
nand U22289 (N_22289,N_17904,N_18278);
nand U22290 (N_22290,N_16042,N_16273);
or U22291 (N_22291,N_16959,N_17197);
and U22292 (N_22292,N_17600,N_17032);
nand U22293 (N_22293,N_17165,N_18200);
or U22294 (N_22294,N_19358,N_19482);
xor U22295 (N_22295,N_17863,N_17968);
xor U22296 (N_22296,N_19323,N_17986);
xor U22297 (N_22297,N_15283,N_17325);
and U22298 (N_22298,N_18249,N_17565);
or U22299 (N_22299,N_15028,N_18969);
xor U22300 (N_22300,N_17893,N_15275);
nor U22301 (N_22301,N_19285,N_19988);
nor U22302 (N_22302,N_16130,N_15758);
nor U22303 (N_22303,N_16174,N_18160);
nor U22304 (N_22304,N_19562,N_19261);
and U22305 (N_22305,N_17709,N_17453);
and U22306 (N_22306,N_18104,N_18193);
nand U22307 (N_22307,N_19624,N_15980);
or U22308 (N_22308,N_16941,N_16810);
or U22309 (N_22309,N_19113,N_16313);
and U22310 (N_22310,N_19803,N_17566);
or U22311 (N_22311,N_19041,N_19700);
nor U22312 (N_22312,N_17293,N_16812);
and U22313 (N_22313,N_15151,N_17462);
or U22314 (N_22314,N_15609,N_15244);
nand U22315 (N_22315,N_16506,N_19162);
xor U22316 (N_22316,N_17742,N_16580);
nor U22317 (N_22317,N_15391,N_17967);
xnor U22318 (N_22318,N_18259,N_17430);
and U22319 (N_22319,N_15620,N_19737);
nand U22320 (N_22320,N_17359,N_16529);
and U22321 (N_22321,N_18999,N_17735);
or U22322 (N_22322,N_19893,N_18459);
and U22323 (N_22323,N_16347,N_19024);
nand U22324 (N_22324,N_17662,N_18493);
nor U22325 (N_22325,N_18516,N_17022);
nor U22326 (N_22326,N_17510,N_17117);
xnor U22327 (N_22327,N_15515,N_16681);
and U22328 (N_22328,N_17652,N_16816);
nand U22329 (N_22329,N_17665,N_17708);
nor U22330 (N_22330,N_16651,N_16405);
nor U22331 (N_22331,N_15514,N_19131);
nand U22332 (N_22332,N_17277,N_17269);
nand U22333 (N_22333,N_19702,N_19837);
nand U22334 (N_22334,N_15117,N_17050);
xor U22335 (N_22335,N_17755,N_19753);
or U22336 (N_22336,N_15187,N_19459);
and U22337 (N_22337,N_17042,N_18284);
nor U22338 (N_22338,N_15037,N_15011);
nor U22339 (N_22339,N_18699,N_19637);
nand U22340 (N_22340,N_16704,N_19583);
xnor U22341 (N_22341,N_16664,N_17737);
nand U22342 (N_22342,N_17750,N_17338);
nand U22343 (N_22343,N_18016,N_16251);
or U22344 (N_22344,N_18212,N_17411);
nor U22345 (N_22345,N_16946,N_17541);
and U22346 (N_22346,N_18819,N_16741);
xnor U22347 (N_22347,N_15191,N_18503);
nand U22348 (N_22348,N_18574,N_15602);
nand U22349 (N_22349,N_18378,N_16604);
and U22350 (N_22350,N_17331,N_18641);
nor U22351 (N_22351,N_19170,N_15833);
nand U22352 (N_22352,N_16811,N_15464);
and U22353 (N_22353,N_18172,N_18761);
nand U22354 (N_22354,N_18749,N_16457);
xnor U22355 (N_22355,N_15124,N_19392);
nand U22356 (N_22356,N_15825,N_16777);
nand U22357 (N_22357,N_15141,N_16254);
nor U22358 (N_22358,N_16469,N_18692);
nand U22359 (N_22359,N_15924,N_19398);
xnor U22360 (N_22360,N_19244,N_15869);
nor U22361 (N_22361,N_17961,N_16385);
and U22362 (N_22362,N_16221,N_15478);
nand U22363 (N_22363,N_18045,N_17617);
nand U22364 (N_22364,N_17594,N_15784);
nor U22365 (N_22365,N_16377,N_17583);
xnor U22366 (N_22366,N_16452,N_15487);
nand U22367 (N_22367,N_15440,N_19468);
nor U22368 (N_22368,N_17751,N_16701);
or U22369 (N_22369,N_16034,N_18569);
or U22370 (N_22370,N_19933,N_18361);
nor U22371 (N_22371,N_18986,N_17133);
or U22372 (N_22372,N_19703,N_19780);
and U22373 (N_22373,N_16303,N_19286);
and U22374 (N_22374,N_15032,N_19360);
nand U22375 (N_22375,N_19977,N_16124);
nand U22376 (N_22376,N_17186,N_19647);
xnor U22377 (N_22377,N_15465,N_19383);
and U22378 (N_22378,N_17874,N_16148);
xor U22379 (N_22379,N_18020,N_15077);
nand U22380 (N_22380,N_15730,N_17545);
xor U22381 (N_22381,N_18822,N_17369);
xor U22382 (N_22382,N_16163,N_18715);
and U22383 (N_22383,N_16863,N_17270);
nor U22384 (N_22384,N_19538,N_18837);
nand U22385 (N_22385,N_16049,N_18706);
and U22386 (N_22386,N_17644,N_15008);
nor U22387 (N_22387,N_16639,N_17443);
or U22388 (N_22388,N_15350,N_18214);
nand U22389 (N_22389,N_18792,N_18672);
nand U22390 (N_22390,N_18954,N_17097);
and U22391 (N_22391,N_16222,N_15512);
nand U22392 (N_22392,N_16952,N_16297);
xnor U22393 (N_22393,N_18595,N_16252);
nor U22394 (N_22394,N_16883,N_19102);
nand U22395 (N_22395,N_18231,N_15125);
or U22396 (N_22396,N_18888,N_15300);
and U22397 (N_22397,N_15686,N_15122);
or U22398 (N_22398,N_19891,N_18814);
nor U22399 (N_22399,N_19774,N_15526);
xor U22400 (N_22400,N_15057,N_15395);
nand U22401 (N_22401,N_19441,N_18507);
xnor U22402 (N_22402,N_18891,N_17418);
nand U22403 (N_22403,N_19226,N_15633);
or U22404 (N_22404,N_18693,N_19862);
xor U22405 (N_22405,N_16383,N_18557);
xor U22406 (N_22406,N_18579,N_16256);
nand U22407 (N_22407,N_17400,N_18098);
xor U22408 (N_22408,N_19800,N_16258);
nor U22409 (N_22409,N_19990,N_18733);
nand U22410 (N_22410,N_18536,N_18832);
nor U22411 (N_22411,N_16044,N_16847);
nor U22412 (N_22412,N_16951,N_17413);
or U22413 (N_22413,N_16086,N_16443);
and U22414 (N_22414,N_16990,N_17820);
xnor U22415 (N_22415,N_15799,N_15036);
nand U22416 (N_22416,N_16830,N_18565);
xnor U22417 (N_22417,N_15597,N_19788);
xnor U22418 (N_22418,N_17796,N_15855);
nor U22419 (N_22419,N_19305,N_15235);
xor U22420 (N_22420,N_18484,N_16493);
xor U22421 (N_22421,N_18199,N_19926);
xor U22422 (N_22422,N_16037,N_18009);
nor U22423 (N_22423,N_18305,N_16445);
and U22424 (N_22424,N_16838,N_17818);
xnor U22425 (N_22425,N_17552,N_16869);
nor U22426 (N_22426,N_16156,N_15341);
nor U22427 (N_22427,N_17273,N_16424);
and U22428 (N_22428,N_16276,N_16112);
and U22429 (N_22429,N_17212,N_17843);
xnor U22430 (N_22430,N_16690,N_17079);
or U22431 (N_22431,N_17229,N_19593);
nor U22432 (N_22432,N_18167,N_18644);
xor U22433 (N_22433,N_19182,N_19331);
nor U22434 (N_22434,N_17658,N_16339);
xnor U22435 (N_22435,N_18068,N_15777);
or U22436 (N_22436,N_15242,N_16642);
xnor U22437 (N_22437,N_16177,N_16500);
and U22438 (N_22438,N_19356,N_16301);
nor U22439 (N_22439,N_16341,N_18246);
or U22440 (N_22440,N_17996,N_19277);
nand U22441 (N_22441,N_18337,N_16245);
nand U22442 (N_22442,N_16903,N_19620);
or U22443 (N_22443,N_19485,N_17450);
xnor U22444 (N_22444,N_15761,N_18480);
nor U22445 (N_22445,N_17295,N_16244);
nor U22446 (N_22446,N_19147,N_15561);
and U22447 (N_22447,N_19980,N_18697);
nor U22448 (N_22448,N_18799,N_15301);
xnor U22449 (N_22449,N_15697,N_17305);
nand U22450 (N_22450,N_16947,N_17215);
and U22451 (N_22451,N_18145,N_19958);
nor U22452 (N_22452,N_18498,N_18067);
and U22453 (N_22453,N_15332,N_15022);
or U22454 (N_22454,N_19350,N_19192);
and U22455 (N_22455,N_16232,N_16359);
xor U22456 (N_22456,N_19553,N_15239);
and U22457 (N_22457,N_15174,N_18255);
nand U22458 (N_22458,N_16069,N_18562);
or U22459 (N_22459,N_17391,N_17946);
and U22460 (N_22460,N_18781,N_16596);
or U22461 (N_22461,N_16542,N_18538);
or U22462 (N_22462,N_15606,N_18915);
nand U22463 (N_22463,N_16048,N_18973);
and U22464 (N_22464,N_18629,N_19607);
nand U22465 (N_22465,N_18926,N_19333);
nand U22466 (N_22466,N_16145,N_19506);
nor U22467 (N_22467,N_15545,N_19535);
or U22468 (N_22468,N_19632,N_15942);
nand U22469 (N_22469,N_15744,N_18647);
xor U22470 (N_22470,N_16397,N_15398);
and U22471 (N_22471,N_16755,N_17569);
xor U22472 (N_22472,N_17445,N_19190);
nand U22473 (N_22473,N_17744,N_15729);
nor U22474 (N_22474,N_18782,N_17831);
and U22475 (N_22475,N_17524,N_15960);
nand U22476 (N_22476,N_15302,N_17128);
nand U22477 (N_22477,N_16326,N_18342);
and U22478 (N_22478,N_16123,N_19551);
xor U22479 (N_22479,N_19090,N_19866);
xnor U22480 (N_22480,N_17795,N_15212);
and U22481 (N_22481,N_15889,N_18972);
nand U22482 (N_22482,N_18071,N_18842);
nor U22483 (N_22483,N_18472,N_19836);
nor U22484 (N_22484,N_15610,N_17911);
or U22485 (N_22485,N_16353,N_17731);
nor U22486 (N_22486,N_18348,N_17372);
and U22487 (N_22487,N_15365,N_15449);
and U22488 (N_22488,N_16323,N_16186);
nor U22489 (N_22489,N_15484,N_17182);
xor U22490 (N_22490,N_15129,N_17876);
or U22491 (N_22491,N_17412,N_15453);
and U22492 (N_22492,N_18149,N_16414);
and U22493 (N_22493,N_17251,N_18515);
nor U22494 (N_22494,N_18079,N_15284);
or U22495 (N_22495,N_17484,N_19016);
xor U22496 (N_22496,N_16813,N_17799);
nand U22497 (N_22497,N_15252,N_17516);
xor U22498 (N_22498,N_16842,N_15598);
nor U22499 (N_22499,N_19758,N_17383);
nor U22500 (N_22500,N_15610,N_15739);
xor U22501 (N_22501,N_19081,N_18816);
xor U22502 (N_22502,N_19602,N_19784);
and U22503 (N_22503,N_18317,N_19843);
nor U22504 (N_22504,N_19503,N_17663);
nor U22505 (N_22505,N_19770,N_16038);
nor U22506 (N_22506,N_15482,N_18150);
nand U22507 (N_22507,N_17950,N_17212);
xnor U22508 (N_22508,N_19941,N_18932);
nand U22509 (N_22509,N_18373,N_15567);
xor U22510 (N_22510,N_19016,N_19886);
nor U22511 (N_22511,N_15478,N_15280);
or U22512 (N_22512,N_16466,N_15535);
or U22513 (N_22513,N_19185,N_19105);
and U22514 (N_22514,N_18696,N_17537);
or U22515 (N_22515,N_15111,N_16188);
nor U22516 (N_22516,N_15996,N_15341);
and U22517 (N_22517,N_18239,N_18698);
nor U22518 (N_22518,N_15844,N_15786);
nor U22519 (N_22519,N_15949,N_15732);
xnor U22520 (N_22520,N_16075,N_16451);
nor U22521 (N_22521,N_16253,N_19571);
xnor U22522 (N_22522,N_19082,N_16993);
or U22523 (N_22523,N_19018,N_17588);
and U22524 (N_22524,N_16729,N_15950);
xnor U22525 (N_22525,N_19401,N_18115);
nand U22526 (N_22526,N_17793,N_17639);
or U22527 (N_22527,N_17706,N_17637);
nor U22528 (N_22528,N_17320,N_17252);
or U22529 (N_22529,N_15363,N_18497);
nor U22530 (N_22530,N_17690,N_17618);
and U22531 (N_22531,N_19489,N_15649);
and U22532 (N_22532,N_18394,N_19325);
and U22533 (N_22533,N_18302,N_18596);
nand U22534 (N_22534,N_17775,N_19800);
xnor U22535 (N_22535,N_18188,N_18652);
nand U22536 (N_22536,N_19166,N_18955);
xor U22537 (N_22537,N_18814,N_17117);
nor U22538 (N_22538,N_16098,N_16200);
nand U22539 (N_22539,N_18109,N_17902);
and U22540 (N_22540,N_19516,N_16313);
or U22541 (N_22541,N_15394,N_15568);
and U22542 (N_22542,N_15534,N_17080);
nor U22543 (N_22543,N_18729,N_16207);
xnor U22544 (N_22544,N_18451,N_18729);
or U22545 (N_22545,N_15186,N_19813);
nand U22546 (N_22546,N_17735,N_16101);
nor U22547 (N_22547,N_17888,N_15871);
and U22548 (N_22548,N_16671,N_15633);
xor U22549 (N_22549,N_17288,N_18367);
nor U22550 (N_22550,N_17196,N_16651);
and U22551 (N_22551,N_19009,N_16777);
nand U22552 (N_22552,N_19793,N_19461);
or U22553 (N_22553,N_19546,N_17882);
xor U22554 (N_22554,N_19078,N_19890);
nor U22555 (N_22555,N_15830,N_18598);
or U22556 (N_22556,N_19735,N_17484);
nand U22557 (N_22557,N_18924,N_15259);
nand U22558 (N_22558,N_17741,N_18865);
nand U22559 (N_22559,N_19217,N_15954);
nand U22560 (N_22560,N_19237,N_19505);
nor U22561 (N_22561,N_17346,N_16709);
xor U22562 (N_22562,N_17488,N_15524);
xor U22563 (N_22563,N_17254,N_18687);
nand U22564 (N_22564,N_19093,N_15859);
nor U22565 (N_22565,N_17067,N_17303);
and U22566 (N_22566,N_16851,N_18653);
or U22567 (N_22567,N_16334,N_16006);
xor U22568 (N_22568,N_19052,N_16041);
nand U22569 (N_22569,N_19025,N_16903);
or U22570 (N_22570,N_18879,N_19991);
xor U22571 (N_22571,N_19613,N_16231);
xnor U22572 (N_22572,N_17118,N_18909);
or U22573 (N_22573,N_19617,N_19695);
and U22574 (N_22574,N_18968,N_17668);
nor U22575 (N_22575,N_17615,N_16237);
and U22576 (N_22576,N_19784,N_18351);
nand U22577 (N_22577,N_17408,N_18006);
nor U22578 (N_22578,N_16940,N_15267);
xor U22579 (N_22579,N_19930,N_15607);
xnor U22580 (N_22580,N_15501,N_17523);
and U22581 (N_22581,N_18510,N_16944);
or U22582 (N_22582,N_17139,N_17673);
and U22583 (N_22583,N_19183,N_19582);
or U22584 (N_22584,N_19078,N_19071);
nor U22585 (N_22585,N_15663,N_15827);
and U22586 (N_22586,N_15752,N_16050);
xor U22587 (N_22587,N_17231,N_19064);
xnor U22588 (N_22588,N_18454,N_17647);
or U22589 (N_22589,N_18243,N_19742);
or U22590 (N_22590,N_18875,N_17833);
nor U22591 (N_22591,N_17955,N_18378);
and U22592 (N_22592,N_15882,N_16730);
or U22593 (N_22593,N_17949,N_18894);
xnor U22594 (N_22594,N_18370,N_15283);
or U22595 (N_22595,N_18948,N_15565);
and U22596 (N_22596,N_19611,N_15642);
or U22597 (N_22597,N_18909,N_19698);
nand U22598 (N_22598,N_19406,N_16382);
and U22599 (N_22599,N_18768,N_19697);
or U22600 (N_22600,N_18075,N_16134);
nand U22601 (N_22601,N_18112,N_19793);
xnor U22602 (N_22602,N_19053,N_16040);
and U22603 (N_22603,N_18879,N_19891);
nand U22604 (N_22604,N_15097,N_17727);
nand U22605 (N_22605,N_17520,N_18264);
and U22606 (N_22606,N_17541,N_17798);
or U22607 (N_22607,N_15655,N_18740);
nand U22608 (N_22608,N_19018,N_17108);
or U22609 (N_22609,N_18469,N_15210);
nand U22610 (N_22610,N_16717,N_15278);
and U22611 (N_22611,N_18556,N_19547);
or U22612 (N_22612,N_19367,N_17702);
and U22613 (N_22613,N_19962,N_15820);
nand U22614 (N_22614,N_16114,N_19801);
xnor U22615 (N_22615,N_15086,N_19544);
xor U22616 (N_22616,N_18205,N_19267);
nor U22617 (N_22617,N_15478,N_15822);
or U22618 (N_22618,N_17064,N_16879);
nor U22619 (N_22619,N_17155,N_15802);
nand U22620 (N_22620,N_15359,N_16548);
xnor U22621 (N_22621,N_15939,N_15947);
nor U22622 (N_22622,N_15250,N_19886);
or U22623 (N_22623,N_16801,N_18459);
nor U22624 (N_22624,N_16049,N_17664);
or U22625 (N_22625,N_17007,N_18678);
and U22626 (N_22626,N_15336,N_18573);
xnor U22627 (N_22627,N_15201,N_15209);
xnor U22628 (N_22628,N_19305,N_19720);
xor U22629 (N_22629,N_15311,N_19560);
or U22630 (N_22630,N_18264,N_18535);
nand U22631 (N_22631,N_15750,N_19150);
nand U22632 (N_22632,N_18634,N_16645);
or U22633 (N_22633,N_17399,N_19256);
or U22634 (N_22634,N_19439,N_17950);
xnor U22635 (N_22635,N_17522,N_17948);
and U22636 (N_22636,N_16323,N_18185);
nand U22637 (N_22637,N_17393,N_15568);
xnor U22638 (N_22638,N_18469,N_18143);
nor U22639 (N_22639,N_18047,N_19180);
nand U22640 (N_22640,N_18818,N_18779);
xor U22641 (N_22641,N_15721,N_18714);
or U22642 (N_22642,N_17949,N_17791);
xnor U22643 (N_22643,N_16783,N_16432);
xnor U22644 (N_22644,N_16574,N_17768);
xor U22645 (N_22645,N_19022,N_19195);
xnor U22646 (N_22646,N_19085,N_18550);
nand U22647 (N_22647,N_16436,N_18036);
or U22648 (N_22648,N_18560,N_17201);
and U22649 (N_22649,N_16311,N_15552);
and U22650 (N_22650,N_19235,N_16664);
xor U22651 (N_22651,N_17506,N_19135);
nand U22652 (N_22652,N_15723,N_17730);
or U22653 (N_22653,N_17250,N_16414);
nand U22654 (N_22654,N_15210,N_17719);
xnor U22655 (N_22655,N_15165,N_15669);
nand U22656 (N_22656,N_18676,N_15726);
nor U22657 (N_22657,N_18235,N_16308);
or U22658 (N_22658,N_19073,N_17073);
and U22659 (N_22659,N_17770,N_17110);
nor U22660 (N_22660,N_16484,N_19157);
nand U22661 (N_22661,N_15025,N_16400);
xnor U22662 (N_22662,N_15805,N_18013);
xnor U22663 (N_22663,N_18480,N_19753);
nand U22664 (N_22664,N_17867,N_17360);
xnor U22665 (N_22665,N_18814,N_19894);
nand U22666 (N_22666,N_19479,N_15581);
and U22667 (N_22667,N_15971,N_18166);
nand U22668 (N_22668,N_19328,N_19337);
nor U22669 (N_22669,N_19379,N_19675);
xnor U22670 (N_22670,N_16125,N_19203);
xnor U22671 (N_22671,N_17507,N_17470);
nor U22672 (N_22672,N_19857,N_17310);
xnor U22673 (N_22673,N_19521,N_18508);
and U22674 (N_22674,N_18181,N_19881);
nand U22675 (N_22675,N_17406,N_19441);
nand U22676 (N_22676,N_18888,N_16333);
nand U22677 (N_22677,N_15648,N_16603);
and U22678 (N_22678,N_17500,N_16282);
xnor U22679 (N_22679,N_16526,N_18757);
nand U22680 (N_22680,N_19782,N_15280);
or U22681 (N_22681,N_17037,N_16321);
or U22682 (N_22682,N_15858,N_16026);
xnor U22683 (N_22683,N_17259,N_15277);
or U22684 (N_22684,N_16008,N_18435);
xnor U22685 (N_22685,N_18005,N_16230);
and U22686 (N_22686,N_17009,N_17829);
or U22687 (N_22687,N_18377,N_19998);
or U22688 (N_22688,N_19337,N_19557);
xor U22689 (N_22689,N_17740,N_16580);
xnor U22690 (N_22690,N_17949,N_18701);
nor U22691 (N_22691,N_15463,N_19867);
and U22692 (N_22692,N_15593,N_17307);
nand U22693 (N_22693,N_16300,N_18018);
xor U22694 (N_22694,N_15909,N_15295);
nor U22695 (N_22695,N_17864,N_15357);
nor U22696 (N_22696,N_18908,N_18941);
nand U22697 (N_22697,N_18373,N_16360);
xnor U22698 (N_22698,N_15403,N_16013);
nand U22699 (N_22699,N_16591,N_18148);
nor U22700 (N_22700,N_19919,N_17042);
nand U22701 (N_22701,N_18923,N_18593);
nor U22702 (N_22702,N_15277,N_16099);
nand U22703 (N_22703,N_19449,N_19104);
nand U22704 (N_22704,N_16720,N_19494);
xor U22705 (N_22705,N_18408,N_18742);
xor U22706 (N_22706,N_16236,N_15648);
xnor U22707 (N_22707,N_17492,N_16946);
nand U22708 (N_22708,N_19191,N_15426);
xor U22709 (N_22709,N_18227,N_18397);
nand U22710 (N_22710,N_16449,N_16674);
or U22711 (N_22711,N_15352,N_18255);
nor U22712 (N_22712,N_18393,N_15587);
nand U22713 (N_22713,N_15151,N_17100);
nand U22714 (N_22714,N_15685,N_17131);
xor U22715 (N_22715,N_15301,N_16836);
nor U22716 (N_22716,N_16214,N_18616);
and U22717 (N_22717,N_18263,N_15138);
and U22718 (N_22718,N_18888,N_17811);
xor U22719 (N_22719,N_19398,N_15194);
xnor U22720 (N_22720,N_19298,N_18337);
xnor U22721 (N_22721,N_15217,N_18890);
nor U22722 (N_22722,N_17945,N_16552);
and U22723 (N_22723,N_19804,N_18294);
nor U22724 (N_22724,N_18055,N_16543);
nor U22725 (N_22725,N_17101,N_15787);
nor U22726 (N_22726,N_15463,N_17051);
or U22727 (N_22727,N_16989,N_18914);
nor U22728 (N_22728,N_17321,N_18809);
nand U22729 (N_22729,N_15348,N_16431);
or U22730 (N_22730,N_15010,N_18793);
nor U22731 (N_22731,N_19353,N_19423);
xnor U22732 (N_22732,N_19397,N_18493);
nor U22733 (N_22733,N_17926,N_18580);
nor U22734 (N_22734,N_18731,N_18036);
or U22735 (N_22735,N_18949,N_15309);
or U22736 (N_22736,N_17768,N_19983);
or U22737 (N_22737,N_16232,N_16856);
xnor U22738 (N_22738,N_19189,N_17930);
and U22739 (N_22739,N_17213,N_15426);
xnor U22740 (N_22740,N_17038,N_19375);
or U22741 (N_22741,N_15291,N_18956);
nor U22742 (N_22742,N_15591,N_16924);
or U22743 (N_22743,N_19321,N_19671);
or U22744 (N_22744,N_16771,N_19818);
nand U22745 (N_22745,N_15033,N_17118);
and U22746 (N_22746,N_17796,N_17146);
or U22747 (N_22747,N_16395,N_17602);
and U22748 (N_22748,N_16733,N_16280);
and U22749 (N_22749,N_15871,N_17425);
xor U22750 (N_22750,N_19887,N_17910);
xor U22751 (N_22751,N_17472,N_16737);
nor U22752 (N_22752,N_16395,N_18794);
xor U22753 (N_22753,N_19708,N_17763);
or U22754 (N_22754,N_17961,N_17134);
and U22755 (N_22755,N_18994,N_17219);
xor U22756 (N_22756,N_16963,N_16945);
or U22757 (N_22757,N_17690,N_16243);
xor U22758 (N_22758,N_15819,N_15692);
nand U22759 (N_22759,N_16169,N_18680);
nand U22760 (N_22760,N_15757,N_16114);
xor U22761 (N_22761,N_15794,N_17132);
nor U22762 (N_22762,N_19552,N_18218);
nor U22763 (N_22763,N_19791,N_17099);
nor U22764 (N_22764,N_18301,N_15558);
and U22765 (N_22765,N_15793,N_16949);
nor U22766 (N_22766,N_15815,N_18989);
or U22767 (N_22767,N_19412,N_19418);
and U22768 (N_22768,N_17571,N_19586);
nand U22769 (N_22769,N_19818,N_18960);
nand U22770 (N_22770,N_19872,N_18352);
nand U22771 (N_22771,N_17386,N_19194);
nand U22772 (N_22772,N_18130,N_16553);
xor U22773 (N_22773,N_18616,N_19395);
nand U22774 (N_22774,N_17982,N_18900);
xor U22775 (N_22775,N_16676,N_17760);
and U22776 (N_22776,N_16954,N_19358);
or U22777 (N_22777,N_19737,N_17038);
nor U22778 (N_22778,N_17177,N_19284);
xnor U22779 (N_22779,N_19240,N_18132);
or U22780 (N_22780,N_15074,N_16176);
xor U22781 (N_22781,N_16018,N_16177);
nor U22782 (N_22782,N_19499,N_19493);
nand U22783 (N_22783,N_15634,N_18230);
nand U22784 (N_22784,N_18890,N_17985);
and U22785 (N_22785,N_19013,N_17741);
and U22786 (N_22786,N_17182,N_19016);
xor U22787 (N_22787,N_15965,N_16830);
nand U22788 (N_22788,N_15372,N_18639);
or U22789 (N_22789,N_15048,N_15378);
nor U22790 (N_22790,N_18464,N_17921);
or U22791 (N_22791,N_17260,N_16614);
and U22792 (N_22792,N_16623,N_15700);
xor U22793 (N_22793,N_19315,N_16338);
and U22794 (N_22794,N_17665,N_17323);
and U22795 (N_22795,N_18042,N_17327);
xnor U22796 (N_22796,N_18104,N_15162);
nand U22797 (N_22797,N_16688,N_17577);
nor U22798 (N_22798,N_18163,N_18707);
xor U22799 (N_22799,N_19729,N_16210);
nor U22800 (N_22800,N_18910,N_18378);
and U22801 (N_22801,N_15392,N_17501);
or U22802 (N_22802,N_16640,N_18560);
xor U22803 (N_22803,N_19764,N_15912);
nand U22804 (N_22804,N_17220,N_18354);
nor U22805 (N_22805,N_18933,N_19334);
or U22806 (N_22806,N_17447,N_17372);
xor U22807 (N_22807,N_19137,N_15989);
xor U22808 (N_22808,N_15947,N_17771);
nand U22809 (N_22809,N_16746,N_15469);
or U22810 (N_22810,N_17086,N_17926);
nand U22811 (N_22811,N_19700,N_17990);
or U22812 (N_22812,N_16086,N_19026);
nand U22813 (N_22813,N_15670,N_18524);
xor U22814 (N_22814,N_18691,N_15467);
xor U22815 (N_22815,N_18449,N_16499);
nand U22816 (N_22816,N_17557,N_16995);
nor U22817 (N_22817,N_16596,N_18337);
nand U22818 (N_22818,N_19401,N_19583);
nor U22819 (N_22819,N_17344,N_19862);
nand U22820 (N_22820,N_17669,N_15572);
nor U22821 (N_22821,N_18547,N_18089);
and U22822 (N_22822,N_17248,N_17522);
nor U22823 (N_22823,N_16049,N_19352);
xnor U22824 (N_22824,N_19147,N_16919);
nor U22825 (N_22825,N_17138,N_17020);
and U22826 (N_22826,N_16663,N_19087);
xnor U22827 (N_22827,N_18915,N_17685);
xor U22828 (N_22828,N_18554,N_18649);
nand U22829 (N_22829,N_17694,N_16853);
and U22830 (N_22830,N_16781,N_15804);
nor U22831 (N_22831,N_16490,N_19446);
nand U22832 (N_22832,N_18484,N_15208);
and U22833 (N_22833,N_18333,N_16667);
or U22834 (N_22834,N_17990,N_16711);
and U22835 (N_22835,N_15156,N_16172);
and U22836 (N_22836,N_19421,N_15771);
nand U22837 (N_22837,N_19271,N_18293);
nor U22838 (N_22838,N_15428,N_16920);
nand U22839 (N_22839,N_19096,N_19047);
or U22840 (N_22840,N_17829,N_19741);
xnor U22841 (N_22841,N_19942,N_17734);
nor U22842 (N_22842,N_18083,N_16636);
or U22843 (N_22843,N_17811,N_16974);
nand U22844 (N_22844,N_17473,N_16113);
or U22845 (N_22845,N_15895,N_19797);
nor U22846 (N_22846,N_15080,N_16631);
nor U22847 (N_22847,N_15271,N_17150);
nor U22848 (N_22848,N_19109,N_19262);
nor U22849 (N_22849,N_16768,N_19008);
xnor U22850 (N_22850,N_19850,N_18221);
xnor U22851 (N_22851,N_18223,N_19290);
xnor U22852 (N_22852,N_19172,N_19463);
and U22853 (N_22853,N_16522,N_16414);
xor U22854 (N_22854,N_17451,N_19598);
nor U22855 (N_22855,N_19650,N_19230);
and U22856 (N_22856,N_16346,N_19073);
nor U22857 (N_22857,N_19371,N_16049);
or U22858 (N_22858,N_15008,N_17541);
nand U22859 (N_22859,N_19762,N_19183);
or U22860 (N_22860,N_15528,N_18842);
xor U22861 (N_22861,N_17760,N_15050);
nor U22862 (N_22862,N_19736,N_19013);
nor U22863 (N_22863,N_16670,N_17097);
or U22864 (N_22864,N_16101,N_18293);
or U22865 (N_22865,N_18174,N_18316);
xor U22866 (N_22866,N_18331,N_15514);
or U22867 (N_22867,N_15520,N_19607);
xor U22868 (N_22868,N_16817,N_15222);
xor U22869 (N_22869,N_19729,N_19785);
or U22870 (N_22870,N_19903,N_17474);
or U22871 (N_22871,N_17086,N_19577);
and U22872 (N_22872,N_15790,N_19220);
and U22873 (N_22873,N_17307,N_15773);
nand U22874 (N_22874,N_17194,N_18172);
xnor U22875 (N_22875,N_15898,N_15536);
nand U22876 (N_22876,N_17776,N_17191);
or U22877 (N_22877,N_15732,N_19076);
xnor U22878 (N_22878,N_19880,N_16913);
xnor U22879 (N_22879,N_17596,N_19813);
nand U22880 (N_22880,N_17910,N_19072);
nand U22881 (N_22881,N_16427,N_18218);
nor U22882 (N_22882,N_18873,N_19227);
nand U22883 (N_22883,N_16658,N_15963);
xnor U22884 (N_22884,N_19226,N_18044);
nor U22885 (N_22885,N_16773,N_17674);
xnor U22886 (N_22886,N_19443,N_15584);
and U22887 (N_22887,N_16963,N_19801);
xor U22888 (N_22888,N_16658,N_16975);
and U22889 (N_22889,N_16307,N_17176);
or U22890 (N_22890,N_15104,N_17327);
or U22891 (N_22891,N_18258,N_19347);
nor U22892 (N_22892,N_19540,N_15696);
nor U22893 (N_22893,N_16470,N_18243);
and U22894 (N_22894,N_19113,N_16590);
nor U22895 (N_22895,N_18613,N_15918);
nand U22896 (N_22896,N_19130,N_15606);
nor U22897 (N_22897,N_17366,N_17373);
and U22898 (N_22898,N_17826,N_19571);
xor U22899 (N_22899,N_16638,N_18413);
nor U22900 (N_22900,N_19757,N_19324);
xnor U22901 (N_22901,N_15401,N_17250);
and U22902 (N_22902,N_18600,N_16948);
or U22903 (N_22903,N_15550,N_19299);
nand U22904 (N_22904,N_18537,N_18118);
xor U22905 (N_22905,N_18385,N_18414);
nand U22906 (N_22906,N_18483,N_17995);
nand U22907 (N_22907,N_17414,N_19885);
or U22908 (N_22908,N_17753,N_19168);
nand U22909 (N_22909,N_18970,N_16944);
xor U22910 (N_22910,N_16054,N_18685);
xor U22911 (N_22911,N_16347,N_19243);
or U22912 (N_22912,N_15069,N_19952);
or U22913 (N_22913,N_15777,N_15977);
nor U22914 (N_22914,N_16385,N_16593);
nand U22915 (N_22915,N_19604,N_19348);
and U22916 (N_22916,N_15627,N_15966);
or U22917 (N_22917,N_16196,N_17530);
nand U22918 (N_22918,N_18323,N_18831);
nand U22919 (N_22919,N_18031,N_17844);
nor U22920 (N_22920,N_15892,N_18744);
nor U22921 (N_22921,N_18666,N_19495);
and U22922 (N_22922,N_15240,N_16100);
nor U22923 (N_22923,N_15413,N_15430);
nand U22924 (N_22924,N_17298,N_15901);
nand U22925 (N_22925,N_19909,N_15774);
xor U22926 (N_22926,N_19266,N_15914);
nand U22927 (N_22927,N_19315,N_15499);
and U22928 (N_22928,N_16565,N_19700);
or U22929 (N_22929,N_17174,N_16984);
or U22930 (N_22930,N_15439,N_16550);
or U22931 (N_22931,N_15850,N_17900);
and U22932 (N_22932,N_15528,N_17964);
xor U22933 (N_22933,N_15884,N_18543);
and U22934 (N_22934,N_17976,N_18821);
nor U22935 (N_22935,N_17485,N_19915);
or U22936 (N_22936,N_18124,N_19217);
nor U22937 (N_22937,N_19772,N_15479);
xnor U22938 (N_22938,N_18618,N_15906);
nand U22939 (N_22939,N_17272,N_19775);
and U22940 (N_22940,N_17800,N_19550);
xnor U22941 (N_22941,N_15736,N_16562);
or U22942 (N_22942,N_19257,N_16022);
nor U22943 (N_22943,N_18408,N_15454);
nand U22944 (N_22944,N_17162,N_16397);
nand U22945 (N_22945,N_15679,N_16407);
or U22946 (N_22946,N_17531,N_18946);
nand U22947 (N_22947,N_19995,N_16215);
nor U22948 (N_22948,N_17407,N_16805);
or U22949 (N_22949,N_19226,N_19681);
and U22950 (N_22950,N_18480,N_18590);
nand U22951 (N_22951,N_15986,N_18883);
xor U22952 (N_22952,N_15938,N_18861);
xnor U22953 (N_22953,N_17541,N_19990);
or U22954 (N_22954,N_17527,N_18327);
nand U22955 (N_22955,N_17616,N_17939);
nand U22956 (N_22956,N_15499,N_18671);
and U22957 (N_22957,N_19058,N_19959);
and U22958 (N_22958,N_19384,N_19141);
nor U22959 (N_22959,N_17140,N_18983);
nand U22960 (N_22960,N_18168,N_18389);
nand U22961 (N_22961,N_17635,N_16486);
xor U22962 (N_22962,N_16396,N_18827);
or U22963 (N_22963,N_19731,N_17142);
xor U22964 (N_22964,N_17396,N_19980);
nor U22965 (N_22965,N_19995,N_17392);
nor U22966 (N_22966,N_16218,N_16959);
and U22967 (N_22967,N_16902,N_17208);
xnor U22968 (N_22968,N_15904,N_17848);
nor U22969 (N_22969,N_15292,N_16947);
and U22970 (N_22970,N_16921,N_15040);
nand U22971 (N_22971,N_15638,N_16069);
or U22972 (N_22972,N_16327,N_16992);
or U22973 (N_22973,N_19823,N_18475);
xnor U22974 (N_22974,N_17835,N_17419);
nor U22975 (N_22975,N_19431,N_19063);
nand U22976 (N_22976,N_18483,N_19443);
or U22977 (N_22977,N_19648,N_19439);
nand U22978 (N_22978,N_16504,N_17745);
and U22979 (N_22979,N_15248,N_17508);
or U22980 (N_22980,N_19230,N_18431);
or U22981 (N_22981,N_19710,N_17330);
and U22982 (N_22982,N_15096,N_19077);
or U22983 (N_22983,N_17343,N_18307);
and U22984 (N_22984,N_19962,N_18842);
or U22985 (N_22985,N_19338,N_17441);
nand U22986 (N_22986,N_15528,N_19467);
and U22987 (N_22987,N_18310,N_17826);
and U22988 (N_22988,N_15439,N_16926);
or U22989 (N_22989,N_19892,N_18745);
xor U22990 (N_22990,N_16227,N_19469);
xnor U22991 (N_22991,N_19698,N_18333);
nand U22992 (N_22992,N_19913,N_16484);
nor U22993 (N_22993,N_16576,N_16353);
nor U22994 (N_22994,N_15942,N_19755);
or U22995 (N_22995,N_15619,N_19989);
nor U22996 (N_22996,N_18414,N_19973);
and U22997 (N_22997,N_15560,N_16757);
nand U22998 (N_22998,N_16647,N_17692);
or U22999 (N_22999,N_16870,N_16176);
xnor U23000 (N_23000,N_18116,N_17833);
xnor U23001 (N_23001,N_16746,N_19044);
nor U23002 (N_23002,N_16400,N_18598);
and U23003 (N_23003,N_15449,N_17547);
or U23004 (N_23004,N_18648,N_15400);
xnor U23005 (N_23005,N_15735,N_19886);
xnor U23006 (N_23006,N_15204,N_15087);
xor U23007 (N_23007,N_15154,N_16034);
nor U23008 (N_23008,N_18884,N_15656);
nand U23009 (N_23009,N_18726,N_15983);
and U23010 (N_23010,N_15796,N_15615);
or U23011 (N_23011,N_19027,N_19315);
or U23012 (N_23012,N_15405,N_16407);
nor U23013 (N_23013,N_18027,N_16926);
and U23014 (N_23014,N_16344,N_15386);
xnor U23015 (N_23015,N_17502,N_16675);
xor U23016 (N_23016,N_19818,N_15639);
or U23017 (N_23017,N_18176,N_16391);
nor U23018 (N_23018,N_18031,N_16416);
or U23019 (N_23019,N_17727,N_15247);
or U23020 (N_23020,N_18654,N_19511);
xor U23021 (N_23021,N_19754,N_19948);
nor U23022 (N_23022,N_19368,N_16137);
xor U23023 (N_23023,N_15605,N_15241);
and U23024 (N_23024,N_17427,N_16254);
and U23025 (N_23025,N_19805,N_16589);
or U23026 (N_23026,N_17553,N_19694);
nand U23027 (N_23027,N_16218,N_15619);
nand U23028 (N_23028,N_17845,N_19608);
or U23029 (N_23029,N_17089,N_15674);
nor U23030 (N_23030,N_16863,N_16028);
and U23031 (N_23031,N_19966,N_19531);
nor U23032 (N_23032,N_17776,N_17733);
nor U23033 (N_23033,N_15149,N_16421);
nand U23034 (N_23034,N_16911,N_15571);
nand U23035 (N_23035,N_17929,N_15594);
nand U23036 (N_23036,N_18870,N_19737);
nand U23037 (N_23037,N_15111,N_18594);
or U23038 (N_23038,N_18489,N_19158);
and U23039 (N_23039,N_18201,N_19503);
or U23040 (N_23040,N_15781,N_18174);
xor U23041 (N_23041,N_18329,N_18729);
or U23042 (N_23042,N_16965,N_18520);
nand U23043 (N_23043,N_19269,N_17160);
nand U23044 (N_23044,N_19334,N_16797);
nor U23045 (N_23045,N_17588,N_17704);
or U23046 (N_23046,N_16983,N_15571);
xor U23047 (N_23047,N_17036,N_19491);
nand U23048 (N_23048,N_17044,N_19749);
nor U23049 (N_23049,N_19159,N_19537);
nor U23050 (N_23050,N_17430,N_16074);
or U23051 (N_23051,N_19258,N_15887);
xnor U23052 (N_23052,N_15747,N_16038);
or U23053 (N_23053,N_15732,N_17168);
and U23054 (N_23054,N_19280,N_18844);
or U23055 (N_23055,N_19585,N_19767);
xor U23056 (N_23056,N_19030,N_17247);
and U23057 (N_23057,N_19293,N_15713);
and U23058 (N_23058,N_19817,N_17084);
xor U23059 (N_23059,N_16679,N_16865);
nand U23060 (N_23060,N_15913,N_16063);
and U23061 (N_23061,N_16293,N_15960);
or U23062 (N_23062,N_17534,N_18112);
or U23063 (N_23063,N_15642,N_15107);
or U23064 (N_23064,N_16157,N_17451);
or U23065 (N_23065,N_19064,N_18331);
and U23066 (N_23066,N_18535,N_17795);
or U23067 (N_23067,N_18650,N_15599);
nand U23068 (N_23068,N_16378,N_19482);
xnor U23069 (N_23069,N_16612,N_17476);
nor U23070 (N_23070,N_17656,N_19938);
or U23071 (N_23071,N_17029,N_15339);
nor U23072 (N_23072,N_15799,N_15104);
nand U23073 (N_23073,N_17426,N_17768);
or U23074 (N_23074,N_15703,N_16242);
and U23075 (N_23075,N_17073,N_18321);
nor U23076 (N_23076,N_18878,N_16393);
and U23077 (N_23077,N_18784,N_15155);
xnor U23078 (N_23078,N_18005,N_19933);
or U23079 (N_23079,N_18638,N_19910);
or U23080 (N_23080,N_18466,N_18493);
nand U23081 (N_23081,N_18462,N_15000);
xor U23082 (N_23082,N_19409,N_18581);
nand U23083 (N_23083,N_15308,N_19492);
nand U23084 (N_23084,N_17602,N_18474);
or U23085 (N_23085,N_15616,N_17664);
nor U23086 (N_23086,N_19847,N_16246);
xnor U23087 (N_23087,N_17826,N_15937);
or U23088 (N_23088,N_15070,N_19013);
nor U23089 (N_23089,N_17343,N_17891);
nor U23090 (N_23090,N_15955,N_17210);
or U23091 (N_23091,N_16086,N_17550);
xnor U23092 (N_23092,N_18491,N_15138);
or U23093 (N_23093,N_18056,N_19002);
or U23094 (N_23094,N_17887,N_16696);
nand U23095 (N_23095,N_17610,N_15758);
or U23096 (N_23096,N_15096,N_19120);
nor U23097 (N_23097,N_16922,N_16475);
or U23098 (N_23098,N_17018,N_15783);
or U23099 (N_23099,N_18342,N_18148);
and U23100 (N_23100,N_18954,N_18962);
nor U23101 (N_23101,N_17817,N_16438);
or U23102 (N_23102,N_15617,N_16242);
nand U23103 (N_23103,N_18539,N_18154);
nor U23104 (N_23104,N_18688,N_19725);
nor U23105 (N_23105,N_19560,N_16076);
xor U23106 (N_23106,N_19255,N_19838);
and U23107 (N_23107,N_18477,N_19742);
xnor U23108 (N_23108,N_15361,N_16683);
and U23109 (N_23109,N_18282,N_18041);
xnor U23110 (N_23110,N_16039,N_17824);
nand U23111 (N_23111,N_15190,N_15889);
nand U23112 (N_23112,N_18131,N_16656);
nand U23113 (N_23113,N_17795,N_18144);
and U23114 (N_23114,N_17572,N_17188);
and U23115 (N_23115,N_16942,N_16280);
nor U23116 (N_23116,N_19903,N_15038);
and U23117 (N_23117,N_16150,N_19075);
xor U23118 (N_23118,N_18012,N_19217);
or U23119 (N_23119,N_19424,N_18372);
or U23120 (N_23120,N_15998,N_17652);
nand U23121 (N_23121,N_19423,N_17102);
nor U23122 (N_23122,N_19838,N_15698);
xor U23123 (N_23123,N_18352,N_16537);
xnor U23124 (N_23124,N_18547,N_15848);
xor U23125 (N_23125,N_17838,N_17587);
nor U23126 (N_23126,N_17429,N_17951);
nand U23127 (N_23127,N_19556,N_18165);
or U23128 (N_23128,N_16196,N_18866);
xnor U23129 (N_23129,N_15613,N_18041);
nor U23130 (N_23130,N_16680,N_18500);
nand U23131 (N_23131,N_15756,N_16203);
nand U23132 (N_23132,N_19651,N_19601);
nor U23133 (N_23133,N_16797,N_15697);
nand U23134 (N_23134,N_17201,N_17899);
and U23135 (N_23135,N_16545,N_15879);
or U23136 (N_23136,N_16832,N_15377);
or U23137 (N_23137,N_17090,N_16721);
and U23138 (N_23138,N_17005,N_18791);
xnor U23139 (N_23139,N_16132,N_18642);
and U23140 (N_23140,N_19931,N_15856);
and U23141 (N_23141,N_18550,N_17857);
nand U23142 (N_23142,N_16569,N_19660);
nor U23143 (N_23143,N_19767,N_16178);
nand U23144 (N_23144,N_15151,N_15854);
nor U23145 (N_23145,N_19769,N_19931);
nand U23146 (N_23146,N_15452,N_16166);
and U23147 (N_23147,N_16678,N_16475);
or U23148 (N_23148,N_19352,N_15816);
and U23149 (N_23149,N_17583,N_16535);
xnor U23150 (N_23150,N_15315,N_17059);
nor U23151 (N_23151,N_17683,N_18961);
nor U23152 (N_23152,N_15404,N_15316);
or U23153 (N_23153,N_18723,N_15065);
and U23154 (N_23154,N_19952,N_18148);
nand U23155 (N_23155,N_19858,N_17928);
nor U23156 (N_23156,N_15151,N_15577);
nor U23157 (N_23157,N_19558,N_16978);
or U23158 (N_23158,N_15617,N_17394);
or U23159 (N_23159,N_15385,N_15819);
and U23160 (N_23160,N_16605,N_18544);
and U23161 (N_23161,N_15620,N_18524);
and U23162 (N_23162,N_17240,N_18186);
xor U23163 (N_23163,N_19857,N_19280);
nor U23164 (N_23164,N_19961,N_18141);
nand U23165 (N_23165,N_18612,N_16490);
nor U23166 (N_23166,N_19330,N_19513);
xnor U23167 (N_23167,N_19544,N_16932);
nor U23168 (N_23168,N_16179,N_17803);
or U23169 (N_23169,N_16732,N_16751);
nand U23170 (N_23170,N_18079,N_17621);
and U23171 (N_23171,N_15606,N_18334);
nand U23172 (N_23172,N_16789,N_15131);
nand U23173 (N_23173,N_16291,N_15501);
nor U23174 (N_23174,N_19291,N_19565);
or U23175 (N_23175,N_19767,N_16220);
and U23176 (N_23176,N_15106,N_18225);
nand U23177 (N_23177,N_16761,N_17709);
or U23178 (N_23178,N_18357,N_18280);
or U23179 (N_23179,N_16096,N_16491);
nand U23180 (N_23180,N_15887,N_16938);
nand U23181 (N_23181,N_18607,N_19538);
xor U23182 (N_23182,N_15432,N_19032);
or U23183 (N_23183,N_19040,N_17957);
or U23184 (N_23184,N_16350,N_19336);
or U23185 (N_23185,N_17465,N_18649);
nor U23186 (N_23186,N_15790,N_16401);
nand U23187 (N_23187,N_18823,N_19584);
nor U23188 (N_23188,N_19965,N_17237);
xnor U23189 (N_23189,N_17289,N_18563);
or U23190 (N_23190,N_16562,N_18592);
nand U23191 (N_23191,N_15071,N_18551);
and U23192 (N_23192,N_18380,N_15782);
nand U23193 (N_23193,N_16996,N_15144);
or U23194 (N_23194,N_17154,N_16110);
nor U23195 (N_23195,N_17963,N_19805);
and U23196 (N_23196,N_15946,N_16123);
nand U23197 (N_23197,N_17061,N_15779);
or U23198 (N_23198,N_19418,N_16235);
nand U23199 (N_23199,N_16629,N_17834);
and U23200 (N_23200,N_19235,N_18005);
and U23201 (N_23201,N_16465,N_15896);
and U23202 (N_23202,N_17910,N_17917);
or U23203 (N_23203,N_16838,N_18362);
nor U23204 (N_23204,N_15300,N_18377);
or U23205 (N_23205,N_19286,N_15849);
nand U23206 (N_23206,N_19956,N_17863);
nor U23207 (N_23207,N_19471,N_17171);
xor U23208 (N_23208,N_19551,N_15405);
or U23209 (N_23209,N_18250,N_16149);
or U23210 (N_23210,N_18857,N_15124);
or U23211 (N_23211,N_17249,N_19950);
or U23212 (N_23212,N_18744,N_17666);
nand U23213 (N_23213,N_19914,N_18448);
nor U23214 (N_23214,N_19859,N_19564);
xor U23215 (N_23215,N_17880,N_16965);
nor U23216 (N_23216,N_15587,N_19694);
nand U23217 (N_23217,N_17306,N_15035);
or U23218 (N_23218,N_17844,N_18128);
nor U23219 (N_23219,N_17719,N_16309);
nand U23220 (N_23220,N_19743,N_18121);
xnor U23221 (N_23221,N_15066,N_15933);
nor U23222 (N_23222,N_17168,N_16752);
nor U23223 (N_23223,N_18297,N_16593);
xnor U23224 (N_23224,N_16110,N_18860);
or U23225 (N_23225,N_19274,N_15395);
or U23226 (N_23226,N_19602,N_18250);
and U23227 (N_23227,N_19449,N_16375);
and U23228 (N_23228,N_17626,N_19222);
xor U23229 (N_23229,N_18188,N_19028);
nor U23230 (N_23230,N_17173,N_18543);
nor U23231 (N_23231,N_17720,N_15830);
xnor U23232 (N_23232,N_18273,N_19728);
nand U23233 (N_23233,N_19700,N_19752);
and U23234 (N_23234,N_15124,N_19145);
and U23235 (N_23235,N_19283,N_18651);
nor U23236 (N_23236,N_15453,N_17980);
and U23237 (N_23237,N_15579,N_15931);
xor U23238 (N_23238,N_15880,N_18243);
and U23239 (N_23239,N_19790,N_16318);
nand U23240 (N_23240,N_17782,N_15632);
and U23241 (N_23241,N_19402,N_16248);
nand U23242 (N_23242,N_17159,N_18274);
or U23243 (N_23243,N_19892,N_16006);
or U23244 (N_23244,N_18134,N_19054);
xor U23245 (N_23245,N_16637,N_15642);
xnor U23246 (N_23246,N_19897,N_17874);
and U23247 (N_23247,N_19005,N_18062);
and U23248 (N_23248,N_18669,N_16561);
nor U23249 (N_23249,N_18763,N_18316);
nor U23250 (N_23250,N_17899,N_15876);
nand U23251 (N_23251,N_18644,N_15039);
and U23252 (N_23252,N_18719,N_18457);
or U23253 (N_23253,N_16005,N_15611);
xor U23254 (N_23254,N_19821,N_19339);
or U23255 (N_23255,N_15480,N_19259);
nand U23256 (N_23256,N_15781,N_16035);
nor U23257 (N_23257,N_17878,N_15671);
nor U23258 (N_23258,N_15439,N_19295);
or U23259 (N_23259,N_15595,N_18276);
nor U23260 (N_23260,N_16040,N_17672);
xor U23261 (N_23261,N_19371,N_15658);
nor U23262 (N_23262,N_19921,N_17688);
nor U23263 (N_23263,N_15185,N_15496);
xnor U23264 (N_23264,N_19718,N_16671);
xor U23265 (N_23265,N_15946,N_19142);
xnor U23266 (N_23266,N_18434,N_17955);
xnor U23267 (N_23267,N_17131,N_15029);
nand U23268 (N_23268,N_16821,N_15991);
nand U23269 (N_23269,N_16318,N_18205);
or U23270 (N_23270,N_19993,N_16324);
nand U23271 (N_23271,N_19033,N_19540);
xnor U23272 (N_23272,N_17860,N_16571);
nor U23273 (N_23273,N_16800,N_19081);
xor U23274 (N_23274,N_16296,N_18065);
xnor U23275 (N_23275,N_15520,N_16717);
nand U23276 (N_23276,N_18891,N_19863);
or U23277 (N_23277,N_18791,N_16682);
and U23278 (N_23278,N_17268,N_19941);
xnor U23279 (N_23279,N_15213,N_19326);
or U23280 (N_23280,N_16157,N_16307);
and U23281 (N_23281,N_15063,N_16636);
nor U23282 (N_23282,N_17555,N_16511);
xnor U23283 (N_23283,N_16538,N_17088);
xnor U23284 (N_23284,N_17430,N_18333);
nor U23285 (N_23285,N_15775,N_15936);
and U23286 (N_23286,N_17514,N_17946);
or U23287 (N_23287,N_16882,N_15951);
nand U23288 (N_23288,N_18356,N_16983);
nor U23289 (N_23289,N_15341,N_15641);
nand U23290 (N_23290,N_16514,N_16725);
xnor U23291 (N_23291,N_15647,N_18642);
nand U23292 (N_23292,N_18723,N_18097);
nor U23293 (N_23293,N_19205,N_15036);
nand U23294 (N_23294,N_15136,N_17769);
nand U23295 (N_23295,N_16612,N_18672);
nand U23296 (N_23296,N_18504,N_16250);
and U23297 (N_23297,N_15788,N_19196);
xor U23298 (N_23298,N_19821,N_19017);
nor U23299 (N_23299,N_16442,N_17872);
xnor U23300 (N_23300,N_15626,N_18357);
xor U23301 (N_23301,N_16261,N_19021);
xor U23302 (N_23302,N_19387,N_18838);
nor U23303 (N_23303,N_19641,N_19212);
or U23304 (N_23304,N_18917,N_15263);
xor U23305 (N_23305,N_15053,N_17478);
or U23306 (N_23306,N_15975,N_18265);
xor U23307 (N_23307,N_18950,N_16638);
xor U23308 (N_23308,N_16485,N_15053);
or U23309 (N_23309,N_17825,N_16531);
nor U23310 (N_23310,N_16621,N_19902);
and U23311 (N_23311,N_17335,N_19558);
and U23312 (N_23312,N_17947,N_17337);
nor U23313 (N_23313,N_17894,N_18056);
xor U23314 (N_23314,N_16333,N_15211);
and U23315 (N_23315,N_19944,N_18074);
and U23316 (N_23316,N_17932,N_16509);
nand U23317 (N_23317,N_15701,N_19683);
nor U23318 (N_23318,N_18089,N_15390);
nor U23319 (N_23319,N_18810,N_17582);
nor U23320 (N_23320,N_19116,N_16426);
nor U23321 (N_23321,N_19766,N_15934);
xor U23322 (N_23322,N_17843,N_17246);
nand U23323 (N_23323,N_19170,N_17750);
or U23324 (N_23324,N_17755,N_18068);
xnor U23325 (N_23325,N_16181,N_15393);
or U23326 (N_23326,N_19563,N_16958);
nand U23327 (N_23327,N_19467,N_15272);
or U23328 (N_23328,N_16510,N_18434);
or U23329 (N_23329,N_16717,N_15544);
or U23330 (N_23330,N_15126,N_17151);
xor U23331 (N_23331,N_19697,N_16379);
or U23332 (N_23332,N_19431,N_15041);
nor U23333 (N_23333,N_19373,N_19215);
nor U23334 (N_23334,N_18551,N_16778);
or U23335 (N_23335,N_17824,N_15776);
xnor U23336 (N_23336,N_17312,N_17444);
and U23337 (N_23337,N_18394,N_16277);
nor U23338 (N_23338,N_18929,N_15767);
nand U23339 (N_23339,N_19820,N_16298);
nor U23340 (N_23340,N_17653,N_17146);
nand U23341 (N_23341,N_18573,N_15269);
xnor U23342 (N_23342,N_15909,N_15955);
xnor U23343 (N_23343,N_19605,N_18780);
nor U23344 (N_23344,N_19221,N_16609);
or U23345 (N_23345,N_19149,N_15227);
nand U23346 (N_23346,N_19895,N_15425);
nor U23347 (N_23347,N_16506,N_19654);
or U23348 (N_23348,N_16927,N_15317);
or U23349 (N_23349,N_16186,N_15160);
nand U23350 (N_23350,N_17622,N_16209);
or U23351 (N_23351,N_18407,N_19566);
or U23352 (N_23352,N_17561,N_19960);
nor U23353 (N_23353,N_15169,N_18699);
or U23354 (N_23354,N_17830,N_16454);
or U23355 (N_23355,N_17225,N_18943);
xor U23356 (N_23356,N_17543,N_19464);
and U23357 (N_23357,N_19242,N_17084);
or U23358 (N_23358,N_19185,N_18600);
or U23359 (N_23359,N_16742,N_18030);
nand U23360 (N_23360,N_16612,N_19326);
xor U23361 (N_23361,N_19943,N_18039);
nor U23362 (N_23362,N_18846,N_17831);
nand U23363 (N_23363,N_16498,N_19760);
and U23364 (N_23364,N_16087,N_18460);
nand U23365 (N_23365,N_17659,N_18594);
xor U23366 (N_23366,N_18895,N_18233);
or U23367 (N_23367,N_15059,N_15816);
nand U23368 (N_23368,N_18044,N_15587);
and U23369 (N_23369,N_16521,N_18749);
xor U23370 (N_23370,N_19057,N_17123);
xnor U23371 (N_23371,N_15400,N_16810);
or U23372 (N_23372,N_17894,N_18110);
and U23373 (N_23373,N_15245,N_16415);
nand U23374 (N_23374,N_17667,N_16499);
and U23375 (N_23375,N_19048,N_17702);
nor U23376 (N_23376,N_18562,N_16260);
xnor U23377 (N_23377,N_15203,N_19288);
or U23378 (N_23378,N_17781,N_15174);
nor U23379 (N_23379,N_18650,N_16600);
nand U23380 (N_23380,N_17954,N_15104);
nor U23381 (N_23381,N_19157,N_15438);
nand U23382 (N_23382,N_16427,N_16841);
nor U23383 (N_23383,N_19721,N_19463);
nand U23384 (N_23384,N_15157,N_17123);
or U23385 (N_23385,N_15805,N_18725);
xor U23386 (N_23386,N_18508,N_16317);
nor U23387 (N_23387,N_15634,N_15978);
or U23388 (N_23388,N_17846,N_19304);
and U23389 (N_23389,N_18295,N_18669);
nor U23390 (N_23390,N_17394,N_15734);
nand U23391 (N_23391,N_19260,N_17698);
and U23392 (N_23392,N_15260,N_16240);
xor U23393 (N_23393,N_17349,N_15713);
xnor U23394 (N_23394,N_18803,N_15117);
xnor U23395 (N_23395,N_16860,N_18192);
or U23396 (N_23396,N_19397,N_18463);
and U23397 (N_23397,N_15286,N_16288);
xnor U23398 (N_23398,N_16401,N_16310);
nand U23399 (N_23399,N_15151,N_18589);
and U23400 (N_23400,N_16188,N_15983);
and U23401 (N_23401,N_15831,N_18004);
or U23402 (N_23402,N_16070,N_18800);
nand U23403 (N_23403,N_16693,N_19729);
xor U23404 (N_23404,N_19039,N_16037);
nand U23405 (N_23405,N_18664,N_16185);
and U23406 (N_23406,N_16212,N_19416);
xor U23407 (N_23407,N_15306,N_15910);
nor U23408 (N_23408,N_18933,N_19572);
nor U23409 (N_23409,N_17811,N_15210);
or U23410 (N_23410,N_19021,N_18484);
nor U23411 (N_23411,N_15055,N_18493);
xnor U23412 (N_23412,N_17138,N_18542);
xor U23413 (N_23413,N_16471,N_16325);
xor U23414 (N_23414,N_15790,N_19182);
nor U23415 (N_23415,N_17802,N_15369);
and U23416 (N_23416,N_19084,N_15878);
nand U23417 (N_23417,N_18872,N_15202);
nor U23418 (N_23418,N_19125,N_17644);
nor U23419 (N_23419,N_17159,N_18666);
xor U23420 (N_23420,N_18825,N_15248);
or U23421 (N_23421,N_17069,N_19853);
and U23422 (N_23422,N_19708,N_19655);
nand U23423 (N_23423,N_17724,N_19850);
nor U23424 (N_23424,N_15828,N_19001);
nand U23425 (N_23425,N_16829,N_15684);
and U23426 (N_23426,N_15639,N_19276);
and U23427 (N_23427,N_19229,N_18195);
or U23428 (N_23428,N_19728,N_16673);
nand U23429 (N_23429,N_15930,N_16626);
xor U23430 (N_23430,N_16797,N_19353);
nand U23431 (N_23431,N_17823,N_19301);
or U23432 (N_23432,N_18220,N_16279);
and U23433 (N_23433,N_19574,N_17629);
nor U23434 (N_23434,N_17658,N_19905);
xor U23435 (N_23435,N_18833,N_17649);
and U23436 (N_23436,N_17415,N_15404);
nand U23437 (N_23437,N_18564,N_16083);
nand U23438 (N_23438,N_16280,N_18036);
nor U23439 (N_23439,N_15709,N_19877);
xnor U23440 (N_23440,N_19094,N_19078);
nor U23441 (N_23441,N_17225,N_19077);
nor U23442 (N_23442,N_19590,N_15546);
nand U23443 (N_23443,N_19045,N_19489);
xnor U23444 (N_23444,N_15839,N_17143);
nor U23445 (N_23445,N_18571,N_15998);
nand U23446 (N_23446,N_15522,N_16529);
and U23447 (N_23447,N_15120,N_16838);
or U23448 (N_23448,N_19979,N_16618);
and U23449 (N_23449,N_17787,N_18432);
xnor U23450 (N_23450,N_19833,N_16609);
nor U23451 (N_23451,N_17701,N_16847);
and U23452 (N_23452,N_17382,N_19748);
nand U23453 (N_23453,N_17894,N_15687);
xor U23454 (N_23454,N_18165,N_15859);
or U23455 (N_23455,N_16418,N_19789);
nor U23456 (N_23456,N_17646,N_15260);
or U23457 (N_23457,N_19042,N_15705);
or U23458 (N_23458,N_16264,N_15451);
xor U23459 (N_23459,N_19190,N_19961);
xnor U23460 (N_23460,N_19318,N_15547);
xnor U23461 (N_23461,N_17011,N_16338);
and U23462 (N_23462,N_19879,N_16470);
and U23463 (N_23463,N_19434,N_19387);
nor U23464 (N_23464,N_17197,N_15128);
or U23465 (N_23465,N_17058,N_17831);
and U23466 (N_23466,N_16726,N_19764);
nor U23467 (N_23467,N_17850,N_18185);
nor U23468 (N_23468,N_16924,N_16214);
xnor U23469 (N_23469,N_18915,N_17064);
and U23470 (N_23470,N_18141,N_19300);
nand U23471 (N_23471,N_16952,N_17081);
xnor U23472 (N_23472,N_15710,N_15607);
nor U23473 (N_23473,N_17165,N_15945);
nor U23474 (N_23474,N_17850,N_16373);
xnor U23475 (N_23475,N_16678,N_17978);
and U23476 (N_23476,N_17404,N_17998);
or U23477 (N_23477,N_18858,N_17279);
nand U23478 (N_23478,N_16989,N_17584);
or U23479 (N_23479,N_17999,N_18935);
and U23480 (N_23480,N_16145,N_17122);
or U23481 (N_23481,N_17257,N_18894);
nand U23482 (N_23482,N_17608,N_16286);
and U23483 (N_23483,N_17567,N_17349);
or U23484 (N_23484,N_15100,N_16224);
or U23485 (N_23485,N_17351,N_19607);
nand U23486 (N_23486,N_16886,N_18606);
nor U23487 (N_23487,N_18453,N_18860);
or U23488 (N_23488,N_17777,N_19031);
or U23489 (N_23489,N_19336,N_16334);
xnor U23490 (N_23490,N_17601,N_17270);
nand U23491 (N_23491,N_19499,N_19529);
or U23492 (N_23492,N_19868,N_17685);
nor U23493 (N_23493,N_17016,N_17305);
or U23494 (N_23494,N_16361,N_15159);
xor U23495 (N_23495,N_16891,N_18978);
and U23496 (N_23496,N_18480,N_17141);
or U23497 (N_23497,N_16581,N_17119);
nand U23498 (N_23498,N_18896,N_19392);
nand U23499 (N_23499,N_15183,N_15116);
xnor U23500 (N_23500,N_15739,N_16097);
nor U23501 (N_23501,N_17059,N_17639);
nor U23502 (N_23502,N_18073,N_19131);
nand U23503 (N_23503,N_19267,N_18275);
and U23504 (N_23504,N_19303,N_19454);
or U23505 (N_23505,N_19515,N_15469);
or U23506 (N_23506,N_16429,N_18321);
or U23507 (N_23507,N_17254,N_17897);
and U23508 (N_23508,N_18012,N_19620);
or U23509 (N_23509,N_17922,N_15064);
nor U23510 (N_23510,N_18967,N_16899);
nand U23511 (N_23511,N_17990,N_18429);
nor U23512 (N_23512,N_18712,N_19757);
or U23513 (N_23513,N_17843,N_18448);
xor U23514 (N_23514,N_19762,N_17287);
nand U23515 (N_23515,N_15779,N_15328);
nor U23516 (N_23516,N_17081,N_18455);
nor U23517 (N_23517,N_19680,N_18231);
or U23518 (N_23518,N_17094,N_19486);
nand U23519 (N_23519,N_16327,N_17773);
nor U23520 (N_23520,N_18905,N_18650);
nand U23521 (N_23521,N_19467,N_17294);
xnor U23522 (N_23522,N_17460,N_17677);
nor U23523 (N_23523,N_16410,N_19003);
or U23524 (N_23524,N_17397,N_19596);
nor U23525 (N_23525,N_19263,N_17429);
and U23526 (N_23526,N_17053,N_16033);
xor U23527 (N_23527,N_19101,N_19434);
nor U23528 (N_23528,N_15893,N_15436);
and U23529 (N_23529,N_15588,N_16999);
nor U23530 (N_23530,N_16896,N_19930);
xor U23531 (N_23531,N_16815,N_16430);
or U23532 (N_23532,N_15315,N_18026);
xnor U23533 (N_23533,N_15198,N_18789);
or U23534 (N_23534,N_19473,N_18551);
and U23535 (N_23535,N_15998,N_19825);
nand U23536 (N_23536,N_17586,N_18075);
and U23537 (N_23537,N_17709,N_18875);
nor U23538 (N_23538,N_15266,N_17003);
and U23539 (N_23539,N_16302,N_19336);
nand U23540 (N_23540,N_19586,N_16817);
and U23541 (N_23541,N_17808,N_17991);
nor U23542 (N_23542,N_18748,N_16354);
or U23543 (N_23543,N_17524,N_16132);
and U23544 (N_23544,N_18211,N_15941);
nand U23545 (N_23545,N_19014,N_15788);
and U23546 (N_23546,N_15129,N_17470);
or U23547 (N_23547,N_19824,N_19318);
or U23548 (N_23548,N_17844,N_16667);
and U23549 (N_23549,N_17108,N_17404);
or U23550 (N_23550,N_16374,N_16899);
or U23551 (N_23551,N_16286,N_19611);
nand U23552 (N_23552,N_19631,N_15580);
nand U23553 (N_23553,N_18827,N_17839);
xor U23554 (N_23554,N_15943,N_18728);
xnor U23555 (N_23555,N_19704,N_15202);
nand U23556 (N_23556,N_15966,N_16057);
or U23557 (N_23557,N_19207,N_18970);
or U23558 (N_23558,N_17427,N_16423);
xor U23559 (N_23559,N_16421,N_17079);
or U23560 (N_23560,N_18079,N_17374);
and U23561 (N_23561,N_16432,N_15812);
nor U23562 (N_23562,N_15267,N_18076);
xnor U23563 (N_23563,N_19548,N_19175);
xnor U23564 (N_23564,N_15296,N_17424);
xnor U23565 (N_23565,N_16754,N_16063);
and U23566 (N_23566,N_16980,N_16184);
nor U23567 (N_23567,N_17013,N_15867);
nand U23568 (N_23568,N_17715,N_16975);
or U23569 (N_23569,N_19564,N_18804);
nor U23570 (N_23570,N_18729,N_19310);
or U23571 (N_23571,N_15838,N_17614);
nor U23572 (N_23572,N_16059,N_17825);
and U23573 (N_23573,N_19400,N_15204);
and U23574 (N_23574,N_16903,N_19626);
xnor U23575 (N_23575,N_19492,N_16254);
xnor U23576 (N_23576,N_18189,N_16544);
nand U23577 (N_23577,N_16370,N_15500);
or U23578 (N_23578,N_16044,N_16717);
or U23579 (N_23579,N_18704,N_16622);
or U23580 (N_23580,N_15547,N_18714);
nor U23581 (N_23581,N_15674,N_16708);
nor U23582 (N_23582,N_19782,N_15570);
or U23583 (N_23583,N_16979,N_17587);
or U23584 (N_23584,N_19765,N_15881);
or U23585 (N_23585,N_15065,N_18515);
xnor U23586 (N_23586,N_16895,N_19416);
and U23587 (N_23587,N_16331,N_16499);
xor U23588 (N_23588,N_19394,N_18437);
nor U23589 (N_23589,N_15714,N_19614);
and U23590 (N_23590,N_18740,N_19020);
xor U23591 (N_23591,N_15621,N_17136);
and U23592 (N_23592,N_19296,N_16844);
or U23593 (N_23593,N_17450,N_15763);
nor U23594 (N_23594,N_17855,N_17342);
and U23595 (N_23595,N_17471,N_17981);
nand U23596 (N_23596,N_16722,N_17307);
or U23597 (N_23597,N_17482,N_17337);
or U23598 (N_23598,N_15044,N_18523);
nand U23599 (N_23599,N_15526,N_16912);
xnor U23600 (N_23600,N_17212,N_15234);
and U23601 (N_23601,N_19377,N_18208);
nand U23602 (N_23602,N_16915,N_18044);
or U23603 (N_23603,N_16965,N_15115);
nand U23604 (N_23604,N_16823,N_16447);
nor U23605 (N_23605,N_18720,N_17653);
and U23606 (N_23606,N_19349,N_19198);
xor U23607 (N_23607,N_17950,N_19948);
xnor U23608 (N_23608,N_18962,N_18765);
or U23609 (N_23609,N_19099,N_18066);
nand U23610 (N_23610,N_17385,N_17287);
or U23611 (N_23611,N_15781,N_18076);
and U23612 (N_23612,N_19563,N_17316);
and U23613 (N_23613,N_17875,N_18335);
nand U23614 (N_23614,N_18471,N_15804);
and U23615 (N_23615,N_19884,N_18165);
or U23616 (N_23616,N_18947,N_16573);
xnor U23617 (N_23617,N_16173,N_17228);
or U23618 (N_23618,N_17624,N_15972);
nand U23619 (N_23619,N_16797,N_18600);
nor U23620 (N_23620,N_17870,N_17863);
nor U23621 (N_23621,N_17538,N_19532);
and U23622 (N_23622,N_16627,N_16931);
nand U23623 (N_23623,N_15357,N_19467);
or U23624 (N_23624,N_17930,N_19355);
and U23625 (N_23625,N_15764,N_15831);
nand U23626 (N_23626,N_15176,N_19640);
or U23627 (N_23627,N_16023,N_18643);
xnor U23628 (N_23628,N_16342,N_19981);
or U23629 (N_23629,N_19194,N_18102);
nand U23630 (N_23630,N_18081,N_15026);
nor U23631 (N_23631,N_18228,N_17977);
and U23632 (N_23632,N_19635,N_16491);
xor U23633 (N_23633,N_18838,N_19315);
xor U23634 (N_23634,N_17728,N_19034);
nor U23635 (N_23635,N_17039,N_17271);
nor U23636 (N_23636,N_15106,N_16446);
xor U23637 (N_23637,N_17813,N_16131);
or U23638 (N_23638,N_17039,N_16628);
nor U23639 (N_23639,N_18197,N_16421);
nor U23640 (N_23640,N_19974,N_16658);
nor U23641 (N_23641,N_16769,N_15336);
and U23642 (N_23642,N_16072,N_18974);
xor U23643 (N_23643,N_15801,N_15105);
nand U23644 (N_23644,N_18041,N_19065);
nor U23645 (N_23645,N_19640,N_15237);
and U23646 (N_23646,N_16929,N_17337);
nor U23647 (N_23647,N_16761,N_17434);
xnor U23648 (N_23648,N_17171,N_18150);
nand U23649 (N_23649,N_16650,N_17677);
nand U23650 (N_23650,N_16856,N_16610);
or U23651 (N_23651,N_18553,N_16948);
and U23652 (N_23652,N_17812,N_17349);
and U23653 (N_23653,N_17491,N_17793);
nand U23654 (N_23654,N_18104,N_19712);
or U23655 (N_23655,N_16156,N_18197);
xnor U23656 (N_23656,N_15460,N_17323);
or U23657 (N_23657,N_18001,N_16669);
nor U23658 (N_23658,N_19452,N_19073);
nor U23659 (N_23659,N_17575,N_16039);
or U23660 (N_23660,N_18708,N_18830);
nand U23661 (N_23661,N_17503,N_15623);
nor U23662 (N_23662,N_15438,N_15733);
and U23663 (N_23663,N_18913,N_15274);
or U23664 (N_23664,N_15519,N_18322);
xnor U23665 (N_23665,N_17722,N_16305);
nand U23666 (N_23666,N_17314,N_19320);
nor U23667 (N_23667,N_16536,N_16912);
or U23668 (N_23668,N_19596,N_17884);
or U23669 (N_23669,N_16804,N_18518);
xnor U23670 (N_23670,N_19661,N_16714);
xnor U23671 (N_23671,N_15121,N_19638);
and U23672 (N_23672,N_18103,N_17992);
xor U23673 (N_23673,N_15991,N_15434);
nor U23674 (N_23674,N_18961,N_18957);
nor U23675 (N_23675,N_15581,N_17836);
or U23676 (N_23676,N_16461,N_15360);
or U23677 (N_23677,N_17984,N_19985);
or U23678 (N_23678,N_16125,N_16530);
xnor U23679 (N_23679,N_17964,N_18191);
nor U23680 (N_23680,N_18856,N_19902);
nand U23681 (N_23681,N_19345,N_18576);
or U23682 (N_23682,N_19498,N_16520);
xnor U23683 (N_23683,N_15750,N_19244);
nand U23684 (N_23684,N_18026,N_19434);
nor U23685 (N_23685,N_19621,N_16123);
nand U23686 (N_23686,N_18090,N_17460);
or U23687 (N_23687,N_16900,N_18772);
xnor U23688 (N_23688,N_17885,N_17040);
or U23689 (N_23689,N_17235,N_18669);
xor U23690 (N_23690,N_17432,N_17001);
or U23691 (N_23691,N_16574,N_15126);
nor U23692 (N_23692,N_15662,N_15864);
xor U23693 (N_23693,N_19474,N_17824);
xor U23694 (N_23694,N_16094,N_19423);
and U23695 (N_23695,N_17467,N_19959);
nor U23696 (N_23696,N_19917,N_17972);
xor U23697 (N_23697,N_15461,N_19365);
nand U23698 (N_23698,N_16094,N_18352);
nor U23699 (N_23699,N_17689,N_16820);
nand U23700 (N_23700,N_16730,N_15620);
xnor U23701 (N_23701,N_19291,N_19040);
or U23702 (N_23702,N_18464,N_18968);
nor U23703 (N_23703,N_16256,N_18912);
xor U23704 (N_23704,N_19883,N_18290);
xor U23705 (N_23705,N_18014,N_15000);
nand U23706 (N_23706,N_19293,N_18581);
xor U23707 (N_23707,N_17053,N_17544);
and U23708 (N_23708,N_18983,N_18793);
or U23709 (N_23709,N_15291,N_19207);
nand U23710 (N_23710,N_15868,N_19626);
and U23711 (N_23711,N_15811,N_19521);
and U23712 (N_23712,N_15480,N_17063);
nand U23713 (N_23713,N_19753,N_18340);
or U23714 (N_23714,N_17597,N_17570);
and U23715 (N_23715,N_15082,N_16374);
xnor U23716 (N_23716,N_18820,N_16115);
or U23717 (N_23717,N_17749,N_16333);
or U23718 (N_23718,N_15722,N_17209);
xor U23719 (N_23719,N_15058,N_19375);
xnor U23720 (N_23720,N_19077,N_15467);
and U23721 (N_23721,N_18735,N_17777);
nor U23722 (N_23722,N_19905,N_19695);
xnor U23723 (N_23723,N_17333,N_15335);
xor U23724 (N_23724,N_15715,N_18926);
or U23725 (N_23725,N_19534,N_16997);
nor U23726 (N_23726,N_15450,N_19024);
and U23727 (N_23727,N_19028,N_16780);
nand U23728 (N_23728,N_19345,N_16954);
or U23729 (N_23729,N_16213,N_15757);
nand U23730 (N_23730,N_18666,N_18936);
xnor U23731 (N_23731,N_15960,N_18328);
nor U23732 (N_23732,N_16317,N_15553);
xor U23733 (N_23733,N_15986,N_18910);
nand U23734 (N_23734,N_19114,N_19201);
xnor U23735 (N_23735,N_17089,N_15260);
nand U23736 (N_23736,N_18704,N_15170);
nor U23737 (N_23737,N_18401,N_19762);
xor U23738 (N_23738,N_17298,N_17169);
and U23739 (N_23739,N_17615,N_15278);
nor U23740 (N_23740,N_17345,N_16983);
nor U23741 (N_23741,N_19619,N_16219);
and U23742 (N_23742,N_18839,N_18508);
xor U23743 (N_23743,N_19781,N_18908);
or U23744 (N_23744,N_19476,N_19392);
nand U23745 (N_23745,N_16382,N_16990);
xor U23746 (N_23746,N_18672,N_16045);
xor U23747 (N_23747,N_18153,N_18768);
and U23748 (N_23748,N_18110,N_19003);
and U23749 (N_23749,N_19701,N_16690);
xor U23750 (N_23750,N_17338,N_19880);
nor U23751 (N_23751,N_19382,N_16806);
xor U23752 (N_23752,N_19432,N_15245);
or U23753 (N_23753,N_15734,N_16757);
or U23754 (N_23754,N_15703,N_17748);
nor U23755 (N_23755,N_15998,N_18624);
nand U23756 (N_23756,N_17167,N_15936);
and U23757 (N_23757,N_19464,N_17709);
and U23758 (N_23758,N_18569,N_19404);
or U23759 (N_23759,N_18005,N_16555);
xnor U23760 (N_23760,N_15864,N_19602);
and U23761 (N_23761,N_19279,N_16061);
and U23762 (N_23762,N_15879,N_16822);
or U23763 (N_23763,N_19121,N_19793);
or U23764 (N_23764,N_17040,N_16862);
nand U23765 (N_23765,N_18044,N_16320);
or U23766 (N_23766,N_16488,N_19895);
or U23767 (N_23767,N_19593,N_19146);
nor U23768 (N_23768,N_16402,N_16117);
xnor U23769 (N_23769,N_18804,N_19602);
or U23770 (N_23770,N_19316,N_17379);
or U23771 (N_23771,N_15068,N_17705);
xnor U23772 (N_23772,N_16566,N_19257);
nor U23773 (N_23773,N_19590,N_17916);
nand U23774 (N_23774,N_18089,N_18341);
and U23775 (N_23775,N_19839,N_18276);
and U23776 (N_23776,N_16711,N_19148);
xor U23777 (N_23777,N_17814,N_19109);
nand U23778 (N_23778,N_18479,N_18943);
and U23779 (N_23779,N_18729,N_17652);
xor U23780 (N_23780,N_15029,N_19386);
or U23781 (N_23781,N_17034,N_15031);
xor U23782 (N_23782,N_18498,N_19960);
and U23783 (N_23783,N_18578,N_19284);
or U23784 (N_23784,N_17084,N_17719);
or U23785 (N_23785,N_16420,N_19474);
nand U23786 (N_23786,N_18270,N_19214);
nor U23787 (N_23787,N_18967,N_15572);
or U23788 (N_23788,N_18363,N_18729);
nor U23789 (N_23789,N_19377,N_17238);
or U23790 (N_23790,N_16080,N_19154);
nand U23791 (N_23791,N_19772,N_19658);
or U23792 (N_23792,N_16312,N_17392);
nand U23793 (N_23793,N_19802,N_18534);
or U23794 (N_23794,N_19731,N_19322);
nor U23795 (N_23795,N_18498,N_17688);
nor U23796 (N_23796,N_19154,N_18108);
nand U23797 (N_23797,N_19959,N_18195);
nor U23798 (N_23798,N_15661,N_18362);
and U23799 (N_23799,N_18273,N_19383);
xnor U23800 (N_23800,N_17915,N_17841);
nor U23801 (N_23801,N_17820,N_15693);
xnor U23802 (N_23802,N_15135,N_18968);
and U23803 (N_23803,N_15715,N_19766);
nor U23804 (N_23804,N_17676,N_16965);
and U23805 (N_23805,N_15046,N_19831);
nand U23806 (N_23806,N_19105,N_18842);
nand U23807 (N_23807,N_18655,N_17239);
nand U23808 (N_23808,N_18720,N_16116);
nor U23809 (N_23809,N_19192,N_18219);
nor U23810 (N_23810,N_17914,N_18019);
and U23811 (N_23811,N_16923,N_19049);
nand U23812 (N_23812,N_16777,N_17001);
nor U23813 (N_23813,N_17873,N_17920);
nand U23814 (N_23814,N_17183,N_15154);
nand U23815 (N_23815,N_15396,N_15365);
xor U23816 (N_23816,N_17823,N_15296);
nor U23817 (N_23817,N_17084,N_17146);
nor U23818 (N_23818,N_18268,N_19871);
xor U23819 (N_23819,N_17295,N_17305);
and U23820 (N_23820,N_16533,N_17770);
nand U23821 (N_23821,N_15248,N_18772);
xnor U23822 (N_23822,N_18368,N_18468);
nand U23823 (N_23823,N_15350,N_15446);
and U23824 (N_23824,N_18779,N_15484);
xor U23825 (N_23825,N_19860,N_16414);
nor U23826 (N_23826,N_16606,N_16096);
nand U23827 (N_23827,N_15367,N_18625);
xnor U23828 (N_23828,N_15558,N_15880);
nand U23829 (N_23829,N_16571,N_16400);
and U23830 (N_23830,N_15359,N_16054);
nor U23831 (N_23831,N_16050,N_16030);
xor U23832 (N_23832,N_19713,N_16395);
xor U23833 (N_23833,N_17826,N_17729);
xnor U23834 (N_23834,N_17319,N_15274);
and U23835 (N_23835,N_16138,N_16358);
xnor U23836 (N_23836,N_16807,N_16046);
nor U23837 (N_23837,N_16998,N_19937);
nor U23838 (N_23838,N_16980,N_19136);
nor U23839 (N_23839,N_19089,N_18172);
and U23840 (N_23840,N_19241,N_18706);
nand U23841 (N_23841,N_15688,N_19074);
xnor U23842 (N_23842,N_16756,N_15750);
xor U23843 (N_23843,N_18658,N_16769);
xnor U23844 (N_23844,N_16116,N_18022);
and U23845 (N_23845,N_17953,N_18676);
or U23846 (N_23846,N_16601,N_15015);
xnor U23847 (N_23847,N_18281,N_18452);
nand U23848 (N_23848,N_19573,N_19727);
or U23849 (N_23849,N_18259,N_17121);
xnor U23850 (N_23850,N_17826,N_19866);
xor U23851 (N_23851,N_17257,N_17797);
and U23852 (N_23852,N_16242,N_19545);
nand U23853 (N_23853,N_17406,N_16292);
and U23854 (N_23854,N_16516,N_19642);
and U23855 (N_23855,N_16565,N_19650);
nor U23856 (N_23856,N_15768,N_15022);
nand U23857 (N_23857,N_15982,N_19267);
nand U23858 (N_23858,N_15166,N_17001);
or U23859 (N_23859,N_17537,N_16743);
and U23860 (N_23860,N_15558,N_18525);
nand U23861 (N_23861,N_19320,N_19890);
xor U23862 (N_23862,N_15411,N_17331);
and U23863 (N_23863,N_19833,N_17322);
or U23864 (N_23864,N_15612,N_16079);
and U23865 (N_23865,N_18035,N_18963);
nand U23866 (N_23866,N_15114,N_15301);
and U23867 (N_23867,N_18680,N_18599);
and U23868 (N_23868,N_19706,N_18649);
and U23869 (N_23869,N_19964,N_17194);
nand U23870 (N_23870,N_17569,N_15931);
nor U23871 (N_23871,N_19193,N_18260);
or U23872 (N_23872,N_19270,N_16718);
and U23873 (N_23873,N_15309,N_18357);
and U23874 (N_23874,N_18226,N_15830);
nor U23875 (N_23875,N_19892,N_19483);
nor U23876 (N_23876,N_18347,N_15792);
and U23877 (N_23877,N_15069,N_17446);
xor U23878 (N_23878,N_16406,N_15604);
and U23879 (N_23879,N_17987,N_19092);
xor U23880 (N_23880,N_15619,N_19189);
nand U23881 (N_23881,N_17639,N_17001);
xor U23882 (N_23882,N_16811,N_16863);
nand U23883 (N_23883,N_15596,N_15323);
or U23884 (N_23884,N_18548,N_15289);
and U23885 (N_23885,N_18883,N_16961);
and U23886 (N_23886,N_15882,N_16651);
and U23887 (N_23887,N_17993,N_17920);
nand U23888 (N_23888,N_15016,N_16134);
or U23889 (N_23889,N_19371,N_17149);
xnor U23890 (N_23890,N_19554,N_17241);
or U23891 (N_23891,N_16665,N_18641);
nand U23892 (N_23892,N_16265,N_19304);
xor U23893 (N_23893,N_18249,N_19538);
nor U23894 (N_23894,N_19925,N_17540);
and U23895 (N_23895,N_16872,N_15403);
xor U23896 (N_23896,N_15911,N_18180);
or U23897 (N_23897,N_16029,N_18369);
or U23898 (N_23898,N_18108,N_19992);
xnor U23899 (N_23899,N_18900,N_19188);
xor U23900 (N_23900,N_18161,N_16895);
and U23901 (N_23901,N_17718,N_18960);
nor U23902 (N_23902,N_17054,N_18287);
xor U23903 (N_23903,N_19199,N_16971);
xor U23904 (N_23904,N_17025,N_18619);
and U23905 (N_23905,N_17732,N_15506);
nor U23906 (N_23906,N_16653,N_19789);
nor U23907 (N_23907,N_17387,N_17993);
nand U23908 (N_23908,N_17802,N_18638);
nand U23909 (N_23909,N_17682,N_18423);
or U23910 (N_23910,N_15103,N_15074);
xnor U23911 (N_23911,N_18460,N_18425);
nand U23912 (N_23912,N_16002,N_18944);
nand U23913 (N_23913,N_16094,N_19143);
nor U23914 (N_23914,N_19232,N_17269);
xnor U23915 (N_23915,N_15318,N_15952);
or U23916 (N_23916,N_16916,N_18539);
nand U23917 (N_23917,N_16951,N_19297);
xor U23918 (N_23918,N_19424,N_15113);
xnor U23919 (N_23919,N_18647,N_19212);
nor U23920 (N_23920,N_18386,N_19319);
and U23921 (N_23921,N_15226,N_18480);
xor U23922 (N_23922,N_15528,N_17378);
or U23923 (N_23923,N_15618,N_19235);
xnor U23924 (N_23924,N_18623,N_17381);
nand U23925 (N_23925,N_17366,N_16794);
xnor U23926 (N_23926,N_18998,N_19553);
and U23927 (N_23927,N_16998,N_18980);
xor U23928 (N_23928,N_18630,N_16204);
or U23929 (N_23929,N_16883,N_16744);
nor U23930 (N_23930,N_16647,N_15260);
xor U23931 (N_23931,N_19279,N_19186);
and U23932 (N_23932,N_17538,N_15723);
and U23933 (N_23933,N_17087,N_15490);
xor U23934 (N_23934,N_15815,N_16269);
or U23935 (N_23935,N_17919,N_19969);
or U23936 (N_23936,N_18403,N_17639);
nand U23937 (N_23937,N_18674,N_18883);
and U23938 (N_23938,N_15885,N_15136);
nor U23939 (N_23939,N_15983,N_19941);
or U23940 (N_23940,N_19134,N_18905);
nor U23941 (N_23941,N_19499,N_18186);
and U23942 (N_23942,N_19761,N_15697);
xor U23943 (N_23943,N_16701,N_17657);
and U23944 (N_23944,N_15689,N_18878);
xnor U23945 (N_23945,N_16385,N_19694);
and U23946 (N_23946,N_17344,N_16202);
nand U23947 (N_23947,N_16120,N_17759);
xnor U23948 (N_23948,N_17273,N_18497);
or U23949 (N_23949,N_17537,N_16854);
xor U23950 (N_23950,N_19477,N_15027);
and U23951 (N_23951,N_19155,N_16288);
or U23952 (N_23952,N_17456,N_16364);
xor U23953 (N_23953,N_19151,N_18455);
nand U23954 (N_23954,N_19083,N_18202);
xnor U23955 (N_23955,N_18625,N_15646);
nand U23956 (N_23956,N_17841,N_19057);
xor U23957 (N_23957,N_15439,N_15827);
or U23958 (N_23958,N_18473,N_15571);
xnor U23959 (N_23959,N_16101,N_18734);
nor U23960 (N_23960,N_15835,N_15446);
and U23961 (N_23961,N_18322,N_15424);
nor U23962 (N_23962,N_16292,N_18343);
xnor U23963 (N_23963,N_17440,N_19093);
and U23964 (N_23964,N_15024,N_15543);
nand U23965 (N_23965,N_18011,N_15938);
nand U23966 (N_23966,N_19053,N_15310);
nor U23967 (N_23967,N_16944,N_18211);
and U23968 (N_23968,N_16200,N_15287);
nor U23969 (N_23969,N_19717,N_15289);
nand U23970 (N_23970,N_17596,N_17044);
nand U23971 (N_23971,N_17734,N_19366);
nand U23972 (N_23972,N_15358,N_16636);
or U23973 (N_23973,N_17725,N_16437);
xnor U23974 (N_23974,N_18723,N_17445);
or U23975 (N_23975,N_19801,N_17954);
xnor U23976 (N_23976,N_19099,N_17652);
nand U23977 (N_23977,N_16515,N_19089);
or U23978 (N_23978,N_17780,N_18298);
xnor U23979 (N_23979,N_19439,N_19320);
nand U23980 (N_23980,N_15974,N_15246);
and U23981 (N_23981,N_19146,N_15733);
and U23982 (N_23982,N_17273,N_16030);
or U23983 (N_23983,N_16551,N_15573);
xor U23984 (N_23984,N_17203,N_15415);
and U23985 (N_23985,N_16306,N_19253);
xor U23986 (N_23986,N_17388,N_15720);
nor U23987 (N_23987,N_16903,N_15775);
or U23988 (N_23988,N_15043,N_19336);
nand U23989 (N_23989,N_15149,N_16763);
and U23990 (N_23990,N_19804,N_17325);
nand U23991 (N_23991,N_15376,N_19742);
nor U23992 (N_23992,N_18735,N_15560);
nand U23993 (N_23993,N_17814,N_15695);
or U23994 (N_23994,N_16513,N_17574);
xnor U23995 (N_23995,N_19341,N_15659);
nand U23996 (N_23996,N_17159,N_19909);
nor U23997 (N_23997,N_17260,N_15905);
nand U23998 (N_23998,N_18082,N_15529);
or U23999 (N_23999,N_16333,N_16903);
xor U24000 (N_24000,N_16182,N_19047);
xor U24001 (N_24001,N_16310,N_15032);
xor U24002 (N_24002,N_17586,N_19000);
xnor U24003 (N_24003,N_17468,N_16381);
xnor U24004 (N_24004,N_17685,N_17986);
and U24005 (N_24005,N_19887,N_19539);
xnor U24006 (N_24006,N_17967,N_19074);
or U24007 (N_24007,N_15448,N_16151);
and U24008 (N_24008,N_18853,N_19964);
xor U24009 (N_24009,N_19643,N_19327);
xnor U24010 (N_24010,N_15674,N_17434);
xnor U24011 (N_24011,N_16284,N_17196);
and U24012 (N_24012,N_19524,N_17638);
or U24013 (N_24013,N_16340,N_16087);
or U24014 (N_24014,N_16941,N_16954);
or U24015 (N_24015,N_15761,N_17387);
xor U24016 (N_24016,N_18052,N_18292);
or U24017 (N_24017,N_17306,N_15554);
or U24018 (N_24018,N_18449,N_16900);
and U24019 (N_24019,N_17418,N_16459);
nor U24020 (N_24020,N_19406,N_17027);
nor U24021 (N_24021,N_17356,N_16512);
nor U24022 (N_24022,N_18051,N_15230);
and U24023 (N_24023,N_15029,N_16518);
or U24024 (N_24024,N_17830,N_16431);
or U24025 (N_24025,N_17805,N_19578);
or U24026 (N_24026,N_18312,N_18698);
and U24027 (N_24027,N_18748,N_17374);
nand U24028 (N_24028,N_19443,N_16800);
nand U24029 (N_24029,N_15508,N_19588);
xnor U24030 (N_24030,N_18364,N_16321);
nor U24031 (N_24031,N_18555,N_19047);
nand U24032 (N_24032,N_19891,N_19320);
nor U24033 (N_24033,N_17969,N_18010);
nor U24034 (N_24034,N_18754,N_17752);
or U24035 (N_24035,N_19263,N_16513);
nand U24036 (N_24036,N_18648,N_16551);
nand U24037 (N_24037,N_15310,N_19376);
xnor U24038 (N_24038,N_18650,N_18800);
nor U24039 (N_24039,N_18476,N_17064);
and U24040 (N_24040,N_17768,N_17746);
nor U24041 (N_24041,N_17952,N_15300);
xnor U24042 (N_24042,N_19536,N_15067);
or U24043 (N_24043,N_17025,N_15552);
nor U24044 (N_24044,N_15590,N_15510);
or U24045 (N_24045,N_16470,N_16465);
nand U24046 (N_24046,N_15674,N_17755);
nor U24047 (N_24047,N_16435,N_15947);
or U24048 (N_24048,N_18135,N_18370);
or U24049 (N_24049,N_15249,N_18240);
or U24050 (N_24050,N_18151,N_19074);
nand U24051 (N_24051,N_16824,N_15245);
and U24052 (N_24052,N_16336,N_18717);
and U24053 (N_24053,N_17343,N_18981);
and U24054 (N_24054,N_17751,N_19905);
or U24055 (N_24055,N_15207,N_15310);
nand U24056 (N_24056,N_17525,N_16158);
and U24057 (N_24057,N_19238,N_15793);
nor U24058 (N_24058,N_18542,N_18252);
xnor U24059 (N_24059,N_16494,N_19607);
xor U24060 (N_24060,N_18917,N_15329);
or U24061 (N_24061,N_16743,N_15018);
or U24062 (N_24062,N_15989,N_15100);
nor U24063 (N_24063,N_17925,N_19308);
xor U24064 (N_24064,N_18351,N_16889);
or U24065 (N_24065,N_15638,N_17569);
nand U24066 (N_24066,N_18854,N_15638);
nor U24067 (N_24067,N_19350,N_16338);
and U24068 (N_24068,N_16781,N_19529);
nor U24069 (N_24069,N_18906,N_16296);
xnor U24070 (N_24070,N_18235,N_19597);
xor U24071 (N_24071,N_16367,N_19187);
or U24072 (N_24072,N_15078,N_18502);
nor U24073 (N_24073,N_18785,N_16249);
nor U24074 (N_24074,N_16600,N_15162);
xor U24075 (N_24075,N_15674,N_17003);
and U24076 (N_24076,N_18294,N_16907);
or U24077 (N_24077,N_15556,N_15251);
xnor U24078 (N_24078,N_18162,N_17006);
and U24079 (N_24079,N_16894,N_19321);
nor U24080 (N_24080,N_18946,N_15502);
nor U24081 (N_24081,N_16862,N_19056);
or U24082 (N_24082,N_19678,N_15333);
nor U24083 (N_24083,N_18095,N_16585);
and U24084 (N_24084,N_15016,N_18626);
or U24085 (N_24085,N_16210,N_16574);
nand U24086 (N_24086,N_17398,N_17212);
xor U24087 (N_24087,N_19629,N_18561);
and U24088 (N_24088,N_19197,N_15476);
xnor U24089 (N_24089,N_18735,N_16465);
xor U24090 (N_24090,N_15884,N_16925);
nand U24091 (N_24091,N_15602,N_16254);
and U24092 (N_24092,N_18896,N_16722);
xnor U24093 (N_24093,N_15728,N_16492);
nor U24094 (N_24094,N_18059,N_15286);
nor U24095 (N_24095,N_16075,N_19408);
and U24096 (N_24096,N_15491,N_15844);
nor U24097 (N_24097,N_17236,N_15243);
nor U24098 (N_24098,N_19311,N_15965);
nand U24099 (N_24099,N_16111,N_18967);
xnor U24100 (N_24100,N_16087,N_15302);
and U24101 (N_24101,N_16152,N_17544);
and U24102 (N_24102,N_19853,N_18525);
nor U24103 (N_24103,N_15215,N_15911);
and U24104 (N_24104,N_17813,N_19929);
nand U24105 (N_24105,N_16210,N_18986);
or U24106 (N_24106,N_16864,N_15051);
and U24107 (N_24107,N_16148,N_18626);
or U24108 (N_24108,N_18379,N_15871);
xnor U24109 (N_24109,N_19568,N_15857);
or U24110 (N_24110,N_16083,N_18316);
nand U24111 (N_24111,N_19297,N_19894);
nor U24112 (N_24112,N_18582,N_19006);
or U24113 (N_24113,N_15383,N_15460);
nand U24114 (N_24114,N_18584,N_19189);
nor U24115 (N_24115,N_18281,N_16531);
nand U24116 (N_24116,N_15084,N_16113);
or U24117 (N_24117,N_19591,N_17740);
xnor U24118 (N_24118,N_16443,N_19031);
and U24119 (N_24119,N_17278,N_17533);
xnor U24120 (N_24120,N_15153,N_18682);
nand U24121 (N_24121,N_17885,N_15304);
and U24122 (N_24122,N_17204,N_15770);
xnor U24123 (N_24123,N_17850,N_18010);
and U24124 (N_24124,N_17271,N_16406);
xor U24125 (N_24125,N_18870,N_19152);
nand U24126 (N_24126,N_17584,N_16035);
and U24127 (N_24127,N_15046,N_18482);
nand U24128 (N_24128,N_18824,N_16025);
or U24129 (N_24129,N_18378,N_15715);
and U24130 (N_24130,N_16317,N_19335);
xor U24131 (N_24131,N_19822,N_15126);
nor U24132 (N_24132,N_17933,N_18891);
nand U24133 (N_24133,N_19257,N_19700);
and U24134 (N_24134,N_17952,N_19002);
xnor U24135 (N_24135,N_16835,N_17428);
and U24136 (N_24136,N_18514,N_19803);
nor U24137 (N_24137,N_17684,N_17203);
xor U24138 (N_24138,N_17822,N_19660);
and U24139 (N_24139,N_18703,N_18693);
nand U24140 (N_24140,N_18560,N_17243);
xor U24141 (N_24141,N_16016,N_16547);
nor U24142 (N_24142,N_19306,N_17096);
and U24143 (N_24143,N_15295,N_15930);
or U24144 (N_24144,N_17500,N_19943);
and U24145 (N_24145,N_19072,N_17051);
xor U24146 (N_24146,N_19085,N_19185);
xor U24147 (N_24147,N_18563,N_19850);
nor U24148 (N_24148,N_18225,N_15482);
or U24149 (N_24149,N_15256,N_19887);
xnor U24150 (N_24150,N_15039,N_18199);
or U24151 (N_24151,N_18560,N_16617);
nor U24152 (N_24152,N_19992,N_18476);
xor U24153 (N_24153,N_19672,N_18007);
nand U24154 (N_24154,N_19986,N_19117);
xnor U24155 (N_24155,N_17553,N_19017);
nand U24156 (N_24156,N_15051,N_18673);
xor U24157 (N_24157,N_16006,N_17451);
and U24158 (N_24158,N_19688,N_15280);
nor U24159 (N_24159,N_16975,N_18504);
nor U24160 (N_24160,N_19396,N_15127);
or U24161 (N_24161,N_16965,N_18867);
or U24162 (N_24162,N_17235,N_16136);
nor U24163 (N_24163,N_15929,N_16565);
xor U24164 (N_24164,N_15789,N_16287);
nor U24165 (N_24165,N_16647,N_17471);
or U24166 (N_24166,N_16199,N_19100);
and U24167 (N_24167,N_19115,N_19023);
xnor U24168 (N_24168,N_17884,N_15377);
and U24169 (N_24169,N_19122,N_19385);
or U24170 (N_24170,N_16683,N_16224);
xnor U24171 (N_24171,N_16840,N_16879);
and U24172 (N_24172,N_16052,N_17659);
or U24173 (N_24173,N_17433,N_16057);
xnor U24174 (N_24174,N_18276,N_17566);
or U24175 (N_24175,N_16899,N_19945);
xor U24176 (N_24176,N_18534,N_16252);
nor U24177 (N_24177,N_15199,N_19655);
or U24178 (N_24178,N_17312,N_17748);
xnor U24179 (N_24179,N_19226,N_16484);
xnor U24180 (N_24180,N_18292,N_17889);
or U24181 (N_24181,N_15324,N_18346);
or U24182 (N_24182,N_18369,N_16096);
and U24183 (N_24183,N_17777,N_17404);
and U24184 (N_24184,N_17571,N_15589);
or U24185 (N_24185,N_17744,N_18408);
nor U24186 (N_24186,N_17537,N_15754);
nor U24187 (N_24187,N_19316,N_17581);
and U24188 (N_24188,N_17471,N_15616);
nor U24189 (N_24189,N_15795,N_17126);
or U24190 (N_24190,N_16217,N_18328);
or U24191 (N_24191,N_18381,N_19704);
nand U24192 (N_24192,N_17144,N_15954);
and U24193 (N_24193,N_18165,N_17376);
or U24194 (N_24194,N_16943,N_16869);
nand U24195 (N_24195,N_15029,N_18437);
xor U24196 (N_24196,N_16559,N_18196);
or U24197 (N_24197,N_19315,N_18132);
nor U24198 (N_24198,N_16094,N_19082);
and U24199 (N_24199,N_15431,N_16836);
nand U24200 (N_24200,N_16356,N_19292);
and U24201 (N_24201,N_16563,N_16320);
xnor U24202 (N_24202,N_15411,N_15673);
and U24203 (N_24203,N_18378,N_15380);
or U24204 (N_24204,N_15474,N_19127);
and U24205 (N_24205,N_18492,N_17281);
and U24206 (N_24206,N_18381,N_18523);
or U24207 (N_24207,N_19190,N_15809);
nor U24208 (N_24208,N_15058,N_15908);
nand U24209 (N_24209,N_16072,N_19582);
or U24210 (N_24210,N_17039,N_18779);
nor U24211 (N_24211,N_18934,N_17185);
xnor U24212 (N_24212,N_19021,N_18316);
and U24213 (N_24213,N_15344,N_17346);
nand U24214 (N_24214,N_19905,N_18990);
nand U24215 (N_24215,N_17739,N_17537);
nand U24216 (N_24216,N_16982,N_15293);
nand U24217 (N_24217,N_16711,N_19600);
or U24218 (N_24218,N_18540,N_18151);
nand U24219 (N_24219,N_17143,N_16267);
and U24220 (N_24220,N_15525,N_17036);
or U24221 (N_24221,N_15206,N_15323);
nand U24222 (N_24222,N_18412,N_19522);
nor U24223 (N_24223,N_17241,N_18712);
nor U24224 (N_24224,N_17351,N_19364);
xor U24225 (N_24225,N_19072,N_17640);
nor U24226 (N_24226,N_15698,N_17310);
nand U24227 (N_24227,N_17098,N_16063);
or U24228 (N_24228,N_16106,N_18724);
nor U24229 (N_24229,N_16690,N_17145);
nand U24230 (N_24230,N_18296,N_18532);
and U24231 (N_24231,N_18027,N_15558);
xor U24232 (N_24232,N_17540,N_19567);
and U24233 (N_24233,N_16434,N_16920);
or U24234 (N_24234,N_15757,N_15559);
or U24235 (N_24235,N_16874,N_17411);
and U24236 (N_24236,N_17617,N_17681);
and U24237 (N_24237,N_15480,N_16636);
and U24238 (N_24238,N_18286,N_18870);
nand U24239 (N_24239,N_17159,N_18397);
nor U24240 (N_24240,N_18722,N_16236);
or U24241 (N_24241,N_18882,N_17813);
nor U24242 (N_24242,N_19841,N_17587);
xor U24243 (N_24243,N_17755,N_16668);
nor U24244 (N_24244,N_17780,N_17936);
or U24245 (N_24245,N_15380,N_16836);
xnor U24246 (N_24246,N_17909,N_18540);
nor U24247 (N_24247,N_15054,N_18367);
or U24248 (N_24248,N_18386,N_17824);
or U24249 (N_24249,N_16522,N_19730);
or U24250 (N_24250,N_16211,N_17378);
nor U24251 (N_24251,N_18081,N_18238);
or U24252 (N_24252,N_17759,N_17668);
or U24253 (N_24253,N_15235,N_18607);
nor U24254 (N_24254,N_17549,N_18028);
xor U24255 (N_24255,N_15279,N_19732);
xor U24256 (N_24256,N_18717,N_15962);
or U24257 (N_24257,N_19732,N_16344);
nand U24258 (N_24258,N_18601,N_18198);
nor U24259 (N_24259,N_16216,N_19508);
nor U24260 (N_24260,N_15195,N_19028);
nand U24261 (N_24261,N_19510,N_17230);
or U24262 (N_24262,N_15362,N_19001);
or U24263 (N_24263,N_19342,N_16553);
xor U24264 (N_24264,N_19835,N_15929);
xnor U24265 (N_24265,N_17377,N_19831);
xnor U24266 (N_24266,N_19838,N_17274);
nand U24267 (N_24267,N_19353,N_18067);
xor U24268 (N_24268,N_17550,N_16838);
or U24269 (N_24269,N_19195,N_18336);
or U24270 (N_24270,N_15958,N_18875);
nand U24271 (N_24271,N_17020,N_15366);
nand U24272 (N_24272,N_15876,N_18849);
nand U24273 (N_24273,N_19401,N_16713);
and U24274 (N_24274,N_15659,N_18542);
nor U24275 (N_24275,N_15885,N_18733);
nor U24276 (N_24276,N_19574,N_19669);
xor U24277 (N_24277,N_18729,N_15988);
nand U24278 (N_24278,N_15934,N_18249);
nor U24279 (N_24279,N_18921,N_19963);
xnor U24280 (N_24280,N_19341,N_19616);
xor U24281 (N_24281,N_15021,N_16467);
and U24282 (N_24282,N_18017,N_16235);
nand U24283 (N_24283,N_16021,N_18091);
nand U24284 (N_24284,N_16052,N_16874);
and U24285 (N_24285,N_16379,N_15179);
nand U24286 (N_24286,N_15335,N_16841);
nand U24287 (N_24287,N_19625,N_16239);
xor U24288 (N_24288,N_18079,N_16032);
nand U24289 (N_24289,N_17026,N_15048);
or U24290 (N_24290,N_16020,N_19986);
and U24291 (N_24291,N_18436,N_17734);
or U24292 (N_24292,N_19300,N_16484);
nor U24293 (N_24293,N_15483,N_18594);
and U24294 (N_24294,N_16832,N_16664);
nor U24295 (N_24295,N_18552,N_15534);
or U24296 (N_24296,N_17390,N_18503);
or U24297 (N_24297,N_15081,N_18413);
and U24298 (N_24298,N_18495,N_15362);
nor U24299 (N_24299,N_17918,N_18142);
nor U24300 (N_24300,N_15233,N_16145);
nor U24301 (N_24301,N_16554,N_18046);
and U24302 (N_24302,N_16785,N_15873);
xor U24303 (N_24303,N_17620,N_18123);
nor U24304 (N_24304,N_17385,N_16697);
or U24305 (N_24305,N_18757,N_19024);
nor U24306 (N_24306,N_17387,N_19407);
and U24307 (N_24307,N_16933,N_15091);
or U24308 (N_24308,N_16666,N_16853);
and U24309 (N_24309,N_15995,N_17458);
or U24310 (N_24310,N_17605,N_16681);
nor U24311 (N_24311,N_19806,N_15762);
nor U24312 (N_24312,N_18452,N_16063);
nor U24313 (N_24313,N_16192,N_19321);
nand U24314 (N_24314,N_16841,N_19747);
and U24315 (N_24315,N_17036,N_18772);
nor U24316 (N_24316,N_15991,N_17882);
nor U24317 (N_24317,N_15105,N_17051);
or U24318 (N_24318,N_15932,N_19580);
or U24319 (N_24319,N_15952,N_16049);
nor U24320 (N_24320,N_19932,N_19773);
or U24321 (N_24321,N_15488,N_17373);
or U24322 (N_24322,N_16354,N_18395);
nand U24323 (N_24323,N_17964,N_18615);
and U24324 (N_24324,N_16932,N_19232);
and U24325 (N_24325,N_18626,N_16670);
xnor U24326 (N_24326,N_16530,N_19459);
and U24327 (N_24327,N_18881,N_18197);
nor U24328 (N_24328,N_19676,N_16257);
or U24329 (N_24329,N_18858,N_19477);
or U24330 (N_24330,N_17888,N_19210);
and U24331 (N_24331,N_17654,N_16412);
or U24332 (N_24332,N_17375,N_18781);
nand U24333 (N_24333,N_15024,N_15176);
nor U24334 (N_24334,N_17001,N_19643);
or U24335 (N_24335,N_15796,N_15743);
nor U24336 (N_24336,N_18227,N_18021);
xnor U24337 (N_24337,N_18885,N_15968);
or U24338 (N_24338,N_17013,N_16937);
and U24339 (N_24339,N_17860,N_19684);
xnor U24340 (N_24340,N_16375,N_19414);
nor U24341 (N_24341,N_17903,N_19795);
xor U24342 (N_24342,N_16515,N_15731);
nor U24343 (N_24343,N_18707,N_18988);
xor U24344 (N_24344,N_19870,N_17219);
nand U24345 (N_24345,N_18381,N_15806);
nand U24346 (N_24346,N_17059,N_18147);
and U24347 (N_24347,N_17041,N_17107);
and U24348 (N_24348,N_15244,N_19237);
or U24349 (N_24349,N_19627,N_19573);
xor U24350 (N_24350,N_19904,N_19622);
nand U24351 (N_24351,N_18158,N_16207);
nand U24352 (N_24352,N_15003,N_17279);
nor U24353 (N_24353,N_17590,N_19130);
and U24354 (N_24354,N_16370,N_18478);
nor U24355 (N_24355,N_16575,N_15211);
nor U24356 (N_24356,N_18630,N_19760);
xor U24357 (N_24357,N_18510,N_16793);
xnor U24358 (N_24358,N_19196,N_18222);
nand U24359 (N_24359,N_15708,N_15703);
nor U24360 (N_24360,N_18790,N_19040);
or U24361 (N_24361,N_16882,N_18567);
or U24362 (N_24362,N_17560,N_19669);
or U24363 (N_24363,N_17787,N_19849);
and U24364 (N_24364,N_16701,N_19918);
xnor U24365 (N_24365,N_19613,N_16402);
nor U24366 (N_24366,N_15226,N_18960);
nor U24367 (N_24367,N_16070,N_16146);
nand U24368 (N_24368,N_19049,N_19112);
nand U24369 (N_24369,N_17551,N_19641);
nand U24370 (N_24370,N_17978,N_17718);
and U24371 (N_24371,N_19792,N_19438);
nor U24372 (N_24372,N_15261,N_16170);
xnor U24373 (N_24373,N_19009,N_19855);
or U24374 (N_24374,N_19694,N_17297);
nor U24375 (N_24375,N_16295,N_17548);
and U24376 (N_24376,N_16395,N_18367);
nor U24377 (N_24377,N_15488,N_15678);
or U24378 (N_24378,N_19058,N_18007);
and U24379 (N_24379,N_17094,N_17476);
nor U24380 (N_24380,N_16244,N_17307);
and U24381 (N_24381,N_16413,N_17593);
nor U24382 (N_24382,N_16415,N_19309);
and U24383 (N_24383,N_16169,N_16240);
nor U24384 (N_24384,N_15568,N_17744);
and U24385 (N_24385,N_17869,N_19478);
nor U24386 (N_24386,N_17818,N_16115);
nand U24387 (N_24387,N_19783,N_18737);
nand U24388 (N_24388,N_19386,N_17219);
nand U24389 (N_24389,N_19556,N_16097);
nor U24390 (N_24390,N_16553,N_18864);
nor U24391 (N_24391,N_19825,N_17003);
nand U24392 (N_24392,N_18932,N_15338);
xnor U24393 (N_24393,N_16239,N_17310);
nand U24394 (N_24394,N_17450,N_15879);
or U24395 (N_24395,N_19642,N_18348);
or U24396 (N_24396,N_18891,N_15057);
nand U24397 (N_24397,N_18369,N_16770);
nor U24398 (N_24398,N_18809,N_17187);
nor U24399 (N_24399,N_17868,N_15440);
xor U24400 (N_24400,N_15131,N_16137);
nand U24401 (N_24401,N_19342,N_16370);
or U24402 (N_24402,N_17938,N_16861);
nand U24403 (N_24403,N_17056,N_16910);
nor U24404 (N_24404,N_15215,N_17594);
or U24405 (N_24405,N_15579,N_17126);
xor U24406 (N_24406,N_16268,N_17714);
nor U24407 (N_24407,N_19623,N_18933);
nand U24408 (N_24408,N_19805,N_15732);
nand U24409 (N_24409,N_15807,N_15668);
nor U24410 (N_24410,N_18056,N_19843);
and U24411 (N_24411,N_15636,N_19325);
and U24412 (N_24412,N_18693,N_15510);
nor U24413 (N_24413,N_18602,N_19191);
nor U24414 (N_24414,N_18951,N_19100);
or U24415 (N_24415,N_16674,N_19072);
and U24416 (N_24416,N_18433,N_16007);
or U24417 (N_24417,N_18128,N_17291);
xor U24418 (N_24418,N_16067,N_19938);
or U24419 (N_24419,N_16440,N_17018);
and U24420 (N_24420,N_18613,N_19586);
nand U24421 (N_24421,N_17040,N_17180);
xnor U24422 (N_24422,N_19867,N_16443);
or U24423 (N_24423,N_19706,N_19384);
and U24424 (N_24424,N_19721,N_17318);
nand U24425 (N_24425,N_19652,N_15058);
nor U24426 (N_24426,N_16792,N_15332);
and U24427 (N_24427,N_15978,N_17745);
nor U24428 (N_24428,N_18974,N_19684);
nor U24429 (N_24429,N_19335,N_15224);
nand U24430 (N_24430,N_16727,N_17196);
nand U24431 (N_24431,N_18875,N_19648);
or U24432 (N_24432,N_15178,N_18298);
or U24433 (N_24433,N_16258,N_18950);
and U24434 (N_24434,N_15579,N_18614);
nor U24435 (N_24435,N_19968,N_17845);
nand U24436 (N_24436,N_18288,N_16358);
nor U24437 (N_24437,N_17114,N_17875);
and U24438 (N_24438,N_18386,N_16255);
and U24439 (N_24439,N_18183,N_19574);
nand U24440 (N_24440,N_16415,N_16493);
nor U24441 (N_24441,N_19216,N_19560);
nand U24442 (N_24442,N_18378,N_15052);
xor U24443 (N_24443,N_15964,N_17179);
nand U24444 (N_24444,N_18824,N_15034);
nor U24445 (N_24445,N_18144,N_15762);
xor U24446 (N_24446,N_15162,N_16961);
nand U24447 (N_24447,N_19232,N_15907);
nor U24448 (N_24448,N_15759,N_16706);
or U24449 (N_24449,N_19331,N_15144);
nor U24450 (N_24450,N_15590,N_17856);
or U24451 (N_24451,N_17096,N_19378);
xor U24452 (N_24452,N_19402,N_18060);
xor U24453 (N_24453,N_19237,N_18387);
xor U24454 (N_24454,N_19590,N_19560);
and U24455 (N_24455,N_16015,N_17752);
nor U24456 (N_24456,N_19275,N_17401);
and U24457 (N_24457,N_16657,N_19565);
nor U24458 (N_24458,N_16182,N_16550);
or U24459 (N_24459,N_17387,N_17700);
or U24460 (N_24460,N_19790,N_18999);
or U24461 (N_24461,N_19461,N_15465);
xnor U24462 (N_24462,N_16093,N_15275);
xnor U24463 (N_24463,N_19520,N_16993);
nor U24464 (N_24464,N_15015,N_16689);
xnor U24465 (N_24465,N_18722,N_16334);
xor U24466 (N_24466,N_18569,N_16291);
xnor U24467 (N_24467,N_16662,N_19968);
or U24468 (N_24468,N_15947,N_15743);
nor U24469 (N_24469,N_17863,N_18274);
or U24470 (N_24470,N_16227,N_17145);
or U24471 (N_24471,N_15232,N_15093);
nor U24472 (N_24472,N_15488,N_16945);
nand U24473 (N_24473,N_17930,N_15450);
nand U24474 (N_24474,N_17847,N_17449);
nor U24475 (N_24475,N_18867,N_15015);
nand U24476 (N_24476,N_19891,N_19642);
nor U24477 (N_24477,N_18947,N_15949);
xor U24478 (N_24478,N_19126,N_16180);
and U24479 (N_24479,N_18738,N_17559);
nand U24480 (N_24480,N_18936,N_15401);
nand U24481 (N_24481,N_18931,N_17716);
and U24482 (N_24482,N_16157,N_16474);
xor U24483 (N_24483,N_18515,N_15743);
and U24484 (N_24484,N_18737,N_17284);
xor U24485 (N_24485,N_19869,N_18447);
xnor U24486 (N_24486,N_19363,N_17446);
xor U24487 (N_24487,N_19356,N_19606);
and U24488 (N_24488,N_17096,N_15579);
nor U24489 (N_24489,N_17411,N_17511);
and U24490 (N_24490,N_17248,N_17456);
or U24491 (N_24491,N_18643,N_15607);
or U24492 (N_24492,N_15351,N_17930);
nand U24493 (N_24493,N_17176,N_16589);
and U24494 (N_24494,N_19695,N_19971);
or U24495 (N_24495,N_19572,N_17937);
and U24496 (N_24496,N_19410,N_17989);
and U24497 (N_24497,N_15890,N_18109);
xnor U24498 (N_24498,N_15120,N_15329);
nor U24499 (N_24499,N_15356,N_19923);
and U24500 (N_24500,N_17123,N_19302);
and U24501 (N_24501,N_15412,N_16074);
nor U24502 (N_24502,N_15771,N_17300);
xor U24503 (N_24503,N_19839,N_16595);
and U24504 (N_24504,N_19292,N_15243);
nand U24505 (N_24505,N_16790,N_18720);
and U24506 (N_24506,N_16154,N_19067);
nand U24507 (N_24507,N_19723,N_19035);
and U24508 (N_24508,N_17145,N_19134);
nor U24509 (N_24509,N_15247,N_16211);
nand U24510 (N_24510,N_17301,N_17417);
nand U24511 (N_24511,N_15776,N_19398);
and U24512 (N_24512,N_16109,N_19215);
xor U24513 (N_24513,N_16091,N_18442);
and U24514 (N_24514,N_15425,N_15946);
nand U24515 (N_24515,N_15300,N_18711);
nor U24516 (N_24516,N_15300,N_17365);
xnor U24517 (N_24517,N_18878,N_19760);
and U24518 (N_24518,N_19780,N_17313);
nor U24519 (N_24519,N_15663,N_19358);
nor U24520 (N_24520,N_19804,N_15468);
nand U24521 (N_24521,N_16343,N_15741);
and U24522 (N_24522,N_15939,N_19650);
nor U24523 (N_24523,N_18933,N_15629);
or U24524 (N_24524,N_18908,N_15167);
nor U24525 (N_24525,N_18593,N_18213);
xor U24526 (N_24526,N_17701,N_19280);
nand U24527 (N_24527,N_16907,N_19912);
xnor U24528 (N_24528,N_17290,N_16720);
nor U24529 (N_24529,N_16902,N_16905);
xnor U24530 (N_24530,N_15249,N_16634);
or U24531 (N_24531,N_15622,N_15025);
xor U24532 (N_24532,N_18379,N_19325);
xor U24533 (N_24533,N_18568,N_15486);
nor U24534 (N_24534,N_15857,N_19080);
xor U24535 (N_24535,N_19430,N_19157);
or U24536 (N_24536,N_16627,N_17873);
nand U24537 (N_24537,N_16832,N_17495);
or U24538 (N_24538,N_16067,N_15902);
nor U24539 (N_24539,N_15542,N_17793);
and U24540 (N_24540,N_17518,N_15205);
nand U24541 (N_24541,N_18590,N_19195);
and U24542 (N_24542,N_19940,N_19270);
nor U24543 (N_24543,N_19485,N_19213);
nand U24544 (N_24544,N_18590,N_17129);
or U24545 (N_24545,N_18491,N_18972);
xor U24546 (N_24546,N_19046,N_16983);
xnor U24547 (N_24547,N_17108,N_19105);
and U24548 (N_24548,N_18740,N_19600);
nor U24549 (N_24549,N_16483,N_17703);
and U24550 (N_24550,N_18853,N_15745);
nand U24551 (N_24551,N_15097,N_18658);
or U24552 (N_24552,N_18755,N_18229);
or U24553 (N_24553,N_16739,N_18683);
nor U24554 (N_24554,N_19789,N_18907);
or U24555 (N_24555,N_19354,N_17172);
xnor U24556 (N_24556,N_18661,N_16184);
xor U24557 (N_24557,N_15007,N_19418);
and U24558 (N_24558,N_19367,N_16523);
nand U24559 (N_24559,N_17007,N_17384);
xor U24560 (N_24560,N_17948,N_19739);
and U24561 (N_24561,N_16633,N_16177);
and U24562 (N_24562,N_16593,N_15095);
nor U24563 (N_24563,N_17544,N_15096);
and U24564 (N_24564,N_16280,N_19955);
or U24565 (N_24565,N_17694,N_17691);
xnor U24566 (N_24566,N_15210,N_16919);
or U24567 (N_24567,N_16054,N_17138);
nor U24568 (N_24568,N_18058,N_17247);
and U24569 (N_24569,N_15688,N_17164);
and U24570 (N_24570,N_19316,N_17613);
nand U24571 (N_24571,N_18015,N_16831);
or U24572 (N_24572,N_18918,N_17529);
nor U24573 (N_24573,N_16283,N_19731);
xor U24574 (N_24574,N_15303,N_17800);
nor U24575 (N_24575,N_16695,N_16120);
nor U24576 (N_24576,N_18379,N_16240);
nand U24577 (N_24577,N_16861,N_18452);
xor U24578 (N_24578,N_19040,N_18594);
nor U24579 (N_24579,N_15080,N_15396);
nor U24580 (N_24580,N_15657,N_16861);
nor U24581 (N_24581,N_17914,N_18223);
or U24582 (N_24582,N_18169,N_15448);
or U24583 (N_24583,N_16923,N_16562);
xnor U24584 (N_24584,N_15609,N_19281);
nor U24585 (N_24585,N_19588,N_17410);
nand U24586 (N_24586,N_18757,N_18950);
xnor U24587 (N_24587,N_16512,N_18950);
or U24588 (N_24588,N_16509,N_15345);
xor U24589 (N_24589,N_16296,N_16289);
xor U24590 (N_24590,N_16304,N_18690);
or U24591 (N_24591,N_19971,N_19183);
nor U24592 (N_24592,N_18526,N_19437);
nor U24593 (N_24593,N_15945,N_15207);
and U24594 (N_24594,N_18694,N_16219);
xnor U24595 (N_24595,N_16837,N_19827);
nand U24596 (N_24596,N_17081,N_18686);
nor U24597 (N_24597,N_18928,N_19221);
nand U24598 (N_24598,N_15549,N_15033);
xnor U24599 (N_24599,N_19954,N_17622);
nand U24600 (N_24600,N_16561,N_16339);
and U24601 (N_24601,N_17482,N_17589);
xnor U24602 (N_24602,N_18529,N_15266);
nor U24603 (N_24603,N_18861,N_16248);
and U24604 (N_24604,N_18664,N_16457);
or U24605 (N_24605,N_15068,N_16354);
nand U24606 (N_24606,N_18491,N_18442);
and U24607 (N_24607,N_19087,N_19539);
xnor U24608 (N_24608,N_17892,N_16905);
xor U24609 (N_24609,N_19913,N_19979);
xor U24610 (N_24610,N_15375,N_18860);
xnor U24611 (N_24611,N_17912,N_18080);
xnor U24612 (N_24612,N_17667,N_16365);
and U24613 (N_24613,N_19267,N_17185);
and U24614 (N_24614,N_15294,N_18589);
nand U24615 (N_24615,N_15984,N_17203);
nor U24616 (N_24616,N_16156,N_15093);
and U24617 (N_24617,N_16063,N_16709);
nor U24618 (N_24618,N_16418,N_16266);
xor U24619 (N_24619,N_17292,N_17142);
nand U24620 (N_24620,N_15030,N_19238);
xor U24621 (N_24621,N_16106,N_19997);
nor U24622 (N_24622,N_19316,N_19295);
or U24623 (N_24623,N_19357,N_16750);
xnor U24624 (N_24624,N_16133,N_17111);
or U24625 (N_24625,N_18884,N_18952);
or U24626 (N_24626,N_15772,N_19784);
nand U24627 (N_24627,N_16283,N_18524);
xor U24628 (N_24628,N_18913,N_16189);
or U24629 (N_24629,N_15870,N_16418);
nor U24630 (N_24630,N_18840,N_15717);
and U24631 (N_24631,N_19170,N_19605);
nor U24632 (N_24632,N_19990,N_17802);
xnor U24633 (N_24633,N_17745,N_16020);
xor U24634 (N_24634,N_16232,N_18942);
and U24635 (N_24635,N_19116,N_17346);
xor U24636 (N_24636,N_18828,N_15621);
and U24637 (N_24637,N_19618,N_15222);
nand U24638 (N_24638,N_17537,N_16466);
or U24639 (N_24639,N_15172,N_15857);
xnor U24640 (N_24640,N_18014,N_17782);
nor U24641 (N_24641,N_18182,N_16311);
nor U24642 (N_24642,N_18707,N_17335);
or U24643 (N_24643,N_15563,N_18492);
xor U24644 (N_24644,N_17561,N_16005);
xor U24645 (N_24645,N_15835,N_18997);
nor U24646 (N_24646,N_15966,N_15587);
or U24647 (N_24647,N_17880,N_15569);
and U24648 (N_24648,N_19034,N_15451);
nand U24649 (N_24649,N_15478,N_18885);
or U24650 (N_24650,N_15886,N_19387);
nor U24651 (N_24651,N_19979,N_19439);
nor U24652 (N_24652,N_18161,N_15843);
xor U24653 (N_24653,N_18002,N_15772);
and U24654 (N_24654,N_15053,N_19434);
or U24655 (N_24655,N_19633,N_16402);
or U24656 (N_24656,N_15230,N_17056);
nor U24657 (N_24657,N_15727,N_16111);
nor U24658 (N_24658,N_16097,N_15742);
nand U24659 (N_24659,N_19769,N_16663);
nor U24660 (N_24660,N_18482,N_19856);
or U24661 (N_24661,N_19800,N_15444);
nor U24662 (N_24662,N_19431,N_15122);
and U24663 (N_24663,N_15795,N_15659);
nor U24664 (N_24664,N_17844,N_15176);
xnor U24665 (N_24665,N_15017,N_17194);
nand U24666 (N_24666,N_19412,N_15903);
nor U24667 (N_24667,N_19003,N_18966);
nor U24668 (N_24668,N_16793,N_15473);
xnor U24669 (N_24669,N_19042,N_19300);
or U24670 (N_24670,N_19255,N_17939);
or U24671 (N_24671,N_17835,N_16854);
and U24672 (N_24672,N_16777,N_15140);
nor U24673 (N_24673,N_19958,N_18869);
nor U24674 (N_24674,N_18585,N_19726);
and U24675 (N_24675,N_16269,N_17251);
and U24676 (N_24676,N_15513,N_16602);
and U24677 (N_24677,N_17089,N_18614);
nor U24678 (N_24678,N_18059,N_18324);
xnor U24679 (N_24679,N_19650,N_16996);
xnor U24680 (N_24680,N_17294,N_16949);
or U24681 (N_24681,N_18690,N_15881);
xnor U24682 (N_24682,N_17668,N_19665);
nor U24683 (N_24683,N_17240,N_19889);
nor U24684 (N_24684,N_17411,N_18615);
and U24685 (N_24685,N_17109,N_17044);
nand U24686 (N_24686,N_19754,N_19513);
nand U24687 (N_24687,N_15281,N_18413);
and U24688 (N_24688,N_18598,N_17121);
nor U24689 (N_24689,N_15066,N_16427);
xor U24690 (N_24690,N_15563,N_15810);
nor U24691 (N_24691,N_15891,N_19494);
xnor U24692 (N_24692,N_16211,N_18279);
nor U24693 (N_24693,N_15724,N_17976);
and U24694 (N_24694,N_18692,N_17469);
nand U24695 (N_24695,N_19012,N_17525);
or U24696 (N_24696,N_19305,N_16668);
or U24697 (N_24697,N_19860,N_17170);
nor U24698 (N_24698,N_18835,N_15051);
xor U24699 (N_24699,N_17275,N_17025);
xor U24700 (N_24700,N_15199,N_18966);
nand U24701 (N_24701,N_15082,N_15871);
nand U24702 (N_24702,N_15255,N_16746);
xor U24703 (N_24703,N_16181,N_19622);
nand U24704 (N_24704,N_17779,N_19482);
nor U24705 (N_24705,N_15173,N_18291);
or U24706 (N_24706,N_19820,N_15184);
nand U24707 (N_24707,N_18644,N_16660);
nand U24708 (N_24708,N_17264,N_19223);
nor U24709 (N_24709,N_15725,N_16407);
or U24710 (N_24710,N_15957,N_15450);
nand U24711 (N_24711,N_16582,N_17567);
or U24712 (N_24712,N_16866,N_18941);
nor U24713 (N_24713,N_19972,N_17235);
nand U24714 (N_24714,N_15279,N_17736);
or U24715 (N_24715,N_16290,N_19995);
nor U24716 (N_24716,N_19414,N_19356);
nand U24717 (N_24717,N_17591,N_18297);
nor U24718 (N_24718,N_19277,N_16557);
nor U24719 (N_24719,N_16208,N_16457);
or U24720 (N_24720,N_16851,N_15914);
nand U24721 (N_24721,N_15320,N_18760);
nor U24722 (N_24722,N_16428,N_16814);
and U24723 (N_24723,N_15446,N_17246);
and U24724 (N_24724,N_16604,N_16607);
xor U24725 (N_24725,N_19882,N_17142);
nand U24726 (N_24726,N_15125,N_17063);
nor U24727 (N_24727,N_17040,N_15256);
and U24728 (N_24728,N_17646,N_15156);
xnor U24729 (N_24729,N_19006,N_15979);
or U24730 (N_24730,N_15370,N_17946);
and U24731 (N_24731,N_16290,N_15398);
and U24732 (N_24732,N_17083,N_19825);
and U24733 (N_24733,N_16759,N_16021);
nand U24734 (N_24734,N_17403,N_19436);
nand U24735 (N_24735,N_15310,N_16827);
xor U24736 (N_24736,N_18142,N_16616);
and U24737 (N_24737,N_17716,N_16707);
nand U24738 (N_24738,N_17602,N_18264);
and U24739 (N_24739,N_19805,N_19299);
nand U24740 (N_24740,N_18539,N_15390);
xnor U24741 (N_24741,N_19598,N_16239);
nand U24742 (N_24742,N_19086,N_15968);
nand U24743 (N_24743,N_17251,N_19617);
nor U24744 (N_24744,N_15413,N_16256);
nand U24745 (N_24745,N_19023,N_15026);
or U24746 (N_24746,N_16474,N_17516);
xor U24747 (N_24747,N_15034,N_17584);
and U24748 (N_24748,N_18012,N_16305);
nor U24749 (N_24749,N_19920,N_17002);
xor U24750 (N_24750,N_16882,N_18024);
xor U24751 (N_24751,N_18863,N_15788);
nor U24752 (N_24752,N_15107,N_18524);
or U24753 (N_24753,N_17981,N_16135);
nand U24754 (N_24754,N_19118,N_19851);
nor U24755 (N_24755,N_17458,N_15215);
xor U24756 (N_24756,N_17738,N_18191);
xor U24757 (N_24757,N_17479,N_18894);
nand U24758 (N_24758,N_19665,N_17295);
xnor U24759 (N_24759,N_16867,N_17550);
nand U24760 (N_24760,N_16230,N_16606);
or U24761 (N_24761,N_15361,N_16761);
or U24762 (N_24762,N_18059,N_19164);
nand U24763 (N_24763,N_16080,N_15131);
or U24764 (N_24764,N_15815,N_16810);
or U24765 (N_24765,N_18100,N_17593);
nand U24766 (N_24766,N_17427,N_16887);
and U24767 (N_24767,N_15342,N_15436);
nor U24768 (N_24768,N_19513,N_17104);
nand U24769 (N_24769,N_19560,N_18219);
xor U24770 (N_24770,N_17378,N_16748);
xor U24771 (N_24771,N_15608,N_18869);
and U24772 (N_24772,N_17591,N_18259);
or U24773 (N_24773,N_17498,N_15818);
and U24774 (N_24774,N_15180,N_16530);
nand U24775 (N_24775,N_17021,N_16726);
and U24776 (N_24776,N_15039,N_18861);
or U24777 (N_24777,N_16377,N_19148);
or U24778 (N_24778,N_17120,N_16046);
and U24779 (N_24779,N_18950,N_16853);
xor U24780 (N_24780,N_17369,N_17241);
nor U24781 (N_24781,N_19680,N_16178);
xnor U24782 (N_24782,N_15058,N_18173);
xnor U24783 (N_24783,N_15967,N_17557);
nor U24784 (N_24784,N_18432,N_15804);
xnor U24785 (N_24785,N_16251,N_18707);
or U24786 (N_24786,N_17537,N_19273);
xor U24787 (N_24787,N_17015,N_17188);
nand U24788 (N_24788,N_16172,N_18993);
nor U24789 (N_24789,N_19493,N_18552);
xnor U24790 (N_24790,N_18809,N_15919);
xnor U24791 (N_24791,N_16220,N_18525);
and U24792 (N_24792,N_19060,N_15334);
nor U24793 (N_24793,N_17791,N_15018);
and U24794 (N_24794,N_19880,N_16836);
nand U24795 (N_24795,N_19357,N_17312);
nor U24796 (N_24796,N_15134,N_16721);
and U24797 (N_24797,N_16130,N_15824);
and U24798 (N_24798,N_19491,N_19713);
or U24799 (N_24799,N_16777,N_17061);
nand U24800 (N_24800,N_16443,N_18498);
xor U24801 (N_24801,N_18651,N_19946);
nor U24802 (N_24802,N_19730,N_17694);
or U24803 (N_24803,N_15260,N_17729);
nand U24804 (N_24804,N_17312,N_19768);
or U24805 (N_24805,N_15728,N_15822);
or U24806 (N_24806,N_17499,N_17520);
or U24807 (N_24807,N_15251,N_17972);
or U24808 (N_24808,N_18389,N_18710);
or U24809 (N_24809,N_16309,N_15419);
nor U24810 (N_24810,N_16748,N_16282);
nor U24811 (N_24811,N_16596,N_15481);
xor U24812 (N_24812,N_17367,N_18316);
xnor U24813 (N_24813,N_18076,N_16177);
or U24814 (N_24814,N_19002,N_19190);
nor U24815 (N_24815,N_18673,N_15268);
xnor U24816 (N_24816,N_15656,N_18590);
nand U24817 (N_24817,N_15100,N_19230);
nand U24818 (N_24818,N_19996,N_15973);
xor U24819 (N_24819,N_18005,N_16360);
and U24820 (N_24820,N_18281,N_16655);
nor U24821 (N_24821,N_17408,N_15062);
or U24822 (N_24822,N_18101,N_16528);
nand U24823 (N_24823,N_16394,N_19930);
nand U24824 (N_24824,N_18315,N_18882);
and U24825 (N_24825,N_15359,N_18514);
nor U24826 (N_24826,N_15440,N_18235);
nand U24827 (N_24827,N_18351,N_17446);
or U24828 (N_24828,N_15884,N_19744);
nand U24829 (N_24829,N_16687,N_16632);
nand U24830 (N_24830,N_19142,N_19516);
xor U24831 (N_24831,N_17762,N_19994);
nor U24832 (N_24832,N_15684,N_15179);
or U24833 (N_24833,N_16932,N_15817);
and U24834 (N_24834,N_19208,N_19657);
or U24835 (N_24835,N_18831,N_17999);
nand U24836 (N_24836,N_16766,N_19004);
and U24837 (N_24837,N_16922,N_16198);
nand U24838 (N_24838,N_17910,N_16726);
or U24839 (N_24839,N_15352,N_18725);
xor U24840 (N_24840,N_18526,N_17277);
xor U24841 (N_24841,N_17401,N_16388);
or U24842 (N_24842,N_16211,N_17274);
nor U24843 (N_24843,N_16402,N_18102);
nor U24844 (N_24844,N_15012,N_17050);
or U24845 (N_24845,N_15344,N_18003);
or U24846 (N_24846,N_16349,N_19248);
nand U24847 (N_24847,N_16978,N_17587);
xor U24848 (N_24848,N_19500,N_15714);
or U24849 (N_24849,N_19223,N_16212);
nor U24850 (N_24850,N_17056,N_16827);
nand U24851 (N_24851,N_18402,N_18304);
and U24852 (N_24852,N_19627,N_17601);
and U24853 (N_24853,N_19113,N_18617);
and U24854 (N_24854,N_16099,N_16238);
xor U24855 (N_24855,N_16462,N_17275);
xnor U24856 (N_24856,N_17787,N_17264);
and U24857 (N_24857,N_15368,N_18146);
xor U24858 (N_24858,N_17276,N_18652);
xnor U24859 (N_24859,N_16259,N_17355);
nand U24860 (N_24860,N_16043,N_16156);
nand U24861 (N_24861,N_19539,N_15970);
and U24862 (N_24862,N_17207,N_19208);
or U24863 (N_24863,N_16768,N_17066);
nand U24864 (N_24864,N_19272,N_17737);
xnor U24865 (N_24865,N_18526,N_17554);
nand U24866 (N_24866,N_19536,N_18244);
and U24867 (N_24867,N_17605,N_17859);
and U24868 (N_24868,N_16727,N_18826);
or U24869 (N_24869,N_15027,N_18417);
or U24870 (N_24870,N_17889,N_15951);
xnor U24871 (N_24871,N_18618,N_18648);
and U24872 (N_24872,N_18144,N_15473);
and U24873 (N_24873,N_19059,N_18799);
or U24874 (N_24874,N_16712,N_18107);
xor U24875 (N_24875,N_18592,N_19781);
nor U24876 (N_24876,N_18954,N_18896);
xor U24877 (N_24877,N_19747,N_15481);
or U24878 (N_24878,N_19807,N_17290);
and U24879 (N_24879,N_17582,N_17863);
xor U24880 (N_24880,N_19590,N_15703);
or U24881 (N_24881,N_17222,N_15126);
nor U24882 (N_24882,N_18142,N_17503);
xor U24883 (N_24883,N_18219,N_16463);
nand U24884 (N_24884,N_19012,N_15138);
nor U24885 (N_24885,N_15248,N_16360);
nor U24886 (N_24886,N_15101,N_19584);
xor U24887 (N_24887,N_17215,N_19169);
xor U24888 (N_24888,N_19728,N_15352);
and U24889 (N_24889,N_15213,N_16825);
and U24890 (N_24890,N_16599,N_15831);
nor U24891 (N_24891,N_19759,N_18291);
or U24892 (N_24892,N_18633,N_18916);
nand U24893 (N_24893,N_17350,N_17551);
xor U24894 (N_24894,N_18607,N_19207);
and U24895 (N_24895,N_17507,N_15586);
nand U24896 (N_24896,N_19323,N_16479);
nand U24897 (N_24897,N_18423,N_15944);
xor U24898 (N_24898,N_19289,N_16046);
nor U24899 (N_24899,N_16240,N_16018);
nand U24900 (N_24900,N_19889,N_19521);
nand U24901 (N_24901,N_19708,N_16279);
nor U24902 (N_24902,N_15830,N_18442);
and U24903 (N_24903,N_18395,N_16029);
and U24904 (N_24904,N_16605,N_19428);
xor U24905 (N_24905,N_17407,N_18701);
nand U24906 (N_24906,N_18989,N_19581);
nor U24907 (N_24907,N_18335,N_16243);
nor U24908 (N_24908,N_16397,N_17985);
or U24909 (N_24909,N_15999,N_19254);
and U24910 (N_24910,N_15429,N_18858);
nand U24911 (N_24911,N_18618,N_18846);
nand U24912 (N_24912,N_18280,N_18738);
nand U24913 (N_24913,N_18507,N_17570);
nand U24914 (N_24914,N_19010,N_16415);
and U24915 (N_24915,N_17943,N_16152);
nor U24916 (N_24916,N_15860,N_19780);
nand U24917 (N_24917,N_19851,N_19727);
nor U24918 (N_24918,N_18651,N_17595);
nand U24919 (N_24919,N_17742,N_17174);
and U24920 (N_24920,N_16061,N_17254);
nand U24921 (N_24921,N_16342,N_18197);
nor U24922 (N_24922,N_16980,N_18806);
xnor U24923 (N_24923,N_17569,N_19103);
xor U24924 (N_24924,N_17215,N_15026);
xnor U24925 (N_24925,N_15656,N_15381);
or U24926 (N_24926,N_19441,N_17605);
xnor U24927 (N_24927,N_16518,N_17055);
nand U24928 (N_24928,N_17778,N_19851);
and U24929 (N_24929,N_16502,N_16415);
nand U24930 (N_24930,N_16298,N_18789);
and U24931 (N_24931,N_16625,N_15160);
nand U24932 (N_24932,N_15773,N_16095);
and U24933 (N_24933,N_15966,N_15896);
xor U24934 (N_24934,N_16352,N_18259);
and U24935 (N_24935,N_16656,N_16072);
nand U24936 (N_24936,N_19953,N_17815);
or U24937 (N_24937,N_17855,N_17776);
nand U24938 (N_24938,N_19956,N_17849);
and U24939 (N_24939,N_18184,N_18634);
and U24940 (N_24940,N_18507,N_16339);
nor U24941 (N_24941,N_18326,N_16719);
xor U24942 (N_24942,N_18878,N_19537);
nand U24943 (N_24943,N_15487,N_19480);
and U24944 (N_24944,N_18237,N_18880);
or U24945 (N_24945,N_18903,N_15050);
nor U24946 (N_24946,N_16836,N_15707);
and U24947 (N_24947,N_15712,N_19058);
or U24948 (N_24948,N_19552,N_16218);
and U24949 (N_24949,N_16357,N_19733);
or U24950 (N_24950,N_17223,N_16230);
xor U24951 (N_24951,N_15717,N_15887);
nor U24952 (N_24952,N_15171,N_15635);
xor U24953 (N_24953,N_19120,N_16842);
nand U24954 (N_24954,N_17622,N_16859);
and U24955 (N_24955,N_19419,N_19099);
or U24956 (N_24956,N_15609,N_18284);
or U24957 (N_24957,N_18777,N_15639);
and U24958 (N_24958,N_18477,N_18028);
or U24959 (N_24959,N_19408,N_17557);
nor U24960 (N_24960,N_15501,N_18123);
nand U24961 (N_24961,N_18670,N_18658);
nand U24962 (N_24962,N_18449,N_15920);
nand U24963 (N_24963,N_17380,N_16878);
and U24964 (N_24964,N_18165,N_19155);
and U24965 (N_24965,N_19300,N_18811);
and U24966 (N_24966,N_18897,N_16501);
nor U24967 (N_24967,N_19082,N_17887);
nor U24968 (N_24968,N_19884,N_18033);
xor U24969 (N_24969,N_17300,N_15058);
and U24970 (N_24970,N_16247,N_19522);
nor U24971 (N_24971,N_16681,N_17162);
xor U24972 (N_24972,N_17469,N_17859);
and U24973 (N_24973,N_17922,N_19897);
and U24974 (N_24974,N_15725,N_15127);
xnor U24975 (N_24975,N_16836,N_17268);
xor U24976 (N_24976,N_19789,N_17121);
nor U24977 (N_24977,N_15907,N_15765);
or U24978 (N_24978,N_15437,N_16256);
or U24979 (N_24979,N_15437,N_15077);
nand U24980 (N_24980,N_18583,N_18644);
and U24981 (N_24981,N_17517,N_17794);
xnor U24982 (N_24982,N_15115,N_18400);
xor U24983 (N_24983,N_19320,N_15769);
or U24984 (N_24984,N_17542,N_19434);
nand U24985 (N_24985,N_18828,N_15654);
and U24986 (N_24986,N_19012,N_18117);
xor U24987 (N_24987,N_19518,N_17272);
and U24988 (N_24988,N_16797,N_18971);
nand U24989 (N_24989,N_18548,N_15854);
nand U24990 (N_24990,N_15863,N_15322);
or U24991 (N_24991,N_17099,N_16061);
or U24992 (N_24992,N_16279,N_15735);
and U24993 (N_24993,N_18407,N_18965);
and U24994 (N_24994,N_17196,N_16162);
nor U24995 (N_24995,N_17174,N_19602);
nor U24996 (N_24996,N_18062,N_15739);
nor U24997 (N_24997,N_19407,N_19429);
or U24998 (N_24998,N_18600,N_15723);
nor U24999 (N_24999,N_15760,N_16207);
nor U25000 (N_25000,N_22077,N_23659);
nand U25001 (N_25001,N_22112,N_21623);
xor U25002 (N_25002,N_24030,N_22211);
and U25003 (N_25003,N_22577,N_21522);
nor U25004 (N_25004,N_22875,N_22068);
nand U25005 (N_25005,N_23405,N_23029);
and U25006 (N_25006,N_21191,N_22969);
or U25007 (N_25007,N_20878,N_21661);
nand U25008 (N_25008,N_24973,N_21095);
or U25009 (N_25009,N_24557,N_23543);
or U25010 (N_25010,N_20436,N_23627);
nor U25011 (N_25011,N_20740,N_23179);
xor U25012 (N_25012,N_21181,N_20872);
or U25013 (N_25013,N_22223,N_24064);
nand U25014 (N_25014,N_24478,N_20724);
nor U25015 (N_25015,N_22162,N_22553);
nand U25016 (N_25016,N_21107,N_20335);
and U25017 (N_25017,N_20081,N_20080);
or U25018 (N_25018,N_21889,N_21658);
and U25019 (N_25019,N_24495,N_24221);
and U25020 (N_25020,N_20836,N_20101);
and U25021 (N_25021,N_23960,N_24648);
and U25022 (N_25022,N_23195,N_21897);
or U25023 (N_25023,N_22871,N_20452);
nand U25024 (N_25024,N_21744,N_20782);
nand U25025 (N_25025,N_24363,N_22096);
nor U25026 (N_25026,N_24271,N_21621);
and U25027 (N_25027,N_21737,N_24901);
and U25028 (N_25028,N_23370,N_23497);
or U25029 (N_25029,N_21323,N_22898);
and U25030 (N_25030,N_20131,N_21740);
xnor U25031 (N_25031,N_20545,N_24402);
or U25032 (N_25032,N_24302,N_20146);
or U25033 (N_25033,N_21784,N_24105);
nand U25034 (N_25034,N_20366,N_24849);
nand U25035 (N_25035,N_22457,N_23315);
nor U25036 (N_25036,N_21531,N_24425);
nand U25037 (N_25037,N_21468,N_21019);
nor U25038 (N_25038,N_23902,N_24250);
xor U25039 (N_25039,N_23621,N_24460);
nor U25040 (N_25040,N_21304,N_21464);
xnor U25041 (N_25041,N_22115,N_21482);
and U25042 (N_25042,N_22637,N_22870);
xor U25043 (N_25043,N_20443,N_24654);
nor U25044 (N_25044,N_21410,N_21388);
xor U25045 (N_25045,N_21115,N_20293);
nand U25046 (N_25046,N_24787,N_21838);
nand U25047 (N_25047,N_20241,N_21617);
and U25048 (N_25048,N_23159,N_24895);
and U25049 (N_25049,N_20446,N_21865);
xor U25050 (N_25050,N_23015,N_22675);
or U25051 (N_25051,N_22347,N_24696);
nand U25052 (N_25052,N_22084,N_21079);
and U25053 (N_25053,N_22722,N_24407);
or U25054 (N_25054,N_24760,N_22177);
and U25055 (N_25055,N_20244,N_24087);
or U25056 (N_25056,N_24524,N_20767);
and U25057 (N_25057,N_22323,N_22657);
xor U25058 (N_25058,N_24333,N_23149);
nand U25059 (N_25059,N_23496,N_21842);
nand U25060 (N_25060,N_24988,N_24780);
and U25061 (N_25061,N_21805,N_20458);
xor U25062 (N_25062,N_24285,N_21277);
nand U25063 (N_25063,N_20199,N_20213);
or U25064 (N_25064,N_22137,N_21519);
nor U25065 (N_25065,N_23866,N_22534);
nand U25066 (N_25066,N_22756,N_21825);
xor U25067 (N_25067,N_22865,N_23601);
nor U25068 (N_25068,N_20262,N_21158);
xnor U25069 (N_25069,N_22779,N_24542);
nor U25070 (N_25070,N_23057,N_21972);
nor U25071 (N_25071,N_22676,N_23792);
and U25072 (N_25072,N_24486,N_21807);
nor U25073 (N_25073,N_20853,N_24739);
xor U25074 (N_25074,N_21993,N_20790);
nor U25075 (N_25075,N_23754,N_23938);
and U25076 (N_25076,N_23335,N_24723);
xnor U25077 (N_25077,N_23797,N_20686);
nor U25078 (N_25078,N_24532,N_24303);
xor U25079 (N_25079,N_20840,N_22951);
nand U25080 (N_25080,N_22046,N_21895);
nor U25081 (N_25081,N_20587,N_20550);
nand U25082 (N_25082,N_24949,N_22488);
nor U25083 (N_25083,N_22814,N_24987);
nand U25084 (N_25084,N_20104,N_21969);
or U25085 (N_25085,N_24931,N_20772);
and U25086 (N_25086,N_23073,N_20763);
or U25087 (N_25087,N_23908,N_20385);
and U25088 (N_25088,N_22655,N_23036);
or U25089 (N_25089,N_20169,N_23889);
or U25090 (N_25090,N_21463,N_20417);
nor U25091 (N_25091,N_23986,N_23401);
xor U25092 (N_25092,N_20312,N_22933);
nor U25093 (N_25093,N_21384,N_22069);
xor U25094 (N_25094,N_23258,N_23012);
nand U25095 (N_25095,N_21274,N_20697);
nand U25096 (N_25096,N_21843,N_22689);
and U25097 (N_25097,N_20832,N_23626);
and U25098 (N_25098,N_20347,N_24602);
nand U25099 (N_25099,N_22558,N_24911);
xor U25100 (N_25100,N_20793,N_23848);
xnor U25101 (N_25101,N_22308,N_21440);
and U25102 (N_25102,N_23502,N_21875);
nor U25103 (N_25103,N_23357,N_22428);
nand U25104 (N_25104,N_23194,N_22330);
nand U25105 (N_25105,N_22463,N_21713);
xor U25106 (N_25106,N_24024,N_21092);
xnor U25107 (N_25107,N_22582,N_22009);
nand U25108 (N_25108,N_21222,N_23577);
xor U25109 (N_25109,N_20970,N_20829);
and U25110 (N_25110,N_20507,N_21885);
and U25111 (N_25111,N_21218,N_24625);
and U25112 (N_25112,N_22809,N_24669);
nand U25113 (N_25113,N_21141,N_20844);
nand U25114 (N_25114,N_22302,N_23612);
and U25115 (N_25115,N_22705,N_21203);
and U25116 (N_25116,N_22060,N_21801);
and U25117 (N_25117,N_23756,N_20180);
nor U25118 (N_25118,N_21930,N_24375);
nand U25119 (N_25119,N_23717,N_21999);
or U25120 (N_25120,N_21917,N_24698);
nand U25121 (N_25121,N_23514,N_23520);
or U25122 (N_25122,N_23956,N_21536);
nor U25123 (N_25123,N_22277,N_24069);
and U25124 (N_25124,N_23487,N_23450);
nand U25125 (N_25125,N_24543,N_20694);
nand U25126 (N_25126,N_21524,N_24481);
or U25127 (N_25127,N_21876,N_20463);
or U25128 (N_25128,N_22087,N_20998);
xnor U25129 (N_25129,N_23298,N_24762);
or U25130 (N_25130,N_22314,N_22994);
xnor U25131 (N_25131,N_22250,N_21105);
xor U25132 (N_25132,N_23834,N_21725);
or U25133 (N_25133,N_21852,N_24392);
xor U25134 (N_25134,N_22189,N_24266);
nor U25135 (N_25135,N_24096,N_22884);
and U25136 (N_25136,N_22480,N_21287);
or U25137 (N_25137,N_20562,N_24045);
or U25138 (N_25138,N_22670,N_20257);
nor U25139 (N_25139,N_22734,N_21403);
and U25140 (N_25140,N_22808,N_21421);
nand U25141 (N_25141,N_24537,N_20392);
and U25142 (N_25142,N_24256,N_24996);
nand U25143 (N_25143,N_24152,N_20026);
or U25144 (N_25144,N_21049,N_22325);
nor U25145 (N_25145,N_22861,N_20828);
and U25146 (N_25146,N_23861,N_20308);
xor U25147 (N_25147,N_23457,N_24245);
xor U25148 (N_25148,N_23019,N_23969);
nor U25149 (N_25149,N_22590,N_22263);
nand U25150 (N_25150,N_24829,N_23837);
nand U25151 (N_25151,N_23638,N_24844);
and U25152 (N_25152,N_22167,N_21698);
and U25153 (N_25153,N_23064,N_21830);
xor U25154 (N_25154,N_24977,N_23417);
nand U25155 (N_25155,N_23273,N_21159);
xnor U25156 (N_25156,N_24730,N_22632);
or U25157 (N_25157,N_23894,N_20179);
or U25158 (N_25158,N_22392,N_20181);
and U25159 (N_25159,N_24210,N_20154);
or U25160 (N_25160,N_24047,N_20904);
and U25161 (N_25161,N_21562,N_23874);
or U25162 (N_25162,N_23527,N_21848);
nand U25163 (N_25163,N_22158,N_23117);
nand U25164 (N_25164,N_20353,N_21899);
nor U25165 (N_25165,N_20886,N_24244);
xor U25166 (N_25166,N_24709,N_20999);
nor U25167 (N_25167,N_23016,N_23504);
nor U25168 (N_25168,N_21321,N_22944);
xnor U25169 (N_25169,N_22486,N_24450);
or U25170 (N_25170,N_23415,N_22171);
nand U25171 (N_25171,N_21393,N_23014);
xnor U25172 (N_25172,N_21090,N_21392);
nand U25173 (N_25173,N_23248,N_21035);
nor U25174 (N_25174,N_22145,N_21634);
and U25175 (N_25175,N_20119,N_23860);
xor U25176 (N_25176,N_21340,N_22608);
nor U25177 (N_25177,N_22617,N_23740);
xor U25178 (N_25178,N_20289,N_22236);
nand U25179 (N_25179,N_24420,N_22134);
and U25180 (N_25180,N_20135,N_21770);
or U25181 (N_25181,N_24902,N_20265);
or U25182 (N_25182,N_24865,N_21777);
or U25183 (N_25183,N_22672,N_23446);
and U25184 (N_25184,N_22749,N_21868);
and U25185 (N_25185,N_24493,N_20093);
xor U25186 (N_25186,N_21366,N_23699);
or U25187 (N_25187,N_21619,N_21127);
xnor U25188 (N_25188,N_22292,N_20382);
or U25189 (N_25189,N_20040,N_21037);
and U25190 (N_25190,N_24139,N_20136);
or U25191 (N_25191,N_21234,N_21592);
nor U25192 (N_25192,N_23851,N_20845);
nor U25193 (N_25193,N_20612,N_24784);
nor U25194 (N_25194,N_20792,N_20727);
and U25195 (N_25195,N_23759,N_23269);
xor U25196 (N_25196,N_21196,N_23210);
xor U25197 (N_25197,N_24428,N_23047);
xnor U25198 (N_25198,N_21541,N_22121);
and U25199 (N_25199,N_22337,N_20705);
nand U25200 (N_25200,N_20687,N_23570);
nand U25201 (N_25201,N_24324,N_21966);
nand U25202 (N_25202,N_24126,N_21017);
nor U25203 (N_25203,N_23259,N_20752);
nand U25204 (N_25204,N_21462,N_21611);
and U25205 (N_25205,N_23686,N_24388);
or U25206 (N_25206,N_23167,N_24222);
or U25207 (N_25207,N_24797,N_20653);
nor U25208 (N_25208,N_24362,N_23979);
nand U25209 (N_25209,N_23827,N_23312);
and U25210 (N_25210,N_21227,N_23286);
nand U25211 (N_25211,N_20590,N_20660);
xnor U25212 (N_25212,N_22980,N_23443);
and U25213 (N_25213,N_23639,N_23785);
xor U25214 (N_25214,N_23013,N_20586);
nand U25215 (N_25215,N_20130,N_21702);
xor U25216 (N_25216,N_22927,N_20654);
xor U25217 (N_25217,N_21820,N_23252);
nor U25218 (N_25218,N_20150,N_23051);
or U25219 (N_25219,N_22587,N_24397);
nor U25220 (N_25220,N_24513,N_24234);
nand U25221 (N_25221,N_24112,N_24611);
nor U25222 (N_25222,N_24062,N_21664);
or U25223 (N_25223,N_22197,N_20977);
nor U25224 (N_25224,N_21850,N_21670);
nor U25225 (N_25225,N_22479,N_24231);
nor U25226 (N_25226,N_20923,N_21282);
and U25227 (N_25227,N_24135,N_22882);
or U25228 (N_25228,N_20006,N_20028);
nand U25229 (N_25229,N_23731,N_20585);
or U25230 (N_25230,N_24395,N_21719);
and U25231 (N_25231,N_23421,N_24377);
nor U25232 (N_25232,N_24845,N_21232);
and U25233 (N_25233,N_20937,N_23566);
or U25234 (N_25234,N_23384,N_20796);
or U25235 (N_25235,N_23964,N_22199);
xor U25236 (N_25236,N_21788,N_20336);
and U25237 (N_25237,N_21004,N_24954);
xnor U25238 (N_25238,N_20144,N_20561);
nor U25239 (N_25239,N_24852,N_22526);
nor U25240 (N_25240,N_24641,N_24485);
or U25241 (N_25241,N_22957,N_23449);
and U25242 (N_25242,N_20574,N_20061);
xnor U25243 (N_25243,N_23327,N_23313);
nand U25244 (N_25244,N_24141,N_22033);
nor U25245 (N_25245,N_20079,N_22748);
nor U25246 (N_25246,N_23316,N_22058);
nand U25247 (N_25247,N_22915,N_21047);
nor U25248 (N_25248,N_24243,N_20641);
and U25249 (N_25249,N_21577,N_20188);
and U25250 (N_25250,N_21046,N_23550);
and U25251 (N_25251,N_22938,N_22713);
nand U25252 (N_25252,N_21109,N_22108);
xor U25253 (N_25253,N_21665,N_21292);
nand U25254 (N_25254,N_21691,N_24410);
nor U25255 (N_25255,N_20221,N_23505);
nand U25256 (N_25256,N_23828,N_23204);
xnor U25257 (N_25257,N_24474,N_23152);
nor U25258 (N_25258,N_22037,N_20487);
and U25259 (N_25259,N_24384,N_21708);
nor U25260 (N_25260,N_23977,N_24389);
xnor U25261 (N_25261,N_23809,N_21439);
nor U25262 (N_25262,N_20295,N_21923);
and U25263 (N_25263,N_23360,N_20126);
nand U25264 (N_25264,N_23276,N_23791);
nand U25265 (N_25265,N_20378,N_21826);
and U25266 (N_25266,N_20598,N_21666);
or U25267 (N_25267,N_23773,N_22328);
or U25268 (N_25268,N_22436,N_23736);
and U25269 (N_25269,N_20432,N_21925);
and U25270 (N_25270,N_23092,N_23083);
nor U25271 (N_25271,N_24693,N_21961);
xnor U25272 (N_25272,N_24079,N_23371);
or U25273 (N_25273,N_23530,N_24970);
nor U25274 (N_25274,N_23649,N_21678);
or U25275 (N_25275,N_22547,N_23491);
nand U25276 (N_25276,N_24885,N_24137);
nand U25277 (N_25277,N_22821,N_24355);
or U25278 (N_25278,N_23741,N_20916);
nand U25279 (N_25279,N_22702,N_22811);
or U25280 (N_25280,N_22209,N_23200);
nand U25281 (N_25281,N_21779,N_21030);
nor U25282 (N_25282,N_23536,N_21609);
and U25283 (N_25283,N_22922,N_22173);
nor U25284 (N_25284,N_22403,N_20622);
xor U25285 (N_25285,N_23030,N_21832);
nor U25286 (N_25286,N_22007,N_20901);
or U25287 (N_25287,N_20311,N_24429);
or U25288 (N_25288,N_22901,N_24744);
nand U25289 (N_25289,N_21310,N_24640);
or U25290 (N_25290,N_20237,N_23905);
and U25291 (N_25291,N_21990,N_24414);
nor U25292 (N_25292,N_23589,N_24813);
nand U25293 (N_25293,N_24861,N_24989);
nand U25294 (N_25294,N_24496,N_21087);
and U25295 (N_25295,N_21921,N_21810);
nand U25296 (N_25296,N_24775,N_23021);
and U25297 (N_25297,N_20978,N_23478);
xor U25298 (N_25298,N_24118,N_22570);
and U25299 (N_25299,N_22303,N_21721);
xor U25300 (N_25300,N_22647,N_20368);
or U25301 (N_25301,N_20332,N_24707);
and U25302 (N_25302,N_22257,N_24461);
and U25303 (N_25303,N_24609,N_20020);
nor U25304 (N_25304,N_22150,N_20468);
and U25305 (N_25305,N_23783,N_22110);
or U25306 (N_25306,N_23533,N_23482);
and U25307 (N_25307,N_24874,N_21627);
xor U25308 (N_25308,N_20220,N_23913);
xnor U25309 (N_25309,N_23281,N_23615);
nand U25310 (N_25310,N_23087,N_23642);
nor U25311 (N_25311,N_21904,N_24074);
nor U25312 (N_25312,N_23148,N_23375);
xnor U25313 (N_25313,N_23600,N_23681);
or U25314 (N_25314,N_21839,N_22109);
xnor U25315 (N_25315,N_24722,N_20616);
and U25316 (N_25316,N_22213,N_24512);
nor U25317 (N_25317,N_22612,N_24624);
and U25318 (N_25318,N_22379,N_21717);
nor U25319 (N_25319,N_24253,N_23723);
xnor U25320 (N_25320,N_23414,N_21612);
and U25321 (N_25321,N_24804,N_22196);
or U25322 (N_25322,N_23279,N_20866);
or U25323 (N_25323,N_24915,N_24751);
nand U25324 (N_25324,N_23843,N_22498);
xor U25325 (N_25325,N_21007,N_21906);
xor U25326 (N_25326,N_21856,N_23939);
or U25327 (N_25327,N_20873,N_21279);
xor U25328 (N_25328,N_21703,N_20320);
and U25329 (N_25329,N_24568,N_20500);
nand U25330 (N_25330,N_22508,N_20594);
nor U25331 (N_25331,N_21135,N_24825);
nor U25332 (N_25332,N_22664,N_22783);
and U25333 (N_25333,N_20214,N_23944);
and U25334 (N_25334,N_23136,N_21437);
or U25335 (N_25335,N_21244,N_23872);
nand U25336 (N_25336,N_23216,N_22846);
nor U25337 (N_25337,N_23169,N_20953);
nand U25338 (N_25338,N_21767,N_23932);
or U25339 (N_25339,N_24867,N_24608);
nor U25340 (N_25340,N_21422,N_20483);
nand U25341 (N_25341,N_24046,N_24835);
or U25342 (N_25342,N_23698,N_21778);
and U25343 (N_25343,N_24431,N_22299);
or U25344 (N_25344,N_22188,N_20551);
nor U25345 (N_25345,N_23277,N_20471);
and U25346 (N_25346,N_22831,N_22304);
and U25347 (N_25347,N_23048,N_23285);
xnor U25348 (N_25348,N_21742,N_24717);
or U25349 (N_25349,N_24948,N_23166);
nor U25350 (N_25350,N_23336,N_22170);
and U25351 (N_25351,N_22184,N_21916);
or U25352 (N_25352,N_20063,N_23150);
nand U25353 (N_25353,N_23321,N_24016);
and U25354 (N_25354,N_20038,N_23374);
or U25355 (N_25355,N_21204,N_21846);
and U25356 (N_25356,N_24765,N_24048);
and U25357 (N_25357,N_21359,N_20636);
or U25358 (N_25358,N_22111,N_20083);
and U25359 (N_25359,N_23614,N_24863);
nand U25360 (N_25360,N_23934,N_23107);
or U25361 (N_25361,N_20331,N_23155);
xnor U25362 (N_25362,N_21579,N_24439);
xor U25363 (N_25363,N_23387,N_23547);
and U25364 (N_25364,N_23024,N_21919);
or U25365 (N_25365,N_23311,N_20802);
or U25366 (N_25366,N_23856,N_22684);
or U25367 (N_25367,N_22414,N_21532);
nor U25368 (N_25368,N_23096,N_22425);
and U25369 (N_25369,N_22646,N_20976);
nand U25370 (N_25370,N_20785,N_21450);
xnor U25371 (N_25371,N_23531,N_22850);
nor U25372 (N_25372,N_23060,N_22371);
xnor U25373 (N_25373,N_21281,N_20429);
or U25374 (N_25374,N_20075,N_23299);
nor U25375 (N_25375,N_20389,N_21589);
nand U25376 (N_25376,N_21419,N_24465);
or U25377 (N_25377,N_22470,N_22475);
nand U25378 (N_25378,N_24349,N_24033);
nor U25379 (N_25379,N_23873,N_20909);
nor U25380 (N_25380,N_20245,N_23924);
and U25381 (N_25381,N_23690,N_21513);
xnor U25382 (N_25382,N_22047,N_22345);
and U25383 (N_25383,N_21759,N_22389);
xor U25384 (N_25384,N_23461,N_23137);
nand U25385 (N_25385,N_24031,N_22653);
nand U25386 (N_25386,N_23199,N_20987);
xnor U25387 (N_25387,N_20486,N_22563);
nand U25388 (N_25388,N_22700,N_24019);
xor U25389 (N_25389,N_20372,N_20750);
and U25390 (N_25390,N_23193,N_20659);
nand U25391 (N_25391,N_21414,N_22910);
and U25392 (N_25392,N_22273,N_22717);
or U25393 (N_25393,N_21153,N_21991);
and U25394 (N_25394,N_23483,N_20924);
xor U25395 (N_25395,N_20008,N_23326);
nor U25396 (N_25396,N_24077,N_22388);
xor U25397 (N_25397,N_24358,N_20548);
or U25398 (N_25398,N_23746,N_20018);
nand U25399 (N_25399,N_24847,N_23126);
nand U25400 (N_25400,N_21256,N_21508);
or U25401 (N_25401,N_24357,N_20175);
nor U25402 (N_25402,N_23814,N_22285);
nand U25403 (N_25403,N_23810,N_20867);
and U25404 (N_25404,N_20068,N_23781);
or U25405 (N_25405,N_21710,N_24866);
nand U25406 (N_25406,N_24567,N_23043);
or U25407 (N_25407,N_21962,N_24583);
xor U25408 (N_25408,N_20954,N_24672);
nor U25409 (N_25409,N_21045,N_24216);
nor U25410 (N_25410,N_21453,N_21834);
nand U25411 (N_25411,N_20291,N_24193);
nand U25412 (N_25412,N_22810,N_24712);
xnor U25413 (N_25413,N_24035,N_24771);
nor U25414 (N_25414,N_20108,N_24904);
or U25415 (N_25415,N_21268,N_20495);
and U25416 (N_25416,N_24889,N_24111);
xor U25417 (N_25417,N_24555,N_23465);
nor U25418 (N_25418,N_23314,N_23996);
xor U25419 (N_25419,N_24589,N_21479);
nand U25420 (N_25420,N_20670,N_24251);
or U25421 (N_25421,N_20158,N_21566);
nand U25422 (N_25422,N_24032,N_24716);
and U25423 (N_25423,N_21913,N_23796);
nand U25424 (N_25424,N_22075,N_21072);
and U25425 (N_25425,N_21510,N_20023);
nand U25426 (N_25426,N_20190,N_22605);
nand U25427 (N_25427,N_23661,N_23474);
or U25428 (N_25428,N_21053,N_23056);
and U25429 (N_25429,N_21616,N_24459);
or U25430 (N_25430,N_22244,N_24345);
or U25431 (N_25431,N_20677,N_21675);
nor U25432 (N_25432,N_22911,N_23629);
nand U25433 (N_25433,N_21251,N_21442);
or U25434 (N_25434,N_23767,N_24790);
nor U25435 (N_25435,N_20920,N_24725);
nor U25436 (N_25436,N_23140,N_24470);
nor U25437 (N_25437,N_20635,N_24212);
nand U25438 (N_25438,N_20688,N_21020);
nor U25439 (N_25439,N_22329,N_22466);
xor U25440 (N_25440,N_22923,N_21647);
and U25441 (N_25441,N_20459,N_24873);
nand U25442 (N_25442,N_24463,N_23282);
nor U25443 (N_25443,N_22286,N_20882);
nor U25444 (N_25444,N_23352,N_23005);
xor U25445 (N_25445,N_23609,N_23693);
nand U25446 (N_25446,N_23617,N_22430);
or U25447 (N_25447,N_23081,N_21455);
and U25448 (N_25448,N_23115,N_22573);
xor U25449 (N_25449,N_23708,N_23270);
and U25450 (N_25450,N_24953,N_24556);
xor U25451 (N_25451,N_23841,N_20222);
xnor U25452 (N_25452,N_24365,N_24014);
or U25453 (N_25453,N_20435,N_20485);
or U25454 (N_25454,N_22863,N_23825);
or U25455 (N_25455,N_24795,N_21835);
nor U25456 (N_25456,N_21174,N_22198);
nor U25457 (N_25457,N_23729,N_21111);
xor U25458 (N_25458,N_20098,N_23309);
nor U25459 (N_25459,N_22505,N_23066);
or U25460 (N_25460,N_20896,N_23607);
and U25461 (N_25461,N_22791,N_21938);
nand U25462 (N_25462,N_24667,N_23662);
and U25463 (N_25463,N_23368,N_24788);
or U25464 (N_25464,N_22950,N_23509);
nand U25465 (N_25465,N_20555,N_21207);
nand U25466 (N_25466,N_23808,N_20810);
xnor U25467 (N_25467,N_23528,N_23422);
nand U25468 (N_25468,N_22954,N_24971);
nand U25469 (N_25469,N_24314,N_24518);
xor U25470 (N_25470,N_22165,N_22409);
nand U25471 (N_25471,N_21382,N_24263);
or U25472 (N_25472,N_22574,N_20690);
nand U25473 (N_25473,N_20082,N_24536);
nor U25474 (N_25474,N_21354,N_23634);
nor U25475 (N_25475,N_23393,N_21803);
nand U25476 (N_25476,N_22694,N_24356);
and U25477 (N_25477,N_21341,N_23963);
and U25478 (N_25478,N_21771,N_24163);
xnor U25479 (N_25479,N_23588,N_24080);
or U25480 (N_25480,N_20152,N_20111);
and U25481 (N_25481,N_23748,N_21747);
and U25482 (N_25482,N_22730,N_21684);
xnor U25483 (N_25483,N_23613,N_24644);
nor U25484 (N_25484,N_23557,N_20593);
or U25485 (N_25485,N_21168,N_20031);
or U25486 (N_25486,N_22906,N_21996);
and U25487 (N_25487,N_22799,N_21029);
or U25488 (N_25488,N_24063,N_20379);
nor U25489 (N_25489,N_22456,N_23998);
nand U25490 (N_25490,N_21569,N_22130);
and U25491 (N_25491,N_21833,N_21027);
nor U25492 (N_25492,N_22829,N_24617);
nor U25493 (N_25493,N_20720,N_24133);
or U25494 (N_25494,N_24480,N_20538);
and U25495 (N_25495,N_23477,N_20890);
nor U25496 (N_25496,N_20666,N_21161);
nor U25497 (N_25497,N_22970,N_20713);
or U25498 (N_25498,N_20974,N_20167);
nand U25499 (N_25499,N_20558,N_20835);
or U25500 (N_25500,N_22500,N_20238);
nand U25501 (N_25501,N_24295,N_22588);
nor U25502 (N_25502,N_23804,N_22815);
nand U25503 (N_25503,N_21346,N_21436);
and U25504 (N_25504,N_21498,N_20854);
or U25505 (N_25505,N_24763,N_20980);
nand U25506 (N_25506,N_22659,N_20667);
nor U25507 (N_25507,N_23685,N_21599);
nor U25508 (N_25508,N_21097,N_23596);
nor U25509 (N_25509,N_24441,N_21413);
nand U25510 (N_25510,N_20386,N_21379);
and U25511 (N_25511,N_23217,N_24299);
nand U25512 (N_25512,N_23124,N_23416);
nand U25513 (N_25513,N_23188,N_20881);
nor U25514 (N_25514,N_24782,N_22258);
nor U25515 (N_25515,N_24142,N_22584);
xnor U25516 (N_25516,N_21098,N_22492);
xor U25517 (N_25517,N_21963,N_24196);
xor U25518 (N_25518,N_24892,N_22073);
and U25519 (N_25519,N_23896,N_24595);
or U25520 (N_25520,N_23683,N_21145);
nand U25521 (N_25521,N_23991,N_22390);
or U25522 (N_25522,N_21016,N_22270);
xor U25523 (N_25523,N_24727,N_20437);
or U25524 (N_25524,N_20683,N_21270);
and U25525 (N_25525,N_21984,N_21061);
xor U25526 (N_25526,N_22971,N_23039);
or U25527 (N_25527,N_22455,N_24191);
nor U25528 (N_25528,N_22999,N_23209);
and U25529 (N_25529,N_20755,N_21223);
or U25530 (N_25530,N_23215,N_22163);
and U25531 (N_25531,N_21014,N_21142);
nor U25532 (N_25532,N_21504,N_21150);
and U25533 (N_25533,N_22288,N_20908);
xnor U25534 (N_25534,N_22718,N_22800);
nand U25535 (N_25535,N_24832,N_23914);
nand U25536 (N_25536,N_22493,N_23758);
or U25537 (N_25537,N_21288,N_24296);
or U25538 (N_25538,N_20255,N_22090);
and U25539 (N_25539,N_24412,N_20066);
or U25540 (N_25540,N_21326,N_24129);
nor U25541 (N_25541,N_20849,N_22918);
nand U25542 (N_25542,N_22266,N_21752);
xnor U25543 (N_25543,N_23032,N_23455);
or U25544 (N_25544,N_20807,N_22651);
nand U25545 (N_25545,N_20718,N_21186);
xor U25546 (N_25546,N_21023,N_20505);
or U25547 (N_25547,N_24993,N_23334);
nor U25548 (N_25548,N_24777,N_20887);
xor U25549 (N_25549,N_24379,N_22504);
or U25550 (N_25550,N_21397,N_24753);
xor U25551 (N_25551,N_22805,N_24718);
nand U25552 (N_25552,N_23055,N_21731);
nand U25553 (N_25553,N_23080,N_21652);
and U25554 (N_25554,N_24172,N_24561);
or U25555 (N_25555,N_20742,N_23592);
and U25556 (N_25556,N_21372,N_24878);
xnor U25557 (N_25557,N_24585,N_22751);
nor U25558 (N_25558,N_22208,N_22298);
and U25559 (N_25559,N_20390,N_22464);
or U25560 (N_25560,N_21473,N_23086);
nor U25561 (N_25561,N_21640,N_21307);
and U25562 (N_25562,N_20818,N_20532);
nand U25563 (N_25563,N_21796,N_22529);
xnor U25564 (N_25564,N_23243,N_21474);
nand U25565 (N_25565,N_24802,N_20360);
nor U25566 (N_25566,N_21760,N_22916);
and U25567 (N_25567,N_21171,N_22120);
and U25568 (N_25568,N_20005,N_20399);
nor U25569 (N_25569,N_20036,N_20838);
and U25570 (N_25570,N_22798,N_22804);
and U25571 (N_25571,N_24520,N_22794);
and U25572 (N_25572,N_22294,N_23095);
nand U25573 (N_25573,N_24743,N_20041);
nor U25574 (N_25574,N_23867,N_23189);
and U25575 (N_25575,N_20968,N_24831);
xor U25576 (N_25576,N_24267,N_22233);
or U25577 (N_25577,N_23970,N_23495);
xnor U25578 (N_25578,N_20957,N_21348);
nand U25579 (N_25579,N_24241,N_23244);
nor U25580 (N_25580,N_23234,N_23500);
and U25581 (N_25581,N_21635,N_20025);
xnor U25582 (N_25582,N_22413,N_20692);
or U25583 (N_25583,N_22660,N_22136);
nor U25584 (N_25584,N_20973,N_20618);
xnor U25585 (N_25585,N_20911,N_24714);
nor U25586 (N_25586,N_23308,N_20084);
nand U25587 (N_25587,N_23337,N_20745);
nor U25588 (N_25588,N_21649,N_24012);
or U25589 (N_25589,N_23331,N_24842);
or U25590 (N_25590,N_21021,N_21732);
nand U25591 (N_25591,N_20699,N_22449);
or U25592 (N_25592,N_21163,N_21553);
or U25593 (N_25593,N_22151,N_22194);
nor U25594 (N_25594,N_20613,N_23236);
nor U25595 (N_25595,N_22454,N_20611);
and U25596 (N_25596,N_20303,N_20990);
or U25597 (N_25597,N_20737,N_23839);
xor U25598 (N_25598,N_22393,N_22622);
xnor U25599 (N_25599,N_21249,N_23362);
nand U25600 (N_25600,N_23516,N_21369);
nor U25601 (N_25601,N_22759,N_21815);
and U25602 (N_25602,N_23510,N_20754);
nand U25603 (N_25603,N_20299,N_21615);
nor U25604 (N_25604,N_21633,N_23444);
or U25605 (N_25605,N_21370,N_20578);
nor U25606 (N_25606,N_24034,N_22267);
or U25607 (N_25607,N_23943,N_24446);
nor U25608 (N_25608,N_21264,N_21394);
xor U25609 (N_25609,N_22521,N_22437);
xor U25610 (N_25610,N_21114,N_24664);
xnor U25611 (N_25611,N_20762,N_22406);
xnor U25612 (N_25612,N_22491,N_22474);
and U25613 (N_25613,N_23883,N_23177);
or U25614 (N_25614,N_22958,N_23481);
and U25615 (N_25615,N_23161,N_21642);
or U25616 (N_25616,N_24330,N_22182);
nor U25617 (N_25617,N_21112,N_24290);
nand U25618 (N_25618,N_22041,N_23116);
xor U25619 (N_25619,N_21728,N_20614);
and U25620 (N_25620,N_24565,N_20416);
nor U25621 (N_25621,N_24374,N_21311);
nand U25622 (N_25622,N_21376,N_23595);
xor U25623 (N_25623,N_20283,N_24124);
or U25624 (N_25624,N_20596,N_22978);
or U25625 (N_25625,N_22019,N_23988);
and U25626 (N_25626,N_21028,N_22094);
or U25627 (N_25627,N_23978,N_23396);
xnor U25628 (N_25628,N_23507,N_23870);
and U25629 (N_25629,N_20029,N_22519);
and U25630 (N_25630,N_22074,N_23436);
nand U25631 (N_25631,N_22638,N_21220);
nand U25632 (N_25632,N_24039,N_23485);
xor U25633 (N_25633,N_24060,N_24144);
nand U25634 (N_25634,N_21428,N_21679);
xor U25635 (N_25635,N_22338,N_24909);
nor U25636 (N_25636,N_24675,N_22416);
nand U25637 (N_25637,N_24626,N_23591);
nor U25638 (N_25638,N_24666,N_20609);
xor U25639 (N_25639,N_23853,N_23388);
xor U25640 (N_25640,N_23668,N_20306);
nand U25641 (N_25641,N_23645,N_22309);
xor U25642 (N_25642,N_20044,N_20466);
xnor U25643 (N_25643,N_23999,N_21175);
xnor U25644 (N_25644,N_21094,N_21544);
or U25645 (N_25645,N_20078,N_24899);
or U25646 (N_25646,N_20711,N_21365);
and U25647 (N_25647,N_24383,N_22830);
or U25648 (N_25648,N_21507,N_21631);
nor U25649 (N_25649,N_20634,N_22753);
xor U25650 (N_25650,N_21353,N_20588);
nand U25651 (N_25651,N_23779,N_23636);
or U25652 (N_25652,N_20497,N_23224);
nor U25653 (N_25653,N_20019,N_24690);
xor U25654 (N_25654,N_20339,N_21648);
nand U25655 (N_25655,N_24366,N_24932);
or U25656 (N_25656,N_22912,N_23735);
and U25657 (N_25657,N_21981,N_20058);
or U25658 (N_25658,N_22373,N_20580);
or U25659 (N_25659,N_21718,N_23701);
and U25660 (N_25660,N_20936,N_23876);
or U25661 (N_25661,N_22501,N_23035);
or U25662 (N_25662,N_24442,N_22363);
nand U25663 (N_25663,N_23774,N_24099);
and U25664 (N_25664,N_24018,N_20067);
and U25665 (N_25665,N_20398,N_22443);
and U25666 (N_25666,N_22613,N_24545);
nor U25667 (N_25667,N_22296,N_21862);
xor U25668 (N_25668,N_24289,N_23105);
or U25669 (N_25669,N_21396,N_24136);
or U25670 (N_25670,N_21484,N_23599);
and U25671 (N_25671,N_20138,N_21712);
nor U25672 (N_25672,N_24505,N_20254);
xor U25673 (N_25673,N_20054,N_21550);
nor U25674 (N_25674,N_24403,N_21010);
xor U25675 (N_25675,N_23802,N_22320);
xor U25676 (N_25676,N_21715,N_23673);
nand U25677 (N_25677,N_22966,N_23941);
and U25678 (N_25678,N_21124,N_24007);
nand U25679 (N_25679,N_22597,N_23511);
nand U25680 (N_25680,N_20479,N_24821);
nand U25681 (N_25681,N_24264,N_23695);
or U25682 (N_25682,N_20370,N_24798);
or U25683 (N_25683,N_22401,N_20408);
nand U25684 (N_25684,N_23128,N_22186);
and U25685 (N_25685,N_21543,N_20883);
nand U25686 (N_25686,N_22940,N_22295);
nand U25687 (N_25687,N_22614,N_24826);
nand U25688 (N_25688,N_20684,N_20330);
nand U25689 (N_25689,N_23845,N_20540);
nand U25690 (N_25690,N_24399,N_24772);
xor U25691 (N_25691,N_24484,N_20848);
and U25692 (N_25692,N_21306,N_22790);
or U25693 (N_25693,N_20274,N_20569);
xor U25694 (N_25694,N_22497,N_21540);
nor U25695 (N_25695,N_20227,N_20271);
xor U25696 (N_25696,N_20850,N_23812);
or U25697 (N_25697,N_22683,N_23078);
or U25698 (N_25698,N_20057,N_20275);
nand U25699 (N_25699,N_20991,N_22787);
or U25700 (N_25700,N_24955,N_24638);
or U25701 (N_25701,N_23878,N_23173);
nor U25702 (N_25702,N_21261,N_22001);
nor U25703 (N_25703,N_22365,N_21083);
xnor U25704 (N_25704,N_20088,N_20695);
or U25705 (N_25705,N_20472,N_21427);
and U25706 (N_25706,N_24121,N_24462);
and U25707 (N_25707,N_20310,N_20301);
or U25708 (N_25708,N_24298,N_20113);
or U25709 (N_25709,N_23038,N_22185);
or U25710 (N_25710,N_20469,N_23213);
nand U25711 (N_25711,N_23182,N_21443);
and U25712 (N_25712,N_24984,N_21015);
and U25713 (N_25713,N_23563,N_20176);
xor U25714 (N_25714,N_23542,N_20689);
nand U25715 (N_25715,N_22595,N_20933);
or U25716 (N_25716,N_22502,N_22116);
nand U25717 (N_25717,N_21780,N_21622);
xnor U25718 (N_25718,N_23682,N_21798);
nor U25719 (N_25719,N_23747,N_20394);
nand U25720 (N_25720,N_20942,N_24213);
and U25721 (N_25721,N_24721,N_20930);
xor U25722 (N_25722,N_21101,N_23262);
and U25723 (N_25723,N_20065,N_20364);
and U25724 (N_25724,N_21795,N_20305);
or U25725 (N_25725,N_23207,N_23582);
or U25726 (N_25726,N_24735,N_21201);
nor U25727 (N_25727,N_23910,N_21182);
and U25728 (N_25728,N_23644,N_22530);
nor U25729 (N_25729,N_21572,N_20794);
nand U25730 (N_25730,N_21603,N_20112);
and U25731 (N_25731,N_23900,N_22207);
and U25732 (N_25732,N_21347,N_21692);
nand U25733 (N_25733,N_20626,N_20444);
nand U25734 (N_25734,N_22141,N_22489);
and U25735 (N_25735,N_22142,N_20884);
nor U25736 (N_25736,N_20278,N_23353);
nor U25737 (N_25737,N_24370,N_22391);
nor U25738 (N_25738,N_20140,N_23183);
and U25739 (N_25739,N_24616,N_24961);
nor U25740 (N_25740,N_20770,N_21783);
or U25741 (N_25741,N_24579,N_22122);
nand U25742 (N_25742,N_20367,N_24740);
and U25743 (N_25743,N_22992,N_24663);
nor U25744 (N_25744,N_20051,N_21985);
nand U25745 (N_25745,N_21130,N_24443);
and U25746 (N_25746,N_23579,N_23573);
nand U25747 (N_25747,N_22143,N_24986);
nor U25748 (N_25748,N_21929,N_22161);
nor U25749 (N_25749,N_23094,N_20431);
or U25750 (N_25750,N_24387,N_24540);
and U25751 (N_25751,N_20323,N_21847);
or U25752 (N_25752,N_23120,N_21447);
or U25753 (N_25753,N_24352,N_24104);
nand U25754 (N_25754,N_23715,N_20281);
xor U25755 (N_25755,N_24947,N_21338);
or U25756 (N_25756,N_23616,N_23711);
xnor U25757 (N_25757,N_22696,N_24890);
xor U25758 (N_25758,N_24539,N_23069);
and U25759 (N_25759,N_23430,N_24005);
and U25760 (N_25760,N_24464,N_21516);
nor U25761 (N_25761,N_23799,N_23121);
nand U25762 (N_25762,N_20234,N_21730);
nor U25763 (N_25763,N_22442,N_22260);
xor U25764 (N_25764,N_22452,N_23343);
xnor U25765 (N_25765,N_20858,N_20151);
and U25766 (N_25766,N_22841,N_20196);
xor U25767 (N_25767,N_23458,N_21548);
and U25768 (N_25768,N_23707,N_20640);
and U25769 (N_25769,N_24685,N_21858);
nor U25770 (N_25770,N_21367,N_23558);
nor U25771 (N_25771,N_20716,N_24169);
nand U25772 (N_25772,N_20002,N_21350);
or U25773 (N_25773,N_21557,N_20219);
and U25774 (N_25774,N_22220,N_20777);
nand U25775 (N_25775,N_20148,N_21869);
nand U25776 (N_25776,N_21146,N_21945);
xnor U25777 (N_25777,N_24910,N_24972);
nor U25778 (N_25778,N_22164,N_20875);
nor U25779 (N_25779,N_21849,N_24805);
nand U25780 (N_25780,N_24082,N_24734);
and U25781 (N_25781,N_23242,N_20917);
and U25782 (N_25782,N_23691,N_22396);
nor U25783 (N_25783,N_24642,N_21246);
nor U25784 (N_25784,N_23317,N_23348);
xor U25785 (N_25785,N_23926,N_20010);
xor U25786 (N_25786,N_21275,N_20035);
xor U25787 (N_25787,N_24021,N_22316);
nor U25788 (N_25788,N_20874,N_23283);
nor U25789 (N_25789,N_20913,N_22816);
nand U25790 (N_25790,N_22862,N_24554);
nor U25791 (N_25791,N_23625,N_21814);
and U25792 (N_25792,N_20069,N_22620);
nand U25793 (N_25793,N_24618,N_22511);
xnor U25794 (N_25794,N_22154,N_21322);
or U25795 (N_25795,N_21821,N_23260);
nand U25796 (N_25796,N_22102,N_23565);
xor U25797 (N_25797,N_24990,N_20907);
nand U25798 (N_25798,N_20356,N_24148);
nand U25799 (N_25799,N_22079,N_24146);
or U25800 (N_25800,N_20333,N_22446);
nand U25801 (N_25801,N_20753,N_23068);
or U25802 (N_25802,N_24704,N_20122);
nand U25803 (N_25803,N_23175,N_20986);
or U25804 (N_25804,N_20107,N_23226);
xor U25805 (N_25805,N_20786,N_20467);
or U25806 (N_25806,N_22545,N_24983);
nand U25807 (N_25807,N_23328,N_20337);
xor U25808 (N_25808,N_20524,N_21958);
or U25809 (N_25809,N_23275,N_21357);
nor U25810 (N_25810,N_21866,N_22826);
xnor U25811 (N_25811,N_21325,N_24305);
and U25812 (N_25812,N_20508,N_24584);
and U25813 (N_25813,N_24571,N_21992);
or U25814 (N_25814,N_20589,N_24688);
xnor U25815 (N_25815,N_21907,N_23622);
or U25816 (N_25816,N_24175,N_22735);
and U25817 (N_25817,N_24541,N_24522);
xnor U25818 (N_25818,N_22952,N_24846);
or U25819 (N_25819,N_20628,N_20984);
nor U25820 (N_25820,N_24952,N_23146);
xor U25821 (N_25821,N_21362,N_21212);
nor U25822 (N_25822,N_23603,N_24497);
xor U25823 (N_25823,N_21892,N_21252);
nor U25824 (N_25824,N_23324,N_24173);
nand U25825 (N_25825,N_21886,N_24436);
nor U25826 (N_25826,N_22152,N_20055);
nor U25827 (N_25827,N_23651,N_23980);
and U25828 (N_25828,N_20204,N_21941);
xnor U25829 (N_25829,N_22044,N_22402);
nor U25830 (N_25830,N_20655,N_21851);
nand U25831 (N_25831,N_23544,N_22985);
xor U25832 (N_25832,N_22307,N_20729);
nor U25833 (N_25833,N_22851,N_21076);
or U25834 (N_25834,N_23280,N_20049);
and U25835 (N_25835,N_23632,N_22411);
nand U25836 (N_25836,N_23237,N_23310);
nand U25837 (N_25837,N_24230,N_20650);
nor U25838 (N_25838,N_20321,N_20559);
and U25839 (N_25839,N_21431,N_20591);
nand U25840 (N_25840,N_23072,N_20355);
nand U25841 (N_25841,N_20373,N_21860);
nor U25842 (N_25842,N_23524,N_22856);
xor U25843 (N_25843,N_24084,N_21539);
or U25844 (N_25844,N_22894,N_20314);
nor U25845 (N_25845,N_22854,N_24065);
nand U25846 (N_25846,N_22598,N_21048);
xnor U25847 (N_25847,N_23654,N_24265);
nor U25848 (N_25848,N_22858,N_22909);
nor U25849 (N_25849,N_20816,N_21769);
nand U25850 (N_25850,N_22042,N_24167);
or U25851 (N_25851,N_23438,N_21052);
xnor U25852 (N_25852,N_24807,N_24677);
nand U25853 (N_25853,N_21118,N_21033);
or U25854 (N_25854,N_22993,N_24501);
xnor U25855 (N_25855,N_23451,N_20902);
and U25856 (N_25856,N_24747,N_22002);
xor U25857 (N_25857,N_21933,N_21660);
nor U25858 (N_25858,N_20395,N_23028);
or U25859 (N_25859,N_23110,N_20189);
nor U25860 (N_25860,N_23838,N_20514);
xor U25861 (N_25861,N_21245,N_22772);
and U25862 (N_25862,N_21641,N_24432);
xor U25863 (N_25863,N_22216,N_23304);
xor U25864 (N_25864,N_20941,N_22902);
nor U25865 (N_25865,N_23898,N_23000);
or U25866 (N_25866,N_22380,N_22349);
or U25867 (N_25867,N_21656,N_23151);
nand U25868 (N_25868,N_22139,N_22781);
or U25869 (N_25869,N_21837,N_23983);
or U25870 (N_25870,N_22225,N_21620);
and U25871 (N_25871,N_20504,N_21529);
nor U25872 (N_25872,N_23733,N_24322);
nand U25873 (N_25873,N_20247,N_22650);
and U25874 (N_25874,N_23091,N_22125);
nand U25875 (N_25875,N_20696,N_21400);
nand U25876 (N_25876,N_20087,N_20448);
nand U25877 (N_25877,N_22282,N_21764);
or U25878 (N_25878,N_22920,N_20357);
nand U25879 (N_25879,N_22232,N_24288);
or U25880 (N_25880,N_24067,N_21687);
or U25881 (N_25881,N_20017,N_21693);
xor U25882 (N_25882,N_21891,N_24249);
xor U25883 (N_25883,N_21166,N_21571);
and U25884 (N_25884,N_20658,N_23253);
xor U25885 (N_25885,N_22027,N_20239);
and U25886 (N_25886,N_22768,N_23863);
nor U25887 (N_25887,N_22407,N_23961);
or U25888 (N_25888,N_22445,N_24020);
nor U25889 (N_25889,N_22157,N_21208);
xnor U25890 (N_25890,N_24097,N_23176);
xnor U25891 (N_25891,N_22983,N_22806);
nand U25892 (N_25892,N_20297,N_23942);
nor U25893 (N_25893,N_24254,N_20732);
xnor U25894 (N_25894,N_20097,N_20177);
nor U25895 (N_25895,N_23663,N_24870);
xnor U25896 (N_25896,N_24128,N_23815);
or U25897 (N_25897,N_23525,N_22631);
nand U25898 (N_25898,N_20365,N_20060);
and U25899 (N_25899,N_23460,N_23537);
or U25900 (N_25900,N_24309,N_23093);
nand U25901 (N_25901,N_23391,N_21351);
or U25902 (N_25902,N_21137,N_21286);
and U25903 (N_25903,N_20186,N_24445);
xnor U25904 (N_25904,N_20259,N_20349);
or U25905 (N_25905,N_24601,N_22562);
xnor U25906 (N_25906,N_20474,N_24229);
xnor U25907 (N_25907,N_24475,N_24656);
xor U25908 (N_25908,N_22658,N_24487);
nor U25909 (N_25909,N_22274,N_20007);
and U25910 (N_25910,N_20997,N_20269);
nor U25911 (N_25911,N_22639,N_23669);
and U25912 (N_25912,N_20393,N_22106);
nand U25913 (N_25913,N_24582,N_20961);
nand U25914 (N_25914,N_23849,N_21398);
and U25915 (N_25915,N_20693,N_23675);
and U25916 (N_25916,N_24122,N_24017);
and U25917 (N_25917,N_23197,N_22648);
nand U25918 (N_25918,N_20090,N_24094);
nor U25919 (N_25919,N_23468,N_20632);
nand U25920 (N_25920,N_22022,N_23325);
nor U25921 (N_25921,N_23665,N_22054);
and U25922 (N_25922,N_22557,N_20012);
or U25923 (N_25923,N_20499,N_22350);
nor U25924 (N_25924,N_23697,N_22867);
xnor U25925 (N_25925,N_22262,N_22478);
or U25926 (N_25926,N_20919,N_23826);
nor U25927 (N_25927,N_22155,N_22180);
or U25928 (N_25928,N_20388,N_21957);
and U25929 (N_25929,N_21226,N_21290);
nor U25930 (N_25930,N_21506,N_20700);
nand U25931 (N_25931,N_23523,N_21108);
and U25932 (N_25932,N_21138,N_24194);
or U25933 (N_25933,N_21651,N_23916);
nand U25934 (N_25934,N_24938,N_24916);
and U25935 (N_25935,N_23408,N_23356);
nand U25936 (N_25936,N_23027,N_20983);
nor U25937 (N_25937,N_24615,N_20529);
nand U25938 (N_25938,N_21828,N_23819);
and U25939 (N_25939,N_24928,N_20243);
xnor U25940 (N_25940,N_24593,N_22681);
nand U25941 (N_25941,N_21964,N_21194);
and U25942 (N_25942,N_21039,N_22200);
nor U25943 (N_25943,N_21444,N_23409);
and U25944 (N_25944,N_24960,N_21637);
or U25945 (N_25945,N_20451,N_24205);
and U25946 (N_25946,N_20918,N_22641);
nand U25947 (N_25947,N_22127,N_20743);
and U25948 (N_25948,N_23658,N_20396);
or U25949 (N_25949,N_21590,N_23089);
and U25950 (N_25950,N_21342,N_20648);
xnor U25951 (N_25951,N_24055,N_24511);
or U25952 (N_25952,N_21976,N_21489);
nand U25953 (N_25953,N_23957,N_20267);
nand U25954 (N_25954,N_23567,N_20050);
and U25955 (N_25955,N_20675,N_24769);
nand U25956 (N_25956,N_24594,N_21983);
nand U25957 (N_25957,N_21711,N_21009);
and U25958 (N_25958,N_20464,N_20296);
xnor U25959 (N_25959,N_21614,N_24371);
nor U25960 (N_25960,N_24042,N_21748);
or U25961 (N_25961,N_22524,N_22812);
nand U25962 (N_25962,N_23583,N_20096);
nor U25963 (N_25963,N_21259,N_22153);
nor U25964 (N_25964,N_20276,N_21116);
and U25965 (N_25965,N_21501,N_21953);
nor U25966 (N_25966,N_24183,N_20125);
or U25967 (N_25967,N_24061,N_24068);
xnor U25968 (N_25968,N_23061,N_22397);
nand U25969 (N_25969,N_22712,N_22317);
and U25970 (N_25970,N_21733,N_21060);
or U25971 (N_25971,N_24054,N_24773);
nand U25972 (N_25972,N_21610,N_22528);
or U25973 (N_25973,N_21179,N_22490);
nor U25974 (N_25974,N_24237,N_21629);
or U25975 (N_25975,N_24050,N_22231);
nor U25976 (N_25976,N_20549,N_24359);
xor U25977 (N_25977,N_22259,N_24998);
nand U25978 (N_25978,N_22005,N_20889);
xnor U25979 (N_25979,N_22752,N_22438);
nor U25980 (N_25980,N_21565,N_24530);
and U25981 (N_25981,N_21242,N_22038);
xor U25982 (N_25982,N_24548,N_21535);
and U25983 (N_25983,N_23232,N_23688);
xnor U25984 (N_25984,N_20975,N_23160);
nand U25985 (N_25985,N_21934,N_23976);
or U25986 (N_25986,N_24232,N_24178);
nand U25987 (N_25987,N_23506,N_23349);
and U25988 (N_25988,N_20465,N_21530);
or U25989 (N_25989,N_21062,N_24877);
xnor U25990 (N_25990,N_23208,N_24531);
nand U25991 (N_25991,N_20014,N_22064);
nand U25992 (N_25992,N_23054,N_23113);
nand U25993 (N_25993,N_24338,N_24514);
nand U25994 (N_25994,N_21667,N_20073);
nor U25995 (N_25995,N_21043,N_24323);
or U25996 (N_25996,N_23720,N_24504);
and U25997 (N_25997,N_23233,N_22802);
or U25998 (N_25998,N_24092,N_23399);
and U25999 (N_25999,N_24095,N_21547);
and U26000 (N_26000,N_24959,N_20506);
and U26001 (N_26001,N_22990,N_23082);
nand U26002 (N_26002,N_22088,N_22886);
xnor U26003 (N_26003,N_23966,N_21727);
xor U26004 (N_26004,N_20218,N_22888);
nand U26005 (N_26005,N_20351,N_24049);
nand U26006 (N_26006,N_20132,N_24670);
and U26007 (N_26007,N_23425,N_22014);
and U26008 (N_26008,N_22523,N_24796);
or U26009 (N_26009,N_22400,N_23046);
or U26010 (N_26010,N_23962,N_23472);
nor U26011 (N_26011,N_22195,N_24449);
or U26012 (N_26012,N_20947,N_22974);
xnor U26013 (N_26013,N_23556,N_21228);
or U26014 (N_26014,N_23852,N_21209);
and U26015 (N_26015,N_20717,N_21231);
and U26016 (N_26016,N_21148,N_23462);
nor U26017 (N_26017,N_23498,N_20576);
xor U26018 (N_26018,N_23555,N_24335);
and U26019 (N_26019,N_24657,N_23052);
and U26020 (N_26020,N_22028,N_24898);
nor U26021 (N_26021,N_23722,N_22386);
xor U26022 (N_26022,N_24001,N_21644);
nor U26023 (N_26023,N_24715,N_22963);
xor U26024 (N_26024,N_20480,N_22516);
xor U26025 (N_26025,N_23714,N_24300);
or U26026 (N_26026,N_21170,N_21591);
nand U26027 (N_26027,N_20103,N_22335);
nor U26028 (N_26028,N_21844,N_24674);
nor U26029 (N_26029,N_24027,N_24386);
nand U26030 (N_26030,N_22499,N_21025);
nand U26031 (N_26031,N_21063,N_23437);
xnor U26032 (N_26032,N_20572,N_22691);
or U26033 (N_26033,N_20324,N_24078);
nand U26034 (N_26034,N_20449,N_23519);
and U26035 (N_26035,N_22450,N_22758);
xor U26036 (N_26036,N_22750,N_24869);
xnor U26037 (N_26037,N_21031,N_24109);
xnor U26038 (N_26038,N_23535,N_21073);
nand U26039 (N_26039,N_23227,N_22434);
nor U26040 (N_26040,N_24703,N_21434);
and U26041 (N_26041,N_22017,N_21375);
and U26042 (N_26042,N_22246,N_24623);
xnor U26043 (N_26043,N_24978,N_22366);
nor U26044 (N_26044,N_20905,N_20153);
nand U26045 (N_26045,N_23598,N_23382);
nand U26046 (N_26046,N_21811,N_22192);
nor U26047 (N_26047,N_21659,N_24914);
nand U26048 (N_26048,N_23102,N_24369);
xor U26049 (N_26049,N_21316,N_23678);
nor U26050 (N_26050,N_21735,N_22052);
and U26051 (N_26051,N_22688,N_22206);
nand U26052 (N_26052,N_20207,N_24502);
and U26053 (N_26053,N_20855,N_23142);
nor U26054 (N_26054,N_24204,N_23835);
or U26055 (N_26055,N_21408,N_22212);
and U26056 (N_26056,N_24170,N_22744);
and U26057 (N_26057,N_20172,N_21908);
nor U26058 (N_26058,N_22615,N_21593);
nor U26059 (N_26059,N_21643,N_24479);
nand U26060 (N_26060,N_20630,N_23158);
nand U26061 (N_26061,N_24630,N_20826);
xor U26062 (N_26062,N_20535,N_23709);
nor U26063 (N_26063,N_23584,N_23694);
xnor U26064 (N_26064,N_20517,N_21581);
and U26065 (N_26065,N_21197,N_21497);
xor U26066 (N_26066,N_23254,N_21495);
nand U26067 (N_26067,N_20706,N_23471);
and U26068 (N_26068,N_20455,N_23235);
or U26069 (N_26069,N_21607,N_24786);
xor U26070 (N_26070,N_20820,N_24976);
nor U26071 (N_26071,N_23597,N_21720);
and U26072 (N_26072,N_20721,N_22773);
xor U26073 (N_26073,N_22514,N_22905);
or U26074 (N_26074,N_21753,N_20163);
and U26075 (N_26075,N_24560,N_22012);
or U26076 (N_26076,N_20888,N_21103);
and U26077 (N_26077,N_22532,N_20402);
xor U26078 (N_26078,N_21790,N_24467);
nand U26079 (N_26079,N_22961,N_20498);
xnor U26080 (N_26080,N_22368,N_24975);
nor U26081 (N_26081,N_23440,N_23131);
nand U26082 (N_26082,N_21688,N_24418);
xnor U26083 (N_26083,N_20651,N_20450);
and U26084 (N_26084,N_22387,N_20595);
nand U26085 (N_26085,N_21685,N_22472);
nor U26086 (N_26086,N_24023,N_21781);
nand U26087 (N_26087,N_24317,N_21949);
and U26088 (N_26088,N_22680,N_24850);
nand U26089 (N_26089,N_22609,N_23893);
or U26090 (N_26090,N_22942,N_21632);
xor U26091 (N_26091,N_20783,N_22226);
and U26092 (N_26092,N_21683,N_21754);
xnor U26093 (N_26093,N_23879,N_24882);
nor U26094 (N_26094,N_21332,N_24334);
nor U26095 (N_26095,N_22721,N_22633);
xor U26096 (N_26096,N_20856,N_22483);
nor U26097 (N_26097,N_24454,N_23411);
xnor U26098 (N_26098,N_22252,N_21152);
nor U26099 (N_26099,N_23534,N_20563);
xor U26100 (N_26100,N_20646,N_22243);
xnor U26101 (N_26101,N_22361,N_23971);
nor U26102 (N_26102,N_22359,N_23323);
nand U26103 (N_26103,N_24329,N_22063);
nand U26104 (N_26104,N_21215,N_23240);
nand U26105 (N_26105,N_23350,N_24051);
xnor U26106 (N_26106,N_20725,N_21345);
xor U26107 (N_26107,N_20198,N_22265);
or U26108 (N_26108,N_20494,N_21294);
nand U26109 (N_26109,N_24326,N_23342);
nand U26110 (N_26110,N_24200,N_23303);
and U26111 (N_26111,N_24761,N_24619);
or U26112 (N_26112,N_23103,N_20592);
nor U26113 (N_26113,N_24851,N_21084);
nand U26114 (N_26114,N_23801,N_20945);
xor U26115 (N_26115,N_22358,N_22276);
xnor U26116 (N_26116,N_24728,N_21472);
and U26117 (N_26117,N_23172,N_21486);
nor U26118 (N_26118,N_22469,N_20915);
or U26119 (N_26119,N_22078,N_20629);
or U26120 (N_26120,N_24799,N_22644);
nor U26121 (N_26121,N_20048,N_21503);
nor U26122 (N_26122,N_22995,N_20992);
nor U26123 (N_26123,N_23385,N_21283);
xor U26124 (N_26124,N_21423,N_23418);
and U26125 (N_26125,N_20560,N_20268);
nor U26126 (N_26126,N_23494,N_23180);
and U26127 (N_26127,N_22278,N_20000);
xor U26128 (N_26128,N_21476,N_22374);
xnor U26129 (N_26129,N_20552,N_21774);
nand U26130 (N_26130,N_22788,N_23734);
xnor U26131 (N_26131,N_24337,N_20139);
xnor U26132 (N_26132,N_20749,N_22774);
and U26133 (N_26133,N_22543,N_20722);
and U26134 (N_26134,N_23025,N_21119);
xor U26135 (N_26135,N_22412,N_21485);
nor U26136 (N_26136,N_22264,N_24622);
nor U26137 (N_26137,N_22941,N_23050);
or U26138 (N_26138,N_24160,N_20834);
nor U26139 (N_26139,N_24491,N_23329);
and U26140 (N_26140,N_23306,N_23037);
xor U26141 (N_26141,N_20120,N_23868);
and U26142 (N_26142,N_23267,N_20619);
xnor U26143 (N_26143,N_24280,N_24995);
xor U26144 (N_26144,N_20944,N_22118);
xor U26145 (N_26145,N_20644,N_22928);
xnor U26146 (N_26146,N_22656,N_24367);
xnor U26147 (N_26147,N_24490,N_24752);
nor U26148 (N_26148,N_23602,N_24770);
or U26149 (N_26149,N_24564,N_24736);
nor U26150 (N_26150,N_22284,N_24188);
nor U26151 (N_26151,N_20709,N_24417);
or U26152 (N_26152,N_23522,N_24523);
or U26153 (N_26153,N_24563,N_21952);
xor U26154 (N_26154,N_21405,N_24699);
or U26155 (N_26155,N_21300,N_20292);
nand U26156 (N_26156,N_23111,N_20253);
or U26157 (N_26157,N_24262,N_21214);
and U26158 (N_26158,N_24327,N_23489);
nand U26159 (N_26159,N_21729,N_22537);
nand U26160 (N_26160,N_21960,N_21864);
xor U26161 (N_26161,N_21418,N_24276);
and U26162 (N_26162,N_24926,N_24754);
and U26163 (N_26163,N_22776,N_21059);
or U26164 (N_26164,N_20765,N_24398);
nor U26165 (N_26165,N_21373,N_22887);
nand U26166 (N_26166,N_21738,N_20811);
or U26167 (N_26167,N_22100,N_21389);
nor U26168 (N_26168,N_21305,N_24659);
or U26169 (N_26169,N_20077,N_22439);
and U26170 (N_26170,N_20704,N_20868);
or U26171 (N_26171,N_24620,N_24576);
nor U26172 (N_26172,N_21538,N_20042);
or U26173 (N_26173,N_20249,N_24219);
and U26174 (N_26174,N_24318,N_24631);
nor U26175 (N_26175,N_24783,N_21149);
xor U26176 (N_26176,N_20428,N_23203);
and U26177 (N_26177,N_20577,N_20427);
or U26178 (N_26178,N_23104,N_21441);
nand U26179 (N_26179,N_21956,N_21881);
nor U26180 (N_26180,N_20877,N_24830);
or U26181 (N_26181,N_20208,N_21352);
xnor U26182 (N_26182,N_21853,N_20460);
and U26183 (N_26183,N_20375,N_22568);
and U26184 (N_26184,N_24580,N_21863);
nand U26185 (N_26185,N_20526,N_21205);
or U26186 (N_26186,N_24855,N_23003);
nor U26187 (N_26187,N_24103,N_20539);
xnor U26188 (N_26188,N_23604,N_23770);
nand U26189 (N_26189,N_22103,N_21178);
xnor U26190 (N_26190,N_21317,N_24922);
nand U26191 (N_26191,N_20680,N_20843);
or U26192 (N_26192,N_23772,N_22578);
or U26193 (N_26193,N_22913,N_22441);
nand U26194 (N_26194,N_22755,N_21582);
xor U26195 (N_26195,N_20870,N_20313);
and U26196 (N_26196,N_21872,N_21696);
nor U26197 (N_26197,N_21520,N_20756);
or U26198 (N_26198,N_22159,N_23147);
nand U26199 (N_26199,N_24321,N_23381);
nor U26200 (N_26200,N_24143,N_21613);
and U26201 (N_26201,N_22071,N_20830);
or U26202 (N_26202,N_20462,N_20216);
nand U26203 (N_26203,N_20719,N_21878);
and U26204 (N_26204,N_20345,N_20768);
nand U26205 (N_26205,N_20897,N_20673);
nor U26206 (N_26206,N_21018,N_21758);
nor U26207 (N_26207,N_20582,N_23829);
and U26208 (N_26208,N_24701,N_24544);
nand U26209 (N_26209,N_20891,N_23365);
or U26210 (N_26210,N_22795,N_21089);
nand U26211 (N_26211,N_20972,N_20946);
nand U26212 (N_26212,N_24858,N_24350);
and U26213 (N_26213,N_21433,N_20085);
or U26214 (N_26214,N_22797,N_22081);
and U26215 (N_26215,N_22554,N_21136);
nor U26216 (N_26216,N_23899,N_23289);
and U26217 (N_26217,N_22319,N_20461);
and U26218 (N_26218,N_22251,N_20114);
and U26219 (N_26219,N_24233,N_22055);
xnor U26220 (N_26220,N_22224,N_24671);
or U26221 (N_26221,N_21585,N_24004);
or U26222 (N_26222,N_22098,N_23854);
and U26223 (N_26223,N_21676,N_20423);
nand U26224 (N_26224,N_21303,N_23920);
nor U26225 (N_26225,N_24888,N_22586);
xnor U26226 (N_26226,N_24073,N_24405);
xnor U26227 (N_26227,N_23459,N_24201);
xnor U26228 (N_26228,N_23641,N_24347);
xnor U26229 (N_26229,N_21289,N_24817);
nand U26230 (N_26230,N_21873,N_24325);
or U26231 (N_26231,N_22931,N_21339);
nand U26232 (N_26232,N_24114,N_21172);
xor U26233 (N_26233,N_24277,N_24293);
nor U26234 (N_26234,N_22807,N_20805);
nor U26235 (N_26235,N_20419,N_22059);
xor U26236 (N_26236,N_21761,N_22035);
nor U26237 (N_26237,N_20657,N_21445);
xnor U26238 (N_26238,N_20266,N_23206);
and U26239 (N_26239,N_24444,N_21195);
and U26240 (N_26240,N_20129,N_23398);
nand U26241 (N_26241,N_21448,N_22793);
nand U26242 (N_26242,N_24015,N_24900);
and U26243 (N_26243,N_22546,N_21879);
or U26244 (N_26244,N_21395,N_21704);
nand U26245 (N_26245,N_21202,N_20166);
or U26246 (N_26246,N_20607,N_23373);
and U26247 (N_26247,N_21598,N_24151);
nand U26248 (N_26248,N_24781,N_23488);
nor U26249 (N_26249,N_20744,N_21093);
nand U26250 (N_26250,N_20159,N_23726);
and U26251 (N_26251,N_21233,N_21238);
xor U26252 (N_26252,N_23886,N_20344);
and U26253 (N_26253,N_24906,N_23703);
nor U26254 (N_26254,N_23670,N_20994);
nor U26255 (N_26255,N_24871,N_23901);
nor U26256 (N_26256,N_24287,N_20053);
or U26257 (N_26257,N_20521,N_22181);
xor U26258 (N_26258,N_23725,N_24434);
or U26259 (N_26259,N_23366,N_24294);
or U26260 (N_26260,N_22091,N_22789);
and U26261 (N_26261,N_23017,N_21831);
xnor U26262 (N_26262,N_22147,N_21185);
nand U26263 (N_26263,N_23338,N_22242);
and U26264 (N_26264,N_22146,N_21680);
or U26265 (N_26265,N_24022,N_21006);
xnor U26266 (N_26266,N_21736,N_22962);
nand U26267 (N_26267,N_24738,N_20568);
nor U26268 (N_26268,N_20354,N_20433);
xor U26269 (N_26269,N_24171,N_21766);
or U26270 (N_26270,N_21278,N_23706);
nor U26271 (N_26271,N_21134,N_21301);
or U26272 (N_26272,N_23517,N_24353);
or U26273 (N_26273,N_20182,N_24894);
or U26274 (N_26274,N_22447,N_23010);
and U26275 (N_26275,N_21940,N_24839);
or U26276 (N_26276,N_23423,N_23127);
and U26277 (N_26277,N_22891,N_22625);
nand U26278 (N_26278,N_23291,N_23927);
and U26279 (N_26279,N_24942,N_22476);
and U26280 (N_26280,N_24834,N_24319);
or U26281 (N_26281,N_20951,N_21900);
xnor U26282 (N_26282,N_22628,N_24380);
or U26283 (N_26283,N_22784,N_22318);
nor U26284 (N_26284,N_23287,N_22695);
xor U26285 (N_26285,N_20338,N_20823);
nand U26286 (N_26286,N_23134,N_24313);
nor U26287 (N_26287,N_22878,N_24115);
or U26288 (N_26288,N_22462,N_24483);
nand U26289 (N_26289,N_24779,N_20963);
nor U26290 (N_26290,N_24072,N_21716);
or U26291 (N_26291,N_22239,N_20286);
nand U26292 (N_26292,N_22105,N_24534);
xnor U26293 (N_26293,N_20210,N_24681);
xor U26294 (N_26294,N_22166,N_22604);
and U26295 (N_26295,N_21705,N_22838);
xor U26296 (N_26296,N_21022,N_23475);
nand U26297 (N_26297,N_22771,N_20964);
nand U26298 (N_26298,N_21902,N_20798);
nor U26299 (N_26299,N_22113,N_21295);
xnor U26300 (N_26300,N_20741,N_24473);
nor U26301 (N_26301,N_22693,N_20898);
nand U26302 (N_26302,N_20735,N_24886);
nor U26303 (N_26303,N_23002,N_21655);
xnor U26304 (N_26304,N_22433,N_22892);
nand U26305 (N_26305,N_22487,N_22204);
and U26306 (N_26306,N_23737,N_22704);
xor U26307 (N_26307,N_22709,N_23952);
or U26308 (N_26308,N_22972,N_20860);
and U26309 (N_26309,N_20702,N_21982);
nand U26310 (N_26310,N_22997,N_20604);
and U26311 (N_26311,N_20072,N_20493);
nand U26312 (N_26312,N_21650,N_23390);
or U26313 (N_26313,N_20791,N_24720);
or U26314 (N_26314,N_20115,N_24635);
nand U26315 (N_26315,N_21836,N_20575);
and U26316 (N_26316,N_22746,N_24713);
xnor U26317 (N_26317,N_23946,N_23635);
nand U26318 (N_26318,N_24310,N_23413);
xor U26319 (N_26319,N_22782,N_22424);
and U26320 (N_26320,N_22549,N_24920);
and U26321 (N_26321,N_20298,N_22967);
or U26322 (N_26322,N_21935,N_24066);
nand U26323 (N_26323,N_24950,N_24155);
and U26324 (N_26324,N_21335,N_23761);
nand U26325 (N_26325,N_22921,N_21987);
and U26326 (N_26326,N_23018,N_22764);
nand U26327 (N_26327,N_22881,N_21371);
and U26328 (N_26328,N_23049,N_23653);
nand U26329 (N_26329,N_22369,N_20380);
and U26330 (N_26330,N_22432,N_20383);
nor U26331 (N_26331,N_20760,N_21586);
or U26332 (N_26332,N_23881,N_23967);
nor U26333 (N_26333,N_22461,N_24964);
nand U26334 (N_26334,N_20956,N_21682);
xnor U26335 (N_26335,N_24057,N_22872);
and U26336 (N_26336,N_21309,N_24924);
nand U26337 (N_26337,N_24838,N_22813);
xnor U26338 (N_26338,N_23546,N_20739);
and U26339 (N_26339,N_21714,N_21745);
or U26340 (N_26340,N_22564,N_20184);
nor U26341 (N_26341,N_24891,N_24958);
nand U26342 (N_26342,N_24433,N_24279);
nor U26343 (N_26343,N_23322,N_24149);
nand U26344 (N_26344,N_24967,N_24979);
xnor U26345 (N_26345,N_20127,N_21587);
or U26346 (N_26346,N_22596,N_21896);
nand U26347 (N_26347,N_20773,N_20879);
nor U26348 (N_26348,N_21380,N_20341);
nor U26349 (N_26349,N_24246,N_23624);
nand U26350 (N_26350,N_22907,N_20260);
xor U26351 (N_26351,N_24009,N_24507);
or U26352 (N_26352,N_20492,N_23257);
nor U26353 (N_26353,N_22729,N_21032);
xnor U26354 (N_26354,N_22763,N_24724);
xor U26355 (N_26355,N_20774,N_20076);
nor U26356 (N_26356,N_22352,N_21040);
or U26357 (N_26357,N_21806,N_21065);
or U26358 (N_26358,N_23467,N_20133);
or U26359 (N_26359,N_23575,N_22667);
nand U26360 (N_26360,N_23154,N_22757);
xor U26361 (N_26361,N_21435,N_22778);
or U26362 (N_26362,N_24166,N_22070);
and U26363 (N_26363,N_22770,N_20359);
nand U26364 (N_26364,N_22477,N_22210);
and U26365 (N_26365,N_24946,N_24755);
nand U26366 (N_26366,N_23251,N_24912);
nor U26367 (N_26367,N_23397,N_21211);
nor U26368 (N_26368,N_23473,N_21800);
xnor U26369 (N_26369,N_24517,N_21457);
nor U26370 (N_26370,N_22370,N_24581);
and U26371 (N_26371,N_21959,N_22747);
xnor U26372 (N_26372,N_22272,N_21663);
nand U26373 (N_26373,N_22986,N_21490);
nor U26374 (N_26374,N_22724,N_20846);
and U26375 (N_26375,N_23585,N_24840);
xnor U26376 (N_26376,N_24566,N_23606);
nor U26377 (N_26377,N_21628,N_21595);
or U26378 (N_26378,N_24719,N_23997);
nand U26379 (N_26379,N_24281,N_24803);
nor U26380 (N_26380,N_22156,N_23830);
xnor U26381 (N_26381,N_22533,N_22925);
nand U26382 (N_26382,N_24002,N_22377);
xor U26383 (N_26383,N_21471,N_24757);
xnor U26384 (N_26384,N_22883,N_21219);
xor U26385 (N_26385,N_22550,N_22538);
nor U26386 (N_26386,N_23097,N_22169);
nor U26387 (N_26387,N_23569,N_21247);
xor U26388 (N_26388,N_20662,N_20736);
nand U26389 (N_26389,N_21267,N_24827);
nand U26390 (N_26390,N_21041,N_20348);
or U26391 (N_26391,N_22191,N_24759);
nand U26392 (N_26392,N_23185,N_21177);
nor U26393 (N_26393,N_21248,N_24157);
xor U26394 (N_26394,N_24162,N_21523);
and U26395 (N_26395,N_22669,N_23786);
xnor U26396 (N_26396,N_20893,N_24692);
or U26397 (N_26397,N_21449,N_22873);
nand U26398 (N_26398,N_20174,N_20894);
nor U26399 (N_26399,N_22531,N_20162);
xor U26400 (N_26400,N_22202,N_20441);
and U26401 (N_26401,N_24815,N_23674);
or U26402 (N_26402,N_21797,N_24492);
or U26403 (N_26403,N_22334,N_20242);
and U26404 (N_26404,N_21947,N_22701);
xor U26405 (N_26405,N_23490,N_23292);
xor U26406 (N_26406,N_23611,N_20606);
or U26407 (N_26407,N_24468,N_22589);
xnor U26408 (N_26408,N_23724,N_21122);
xor U26409 (N_26409,N_20812,N_22703);
nor U26410 (N_26410,N_21096,N_23201);
or U26411 (N_26411,N_20043,N_21903);
and U26412 (N_26412,N_21533,N_20202);
and U26413 (N_26413,N_24282,N_20263);
nand U26414 (N_26414,N_22606,N_21817);
nor U26415 (N_26415,N_20272,N_22149);
xor U26416 (N_26416,N_23118,N_22948);
nor U26417 (N_26417,N_23264,N_22394);
nand U26418 (N_26418,N_24965,N_20376);
nor U26419 (N_26419,N_22692,N_23354);
xor U26420 (N_26420,N_22214,N_21131);
nand U26421 (N_26421,N_22114,N_20192);
xnor U26422 (N_26422,N_22792,N_21458);
xor U26423 (N_26423,N_24857,N_21075);
xor U26424 (N_26424,N_20603,N_23023);
or U26425 (N_26425,N_20726,N_23666);
or U26426 (N_26426,N_20258,N_22040);
and U26427 (N_26427,N_21480,N_23719);
nand U26428 (N_26428,N_23402,N_22512);
nor U26429 (N_26429,N_21580,N_24726);
nand U26430 (N_26430,N_24935,N_23728);
nor U26431 (N_26431,N_24525,N_21657);
nor U26432 (N_26432,N_24192,N_23499);
nor U26433 (N_26433,N_23862,N_20542);
and U26434 (N_26434,N_23022,N_21726);
nor U26435 (N_26435,N_24190,N_24519);
or U26436 (N_26436,N_21262,N_22313);
and U26437 (N_26437,N_24260,N_21154);
and U26438 (N_26438,N_23501,N_22431);
or U26439 (N_26439,N_20476,N_20573);
nand U26440 (N_26440,N_21997,N_22610);
nor U26441 (N_26441,N_24945,N_23070);
and U26442 (N_26442,N_20788,N_21364);
nor U26443 (N_26443,N_21478,N_24010);
or U26444 (N_26444,N_23090,N_21493);
xor U26445 (N_26445,N_20608,N_20962);
nand U26446 (N_26446,N_23895,N_22585);
or U26447 (N_26447,N_23006,N_20034);
nand U26448 (N_26448,N_24059,N_23076);
nor U26449 (N_26449,N_22448,N_23272);
and U26450 (N_26450,N_24604,N_24003);
nand U26451 (N_26451,N_20600,N_22825);
or U26452 (N_26452,N_21928,N_23186);
nand U26453 (N_26453,N_24646,N_21584);
and U26454 (N_26454,N_20178,N_21024);
xnor U26455 (N_26455,N_20597,N_21901);
and U26456 (N_26456,N_23743,N_23219);
or U26457 (N_26457,N_22031,N_23223);
nand U26458 (N_26458,N_22051,N_23739);
nand U26459 (N_26459,N_24546,N_23435);
nand U26460 (N_26460,N_21601,N_22885);
and U26461 (N_26461,N_21193,N_21225);
and U26462 (N_26462,N_21237,N_21799);
nor U26463 (N_26463,N_23664,N_23339);
and U26464 (N_26464,N_22020,N_22072);
or U26465 (N_26465,N_23231,N_23580);
or U26466 (N_26466,N_21068,N_24968);
nor U26467 (N_26467,N_21662,N_22527);
xnor U26468 (N_26468,N_21452,N_24411);
or U26469 (N_26469,N_21808,N_23984);
or U26470 (N_26470,N_20106,N_22183);
nor U26471 (N_26471,N_22900,N_23564);
or U26472 (N_26472,N_23992,N_20343);
and U26473 (N_26473,N_22869,N_24426);
or U26474 (N_26474,N_23700,N_21199);
nand U26475 (N_26475,N_22293,N_24767);
and U26476 (N_26476,N_23153,N_24941);
xor U26477 (N_26477,N_24421,N_21167);
nand U26478 (N_26478,N_23318,N_21526);
nor U26479 (N_26479,N_20205,N_21624);
or U26480 (N_26480,N_22346,N_23738);
or U26481 (N_26481,N_23936,N_20955);
xnor U26482 (N_26482,N_23268,N_20715);
xnor U26483 (N_26483,N_20759,N_23300);
nand U26484 (N_26484,N_21085,N_21794);
nand U26485 (N_26485,N_20769,N_20800);
or U26486 (N_26486,N_24668,N_21318);
or U26487 (N_26487,N_24382,N_21120);
and U26488 (N_26488,N_24236,N_21164);
nand U26489 (N_26489,N_24482,N_21200);
nor U26490 (N_26490,N_24841,N_23750);
and U26491 (N_26491,N_21026,N_20967);
xor U26492 (N_26492,N_20789,N_21567);
nor U26493 (N_26493,N_23672,N_22341);
or U26494 (N_26494,N_20256,N_22364);
or U26495 (N_26495,N_22281,N_23290);
nor U26496 (N_26496,N_22026,N_24923);
or U26497 (N_26497,N_24746,N_23631);
or U26498 (N_26498,N_20156,N_20056);
or U26499 (N_26499,N_21918,N_22008);
nand U26500 (N_26500,N_21517,N_22049);
nor U26501 (N_26501,N_21360,N_24041);
and U26502 (N_26502,N_24809,N_22844);
or U26503 (N_26503,N_20639,N_24810);
nand U26504 (N_26504,N_22848,N_20511);
and U26505 (N_26505,N_21487,N_23463);
nor U26506 (N_26506,N_24574,N_22240);
and U26507 (N_26507,N_24503,N_24110);
xor U26508 (N_26508,N_22859,N_23278);
nor U26509 (N_26509,N_22668,N_22215);
nand U26510 (N_26510,N_21792,N_20164);
and U26511 (N_26511,N_24248,N_23196);
nand U26512 (N_26512,N_20287,N_21880);
nand U26513 (N_26513,N_22988,N_24156);
and U26514 (N_26514,N_20674,N_21319);
nand U26515 (N_26515,N_24011,N_24476);
and U26516 (N_26516,N_20322,N_22238);
nand U26517 (N_26517,N_24106,N_21668);
and U26518 (N_26518,N_20723,N_22630);
nor U26519 (N_26519,N_20547,N_21975);
nor U26520 (N_26520,N_24238,N_23657);
nand U26521 (N_26521,N_22289,N_24818);
and U26522 (N_26522,N_22291,N_24705);
or U26523 (N_26523,N_21081,N_23784);
nand U26524 (N_26524,N_24575,N_20565);
nor U26525 (N_26525,N_24258,N_22895);
and U26526 (N_26526,N_23406,N_22255);
and U26527 (N_26527,N_23100,N_23540);
or U26528 (N_26528,N_22824,N_24026);
or U26529 (N_26529,N_20013,N_23935);
xnor U26530 (N_26530,N_22743,N_20625);
nor U26531 (N_26531,N_20996,N_20264);
nand U26532 (N_26532,N_21333,N_24342);
xor U26533 (N_26533,N_23753,N_21329);
or U26534 (N_26534,N_21374,N_22559);
nand U26535 (N_26535,N_24466,N_24697);
and U26536 (N_26536,N_23742,N_22097);
nand U26537 (N_26537,N_20410,N_22254);
nor U26538 (N_26538,N_22305,N_20821);
and U26539 (N_26539,N_24416,N_20971);
or U26540 (N_26540,N_24603,N_23432);
xor U26541 (N_26541,N_21791,N_23846);
nand U26542 (N_26542,N_24240,N_24811);
or U26543 (N_26543,N_23297,N_22248);
nor U26544 (N_26544,N_22333,N_24732);
nor U26545 (N_26545,N_23214,N_23130);
nor U26546 (N_26546,N_21327,N_21528);
and U26547 (N_26547,N_22908,N_20643);
nor U26548 (N_26548,N_20537,N_24437);
nor U26549 (N_26549,N_24186,N_20714);
or U26550 (N_26550,N_20121,N_23062);
and U26551 (N_26551,N_22876,N_20922);
nor U26552 (N_26552,N_20197,N_21707);
nor U26553 (N_26553,N_23836,N_21756);
or U26554 (N_26554,N_24634,N_23320);
and U26555 (N_26555,N_21411,N_23170);
or U26556 (N_26556,N_21308,N_23824);
or U26557 (N_26557,N_21859,N_20799);
or U26558 (N_26558,N_20982,N_22036);
and U26559 (N_26559,N_20581,N_24862);
nand U26560 (N_26560,N_20421,N_22473);
or U26561 (N_26561,N_24884,N_20160);
nor U26562 (N_26562,N_21401,N_21187);
or U26563 (N_26563,N_22552,N_22687);
xnor U26564 (N_26564,N_24929,N_23646);
nor U26565 (N_26565,N_23526,N_24159);
or U26566 (N_26566,N_22932,N_20627);
or U26567 (N_26567,N_20400,N_20681);
and U26568 (N_26568,N_20676,N_20191);
nand U26569 (N_26569,N_22228,N_21995);
xnor U26570 (N_26570,N_22222,N_24090);
nor U26571 (N_26571,N_21965,N_24774);
nor U26572 (N_26572,N_24516,N_21980);
or U26573 (N_26573,N_21402,N_21690);
and U26574 (N_26574,N_23302,N_24225);
and U26575 (N_26575,N_24422,N_21749);
xnor U26576 (N_26576,N_22444,N_23099);
xnor U26577 (N_26577,N_20633,N_24836);
nand U26578 (N_26578,N_24897,N_21206);
nand U26579 (N_26579,N_24653,N_21905);
nor U26580 (N_26580,N_21363,N_23171);
or U26581 (N_26581,N_23757,N_24764);
and U26582 (N_26582,N_21512,N_23042);
nand U26583 (N_26583,N_22762,N_22663);
or U26584 (N_26584,N_22973,N_24435);
nor U26585 (N_26585,N_20358,N_20318);
xnor U26586 (N_26586,N_21064,N_24331);
or U26587 (N_26587,N_23764,N_20841);
xor U26588 (N_26588,N_20712,N_20624);
or U26589 (N_26589,N_24533,N_24270);
nor U26590 (N_26590,N_22076,N_20407);
or U26591 (N_26591,N_22420,N_21948);
nand U26592 (N_26592,N_24187,N_23749);
nand U26593 (N_26593,N_21235,N_22312);
and U26594 (N_26594,N_21626,N_22011);
and U26595 (N_26595,N_21276,N_22507);
or U26596 (N_26596,N_24934,N_22818);
nand U26597 (N_26597,N_20852,N_24528);
or U26598 (N_26598,N_23448,N_23857);
nor U26599 (N_26599,N_22384,N_20316);
and U26600 (N_26600,N_23660,N_22301);
nand U26601 (N_26601,N_20672,N_20233);
nor U26602 (N_26602,N_24123,N_21424);
nor U26603 (N_26603,N_24992,N_22565);
nand U26604 (N_26604,N_22728,N_21911);
nand U26605 (N_26605,N_20869,N_21967);
nand U26606 (N_26606,N_23648,N_21314);
and U26607 (N_26607,N_23202,N_22117);
nand U26608 (N_26608,N_22964,N_20806);
xor U26609 (N_26609,N_22356,N_24088);
nor U26610 (N_26610,N_23347,N_23452);
nand U26611 (N_26611,N_20261,N_22083);
or U26612 (N_26612,N_24649,N_22383);
or U26613 (N_26613,N_22029,N_20001);
and U26614 (N_26614,N_22833,N_20195);
xor U26615 (N_26615,N_24209,N_22903);
xor U26616 (N_26616,N_21813,N_20325);
xor U26617 (N_26617,N_22405,N_20859);
nor U26618 (N_26618,N_23777,N_21874);
and U26619 (N_26619,N_21456,N_24228);
nand U26620 (N_26620,N_23238,N_22018);
nand U26621 (N_26621,N_21511,N_24195);
nand U26622 (N_26622,N_21699,N_21102);
and U26623 (N_26623,N_22168,N_24535);
and U26624 (N_26624,N_22095,N_20661);
or U26625 (N_26625,N_21126,N_23288);
nor U26626 (N_26626,N_21681,N_22515);
and U26627 (N_26627,N_22481,N_21147);
xor U26628 (N_26628,N_23518,N_24547);
and U26629 (N_26629,N_22279,N_21525);
or U26630 (N_26630,N_24907,N_22720);
and U26631 (N_26631,N_24268,N_21936);
and U26632 (N_26632,N_23817,N_23265);
or U26633 (N_26633,N_23803,N_20784);
and U26634 (N_26634,N_20847,N_24658);
xnor U26635 (N_26635,N_21950,N_20288);
nor U26636 (N_26636,N_23752,N_24131);
or U26637 (N_26637,N_24419,N_21898);
xnor U26638 (N_26638,N_23911,N_20903);
nor U26639 (N_26639,N_24745,N_23538);
xor U26640 (N_26640,N_23553,N_21066);
nor U26641 (N_26641,N_20570,N_22021);
and U26642 (N_26642,N_22034,N_23965);
xnor U26643 (N_26643,N_23135,N_24223);
nor U26644 (N_26644,N_24053,N_22237);
nand U26645 (N_26645,N_24588,N_20979);
nor U26646 (N_26646,N_24791,N_21636);
nand U26647 (N_26647,N_20809,N_20187);
xnor U26648 (N_26648,N_20825,N_20235);
and U26649 (N_26649,N_21190,N_22093);
xnor U26650 (N_26650,N_20095,N_22956);
xor U26651 (N_26651,N_20211,N_23476);
nand U26652 (N_26652,N_23181,N_24093);
nand U26653 (N_26653,N_21192,N_23341);
or U26654 (N_26654,N_20290,N_24499);
xor U26655 (N_26655,N_21054,N_21509);
and U26656 (N_26656,N_21038,N_23840);
xor U26657 (N_26657,N_23404,N_24168);
and U26658 (N_26658,N_21313,N_24650);
or U26659 (N_26659,N_24691,N_24962);
nand U26660 (N_26660,N_21416,N_21012);
xor U26661 (N_26661,N_24883,N_21240);
and U26662 (N_26662,N_22690,N_20934);
xnor U26663 (N_26663,N_22542,N_22065);
nor U26664 (N_26664,N_23445,N_21113);
xnor U26665 (N_26665,N_20406,N_22193);
and U26666 (N_26666,N_24274,N_22877);
nand U26667 (N_26667,N_20456,N_20309);
nand U26668 (N_26668,N_22190,N_24665);
nor U26669 (N_26669,N_20664,N_22823);
nor U26670 (N_26670,N_22860,N_20571);
and U26671 (N_26671,N_20032,N_23539);
xnor U26672 (N_26672,N_20212,N_20371);
nand U26673 (N_26673,N_20748,N_22518);
nand U26674 (N_26674,N_20384,N_23721);
nor U26675 (N_26675,N_23222,N_20342);
nor U26676 (N_26676,N_23858,N_21625);
nor U26677 (N_26677,N_20496,N_23552);
xor U26678 (N_26678,N_22600,N_21143);
xnor U26679 (N_26679,N_20128,N_24908);
and U26680 (N_26680,N_21755,N_20326);
xor U26681 (N_26681,N_20665,N_23930);
and U26682 (N_26682,N_24980,N_22398);
nand U26683 (N_26683,N_24404,N_24145);
and U26684 (N_26684,N_21890,N_23919);
or U26685 (N_26685,N_24521,N_21454);
or U26686 (N_26686,N_23869,N_20412);
nand U26687 (N_26687,N_20566,N_21324);
or U26688 (N_26688,N_23705,N_21845);
and U26689 (N_26689,N_21973,N_20671);
or U26690 (N_26690,N_20362,N_22943);
or U26691 (N_26691,N_20091,N_24655);
and U26692 (N_26692,N_21701,N_21386);
and U26693 (N_26693,N_20926,N_21139);
xnor U26694 (N_26694,N_24572,N_22382);
xor U26695 (N_26695,N_20536,N_21162);
and U26696 (N_26696,N_21243,N_24506);
and U26697 (N_26697,N_21706,N_24801);
nor U26698 (N_26698,N_22836,N_20817);
or U26699 (N_26699,N_20477,N_22714);
and U26700 (N_26700,N_20927,N_23940);
and U26701 (N_26701,N_21514,N_24812);
nand U26702 (N_26702,N_21527,N_20230);
nor U26703 (N_26703,N_24749,N_20533);
and U26704 (N_26704,N_22738,N_23945);
and U26705 (N_26705,N_24153,N_22741);
or U26706 (N_26706,N_22919,N_20059);
or U26707 (N_26707,N_22726,N_21884);
xnor U26708 (N_26708,N_22510,N_22880);
xnor U26709 (N_26709,N_23954,N_24896);
or U26710 (N_26710,N_21383,N_22636);
xor U26711 (N_26711,N_24283,N_24785);
xnor U26712 (N_26712,N_24185,N_21071);
xnor U26713 (N_26713,N_20758,N_23512);
nor U26714 (N_26714,N_20482,N_23026);
xnor U26715 (N_26715,N_24406,N_23034);
and U26716 (N_26716,N_22635,N_24284);
nand U26717 (N_26717,N_22736,N_22174);
or U26718 (N_26718,N_22099,N_22517);
nor U26719 (N_26719,N_23716,N_24451);
nor U26720 (N_26720,N_24453,N_23887);
or U26721 (N_26721,N_24605,N_22899);
nand U26722 (N_26722,N_21230,N_20776);
xor U26723 (N_26723,N_23156,N_23139);
nor U26724 (N_26724,N_20876,N_22591);
nand U26725 (N_26725,N_22976,N_22780);
xor U26726 (N_26726,N_20556,N_23855);
nor U26727 (N_26727,N_21477,N_20418);
xnor U26728 (N_26728,N_21466,N_22640);
nand U26729 (N_26729,N_21689,N_20546);
xor U26730 (N_26730,N_23101,N_22626);
or U26731 (N_26731,N_20425,N_20771);
nor U26732 (N_26732,N_22144,N_20801);
or U26733 (N_26733,N_21000,N_24176);
and U26734 (N_26734,N_24278,N_24292);
xnor U26735 (N_26735,N_21250,N_23586);
xor U26736 (N_26736,N_21368,N_24308);
nand U26737 (N_26737,N_21221,N_21217);
and U26738 (N_26738,N_21560,N_23033);
and U26739 (N_26739,N_24872,N_21709);
and U26740 (N_26740,N_21827,N_22946);
xnor U26741 (N_26741,N_20300,N_23745);
or U26742 (N_26742,N_23221,N_21932);
xor U26743 (N_26743,N_23011,N_20024);
and U26744 (N_26744,N_23256,N_21602);
nor U26745 (N_26745,N_23228,N_21429);
or U26746 (N_26746,N_23439,N_24936);
and U26747 (N_26747,N_20824,N_21330);
nand U26748 (N_26748,N_23020,N_21673);
and U26749 (N_26749,N_22300,N_23380);
nor U26750 (N_26750,N_21576,N_20173);
or U26751 (N_26751,N_22378,N_23284);
or U26752 (N_26752,N_21870,N_22003);
nor U26753 (N_26753,N_23191,N_24348);
nor U26754 (N_26754,N_20102,N_23225);
xor U26755 (N_26755,N_20363,N_23395);
nor U26756 (N_26756,N_22996,N_22032);
and U26757 (N_26757,N_22217,N_22548);
xor U26758 (N_26758,N_22616,N_20543);
nor U26759 (N_26759,N_21121,N_23730);
nor U26760 (N_26760,N_23549,N_21328);
or U26761 (N_26761,N_22187,N_22579);
nor U26762 (N_26762,N_21804,N_22711);
nand U26763 (N_26763,N_23004,N_20679);
xor U26764 (N_26764,N_23953,N_23075);
nor U26765 (N_26765,N_23950,N_23420);
xor U26766 (N_26766,N_24637,N_23628);
or U26767 (N_26767,N_20003,N_24312);
and U26768 (N_26768,N_23198,N_20554);
nor U26769 (N_26769,N_22583,N_20892);
xor U26770 (N_26770,N_21488,N_24469);
or U26771 (N_26771,N_23667,N_21404);
nor U26772 (N_26772,N_20315,N_24758);
nor U26773 (N_26773,N_21563,N_24075);
nand U26774 (N_26774,N_22013,N_21086);
or U26775 (N_26775,N_24373,N_20064);
or U26776 (N_26776,N_21343,N_22864);
and U26777 (N_26777,N_24189,N_23652);
nand U26778 (N_26778,N_22006,N_22843);
and U26779 (N_26779,N_22959,N_20615);
or U26780 (N_26780,N_23133,N_22581);
xnor U26781 (N_26781,N_20649,N_23806);
xor U26782 (N_26782,N_24494,N_23274);
xor U26783 (N_26783,N_20520,N_22460);
xor U26784 (N_26784,N_22893,N_23831);
nand U26785 (N_26785,N_22739,N_21280);
nand U26786 (N_26786,N_20925,N_21750);
xnor U26787 (N_26787,N_24994,N_23230);
nor U26788 (N_26788,N_20328,N_21412);
or U26789 (N_26789,N_23805,N_23871);
nor U26790 (N_26790,N_22914,N_24217);
and U26791 (N_26791,N_22024,N_20155);
nor U26792 (N_26792,N_20248,N_23833);
or U26793 (N_26793,N_22271,N_22129);
xor U26794 (N_26794,N_21100,N_21013);
or U26795 (N_26795,N_22947,N_20201);
nand U26796 (N_26796,N_23755,N_24710);
xor U26797 (N_26797,N_24647,N_24676);
nand U26798 (N_26798,N_21069,N_20842);
xor U26799 (N_26799,N_22842,N_23554);
and U26800 (N_26800,N_23541,N_24089);
or U26801 (N_26801,N_21465,N_20620);
and U26802 (N_26802,N_22050,N_23581);
and U26803 (N_26803,N_21355,N_21381);
nand U26804 (N_26804,N_24879,N_20567);
and U26805 (N_26805,N_22085,N_20731);
and U26806 (N_26806,N_22949,N_22929);
xor U26807 (N_26807,N_21210,N_23344);
or U26808 (N_26808,N_20839,N_20819);
nand U26809 (N_26809,N_24700,N_23776);
and U26810 (N_26810,N_23508,N_24125);
nor U26811 (N_26811,N_20775,N_24596);
nor U26812 (N_26812,N_22737,N_20527);
xnor U26813 (N_26813,N_24636,N_23466);
nor U26814 (N_26814,N_24621,N_20434);
nand U26815 (N_26815,N_20161,N_21578);
nor U26816 (N_26816,N_22256,N_23293);
and U26817 (N_26817,N_21128,N_22418);
nand U26818 (N_26818,N_21877,N_22131);
nand U26819 (N_26819,N_20708,N_21438);
nor U26820 (N_26820,N_20409,N_20814);
or U26821 (N_26821,N_20170,N_21034);
and U26822 (N_26822,N_20678,N_24091);
and U26823 (N_26823,N_22000,N_24455);
nor U26824 (N_26824,N_22679,N_22495);
nor U26825 (N_26825,N_21739,N_24207);
xnor U26826 (N_26826,N_22395,N_21974);
and U26827 (N_26827,N_20519,N_22619);
nor U26828 (N_26828,N_24107,N_21822);
xnor U26829 (N_26829,N_24508,N_22082);
nand U26830 (N_26830,N_21213,N_21638);
xor U26831 (N_26831,N_20250,N_22775);
or U26832 (N_26832,N_21125,N_21432);
or U26833 (N_26833,N_21787,N_20401);
or U26834 (N_26834,N_21110,N_21608);
and U26835 (N_26835,N_22421,N_22984);
and U26836 (N_26836,N_20938,N_21855);
nor U26837 (N_26837,N_20027,N_20668);
nor U26838 (N_26838,N_21157,N_24116);
and U26839 (N_26839,N_20871,N_22280);
or U26840 (N_26840,N_22126,N_22261);
and U26841 (N_26841,N_22968,N_21198);
or U26842 (N_26842,N_21537,N_20165);
and U26843 (N_26843,N_23679,N_23987);
nor U26844 (N_26844,N_20475,N_24440);
or U26845 (N_26845,N_24687,N_21583);
and U26846 (N_26846,N_22868,N_24456);
xnor U26847 (N_26847,N_22904,N_21044);
nor U26848 (N_26848,N_20270,N_24132);
nor U26849 (N_26849,N_21499,N_24930);
or U26850 (N_26850,N_21496,N_24793);
xnor U26851 (N_26851,N_20439,N_21011);
and U26852 (N_26852,N_21377,N_23088);
and U26853 (N_26853,N_21451,N_22594);
nand U26854 (N_26854,N_22355,N_24800);
xor U26855 (N_26855,N_24549,N_21986);
and U26856 (N_26856,N_23671,N_20950);
and U26857 (N_26857,N_22148,N_22785);
xor U26858 (N_26858,N_21312,N_21723);
nor U26859 (N_26859,N_24286,N_23184);
xnor U26860 (N_26860,N_20447,N_21055);
nor U26861 (N_26861,N_23162,N_22135);
or U26862 (N_26862,N_22423,N_23532);
xor U26863 (N_26863,N_24489,N_22399);
xor U26864 (N_26864,N_20457,N_22754);
and U26865 (N_26865,N_22080,N_24150);
or U26866 (N_26866,N_24273,N_21882);
and U26867 (N_26867,N_24550,N_23995);
nand U26868 (N_26868,N_21315,N_21867);
nand U26869 (N_26869,N_21606,N_24607);
xor U26870 (N_26870,N_24887,N_22539);
nand U26871 (N_26871,N_24413,N_20490);
xor U26872 (N_26872,N_20369,N_24859);
or U26873 (N_26873,N_23610,N_21630);
nand U26874 (N_26874,N_20052,N_21430);
or U26875 (N_26875,N_23821,N_23486);
nor U26876 (N_26876,N_22048,N_24893);
nor U26877 (N_26877,N_21446,N_23763);
or U26878 (N_26878,N_20939,N_20645);
or U26879 (N_26879,N_22245,N_23484);
nand U26880 (N_26880,N_24390,N_23684);
nand U26881 (N_26881,N_20319,N_24737);
nand U26882 (N_26882,N_23775,N_24393);
nand U26883 (N_26883,N_22326,N_22645);
nor U26884 (N_26884,N_22917,N_22408);
nand U26885 (N_26885,N_24083,N_21946);
or U26886 (N_26886,N_20605,N_21224);
or U26887 (N_26887,N_24208,N_23355);
and U26888 (N_26888,N_22822,N_22010);
and U26889 (N_26889,N_21334,N_24203);
xor U26890 (N_26890,N_22945,N_23568);
and U26891 (N_26891,N_24158,N_23921);
nor U26892 (N_26892,N_24590,N_23247);
nor U26893 (N_26893,N_24372,N_23620);
or U26894 (N_26894,N_22566,N_20531);
and U26895 (N_26895,N_23109,N_20157);
or U26896 (N_26896,N_22840,N_20149);
xnor U26897 (N_26897,N_22221,N_20864);
nor U26898 (N_26898,N_23085,N_20757);
nand U26899 (N_26899,N_24361,N_24360);
nand U26900 (N_26900,N_23045,N_21840);
nand U26901 (N_26901,N_20863,N_22427);
nand U26902 (N_26902,N_24471,N_24933);
xor U26903 (N_26903,N_20861,N_21106);
xnor U26904 (N_26904,N_24816,N_23778);
nor U26905 (N_26905,N_20327,N_21151);
or U26906 (N_26906,N_24573,N_23909);
or U26907 (N_26907,N_21385,N_22732);
and U26908 (N_26908,N_23419,N_22133);
nand U26909 (N_26909,N_23751,N_20387);
and U26910 (N_26910,N_20105,N_20734);
nor U26911 (N_26911,N_20780,N_21857);
nor U26912 (N_26912,N_20501,N_24643);
and U26913 (N_26913,N_23424,N_23888);
and U26914 (N_26914,N_22160,N_22351);
nor U26915 (N_26915,N_23650,N_24457);
or U26916 (N_26916,N_24029,N_23428);
nor U26917 (N_26917,N_21051,N_22981);
or U26918 (N_26918,N_21951,N_23904);
or U26919 (N_26919,N_23263,N_24881);
or U26920 (N_26920,N_23255,N_20512);
and U26921 (N_26921,N_21387,N_22556);
xnor U26922 (N_26922,N_23249,N_20377);
xor U26923 (N_26923,N_23129,N_20484);
nor U26924 (N_26924,N_23426,N_23925);
and U26925 (N_26925,N_23410,N_24174);
xor U26926 (N_26926,N_22372,N_22415);
xnor U26927 (N_26927,N_23732,N_22837);
nor U26928 (N_26928,N_22849,N_24396);
and U26929 (N_26929,N_23951,N_23218);
or U26930 (N_26930,N_21773,N_20960);
nand U26931 (N_26931,N_22652,N_24854);
nand U26932 (N_26932,N_22618,N_21861);
or U26933 (N_26933,N_24448,N_24612);
nor U26934 (N_26934,N_23145,N_24202);
or U26935 (N_26935,N_20232,N_23676);
xor U26936 (N_26936,N_24943,N_24220);
nand U26937 (N_26937,N_24628,N_20728);
nor U26938 (N_26938,N_22230,N_20142);
nor U26939 (N_26939,N_22857,N_20414);
xnor U26940 (N_26940,N_23655,N_20518);
nand U26941 (N_26941,N_22834,N_24731);
and U26942 (N_26942,N_22716,N_21104);
nand U26943 (N_26943,N_22520,N_24711);
nor U26944 (N_26944,N_23456,N_22360);
and U26945 (N_26945,N_23637,N_23702);
nor U26946 (N_26946,N_23363,N_22733);
and U26947 (N_26947,N_20011,N_22897);
xor U26948 (N_26948,N_22482,N_23823);
or U26949 (N_26949,N_20110,N_20602);
xor U26950 (N_26950,N_22890,N_23587);
xnor U26951 (N_26951,N_20766,N_23929);
nand U26952 (N_26952,N_22710,N_22936);
and U26953 (N_26953,N_23453,N_23574);
xnor U26954 (N_26954,N_24226,N_20470);
xor U26955 (N_26955,N_24119,N_20037);
nand U26956 (N_26956,N_20381,N_20422);
nor U26957 (N_26957,N_21931,N_20445);
nor U26958 (N_26958,N_21549,N_21977);
nor U26959 (N_26959,N_23630,N_24974);
and U26960 (N_26960,N_24340,N_20047);
nand U26961 (N_26961,N_21160,N_20404);
nor U26962 (N_26962,N_24515,N_20995);
nor U26963 (N_26963,N_22674,N_22953);
nor U26964 (N_26964,N_23593,N_22765);
and U26965 (N_26965,N_24706,N_21001);
or U26966 (N_26966,N_22203,N_24627);
xor U26967 (N_26967,N_24108,N_20865);
xor U26968 (N_26968,N_24778,N_23503);
nor U26969 (N_26969,N_21391,N_23122);
or U26970 (N_26970,N_21082,N_24215);
nand U26971 (N_26971,N_21258,N_20413);
or U26972 (N_26972,N_20621,N_24833);
nor U26973 (N_26973,N_23890,N_23790);
nand U26974 (N_26974,N_21979,N_23427);
or U26975 (N_26975,N_21005,N_21070);
nor U26976 (N_26976,N_22561,N_20534);
nor U26977 (N_26977,N_24940,N_23229);
nor U26978 (N_26978,N_24341,N_24599);
or U26979 (N_26979,N_20599,N_21255);
xor U26980 (N_26980,N_20993,N_20294);
nand U26981 (N_26981,N_22525,N_23864);
nand U26982 (N_26982,N_24822,N_24165);
xor U26983 (N_26983,N_21793,N_20827);
or U26984 (N_26984,N_22666,N_20285);
xor U26985 (N_26985,N_20240,N_23433);
and U26986 (N_26986,N_22342,N_21067);
and U26987 (N_26987,N_21156,N_20109);
xnor U26988 (N_26988,N_23464,N_23168);
and U26989 (N_26989,N_23578,N_23820);
and U26990 (N_26990,N_24134,N_24218);
xor U26991 (N_26991,N_22654,N_24235);
nor U26992 (N_26992,N_20985,N_22685);
or U26993 (N_26993,N_23340,N_20021);
xnor U26994 (N_26994,N_23696,N_21500);
and U26995 (N_26995,N_23119,N_21697);
or U26996 (N_26996,N_24828,N_23680);
xnor U26997 (N_26997,N_20831,N_23515);
and U26998 (N_26998,N_22767,N_23891);
xnor U26999 (N_26999,N_22348,N_23793);
or U27000 (N_27000,N_21505,N_24806);
and U27001 (N_27001,N_22376,N_23429);
or U27002 (N_27002,N_21746,N_24301);
nor U27003 (N_27003,N_24038,N_24660);
nand U27004 (N_27004,N_22536,N_21671);
and U27005 (N_27005,N_21008,N_23077);
nand U27006 (N_27006,N_22092,N_24311);
or U27007 (N_27007,N_24101,N_24040);
nor U27008 (N_27008,N_23359,N_24415);
nor U27009 (N_27009,N_20317,N_20089);
nor U27010 (N_27010,N_20147,N_21887);
nor U27011 (N_27011,N_21994,N_24037);
and U27012 (N_27012,N_24306,N_20094);
nand U27013 (N_27013,N_21058,N_22803);
and U27014 (N_27014,N_22623,N_21943);
or U27015 (N_27015,N_22592,N_20663);
and U27016 (N_27016,N_22715,N_24860);
or U27017 (N_27017,N_23239,N_22332);
and U27018 (N_27018,N_20981,N_22172);
or U27019 (N_27019,N_24843,N_23994);
nand U27020 (N_27020,N_23850,N_22535);
nand U27021 (N_27021,N_22673,N_24919);
or U27022 (N_27022,N_21284,N_20808);
and U27023 (N_27023,N_24868,N_23074);
or U27024 (N_27024,N_22485,N_24500);
and U27025 (N_27025,N_21645,N_24100);
xor U27026 (N_27026,N_23031,N_23394);
and U27027 (N_27027,N_23164,N_21265);
nand U27028 (N_27028,N_21469,N_20764);
xnor U27029 (N_27029,N_24307,N_20284);
and U27030 (N_27030,N_23915,N_23479);
nor U27031 (N_27031,N_21763,N_20282);
nand U27032 (N_27032,N_23972,N_23071);
and U27033 (N_27033,N_20346,N_23788);
nand U27034 (N_27034,N_22706,N_23220);
xor U27035 (N_27035,N_22719,N_24259);
nor U27036 (N_27036,N_23771,N_24562);
nor U27037 (N_27037,N_20912,N_23386);
xnor U27038 (N_27038,N_22896,N_21358);
nor U27039 (N_27039,N_24966,N_24401);
nand U27040 (N_27040,N_24981,N_24766);
xnor U27041 (N_27041,N_22607,N_20949);
or U27042 (N_27042,N_23989,N_24472);
xor U27043 (N_27043,N_21922,N_20510);
nor U27044 (N_27044,N_21481,N_21050);
nor U27045 (N_27045,N_23795,N_24269);
nand U27046 (N_27046,N_24197,N_23947);
or U27047 (N_27047,N_24553,N_22331);
and U27048 (N_27048,N_20225,N_23931);
and U27049 (N_27049,N_22796,N_20943);
and U27050 (N_27050,N_23212,N_22939);
and U27051 (N_27051,N_24316,N_22853);
or U27052 (N_27052,N_24394,N_24154);
or U27053 (N_27053,N_22777,N_23059);
or U27054 (N_27054,N_22496,N_24013);
nand U27055 (N_27055,N_21776,N_24447);
or U27056 (N_27056,N_22067,N_20062);
and U27057 (N_27057,N_24354,N_22030);
xnor U27058 (N_27058,N_24875,N_21155);
or U27059 (N_27059,N_22924,N_21459);
or U27060 (N_27060,N_24255,N_22205);
nor U27061 (N_27061,N_23973,N_20224);
nand U27062 (N_27062,N_20033,N_24997);
nand U27063 (N_27063,N_20099,N_23562);
or U27064 (N_27064,N_20424,N_23623);
xor U27065 (N_27065,N_24689,N_23470);
or U27066 (N_27066,N_23713,N_21144);
or U27067 (N_27067,N_24127,N_22429);
nand U27068 (N_27068,N_22682,N_24794);
and U27069 (N_27069,N_23112,N_24597);
or U27070 (N_27070,N_21337,N_21818);
xor U27071 (N_27071,N_20738,N_20502);
nor U27072 (N_27072,N_21545,N_21724);
and U27073 (N_27073,N_22219,N_23307);
nand U27074 (N_27074,N_23571,N_24629);
or U27075 (N_27075,N_24526,N_23098);
nor U27076 (N_27076,N_24951,N_20046);
nand U27077 (N_27077,N_24070,N_24477);
xor U27078 (N_27078,N_22569,N_22677);
nor U27079 (N_27079,N_20229,N_21910);
or U27080 (N_27080,N_20781,N_21123);
nand U27081 (N_27081,N_21331,N_23492);
or U27082 (N_27082,N_22662,N_24098);
and U27083 (N_27083,N_24729,N_22253);
xnor U27084 (N_27084,N_20515,N_23143);
nand U27085 (N_27085,N_22766,N_23865);
and U27086 (N_27086,N_21297,N_22016);
xor U27087 (N_27087,N_20185,N_21772);
and U27088 (N_27088,N_22354,N_24679);
or U27089 (N_27089,N_23379,N_20730);
xnor U27090 (N_27090,N_21618,N_23643);
xnor U27091 (N_27091,N_20584,N_22025);
and U27092 (N_27092,N_23246,N_20503);
nand U27093 (N_27093,N_21273,N_21293);
or U27094 (N_27094,N_21399,N_20183);
and U27095 (N_27095,N_23949,N_22453);
xor U27096 (N_27096,N_20803,N_23333);
or U27097 (N_27097,N_20403,N_21077);
nand U27098 (N_27098,N_23762,N_23959);
and U27099 (N_27099,N_21988,N_22551);
nand U27100 (N_27100,N_23907,N_20478);
and U27101 (N_27101,N_22426,N_21920);
xnor U27102 (N_27102,N_20117,N_22998);
xor U27103 (N_27103,N_23442,N_21871);
and U27104 (N_27104,N_22665,N_20374);
xnor U27105 (N_27105,N_24000,N_24085);
nor U27106 (N_27106,N_22123,N_21117);
xnor U27107 (N_27107,N_22627,N_24551);
xor U27108 (N_27108,N_21216,N_24008);
or U27109 (N_27109,N_24409,N_21816);
nand U27110 (N_27110,N_20698,N_24733);
or U27111 (N_27111,N_20277,N_21686);
xor U27112 (N_27112,N_20206,N_21542);
and U27113 (N_27113,N_20900,N_24819);
and U27114 (N_27114,N_20100,N_22513);
or U27115 (N_27115,N_23364,N_21768);
and U27116 (N_27116,N_21417,N_24808);
nand U27117 (N_27117,N_21939,N_21406);
xor U27118 (N_27118,N_20669,N_21271);
and U27119 (N_27119,N_21091,N_20822);
xnor U27120 (N_27120,N_24242,N_22062);
or U27121 (N_27121,N_23844,N_20959);
xnor U27122 (N_27122,N_24071,N_21674);
xor U27123 (N_27123,N_23832,N_20307);
nand U27124 (N_27124,N_23545,N_20168);
or U27125 (N_27125,N_20761,N_23548);
nor U27126 (N_27126,N_22176,N_22175);
nor U27127 (N_27127,N_24661,N_23633);
and U27128 (N_27128,N_21782,N_24742);
nor U27129 (N_27129,N_21494,N_24036);
and U27130 (N_27130,N_21229,N_21425);
nor U27131 (N_27131,N_21588,N_23441);
xor U27132 (N_27132,N_22576,N_22435);
xnor U27133 (N_27133,N_23529,N_21970);
nand U27134 (N_27134,N_20203,N_21888);
nor U27135 (N_27135,N_24606,N_21056);
nand U27136 (N_27136,N_24315,N_22634);
and U27137 (N_27137,N_23884,N_22494);
nor U27138 (N_27138,N_23656,N_23782);
xor U27139 (N_27139,N_20215,N_24905);
or U27140 (N_27140,N_22101,N_23376);
xnor U27141 (N_27141,N_20528,N_23704);
or U27142 (N_27142,N_20928,N_22417);
xnor U27143 (N_27143,N_24424,N_23392);
or U27144 (N_27144,N_23008,N_24552);
and U27145 (N_27145,N_21694,N_22819);
xnor U27146 (N_27146,N_21596,N_21757);
nor U27147 (N_27147,N_21460,N_23330);
nor U27148 (N_27148,N_20544,N_23266);
or U27149 (N_27149,N_22290,N_21978);
or U27150 (N_27150,N_20948,N_22621);
or U27151 (N_27151,N_22178,N_21573);
nor U27152 (N_27152,N_21883,N_23084);
nor U27153 (N_27153,N_22661,N_24991);
nand U27154 (N_27154,N_20623,N_23928);
xor U27155 (N_27155,N_24957,N_21515);
nand U27156 (N_27156,N_24239,N_22723);
xor U27157 (N_27157,N_22769,N_20564);
nor U27158 (N_27158,N_22119,N_20430);
and U27159 (N_27159,N_24147,N_21604);
xnor U27160 (N_27160,N_24498,N_24600);
nor U27161 (N_27161,N_20530,N_21521);
and U27162 (N_27162,N_20411,N_20426);
nand U27163 (N_27163,N_23108,N_22707);
xnor U27164 (N_27164,N_21254,N_22385);
nor U27165 (N_27165,N_20921,N_23400);
and U27166 (N_27166,N_24695,N_22471);
nor U27167 (N_27167,N_24598,N_22340);
or U27168 (N_27168,N_20851,N_21564);
nor U27169 (N_27169,N_21298,N_21605);
nand U27170 (N_27170,N_23875,N_21812);
and U27171 (N_27171,N_22786,N_21467);
nor U27172 (N_27172,N_23787,N_24592);
nand U27173 (N_27173,N_24750,N_20910);
xnor U27174 (N_27174,N_20143,N_21955);
nand U27175 (N_27175,N_23241,N_22761);
nor U27176 (N_27176,N_24275,N_22089);
nor U27177 (N_27177,N_21942,N_20691);
or U27178 (N_27178,N_24006,N_20778);
nand U27179 (N_27179,N_23205,N_22503);
nor U27180 (N_27180,N_24529,N_22467);
nand U27181 (N_27181,N_21236,N_22310);
and U27182 (N_27182,N_23187,N_24400);
or U27183 (N_27183,N_20525,N_22234);
nand U27184 (N_27184,N_23007,N_22327);
and U27185 (N_27185,N_24558,N_24864);
and U27186 (N_27186,N_24633,N_21356);
nor U27187 (N_27187,N_23434,N_20252);
nand U27188 (N_27188,N_21944,N_24917);
xnor U27189 (N_27189,N_21556,N_22602);
nand U27190 (N_27190,N_20647,N_20116);
nand U27191 (N_27191,N_20940,N_20145);
and U27192 (N_27192,N_24776,N_24452);
xor U27193 (N_27193,N_20491,N_21302);
nor U27194 (N_27194,N_24181,N_23918);
nor U27195 (N_27195,N_23794,N_21554);
xnor U27196 (N_27196,N_24673,N_24913);
xor U27197 (N_27197,N_22179,N_24509);
nand U27198 (N_27198,N_23859,N_21057);
nand U27199 (N_27199,N_23551,N_22572);
nor U27200 (N_27200,N_22889,N_22381);
xor U27201 (N_27201,N_22847,N_20952);
xor U27202 (N_27202,N_23968,N_24385);
or U27203 (N_27203,N_22353,N_23906);
or U27204 (N_27204,N_22544,N_22835);
nand U27205 (N_27205,N_21088,N_24680);
xor U27206 (N_27206,N_21078,N_20304);
xnor U27207 (N_27207,N_24130,N_21823);
nand U27208 (N_27208,N_24587,N_21344);
or U27209 (N_27209,N_24918,N_21594);
nand U27210 (N_27210,N_20541,N_21570);
and U27211 (N_27211,N_20929,N_23332);
nor U27212 (N_27212,N_23937,N_22522);
and U27213 (N_27213,N_21600,N_22249);
nand U27214 (N_27214,N_24076,N_23301);
nand U27215 (N_27215,N_22440,N_22509);
and U27216 (N_27216,N_22506,N_20022);
nand U27217 (N_27217,N_24164,N_22362);
and U27218 (N_27218,N_20015,N_21561);
nand U27219 (N_27219,N_22107,N_21184);
xnor U27220 (N_27220,N_24939,N_24741);
nand U27221 (N_27221,N_21470,N_24694);
or U27222 (N_27222,N_21893,N_20557);
nor U27223 (N_27223,N_20656,N_23727);
or U27224 (N_27224,N_23687,N_21775);
or U27225 (N_27225,N_22321,N_20638);
and U27226 (N_27226,N_24304,N_20438);
or U27227 (N_27227,N_23594,N_21765);
nor U27228 (N_27228,N_21169,N_21296);
nor U27229 (N_27229,N_20280,N_23132);
and U27230 (N_27230,N_20509,N_20965);
or U27231 (N_27231,N_22989,N_20092);
and U27232 (N_27232,N_23933,N_21743);
or U27233 (N_27233,N_23063,N_20420);
and U27234 (N_27234,N_23647,N_23294);
xor U27235 (N_27235,N_24559,N_20352);
and U27236 (N_27236,N_24823,N_20074);
xor U27237 (N_27237,N_21239,N_23608);
and U27238 (N_27238,N_24261,N_22268);
or U27239 (N_27239,N_24182,N_21968);
and U27240 (N_27240,N_23923,N_21653);
and U27241 (N_27241,N_20516,N_22926);
and U27242 (N_27242,N_24140,N_21574);
or U27243 (N_27243,N_20009,N_21734);
nand U27244 (N_27244,N_22832,N_20862);
xor U27245 (N_27245,N_20804,N_22975);
nand U27246 (N_27246,N_24662,N_23372);
nand U27247 (N_27247,N_23163,N_24058);
xnor U27248 (N_27248,N_23431,N_23619);
or U27249 (N_27249,N_24837,N_20223);
or U27250 (N_27250,N_22039,N_20958);
nor U27251 (N_27251,N_22575,N_22315);
nand U27252 (N_27252,N_21555,N_24177);
xnor U27253 (N_27253,N_22855,N_20703);
and U27254 (N_27254,N_22269,N_21257);
and U27255 (N_27255,N_24179,N_20682);
nor U27256 (N_27256,N_24748,N_21954);
or U27257 (N_27257,N_24982,N_20966);
nand U27258 (N_27258,N_24297,N_21002);
nand U27259 (N_27259,N_23407,N_21461);
xnor U27260 (N_27260,N_23605,N_24639);
and U27261 (N_27261,N_24488,N_22845);
nand U27262 (N_27262,N_22410,N_20137);
xor U27263 (N_27263,N_20228,N_21299);
nand U27264 (N_27264,N_21786,N_23469);
and U27265 (N_27265,N_20415,N_21646);
and U27266 (N_27266,N_22934,N_23001);
xor U27267 (N_27267,N_23058,N_22629);
xor U27268 (N_27268,N_21407,N_21751);
nor U27269 (N_27269,N_21133,N_23521);
and U27270 (N_27270,N_24332,N_23712);
nand U27271 (N_27271,N_23768,N_24814);
nand U27272 (N_27272,N_24937,N_21074);
nand U27273 (N_27273,N_23079,N_24577);
or U27274 (N_27274,N_23692,N_24368);
and U27275 (N_27275,N_23897,N_20795);
or U27276 (N_27276,N_23295,N_20779);
or U27277 (N_27277,N_24956,N_20200);
nand U27278 (N_27278,N_22982,N_22571);
xnor U27279 (N_27279,N_20899,N_20989);
xnor U27280 (N_27280,N_24120,N_20489);
and U27281 (N_27281,N_23513,N_20935);
nor U27282 (N_27282,N_24527,N_23955);
nand U27283 (N_27283,N_24569,N_21695);
nand U27284 (N_27284,N_22727,N_21546);
and U27285 (N_27285,N_23041,N_20361);
nor U27286 (N_27286,N_21260,N_20118);
nor U27287 (N_27287,N_22935,N_23560);
or U27288 (N_27288,N_23993,N_24684);
nor U27289 (N_27289,N_22960,N_22977);
xor U27290 (N_27290,N_22567,N_23885);
nand U27291 (N_27291,N_20631,N_21269);
or U27292 (N_27292,N_22140,N_23367);
xnor U27293 (N_27293,N_22955,N_22357);
or U27294 (N_27294,N_21285,N_24586);
nor U27295 (N_27295,N_23559,N_21672);
nor U27296 (N_27296,N_21349,N_23800);
and U27297 (N_27297,N_23403,N_23141);
and U27298 (N_27298,N_22247,N_22593);
and U27299 (N_27299,N_20797,N_24028);
xor U27300 (N_27300,N_22045,N_24214);
nand U27301 (N_27301,N_20652,N_24339);
xor U27302 (N_27302,N_23990,N_20391);
or U27303 (N_27303,N_23377,N_24081);
and U27304 (N_27304,N_22056,N_23576);
and U27305 (N_27305,N_22745,N_22820);
nand U27306 (N_27306,N_23157,N_21132);
and U27307 (N_27307,N_20004,N_22235);
nand U27308 (N_27308,N_23412,N_22311);
xor U27309 (N_27309,N_20481,N_20931);
or U27310 (N_27310,N_23811,N_24999);
nor U27311 (N_27311,N_21176,N_22708);
and U27312 (N_27312,N_21722,N_24591);
nand U27313 (N_27313,N_24969,N_22580);
nand U27314 (N_27314,N_21654,N_24921);
and U27315 (N_27315,N_23351,N_21909);
and U27316 (N_27316,N_24180,N_21971);
and U27317 (N_27317,N_21320,N_20279);
and U27318 (N_27318,N_20039,N_22699);
or U27319 (N_27319,N_20217,N_23378);
nor U27320 (N_27320,N_24052,N_20488);
nand U27321 (N_27321,N_22218,N_20302);
xnor U27322 (N_27322,N_24510,N_21829);
or U27323 (N_27323,N_21241,N_20969);
and U27324 (N_27324,N_21080,N_22698);
xor U27325 (N_27325,N_21129,N_23319);
nand U27326 (N_27326,N_22965,N_21036);
nand U27327 (N_27327,N_23192,N_23271);
or U27328 (N_27328,N_22015,N_22624);
xor U27329 (N_27329,N_24682,N_20397);
nand U27330 (N_27330,N_21998,N_22649);
xor U27331 (N_27331,N_20553,N_24578);
and U27332 (N_27332,N_23822,N_23892);
nor U27333 (N_27333,N_22066,N_21188);
nand U27334 (N_27334,N_22671,N_21165);
nand U27335 (N_27335,N_23009,N_23816);
nor U27336 (N_27336,N_21492,N_20906);
and U27337 (N_27337,N_21894,N_23640);
and U27338 (N_27338,N_20030,N_21426);
or U27339 (N_27339,N_20746,N_23053);
and U27340 (N_27340,N_23903,N_24768);
nor U27341 (N_27341,N_20473,N_21914);
nand U27342 (N_27342,N_20071,N_24138);
nand U27343 (N_27343,N_23982,N_24376);
and U27344 (N_27344,N_22874,N_21409);
nand U27345 (N_27345,N_23766,N_22367);
nor U27346 (N_27346,N_21558,N_22053);
xnor U27347 (N_27347,N_24686,N_20350);
xnor U27348 (N_27348,N_23178,N_20251);
nor U27349 (N_27349,N_20747,N_22852);
nor U27350 (N_27350,N_24538,N_20273);
nor U27351 (N_27351,N_20171,N_20701);
nor U27352 (N_27352,N_24257,N_20209);
xnor U27353 (N_27353,N_21361,N_22419);
xor U27354 (N_27354,N_20895,N_21741);
nand U27355 (N_27355,N_20833,N_23974);
xnor U27356 (N_27356,N_24613,N_22458);
xor U27357 (N_27357,N_22801,N_24025);
or U27358 (N_27358,N_23040,N_20914);
nor U27359 (N_27359,N_21924,N_22057);
or U27360 (N_27360,N_22817,N_20707);
or U27361 (N_27361,N_23044,N_24430);
xor U27362 (N_27362,N_22678,N_24702);
or U27363 (N_27363,N_24043,N_21336);
nand U27364 (N_27364,N_20440,N_21253);
and U27365 (N_27365,N_22023,N_23250);
or U27366 (N_27366,N_22086,N_22827);
or U27367 (N_27367,N_24438,N_22555);
xor U27368 (N_27368,N_20880,N_23383);
or U27369 (N_27369,N_21762,N_24985);
nor U27370 (N_27370,N_22336,N_24364);
and U27371 (N_27371,N_24708,N_22866);
nor U27372 (N_27372,N_20340,N_24614);
nand U27373 (N_27373,N_20453,N_20583);
xnor U27374 (N_27374,N_24247,N_24820);
nand U27375 (N_27375,N_23245,N_24391);
or U27376 (N_27376,N_23106,N_23261);
xor U27377 (N_27377,N_20685,N_20123);
or U27378 (N_27378,N_22879,N_24652);
and U27379 (N_27379,N_23975,N_22541);
or U27380 (N_27380,N_23618,N_23710);
and U27381 (N_27381,N_20442,N_24161);
nand U27382 (N_27382,N_22484,N_24344);
xor U27383 (N_27383,N_24927,N_24320);
nand U27384 (N_27384,N_22742,N_21854);
xnor U27385 (N_27385,N_23798,N_23480);
nor U27386 (N_27386,N_23689,N_20329);
nor U27387 (N_27387,N_21802,N_22601);
and U27388 (N_27388,N_23769,N_22987);
xnor U27389 (N_27389,N_24423,N_21677);
and U27390 (N_27390,N_23922,N_20045);
xnor U27391 (N_27391,N_24903,N_22930);
or U27392 (N_27392,N_20194,N_20885);
and U27393 (N_27393,N_20751,N_20837);
or U27394 (N_27394,N_23165,N_24645);
nand U27395 (N_27395,N_23305,N_24378);
nor U27396 (N_27396,N_23114,N_23765);
nor U27397 (N_27397,N_23958,N_24381);
nor U27398 (N_27398,N_20246,N_20193);
nor U27399 (N_27399,N_22138,N_24113);
xnor U27400 (N_27400,N_24678,N_22560);
and U27401 (N_27401,N_24876,N_20523);
and U27402 (N_27402,N_24683,N_20134);
nor U27403 (N_27403,N_23882,N_21575);
nand U27404 (N_27404,N_23296,N_24856);
nand U27405 (N_27405,N_23917,N_23493);
nand U27406 (N_27406,N_22725,N_20787);
and U27407 (N_27407,N_21669,N_23123);
nor U27408 (N_27408,N_20857,N_21927);
nand U27409 (N_27409,N_24570,N_22603);
nor U27410 (N_27410,N_24632,N_22686);
or U27411 (N_27411,N_24252,N_23561);
nor U27412 (N_27412,N_21272,N_24756);
nor U27413 (N_27413,N_22061,N_23138);
nor U27414 (N_27414,N_21926,N_21390);
and U27415 (N_27415,N_24792,N_22124);
nor U27416 (N_27416,N_22322,N_20932);
nand U27417 (N_27417,N_20522,N_22343);
xnor U27418 (N_27418,N_23358,N_23780);
or U27419 (N_27419,N_22611,N_20226);
and U27420 (N_27420,N_21491,N_24211);
nor U27421 (N_27421,N_20334,N_24117);
and U27422 (N_27422,N_21937,N_23813);
nand U27423 (N_27423,N_24944,N_22201);
xor U27424 (N_27424,N_22043,N_22104);
xor U27425 (N_27425,N_20710,N_20231);
or U27426 (N_27426,N_23361,N_23345);
nor U27427 (N_27427,N_24848,N_23346);
or U27428 (N_27428,N_22937,N_22132);
and U27429 (N_27429,N_24408,N_21183);
xnor U27430 (N_27430,N_22287,N_24346);
nor U27431 (N_27431,N_23880,N_24925);
nand U27432 (N_27432,N_22465,N_22991);
and U27433 (N_27433,N_22451,N_24206);
nor U27434 (N_27434,N_22459,N_21099);
and U27435 (N_27435,N_23454,N_21915);
and U27436 (N_27436,N_20988,N_20405);
or U27437 (N_27437,N_22599,N_21483);
and U27438 (N_27438,N_23847,N_24651);
xnor U27439 (N_27439,N_20236,N_23807);
xnor U27440 (N_27440,N_22731,N_22275);
nand U27441 (N_27441,N_21263,N_21420);
nor U27442 (N_27442,N_22344,N_21415);
or U27443 (N_27443,N_23211,N_24056);
or U27444 (N_27444,N_20141,N_21841);
nand U27445 (N_27445,N_24224,N_22229);
or U27446 (N_27446,N_21189,N_21824);
and U27447 (N_27447,N_23718,N_23190);
nor U27448 (N_27448,N_23842,N_21502);
and U27449 (N_27449,N_22979,N_21266);
and U27450 (N_27450,N_24102,N_24291);
xor U27451 (N_27451,N_21639,N_24328);
nor U27452 (N_27452,N_24227,N_24184);
and U27453 (N_27453,N_22339,N_23818);
nand U27454 (N_27454,N_21559,N_23174);
or U27455 (N_27455,N_22468,N_23877);
and U27456 (N_27456,N_23572,N_21475);
xor U27457 (N_27457,N_24824,N_23981);
or U27458 (N_27458,N_23948,N_24044);
xor U27459 (N_27459,N_24880,N_24789);
nand U27460 (N_27460,N_21568,N_21180);
nand U27461 (N_27461,N_24343,N_20815);
nor U27462 (N_27462,N_22241,N_23985);
nand U27463 (N_27463,N_22375,N_20070);
and U27464 (N_27464,N_20813,N_24086);
or U27465 (N_27465,N_22297,N_23447);
nand U27466 (N_27466,N_20454,N_20016);
or U27467 (N_27467,N_22760,N_23760);
nand U27468 (N_27468,N_22422,N_21912);
xnor U27469 (N_27469,N_23744,N_22740);
nand U27470 (N_27470,N_24336,N_20637);
nor U27471 (N_27471,N_22540,N_21819);
xor U27472 (N_27472,N_24458,N_23389);
and U27473 (N_27473,N_20086,N_23912);
or U27474 (N_27474,N_23677,N_21378);
nor U27475 (N_27475,N_23067,N_24198);
or U27476 (N_27476,N_21597,N_23369);
nor U27477 (N_27477,N_23065,N_20617);
nand U27478 (N_27478,N_21552,N_22828);
nor U27479 (N_27479,N_21173,N_21700);
xor U27480 (N_27480,N_21989,N_21785);
or U27481 (N_27481,N_20601,N_21042);
or U27482 (N_27482,N_22839,N_24963);
and U27483 (N_27483,N_23125,N_21534);
nand U27484 (N_27484,N_22643,N_24272);
and U27485 (N_27485,N_21003,N_23590);
and U27486 (N_27486,N_22004,N_22404);
nor U27487 (N_27487,N_21809,N_22128);
and U27488 (N_27488,N_22642,N_23144);
xor U27489 (N_27489,N_23789,N_21291);
and U27490 (N_27490,N_24351,N_22324);
xnor U27491 (N_27491,N_21789,N_24853);
and U27492 (N_27492,N_22283,N_20513);
nor U27493 (N_27493,N_20124,N_20642);
and U27494 (N_27494,N_22306,N_24427);
and U27495 (N_27495,N_24610,N_21551);
nand U27496 (N_27496,N_20579,N_20733);
nand U27497 (N_27497,N_21140,N_22227);
nand U27498 (N_27498,N_22697,N_20610);
nor U27499 (N_27499,N_21518,N_24199);
xnor U27500 (N_27500,N_24346,N_24746);
or U27501 (N_27501,N_20013,N_24944);
nor U27502 (N_27502,N_24777,N_22695);
xor U27503 (N_27503,N_21827,N_20869);
nor U27504 (N_27504,N_20490,N_23561);
nor U27505 (N_27505,N_23597,N_23176);
or U27506 (N_27506,N_22215,N_23927);
nor U27507 (N_27507,N_23102,N_22476);
and U27508 (N_27508,N_20342,N_21176);
and U27509 (N_27509,N_24991,N_22441);
nor U27510 (N_27510,N_20662,N_21282);
and U27511 (N_27511,N_24309,N_20028);
nor U27512 (N_27512,N_22838,N_21139);
nand U27513 (N_27513,N_24191,N_23134);
nand U27514 (N_27514,N_24306,N_20759);
nand U27515 (N_27515,N_22927,N_23869);
nand U27516 (N_27516,N_21398,N_22451);
xor U27517 (N_27517,N_22511,N_23685);
nor U27518 (N_27518,N_23122,N_23318);
and U27519 (N_27519,N_20245,N_22734);
and U27520 (N_27520,N_21126,N_24135);
or U27521 (N_27521,N_22265,N_23131);
xnor U27522 (N_27522,N_24640,N_24216);
or U27523 (N_27523,N_22424,N_20185);
or U27524 (N_27524,N_24251,N_22514);
and U27525 (N_27525,N_20859,N_24397);
nand U27526 (N_27526,N_21529,N_20958);
xnor U27527 (N_27527,N_21890,N_23483);
and U27528 (N_27528,N_23880,N_23287);
xnor U27529 (N_27529,N_23403,N_22436);
xor U27530 (N_27530,N_24900,N_22691);
nor U27531 (N_27531,N_22501,N_21214);
nor U27532 (N_27532,N_22455,N_22253);
and U27533 (N_27533,N_23264,N_24096);
or U27534 (N_27534,N_23774,N_24594);
nor U27535 (N_27535,N_21745,N_20520);
xor U27536 (N_27536,N_21056,N_24197);
or U27537 (N_27537,N_24518,N_22956);
xor U27538 (N_27538,N_23592,N_22219);
xor U27539 (N_27539,N_22006,N_24662);
nor U27540 (N_27540,N_22000,N_22768);
nand U27541 (N_27541,N_23899,N_24330);
xor U27542 (N_27542,N_20413,N_22024);
and U27543 (N_27543,N_20601,N_21983);
and U27544 (N_27544,N_22190,N_23060);
nand U27545 (N_27545,N_21409,N_23727);
xor U27546 (N_27546,N_24538,N_20237);
and U27547 (N_27547,N_24360,N_20171);
nand U27548 (N_27548,N_20165,N_21502);
nor U27549 (N_27549,N_24256,N_24222);
and U27550 (N_27550,N_23662,N_23649);
nand U27551 (N_27551,N_23173,N_22984);
xor U27552 (N_27552,N_22611,N_23727);
nor U27553 (N_27553,N_20163,N_22782);
nand U27554 (N_27554,N_22690,N_23026);
xnor U27555 (N_27555,N_24814,N_20524);
nor U27556 (N_27556,N_20525,N_22375);
nand U27557 (N_27557,N_20801,N_21035);
nor U27558 (N_27558,N_22303,N_23129);
nor U27559 (N_27559,N_22031,N_20437);
or U27560 (N_27560,N_20310,N_23674);
and U27561 (N_27561,N_22506,N_21042);
and U27562 (N_27562,N_24895,N_24606);
and U27563 (N_27563,N_20307,N_23838);
nand U27564 (N_27564,N_22151,N_23102);
nand U27565 (N_27565,N_20073,N_21384);
or U27566 (N_27566,N_23246,N_23828);
nand U27567 (N_27567,N_22246,N_24099);
nand U27568 (N_27568,N_22215,N_24976);
and U27569 (N_27569,N_21887,N_20405);
or U27570 (N_27570,N_21968,N_21538);
xnor U27571 (N_27571,N_22105,N_24150);
and U27572 (N_27572,N_23813,N_20004);
or U27573 (N_27573,N_23096,N_22620);
nand U27574 (N_27574,N_21729,N_23822);
or U27575 (N_27575,N_23712,N_23133);
xor U27576 (N_27576,N_23205,N_21924);
nor U27577 (N_27577,N_23794,N_21891);
nand U27578 (N_27578,N_21463,N_22390);
nor U27579 (N_27579,N_20092,N_22802);
and U27580 (N_27580,N_22325,N_22114);
or U27581 (N_27581,N_21773,N_22872);
or U27582 (N_27582,N_23021,N_23376);
and U27583 (N_27583,N_24099,N_23657);
or U27584 (N_27584,N_23727,N_21827);
xor U27585 (N_27585,N_23392,N_23399);
or U27586 (N_27586,N_22735,N_21453);
nand U27587 (N_27587,N_24315,N_22233);
nand U27588 (N_27588,N_24122,N_24764);
and U27589 (N_27589,N_22351,N_22871);
xor U27590 (N_27590,N_22582,N_23545);
xor U27591 (N_27591,N_24890,N_24907);
xnor U27592 (N_27592,N_21642,N_23565);
xnor U27593 (N_27593,N_20984,N_24003);
and U27594 (N_27594,N_23257,N_21862);
or U27595 (N_27595,N_22587,N_21174);
nor U27596 (N_27596,N_24411,N_22791);
nand U27597 (N_27597,N_24752,N_20059);
or U27598 (N_27598,N_22396,N_21831);
or U27599 (N_27599,N_21711,N_24241);
xor U27600 (N_27600,N_23247,N_24501);
and U27601 (N_27601,N_22939,N_24122);
or U27602 (N_27602,N_20801,N_21603);
nor U27603 (N_27603,N_20235,N_22418);
nand U27604 (N_27604,N_24773,N_24176);
xor U27605 (N_27605,N_23846,N_23538);
or U27606 (N_27606,N_24835,N_20897);
or U27607 (N_27607,N_23639,N_22797);
xnor U27608 (N_27608,N_20274,N_23021);
xnor U27609 (N_27609,N_24571,N_21433);
nand U27610 (N_27610,N_22447,N_21505);
xor U27611 (N_27611,N_21747,N_23118);
and U27612 (N_27612,N_20641,N_20343);
xor U27613 (N_27613,N_24003,N_20845);
xor U27614 (N_27614,N_20837,N_21840);
nand U27615 (N_27615,N_23431,N_23901);
and U27616 (N_27616,N_24463,N_20447);
or U27617 (N_27617,N_23785,N_20229);
xnor U27618 (N_27618,N_22239,N_23277);
nor U27619 (N_27619,N_22069,N_22738);
and U27620 (N_27620,N_21241,N_23358);
xnor U27621 (N_27621,N_21294,N_21710);
and U27622 (N_27622,N_20877,N_22265);
and U27623 (N_27623,N_23105,N_22322);
and U27624 (N_27624,N_20230,N_22212);
nand U27625 (N_27625,N_20941,N_20358);
nor U27626 (N_27626,N_22134,N_24432);
nand U27627 (N_27627,N_22200,N_22681);
nand U27628 (N_27628,N_22266,N_23488);
xnor U27629 (N_27629,N_20644,N_23867);
nand U27630 (N_27630,N_24604,N_23986);
and U27631 (N_27631,N_22311,N_24057);
or U27632 (N_27632,N_21162,N_22025);
xnor U27633 (N_27633,N_21504,N_23706);
and U27634 (N_27634,N_22347,N_24823);
or U27635 (N_27635,N_21228,N_21633);
and U27636 (N_27636,N_24843,N_23093);
and U27637 (N_27637,N_20621,N_21735);
and U27638 (N_27638,N_24062,N_23541);
and U27639 (N_27639,N_21192,N_22702);
nor U27640 (N_27640,N_23697,N_24432);
xnor U27641 (N_27641,N_23517,N_24766);
xor U27642 (N_27642,N_20215,N_23082);
nor U27643 (N_27643,N_20313,N_24015);
nand U27644 (N_27644,N_24104,N_21105);
or U27645 (N_27645,N_23579,N_21156);
xor U27646 (N_27646,N_24727,N_21930);
nor U27647 (N_27647,N_23189,N_24108);
nand U27648 (N_27648,N_22914,N_23842);
or U27649 (N_27649,N_21020,N_22998);
or U27650 (N_27650,N_22456,N_23382);
and U27651 (N_27651,N_23093,N_24048);
xor U27652 (N_27652,N_20043,N_24104);
nor U27653 (N_27653,N_24626,N_22336);
nor U27654 (N_27654,N_24091,N_21125);
or U27655 (N_27655,N_22414,N_20951);
xor U27656 (N_27656,N_24317,N_20619);
and U27657 (N_27657,N_24334,N_20953);
nor U27658 (N_27658,N_23194,N_23808);
or U27659 (N_27659,N_20274,N_23806);
or U27660 (N_27660,N_24329,N_23746);
nand U27661 (N_27661,N_21049,N_22046);
nand U27662 (N_27662,N_21675,N_23810);
nor U27663 (N_27663,N_22275,N_24944);
xnor U27664 (N_27664,N_20537,N_23116);
and U27665 (N_27665,N_21298,N_21034);
xor U27666 (N_27666,N_20256,N_23522);
or U27667 (N_27667,N_23294,N_21468);
xnor U27668 (N_27668,N_24243,N_22153);
nor U27669 (N_27669,N_21307,N_22760);
or U27670 (N_27670,N_20970,N_23882);
nor U27671 (N_27671,N_23255,N_23711);
and U27672 (N_27672,N_23332,N_21782);
nor U27673 (N_27673,N_22441,N_23407);
or U27674 (N_27674,N_21908,N_21498);
and U27675 (N_27675,N_20930,N_24650);
or U27676 (N_27676,N_24621,N_20258);
and U27677 (N_27677,N_22586,N_24469);
or U27678 (N_27678,N_23597,N_20507);
nor U27679 (N_27679,N_22695,N_23944);
or U27680 (N_27680,N_23465,N_22295);
nor U27681 (N_27681,N_23724,N_20080);
or U27682 (N_27682,N_21111,N_24592);
nand U27683 (N_27683,N_21794,N_24720);
nand U27684 (N_27684,N_23423,N_20683);
xnor U27685 (N_27685,N_20014,N_22282);
nand U27686 (N_27686,N_20546,N_24762);
nor U27687 (N_27687,N_22293,N_21057);
nor U27688 (N_27688,N_23702,N_23042);
xor U27689 (N_27689,N_22821,N_23660);
nand U27690 (N_27690,N_24112,N_24818);
or U27691 (N_27691,N_21393,N_20413);
nand U27692 (N_27692,N_22980,N_21065);
or U27693 (N_27693,N_24880,N_22150);
nor U27694 (N_27694,N_20826,N_23251);
xor U27695 (N_27695,N_23451,N_24564);
xor U27696 (N_27696,N_24140,N_20282);
nand U27697 (N_27697,N_20996,N_24351);
xor U27698 (N_27698,N_20893,N_24823);
and U27699 (N_27699,N_20359,N_22724);
and U27700 (N_27700,N_20357,N_20485);
and U27701 (N_27701,N_22181,N_24092);
xnor U27702 (N_27702,N_24147,N_24768);
or U27703 (N_27703,N_23614,N_23394);
or U27704 (N_27704,N_21688,N_21109);
nor U27705 (N_27705,N_20065,N_21219);
xor U27706 (N_27706,N_23228,N_20011);
xor U27707 (N_27707,N_21348,N_23246);
nand U27708 (N_27708,N_23067,N_20105);
nor U27709 (N_27709,N_20927,N_22280);
xor U27710 (N_27710,N_24078,N_20607);
and U27711 (N_27711,N_23121,N_20296);
and U27712 (N_27712,N_22467,N_24450);
nor U27713 (N_27713,N_21361,N_24233);
nor U27714 (N_27714,N_21015,N_20651);
xor U27715 (N_27715,N_24244,N_24461);
or U27716 (N_27716,N_22915,N_23352);
and U27717 (N_27717,N_24675,N_20706);
or U27718 (N_27718,N_23633,N_21048);
or U27719 (N_27719,N_20713,N_24403);
nor U27720 (N_27720,N_22343,N_20985);
or U27721 (N_27721,N_21367,N_23682);
xor U27722 (N_27722,N_21178,N_21796);
nor U27723 (N_27723,N_20075,N_22043);
nand U27724 (N_27724,N_24178,N_22785);
and U27725 (N_27725,N_23532,N_24840);
or U27726 (N_27726,N_20938,N_24797);
and U27727 (N_27727,N_23436,N_21784);
nand U27728 (N_27728,N_23231,N_21889);
xor U27729 (N_27729,N_23712,N_21464);
nor U27730 (N_27730,N_21824,N_22491);
nor U27731 (N_27731,N_22545,N_21565);
and U27732 (N_27732,N_24684,N_24983);
or U27733 (N_27733,N_20299,N_21343);
or U27734 (N_27734,N_24360,N_20628);
or U27735 (N_27735,N_21934,N_20993);
nor U27736 (N_27736,N_22047,N_23705);
nand U27737 (N_27737,N_20227,N_22080);
nand U27738 (N_27738,N_24915,N_21792);
or U27739 (N_27739,N_21654,N_20438);
nand U27740 (N_27740,N_23296,N_20360);
xor U27741 (N_27741,N_21159,N_21558);
nor U27742 (N_27742,N_24329,N_22995);
or U27743 (N_27743,N_23791,N_21863);
nand U27744 (N_27744,N_20283,N_21279);
nor U27745 (N_27745,N_24205,N_20318);
nor U27746 (N_27746,N_21266,N_22689);
nor U27747 (N_27747,N_21226,N_23343);
nand U27748 (N_27748,N_24149,N_23302);
or U27749 (N_27749,N_22931,N_22525);
nand U27750 (N_27750,N_23349,N_22061);
xnor U27751 (N_27751,N_20496,N_24009);
xor U27752 (N_27752,N_20794,N_24455);
or U27753 (N_27753,N_22307,N_21860);
nand U27754 (N_27754,N_21571,N_20500);
and U27755 (N_27755,N_21071,N_22705);
nor U27756 (N_27756,N_20825,N_23029);
xnor U27757 (N_27757,N_23052,N_22750);
and U27758 (N_27758,N_23400,N_21886);
nor U27759 (N_27759,N_23822,N_24827);
nor U27760 (N_27760,N_22014,N_20952);
xor U27761 (N_27761,N_21693,N_20920);
nor U27762 (N_27762,N_23912,N_23469);
nor U27763 (N_27763,N_24824,N_21577);
and U27764 (N_27764,N_23430,N_22408);
nor U27765 (N_27765,N_23267,N_21252);
nand U27766 (N_27766,N_22008,N_24385);
and U27767 (N_27767,N_23196,N_23531);
and U27768 (N_27768,N_23026,N_20093);
and U27769 (N_27769,N_24946,N_20553);
xnor U27770 (N_27770,N_22787,N_24780);
and U27771 (N_27771,N_24861,N_24475);
nor U27772 (N_27772,N_22370,N_24958);
nand U27773 (N_27773,N_22608,N_20228);
nor U27774 (N_27774,N_24415,N_21662);
or U27775 (N_27775,N_24197,N_23079);
or U27776 (N_27776,N_21371,N_24401);
nand U27777 (N_27777,N_21520,N_20076);
and U27778 (N_27778,N_21758,N_24407);
nand U27779 (N_27779,N_21236,N_23059);
nand U27780 (N_27780,N_23457,N_24925);
nor U27781 (N_27781,N_24547,N_23257);
nand U27782 (N_27782,N_20634,N_23789);
xnor U27783 (N_27783,N_23350,N_23933);
and U27784 (N_27784,N_21859,N_20665);
or U27785 (N_27785,N_21443,N_23796);
and U27786 (N_27786,N_23124,N_23633);
and U27787 (N_27787,N_24401,N_20793);
and U27788 (N_27788,N_22702,N_20168);
and U27789 (N_27789,N_20816,N_20140);
nor U27790 (N_27790,N_20779,N_21745);
and U27791 (N_27791,N_21458,N_22807);
nor U27792 (N_27792,N_22631,N_22821);
xnor U27793 (N_27793,N_24022,N_20853);
or U27794 (N_27794,N_21668,N_20148);
nor U27795 (N_27795,N_24199,N_22689);
nand U27796 (N_27796,N_22393,N_20628);
and U27797 (N_27797,N_24114,N_20021);
or U27798 (N_27798,N_23665,N_20113);
xor U27799 (N_27799,N_22697,N_24165);
nand U27800 (N_27800,N_22368,N_21069);
or U27801 (N_27801,N_24994,N_23556);
nand U27802 (N_27802,N_21016,N_21720);
or U27803 (N_27803,N_21963,N_24448);
and U27804 (N_27804,N_23159,N_20511);
or U27805 (N_27805,N_24107,N_24414);
and U27806 (N_27806,N_22098,N_23950);
nor U27807 (N_27807,N_24892,N_20051);
or U27808 (N_27808,N_20029,N_23448);
and U27809 (N_27809,N_22238,N_22094);
or U27810 (N_27810,N_21235,N_23784);
xnor U27811 (N_27811,N_23156,N_23388);
xnor U27812 (N_27812,N_24003,N_21829);
xnor U27813 (N_27813,N_21506,N_24979);
xnor U27814 (N_27814,N_24345,N_23498);
xor U27815 (N_27815,N_20516,N_23721);
or U27816 (N_27816,N_20249,N_21306);
nand U27817 (N_27817,N_23954,N_23199);
xnor U27818 (N_27818,N_21750,N_24907);
and U27819 (N_27819,N_20870,N_23239);
and U27820 (N_27820,N_21545,N_23999);
nor U27821 (N_27821,N_22096,N_21467);
and U27822 (N_27822,N_24411,N_22709);
xnor U27823 (N_27823,N_20918,N_22948);
or U27824 (N_27824,N_20138,N_24642);
xor U27825 (N_27825,N_24820,N_22004);
nand U27826 (N_27826,N_22975,N_24416);
xnor U27827 (N_27827,N_22959,N_20888);
and U27828 (N_27828,N_20102,N_24576);
or U27829 (N_27829,N_23377,N_23762);
nand U27830 (N_27830,N_24683,N_22670);
and U27831 (N_27831,N_24148,N_21311);
nand U27832 (N_27832,N_24836,N_20542);
or U27833 (N_27833,N_24881,N_24318);
xor U27834 (N_27834,N_20715,N_21594);
nand U27835 (N_27835,N_22236,N_20287);
or U27836 (N_27836,N_21430,N_23899);
nor U27837 (N_27837,N_21140,N_24962);
xnor U27838 (N_27838,N_21833,N_22729);
or U27839 (N_27839,N_22138,N_22190);
nor U27840 (N_27840,N_20688,N_21290);
xor U27841 (N_27841,N_24073,N_22894);
or U27842 (N_27842,N_21045,N_23390);
nor U27843 (N_27843,N_22216,N_20607);
or U27844 (N_27844,N_24065,N_22587);
or U27845 (N_27845,N_21575,N_21358);
and U27846 (N_27846,N_24223,N_21183);
and U27847 (N_27847,N_24715,N_21863);
or U27848 (N_27848,N_20868,N_24898);
nand U27849 (N_27849,N_20380,N_22176);
xnor U27850 (N_27850,N_23190,N_20278);
or U27851 (N_27851,N_22293,N_22692);
and U27852 (N_27852,N_24353,N_23788);
nor U27853 (N_27853,N_22498,N_21445);
nand U27854 (N_27854,N_22024,N_22918);
xnor U27855 (N_27855,N_23105,N_20996);
and U27856 (N_27856,N_24361,N_21369);
and U27857 (N_27857,N_23300,N_20461);
xnor U27858 (N_27858,N_24303,N_22187);
nand U27859 (N_27859,N_20763,N_24874);
nand U27860 (N_27860,N_20093,N_21539);
nand U27861 (N_27861,N_21390,N_20061);
and U27862 (N_27862,N_24183,N_24230);
nor U27863 (N_27863,N_20632,N_22171);
and U27864 (N_27864,N_23553,N_22013);
and U27865 (N_27865,N_24706,N_23118);
nor U27866 (N_27866,N_24349,N_24828);
xor U27867 (N_27867,N_23656,N_23408);
nand U27868 (N_27868,N_21687,N_20577);
xnor U27869 (N_27869,N_22768,N_24565);
and U27870 (N_27870,N_24470,N_22404);
nand U27871 (N_27871,N_20805,N_22179);
nand U27872 (N_27872,N_24714,N_23263);
xor U27873 (N_27873,N_20859,N_21190);
xnor U27874 (N_27874,N_24134,N_21155);
xor U27875 (N_27875,N_23288,N_23141);
nor U27876 (N_27876,N_20724,N_23183);
or U27877 (N_27877,N_23985,N_23068);
nor U27878 (N_27878,N_20493,N_22826);
xnor U27879 (N_27879,N_23749,N_21147);
xor U27880 (N_27880,N_23640,N_24287);
nor U27881 (N_27881,N_21259,N_21216);
nand U27882 (N_27882,N_22782,N_20412);
and U27883 (N_27883,N_24522,N_21660);
nor U27884 (N_27884,N_20505,N_21170);
and U27885 (N_27885,N_21739,N_22672);
xnor U27886 (N_27886,N_24494,N_24740);
and U27887 (N_27887,N_22393,N_20236);
and U27888 (N_27888,N_24640,N_24094);
xor U27889 (N_27889,N_20516,N_20870);
or U27890 (N_27890,N_21527,N_21495);
or U27891 (N_27891,N_23792,N_22648);
xor U27892 (N_27892,N_22478,N_23948);
nor U27893 (N_27893,N_20434,N_21105);
nand U27894 (N_27894,N_21611,N_20120);
nand U27895 (N_27895,N_24454,N_21688);
nor U27896 (N_27896,N_21941,N_24657);
or U27897 (N_27897,N_22132,N_24044);
and U27898 (N_27898,N_22039,N_24048);
xnor U27899 (N_27899,N_20487,N_23031);
nor U27900 (N_27900,N_20032,N_21929);
xnor U27901 (N_27901,N_23108,N_22441);
nor U27902 (N_27902,N_21493,N_24926);
nor U27903 (N_27903,N_23919,N_23365);
xnor U27904 (N_27904,N_20969,N_22935);
nor U27905 (N_27905,N_23411,N_20616);
nand U27906 (N_27906,N_22536,N_21732);
xor U27907 (N_27907,N_24935,N_20700);
xor U27908 (N_27908,N_23929,N_23022);
nor U27909 (N_27909,N_23198,N_20526);
xnor U27910 (N_27910,N_20771,N_20645);
nand U27911 (N_27911,N_21984,N_21907);
and U27912 (N_27912,N_24400,N_23225);
or U27913 (N_27913,N_23654,N_24151);
or U27914 (N_27914,N_24146,N_21466);
and U27915 (N_27915,N_21513,N_20704);
xor U27916 (N_27916,N_24382,N_21483);
or U27917 (N_27917,N_21507,N_23117);
nand U27918 (N_27918,N_22006,N_23781);
nand U27919 (N_27919,N_23225,N_23180);
or U27920 (N_27920,N_23291,N_24247);
nor U27921 (N_27921,N_23545,N_22218);
or U27922 (N_27922,N_20173,N_20123);
nor U27923 (N_27923,N_21385,N_24638);
nand U27924 (N_27924,N_20742,N_23209);
xnor U27925 (N_27925,N_23532,N_22841);
and U27926 (N_27926,N_22637,N_22514);
or U27927 (N_27927,N_22418,N_24528);
xnor U27928 (N_27928,N_22597,N_22063);
and U27929 (N_27929,N_24730,N_20046);
and U27930 (N_27930,N_24985,N_24184);
and U27931 (N_27931,N_22748,N_22701);
nand U27932 (N_27932,N_24238,N_22586);
or U27933 (N_27933,N_24602,N_23669);
and U27934 (N_27934,N_24558,N_20066);
xnor U27935 (N_27935,N_22847,N_23157);
nor U27936 (N_27936,N_24575,N_20624);
nor U27937 (N_27937,N_23512,N_24288);
and U27938 (N_27938,N_20181,N_21680);
and U27939 (N_27939,N_23920,N_24372);
or U27940 (N_27940,N_21673,N_22523);
and U27941 (N_27941,N_23722,N_21622);
nor U27942 (N_27942,N_22091,N_21169);
and U27943 (N_27943,N_23038,N_23352);
and U27944 (N_27944,N_20063,N_22374);
and U27945 (N_27945,N_21977,N_22218);
nor U27946 (N_27946,N_21926,N_23576);
nand U27947 (N_27947,N_21144,N_24688);
and U27948 (N_27948,N_21319,N_20542);
and U27949 (N_27949,N_21006,N_20533);
nand U27950 (N_27950,N_22998,N_22152);
xnor U27951 (N_27951,N_24723,N_24638);
nand U27952 (N_27952,N_23933,N_24016);
nor U27953 (N_27953,N_20884,N_24555);
xor U27954 (N_27954,N_20107,N_22647);
nor U27955 (N_27955,N_21426,N_24371);
xnor U27956 (N_27956,N_22710,N_21335);
or U27957 (N_27957,N_24728,N_20547);
nor U27958 (N_27958,N_22785,N_20869);
or U27959 (N_27959,N_24354,N_23245);
nand U27960 (N_27960,N_22229,N_21543);
xnor U27961 (N_27961,N_22853,N_22939);
xnor U27962 (N_27962,N_24284,N_20842);
nand U27963 (N_27963,N_20825,N_20156);
xor U27964 (N_27964,N_24052,N_20598);
nand U27965 (N_27965,N_24021,N_20278);
nor U27966 (N_27966,N_21183,N_22881);
nand U27967 (N_27967,N_21985,N_21530);
or U27968 (N_27968,N_22392,N_22805);
nand U27969 (N_27969,N_24489,N_23487);
nand U27970 (N_27970,N_24805,N_24182);
nand U27971 (N_27971,N_21892,N_23070);
nor U27972 (N_27972,N_23126,N_21197);
nor U27973 (N_27973,N_21921,N_24688);
nand U27974 (N_27974,N_21195,N_22695);
and U27975 (N_27975,N_22262,N_22025);
nand U27976 (N_27976,N_23744,N_20408);
and U27977 (N_27977,N_23119,N_22585);
nor U27978 (N_27978,N_23486,N_22414);
nor U27979 (N_27979,N_22042,N_22149);
and U27980 (N_27980,N_24390,N_21220);
nand U27981 (N_27981,N_20377,N_21729);
xor U27982 (N_27982,N_22362,N_22745);
nor U27983 (N_27983,N_23130,N_20470);
or U27984 (N_27984,N_24271,N_21896);
and U27985 (N_27985,N_23514,N_21233);
and U27986 (N_27986,N_21322,N_23932);
nand U27987 (N_27987,N_23158,N_21589);
or U27988 (N_27988,N_20244,N_23720);
xor U27989 (N_27989,N_24908,N_20403);
or U27990 (N_27990,N_21179,N_22649);
nand U27991 (N_27991,N_24864,N_20967);
nor U27992 (N_27992,N_21813,N_20377);
or U27993 (N_27993,N_22722,N_23440);
xnor U27994 (N_27994,N_21205,N_24630);
or U27995 (N_27995,N_24524,N_23182);
nor U27996 (N_27996,N_23450,N_22431);
nor U27997 (N_27997,N_22800,N_22012);
xor U27998 (N_27998,N_23321,N_21886);
nand U27999 (N_27999,N_22764,N_21347);
nor U28000 (N_28000,N_21381,N_24685);
and U28001 (N_28001,N_24841,N_22126);
nor U28002 (N_28002,N_24454,N_22314);
and U28003 (N_28003,N_23553,N_22760);
nor U28004 (N_28004,N_22673,N_24973);
nand U28005 (N_28005,N_24631,N_22126);
nor U28006 (N_28006,N_21580,N_22808);
and U28007 (N_28007,N_22182,N_23128);
xnor U28008 (N_28008,N_21067,N_20740);
and U28009 (N_28009,N_23200,N_20547);
and U28010 (N_28010,N_21068,N_24130);
nor U28011 (N_28011,N_22040,N_24891);
nand U28012 (N_28012,N_21848,N_23311);
nor U28013 (N_28013,N_22934,N_23174);
nand U28014 (N_28014,N_24806,N_22362);
nand U28015 (N_28015,N_24750,N_23598);
or U28016 (N_28016,N_23013,N_20746);
nor U28017 (N_28017,N_22015,N_24014);
xnor U28018 (N_28018,N_22448,N_21865);
and U28019 (N_28019,N_21248,N_20562);
and U28020 (N_28020,N_24817,N_24694);
nor U28021 (N_28021,N_23484,N_20872);
nor U28022 (N_28022,N_20082,N_24184);
nand U28023 (N_28023,N_21845,N_23503);
xnor U28024 (N_28024,N_20835,N_22749);
xnor U28025 (N_28025,N_21749,N_20066);
nand U28026 (N_28026,N_23166,N_21498);
xnor U28027 (N_28027,N_24871,N_21916);
xor U28028 (N_28028,N_22862,N_21785);
or U28029 (N_28029,N_21553,N_21229);
xor U28030 (N_28030,N_21872,N_22532);
nor U28031 (N_28031,N_24911,N_24148);
and U28032 (N_28032,N_24368,N_23422);
or U28033 (N_28033,N_22573,N_21618);
nor U28034 (N_28034,N_20051,N_21811);
nor U28035 (N_28035,N_21315,N_24919);
xor U28036 (N_28036,N_24520,N_21583);
nor U28037 (N_28037,N_23415,N_22556);
nor U28038 (N_28038,N_21511,N_24952);
or U28039 (N_28039,N_22448,N_20589);
nand U28040 (N_28040,N_21158,N_20005);
xnor U28041 (N_28041,N_24532,N_20700);
nand U28042 (N_28042,N_24610,N_23220);
or U28043 (N_28043,N_24151,N_22598);
and U28044 (N_28044,N_21411,N_21914);
nor U28045 (N_28045,N_20000,N_24046);
or U28046 (N_28046,N_24414,N_23275);
xor U28047 (N_28047,N_20173,N_20691);
and U28048 (N_28048,N_21291,N_24182);
and U28049 (N_28049,N_24431,N_20150);
xor U28050 (N_28050,N_24160,N_23833);
and U28051 (N_28051,N_22940,N_24193);
nand U28052 (N_28052,N_24366,N_22058);
nor U28053 (N_28053,N_21412,N_21084);
nand U28054 (N_28054,N_22789,N_20328);
or U28055 (N_28055,N_22970,N_22457);
nor U28056 (N_28056,N_22867,N_23089);
and U28057 (N_28057,N_23250,N_23134);
nor U28058 (N_28058,N_21459,N_23506);
nor U28059 (N_28059,N_22759,N_24062);
nor U28060 (N_28060,N_22869,N_23729);
or U28061 (N_28061,N_23489,N_23056);
or U28062 (N_28062,N_24813,N_22546);
nor U28063 (N_28063,N_21295,N_22787);
nor U28064 (N_28064,N_24685,N_24125);
xor U28065 (N_28065,N_22226,N_24618);
or U28066 (N_28066,N_20093,N_24737);
and U28067 (N_28067,N_24005,N_20672);
nor U28068 (N_28068,N_22200,N_21604);
nor U28069 (N_28069,N_23228,N_24089);
and U28070 (N_28070,N_24306,N_20704);
nand U28071 (N_28071,N_24169,N_21835);
nand U28072 (N_28072,N_24548,N_24842);
and U28073 (N_28073,N_20936,N_24397);
nor U28074 (N_28074,N_22828,N_23268);
nor U28075 (N_28075,N_22869,N_23870);
xnor U28076 (N_28076,N_20513,N_23731);
and U28077 (N_28077,N_22244,N_24424);
nand U28078 (N_28078,N_20030,N_21178);
or U28079 (N_28079,N_23157,N_24317);
xnor U28080 (N_28080,N_20457,N_24908);
xnor U28081 (N_28081,N_24815,N_20517);
or U28082 (N_28082,N_24789,N_24031);
and U28083 (N_28083,N_23497,N_23424);
nor U28084 (N_28084,N_22059,N_23538);
xnor U28085 (N_28085,N_22507,N_21562);
or U28086 (N_28086,N_22435,N_24017);
xnor U28087 (N_28087,N_21638,N_21271);
xnor U28088 (N_28088,N_21858,N_24719);
and U28089 (N_28089,N_24088,N_22229);
and U28090 (N_28090,N_21974,N_23735);
or U28091 (N_28091,N_20749,N_23459);
xor U28092 (N_28092,N_23705,N_20924);
or U28093 (N_28093,N_21854,N_22544);
xor U28094 (N_28094,N_24456,N_24320);
xor U28095 (N_28095,N_21500,N_23145);
and U28096 (N_28096,N_22314,N_22906);
nor U28097 (N_28097,N_23031,N_22280);
xnor U28098 (N_28098,N_20369,N_23735);
nand U28099 (N_28099,N_20528,N_22568);
nor U28100 (N_28100,N_24197,N_24107);
nor U28101 (N_28101,N_20255,N_22209);
and U28102 (N_28102,N_22571,N_23076);
xnor U28103 (N_28103,N_23737,N_22435);
or U28104 (N_28104,N_23433,N_21600);
and U28105 (N_28105,N_21376,N_21771);
nor U28106 (N_28106,N_21648,N_23580);
nand U28107 (N_28107,N_23004,N_20007);
and U28108 (N_28108,N_23510,N_23052);
nor U28109 (N_28109,N_20197,N_21801);
or U28110 (N_28110,N_22622,N_20817);
or U28111 (N_28111,N_23693,N_20076);
and U28112 (N_28112,N_21081,N_24468);
xnor U28113 (N_28113,N_20424,N_23784);
nand U28114 (N_28114,N_22311,N_23521);
nor U28115 (N_28115,N_23796,N_21022);
and U28116 (N_28116,N_23353,N_23688);
nor U28117 (N_28117,N_20271,N_22484);
and U28118 (N_28118,N_20671,N_21275);
xnor U28119 (N_28119,N_23931,N_23831);
nand U28120 (N_28120,N_23900,N_21966);
nor U28121 (N_28121,N_23309,N_22980);
xor U28122 (N_28122,N_22551,N_24722);
and U28123 (N_28123,N_22266,N_21697);
xor U28124 (N_28124,N_22285,N_21579);
or U28125 (N_28125,N_24323,N_22067);
nor U28126 (N_28126,N_22189,N_20094);
nor U28127 (N_28127,N_23334,N_23798);
xor U28128 (N_28128,N_24267,N_21016);
and U28129 (N_28129,N_23329,N_24374);
xnor U28130 (N_28130,N_24220,N_24685);
and U28131 (N_28131,N_21323,N_23114);
nand U28132 (N_28132,N_22978,N_22833);
and U28133 (N_28133,N_20364,N_23685);
or U28134 (N_28134,N_21039,N_24248);
xnor U28135 (N_28135,N_22936,N_21283);
or U28136 (N_28136,N_21626,N_21938);
xnor U28137 (N_28137,N_24151,N_22421);
or U28138 (N_28138,N_22631,N_20598);
xor U28139 (N_28139,N_24639,N_21284);
and U28140 (N_28140,N_23772,N_21137);
or U28141 (N_28141,N_23003,N_20378);
nand U28142 (N_28142,N_20433,N_23625);
or U28143 (N_28143,N_24409,N_20960);
nor U28144 (N_28144,N_20626,N_23892);
and U28145 (N_28145,N_22348,N_21063);
or U28146 (N_28146,N_20627,N_23099);
xnor U28147 (N_28147,N_20738,N_24014);
xnor U28148 (N_28148,N_22637,N_21085);
nor U28149 (N_28149,N_22016,N_21319);
xor U28150 (N_28150,N_22472,N_24998);
nor U28151 (N_28151,N_22101,N_21384);
or U28152 (N_28152,N_24090,N_23701);
or U28153 (N_28153,N_24657,N_21552);
nand U28154 (N_28154,N_21951,N_23658);
or U28155 (N_28155,N_23259,N_21168);
and U28156 (N_28156,N_24434,N_21222);
nand U28157 (N_28157,N_20382,N_21406);
or U28158 (N_28158,N_23366,N_23291);
nor U28159 (N_28159,N_20988,N_20703);
or U28160 (N_28160,N_24956,N_23931);
nand U28161 (N_28161,N_20551,N_20948);
xnor U28162 (N_28162,N_21124,N_21582);
nand U28163 (N_28163,N_22705,N_24647);
xnor U28164 (N_28164,N_23252,N_22904);
or U28165 (N_28165,N_21051,N_20903);
nand U28166 (N_28166,N_24152,N_22962);
or U28167 (N_28167,N_20600,N_22912);
nand U28168 (N_28168,N_24244,N_21723);
and U28169 (N_28169,N_23192,N_23354);
xnor U28170 (N_28170,N_22223,N_20088);
xnor U28171 (N_28171,N_21055,N_23897);
nand U28172 (N_28172,N_20025,N_22356);
or U28173 (N_28173,N_24085,N_24914);
xor U28174 (N_28174,N_20180,N_20554);
and U28175 (N_28175,N_21485,N_21162);
nand U28176 (N_28176,N_20079,N_22185);
xnor U28177 (N_28177,N_23608,N_23140);
xor U28178 (N_28178,N_22418,N_23263);
nand U28179 (N_28179,N_24724,N_24526);
and U28180 (N_28180,N_23648,N_21413);
nor U28181 (N_28181,N_22592,N_21391);
and U28182 (N_28182,N_24069,N_23038);
xnor U28183 (N_28183,N_20877,N_23299);
and U28184 (N_28184,N_21861,N_20037);
or U28185 (N_28185,N_21054,N_21756);
nand U28186 (N_28186,N_23891,N_22313);
nor U28187 (N_28187,N_24767,N_22965);
or U28188 (N_28188,N_22420,N_21829);
nand U28189 (N_28189,N_24860,N_21599);
xnor U28190 (N_28190,N_23196,N_21701);
and U28191 (N_28191,N_22293,N_24094);
or U28192 (N_28192,N_20121,N_22775);
or U28193 (N_28193,N_21706,N_21283);
nand U28194 (N_28194,N_24633,N_22981);
or U28195 (N_28195,N_20290,N_20118);
nor U28196 (N_28196,N_23667,N_24354);
and U28197 (N_28197,N_23996,N_21444);
or U28198 (N_28198,N_20415,N_20549);
or U28199 (N_28199,N_24480,N_22350);
xnor U28200 (N_28200,N_20599,N_22797);
and U28201 (N_28201,N_20382,N_24653);
nand U28202 (N_28202,N_24552,N_20553);
nand U28203 (N_28203,N_23215,N_20781);
and U28204 (N_28204,N_22010,N_21839);
nor U28205 (N_28205,N_22658,N_22070);
and U28206 (N_28206,N_21292,N_20608);
or U28207 (N_28207,N_22125,N_21786);
nor U28208 (N_28208,N_20506,N_24341);
nand U28209 (N_28209,N_20063,N_20795);
or U28210 (N_28210,N_21644,N_22251);
xnor U28211 (N_28211,N_24437,N_20643);
and U28212 (N_28212,N_21706,N_23119);
xnor U28213 (N_28213,N_24806,N_24889);
nand U28214 (N_28214,N_22819,N_23421);
nand U28215 (N_28215,N_22007,N_21546);
nor U28216 (N_28216,N_23418,N_24703);
and U28217 (N_28217,N_21888,N_21442);
and U28218 (N_28218,N_20953,N_24961);
or U28219 (N_28219,N_24204,N_20776);
or U28220 (N_28220,N_20365,N_23369);
nand U28221 (N_28221,N_21615,N_20630);
nor U28222 (N_28222,N_24485,N_24701);
or U28223 (N_28223,N_21837,N_22826);
nor U28224 (N_28224,N_20176,N_23816);
nor U28225 (N_28225,N_23550,N_22578);
or U28226 (N_28226,N_20323,N_21808);
xor U28227 (N_28227,N_24884,N_24472);
nor U28228 (N_28228,N_22662,N_23565);
and U28229 (N_28229,N_24363,N_23587);
or U28230 (N_28230,N_23401,N_24487);
nor U28231 (N_28231,N_20533,N_20826);
nand U28232 (N_28232,N_23835,N_22020);
nand U28233 (N_28233,N_21018,N_24211);
and U28234 (N_28234,N_21609,N_21256);
nand U28235 (N_28235,N_23027,N_23239);
nand U28236 (N_28236,N_21813,N_24546);
nor U28237 (N_28237,N_22651,N_20015);
and U28238 (N_28238,N_21314,N_24652);
xor U28239 (N_28239,N_22756,N_23241);
nor U28240 (N_28240,N_23921,N_22673);
nand U28241 (N_28241,N_21851,N_22883);
nor U28242 (N_28242,N_23741,N_22548);
xor U28243 (N_28243,N_20096,N_22131);
nor U28244 (N_28244,N_21355,N_23282);
and U28245 (N_28245,N_23572,N_21539);
nand U28246 (N_28246,N_23537,N_20015);
xor U28247 (N_28247,N_24445,N_22899);
xor U28248 (N_28248,N_20839,N_20442);
xnor U28249 (N_28249,N_24183,N_24261);
or U28250 (N_28250,N_24519,N_23986);
nor U28251 (N_28251,N_22042,N_24197);
xnor U28252 (N_28252,N_21005,N_22852);
xnor U28253 (N_28253,N_23200,N_23609);
nand U28254 (N_28254,N_22956,N_20257);
nand U28255 (N_28255,N_20217,N_24710);
xor U28256 (N_28256,N_23252,N_22068);
or U28257 (N_28257,N_21359,N_23465);
and U28258 (N_28258,N_24825,N_23928);
xor U28259 (N_28259,N_24886,N_24411);
nand U28260 (N_28260,N_21212,N_20855);
xor U28261 (N_28261,N_23297,N_20729);
and U28262 (N_28262,N_20774,N_23502);
and U28263 (N_28263,N_23041,N_21933);
and U28264 (N_28264,N_20109,N_24523);
or U28265 (N_28265,N_20801,N_23392);
nand U28266 (N_28266,N_21517,N_22175);
and U28267 (N_28267,N_23752,N_23931);
nor U28268 (N_28268,N_24947,N_23918);
nand U28269 (N_28269,N_20033,N_20182);
and U28270 (N_28270,N_20894,N_24977);
and U28271 (N_28271,N_24073,N_24555);
nand U28272 (N_28272,N_22589,N_22094);
or U28273 (N_28273,N_22825,N_22583);
nor U28274 (N_28274,N_21404,N_23625);
and U28275 (N_28275,N_22576,N_21609);
xnor U28276 (N_28276,N_20463,N_24528);
nor U28277 (N_28277,N_21903,N_23773);
xnor U28278 (N_28278,N_21044,N_22679);
or U28279 (N_28279,N_22859,N_20697);
or U28280 (N_28280,N_22343,N_21118);
or U28281 (N_28281,N_23050,N_23600);
or U28282 (N_28282,N_24577,N_22336);
or U28283 (N_28283,N_24560,N_21440);
xnor U28284 (N_28284,N_20705,N_21066);
or U28285 (N_28285,N_22743,N_24140);
nor U28286 (N_28286,N_23881,N_21736);
nor U28287 (N_28287,N_21696,N_20272);
xnor U28288 (N_28288,N_20922,N_21400);
nor U28289 (N_28289,N_21215,N_24478);
or U28290 (N_28290,N_20240,N_21768);
nor U28291 (N_28291,N_23918,N_21851);
and U28292 (N_28292,N_23557,N_24313);
nand U28293 (N_28293,N_20168,N_21263);
and U28294 (N_28294,N_21562,N_20144);
xnor U28295 (N_28295,N_22931,N_22627);
xnor U28296 (N_28296,N_23990,N_22571);
nand U28297 (N_28297,N_22479,N_24370);
nand U28298 (N_28298,N_21744,N_21292);
nand U28299 (N_28299,N_20111,N_24362);
nand U28300 (N_28300,N_23301,N_24158);
xnor U28301 (N_28301,N_24140,N_21052);
nand U28302 (N_28302,N_20829,N_23531);
or U28303 (N_28303,N_21809,N_21664);
and U28304 (N_28304,N_22276,N_23907);
nor U28305 (N_28305,N_23785,N_20300);
or U28306 (N_28306,N_20323,N_23122);
nand U28307 (N_28307,N_23133,N_23403);
xor U28308 (N_28308,N_24788,N_23507);
nand U28309 (N_28309,N_20676,N_22163);
or U28310 (N_28310,N_21519,N_24856);
xnor U28311 (N_28311,N_20160,N_22033);
and U28312 (N_28312,N_22509,N_22499);
xor U28313 (N_28313,N_20357,N_22267);
nor U28314 (N_28314,N_20386,N_23611);
nand U28315 (N_28315,N_20082,N_20498);
xnor U28316 (N_28316,N_24907,N_23441);
xor U28317 (N_28317,N_21158,N_20634);
xor U28318 (N_28318,N_24727,N_22500);
and U28319 (N_28319,N_20009,N_21001);
nor U28320 (N_28320,N_23452,N_22395);
or U28321 (N_28321,N_21383,N_24473);
nand U28322 (N_28322,N_21729,N_20507);
xor U28323 (N_28323,N_22965,N_20708);
or U28324 (N_28324,N_23867,N_23182);
and U28325 (N_28325,N_20431,N_22077);
xor U28326 (N_28326,N_24398,N_22954);
or U28327 (N_28327,N_20341,N_23108);
xor U28328 (N_28328,N_23103,N_23022);
nor U28329 (N_28329,N_20187,N_20396);
xor U28330 (N_28330,N_20609,N_20369);
nand U28331 (N_28331,N_22794,N_22610);
nand U28332 (N_28332,N_20601,N_23277);
nand U28333 (N_28333,N_22345,N_20742);
nor U28334 (N_28334,N_22244,N_24822);
nand U28335 (N_28335,N_23195,N_24353);
xnor U28336 (N_28336,N_22641,N_24710);
and U28337 (N_28337,N_20903,N_23917);
and U28338 (N_28338,N_23942,N_20377);
and U28339 (N_28339,N_23069,N_21931);
and U28340 (N_28340,N_21969,N_23208);
xnor U28341 (N_28341,N_22923,N_23685);
or U28342 (N_28342,N_24275,N_24736);
or U28343 (N_28343,N_24264,N_22602);
nand U28344 (N_28344,N_24210,N_20380);
nand U28345 (N_28345,N_24820,N_21190);
nor U28346 (N_28346,N_23857,N_22105);
xnor U28347 (N_28347,N_21455,N_23374);
xnor U28348 (N_28348,N_20358,N_23384);
or U28349 (N_28349,N_21170,N_23778);
or U28350 (N_28350,N_23270,N_24116);
or U28351 (N_28351,N_20728,N_24838);
and U28352 (N_28352,N_23943,N_22707);
and U28353 (N_28353,N_23777,N_24570);
and U28354 (N_28354,N_22221,N_24581);
and U28355 (N_28355,N_24019,N_22261);
and U28356 (N_28356,N_24888,N_22132);
nand U28357 (N_28357,N_22282,N_23784);
nand U28358 (N_28358,N_23857,N_23961);
or U28359 (N_28359,N_22739,N_21958);
nand U28360 (N_28360,N_24174,N_21790);
or U28361 (N_28361,N_24339,N_24454);
nand U28362 (N_28362,N_24759,N_21807);
and U28363 (N_28363,N_21257,N_23225);
xnor U28364 (N_28364,N_24331,N_24302);
xor U28365 (N_28365,N_22920,N_24437);
nor U28366 (N_28366,N_21876,N_22706);
nand U28367 (N_28367,N_22282,N_22840);
xor U28368 (N_28368,N_21746,N_20316);
or U28369 (N_28369,N_20031,N_24519);
xnor U28370 (N_28370,N_24941,N_20904);
nor U28371 (N_28371,N_20446,N_24493);
and U28372 (N_28372,N_20695,N_22747);
nand U28373 (N_28373,N_24375,N_20740);
xnor U28374 (N_28374,N_20947,N_24523);
xor U28375 (N_28375,N_20746,N_24669);
xnor U28376 (N_28376,N_24986,N_20233);
xor U28377 (N_28377,N_22277,N_23643);
and U28378 (N_28378,N_21488,N_22169);
or U28379 (N_28379,N_23492,N_21730);
or U28380 (N_28380,N_22779,N_24249);
nor U28381 (N_28381,N_20123,N_22606);
and U28382 (N_28382,N_21107,N_24342);
nor U28383 (N_28383,N_22085,N_23390);
xnor U28384 (N_28384,N_20675,N_21268);
nor U28385 (N_28385,N_21181,N_24648);
or U28386 (N_28386,N_21666,N_20696);
nand U28387 (N_28387,N_24809,N_24908);
xor U28388 (N_28388,N_21301,N_24293);
and U28389 (N_28389,N_24289,N_20309);
nand U28390 (N_28390,N_22361,N_23333);
xor U28391 (N_28391,N_21788,N_22900);
and U28392 (N_28392,N_22064,N_21590);
or U28393 (N_28393,N_20620,N_21074);
nor U28394 (N_28394,N_22624,N_21264);
or U28395 (N_28395,N_21078,N_22631);
xnor U28396 (N_28396,N_24032,N_23683);
nand U28397 (N_28397,N_24602,N_22192);
nor U28398 (N_28398,N_22860,N_21822);
nand U28399 (N_28399,N_22369,N_20065);
nand U28400 (N_28400,N_21975,N_24661);
nor U28401 (N_28401,N_22638,N_23270);
or U28402 (N_28402,N_20947,N_20702);
xor U28403 (N_28403,N_20348,N_21388);
nand U28404 (N_28404,N_20042,N_22629);
and U28405 (N_28405,N_24341,N_24734);
or U28406 (N_28406,N_20089,N_23774);
or U28407 (N_28407,N_20374,N_20475);
xnor U28408 (N_28408,N_21068,N_22468);
nor U28409 (N_28409,N_22194,N_24755);
and U28410 (N_28410,N_24000,N_21953);
or U28411 (N_28411,N_23531,N_22635);
and U28412 (N_28412,N_23663,N_21140);
nand U28413 (N_28413,N_24244,N_20018);
or U28414 (N_28414,N_24130,N_24221);
nand U28415 (N_28415,N_23257,N_20696);
nand U28416 (N_28416,N_21016,N_20265);
and U28417 (N_28417,N_22079,N_20019);
nor U28418 (N_28418,N_21375,N_20887);
nor U28419 (N_28419,N_21003,N_24731);
nand U28420 (N_28420,N_21740,N_24234);
or U28421 (N_28421,N_20683,N_20065);
xor U28422 (N_28422,N_20284,N_24391);
nor U28423 (N_28423,N_21735,N_20357);
xnor U28424 (N_28424,N_20600,N_22683);
nand U28425 (N_28425,N_23333,N_23919);
and U28426 (N_28426,N_24600,N_24777);
or U28427 (N_28427,N_24383,N_23097);
and U28428 (N_28428,N_23843,N_22758);
or U28429 (N_28429,N_23306,N_20503);
xnor U28430 (N_28430,N_22304,N_23277);
nand U28431 (N_28431,N_21342,N_20747);
and U28432 (N_28432,N_21942,N_22214);
or U28433 (N_28433,N_22985,N_21448);
and U28434 (N_28434,N_21623,N_21162);
and U28435 (N_28435,N_23024,N_22376);
and U28436 (N_28436,N_21935,N_23442);
nand U28437 (N_28437,N_23174,N_21619);
xnor U28438 (N_28438,N_23044,N_24474);
or U28439 (N_28439,N_22753,N_22945);
nand U28440 (N_28440,N_24450,N_23883);
or U28441 (N_28441,N_20190,N_20865);
and U28442 (N_28442,N_21677,N_22307);
and U28443 (N_28443,N_22413,N_22459);
nand U28444 (N_28444,N_23628,N_21638);
nor U28445 (N_28445,N_20625,N_22201);
or U28446 (N_28446,N_22139,N_22172);
or U28447 (N_28447,N_24171,N_22932);
xor U28448 (N_28448,N_24100,N_22383);
and U28449 (N_28449,N_21130,N_23137);
and U28450 (N_28450,N_21306,N_20253);
nor U28451 (N_28451,N_22496,N_20027);
and U28452 (N_28452,N_23827,N_24041);
nor U28453 (N_28453,N_22272,N_21148);
xor U28454 (N_28454,N_22195,N_23358);
or U28455 (N_28455,N_21642,N_20940);
and U28456 (N_28456,N_24050,N_20666);
nor U28457 (N_28457,N_21474,N_21321);
or U28458 (N_28458,N_21716,N_21571);
or U28459 (N_28459,N_23425,N_20716);
or U28460 (N_28460,N_23969,N_21387);
and U28461 (N_28461,N_24389,N_23107);
or U28462 (N_28462,N_23455,N_20822);
nor U28463 (N_28463,N_24583,N_22737);
or U28464 (N_28464,N_24576,N_22869);
nand U28465 (N_28465,N_21576,N_24453);
or U28466 (N_28466,N_24372,N_21429);
and U28467 (N_28467,N_24932,N_20725);
and U28468 (N_28468,N_21169,N_20943);
nor U28469 (N_28469,N_20257,N_22755);
or U28470 (N_28470,N_24493,N_23147);
nand U28471 (N_28471,N_24631,N_22640);
and U28472 (N_28472,N_21757,N_20127);
nor U28473 (N_28473,N_24073,N_20187);
nor U28474 (N_28474,N_21625,N_22669);
nand U28475 (N_28475,N_22210,N_20404);
nand U28476 (N_28476,N_20950,N_20064);
or U28477 (N_28477,N_20935,N_24979);
nand U28478 (N_28478,N_22858,N_20546);
xnor U28479 (N_28479,N_23395,N_22702);
and U28480 (N_28480,N_21173,N_22989);
xnor U28481 (N_28481,N_24779,N_24087);
and U28482 (N_28482,N_24383,N_22033);
or U28483 (N_28483,N_23940,N_21066);
nand U28484 (N_28484,N_24419,N_23672);
or U28485 (N_28485,N_22256,N_21127);
nor U28486 (N_28486,N_24553,N_21422);
nor U28487 (N_28487,N_23528,N_24947);
xor U28488 (N_28488,N_24522,N_21065);
nand U28489 (N_28489,N_22636,N_24446);
xnor U28490 (N_28490,N_22595,N_22634);
nor U28491 (N_28491,N_23400,N_24502);
nand U28492 (N_28492,N_23592,N_20194);
and U28493 (N_28493,N_20333,N_21539);
nand U28494 (N_28494,N_24009,N_20215);
or U28495 (N_28495,N_21481,N_23698);
or U28496 (N_28496,N_24346,N_22649);
and U28497 (N_28497,N_20643,N_22810);
nor U28498 (N_28498,N_23343,N_24281);
xor U28499 (N_28499,N_20340,N_22234);
and U28500 (N_28500,N_20486,N_22661);
xnor U28501 (N_28501,N_23145,N_21792);
or U28502 (N_28502,N_20029,N_21620);
or U28503 (N_28503,N_22679,N_22162);
nand U28504 (N_28504,N_20917,N_24493);
nand U28505 (N_28505,N_20753,N_23326);
xnor U28506 (N_28506,N_20327,N_24795);
or U28507 (N_28507,N_23733,N_23384);
and U28508 (N_28508,N_24880,N_23350);
nand U28509 (N_28509,N_20741,N_20589);
nand U28510 (N_28510,N_23493,N_20869);
xnor U28511 (N_28511,N_21708,N_21894);
nor U28512 (N_28512,N_22363,N_22495);
or U28513 (N_28513,N_23311,N_20485);
nand U28514 (N_28514,N_21266,N_22809);
xnor U28515 (N_28515,N_22846,N_21642);
or U28516 (N_28516,N_24190,N_24549);
or U28517 (N_28517,N_23680,N_21325);
and U28518 (N_28518,N_23942,N_24708);
or U28519 (N_28519,N_23010,N_23269);
nand U28520 (N_28520,N_24317,N_22635);
or U28521 (N_28521,N_20197,N_24035);
and U28522 (N_28522,N_23144,N_24973);
nor U28523 (N_28523,N_23919,N_22418);
and U28524 (N_28524,N_24242,N_23604);
nand U28525 (N_28525,N_20939,N_21548);
xor U28526 (N_28526,N_24108,N_24102);
nand U28527 (N_28527,N_20411,N_21000);
xnor U28528 (N_28528,N_24576,N_24675);
and U28529 (N_28529,N_22725,N_21122);
or U28530 (N_28530,N_22726,N_22261);
and U28531 (N_28531,N_20321,N_22488);
nand U28532 (N_28532,N_20697,N_21671);
nor U28533 (N_28533,N_23934,N_23573);
nor U28534 (N_28534,N_22683,N_22162);
nor U28535 (N_28535,N_20390,N_20749);
or U28536 (N_28536,N_22154,N_21025);
or U28537 (N_28537,N_22098,N_21710);
nand U28538 (N_28538,N_23319,N_22764);
nor U28539 (N_28539,N_24746,N_24157);
xor U28540 (N_28540,N_20501,N_21004);
and U28541 (N_28541,N_22609,N_21409);
nand U28542 (N_28542,N_21550,N_21054);
or U28543 (N_28543,N_22322,N_20316);
nand U28544 (N_28544,N_23425,N_21461);
nor U28545 (N_28545,N_23256,N_21756);
nor U28546 (N_28546,N_24756,N_23436);
nand U28547 (N_28547,N_21970,N_20878);
nor U28548 (N_28548,N_20864,N_23101);
nor U28549 (N_28549,N_23580,N_23687);
and U28550 (N_28550,N_22087,N_22393);
xor U28551 (N_28551,N_23714,N_20274);
xor U28552 (N_28552,N_24564,N_22028);
nor U28553 (N_28553,N_23495,N_20477);
nand U28554 (N_28554,N_22639,N_24362);
and U28555 (N_28555,N_21927,N_21500);
nor U28556 (N_28556,N_21521,N_24119);
or U28557 (N_28557,N_24868,N_20264);
nor U28558 (N_28558,N_20350,N_20679);
xor U28559 (N_28559,N_20924,N_22926);
and U28560 (N_28560,N_21045,N_21267);
nand U28561 (N_28561,N_24094,N_23695);
nand U28562 (N_28562,N_21656,N_21861);
nor U28563 (N_28563,N_20522,N_22118);
or U28564 (N_28564,N_24789,N_24589);
or U28565 (N_28565,N_24760,N_22853);
xnor U28566 (N_28566,N_22801,N_24019);
xnor U28567 (N_28567,N_21259,N_21344);
xnor U28568 (N_28568,N_24224,N_23438);
or U28569 (N_28569,N_24305,N_23898);
and U28570 (N_28570,N_24169,N_21466);
or U28571 (N_28571,N_21122,N_23889);
nand U28572 (N_28572,N_21432,N_21420);
xnor U28573 (N_28573,N_24046,N_20132);
nand U28574 (N_28574,N_23944,N_23338);
and U28575 (N_28575,N_23252,N_23916);
xor U28576 (N_28576,N_20133,N_20436);
xnor U28577 (N_28577,N_24472,N_20547);
nand U28578 (N_28578,N_20139,N_22428);
or U28579 (N_28579,N_21457,N_21510);
xor U28580 (N_28580,N_20886,N_23310);
nand U28581 (N_28581,N_22926,N_24769);
or U28582 (N_28582,N_21881,N_23032);
nand U28583 (N_28583,N_24954,N_23114);
or U28584 (N_28584,N_24611,N_21354);
or U28585 (N_28585,N_21884,N_24860);
or U28586 (N_28586,N_24388,N_22942);
or U28587 (N_28587,N_21623,N_24388);
nand U28588 (N_28588,N_24951,N_23840);
or U28589 (N_28589,N_24309,N_22401);
xor U28590 (N_28590,N_23954,N_21429);
xor U28591 (N_28591,N_23652,N_20503);
nand U28592 (N_28592,N_24105,N_23220);
nor U28593 (N_28593,N_22795,N_24051);
and U28594 (N_28594,N_23388,N_20103);
or U28595 (N_28595,N_22347,N_20806);
nand U28596 (N_28596,N_23178,N_20147);
and U28597 (N_28597,N_21945,N_24915);
xnor U28598 (N_28598,N_24472,N_20712);
and U28599 (N_28599,N_23629,N_20488);
xor U28600 (N_28600,N_21776,N_23853);
xor U28601 (N_28601,N_24628,N_24333);
and U28602 (N_28602,N_21300,N_20495);
or U28603 (N_28603,N_24091,N_22504);
xnor U28604 (N_28604,N_23450,N_22879);
and U28605 (N_28605,N_24543,N_23035);
nor U28606 (N_28606,N_22871,N_22326);
nand U28607 (N_28607,N_21503,N_23393);
nand U28608 (N_28608,N_22640,N_20022);
nor U28609 (N_28609,N_23430,N_23364);
or U28610 (N_28610,N_22768,N_22014);
xor U28611 (N_28611,N_21961,N_22107);
or U28612 (N_28612,N_20678,N_22216);
and U28613 (N_28613,N_22393,N_22691);
nor U28614 (N_28614,N_24454,N_20869);
nand U28615 (N_28615,N_20097,N_24480);
nand U28616 (N_28616,N_24093,N_23108);
nand U28617 (N_28617,N_23964,N_21947);
xnor U28618 (N_28618,N_22894,N_24592);
or U28619 (N_28619,N_22573,N_20843);
or U28620 (N_28620,N_22131,N_22996);
nor U28621 (N_28621,N_22377,N_21728);
nand U28622 (N_28622,N_24635,N_23000);
nand U28623 (N_28623,N_20513,N_23152);
or U28624 (N_28624,N_23082,N_21770);
xor U28625 (N_28625,N_20612,N_20845);
nor U28626 (N_28626,N_23793,N_22463);
nor U28627 (N_28627,N_21782,N_22980);
and U28628 (N_28628,N_24212,N_23597);
or U28629 (N_28629,N_23003,N_21733);
nand U28630 (N_28630,N_21694,N_23593);
and U28631 (N_28631,N_21365,N_20790);
and U28632 (N_28632,N_20977,N_20218);
nand U28633 (N_28633,N_24100,N_20445);
nand U28634 (N_28634,N_24261,N_21463);
xor U28635 (N_28635,N_20762,N_22346);
and U28636 (N_28636,N_22104,N_20955);
xnor U28637 (N_28637,N_21064,N_22812);
and U28638 (N_28638,N_23950,N_24927);
nor U28639 (N_28639,N_21500,N_24863);
and U28640 (N_28640,N_22133,N_24278);
nand U28641 (N_28641,N_20471,N_24823);
or U28642 (N_28642,N_24042,N_21256);
or U28643 (N_28643,N_20763,N_20018);
nor U28644 (N_28644,N_22698,N_22346);
or U28645 (N_28645,N_20010,N_24340);
or U28646 (N_28646,N_22868,N_23765);
nor U28647 (N_28647,N_20562,N_20359);
nor U28648 (N_28648,N_24247,N_24824);
nand U28649 (N_28649,N_24464,N_24195);
and U28650 (N_28650,N_20939,N_21177);
and U28651 (N_28651,N_20004,N_20929);
or U28652 (N_28652,N_24958,N_22807);
or U28653 (N_28653,N_23644,N_21494);
or U28654 (N_28654,N_20073,N_20232);
and U28655 (N_28655,N_24762,N_21860);
nor U28656 (N_28656,N_24771,N_22237);
xor U28657 (N_28657,N_21323,N_23931);
nor U28658 (N_28658,N_22788,N_21686);
nor U28659 (N_28659,N_22384,N_21162);
xnor U28660 (N_28660,N_24833,N_24174);
and U28661 (N_28661,N_21648,N_23687);
nor U28662 (N_28662,N_22856,N_21017);
xnor U28663 (N_28663,N_24005,N_23209);
and U28664 (N_28664,N_20623,N_22983);
and U28665 (N_28665,N_23239,N_22025);
or U28666 (N_28666,N_21331,N_23489);
and U28667 (N_28667,N_23364,N_22914);
xnor U28668 (N_28668,N_22869,N_22286);
or U28669 (N_28669,N_24577,N_23105);
xor U28670 (N_28670,N_24914,N_24927);
and U28671 (N_28671,N_24164,N_24028);
or U28672 (N_28672,N_23347,N_24824);
or U28673 (N_28673,N_20153,N_20170);
nor U28674 (N_28674,N_20451,N_21189);
nand U28675 (N_28675,N_24247,N_23238);
xnor U28676 (N_28676,N_24845,N_23710);
xnor U28677 (N_28677,N_20770,N_21200);
xnor U28678 (N_28678,N_22220,N_22801);
or U28679 (N_28679,N_24899,N_22558);
nor U28680 (N_28680,N_24087,N_20602);
and U28681 (N_28681,N_24495,N_22426);
nand U28682 (N_28682,N_20566,N_23350);
xnor U28683 (N_28683,N_20295,N_22160);
xnor U28684 (N_28684,N_23065,N_22361);
or U28685 (N_28685,N_22657,N_22018);
and U28686 (N_28686,N_22075,N_22942);
nor U28687 (N_28687,N_20681,N_22634);
nand U28688 (N_28688,N_22372,N_20962);
and U28689 (N_28689,N_22830,N_22463);
and U28690 (N_28690,N_21078,N_22679);
nand U28691 (N_28691,N_22205,N_23264);
or U28692 (N_28692,N_21394,N_24122);
and U28693 (N_28693,N_24712,N_23255);
xor U28694 (N_28694,N_24006,N_22811);
nand U28695 (N_28695,N_20539,N_21365);
or U28696 (N_28696,N_23865,N_20385);
and U28697 (N_28697,N_22085,N_23258);
nor U28698 (N_28698,N_22797,N_21608);
or U28699 (N_28699,N_21360,N_23387);
nor U28700 (N_28700,N_24034,N_23649);
xor U28701 (N_28701,N_22932,N_24842);
xnor U28702 (N_28702,N_24670,N_20953);
or U28703 (N_28703,N_22227,N_20704);
nor U28704 (N_28704,N_24949,N_24297);
xnor U28705 (N_28705,N_22305,N_23068);
nand U28706 (N_28706,N_24198,N_20723);
or U28707 (N_28707,N_22464,N_24600);
nor U28708 (N_28708,N_22415,N_24358);
nand U28709 (N_28709,N_23268,N_21459);
nor U28710 (N_28710,N_22372,N_20843);
or U28711 (N_28711,N_20849,N_23753);
or U28712 (N_28712,N_23198,N_24371);
nor U28713 (N_28713,N_22304,N_21443);
nor U28714 (N_28714,N_23843,N_21706);
or U28715 (N_28715,N_23497,N_22223);
nand U28716 (N_28716,N_22223,N_20868);
nor U28717 (N_28717,N_23345,N_22209);
nand U28718 (N_28718,N_24317,N_23116);
nor U28719 (N_28719,N_23722,N_24682);
and U28720 (N_28720,N_21515,N_23139);
xor U28721 (N_28721,N_22030,N_23245);
nand U28722 (N_28722,N_22910,N_21250);
and U28723 (N_28723,N_23440,N_24535);
or U28724 (N_28724,N_24013,N_20884);
nor U28725 (N_28725,N_20308,N_23102);
nand U28726 (N_28726,N_23596,N_21959);
nor U28727 (N_28727,N_23025,N_20261);
or U28728 (N_28728,N_24661,N_24395);
xnor U28729 (N_28729,N_21274,N_22614);
or U28730 (N_28730,N_23092,N_23966);
nand U28731 (N_28731,N_20271,N_21050);
nor U28732 (N_28732,N_24562,N_24629);
nand U28733 (N_28733,N_21614,N_21713);
nand U28734 (N_28734,N_21961,N_20638);
and U28735 (N_28735,N_22432,N_23045);
xor U28736 (N_28736,N_20038,N_20178);
nand U28737 (N_28737,N_24798,N_20712);
and U28738 (N_28738,N_22496,N_20699);
nor U28739 (N_28739,N_20241,N_21728);
nand U28740 (N_28740,N_24212,N_23567);
and U28741 (N_28741,N_23178,N_20512);
and U28742 (N_28742,N_23049,N_24156);
xnor U28743 (N_28743,N_22624,N_20868);
or U28744 (N_28744,N_23908,N_23915);
and U28745 (N_28745,N_24368,N_20949);
nand U28746 (N_28746,N_22153,N_23404);
nor U28747 (N_28747,N_24182,N_20996);
or U28748 (N_28748,N_20694,N_24778);
and U28749 (N_28749,N_22576,N_24065);
and U28750 (N_28750,N_21161,N_20335);
nor U28751 (N_28751,N_22040,N_22660);
xnor U28752 (N_28752,N_23765,N_24365);
nand U28753 (N_28753,N_21195,N_24321);
nand U28754 (N_28754,N_24859,N_20139);
xnor U28755 (N_28755,N_20348,N_21877);
nor U28756 (N_28756,N_22423,N_21874);
nand U28757 (N_28757,N_23891,N_23226);
xor U28758 (N_28758,N_23452,N_20480);
and U28759 (N_28759,N_24755,N_22730);
xor U28760 (N_28760,N_21029,N_24690);
nand U28761 (N_28761,N_20997,N_21569);
nor U28762 (N_28762,N_21658,N_24105);
or U28763 (N_28763,N_21246,N_23983);
xnor U28764 (N_28764,N_23274,N_21250);
nand U28765 (N_28765,N_22310,N_23698);
and U28766 (N_28766,N_22267,N_23130);
or U28767 (N_28767,N_20999,N_23339);
xor U28768 (N_28768,N_23581,N_23406);
or U28769 (N_28769,N_24644,N_24668);
and U28770 (N_28770,N_22680,N_21665);
xnor U28771 (N_28771,N_23099,N_20769);
nor U28772 (N_28772,N_23679,N_23427);
xor U28773 (N_28773,N_24509,N_22133);
nand U28774 (N_28774,N_23511,N_23903);
nand U28775 (N_28775,N_22704,N_20862);
nor U28776 (N_28776,N_23042,N_24598);
or U28777 (N_28777,N_20443,N_21915);
nand U28778 (N_28778,N_24739,N_21497);
nor U28779 (N_28779,N_24629,N_22061);
nor U28780 (N_28780,N_20060,N_22209);
and U28781 (N_28781,N_21320,N_20479);
or U28782 (N_28782,N_24276,N_23374);
nor U28783 (N_28783,N_22667,N_24544);
nand U28784 (N_28784,N_24823,N_24908);
or U28785 (N_28785,N_24961,N_22692);
or U28786 (N_28786,N_20871,N_23877);
or U28787 (N_28787,N_22530,N_20893);
nand U28788 (N_28788,N_22343,N_24076);
and U28789 (N_28789,N_22739,N_24395);
nor U28790 (N_28790,N_20982,N_22887);
nor U28791 (N_28791,N_20950,N_20063);
nand U28792 (N_28792,N_22216,N_24860);
xor U28793 (N_28793,N_22070,N_20825);
or U28794 (N_28794,N_24440,N_22040);
nand U28795 (N_28795,N_23792,N_22691);
nor U28796 (N_28796,N_23415,N_24293);
nor U28797 (N_28797,N_20975,N_20733);
nand U28798 (N_28798,N_21034,N_24397);
and U28799 (N_28799,N_24687,N_21459);
or U28800 (N_28800,N_21860,N_23119);
xnor U28801 (N_28801,N_21104,N_20049);
or U28802 (N_28802,N_21980,N_23364);
and U28803 (N_28803,N_24224,N_22872);
xnor U28804 (N_28804,N_21459,N_24464);
or U28805 (N_28805,N_20209,N_20745);
xor U28806 (N_28806,N_20129,N_22651);
or U28807 (N_28807,N_24147,N_24656);
xnor U28808 (N_28808,N_22202,N_24864);
nor U28809 (N_28809,N_20063,N_23913);
xnor U28810 (N_28810,N_23711,N_22732);
and U28811 (N_28811,N_21336,N_20948);
nor U28812 (N_28812,N_23273,N_23885);
xnor U28813 (N_28813,N_22966,N_24662);
or U28814 (N_28814,N_22122,N_23687);
or U28815 (N_28815,N_24436,N_24747);
and U28816 (N_28816,N_22976,N_21792);
nor U28817 (N_28817,N_24133,N_24174);
nand U28818 (N_28818,N_23887,N_24106);
or U28819 (N_28819,N_22075,N_24269);
nand U28820 (N_28820,N_23031,N_21813);
or U28821 (N_28821,N_20796,N_22736);
nor U28822 (N_28822,N_22746,N_20176);
xnor U28823 (N_28823,N_24844,N_20670);
nor U28824 (N_28824,N_20183,N_21220);
and U28825 (N_28825,N_23773,N_23095);
and U28826 (N_28826,N_24714,N_23590);
and U28827 (N_28827,N_20405,N_20396);
or U28828 (N_28828,N_21972,N_21313);
and U28829 (N_28829,N_22708,N_20148);
nor U28830 (N_28830,N_21978,N_21395);
xor U28831 (N_28831,N_21956,N_22347);
xor U28832 (N_28832,N_24445,N_24817);
or U28833 (N_28833,N_23342,N_21526);
xor U28834 (N_28834,N_23895,N_20338);
and U28835 (N_28835,N_23502,N_24052);
or U28836 (N_28836,N_22176,N_22545);
or U28837 (N_28837,N_24672,N_21958);
and U28838 (N_28838,N_23730,N_20949);
nand U28839 (N_28839,N_24116,N_21063);
nand U28840 (N_28840,N_24338,N_22846);
nand U28841 (N_28841,N_20117,N_24728);
nand U28842 (N_28842,N_21837,N_21645);
and U28843 (N_28843,N_24068,N_21662);
nand U28844 (N_28844,N_20947,N_21686);
and U28845 (N_28845,N_23106,N_23322);
xnor U28846 (N_28846,N_24987,N_23150);
and U28847 (N_28847,N_24010,N_22056);
xnor U28848 (N_28848,N_24275,N_20478);
nor U28849 (N_28849,N_23960,N_22854);
and U28850 (N_28850,N_20057,N_20657);
or U28851 (N_28851,N_22491,N_24467);
xnor U28852 (N_28852,N_24309,N_23788);
and U28853 (N_28853,N_24731,N_21707);
or U28854 (N_28854,N_21701,N_24550);
nand U28855 (N_28855,N_20486,N_20613);
nand U28856 (N_28856,N_20797,N_23938);
or U28857 (N_28857,N_22283,N_24834);
or U28858 (N_28858,N_21992,N_21202);
xor U28859 (N_28859,N_21509,N_24081);
xnor U28860 (N_28860,N_22473,N_20552);
and U28861 (N_28861,N_20857,N_24178);
xor U28862 (N_28862,N_21268,N_24550);
or U28863 (N_28863,N_22583,N_22843);
or U28864 (N_28864,N_22294,N_21196);
and U28865 (N_28865,N_22767,N_21685);
nor U28866 (N_28866,N_23335,N_20731);
nor U28867 (N_28867,N_20960,N_23256);
and U28868 (N_28868,N_20113,N_21965);
or U28869 (N_28869,N_21499,N_22096);
nor U28870 (N_28870,N_20484,N_20859);
nand U28871 (N_28871,N_20909,N_24273);
or U28872 (N_28872,N_22370,N_22810);
and U28873 (N_28873,N_22217,N_24888);
or U28874 (N_28874,N_22975,N_22846);
xnor U28875 (N_28875,N_24990,N_20064);
xnor U28876 (N_28876,N_22323,N_20441);
nor U28877 (N_28877,N_22662,N_24444);
or U28878 (N_28878,N_22689,N_23941);
nand U28879 (N_28879,N_23189,N_24730);
and U28880 (N_28880,N_23844,N_23842);
nand U28881 (N_28881,N_20186,N_20978);
xor U28882 (N_28882,N_20065,N_24446);
and U28883 (N_28883,N_23691,N_24927);
nor U28884 (N_28884,N_21481,N_23098);
xnor U28885 (N_28885,N_23497,N_21506);
nand U28886 (N_28886,N_20272,N_24127);
nor U28887 (N_28887,N_20848,N_21069);
nand U28888 (N_28888,N_22104,N_20345);
or U28889 (N_28889,N_21041,N_21817);
or U28890 (N_28890,N_24785,N_20413);
nor U28891 (N_28891,N_21324,N_22310);
nor U28892 (N_28892,N_20450,N_23687);
or U28893 (N_28893,N_20362,N_23661);
nor U28894 (N_28894,N_20256,N_23475);
nor U28895 (N_28895,N_22776,N_23278);
and U28896 (N_28896,N_20302,N_21328);
nor U28897 (N_28897,N_23388,N_23516);
or U28898 (N_28898,N_24460,N_20663);
or U28899 (N_28899,N_23378,N_24886);
nand U28900 (N_28900,N_20430,N_23186);
or U28901 (N_28901,N_20296,N_21126);
nor U28902 (N_28902,N_22597,N_23600);
xnor U28903 (N_28903,N_22723,N_21844);
and U28904 (N_28904,N_23656,N_21619);
nand U28905 (N_28905,N_22763,N_21977);
nand U28906 (N_28906,N_21498,N_20095);
and U28907 (N_28907,N_20640,N_24979);
nor U28908 (N_28908,N_24054,N_24177);
nand U28909 (N_28909,N_21542,N_21318);
nand U28910 (N_28910,N_20555,N_22934);
nand U28911 (N_28911,N_23728,N_23846);
or U28912 (N_28912,N_20942,N_23601);
nor U28913 (N_28913,N_21622,N_24995);
and U28914 (N_28914,N_23863,N_21629);
and U28915 (N_28915,N_21436,N_22396);
and U28916 (N_28916,N_24678,N_23935);
nand U28917 (N_28917,N_23457,N_20723);
and U28918 (N_28918,N_22884,N_20765);
and U28919 (N_28919,N_22943,N_24977);
or U28920 (N_28920,N_24424,N_23508);
xnor U28921 (N_28921,N_24373,N_20927);
xnor U28922 (N_28922,N_20230,N_22609);
or U28923 (N_28923,N_24025,N_21260);
nand U28924 (N_28924,N_23891,N_24538);
nor U28925 (N_28925,N_22530,N_20074);
xnor U28926 (N_28926,N_24647,N_21959);
nor U28927 (N_28927,N_24191,N_24906);
or U28928 (N_28928,N_24575,N_20595);
or U28929 (N_28929,N_21539,N_24883);
nand U28930 (N_28930,N_24263,N_20050);
nand U28931 (N_28931,N_23316,N_24253);
nor U28932 (N_28932,N_20691,N_21874);
and U28933 (N_28933,N_20410,N_24527);
and U28934 (N_28934,N_21924,N_21593);
xor U28935 (N_28935,N_21198,N_20873);
or U28936 (N_28936,N_24116,N_24189);
or U28937 (N_28937,N_20066,N_23575);
nand U28938 (N_28938,N_22661,N_24201);
or U28939 (N_28939,N_22140,N_23030);
nand U28940 (N_28940,N_22748,N_20826);
nor U28941 (N_28941,N_23703,N_24496);
nor U28942 (N_28942,N_22324,N_23263);
and U28943 (N_28943,N_24862,N_24609);
nand U28944 (N_28944,N_22762,N_20195);
nand U28945 (N_28945,N_23681,N_24849);
or U28946 (N_28946,N_23683,N_21355);
or U28947 (N_28947,N_22300,N_24421);
nand U28948 (N_28948,N_24187,N_22362);
nand U28949 (N_28949,N_21202,N_23568);
or U28950 (N_28950,N_22503,N_23954);
xnor U28951 (N_28951,N_23680,N_22670);
nor U28952 (N_28952,N_24462,N_24551);
or U28953 (N_28953,N_20600,N_20990);
and U28954 (N_28954,N_21662,N_23791);
and U28955 (N_28955,N_21504,N_20189);
nand U28956 (N_28956,N_22214,N_23011);
xnor U28957 (N_28957,N_21322,N_22973);
xnor U28958 (N_28958,N_23177,N_23711);
or U28959 (N_28959,N_23063,N_21594);
nor U28960 (N_28960,N_21125,N_20176);
nor U28961 (N_28961,N_20706,N_21043);
xnor U28962 (N_28962,N_22701,N_22388);
or U28963 (N_28963,N_23864,N_20451);
and U28964 (N_28964,N_23360,N_21844);
nor U28965 (N_28965,N_23709,N_21898);
or U28966 (N_28966,N_23248,N_21143);
xnor U28967 (N_28967,N_21627,N_20526);
and U28968 (N_28968,N_23635,N_24315);
nor U28969 (N_28969,N_21645,N_24010);
nand U28970 (N_28970,N_20920,N_22569);
xnor U28971 (N_28971,N_20628,N_21428);
or U28972 (N_28972,N_21495,N_24770);
xor U28973 (N_28973,N_21613,N_23951);
or U28974 (N_28974,N_20767,N_23726);
xor U28975 (N_28975,N_24695,N_21138);
and U28976 (N_28976,N_20360,N_21507);
nand U28977 (N_28977,N_22142,N_23546);
or U28978 (N_28978,N_24869,N_24336);
xnor U28979 (N_28979,N_20526,N_22906);
nand U28980 (N_28980,N_24163,N_23523);
or U28981 (N_28981,N_23568,N_24154);
xor U28982 (N_28982,N_24757,N_21627);
nand U28983 (N_28983,N_23119,N_23075);
nand U28984 (N_28984,N_23434,N_24880);
xor U28985 (N_28985,N_23839,N_23383);
nand U28986 (N_28986,N_21474,N_23031);
nand U28987 (N_28987,N_21178,N_20426);
and U28988 (N_28988,N_24305,N_22798);
nor U28989 (N_28989,N_20479,N_22421);
xor U28990 (N_28990,N_23571,N_20604);
xnor U28991 (N_28991,N_22399,N_21842);
xnor U28992 (N_28992,N_22431,N_22498);
and U28993 (N_28993,N_22507,N_24128);
nand U28994 (N_28994,N_20818,N_22889);
or U28995 (N_28995,N_22987,N_24122);
or U28996 (N_28996,N_22811,N_22950);
xor U28997 (N_28997,N_23314,N_22717);
nand U28998 (N_28998,N_24789,N_21715);
and U28999 (N_28999,N_21766,N_20658);
nand U29000 (N_29000,N_24858,N_22682);
xnor U29001 (N_29001,N_22065,N_21369);
or U29002 (N_29002,N_21423,N_20669);
nor U29003 (N_29003,N_24603,N_23643);
nor U29004 (N_29004,N_23654,N_22896);
xnor U29005 (N_29005,N_23432,N_24686);
nand U29006 (N_29006,N_22562,N_23629);
xor U29007 (N_29007,N_21394,N_23659);
xor U29008 (N_29008,N_23843,N_22224);
and U29009 (N_29009,N_23513,N_22405);
or U29010 (N_29010,N_21389,N_24308);
nor U29011 (N_29011,N_23086,N_21713);
nand U29012 (N_29012,N_22322,N_21547);
xnor U29013 (N_29013,N_20734,N_22046);
nand U29014 (N_29014,N_21162,N_22522);
xnor U29015 (N_29015,N_20635,N_21646);
or U29016 (N_29016,N_23673,N_20971);
and U29017 (N_29017,N_21943,N_20135);
xnor U29018 (N_29018,N_21861,N_22215);
xnor U29019 (N_29019,N_24196,N_20965);
and U29020 (N_29020,N_24051,N_20193);
and U29021 (N_29021,N_24746,N_21702);
nand U29022 (N_29022,N_20546,N_24307);
nand U29023 (N_29023,N_24409,N_21156);
nand U29024 (N_29024,N_20258,N_24495);
nand U29025 (N_29025,N_22553,N_20871);
nor U29026 (N_29026,N_20341,N_23802);
xnor U29027 (N_29027,N_24395,N_23404);
and U29028 (N_29028,N_21645,N_23045);
and U29029 (N_29029,N_20292,N_23947);
nand U29030 (N_29030,N_22428,N_24398);
xor U29031 (N_29031,N_23522,N_20379);
nand U29032 (N_29032,N_20076,N_20088);
and U29033 (N_29033,N_21916,N_21515);
nor U29034 (N_29034,N_21916,N_24969);
xnor U29035 (N_29035,N_23839,N_22924);
or U29036 (N_29036,N_23739,N_22217);
nand U29037 (N_29037,N_20120,N_22230);
nor U29038 (N_29038,N_21149,N_23349);
and U29039 (N_29039,N_24371,N_22392);
or U29040 (N_29040,N_24788,N_21795);
and U29041 (N_29041,N_20184,N_23601);
nor U29042 (N_29042,N_22815,N_20542);
nand U29043 (N_29043,N_20483,N_21999);
nor U29044 (N_29044,N_20769,N_20829);
and U29045 (N_29045,N_22320,N_20584);
nor U29046 (N_29046,N_21276,N_23001);
and U29047 (N_29047,N_24430,N_21633);
xor U29048 (N_29048,N_24927,N_20932);
nor U29049 (N_29049,N_24248,N_21082);
nand U29050 (N_29050,N_22376,N_23824);
nand U29051 (N_29051,N_20294,N_23360);
xnor U29052 (N_29052,N_24947,N_22950);
nand U29053 (N_29053,N_20768,N_24953);
or U29054 (N_29054,N_22301,N_22029);
nor U29055 (N_29055,N_23799,N_21422);
or U29056 (N_29056,N_20887,N_20124);
xor U29057 (N_29057,N_20535,N_20927);
nor U29058 (N_29058,N_22627,N_23870);
xor U29059 (N_29059,N_21151,N_21000);
xnor U29060 (N_29060,N_23439,N_20408);
and U29061 (N_29061,N_23174,N_23316);
xor U29062 (N_29062,N_23203,N_24224);
or U29063 (N_29063,N_23377,N_20076);
xor U29064 (N_29064,N_21980,N_23603);
xnor U29065 (N_29065,N_23755,N_20086);
nor U29066 (N_29066,N_22673,N_23521);
and U29067 (N_29067,N_22234,N_24320);
nor U29068 (N_29068,N_22875,N_22557);
xor U29069 (N_29069,N_21512,N_20326);
xnor U29070 (N_29070,N_20707,N_24997);
and U29071 (N_29071,N_23408,N_21818);
xnor U29072 (N_29072,N_20393,N_22841);
or U29073 (N_29073,N_24857,N_20816);
nand U29074 (N_29074,N_23979,N_24491);
nand U29075 (N_29075,N_22624,N_24695);
xor U29076 (N_29076,N_20053,N_21200);
xnor U29077 (N_29077,N_21497,N_24026);
xnor U29078 (N_29078,N_22589,N_20792);
nor U29079 (N_29079,N_22859,N_21682);
or U29080 (N_29080,N_22806,N_24774);
and U29081 (N_29081,N_23168,N_20874);
or U29082 (N_29082,N_21428,N_22913);
nor U29083 (N_29083,N_20666,N_23790);
xor U29084 (N_29084,N_22581,N_21641);
nor U29085 (N_29085,N_20958,N_23081);
nor U29086 (N_29086,N_22664,N_22219);
nand U29087 (N_29087,N_20398,N_21975);
nor U29088 (N_29088,N_24445,N_22707);
or U29089 (N_29089,N_24820,N_20589);
xor U29090 (N_29090,N_22764,N_22759);
or U29091 (N_29091,N_23213,N_22022);
nand U29092 (N_29092,N_20381,N_21921);
and U29093 (N_29093,N_24905,N_24128);
or U29094 (N_29094,N_20560,N_21694);
or U29095 (N_29095,N_24594,N_20381);
or U29096 (N_29096,N_22753,N_23411);
nor U29097 (N_29097,N_23245,N_21113);
or U29098 (N_29098,N_21981,N_21092);
nor U29099 (N_29099,N_22626,N_21283);
xnor U29100 (N_29100,N_20218,N_24913);
or U29101 (N_29101,N_24403,N_21773);
or U29102 (N_29102,N_24668,N_20556);
nand U29103 (N_29103,N_21513,N_20877);
xnor U29104 (N_29104,N_24908,N_20496);
nor U29105 (N_29105,N_21429,N_20546);
or U29106 (N_29106,N_23148,N_23678);
nor U29107 (N_29107,N_21763,N_20224);
and U29108 (N_29108,N_22697,N_21111);
or U29109 (N_29109,N_21936,N_20767);
nand U29110 (N_29110,N_21439,N_22684);
nor U29111 (N_29111,N_24914,N_22661);
or U29112 (N_29112,N_23349,N_21737);
nand U29113 (N_29113,N_22223,N_24561);
or U29114 (N_29114,N_23303,N_24678);
xnor U29115 (N_29115,N_20726,N_23628);
and U29116 (N_29116,N_20169,N_24371);
or U29117 (N_29117,N_20267,N_21750);
and U29118 (N_29118,N_22398,N_23542);
nor U29119 (N_29119,N_22919,N_22038);
and U29120 (N_29120,N_23945,N_24705);
or U29121 (N_29121,N_23123,N_23768);
and U29122 (N_29122,N_23192,N_20909);
nor U29123 (N_29123,N_22557,N_21879);
xnor U29124 (N_29124,N_22580,N_20303);
and U29125 (N_29125,N_20936,N_23023);
nand U29126 (N_29126,N_22383,N_24375);
or U29127 (N_29127,N_24054,N_22705);
and U29128 (N_29128,N_21767,N_23821);
xnor U29129 (N_29129,N_20100,N_24495);
or U29130 (N_29130,N_24556,N_20545);
nor U29131 (N_29131,N_24697,N_24210);
nor U29132 (N_29132,N_22688,N_24472);
xnor U29133 (N_29133,N_24006,N_21779);
and U29134 (N_29134,N_24351,N_23197);
and U29135 (N_29135,N_20764,N_20949);
and U29136 (N_29136,N_23762,N_23868);
and U29137 (N_29137,N_23067,N_22945);
and U29138 (N_29138,N_24033,N_22343);
or U29139 (N_29139,N_22322,N_20226);
and U29140 (N_29140,N_23975,N_21267);
and U29141 (N_29141,N_24553,N_21111);
xor U29142 (N_29142,N_22496,N_23284);
or U29143 (N_29143,N_24962,N_24701);
and U29144 (N_29144,N_20836,N_21033);
or U29145 (N_29145,N_20790,N_23442);
xnor U29146 (N_29146,N_24908,N_20473);
or U29147 (N_29147,N_20723,N_24915);
xor U29148 (N_29148,N_21322,N_20964);
nor U29149 (N_29149,N_22893,N_21014);
xor U29150 (N_29150,N_20400,N_22122);
xnor U29151 (N_29151,N_20105,N_23515);
nand U29152 (N_29152,N_20034,N_23818);
xnor U29153 (N_29153,N_23762,N_21860);
xor U29154 (N_29154,N_20521,N_21932);
nand U29155 (N_29155,N_23723,N_23054);
xor U29156 (N_29156,N_23197,N_21874);
or U29157 (N_29157,N_23848,N_21761);
xor U29158 (N_29158,N_20588,N_23182);
nor U29159 (N_29159,N_24613,N_20528);
nand U29160 (N_29160,N_24920,N_21610);
nand U29161 (N_29161,N_24068,N_21322);
and U29162 (N_29162,N_22168,N_22232);
and U29163 (N_29163,N_24358,N_22967);
nor U29164 (N_29164,N_22984,N_23559);
nand U29165 (N_29165,N_20426,N_21965);
and U29166 (N_29166,N_21311,N_21553);
nor U29167 (N_29167,N_24029,N_22167);
nand U29168 (N_29168,N_23802,N_24585);
or U29169 (N_29169,N_22882,N_20290);
and U29170 (N_29170,N_21329,N_22326);
xor U29171 (N_29171,N_23925,N_20589);
and U29172 (N_29172,N_21809,N_24974);
nand U29173 (N_29173,N_20714,N_23452);
xor U29174 (N_29174,N_24354,N_21299);
and U29175 (N_29175,N_20402,N_21865);
nand U29176 (N_29176,N_24837,N_20494);
or U29177 (N_29177,N_23254,N_23669);
nand U29178 (N_29178,N_22451,N_23145);
nand U29179 (N_29179,N_21162,N_21901);
or U29180 (N_29180,N_21334,N_23971);
xor U29181 (N_29181,N_24675,N_24212);
nand U29182 (N_29182,N_24011,N_23779);
nor U29183 (N_29183,N_24995,N_20531);
nor U29184 (N_29184,N_23471,N_21475);
nor U29185 (N_29185,N_23399,N_21513);
and U29186 (N_29186,N_23093,N_23829);
and U29187 (N_29187,N_23655,N_22433);
xnor U29188 (N_29188,N_24327,N_24792);
nand U29189 (N_29189,N_20528,N_22664);
nand U29190 (N_29190,N_21069,N_21118);
nor U29191 (N_29191,N_20549,N_21802);
nand U29192 (N_29192,N_24641,N_20328);
nor U29193 (N_29193,N_21834,N_24987);
xor U29194 (N_29194,N_22345,N_20192);
and U29195 (N_29195,N_23181,N_21443);
nand U29196 (N_29196,N_24206,N_24276);
and U29197 (N_29197,N_23688,N_23833);
xnor U29198 (N_29198,N_24170,N_24984);
xnor U29199 (N_29199,N_23208,N_24382);
nor U29200 (N_29200,N_20320,N_20016);
nor U29201 (N_29201,N_22327,N_23226);
xnor U29202 (N_29202,N_24046,N_22529);
or U29203 (N_29203,N_21577,N_22485);
xnor U29204 (N_29204,N_23004,N_21803);
or U29205 (N_29205,N_20286,N_22229);
nor U29206 (N_29206,N_24118,N_21411);
nand U29207 (N_29207,N_20985,N_23083);
nand U29208 (N_29208,N_23905,N_24489);
and U29209 (N_29209,N_22112,N_22280);
nand U29210 (N_29210,N_21089,N_24213);
nor U29211 (N_29211,N_23747,N_21516);
nor U29212 (N_29212,N_21412,N_21092);
and U29213 (N_29213,N_20674,N_21109);
and U29214 (N_29214,N_21485,N_23804);
nor U29215 (N_29215,N_22842,N_20214);
nand U29216 (N_29216,N_23368,N_20974);
xnor U29217 (N_29217,N_24317,N_23670);
or U29218 (N_29218,N_20574,N_21341);
and U29219 (N_29219,N_23146,N_20018);
nor U29220 (N_29220,N_24349,N_24558);
and U29221 (N_29221,N_22978,N_22542);
xnor U29222 (N_29222,N_22949,N_23136);
nand U29223 (N_29223,N_23385,N_21904);
or U29224 (N_29224,N_22423,N_22223);
nor U29225 (N_29225,N_21399,N_20164);
xor U29226 (N_29226,N_22470,N_21212);
or U29227 (N_29227,N_20347,N_21028);
and U29228 (N_29228,N_21713,N_24140);
xor U29229 (N_29229,N_23704,N_24742);
nand U29230 (N_29230,N_23330,N_21447);
xnor U29231 (N_29231,N_24354,N_22352);
nand U29232 (N_29232,N_23891,N_20408);
and U29233 (N_29233,N_21209,N_22333);
xnor U29234 (N_29234,N_21687,N_24493);
nand U29235 (N_29235,N_22221,N_22682);
nor U29236 (N_29236,N_20237,N_21138);
xor U29237 (N_29237,N_22951,N_24120);
nand U29238 (N_29238,N_23205,N_20568);
and U29239 (N_29239,N_20836,N_23412);
nand U29240 (N_29240,N_24652,N_21980);
xor U29241 (N_29241,N_20536,N_24547);
xor U29242 (N_29242,N_23147,N_20099);
nor U29243 (N_29243,N_20493,N_21505);
xor U29244 (N_29244,N_21560,N_21559);
nor U29245 (N_29245,N_22593,N_21139);
xor U29246 (N_29246,N_24061,N_24495);
and U29247 (N_29247,N_24503,N_20229);
nand U29248 (N_29248,N_21098,N_22247);
and U29249 (N_29249,N_24450,N_24318);
or U29250 (N_29250,N_21417,N_23357);
and U29251 (N_29251,N_22043,N_21804);
and U29252 (N_29252,N_24402,N_22308);
and U29253 (N_29253,N_21630,N_20095);
xnor U29254 (N_29254,N_22189,N_23191);
and U29255 (N_29255,N_24688,N_22643);
nor U29256 (N_29256,N_22092,N_23500);
or U29257 (N_29257,N_20832,N_22476);
nand U29258 (N_29258,N_20614,N_23977);
nor U29259 (N_29259,N_23225,N_24010);
xnor U29260 (N_29260,N_22036,N_24595);
nand U29261 (N_29261,N_20572,N_20228);
nand U29262 (N_29262,N_23647,N_23439);
and U29263 (N_29263,N_24543,N_23742);
nor U29264 (N_29264,N_23389,N_21907);
and U29265 (N_29265,N_20877,N_23748);
or U29266 (N_29266,N_20770,N_22522);
nor U29267 (N_29267,N_20171,N_22418);
nor U29268 (N_29268,N_23324,N_22814);
nand U29269 (N_29269,N_23710,N_23713);
or U29270 (N_29270,N_23906,N_20826);
and U29271 (N_29271,N_24604,N_20462);
nand U29272 (N_29272,N_23012,N_22154);
xor U29273 (N_29273,N_22902,N_20874);
nor U29274 (N_29274,N_24502,N_24588);
and U29275 (N_29275,N_24934,N_21653);
and U29276 (N_29276,N_21982,N_21916);
nor U29277 (N_29277,N_24542,N_23110);
nor U29278 (N_29278,N_24445,N_22683);
nand U29279 (N_29279,N_21602,N_20578);
nand U29280 (N_29280,N_24476,N_24390);
and U29281 (N_29281,N_22171,N_23679);
nor U29282 (N_29282,N_20942,N_23351);
and U29283 (N_29283,N_22379,N_23810);
and U29284 (N_29284,N_23932,N_22596);
xor U29285 (N_29285,N_20358,N_24826);
nand U29286 (N_29286,N_24928,N_22813);
and U29287 (N_29287,N_24896,N_23371);
nand U29288 (N_29288,N_21092,N_21730);
and U29289 (N_29289,N_23321,N_23854);
or U29290 (N_29290,N_23461,N_21383);
or U29291 (N_29291,N_22827,N_23751);
or U29292 (N_29292,N_21793,N_21295);
and U29293 (N_29293,N_23180,N_20413);
nor U29294 (N_29294,N_22861,N_23888);
xnor U29295 (N_29295,N_24358,N_21310);
nor U29296 (N_29296,N_20328,N_22693);
xnor U29297 (N_29297,N_24173,N_22839);
and U29298 (N_29298,N_21340,N_21880);
nand U29299 (N_29299,N_22612,N_20874);
and U29300 (N_29300,N_20761,N_21647);
nand U29301 (N_29301,N_23891,N_20657);
nor U29302 (N_29302,N_22190,N_21338);
nor U29303 (N_29303,N_21863,N_23111);
xor U29304 (N_29304,N_21930,N_24621);
nor U29305 (N_29305,N_24423,N_22459);
xor U29306 (N_29306,N_21307,N_20242);
nand U29307 (N_29307,N_23130,N_24229);
nor U29308 (N_29308,N_23286,N_24699);
and U29309 (N_29309,N_22651,N_24473);
or U29310 (N_29310,N_22804,N_22149);
xnor U29311 (N_29311,N_21795,N_23233);
nand U29312 (N_29312,N_24841,N_24236);
xnor U29313 (N_29313,N_21801,N_22324);
xnor U29314 (N_29314,N_21161,N_22701);
and U29315 (N_29315,N_21363,N_23098);
xnor U29316 (N_29316,N_20304,N_23869);
or U29317 (N_29317,N_24896,N_21408);
and U29318 (N_29318,N_22085,N_22176);
or U29319 (N_29319,N_23398,N_22198);
nand U29320 (N_29320,N_23181,N_22932);
or U29321 (N_29321,N_21148,N_21445);
or U29322 (N_29322,N_23226,N_24612);
nor U29323 (N_29323,N_24241,N_22698);
nor U29324 (N_29324,N_22730,N_22100);
xnor U29325 (N_29325,N_23053,N_20764);
nand U29326 (N_29326,N_21054,N_22691);
xor U29327 (N_29327,N_21121,N_20356);
and U29328 (N_29328,N_24973,N_23500);
nand U29329 (N_29329,N_22044,N_24088);
xnor U29330 (N_29330,N_21256,N_20109);
nand U29331 (N_29331,N_20811,N_23439);
xor U29332 (N_29332,N_20024,N_23399);
nor U29333 (N_29333,N_22195,N_23466);
nand U29334 (N_29334,N_24598,N_21428);
nor U29335 (N_29335,N_20823,N_22161);
xor U29336 (N_29336,N_20236,N_22372);
xor U29337 (N_29337,N_23683,N_22637);
xnor U29338 (N_29338,N_22722,N_22963);
xor U29339 (N_29339,N_21180,N_23445);
or U29340 (N_29340,N_21177,N_23254);
nand U29341 (N_29341,N_22412,N_22253);
xor U29342 (N_29342,N_21712,N_24644);
xnor U29343 (N_29343,N_22808,N_21254);
or U29344 (N_29344,N_22172,N_24407);
or U29345 (N_29345,N_21067,N_24000);
and U29346 (N_29346,N_21566,N_20915);
nand U29347 (N_29347,N_22515,N_21615);
nand U29348 (N_29348,N_21214,N_23829);
nand U29349 (N_29349,N_24743,N_23437);
and U29350 (N_29350,N_20200,N_23987);
or U29351 (N_29351,N_23321,N_22899);
nor U29352 (N_29352,N_24385,N_23460);
or U29353 (N_29353,N_23079,N_20657);
nand U29354 (N_29354,N_24446,N_23907);
or U29355 (N_29355,N_23742,N_21044);
xor U29356 (N_29356,N_22561,N_22676);
xnor U29357 (N_29357,N_23275,N_24600);
nor U29358 (N_29358,N_20194,N_21681);
xnor U29359 (N_29359,N_23376,N_20082);
nor U29360 (N_29360,N_22688,N_20133);
nand U29361 (N_29361,N_20535,N_21459);
nand U29362 (N_29362,N_24688,N_23344);
or U29363 (N_29363,N_21724,N_24801);
nand U29364 (N_29364,N_23770,N_24054);
xnor U29365 (N_29365,N_21776,N_20193);
or U29366 (N_29366,N_24458,N_22892);
nand U29367 (N_29367,N_23737,N_24866);
nor U29368 (N_29368,N_21678,N_21439);
xnor U29369 (N_29369,N_23592,N_23825);
or U29370 (N_29370,N_24775,N_20179);
or U29371 (N_29371,N_20504,N_20476);
or U29372 (N_29372,N_24539,N_21930);
nor U29373 (N_29373,N_21950,N_24614);
nand U29374 (N_29374,N_21778,N_21075);
nor U29375 (N_29375,N_24993,N_21753);
nor U29376 (N_29376,N_23660,N_20483);
and U29377 (N_29377,N_22591,N_23039);
nor U29378 (N_29378,N_21014,N_20125);
and U29379 (N_29379,N_24368,N_21408);
nor U29380 (N_29380,N_20984,N_22230);
and U29381 (N_29381,N_23567,N_21827);
or U29382 (N_29382,N_22235,N_20602);
or U29383 (N_29383,N_20240,N_21228);
xor U29384 (N_29384,N_23731,N_23591);
nor U29385 (N_29385,N_20682,N_20385);
or U29386 (N_29386,N_21973,N_22997);
and U29387 (N_29387,N_24139,N_24129);
and U29388 (N_29388,N_22309,N_20837);
or U29389 (N_29389,N_20149,N_22822);
nor U29390 (N_29390,N_23044,N_20078);
nor U29391 (N_29391,N_22584,N_20975);
or U29392 (N_29392,N_21905,N_23291);
or U29393 (N_29393,N_20834,N_22291);
and U29394 (N_29394,N_23386,N_21553);
nand U29395 (N_29395,N_23694,N_24348);
nand U29396 (N_29396,N_20612,N_24544);
and U29397 (N_29397,N_21003,N_20398);
xor U29398 (N_29398,N_23556,N_22845);
nand U29399 (N_29399,N_20250,N_24377);
xnor U29400 (N_29400,N_21476,N_23030);
xor U29401 (N_29401,N_24927,N_22399);
nor U29402 (N_29402,N_21617,N_21392);
and U29403 (N_29403,N_21117,N_24699);
nor U29404 (N_29404,N_23827,N_22372);
nor U29405 (N_29405,N_22242,N_24751);
xor U29406 (N_29406,N_20703,N_22799);
and U29407 (N_29407,N_22457,N_24225);
and U29408 (N_29408,N_20383,N_21600);
nand U29409 (N_29409,N_22389,N_22697);
nor U29410 (N_29410,N_21473,N_24796);
nor U29411 (N_29411,N_20627,N_24978);
and U29412 (N_29412,N_20239,N_21888);
or U29413 (N_29413,N_23461,N_23070);
xnor U29414 (N_29414,N_20944,N_20828);
xor U29415 (N_29415,N_21199,N_21654);
and U29416 (N_29416,N_20752,N_22474);
or U29417 (N_29417,N_21639,N_22527);
nand U29418 (N_29418,N_20500,N_22764);
or U29419 (N_29419,N_22013,N_23692);
nor U29420 (N_29420,N_20967,N_24776);
nand U29421 (N_29421,N_23905,N_20333);
nand U29422 (N_29422,N_20220,N_22682);
or U29423 (N_29423,N_21715,N_24081);
nand U29424 (N_29424,N_22212,N_23332);
xnor U29425 (N_29425,N_24107,N_21303);
or U29426 (N_29426,N_24349,N_22311);
and U29427 (N_29427,N_22371,N_23410);
nor U29428 (N_29428,N_23926,N_22096);
nor U29429 (N_29429,N_21688,N_24401);
and U29430 (N_29430,N_21169,N_21285);
nand U29431 (N_29431,N_21961,N_22392);
nor U29432 (N_29432,N_22990,N_24267);
and U29433 (N_29433,N_21671,N_21295);
nand U29434 (N_29434,N_23561,N_22857);
nand U29435 (N_29435,N_24468,N_24249);
and U29436 (N_29436,N_20230,N_20449);
xor U29437 (N_29437,N_20961,N_23685);
and U29438 (N_29438,N_24584,N_22940);
or U29439 (N_29439,N_20573,N_21431);
xor U29440 (N_29440,N_24743,N_24088);
or U29441 (N_29441,N_22008,N_24177);
nand U29442 (N_29442,N_22364,N_21703);
or U29443 (N_29443,N_24640,N_22968);
or U29444 (N_29444,N_22874,N_24270);
xnor U29445 (N_29445,N_20576,N_24915);
nand U29446 (N_29446,N_21903,N_20629);
nor U29447 (N_29447,N_20404,N_22993);
and U29448 (N_29448,N_23349,N_23113);
nor U29449 (N_29449,N_24178,N_22962);
or U29450 (N_29450,N_21243,N_20682);
and U29451 (N_29451,N_23196,N_24541);
nand U29452 (N_29452,N_22245,N_21165);
nor U29453 (N_29453,N_24750,N_23390);
nand U29454 (N_29454,N_23296,N_23743);
or U29455 (N_29455,N_23613,N_20171);
or U29456 (N_29456,N_24720,N_23436);
xnor U29457 (N_29457,N_24869,N_24388);
nor U29458 (N_29458,N_24274,N_23204);
xor U29459 (N_29459,N_21748,N_23581);
xor U29460 (N_29460,N_21338,N_23963);
xnor U29461 (N_29461,N_21500,N_23235);
or U29462 (N_29462,N_20926,N_24686);
nand U29463 (N_29463,N_20033,N_22537);
nand U29464 (N_29464,N_22582,N_21905);
or U29465 (N_29465,N_23632,N_24355);
nand U29466 (N_29466,N_21032,N_21156);
or U29467 (N_29467,N_24822,N_24156);
or U29468 (N_29468,N_22108,N_22196);
and U29469 (N_29469,N_21431,N_21127);
nand U29470 (N_29470,N_20039,N_22309);
nor U29471 (N_29471,N_22498,N_21918);
or U29472 (N_29472,N_23556,N_20610);
and U29473 (N_29473,N_22340,N_21156);
nand U29474 (N_29474,N_22566,N_23680);
xnor U29475 (N_29475,N_23765,N_20318);
and U29476 (N_29476,N_23814,N_20121);
nand U29477 (N_29477,N_23312,N_22376);
or U29478 (N_29478,N_20123,N_23462);
xnor U29479 (N_29479,N_24320,N_24206);
xnor U29480 (N_29480,N_24604,N_22249);
nor U29481 (N_29481,N_20524,N_24233);
and U29482 (N_29482,N_24656,N_21695);
and U29483 (N_29483,N_20468,N_23928);
nor U29484 (N_29484,N_23095,N_20632);
nand U29485 (N_29485,N_21102,N_21794);
or U29486 (N_29486,N_24391,N_20136);
or U29487 (N_29487,N_22336,N_24072);
nand U29488 (N_29488,N_24591,N_24102);
or U29489 (N_29489,N_23361,N_21861);
and U29490 (N_29490,N_23116,N_21073);
nand U29491 (N_29491,N_20449,N_22697);
nand U29492 (N_29492,N_24817,N_23861);
nand U29493 (N_29493,N_21299,N_20800);
nand U29494 (N_29494,N_21071,N_21915);
and U29495 (N_29495,N_23994,N_24079);
xor U29496 (N_29496,N_22121,N_24260);
or U29497 (N_29497,N_21017,N_23762);
nand U29498 (N_29498,N_23860,N_24741);
or U29499 (N_29499,N_21103,N_23540);
nand U29500 (N_29500,N_24609,N_22336);
xnor U29501 (N_29501,N_21582,N_20427);
nand U29502 (N_29502,N_21546,N_23784);
xor U29503 (N_29503,N_22903,N_20897);
nor U29504 (N_29504,N_24004,N_22270);
nand U29505 (N_29505,N_23821,N_20958);
nor U29506 (N_29506,N_23345,N_22335);
nor U29507 (N_29507,N_22471,N_23398);
nor U29508 (N_29508,N_20353,N_21213);
nand U29509 (N_29509,N_22938,N_22159);
nand U29510 (N_29510,N_22940,N_22281);
and U29511 (N_29511,N_21640,N_20146);
or U29512 (N_29512,N_21269,N_21957);
and U29513 (N_29513,N_24604,N_24005);
xor U29514 (N_29514,N_22555,N_21007);
or U29515 (N_29515,N_24456,N_22625);
nand U29516 (N_29516,N_21164,N_24168);
xor U29517 (N_29517,N_21498,N_24736);
or U29518 (N_29518,N_21650,N_22327);
nor U29519 (N_29519,N_22893,N_21153);
or U29520 (N_29520,N_23623,N_20714);
nor U29521 (N_29521,N_23374,N_22822);
nand U29522 (N_29522,N_21641,N_20123);
xnor U29523 (N_29523,N_21786,N_23823);
or U29524 (N_29524,N_20604,N_21659);
nor U29525 (N_29525,N_24470,N_21400);
nand U29526 (N_29526,N_22560,N_24650);
nand U29527 (N_29527,N_20093,N_21500);
xnor U29528 (N_29528,N_22627,N_20240);
xnor U29529 (N_29529,N_20036,N_21563);
and U29530 (N_29530,N_22936,N_21729);
and U29531 (N_29531,N_22327,N_24755);
and U29532 (N_29532,N_20076,N_23044);
and U29533 (N_29533,N_22408,N_21832);
nor U29534 (N_29534,N_24422,N_23868);
xnor U29535 (N_29535,N_20355,N_21052);
xor U29536 (N_29536,N_24506,N_21217);
nand U29537 (N_29537,N_21177,N_23388);
nor U29538 (N_29538,N_20535,N_21432);
nand U29539 (N_29539,N_21151,N_23061);
or U29540 (N_29540,N_22948,N_23420);
nand U29541 (N_29541,N_24447,N_24371);
xor U29542 (N_29542,N_20979,N_22808);
and U29543 (N_29543,N_22144,N_22936);
and U29544 (N_29544,N_24397,N_24550);
nor U29545 (N_29545,N_22045,N_21225);
nor U29546 (N_29546,N_22610,N_24498);
or U29547 (N_29547,N_23394,N_23958);
xor U29548 (N_29548,N_22861,N_24996);
and U29549 (N_29549,N_20911,N_21811);
xnor U29550 (N_29550,N_20485,N_23634);
xnor U29551 (N_29551,N_22855,N_24243);
nand U29552 (N_29552,N_23864,N_20517);
or U29553 (N_29553,N_20897,N_24724);
nor U29554 (N_29554,N_24084,N_24019);
or U29555 (N_29555,N_21700,N_22194);
and U29556 (N_29556,N_23569,N_22337);
or U29557 (N_29557,N_21650,N_21069);
nand U29558 (N_29558,N_21089,N_22617);
xnor U29559 (N_29559,N_23196,N_23317);
or U29560 (N_29560,N_21047,N_23399);
nand U29561 (N_29561,N_21027,N_21162);
nand U29562 (N_29562,N_22556,N_22111);
xnor U29563 (N_29563,N_21994,N_23322);
xnor U29564 (N_29564,N_20097,N_20129);
or U29565 (N_29565,N_20791,N_23794);
nor U29566 (N_29566,N_22822,N_23314);
nand U29567 (N_29567,N_23627,N_24211);
nand U29568 (N_29568,N_22472,N_22523);
nand U29569 (N_29569,N_22679,N_23808);
nand U29570 (N_29570,N_22501,N_24713);
nor U29571 (N_29571,N_20310,N_22159);
nor U29572 (N_29572,N_23208,N_24287);
nand U29573 (N_29573,N_24858,N_21615);
nor U29574 (N_29574,N_24222,N_20862);
xnor U29575 (N_29575,N_21829,N_24088);
nand U29576 (N_29576,N_22152,N_20718);
nand U29577 (N_29577,N_20327,N_20306);
nand U29578 (N_29578,N_24130,N_20515);
or U29579 (N_29579,N_23950,N_22038);
or U29580 (N_29580,N_20422,N_23202);
nand U29581 (N_29581,N_20820,N_20090);
xnor U29582 (N_29582,N_23513,N_23097);
nand U29583 (N_29583,N_24989,N_22768);
nand U29584 (N_29584,N_21081,N_24241);
nor U29585 (N_29585,N_24406,N_22861);
and U29586 (N_29586,N_21728,N_23191);
and U29587 (N_29587,N_24371,N_23835);
nand U29588 (N_29588,N_23093,N_22070);
nand U29589 (N_29589,N_24688,N_23817);
nor U29590 (N_29590,N_23028,N_24672);
nand U29591 (N_29591,N_24094,N_21996);
and U29592 (N_29592,N_21298,N_20560);
nor U29593 (N_29593,N_20087,N_22100);
nor U29594 (N_29594,N_22485,N_20522);
xor U29595 (N_29595,N_21396,N_23512);
nand U29596 (N_29596,N_24199,N_21905);
nand U29597 (N_29597,N_20068,N_24946);
nor U29598 (N_29598,N_21029,N_22131);
and U29599 (N_29599,N_23530,N_21415);
or U29600 (N_29600,N_22047,N_21509);
nand U29601 (N_29601,N_24923,N_23757);
and U29602 (N_29602,N_22670,N_20361);
or U29603 (N_29603,N_24171,N_23066);
nor U29604 (N_29604,N_23111,N_20954);
nor U29605 (N_29605,N_22282,N_21750);
xnor U29606 (N_29606,N_20378,N_24881);
xnor U29607 (N_29607,N_22667,N_23718);
or U29608 (N_29608,N_22948,N_22535);
xnor U29609 (N_29609,N_22053,N_24132);
nand U29610 (N_29610,N_21481,N_20458);
nand U29611 (N_29611,N_24367,N_20978);
or U29612 (N_29612,N_24230,N_21995);
xnor U29613 (N_29613,N_24483,N_24426);
xor U29614 (N_29614,N_24030,N_24228);
nand U29615 (N_29615,N_24700,N_20220);
or U29616 (N_29616,N_23260,N_23425);
nor U29617 (N_29617,N_22574,N_24260);
xnor U29618 (N_29618,N_24843,N_24333);
xor U29619 (N_29619,N_21555,N_22842);
nor U29620 (N_29620,N_20054,N_22271);
and U29621 (N_29621,N_24733,N_23997);
xor U29622 (N_29622,N_21683,N_24091);
xor U29623 (N_29623,N_22439,N_22456);
xor U29624 (N_29624,N_24384,N_22788);
xor U29625 (N_29625,N_24095,N_22133);
xor U29626 (N_29626,N_21264,N_22123);
nand U29627 (N_29627,N_22212,N_21703);
xor U29628 (N_29628,N_22036,N_20422);
and U29629 (N_29629,N_21511,N_20660);
xnor U29630 (N_29630,N_20818,N_20417);
nand U29631 (N_29631,N_21982,N_21140);
nor U29632 (N_29632,N_20359,N_22800);
or U29633 (N_29633,N_24311,N_21019);
xnor U29634 (N_29634,N_24250,N_21164);
nor U29635 (N_29635,N_24355,N_23375);
and U29636 (N_29636,N_21173,N_20074);
nor U29637 (N_29637,N_20084,N_20109);
and U29638 (N_29638,N_23665,N_24229);
nand U29639 (N_29639,N_24563,N_23840);
or U29640 (N_29640,N_21333,N_23941);
and U29641 (N_29641,N_24367,N_21031);
and U29642 (N_29642,N_21588,N_22066);
or U29643 (N_29643,N_23664,N_24479);
xnor U29644 (N_29644,N_23349,N_23613);
nand U29645 (N_29645,N_22525,N_20527);
and U29646 (N_29646,N_23086,N_23849);
and U29647 (N_29647,N_23283,N_21466);
and U29648 (N_29648,N_24708,N_21045);
xnor U29649 (N_29649,N_23976,N_24723);
nor U29650 (N_29650,N_22797,N_24852);
nor U29651 (N_29651,N_24170,N_22295);
nand U29652 (N_29652,N_21440,N_23956);
xor U29653 (N_29653,N_22104,N_24743);
xor U29654 (N_29654,N_24721,N_20894);
xor U29655 (N_29655,N_20750,N_24043);
or U29656 (N_29656,N_23487,N_20188);
or U29657 (N_29657,N_23527,N_21077);
nand U29658 (N_29658,N_24900,N_24887);
xnor U29659 (N_29659,N_21828,N_20724);
nand U29660 (N_29660,N_21161,N_20309);
nor U29661 (N_29661,N_22832,N_24295);
nand U29662 (N_29662,N_23189,N_21525);
nor U29663 (N_29663,N_20157,N_23306);
nand U29664 (N_29664,N_20916,N_24935);
nand U29665 (N_29665,N_21154,N_21808);
nor U29666 (N_29666,N_20870,N_20915);
nor U29667 (N_29667,N_20743,N_23703);
or U29668 (N_29668,N_22933,N_21475);
xor U29669 (N_29669,N_24657,N_20357);
or U29670 (N_29670,N_20430,N_20788);
or U29671 (N_29671,N_22795,N_24194);
nor U29672 (N_29672,N_21559,N_21811);
or U29673 (N_29673,N_22972,N_21060);
and U29674 (N_29674,N_22824,N_20663);
nor U29675 (N_29675,N_23027,N_20832);
nand U29676 (N_29676,N_21835,N_24415);
nor U29677 (N_29677,N_21082,N_24503);
and U29678 (N_29678,N_22123,N_24923);
or U29679 (N_29679,N_23205,N_23231);
xnor U29680 (N_29680,N_21441,N_22916);
nor U29681 (N_29681,N_20207,N_22323);
and U29682 (N_29682,N_20644,N_23557);
or U29683 (N_29683,N_23154,N_23183);
or U29684 (N_29684,N_23564,N_21973);
nor U29685 (N_29685,N_22677,N_21724);
or U29686 (N_29686,N_20798,N_23293);
or U29687 (N_29687,N_22216,N_22824);
xor U29688 (N_29688,N_21843,N_23972);
nand U29689 (N_29689,N_20914,N_20040);
or U29690 (N_29690,N_20088,N_23755);
or U29691 (N_29691,N_23572,N_23104);
or U29692 (N_29692,N_23809,N_24535);
nand U29693 (N_29693,N_24003,N_24758);
and U29694 (N_29694,N_22223,N_20795);
xnor U29695 (N_29695,N_24307,N_23534);
nor U29696 (N_29696,N_21889,N_21555);
nor U29697 (N_29697,N_24059,N_24401);
nor U29698 (N_29698,N_21438,N_23548);
nor U29699 (N_29699,N_24845,N_24864);
or U29700 (N_29700,N_21206,N_22911);
nand U29701 (N_29701,N_23137,N_22272);
xnor U29702 (N_29702,N_24875,N_20599);
and U29703 (N_29703,N_20578,N_21529);
or U29704 (N_29704,N_20658,N_22667);
nand U29705 (N_29705,N_22960,N_20754);
nand U29706 (N_29706,N_22844,N_20974);
nand U29707 (N_29707,N_21354,N_24358);
nor U29708 (N_29708,N_22667,N_20307);
nand U29709 (N_29709,N_24280,N_20348);
or U29710 (N_29710,N_20467,N_20339);
and U29711 (N_29711,N_24037,N_22543);
xor U29712 (N_29712,N_24469,N_21741);
nor U29713 (N_29713,N_24721,N_21003);
and U29714 (N_29714,N_20242,N_20385);
nor U29715 (N_29715,N_22100,N_22549);
nand U29716 (N_29716,N_20637,N_22628);
xnor U29717 (N_29717,N_22805,N_20502);
xor U29718 (N_29718,N_22884,N_20681);
xor U29719 (N_29719,N_21951,N_22153);
and U29720 (N_29720,N_21830,N_21458);
nand U29721 (N_29721,N_21453,N_24326);
and U29722 (N_29722,N_22088,N_24967);
and U29723 (N_29723,N_22643,N_20989);
nand U29724 (N_29724,N_22137,N_22539);
or U29725 (N_29725,N_20870,N_21145);
xnor U29726 (N_29726,N_21107,N_21225);
xnor U29727 (N_29727,N_24726,N_20566);
nor U29728 (N_29728,N_24813,N_22352);
nor U29729 (N_29729,N_20930,N_22679);
nor U29730 (N_29730,N_20025,N_21227);
xnor U29731 (N_29731,N_23245,N_23359);
and U29732 (N_29732,N_21517,N_20355);
nand U29733 (N_29733,N_24714,N_24158);
nand U29734 (N_29734,N_20637,N_22009);
xor U29735 (N_29735,N_22855,N_24222);
nand U29736 (N_29736,N_23845,N_22201);
nand U29737 (N_29737,N_20670,N_21648);
or U29738 (N_29738,N_20475,N_20714);
and U29739 (N_29739,N_23916,N_23803);
nor U29740 (N_29740,N_23372,N_22202);
nor U29741 (N_29741,N_22438,N_22714);
and U29742 (N_29742,N_23567,N_24460);
and U29743 (N_29743,N_24492,N_21516);
and U29744 (N_29744,N_24659,N_24431);
and U29745 (N_29745,N_22956,N_24120);
and U29746 (N_29746,N_20847,N_24001);
xnor U29747 (N_29747,N_23061,N_21183);
nand U29748 (N_29748,N_22015,N_21978);
nand U29749 (N_29749,N_24243,N_22280);
nor U29750 (N_29750,N_24143,N_20348);
xor U29751 (N_29751,N_22349,N_21456);
nor U29752 (N_29752,N_22640,N_22154);
xnor U29753 (N_29753,N_22612,N_20796);
and U29754 (N_29754,N_21615,N_22259);
nor U29755 (N_29755,N_21420,N_22072);
or U29756 (N_29756,N_23675,N_21282);
nor U29757 (N_29757,N_21919,N_24107);
xor U29758 (N_29758,N_21954,N_20955);
and U29759 (N_29759,N_23503,N_22670);
xor U29760 (N_29760,N_22635,N_20166);
xnor U29761 (N_29761,N_24628,N_24947);
nor U29762 (N_29762,N_20070,N_23967);
nand U29763 (N_29763,N_20679,N_20355);
and U29764 (N_29764,N_23449,N_23997);
or U29765 (N_29765,N_24673,N_24259);
and U29766 (N_29766,N_21471,N_23749);
and U29767 (N_29767,N_22163,N_24836);
and U29768 (N_29768,N_23417,N_22410);
or U29769 (N_29769,N_20260,N_21527);
and U29770 (N_29770,N_20127,N_21659);
and U29771 (N_29771,N_23108,N_23685);
nand U29772 (N_29772,N_21677,N_24318);
nor U29773 (N_29773,N_23841,N_21500);
or U29774 (N_29774,N_23658,N_22650);
or U29775 (N_29775,N_24324,N_24455);
xor U29776 (N_29776,N_22046,N_21772);
or U29777 (N_29777,N_24888,N_23538);
xor U29778 (N_29778,N_21250,N_20422);
nand U29779 (N_29779,N_23765,N_22842);
and U29780 (N_29780,N_23346,N_22001);
nor U29781 (N_29781,N_20579,N_22613);
xnor U29782 (N_29782,N_22463,N_21858);
or U29783 (N_29783,N_22587,N_20772);
xor U29784 (N_29784,N_24154,N_23905);
or U29785 (N_29785,N_20341,N_21377);
and U29786 (N_29786,N_21718,N_24470);
nand U29787 (N_29787,N_24415,N_21231);
xor U29788 (N_29788,N_20835,N_23876);
xnor U29789 (N_29789,N_21369,N_23953);
nand U29790 (N_29790,N_24948,N_20616);
xor U29791 (N_29791,N_23195,N_21594);
and U29792 (N_29792,N_24726,N_23829);
and U29793 (N_29793,N_21074,N_22333);
xor U29794 (N_29794,N_20882,N_21250);
nor U29795 (N_29795,N_24737,N_24815);
and U29796 (N_29796,N_24522,N_24476);
nand U29797 (N_29797,N_22601,N_24246);
nand U29798 (N_29798,N_20810,N_22664);
nand U29799 (N_29799,N_20946,N_21036);
and U29800 (N_29800,N_22154,N_22079);
nor U29801 (N_29801,N_21872,N_22541);
and U29802 (N_29802,N_24739,N_20280);
and U29803 (N_29803,N_23436,N_20273);
xor U29804 (N_29804,N_23032,N_22140);
and U29805 (N_29805,N_20340,N_22001);
and U29806 (N_29806,N_24219,N_21781);
nand U29807 (N_29807,N_20076,N_24095);
or U29808 (N_29808,N_23635,N_24564);
or U29809 (N_29809,N_22609,N_22838);
or U29810 (N_29810,N_23584,N_21182);
nor U29811 (N_29811,N_20916,N_21852);
or U29812 (N_29812,N_23030,N_20487);
nor U29813 (N_29813,N_21284,N_22828);
and U29814 (N_29814,N_23063,N_20896);
and U29815 (N_29815,N_21850,N_21947);
nand U29816 (N_29816,N_22063,N_21568);
and U29817 (N_29817,N_22330,N_21069);
xor U29818 (N_29818,N_21882,N_20006);
nand U29819 (N_29819,N_20794,N_22941);
nand U29820 (N_29820,N_23994,N_22330);
and U29821 (N_29821,N_23297,N_20817);
or U29822 (N_29822,N_20117,N_22480);
xnor U29823 (N_29823,N_24652,N_23320);
or U29824 (N_29824,N_20789,N_23752);
nand U29825 (N_29825,N_24721,N_23120);
xor U29826 (N_29826,N_21926,N_21768);
or U29827 (N_29827,N_23964,N_21931);
nor U29828 (N_29828,N_22840,N_24799);
and U29829 (N_29829,N_21403,N_21846);
or U29830 (N_29830,N_23994,N_20215);
nor U29831 (N_29831,N_24260,N_24377);
and U29832 (N_29832,N_21528,N_21903);
xnor U29833 (N_29833,N_21213,N_23322);
nor U29834 (N_29834,N_21787,N_23093);
nand U29835 (N_29835,N_23638,N_21857);
or U29836 (N_29836,N_21725,N_23039);
nor U29837 (N_29837,N_22950,N_24211);
and U29838 (N_29838,N_22478,N_21979);
and U29839 (N_29839,N_20396,N_22528);
nor U29840 (N_29840,N_20226,N_21306);
nor U29841 (N_29841,N_20200,N_24462);
nand U29842 (N_29842,N_22334,N_24548);
nand U29843 (N_29843,N_22686,N_20768);
or U29844 (N_29844,N_20394,N_21548);
or U29845 (N_29845,N_24562,N_24851);
nand U29846 (N_29846,N_21037,N_24332);
nor U29847 (N_29847,N_23761,N_23855);
xor U29848 (N_29848,N_24040,N_22457);
and U29849 (N_29849,N_21617,N_24321);
nand U29850 (N_29850,N_20941,N_22162);
or U29851 (N_29851,N_21108,N_23278);
xor U29852 (N_29852,N_24637,N_23503);
and U29853 (N_29853,N_20004,N_20940);
and U29854 (N_29854,N_23867,N_20026);
xor U29855 (N_29855,N_23036,N_23729);
or U29856 (N_29856,N_24217,N_20378);
xor U29857 (N_29857,N_24424,N_22481);
or U29858 (N_29858,N_21189,N_22530);
nand U29859 (N_29859,N_22865,N_21012);
or U29860 (N_29860,N_24039,N_21133);
or U29861 (N_29861,N_20991,N_23155);
nand U29862 (N_29862,N_23626,N_24489);
or U29863 (N_29863,N_22756,N_22162);
and U29864 (N_29864,N_23837,N_24687);
xor U29865 (N_29865,N_22440,N_23719);
nor U29866 (N_29866,N_20451,N_23501);
and U29867 (N_29867,N_21554,N_22837);
nor U29868 (N_29868,N_24276,N_24146);
nand U29869 (N_29869,N_20558,N_22298);
nor U29870 (N_29870,N_21121,N_22771);
nand U29871 (N_29871,N_20422,N_20168);
nand U29872 (N_29872,N_20646,N_24130);
nand U29873 (N_29873,N_23278,N_21111);
nor U29874 (N_29874,N_24967,N_22214);
xnor U29875 (N_29875,N_21793,N_20161);
nand U29876 (N_29876,N_21291,N_24646);
and U29877 (N_29877,N_21317,N_20271);
nand U29878 (N_29878,N_24533,N_23504);
nand U29879 (N_29879,N_21539,N_22032);
nor U29880 (N_29880,N_20977,N_20382);
or U29881 (N_29881,N_23656,N_23821);
nor U29882 (N_29882,N_24261,N_23026);
and U29883 (N_29883,N_20712,N_21736);
nor U29884 (N_29884,N_24083,N_21720);
nor U29885 (N_29885,N_22862,N_20442);
nor U29886 (N_29886,N_22490,N_23000);
or U29887 (N_29887,N_22767,N_20650);
nand U29888 (N_29888,N_24996,N_21691);
nor U29889 (N_29889,N_23836,N_23800);
and U29890 (N_29890,N_22277,N_20709);
nand U29891 (N_29891,N_24354,N_20907);
nand U29892 (N_29892,N_21430,N_22562);
xnor U29893 (N_29893,N_24067,N_22259);
and U29894 (N_29894,N_20361,N_21052);
nor U29895 (N_29895,N_21974,N_23643);
xor U29896 (N_29896,N_21106,N_23408);
or U29897 (N_29897,N_23414,N_23163);
nand U29898 (N_29898,N_21459,N_22814);
or U29899 (N_29899,N_21400,N_20176);
xnor U29900 (N_29900,N_22801,N_23342);
or U29901 (N_29901,N_23960,N_22163);
xnor U29902 (N_29902,N_23626,N_21569);
xnor U29903 (N_29903,N_22107,N_24093);
nand U29904 (N_29904,N_20204,N_24676);
xnor U29905 (N_29905,N_23524,N_24746);
or U29906 (N_29906,N_21691,N_22340);
and U29907 (N_29907,N_23060,N_20859);
nor U29908 (N_29908,N_21669,N_24069);
or U29909 (N_29909,N_20455,N_24643);
xor U29910 (N_29910,N_21675,N_24409);
and U29911 (N_29911,N_24631,N_22850);
and U29912 (N_29912,N_23136,N_22951);
xor U29913 (N_29913,N_21047,N_21396);
xor U29914 (N_29914,N_23769,N_20985);
nor U29915 (N_29915,N_20472,N_21014);
nor U29916 (N_29916,N_21279,N_23627);
or U29917 (N_29917,N_22517,N_24385);
xor U29918 (N_29918,N_24526,N_24850);
or U29919 (N_29919,N_22947,N_23029);
nand U29920 (N_29920,N_21723,N_23128);
xor U29921 (N_29921,N_24075,N_20112);
or U29922 (N_29922,N_23833,N_22521);
and U29923 (N_29923,N_22947,N_20895);
nand U29924 (N_29924,N_23958,N_22783);
nand U29925 (N_29925,N_23214,N_23389);
and U29926 (N_29926,N_20793,N_24614);
nand U29927 (N_29927,N_23906,N_22509);
xnor U29928 (N_29928,N_22905,N_20017);
nand U29929 (N_29929,N_21182,N_21852);
or U29930 (N_29930,N_21661,N_20168);
xor U29931 (N_29931,N_23044,N_20372);
nor U29932 (N_29932,N_24829,N_22468);
xnor U29933 (N_29933,N_21800,N_20392);
xor U29934 (N_29934,N_23170,N_20796);
or U29935 (N_29935,N_24243,N_24602);
and U29936 (N_29936,N_22824,N_20109);
nand U29937 (N_29937,N_22598,N_21581);
xnor U29938 (N_29938,N_21275,N_21662);
xnor U29939 (N_29939,N_20321,N_21465);
xnor U29940 (N_29940,N_20000,N_20222);
and U29941 (N_29941,N_23408,N_23860);
nor U29942 (N_29942,N_23707,N_22534);
or U29943 (N_29943,N_23661,N_21393);
or U29944 (N_29944,N_23692,N_21359);
or U29945 (N_29945,N_21634,N_21266);
xnor U29946 (N_29946,N_24550,N_22306);
nand U29947 (N_29947,N_22866,N_23939);
nand U29948 (N_29948,N_22996,N_21809);
or U29949 (N_29949,N_23717,N_21071);
and U29950 (N_29950,N_23937,N_22316);
nor U29951 (N_29951,N_24761,N_20414);
nor U29952 (N_29952,N_22580,N_22085);
and U29953 (N_29953,N_21776,N_24515);
and U29954 (N_29954,N_20521,N_20909);
nand U29955 (N_29955,N_23603,N_21443);
nand U29956 (N_29956,N_22182,N_22756);
and U29957 (N_29957,N_21431,N_22918);
and U29958 (N_29958,N_22061,N_21843);
nor U29959 (N_29959,N_20828,N_21666);
nand U29960 (N_29960,N_24796,N_24806);
or U29961 (N_29961,N_24531,N_22934);
or U29962 (N_29962,N_24556,N_22823);
and U29963 (N_29963,N_23298,N_22909);
nand U29964 (N_29964,N_24906,N_22858);
nor U29965 (N_29965,N_20439,N_23408);
or U29966 (N_29966,N_24546,N_21641);
xor U29967 (N_29967,N_24655,N_20815);
or U29968 (N_29968,N_22092,N_21650);
nand U29969 (N_29969,N_22064,N_24033);
nor U29970 (N_29970,N_23436,N_22696);
and U29971 (N_29971,N_23504,N_24992);
xnor U29972 (N_29972,N_21396,N_22215);
or U29973 (N_29973,N_21007,N_21406);
or U29974 (N_29974,N_22504,N_22045);
nand U29975 (N_29975,N_23133,N_22224);
nor U29976 (N_29976,N_20691,N_21687);
xnor U29977 (N_29977,N_22588,N_24881);
nand U29978 (N_29978,N_21391,N_21202);
or U29979 (N_29979,N_21151,N_24059);
nor U29980 (N_29980,N_20046,N_23328);
nand U29981 (N_29981,N_23690,N_20309);
and U29982 (N_29982,N_21154,N_21965);
xnor U29983 (N_29983,N_22490,N_23590);
xor U29984 (N_29984,N_20006,N_22855);
nor U29985 (N_29985,N_24434,N_21142);
nor U29986 (N_29986,N_20402,N_24996);
nor U29987 (N_29987,N_20202,N_22408);
or U29988 (N_29988,N_23747,N_23597);
nand U29989 (N_29989,N_24989,N_21798);
nor U29990 (N_29990,N_23841,N_21166);
and U29991 (N_29991,N_23813,N_23240);
xnor U29992 (N_29992,N_20853,N_20258);
or U29993 (N_29993,N_24416,N_20865);
nor U29994 (N_29994,N_21563,N_24140);
and U29995 (N_29995,N_22874,N_20271);
or U29996 (N_29996,N_23045,N_21518);
nor U29997 (N_29997,N_23655,N_24775);
or U29998 (N_29998,N_24440,N_24237);
and U29999 (N_29999,N_24974,N_21266);
xor UO_0 (O_0,N_28893,N_28169);
xor UO_1 (O_1,N_25646,N_25260);
xor UO_2 (O_2,N_28482,N_25842);
xnor UO_3 (O_3,N_27619,N_25048);
xor UO_4 (O_4,N_25485,N_29585);
nor UO_5 (O_5,N_26989,N_27068);
nand UO_6 (O_6,N_28718,N_26119);
nor UO_7 (O_7,N_26686,N_25429);
nand UO_8 (O_8,N_26205,N_27349);
or UO_9 (O_9,N_29087,N_29647);
xor UO_10 (O_10,N_29637,N_25274);
nor UO_11 (O_11,N_29706,N_26295);
nor UO_12 (O_12,N_29006,N_27576);
nor UO_13 (O_13,N_25720,N_26706);
and UO_14 (O_14,N_25947,N_26136);
xor UO_15 (O_15,N_26442,N_25359);
and UO_16 (O_16,N_28556,N_28872);
nand UO_17 (O_17,N_29520,N_27949);
nor UO_18 (O_18,N_29281,N_29317);
nor UO_19 (O_19,N_26407,N_29055);
nand UO_20 (O_20,N_29711,N_28121);
xor UO_21 (O_21,N_29673,N_25316);
nand UO_22 (O_22,N_28365,N_25886);
and UO_23 (O_23,N_26805,N_25630);
or UO_24 (O_24,N_29227,N_29631);
xnor UO_25 (O_25,N_29265,N_27411);
nor UO_26 (O_26,N_29464,N_29306);
xor UO_27 (O_27,N_25970,N_28749);
or UO_28 (O_28,N_25869,N_29714);
and UO_29 (O_29,N_27206,N_25540);
or UO_30 (O_30,N_29870,N_29615);
and UO_31 (O_31,N_25236,N_27158);
xor UO_32 (O_32,N_29307,N_25439);
nor UO_33 (O_33,N_29091,N_26497);
nor UO_34 (O_34,N_28554,N_29686);
xnor UO_35 (O_35,N_27396,N_27702);
and UO_36 (O_36,N_27503,N_28447);
xnor UO_37 (O_37,N_25923,N_25061);
nand UO_38 (O_38,N_26670,N_27104);
xnor UO_39 (O_39,N_29251,N_29429);
xor UO_40 (O_40,N_29385,N_27355);
or UO_41 (O_41,N_29873,N_29191);
nor UO_42 (O_42,N_27175,N_25373);
nor UO_43 (O_43,N_27638,N_29557);
xnor UO_44 (O_44,N_27775,N_26541);
and UO_45 (O_45,N_28859,N_29024);
xnor UO_46 (O_46,N_27896,N_27011);
and UO_47 (O_47,N_26215,N_27688);
and UO_48 (O_48,N_29021,N_27826);
nor UO_49 (O_49,N_25560,N_26879);
xnor UO_50 (O_50,N_26786,N_26367);
nor UO_51 (O_51,N_26612,N_25418);
xor UO_52 (O_52,N_29952,N_29488);
and UO_53 (O_53,N_29405,N_29209);
and UO_54 (O_54,N_26108,N_29819);
or UO_55 (O_55,N_25332,N_25212);
and UO_56 (O_56,N_25749,N_26198);
xor UO_57 (O_57,N_25997,N_28319);
or UO_58 (O_58,N_25665,N_25634);
xnor UO_59 (O_59,N_28467,N_29401);
nand UO_60 (O_60,N_27436,N_28255);
and UO_61 (O_61,N_25085,N_28524);
nor UO_62 (O_62,N_28399,N_29927);
nor UO_63 (O_63,N_25833,N_25189);
xor UO_64 (O_64,N_28147,N_28750);
nor UO_65 (O_65,N_26019,N_25738);
nor UO_66 (O_66,N_28136,N_26249);
and UO_67 (O_67,N_25153,N_26269);
and UO_68 (O_68,N_25571,N_29619);
nor UO_69 (O_69,N_26032,N_29343);
or UO_70 (O_70,N_26861,N_29574);
xor UO_71 (O_71,N_28901,N_27839);
xnor UO_72 (O_72,N_27305,N_28907);
or UO_73 (O_73,N_26624,N_29509);
or UO_74 (O_74,N_28009,N_26993);
nor UO_75 (O_75,N_28200,N_27832);
nand UO_76 (O_76,N_26838,N_29215);
and UO_77 (O_77,N_28496,N_25534);
nand UO_78 (O_78,N_25919,N_28838);
nor UO_79 (O_79,N_29526,N_27053);
and UO_80 (O_80,N_26485,N_28756);
nand UO_81 (O_81,N_29189,N_26042);
nor UO_82 (O_82,N_27549,N_25039);
nor UO_83 (O_83,N_25060,N_27783);
nor UO_84 (O_84,N_26960,N_29579);
or UO_85 (O_85,N_26554,N_26446);
nor UO_86 (O_86,N_29442,N_25849);
nand UO_87 (O_87,N_25371,N_26878);
nand UO_88 (O_88,N_26320,N_26823);
and UO_89 (O_89,N_26789,N_27891);
nor UO_90 (O_90,N_26317,N_26869);
nand UO_91 (O_91,N_27048,N_27142);
and UO_92 (O_92,N_27451,N_28353);
nor UO_93 (O_93,N_27331,N_26049);
xor UO_94 (O_94,N_29158,N_29296);
nor UO_95 (O_95,N_28818,N_29816);
nor UO_96 (O_96,N_26462,N_27185);
or UO_97 (O_97,N_25132,N_29333);
nand UO_98 (O_98,N_28313,N_25312);
nor UO_99 (O_99,N_27279,N_25953);
xnor UO_100 (O_100,N_27022,N_29116);
or UO_101 (O_101,N_28745,N_27587);
or UO_102 (O_102,N_27192,N_29182);
nand UO_103 (O_103,N_26106,N_29228);
and UO_104 (O_104,N_26752,N_27985);
nand UO_105 (O_105,N_27536,N_26586);
nor UO_106 (O_106,N_25319,N_27534);
and UO_107 (O_107,N_28646,N_25896);
nor UO_108 (O_108,N_26236,N_28805);
nor UO_109 (O_109,N_27584,N_25469);
nand UO_110 (O_110,N_25237,N_29008);
nand UO_111 (O_111,N_25504,N_29079);
nor UO_112 (O_112,N_28377,N_29436);
nand UO_113 (O_113,N_25370,N_29869);
nand UO_114 (O_114,N_28285,N_29144);
xnor UO_115 (O_115,N_26949,N_29976);
xnor UO_116 (O_116,N_25426,N_29463);
xnor UO_117 (O_117,N_29492,N_29097);
nand UO_118 (O_118,N_27656,N_26769);
nand UO_119 (O_119,N_26226,N_28110);
nor UO_120 (O_120,N_25839,N_29907);
or UO_121 (O_121,N_28519,N_29568);
nand UO_122 (O_122,N_26966,N_29051);
nand UO_123 (O_123,N_27473,N_28485);
and UO_124 (O_124,N_26221,N_29115);
and UO_125 (O_125,N_27790,N_29199);
nand UO_126 (O_126,N_27504,N_27021);
and UO_127 (O_127,N_29473,N_26073);
nand UO_128 (O_128,N_27393,N_28952);
nand UO_129 (O_129,N_27098,N_29314);
xnor UO_130 (O_130,N_25673,N_29198);
nand UO_131 (O_131,N_28663,N_26309);
nand UO_132 (O_132,N_27294,N_28426);
and UO_133 (O_133,N_29733,N_25457);
nand UO_134 (O_134,N_27151,N_25337);
and UO_135 (O_135,N_29226,N_25487);
and UO_136 (O_136,N_25003,N_27248);
or UO_137 (O_137,N_28533,N_27663);
and UO_138 (O_138,N_29774,N_27486);
and UO_139 (O_139,N_27367,N_26053);
or UO_140 (O_140,N_29025,N_25577);
nand UO_141 (O_141,N_27467,N_25706);
or UO_142 (O_142,N_27395,N_26086);
and UO_143 (O_143,N_28954,N_29089);
xor UO_144 (O_144,N_25561,N_29503);
xnor UO_145 (O_145,N_27258,N_28509);
nor UO_146 (O_146,N_28022,N_28576);
and UO_147 (O_147,N_28483,N_27023);
xnor UO_148 (O_148,N_28317,N_28171);
and UO_149 (O_149,N_25361,N_26658);
and UO_150 (O_150,N_29220,N_26833);
nor UO_151 (O_151,N_29812,N_29135);
nor UO_152 (O_152,N_26804,N_27768);
xnor UO_153 (O_153,N_27830,N_29664);
and UO_154 (O_154,N_28624,N_28058);
or UO_155 (O_155,N_28106,N_29943);
nor UO_156 (O_156,N_28234,N_28575);
nand UO_157 (O_157,N_25360,N_29868);
or UO_158 (O_158,N_28792,N_27244);
xnor UO_159 (O_159,N_28677,N_27567);
xnor UO_160 (O_160,N_25489,N_28462);
and UO_161 (O_161,N_27416,N_28812);
nor UO_162 (O_162,N_28763,N_25216);
and UO_163 (O_163,N_25968,N_29207);
xnor UO_164 (O_164,N_27629,N_25606);
nand UO_165 (O_165,N_26832,N_27550);
or UO_166 (O_166,N_29478,N_28248);
nand UO_167 (O_167,N_25270,N_25547);
xnor UO_168 (O_168,N_26599,N_25357);
or UO_169 (O_169,N_27876,N_26591);
or UO_170 (O_170,N_25082,N_27227);
and UO_171 (O_171,N_25773,N_25697);
xnor UO_172 (O_172,N_27535,N_29888);
or UO_173 (O_173,N_28804,N_26550);
and UO_174 (O_174,N_27062,N_26742);
or UO_175 (O_175,N_25403,N_26493);
nor UO_176 (O_176,N_27323,N_26260);
or UO_177 (O_177,N_25340,N_25572);
nand UO_178 (O_178,N_27910,N_26449);
xnor UO_179 (O_179,N_26441,N_28175);
or UO_180 (O_180,N_26375,N_27223);
or UO_181 (O_181,N_28358,N_27815);
or UO_182 (O_182,N_26154,N_29107);
nor UO_183 (O_183,N_28260,N_25036);
or UO_184 (O_184,N_26498,N_28985);
or UO_185 (O_185,N_26963,N_27037);
xor UO_186 (O_186,N_27383,N_27738);
xor UO_187 (O_187,N_28505,N_25442);
nand UO_188 (O_188,N_26731,N_29605);
or UO_189 (O_189,N_26836,N_27528);
xnor UO_190 (O_190,N_27615,N_25303);
and UO_191 (O_191,N_27715,N_25927);
and UO_192 (O_192,N_26327,N_28087);
xor UO_193 (O_193,N_27407,N_28210);
nand UO_194 (O_194,N_26669,N_25602);
xnor UO_195 (O_195,N_28222,N_27514);
nand UO_196 (O_196,N_26715,N_27443);
xnor UO_197 (O_197,N_27811,N_27621);
xor UO_198 (O_198,N_29528,N_25088);
xor UO_199 (O_199,N_26166,N_28359);
nand UO_200 (O_200,N_25354,N_25565);
or UO_201 (O_201,N_29577,N_29065);
nor UO_202 (O_202,N_27623,N_25820);
xor UO_203 (O_203,N_26425,N_29687);
nand UO_204 (O_204,N_29009,N_29569);
or UO_205 (O_205,N_27292,N_26971);
or UO_206 (O_206,N_26928,N_27828);
xor UO_207 (O_207,N_28207,N_25811);
or UO_208 (O_208,N_28468,N_29018);
or UO_209 (O_209,N_28033,N_25087);
nor UO_210 (O_210,N_27975,N_27445);
nor UO_211 (O_211,N_27533,N_28719);
nor UO_212 (O_212,N_28439,N_28738);
and UO_213 (O_213,N_27626,N_25247);
nor UO_214 (O_214,N_27662,N_27610);
or UO_215 (O_215,N_25201,N_27599);
xnor UO_216 (O_216,N_28654,N_28112);
nand UO_217 (O_217,N_25139,N_27878);
xor UO_218 (O_218,N_28866,N_26464);
or UO_219 (O_219,N_27952,N_29529);
xor UO_220 (O_220,N_26958,N_26028);
nor UO_221 (O_221,N_26470,N_25386);
nor UO_222 (O_222,N_28568,N_28645);
nor UO_223 (O_223,N_28461,N_26735);
or UO_224 (O_224,N_26360,N_25168);
and UO_225 (O_225,N_27564,N_29556);
nor UO_226 (O_226,N_29042,N_27287);
xnor UO_227 (O_227,N_29337,N_26620);
nor UO_228 (O_228,N_29358,N_27427);
or UO_229 (O_229,N_26180,N_26057);
nor UO_230 (O_230,N_28672,N_26622);
nand UO_231 (O_231,N_28975,N_25650);
or UO_232 (O_232,N_26834,N_25631);
xor UO_233 (O_233,N_27991,N_27356);
nor UO_234 (O_234,N_27007,N_26936);
xor UO_235 (O_235,N_29852,N_25242);
nor UO_236 (O_236,N_26068,N_26209);
or UO_237 (O_237,N_27850,N_29895);
xnor UO_238 (O_238,N_28717,N_26107);
xnor UO_239 (O_239,N_29783,N_25299);
nor UO_240 (O_240,N_25728,N_28465);
nor UO_241 (O_241,N_25541,N_26561);
or UO_242 (O_242,N_27482,N_27485);
nor UO_243 (O_243,N_26531,N_27980);
and UO_244 (O_244,N_27899,N_27620);
nor UO_245 (O_245,N_25494,N_29034);
nor UO_246 (O_246,N_25350,N_28927);
and UO_247 (O_247,N_27718,N_29519);
nand UO_248 (O_248,N_29809,N_26137);
nand UO_249 (O_249,N_28660,N_27253);
nand UO_250 (O_250,N_25273,N_29186);
xnor UO_251 (O_251,N_29997,N_25416);
or UO_252 (O_252,N_28469,N_29933);
nor UO_253 (O_253,N_28597,N_25329);
xnor UO_254 (O_254,N_27137,N_29440);
nor UO_255 (O_255,N_29621,N_25855);
and UO_256 (O_256,N_25887,N_26743);
and UO_257 (O_257,N_26120,N_26328);
nand UO_258 (O_258,N_29471,N_28449);
and UO_259 (O_259,N_25978,N_27057);
nor UO_260 (O_260,N_26457,N_25748);
nor UO_261 (O_261,N_29962,N_28497);
xnor UO_262 (O_262,N_27820,N_29902);
nor UO_263 (O_263,N_28860,N_25279);
and UO_264 (O_264,N_27459,N_26573);
nor UO_265 (O_265,N_28555,N_29530);
or UO_266 (O_266,N_26794,N_27522);
and UO_267 (O_267,N_25548,N_27505);
or UO_268 (O_268,N_25834,N_28811);
or UO_269 (O_269,N_25711,N_28902);
or UO_270 (O_270,N_29964,N_26520);
or UO_271 (O_271,N_28571,N_26835);
nand UO_272 (O_272,N_25532,N_27444);
or UO_273 (O_273,N_25815,N_29742);
nor UO_274 (O_274,N_27732,N_28266);
nand UO_275 (O_275,N_28354,N_27114);
or UO_276 (O_276,N_25344,N_25476);
or UO_277 (O_277,N_26986,N_29369);
xnor UO_278 (O_278,N_29656,N_29521);
or UO_279 (O_279,N_26718,N_29225);
nand UO_280 (O_280,N_26808,N_25217);
and UO_281 (O_281,N_28041,N_27280);
and UO_282 (O_282,N_27370,N_29630);
and UO_283 (O_283,N_27546,N_25077);
nand UO_284 (O_284,N_29623,N_25045);
and UO_285 (O_285,N_29004,N_25567);
nor UO_286 (O_286,N_28173,N_28986);
and UO_287 (O_287,N_25982,N_26456);
and UO_288 (O_288,N_27933,N_26852);
xor UO_289 (O_289,N_28869,N_29743);
and UO_290 (O_290,N_25766,N_27679);
and UO_291 (O_291,N_29030,N_27651);
xnor UO_292 (O_292,N_27088,N_26699);
xnor UO_293 (O_293,N_25911,N_27178);
and UO_294 (O_294,N_28127,N_28400);
nor UO_295 (O_295,N_26614,N_27089);
xor UO_296 (O_296,N_29078,N_25383);
xor UO_297 (O_297,N_29177,N_27959);
and UO_298 (O_298,N_29164,N_28458);
nand UO_299 (O_299,N_29154,N_29893);
and UO_300 (O_300,N_28402,N_29470);
xor UO_301 (O_301,N_29787,N_26817);
and UO_302 (O_302,N_25991,N_27747);
and UO_303 (O_303,N_25629,N_27707);
xor UO_304 (O_304,N_26499,N_29272);
or UO_305 (O_305,N_27483,N_27471);
and UO_306 (O_306,N_28101,N_29772);
nor UO_307 (O_307,N_25050,N_29214);
nor UO_308 (O_308,N_26130,N_29134);
xnor UO_309 (O_309,N_27364,N_25551);
xor UO_310 (O_310,N_25218,N_28238);
or UO_311 (O_311,N_29074,N_27851);
or UO_312 (O_312,N_29906,N_26024);
or UO_313 (O_313,N_25215,N_26719);
and UO_314 (O_314,N_29833,N_26812);
xor UO_315 (O_315,N_25222,N_28129);
or UO_316 (O_316,N_27424,N_26807);
xnor UO_317 (O_317,N_25544,N_27273);
nand UO_318 (O_318,N_29644,N_27800);
nand UO_319 (O_319,N_28998,N_28612);
and UO_320 (O_320,N_29286,N_25325);
or UO_321 (O_321,N_29183,N_27853);
nor UO_322 (O_322,N_25349,N_29766);
and UO_323 (O_323,N_29834,N_27472);
nand UO_324 (O_324,N_28513,N_26583);
or UO_325 (O_325,N_28375,N_26748);
nand UO_326 (O_326,N_26310,N_27574);
nand UO_327 (O_327,N_26113,N_25958);
xnor UO_328 (O_328,N_29865,N_25098);
nor UO_329 (O_329,N_26129,N_29562);
xnor UO_330 (O_330,N_27598,N_26605);
nand UO_331 (O_331,N_29961,N_27817);
or UO_332 (O_332,N_29323,N_26896);
xnor UO_333 (O_333,N_25961,N_28066);
or UO_334 (O_334,N_25172,N_28681);
nand UO_335 (O_335,N_25611,N_28059);
nor UO_336 (O_336,N_25717,N_29864);
and UO_337 (O_337,N_29671,N_29432);
and UO_338 (O_338,N_27887,N_26292);
xnor UO_339 (O_339,N_25230,N_25873);
nand UO_340 (O_340,N_25628,N_28079);
or UO_341 (O_341,N_25455,N_27593);
nand UO_342 (O_342,N_26004,N_25134);
nor UO_343 (O_343,N_29054,N_29632);
and UO_344 (O_344,N_28417,N_28620);
xnor UO_345 (O_345,N_28931,N_27211);
or UO_346 (O_346,N_26430,N_25674);
xor UO_347 (O_347,N_27769,N_28710);
nor UO_348 (O_348,N_29604,N_28451);
and UO_349 (O_349,N_28393,N_25019);
or UO_350 (O_350,N_28284,N_26785);
nand UO_351 (O_351,N_25778,N_26160);
xor UO_352 (O_352,N_25179,N_28583);
and UO_353 (O_353,N_25355,N_27901);
and UO_354 (O_354,N_25688,N_27698);
or UO_355 (O_355,N_25760,N_27888);
nand UO_356 (O_356,N_25497,N_25684);
nand UO_357 (O_357,N_26156,N_27784);
and UO_358 (O_358,N_29938,N_25810);
nand UO_359 (O_359,N_29827,N_29598);
and UO_360 (O_360,N_25417,N_29900);
xnor UO_361 (O_361,N_25318,N_25871);
xnor UO_362 (O_362,N_28262,N_28622);
and UO_363 (O_363,N_27753,N_29591);
or UO_364 (O_364,N_27898,N_27986);
nor UO_365 (O_365,N_29178,N_29588);
nand UO_366 (O_366,N_29941,N_26764);
and UO_367 (O_367,N_26749,N_28661);
xor UO_368 (O_368,N_29094,N_29016);
xnor UO_369 (O_369,N_25415,N_25704);
or UO_370 (O_370,N_25696,N_25928);
and UO_371 (O_371,N_25166,N_28606);
nand UO_372 (O_372,N_26631,N_28566);
xnor UO_373 (O_373,N_29691,N_28650);
and UO_374 (O_374,N_29156,N_29756);
and UO_375 (O_375,N_27777,N_29689);
nor UO_376 (O_376,N_27064,N_28126);
nor UO_377 (O_377,N_27762,N_25335);
xnor UO_378 (O_378,N_29603,N_28735);
nand UO_379 (O_379,N_26268,N_29719);
xnor UO_380 (O_380,N_27054,N_26332);
nand UO_381 (O_381,N_25155,N_27460);
or UO_382 (O_382,N_26347,N_29035);
xor UO_383 (O_383,N_28563,N_27386);
nand UO_384 (O_384,N_27469,N_27760);
nor UO_385 (O_385,N_25389,N_26151);
and UO_386 (O_386,N_29354,N_26210);
nand UO_387 (O_387,N_25980,N_29020);
nand UO_388 (O_388,N_26746,N_25280);
nor UO_389 (O_389,N_27464,N_29684);
and UO_390 (O_390,N_28137,N_28787);
and UO_391 (O_391,N_25715,N_27672);
nor UO_392 (O_392,N_27999,N_27968);
nand UO_393 (O_393,N_29146,N_29657);
and UO_394 (O_394,N_25365,N_29871);
nor UO_395 (O_395,N_25092,N_28688);
and UO_396 (O_396,N_25183,N_25814);
nand UO_397 (O_397,N_28490,N_27002);
nand UO_398 (O_398,N_26562,N_27454);
xor UO_399 (O_399,N_28236,N_29181);
nand UO_400 (O_400,N_29150,N_27819);
or UO_401 (O_401,N_26941,N_27220);
nor UO_402 (O_402,N_27600,N_25081);
nand UO_403 (O_403,N_29669,N_25755);
and UO_404 (O_404,N_29411,N_29775);
or UO_405 (O_405,N_25922,N_29947);
and UO_406 (O_406,N_28899,N_29259);
and UO_407 (O_407,N_25419,N_26518);
nand UO_408 (O_408,N_27491,N_27366);
and UO_409 (O_409,N_25459,N_28586);
nand UO_410 (O_410,N_29081,N_28746);
and UO_411 (O_411,N_25683,N_28336);
and UO_412 (O_412,N_28132,N_29650);
xor UO_413 (O_413,N_29212,N_27035);
or UO_414 (O_414,N_25671,N_27265);
nor UO_415 (O_415,N_27345,N_28167);
xnor UO_416 (O_416,N_28897,N_28435);
nand UO_417 (O_417,N_26766,N_28648);
nand UO_418 (O_418,N_25808,N_28088);
nand UO_419 (O_419,N_29174,N_26409);
or UO_420 (O_420,N_28871,N_25413);
nor UO_421 (O_421,N_29184,N_26714);
xnor UO_422 (O_422,N_28289,N_27511);
and UO_423 (O_423,N_27232,N_29512);
xor UO_424 (O_424,N_26377,N_26293);
and UO_425 (O_425,N_25470,N_25465);
xnor UO_426 (O_426,N_27010,N_28836);
and UO_427 (O_427,N_27374,N_28988);
and UO_428 (O_428,N_29913,N_25788);
or UO_429 (O_429,N_29677,N_29702);
nand UO_430 (O_430,N_26104,N_27299);
and UO_431 (O_431,N_27521,N_26738);
nand UO_432 (O_432,N_28291,N_26828);
nor UO_433 (O_433,N_28821,N_29233);
xnor UO_434 (O_434,N_28351,N_29860);
nand UO_435 (O_435,N_27967,N_25104);
xnor UO_436 (O_436,N_29216,N_25265);
nand UO_437 (O_437,N_25441,N_25669);
or UO_438 (O_438,N_29708,N_29570);
xnor UO_439 (O_439,N_26085,N_28333);
and UO_440 (O_440,N_25313,N_26813);
nor UO_441 (O_441,N_29533,N_29359);
or UO_442 (O_442,N_28923,N_29908);
xnor UO_443 (O_443,N_26267,N_25009);
nand UO_444 (O_444,N_29229,N_28537);
or UO_445 (O_445,N_27866,N_28003);
xnor UO_446 (O_446,N_27660,N_29010);
nor UO_447 (O_447,N_28054,N_25557);
nand UO_448 (O_448,N_29814,N_25816);
nor UO_449 (O_449,N_27008,N_28630);
nand UO_450 (O_450,N_29142,N_27737);
or UO_451 (O_451,N_27278,N_29840);
nor UO_452 (O_452,N_29748,N_25073);
nand UO_453 (O_453,N_27776,N_29678);
nor UO_454 (O_454,N_28771,N_25654);
xnor UO_455 (O_455,N_26133,N_27180);
xor UO_456 (O_456,N_27518,N_25402);
or UO_457 (O_457,N_26643,N_27588);
or UO_458 (O_458,N_26152,N_27654);
or UO_459 (O_459,N_26455,N_27920);
xnor UO_460 (O_460,N_27708,N_29494);
nand UO_461 (O_461,N_27647,N_28492);
xor UO_462 (O_462,N_25708,N_28094);
nand UO_463 (O_463,N_28437,N_26431);
or UO_464 (O_464,N_25352,N_27818);
and UO_465 (O_465,N_28702,N_27016);
xnor UO_466 (O_466,N_28012,N_28637);
and UO_467 (O_467,N_26373,N_26517);
xor UO_468 (O_468,N_25616,N_25493);
xor UO_469 (O_469,N_25533,N_26590);
nand UO_470 (O_470,N_29974,N_29837);
nand UO_471 (O_471,N_28316,N_26703);
nor UO_472 (O_472,N_27788,N_26444);
nand UO_473 (O_473,N_28765,N_25138);
and UO_474 (O_474,N_28679,N_27208);
and UO_475 (O_475,N_28356,N_29720);
and UO_476 (O_476,N_25897,N_25806);
nor UO_477 (O_477,N_26810,N_25185);
and UO_478 (O_478,N_25826,N_26352);
xnor UO_479 (O_479,N_27448,N_29293);
xor UO_480 (O_480,N_25458,N_29892);
or UO_481 (O_481,N_28632,N_29612);
and UO_482 (O_482,N_29362,N_29486);
or UO_483 (O_483,N_27844,N_27979);
and UO_484 (O_484,N_29994,N_27428);
xor UO_485 (O_485,N_26551,N_29434);
nor UO_486 (O_486,N_26571,N_27105);
or UO_487 (O_487,N_29608,N_25324);
nand UO_488 (O_488,N_28223,N_26117);
xor UO_489 (O_489,N_26316,N_25932);
or UO_490 (O_490,N_28241,N_27510);
xor UO_491 (O_491,N_29957,N_27456);
xor UO_492 (O_492,N_25178,N_25946);
nor UO_493 (O_493,N_28751,N_28495);
nand UO_494 (O_494,N_27316,N_25879);
and UO_495 (O_495,N_25289,N_28916);
and UO_496 (O_496,N_28168,N_26939);
and UO_497 (O_497,N_25503,N_26420);
or UO_498 (O_498,N_27059,N_27658);
xnor UO_499 (O_499,N_27578,N_28900);
nand UO_500 (O_500,N_29820,N_27298);
nand UO_501 (O_501,N_26871,N_29716);
and UO_502 (O_502,N_27197,N_25204);
and UO_503 (O_503,N_26083,N_29986);
or UO_504 (O_504,N_29878,N_27908);
or UO_505 (O_505,N_29137,N_28842);
nor UO_506 (O_506,N_25714,N_27249);
xnor UO_507 (O_507,N_29302,N_26589);
xnor UO_508 (O_508,N_26982,N_27375);
or UO_509 (O_509,N_29535,N_28172);
and UO_510 (O_510,N_25575,N_28607);
or UO_511 (O_511,N_29378,N_26237);
or UO_512 (O_512,N_28511,N_26572);
and UO_513 (O_513,N_28919,N_26625);
nand UO_514 (O_514,N_28728,N_26401);
or UO_515 (O_515,N_26897,N_25320);
nor UO_516 (O_516,N_29980,N_26502);
or UO_517 (O_517,N_27706,N_28535);
xor UO_518 (O_518,N_28943,N_25604);
and UO_519 (O_519,N_27177,N_26251);
and UO_520 (O_520,N_29430,N_25151);
and UO_521 (O_521,N_25075,N_25894);
xnor UO_522 (O_522,N_27263,N_26288);
or UO_523 (O_523,N_28956,N_29939);
and UO_524 (O_524,N_28834,N_26623);
nand UO_525 (O_525,N_27187,N_26078);
nor UO_526 (O_526,N_29755,N_25827);
nor UO_527 (O_527,N_25678,N_26335);
nor UO_528 (O_528,N_28990,N_27502);
nor UO_529 (O_529,N_25859,N_27246);
nand UO_530 (O_530,N_27722,N_27418);
xor UO_531 (O_531,N_28516,N_25774);
or UO_532 (O_532,N_26186,N_28546);
nand UO_533 (O_533,N_29095,N_26917);
nand UO_534 (O_534,N_27860,N_26406);
nor UO_535 (O_535,N_28194,N_26851);
nor UO_536 (O_536,N_26282,N_26870);
nand UO_537 (O_537,N_25328,N_26170);
xnor UO_538 (O_538,N_25942,N_27696);
and UO_539 (O_539,N_26333,N_28179);
and UO_540 (O_540,N_28529,N_27537);
xnor UO_541 (O_541,N_27988,N_28329);
and UO_542 (O_542,N_25395,N_28474);
or UO_543 (O_543,N_25852,N_26285);
or UO_544 (O_544,N_27083,N_28981);
xnor UO_545 (O_545,N_29613,N_27756);
nand UO_546 (O_546,N_29490,N_27308);
or UO_547 (O_547,N_26356,N_26182);
and UO_548 (O_548,N_27905,N_25323);
or UO_549 (O_549,N_25390,N_28669);
xor UO_550 (O_550,N_25059,N_28915);
and UO_551 (O_551,N_26592,N_28689);
xor UO_552 (O_552,N_27804,N_25154);
nand UO_553 (O_553,N_27594,N_28743);
nand UO_554 (O_554,N_27875,N_25135);
nand UO_555 (O_555,N_29426,N_28114);
or UO_556 (O_556,N_27025,N_29666);
nand UO_557 (O_557,N_29617,N_25587);
or UO_558 (O_558,N_25232,N_25233);
nand UO_559 (O_559,N_26519,N_26365);
or UO_560 (O_560,N_27138,N_29260);
xor UO_561 (O_561,N_29437,N_27923);
nand UO_562 (O_562,N_28153,N_29622);
and UO_563 (O_563,N_26781,N_28457);
or UO_564 (O_564,N_25566,N_27873);
xnor UO_565 (O_565,N_28338,N_28027);
nand UO_566 (O_566,N_29263,N_27964);
nand UO_567 (O_567,N_28189,N_25254);
or UO_568 (O_568,N_27289,N_26142);
xnor UO_569 (O_569,N_26618,N_25181);
and UO_570 (O_570,N_28557,N_28042);
nand UO_571 (O_571,N_28026,N_27982);
and UO_572 (O_572,N_27801,N_28824);
and UO_573 (O_573,N_28091,N_29360);
or UO_574 (O_574,N_27166,N_27470);
xnor UO_575 (O_575,N_28104,N_27394);
and UO_576 (O_576,N_25655,N_25028);
nor UO_577 (O_577,N_26257,N_27234);
nor UO_578 (O_578,N_28764,N_29909);
or UO_579 (O_579,N_26240,N_25012);
xor UO_580 (O_580,N_27382,N_27532);
and UO_581 (O_581,N_27517,N_26099);
xor UO_582 (O_582,N_27196,N_29979);
nand UO_583 (O_583,N_27019,N_29484);
xor UO_584 (O_584,N_29821,N_27617);
or UO_585 (O_585,N_25491,N_26248);
nand UO_586 (O_586,N_26626,N_26021);
xor UO_587 (O_587,N_27169,N_27682);
xor UO_588 (O_588,N_28456,N_27141);
xnor UO_589 (O_589,N_29731,N_26200);
or UO_590 (O_590,N_29914,N_28381);
nor UO_591 (O_591,N_26568,N_25558);
and UO_592 (O_592,N_29828,N_28401);
or UO_593 (O_593,N_29954,N_26270);
or UO_594 (O_594,N_29648,N_26514);
or UO_595 (O_595,N_27313,N_26616);
xnor UO_596 (O_596,N_25144,N_29280);
and UO_597 (O_597,N_29825,N_29773);
nand UO_598 (O_598,N_29266,N_29131);
and UO_599 (O_599,N_25651,N_26211);
or UO_600 (O_600,N_28430,N_25823);
nor UO_601 (O_601,N_27724,N_25020);
nand UO_602 (O_602,N_26468,N_28525);
xor UO_603 (O_603,N_25071,N_27183);
nor UO_604 (O_604,N_25698,N_26983);
xor UO_605 (O_605,N_25380,N_29277);
nand UO_606 (O_606,N_25789,N_28095);
and UO_607 (O_607,N_28657,N_29596);
nand UO_608 (O_608,N_26856,N_28993);
or UO_609 (O_609,N_29752,N_27224);
nand UO_610 (O_610,N_27805,N_25605);
xor UO_611 (O_611,N_27846,N_27690);
xor UO_612 (O_612,N_25642,N_25783);
xor UO_613 (O_613,N_29357,N_27604);
and UO_614 (O_614,N_26150,N_26418);
or UO_615 (O_615,N_27631,N_26475);
nor UO_616 (O_616,N_28957,N_26416);
and UO_617 (O_617,N_27757,N_26097);
nor UO_618 (O_618,N_27239,N_29396);
nor UO_619 (O_619,N_27174,N_29792);
nor UO_620 (O_620,N_27595,N_27857);
or UO_621 (O_621,N_26884,N_25187);
nor UO_622 (O_622,N_28187,N_25737);
nand UO_623 (O_623,N_29981,N_25941);
nor UO_624 (O_624,N_27121,N_29601);
or UO_625 (O_625,N_27100,N_29428);
or UO_626 (O_626,N_27139,N_25268);
nor UO_627 (O_627,N_27111,N_26175);
or UO_628 (O_628,N_25207,N_26114);
and UO_629 (O_629,N_29153,N_25142);
xnor UO_630 (O_630,N_27739,N_28877);
or UO_631 (O_631,N_27080,N_27838);
or UO_632 (O_632,N_29504,N_29790);
xor UO_633 (O_633,N_29823,N_29022);
and UO_634 (O_634,N_29759,N_26147);
and UO_635 (O_635,N_26908,N_28043);
or UO_636 (O_636,N_28322,N_29867);
or UO_637 (O_637,N_25026,N_26296);
or UO_638 (O_638,N_25130,N_27328);
and UO_639 (O_639,N_28775,N_27184);
xnor UO_640 (O_640,N_28589,N_26671);
xor UO_641 (O_641,N_26680,N_28974);
or UO_642 (O_642,N_28857,N_26740);
or UO_643 (O_643,N_27466,N_29127);
xor UO_644 (O_644,N_29236,N_27643);
or UO_645 (O_645,N_26040,N_27854);
nor UO_646 (O_646,N_25785,N_27648);
nor UO_647 (O_647,N_26010,N_28138);
or UO_648 (O_648,N_28656,N_25175);
nor UO_649 (O_649,N_28531,N_25906);
nand UO_650 (O_650,N_27721,N_25225);
and UO_651 (O_651,N_25286,N_25756);
or UO_652 (O_652,N_28452,N_29015);
nor UO_653 (O_653,N_29534,N_28647);
xnor UO_654 (O_654,N_25510,N_29168);
or UO_655 (O_655,N_27274,N_28340);
xnor UO_656 (O_656,N_27400,N_27795);
or UO_657 (O_657,N_26228,N_28802);
or UO_658 (O_658,N_25391,N_26438);
and UO_659 (O_659,N_27545,N_26560);
xnor UO_660 (O_660,N_27020,N_27406);
nand UO_661 (O_661,N_29407,N_28725);
nand UO_662 (O_662,N_25096,N_26563);
and UO_663 (O_663,N_25905,N_25645);
or UO_664 (O_664,N_25902,N_26895);
xnor UO_665 (O_665,N_26820,N_27476);
nor UO_666 (O_666,N_28784,N_25574);
or UO_667 (O_667,N_27892,N_27207);
or UO_668 (O_668,N_25300,N_26632);
nor UO_669 (O_669,N_26973,N_28086);
or UO_670 (O_670,N_29727,N_26645);
and UO_671 (O_671,N_26959,N_25310);
nor UO_672 (O_672,N_26165,N_28603);
and UO_673 (O_673,N_25841,N_27429);
and UO_674 (O_674,N_25084,N_28963);
xor UO_675 (O_675,N_25750,N_28909);
nor UO_676 (O_676,N_27608,N_26345);
or UO_677 (O_677,N_25619,N_28701);
xnor UO_678 (O_678,N_29423,N_29811);
or UO_679 (O_679,N_26189,N_25751);
nand UO_680 (O_680,N_28201,N_27094);
or UO_681 (O_681,N_28534,N_26387);
xor UO_682 (O_682,N_25192,N_29841);
xnor UO_683 (O_683,N_29060,N_29890);
xor UO_684 (O_684,N_26526,N_29090);
nor UO_685 (O_685,N_28935,N_29201);
nor UO_686 (O_686,N_29468,N_25501);
nand UO_687 (O_687,N_28267,N_28649);
xor UO_688 (O_688,N_26417,N_29053);
nand UO_689 (O_689,N_26331,N_28662);
nand UO_690 (O_690,N_27372,N_29680);
xnor UO_691 (O_691,N_28550,N_29698);
or UO_692 (O_692,N_27012,N_25379);
or UO_693 (O_693,N_25231,N_26937);
xor UO_694 (O_694,N_26535,N_29722);
and UO_695 (O_695,N_29918,N_28368);
nor UO_696 (O_696,N_25269,N_29950);
or UO_697 (O_697,N_27639,N_28800);
nand UO_698 (O_698,N_28785,N_25691);
xor UO_699 (O_699,N_28816,N_28388);
nor UO_700 (O_700,N_27508,N_27171);
or UO_701 (O_701,N_29482,N_28741);
or UO_702 (O_702,N_29170,N_26437);
and UO_703 (O_703,N_29414,N_28769);
and UO_704 (O_704,N_28712,N_28890);
and UO_705 (O_705,N_27433,N_29487);
xor UO_706 (O_706,N_27346,N_29524);
or UO_707 (O_707,N_27734,N_25462);
nor UO_708 (O_708,N_28001,N_27049);
nand UO_709 (O_709,N_29310,N_28293);
nor UO_710 (O_710,N_25495,N_28958);
nand UO_711 (O_711,N_28069,N_26298);
xor UO_712 (O_712,N_26286,N_25388);
nor UO_713 (O_713,N_25109,N_29508);
xor UO_714 (O_714,N_28111,N_28265);
or UO_715 (O_715,N_25381,N_28948);
nand UO_716 (O_716,N_29321,N_29642);
or UO_717 (O_717,N_26978,N_26448);
nand UO_718 (O_718,N_28530,N_29844);
or UO_719 (O_719,N_25498,N_29133);
nand UO_720 (O_720,N_26607,N_29450);
nor UO_721 (O_721,N_29443,N_28232);
and UO_722 (O_722,N_25305,N_29173);
nand UO_723 (O_723,N_25430,N_26326);
nor UO_724 (O_724,N_27560,N_27384);
nor UO_725 (O_725,N_27893,N_26290);
or UO_726 (O_726,N_28446,N_29166);
or UO_727 (O_727,N_29626,N_25759);
and UO_728 (O_728,N_25858,N_28191);
or UO_729 (O_729,N_29175,N_25351);
nor UO_730 (O_730,N_26544,N_29056);
nand UO_731 (O_731,N_25102,N_29910);
xor UO_732 (O_732,N_26105,N_26919);
or UO_733 (O_733,N_27074,N_25129);
or UO_734 (O_734,N_28972,N_27685);
nor UO_735 (O_735,N_27493,N_26651);
xor UO_736 (O_736,N_27625,N_26344);
nor UO_737 (O_737,N_29451,N_26172);
xnor UO_738 (O_738,N_28097,N_25200);
and UO_739 (O_739,N_28671,N_26753);
or UO_740 (O_740,N_25086,N_29651);
or UO_741 (O_741,N_29398,N_29238);
and UO_742 (O_742,N_27478,N_29300);
nand UO_743 (O_743,N_29750,N_26818);
xor UO_744 (O_744,N_28825,N_27765);
xor UO_745 (O_745,N_26829,N_26727);
xnor UO_746 (O_746,N_25235,N_27902);
nand UO_747 (O_747,N_25257,N_27509);
nand UO_748 (O_748,N_29889,N_26630);
and UO_749 (O_749,N_26100,N_28298);
nor UO_750 (O_750,N_29998,N_25211);
and UO_751 (O_751,N_28360,N_25213);
nand UO_752 (O_752,N_26745,N_26324);
nor UO_753 (O_753,N_28311,N_28036);
nor UO_754 (O_754,N_29084,N_29866);
or UO_755 (O_755,N_27350,N_26301);
xor UO_756 (O_756,N_25518,N_26102);
or UO_757 (O_757,N_25226,N_26883);
nand UO_758 (O_758,N_28983,N_29179);
or UO_759 (O_759,N_25291,N_26628);
or UO_760 (O_760,N_28618,N_25578);
and UO_761 (O_761,N_27931,N_26688);
or UO_762 (O_762,N_26319,N_26681);
xnor UO_763 (O_763,N_28826,N_28139);
or UO_764 (O_764,N_29377,N_28310);
or UO_765 (O_765,N_26931,N_25845);
or UO_766 (O_766,N_28744,N_28416);
nor UO_767 (O_767,N_26953,N_26600);
or UO_768 (O_768,N_27487,N_25209);
or UO_769 (O_769,N_29472,N_26640);
or UO_770 (O_770,N_27027,N_26481);
nand UO_771 (O_771,N_26063,N_29660);
xor UO_772 (O_772,N_28020,N_25097);
and UO_773 (O_773,N_26044,N_29966);
nand UO_774 (O_774,N_29033,N_26755);
nand UO_775 (O_775,N_28436,N_26266);
nor UO_776 (O_776,N_25609,N_29045);
or UO_777 (O_777,N_28694,N_27042);
or UO_778 (O_778,N_27262,N_26025);
xnor UO_779 (O_779,N_26933,N_25527);
or UO_780 (O_780,N_27772,N_29646);
or UO_781 (O_781,N_28770,N_29757);
xor UO_782 (O_782,N_26039,N_28004);
nor UO_783 (O_783,N_25263,N_26575);
and UO_784 (O_784,N_26369,N_28808);
xor UO_785 (O_785,N_27412,N_28881);
nand UO_786 (O_786,N_29949,N_28615);
nor UO_787 (O_787,N_25682,N_29595);
nor UO_788 (O_788,N_26708,N_26521);
or UO_789 (O_789,N_26893,N_26340);
or UO_790 (O_790,N_28999,N_29145);
nor UO_791 (O_791,N_27282,N_25610);
nor UO_792 (O_792,N_25307,N_29388);
xor UO_793 (O_793,N_27919,N_27055);
xnor UO_794 (O_794,N_29707,N_26361);
xnor UO_795 (O_795,N_27691,N_26023);
nand UO_796 (O_796,N_27179,N_25934);
and UO_797 (O_797,N_25290,N_26802);
nand UO_798 (O_798,N_27513,N_28408);
nor UO_799 (O_799,N_25034,N_25002);
xnor UO_800 (O_800,N_29194,N_29368);
and UO_801 (O_801,N_26474,N_28411);
and UO_802 (O_802,N_28696,N_25001);
xnor UO_803 (O_803,N_26556,N_29953);
or UO_804 (O_804,N_26394,N_26061);
xor UO_805 (O_805,N_25781,N_29555);
and UO_806 (O_806,N_27369,N_27544);
nor UO_807 (O_807,N_28130,N_25612);
xnor UO_808 (O_808,N_26867,N_27791);
and UO_809 (O_809,N_29005,N_26904);
or UO_810 (O_810,N_25244,N_26553);
nand UO_811 (O_811,N_26976,N_29433);
xor UO_812 (O_812,N_25726,N_25475);
nand UO_813 (O_813,N_26022,N_25687);
xnor UO_814 (O_814,N_25327,N_29242);
or UO_815 (O_815,N_27516,N_25656);
nor UO_816 (O_816,N_28673,N_28994);
or UO_817 (O_817,N_28797,N_29273);
xor UO_818 (O_818,N_26111,N_29663);
nand UO_819 (O_819,N_26603,N_29653);
or UO_820 (O_820,N_26503,N_28257);
nand UO_821 (O_821,N_29929,N_25272);
nor UO_822 (O_822,N_26830,N_29249);
nor UO_823 (O_823,N_29455,N_25221);
or UO_824 (O_824,N_25929,N_28133);
nor UO_825 (O_825,N_25302,N_26325);
nand UO_826 (O_826,N_29661,N_28300);
nor UO_827 (O_827,N_27703,N_29818);
nor UO_828 (O_828,N_28404,N_27961);
nor UO_829 (O_829,N_25509,N_25018);
nand UO_830 (O_830,N_29985,N_26523);
nand UO_831 (O_831,N_26007,N_27929);
or UO_832 (O_832,N_26682,N_27235);
or UO_833 (O_833,N_28666,N_26255);
and UO_834 (O_834,N_27976,N_26952);
xor UO_835 (O_835,N_29848,N_25293);
and UO_836 (O_836,N_29283,N_27015);
and UO_837 (O_837,N_29594,N_26677);
xnor UO_838 (O_838,N_29327,N_28995);
nor UO_839 (O_839,N_26529,N_29559);
xnor UO_840 (O_840,N_28448,N_27692);
or UO_841 (O_841,N_29649,N_29493);
and UO_842 (O_842,N_26477,N_25707);
and UO_843 (O_843,N_28527,N_29782);
nor UO_844 (O_844,N_27236,N_28538);
nor UO_845 (O_845,N_26581,N_29002);
nor UO_846 (O_846,N_28870,N_26905);
nor UO_847 (O_847,N_27761,N_25734);
xnor UO_848 (O_848,N_29881,N_26243);
nor UO_849 (O_849,N_28973,N_28506);
xnor UO_850 (O_850,N_25125,N_28149);
nand UO_851 (O_851,N_26629,N_26219);
and UO_852 (O_852,N_26793,N_25798);
nand UO_853 (O_853,N_25011,N_27627);
nor UO_854 (O_854,N_29607,N_28693);
xor UO_855 (O_855,N_27833,N_26854);
or UO_856 (O_856,N_29767,N_25570);
xnor UO_857 (O_857,N_26863,N_26355);
xor UO_858 (O_858,N_27577,N_25433);
or UO_859 (O_859,N_27835,N_29558);
nand UO_860 (O_860,N_27195,N_29830);
and UO_861 (O_861,N_27680,N_27938);
xor UO_862 (O_862,N_26938,N_26683);
and UO_863 (O_863,N_27940,N_26796);
nor UO_864 (O_864,N_26822,N_29713);
nor UO_865 (O_865,N_27130,N_26737);
nand UO_866 (O_866,N_28991,N_26397);
nand UO_867 (O_867,N_28562,N_26030);
or UO_868 (O_868,N_29693,N_28928);
nor UO_869 (O_869,N_25214,N_27309);
or UO_870 (O_870,N_29062,N_25915);
xor UO_871 (O_871,N_25637,N_28190);
nor UO_872 (O_872,N_27515,N_27455);
or UO_873 (O_873,N_25992,N_28214);
xor UO_874 (O_874,N_29379,N_28713);
nand UO_875 (O_875,N_27889,N_29506);
or UO_876 (O_876,N_25472,N_28174);
nor UO_877 (O_877,N_26776,N_26667);
nor UO_878 (O_878,N_26524,N_28766);
xor UO_879 (O_879,N_29536,N_25519);
nor UO_880 (O_880,N_25556,N_25736);
xor UO_881 (O_881,N_28945,N_28048);
nand UO_882 (O_882,N_26034,N_25835);
or UO_883 (O_883,N_27998,N_29104);
and UO_884 (O_884,N_26008,N_29497);
or UO_885 (O_885,N_29972,N_25675);
xnor UO_886 (O_886,N_29318,N_27069);
or UO_887 (O_887,N_28342,N_26092);
nor UO_888 (O_888,N_26088,N_28658);
or UO_889 (O_889,N_25309,N_25973);
and UO_890 (O_890,N_28253,N_25250);
nand UO_891 (O_891,N_26187,N_28061);
or UO_892 (O_892,N_25219,N_26103);
xnor UO_893 (O_893,N_29959,N_29924);
and UO_894 (O_894,N_29319,N_29638);
xor UO_895 (O_895,N_26005,N_28585);
xnor UO_896 (O_896,N_29467,N_26713);
xor UO_897 (O_897,N_27816,N_28697);
or UO_898 (O_898,N_25856,N_28858);
nor UO_899 (O_899,N_29798,N_26981);
and UO_900 (O_900,N_29537,N_29560);
nor UO_901 (O_901,N_25890,N_26641);
nand UO_902 (O_902,N_26239,N_28141);
nor UO_903 (O_903,N_29518,N_29301);
nand UO_904 (O_904,N_27066,N_28790);
or UO_905 (O_905,N_28941,N_29522);
nand UO_906 (O_906,N_28619,N_28574);
or UO_907 (O_907,N_27507,N_29088);
and UO_908 (O_908,N_26002,N_28050);
and UO_909 (O_909,N_26799,N_28795);
and UO_910 (O_910,N_27970,N_27989);
and UO_911 (O_911,N_27135,N_27879);
xnor UO_912 (O_912,N_28055,N_29826);
or UO_913 (O_913,N_29108,N_28540);
and UO_914 (O_914,N_26578,N_25639);
and UO_915 (O_915,N_25450,N_27547);
and UO_916 (O_916,N_27568,N_27771);
xor UO_917 (O_917,N_27565,N_27216);
nand UO_918 (O_918,N_28413,N_26087);
xor UO_919 (O_919,N_27045,N_26844);
nand UO_920 (O_920,N_25821,N_28863);
nand UO_921 (O_921,N_28580,N_26214);
nand UO_922 (O_922,N_26914,N_28906);
xnor UO_923 (O_923,N_28315,N_25240);
nor UO_924 (O_924,N_28166,N_29847);
nor UO_925 (O_925,N_29417,N_27432);
and UO_926 (O_926,N_28350,N_26432);
and UO_927 (O_927,N_28225,N_27440);
and UO_928 (O_928,N_26574,N_27150);
and UO_929 (O_929,N_28391,N_29279);
nor UO_930 (O_930,N_26000,N_28936);
or UO_931 (O_931,N_28292,N_29926);
xor UO_932 (O_932,N_25137,N_25348);
or UO_933 (O_933,N_27118,N_25794);
nand UO_934 (O_934,N_26056,N_26721);
nand UO_935 (O_935,N_29624,N_29960);
xor UO_936 (O_936,N_27422,N_28102);
xnor UO_937 (O_937,N_26067,N_28989);
and UO_938 (O_938,N_27652,N_29000);
and UO_939 (O_939,N_28049,N_28454);
or UO_940 (O_940,N_29978,N_29412);
or UO_941 (O_941,N_29485,N_26199);
or UO_942 (O_942,N_27162,N_26948);
nor UO_943 (O_943,N_27161,N_28714);
nor UO_944 (O_944,N_27450,N_28910);
or UO_945 (O_945,N_28242,N_29897);
nor UO_946 (O_946,N_28025,N_29872);
xnor UO_947 (O_947,N_26984,N_27990);
nor UO_948 (O_948,N_25925,N_25819);
nand UO_949 (O_949,N_26357,N_26545);
and UO_950 (O_950,N_25069,N_29257);
xnor UO_951 (O_951,N_28926,N_27112);
nor UO_952 (O_952,N_26066,N_27004);
or UO_953 (O_953,N_27634,N_29794);
nor UO_954 (O_954,N_26434,N_29667);
nand UO_955 (O_955,N_27694,N_27597);
and UO_956 (O_956,N_26126,N_26921);
nand UO_957 (O_957,N_27897,N_26827);
or UO_958 (O_958,N_27993,N_29725);
nand UO_959 (O_959,N_27490,N_27530);
and UO_960 (O_960,N_28788,N_29781);
and UO_961 (O_961,N_28307,N_27726);
and UO_962 (O_962,N_28779,N_26975);
and UO_963 (O_963,N_29859,N_27391);
and UO_964 (O_964,N_26913,N_28814);
or UO_965 (O_965,N_25971,N_26020);
nand UO_966 (O_966,N_29643,N_27267);
and UO_967 (O_967,N_29341,N_27176);
or UO_968 (O_968,N_29185,N_29636);
nand UO_969 (O_969,N_26465,N_28992);
or UO_970 (O_970,N_25256,N_26668);
or UO_971 (O_971,N_29151,N_29842);
or UO_972 (O_972,N_29540,N_28594);
xor UO_973 (O_973,N_29715,N_29970);
nor UO_974 (O_974,N_29041,N_29838);
nor UO_975 (O_975,N_25761,N_25853);
and UO_976 (O_976,N_27797,N_26163);
xor UO_977 (O_977,N_25779,N_27073);
and UO_978 (O_978,N_27205,N_26222);
or UO_979 (O_979,N_26471,N_28882);
xnor UO_980 (O_980,N_28481,N_27573);
or UO_981 (O_981,N_29340,N_25004);
nor UO_982 (O_982,N_27189,N_29836);
nor UO_983 (O_983,N_25049,N_27495);
or UO_984 (O_984,N_28740,N_27512);
nor UO_985 (O_985,N_28668,N_28473);
and UO_986 (O_986,N_28283,N_29723);
or UO_987 (O_987,N_26875,N_27254);
and UO_988 (O_988,N_28251,N_25460);
nand UO_989 (O_989,N_27774,N_26181);
nand UO_990 (O_990,N_28747,N_27006);
xnor UO_991 (O_991,N_25670,N_26927);
and UO_992 (O_992,N_26265,N_29329);
and UO_993 (O_993,N_27222,N_29112);
xor UO_994 (O_994,N_29734,N_29789);
or UO_995 (O_995,N_27209,N_29763);
or UO_996 (O_996,N_26478,N_26906);
nand UO_997 (O_997,N_29072,N_26555);
nor UO_998 (O_998,N_28299,N_28703);
xnor UO_999 (O_999,N_29309,N_28305);
nand UO_1000 (O_1000,N_26587,N_25404);
or UO_1001 (O_1001,N_28034,N_28453);
or UO_1002 (O_1002,N_29044,N_28099);
nand UO_1003 (O_1003,N_26758,N_27735);
nand UO_1004 (O_1004,N_27181,N_25174);
nand UO_1005 (O_1005,N_25694,N_29581);
or UO_1006 (O_1006,N_29514,N_25550);
nor UO_1007 (O_1007,N_28044,N_25770);
nor UO_1008 (O_1008,N_29491,N_25047);
nor UO_1009 (O_1009,N_27065,N_26334);
xnor UO_1010 (O_1010,N_29067,N_27855);
nor UO_1011 (O_1011,N_26079,N_26148);
xor UO_1012 (O_1012,N_28822,N_28203);
xnor UO_1013 (O_1013,N_29547,N_28664);
nor UO_1014 (O_1014,N_26258,N_26543);
or UO_1015 (O_1015,N_26792,N_26112);
nor UO_1016 (O_1016,N_25899,N_25812);
or UO_1017 (O_1017,N_27637,N_25330);
xor UO_1018 (O_1018,N_25528,N_27661);
nor UO_1019 (O_1019,N_25590,N_26321);
or UO_1020 (O_1020,N_28080,N_25700);
nor UO_1021 (O_1021,N_27468,N_25964);
nand UO_1022 (O_1022,N_28100,N_29709);
xnor UO_1023 (O_1023,N_25454,N_26841);
or UO_1024 (O_1024,N_26311,N_25977);
or UO_1025 (O_1025,N_27605,N_26427);
nand UO_1026 (O_1026,N_28051,N_28700);
xnor UO_1027 (O_1027,N_27186,N_29222);
nor UO_1028 (O_1028,N_29566,N_27705);
xnor UO_1029 (O_1029,N_29882,N_28684);
nand UO_1030 (O_1030,N_25955,N_27580);
nor UO_1031 (O_1031,N_27238,N_27984);
xor UO_1032 (O_1032,N_28093,N_26071);
and UO_1033 (O_1033,N_26422,N_28263);
nor UO_1034 (O_1034,N_25988,N_25136);
xor UO_1035 (O_1035,N_25516,N_26077);
nor UO_1036 (O_1036,N_26379,N_28376);
nand UO_1037 (O_1037,N_28971,N_26177);
nand UO_1038 (O_1038,N_25468,N_28011);
nand UO_1039 (O_1039,N_28828,N_26363);
and UO_1040 (O_1040,N_26245,N_25872);
or UO_1041 (O_1041,N_29162,N_28076);
or UO_1042 (O_1042,N_28898,N_28412);
nor UO_1043 (O_1043,N_28124,N_29211);
nand UO_1044 (O_1044,N_28245,N_27559);
nand UO_1045 (O_1045,N_29205,N_26757);
nand UO_1046 (O_1046,N_27716,N_25876);
or UO_1047 (O_1047,N_29118,N_29410);
or UO_1048 (O_1048,N_28864,N_25021);
nor UO_1049 (O_1049,N_28030,N_27955);
xnor UO_1050 (O_1050,N_26809,N_27492);
and UO_1051 (O_1051,N_29292,N_27373);
nand UO_1052 (O_1052,N_29040,N_29124);
and UO_1053 (O_1053,N_29483,N_29243);
nor UO_1054 (O_1054,N_25805,N_29052);
xnor UO_1055 (O_1055,N_28853,N_26197);
nor UO_1056 (O_1056,N_27572,N_28240);
or UO_1057 (O_1057,N_26313,N_28865);
xor UO_1058 (O_1058,N_26217,N_28334);
xor UO_1059 (O_1059,N_26987,N_29945);
nand UO_1060 (O_1060,N_25376,N_29583);
xnor UO_1061 (O_1061,N_25188,N_27748);
nand UO_1062 (O_1062,N_28774,N_25238);
xnor UO_1063 (O_1063,N_26565,N_29389);
xnor UO_1064 (O_1064,N_25106,N_25156);
or UO_1065 (O_1065,N_27664,N_26725);
nor UO_1066 (O_1066,N_28653,N_25866);
xor UO_1067 (O_1067,N_25523,N_26469);
nand UO_1068 (O_1068,N_26428,N_27480);
or UO_1069 (O_1069,N_28421,N_26299);
and UO_1070 (O_1070,N_27529,N_27883);
or UO_1071 (O_1071,N_25898,N_26035);
nor UO_1072 (O_1072,N_25514,N_26436);
nand UO_1073 (O_1073,N_25119,N_29590);
or UO_1074 (O_1074,N_25638,N_27430);
nand UO_1075 (O_1075,N_26169,N_26378);
xor UO_1076 (O_1076,N_25124,N_27426);
xnor UO_1077 (O_1077,N_26501,N_25409);
xor UO_1078 (O_1078,N_28226,N_26091);
or UO_1079 (O_1079,N_28517,N_27645);
or UO_1080 (O_1080,N_27397,N_25194);
or UO_1081 (O_1081,N_29705,N_28244);
nor UO_1082 (O_1082,N_26704,N_26204);
and UO_1083 (O_1083,N_26726,N_29395);
nor UO_1084 (O_1084,N_25730,N_28791);
nand UO_1085 (O_1085,N_28734,N_27941);
or UO_1086 (O_1086,N_25095,N_26765);
xnor UO_1087 (O_1087,N_27203,N_25264);
nor UO_1088 (O_1088,N_26846,N_27746);
and UO_1089 (O_1089,N_28539,N_26661);
nand UO_1090 (O_1090,N_25434,N_25530);
nor UO_1091 (O_1091,N_29406,N_27731);
or UO_1092 (O_1092,N_25614,N_25666);
or UO_1093 (O_1093,N_25322,N_29824);
and UO_1094 (O_1094,N_25298,N_28518);
nor UO_1095 (O_1095,N_25652,N_25939);
and UO_1096 (O_1096,N_29363,N_27170);
or UO_1097 (O_1097,N_27673,N_27780);
nand UO_1098 (O_1098,N_27842,N_25284);
nand UO_1099 (O_1099,N_27336,N_29415);
and UO_1100 (O_1100,N_26945,N_26761);
nor UO_1101 (O_1101,N_25603,N_25640);
or UO_1102 (O_1102,N_26522,N_29545);
nand UO_1103 (O_1103,N_25296,N_29447);
and UO_1104 (O_1104,N_27296,N_25521);
nand UO_1105 (O_1105,N_25889,N_29449);
nor UO_1106 (O_1106,N_27953,N_25111);
or UO_1107 (O_1107,N_29877,N_27217);
and UO_1108 (O_1108,N_28010,N_29057);
xnor UO_1109 (O_1109,N_26370,N_28565);
and UO_1110 (O_1110,N_25432,N_27675);
xor UO_1111 (O_1111,N_26246,N_27090);
xor UO_1112 (O_1112,N_25757,N_26664);
nor UO_1113 (O_1113,N_26146,N_29221);
nor UO_1114 (O_1114,N_27132,N_25729);
nor UO_1115 (O_1115,N_28096,N_29550);
nand UO_1116 (O_1116,N_27884,N_29652);
and UO_1117 (O_1117,N_27013,N_29098);
nand UO_1118 (O_1118,N_26968,N_27745);
nor UO_1119 (O_1119,N_28844,N_27488);
or UO_1120 (O_1120,N_27687,N_29739);
nor UO_1121 (O_1121,N_28883,N_26955);
and UO_1122 (O_1122,N_28193,N_29563);
or UO_1123 (O_1123,N_29372,N_28634);
nand UO_1124 (O_1124,N_29176,N_27730);
or UO_1125 (O_1125,N_26998,N_28724);
xor UO_1126 (O_1126,N_29171,N_25421);
nand UO_1127 (O_1127,N_26892,N_29352);
nor UO_1128 (O_1128,N_26341,N_27864);
nor UO_1129 (O_1129,N_27122,N_28934);
xor UO_1130 (O_1130,N_26611,N_28085);
nor UO_1131 (O_1131,N_28369,N_29155);
xnor UO_1132 (O_1132,N_27099,N_29241);
nor UO_1133 (O_1133,N_29817,N_27958);
xor UO_1134 (O_1134,N_29751,N_29899);
xnor UO_1135 (O_1135,N_27882,N_27032);
or UO_1136 (O_1136,N_29190,N_29391);
nor UO_1137 (O_1137,N_27553,N_25596);
nor UO_1138 (O_1138,N_27252,N_29765);
nor UO_1139 (O_1139,N_29313,N_26473);
or UO_1140 (O_1140,N_27438,N_25626);
nand UO_1141 (O_1141,N_27789,N_27543);
or UO_1142 (O_1142,N_25888,N_27684);
nand UO_1143 (O_1143,N_25813,N_26134);
or UO_1144 (O_1144,N_29510,N_26894);
nand UO_1145 (O_1145,N_28635,N_27569);
and UO_1146 (O_1146,N_28239,N_29641);
and UO_1147 (O_1147,N_25883,N_29635);
nand UO_1148 (O_1148,N_27525,N_29544);
nor UO_1149 (O_1149,N_25692,N_28432);
and UO_1150 (O_1150,N_26128,N_26149);
nor UO_1151 (O_1151,N_27966,N_29109);
or UO_1152 (O_1152,N_29851,N_27585);
xnor UO_1153 (O_1153,N_25382,N_26196);
or UO_1154 (O_1154,N_26576,N_25398);
and UO_1155 (O_1155,N_28593,N_27689);
and UO_1156 (O_1156,N_26940,N_25058);
xor UO_1157 (O_1157,N_26001,N_27327);
xnor UO_1158 (O_1158,N_28512,N_26201);
or UO_1159 (O_1159,N_26192,N_28024);
or UO_1160 (O_1160,N_26510,N_29967);
nor UO_1161 (O_1161,N_26532,N_28219);
or UO_1162 (O_1162,N_28809,N_25241);
or UO_1163 (O_1163,N_27602,N_26362);
and UO_1164 (O_1164,N_29760,N_26135);
and UO_1165 (O_1165,N_28984,N_28578);
and UO_1166 (O_1166,N_28982,N_27750);
nand UO_1167 (O_1167,N_29083,N_26685);
nand UO_1168 (O_1168,N_26774,N_28148);
or UO_1169 (O_1169,N_29439,N_29946);
and UO_1170 (O_1170,N_26542,N_27582);
or UO_1171 (O_1171,N_28072,N_27792);
and UO_1172 (O_1172,N_29456,N_27257);
or UO_1173 (O_1173,N_29592,N_25094);
nand UO_1174 (O_1174,N_25170,N_26540);
xnor UO_1175 (O_1175,N_25079,N_26412);
xor UO_1176 (O_1176,N_26354,N_27858);
and UO_1177 (O_1177,N_29046,N_28682);
or UO_1178 (O_1178,N_25576,N_26329);
and UO_1179 (O_1179,N_27779,N_25055);
and UO_1180 (O_1180,N_28296,N_28567);
and UO_1181 (O_1181,N_28339,N_29370);
xnor UO_1182 (O_1182,N_29564,N_25681);
and UO_1183 (O_1183,N_25712,N_25447);
and UO_1184 (O_1184,N_29435,N_28158);
nor UO_1185 (O_1185,N_26798,N_26242);
and UO_1186 (O_1186,N_26548,N_25145);
nor UO_1187 (O_1187,N_28279,N_28912);
xor UO_1188 (O_1188,N_28726,N_29863);
xor UO_1189 (O_1189,N_26054,N_29063);
and UO_1190 (O_1190,N_27160,N_28277);
xnor UO_1191 (O_1191,N_25769,N_25308);
xnor UO_1192 (O_1192,N_27947,N_25032);
nor UO_1193 (O_1193,N_25522,N_27277);
nand UO_1194 (O_1194,N_28206,N_29304);
nand UO_1195 (O_1195,N_27880,N_28803);
or UO_1196 (O_1196,N_28856,N_28098);
or UO_1197 (O_1197,N_28861,N_29628);
nand UO_1198 (O_1198,N_26570,N_27921);
xnor UO_1199 (O_1199,N_27325,N_26405);
nand UO_1200 (O_1200,N_28855,N_25701);
xor UO_1201 (O_1201,N_27072,N_26773);
xor UO_1202 (O_1202,N_29777,N_28215);
or UO_1203 (O_1203,N_29400,N_27034);
nor UO_1204 (O_1204,N_29741,N_28108);
xor UO_1205 (O_1205,N_28843,N_25262);
nor UO_1206 (O_1206,N_27796,N_25710);
nor UO_1207 (O_1207,N_25267,N_28117);
nor UO_1208 (O_1208,N_29459,N_28614);
xor UO_1209 (O_1209,N_25893,N_25375);
nand UO_1210 (O_1210,N_28345,N_27720);
and UO_1211 (O_1211,N_28143,N_25830);
xnor UO_1212 (O_1212,N_26491,N_28438);
xor UO_1213 (O_1213,N_25624,N_28794);
nor UO_1214 (O_1214,N_25969,N_27437);
xor UO_1215 (O_1215,N_29113,N_29553);
or UO_1216 (O_1216,N_26674,N_29246);
or UO_1217 (O_1217,N_26882,N_28727);
nor UO_1218 (O_1218,N_26124,N_28762);
or UO_1219 (O_1219,N_27247,N_26159);
or UO_1220 (O_1220,N_25110,N_26868);
nand UO_1221 (O_1221,N_26395,N_25972);
nor UO_1222 (O_1222,N_26741,N_28445);
or UO_1223 (O_1223,N_27678,N_27589);
nand UO_1224 (O_1224,N_27115,N_28212);
nor UO_1225 (O_1225,N_27928,N_27686);
nor UO_1226 (O_1226,N_27484,N_26734);
nand UO_1227 (O_1227,N_28911,N_28605);
or UO_1228 (O_1228,N_29898,N_26500);
nor UO_1229 (O_1229,N_29948,N_28349);
nor UO_1230 (O_1230,N_27538,N_25524);
xor UO_1231 (O_1231,N_25920,N_28103);
nor UO_1232 (O_1232,N_27773,N_27043);
nor UO_1233 (O_1233,N_28949,N_27303);
nor UO_1234 (O_1234,N_29172,N_27847);
and UO_1235 (O_1235,N_28639,N_27018);
nor UO_1236 (O_1236,N_26654,N_29513);
and UO_1237 (O_1237,N_29353,N_25594);
nor UO_1238 (O_1238,N_26997,N_27736);
nor UO_1239 (O_1239,N_29589,N_27338);
or UO_1240 (O_1240,N_28667,N_25425);
and UO_1241 (O_1241,N_25986,N_27603);
or UO_1242 (O_1242,N_25167,N_29036);
xnor UO_1243 (O_1243,N_28362,N_29832);
nand UO_1244 (O_1244,N_25952,N_28157);
and UO_1245 (O_1245,N_25951,N_29894);
nand UO_1246 (O_1246,N_28424,N_26081);
and UO_1247 (O_1247,N_28514,N_25007);
nor UO_1248 (O_1248,N_28182,N_28455);
nor UO_1249 (O_1249,N_27699,N_26932);
and UO_1250 (O_1250,N_25822,N_25486);
and UO_1251 (O_1251,N_29334,N_29461);
or UO_1252 (O_1252,N_29100,N_29549);
xor UO_1253 (O_1253,N_27727,N_25542);
or UO_1254 (O_1254,N_26815,N_27922);
and UO_1255 (O_1255,N_27479,N_28628);
xnor UO_1256 (O_1256,N_25851,N_25505);
nand UO_1257 (O_1257,N_29294,N_28199);
xor UO_1258 (O_1258,N_27946,N_26593);
nor UO_1259 (O_1259,N_25793,N_26964);
or UO_1260 (O_1260,N_27950,N_29161);
nor UO_1261 (O_1261,N_28204,N_28918);
nor UO_1262 (O_1262,N_26819,N_27934);
nor UO_1263 (O_1263,N_29931,N_25116);
nor UO_1264 (O_1264,N_26970,N_29316);
and UO_1265 (O_1265,N_25334,N_26018);
nand UO_1266 (O_1266,N_25401,N_25949);
or UO_1267 (O_1267,N_26116,N_25787);
nand UO_1268 (O_1268,N_26036,N_29921);
or UO_1269 (O_1269,N_27871,N_29726);
xor UO_1270 (O_1270,N_28163,N_29206);
and UO_1271 (O_1271,N_26803,N_25143);
nor UO_1272 (O_1272,N_26230,N_29915);
nor UO_1273 (O_1273,N_29712,N_26676);
nor UO_1274 (O_1274,N_27579,N_29806);
and UO_1275 (O_1275,N_28008,N_28420);
nand UO_1276 (O_1276,N_29969,N_27563);
and UO_1277 (O_1277,N_25742,N_27810);
or UO_1278 (O_1278,N_26779,N_26694);
nor UO_1279 (O_1279,N_29676,N_28188);
or UO_1280 (O_1280,N_28504,N_29668);
xor UO_1281 (O_1281,N_29130,N_28144);
nand UO_1282 (O_1282,N_29849,N_29688);
or UO_1283 (O_1283,N_27159,N_25294);
nor UO_1284 (O_1284,N_28867,N_29122);
or UO_1285 (O_1285,N_28545,N_27398);
and UO_1286 (O_1286,N_29835,N_29797);
xor UO_1287 (O_1287,N_25121,N_27912);
nand UO_1288 (O_1288,N_25161,N_26689);
and UO_1289 (O_1289,N_26579,N_29499);
and UO_1290 (O_1290,N_25719,N_29618);
and UO_1291 (O_1291,N_26353,N_29879);
nor UO_1292 (O_1292,N_28904,N_26736);
or UO_1293 (O_1293,N_28387,N_28005);
nand UO_1294 (O_1294,N_27458,N_29887);
nand UO_1295 (O_1295,N_27075,N_26303);
or UO_1296 (O_1296,N_25954,N_29469);
and UO_1297 (O_1297,N_26213,N_27640);
nor UO_1298 (O_1298,N_28781,N_29861);
or UO_1299 (O_1299,N_28611,N_28007);
xnor UO_1300 (O_1300,N_25304,N_27047);
or UO_1301 (O_1301,N_29270,N_26484);
nand UO_1302 (O_1302,N_28131,N_28014);
nor UO_1303 (O_1303,N_28799,N_25517);
or UO_1304 (O_1304,N_28304,N_29717);
or UO_1305 (O_1305,N_27155,N_27695);
or UO_1306 (O_1306,N_27868,N_29788);
xnor UO_1307 (O_1307,N_25027,N_28160);
or UO_1308 (O_1308,N_27210,N_28364);
nor UO_1309 (O_1309,N_27609,N_27520);
xor UO_1310 (O_1310,N_25013,N_26256);
and UO_1311 (O_1311,N_27332,N_28070);
nand UO_1312 (O_1312,N_26657,N_26886);
xnor UO_1313 (O_1313,N_28314,N_27193);
nand UO_1314 (O_1314,N_25895,N_29735);
nor UO_1315 (O_1315,N_25173,N_29905);
xor UO_1316 (O_1316,N_27932,N_26885);
and UO_1317 (O_1317,N_26816,N_25537);
or UO_1318 (O_1318,N_28891,N_25199);
nand UO_1319 (O_1319,N_27763,N_29850);
xnor UO_1320 (O_1320,N_29136,N_29704);
and UO_1321 (O_1321,N_29498,N_27199);
xnor UO_1322 (O_1322,N_27717,N_29575);
nor UO_1323 (O_1323,N_26795,N_28065);
and UO_1324 (O_1324,N_28231,N_25220);
and UO_1325 (O_1325,N_26229,N_28691);
nand UO_1326 (O_1326,N_27794,N_29610);
and UO_1327 (O_1327,N_28367,N_29125);
nor UO_1328 (O_1328,N_28705,N_27942);
xor UO_1329 (O_1329,N_29371,N_25621);
nand UO_1330 (O_1330,N_25243,N_27275);
or UO_1331 (O_1331,N_28708,N_25427);
or UO_1332 (O_1332,N_29059,N_26090);
or UO_1333 (O_1333,N_29940,N_26350);
or UO_1334 (O_1334,N_25758,N_29290);
xor UO_1335 (O_1335,N_28616,N_25862);
and UO_1336 (O_1336,N_25739,N_25938);
xnor UO_1337 (O_1337,N_29408,N_29285);
and UO_1338 (O_1338,N_26173,N_26811);
xor UO_1339 (O_1339,N_27644,N_26062);
or UO_1340 (O_1340,N_26527,N_26391);
nand UO_1341 (O_1341,N_27086,N_28754);
and UO_1342 (O_1342,N_29779,N_25543);
or UO_1343 (O_1343,N_28950,N_28414);
and UO_1344 (O_1344,N_25967,N_29431);
or UO_1345 (O_1345,N_27061,N_26900);
and UO_1346 (O_1346,N_29465,N_27895);
nor UO_1347 (O_1347,N_29393,N_25583);
or UO_1348 (O_1348,N_26451,N_26837);
nand UO_1349 (O_1349,N_25563,N_28623);
nand UO_1350 (O_1350,N_29542,N_25994);
or UO_1351 (O_1351,N_26538,N_27915);
and UO_1352 (O_1352,N_26516,N_26366);
or UO_1353 (O_1353,N_25063,N_29232);
xnor UO_1354 (O_1354,N_27110,N_29424);
xnor UO_1355 (O_1355,N_27399,N_28964);
and UO_1356 (O_1356,N_27291,N_25985);
nor UO_1357 (O_1357,N_27713,N_27701);
or UO_1358 (O_1358,N_27251,N_29367);
xnor UO_1359 (O_1359,N_29195,N_27996);
nor UO_1360 (O_1360,N_25396,N_26806);
nor UO_1361 (O_1361,N_25880,N_26733);
nor UO_1362 (O_1362,N_28685,N_25618);
xnor UO_1363 (O_1363,N_29192,N_29843);
nand UO_1364 (O_1364,N_29076,N_26801);
and UO_1365 (O_1365,N_26767,N_29267);
nor UO_1366 (O_1366,N_28500,N_25040);
and UO_1367 (O_1367,N_25062,N_28920);
and UO_1368 (O_1368,N_29394,N_29496);
and UO_1369 (O_1369,N_25892,N_26638);
nor UO_1370 (O_1370,N_29699,N_29322);
and UO_1371 (O_1371,N_25767,N_25664);
xor UO_1372 (O_1372,N_26297,N_25507);
xor UO_1373 (O_1373,N_26967,N_26421);
xor UO_1374 (O_1374,N_26487,N_28275);
nand UO_1375 (O_1375,N_29262,N_26866);
nand UO_1376 (O_1376,N_29282,N_26992);
nand UO_1377 (O_1377,N_25281,N_25996);
and UO_1378 (O_1378,N_25101,N_26075);
nor UO_1379 (O_1379,N_28060,N_25554);
and UO_1380 (O_1380,N_25152,N_29593);
and UO_1381 (O_1381,N_26231,N_27937);
and UO_1382 (O_1382,N_26717,N_26876);
and UO_1383 (O_1383,N_27969,N_26390);
nor UO_1384 (O_1384,N_28896,N_26881);
and UO_1385 (O_1385,N_28297,N_27807);
xnor UO_1386 (O_1386,N_26642,N_26411);
or UO_1387 (O_1387,N_27163,N_25445);
xnor UO_1388 (O_1388,N_27307,N_29441);
nor UO_1389 (O_1389,N_28595,N_26843);
and UO_1390 (O_1390,N_26505,N_28507);
nand UO_1391 (O_1391,N_29284,N_28813);
xnor UO_1392 (O_1392,N_26308,N_25647);
nand UO_1393 (O_1393,N_26318,N_26480);
or UO_1394 (O_1394,N_29539,N_27907);
nor UO_1395 (O_1395,N_26716,N_28252);
and UO_1396 (O_1396,N_28807,N_28276);
nor UO_1397 (O_1397,N_27060,N_28357);
nand UO_1398 (O_1398,N_29732,N_29747);
and UO_1399 (O_1399,N_25484,N_29987);
nor UO_1400 (O_1400,N_29460,N_26613);
nor UO_1401 (O_1401,N_28135,N_26627);
xor UO_1402 (O_1402,N_28521,N_29332);
nand UO_1403 (O_1403,N_25078,N_26609);
xnor UO_1404 (O_1404,N_25735,N_28221);
nor UO_1405 (O_1405,N_25539,N_26839);
nor UO_1406 (O_1406,N_26698,N_26424);
or UO_1407 (O_1407,N_27264,N_28450);
xnor UO_1408 (O_1408,N_26957,N_29662);
and UO_1409 (O_1409,N_25625,N_25483);
xnor UO_1410 (O_1410,N_26509,N_28946);
nor UO_1411 (O_1411,N_29988,N_26089);
xnor UO_1412 (O_1412,N_26241,N_29516);
or UO_1413 (O_1413,N_26031,N_28406);
or UO_1414 (O_1414,N_29031,N_28463);
xnor UO_1415 (O_1415,N_29973,N_27917);
nor UO_1416 (O_1416,N_28845,N_29421);
nand UO_1417 (O_1417,N_29308,N_27916);
xnor UO_1418 (O_1418,N_25347,N_29288);
xor UO_1419 (O_1419,N_29159,N_29770);
nor UO_1420 (O_1420,N_29248,N_28885);
or UO_1421 (O_1421,N_25015,N_29117);
xor UO_1422 (O_1422,N_27886,N_25099);
or UO_1423 (O_1423,N_26191,N_25252);
nor UO_1424 (O_1424,N_27165,N_28218);
xor UO_1425 (O_1425,N_27250,N_27987);
nor UO_1426 (O_1426,N_27028,N_28146);
nand UO_1427 (O_1427,N_29239,N_28046);
nand UO_1428 (O_1428,N_29276,N_26376);
xor UO_1429 (O_1429,N_26965,N_28875);
or UO_1430 (O_1430,N_29479,N_27741);
and UO_1431 (O_1431,N_28777,N_26176);
nand UO_1432 (O_1432,N_29254,N_26276);
and UO_1433 (O_1433,N_26705,N_28475);
nand UO_1434 (O_1434,N_29552,N_26388);
nor UO_1435 (O_1435,N_29578,N_27168);
xnor UO_1436 (O_1436,N_25428,N_29531);
xnor UO_1437 (O_1437,N_27729,N_28652);
xor UO_1438 (O_1438,N_25407,N_26771);
nor UO_1439 (O_1439,N_27256,N_25275);
or UO_1440 (O_1440,N_27744,N_25790);
or UO_1441 (O_1441,N_25868,N_28959);
and UO_1442 (O_1442,N_26323,N_26358);
xor UO_1443 (O_1443,N_28880,N_28017);
and UO_1444 (O_1444,N_27225,N_29955);
and UO_1445 (O_1445,N_28347,N_28520);
or UO_1446 (O_1446,N_26649,N_27674);
or UO_1447 (O_1447,N_26439,N_25854);
nand UO_1448 (O_1448,N_29675,N_26775);
nor UO_1449 (O_1449,N_29917,N_25072);
and UO_1450 (O_1450,N_27354,N_26359);
and UO_1451 (O_1451,N_27494,N_26901);
and UO_1452 (O_1452,N_26712,N_27191);
and UO_1453 (O_1453,N_25529,N_29856);
or UO_1454 (O_1454,N_29017,N_29477);
nor UO_1455 (O_1455,N_27315,N_29991);
nor UO_1456 (O_1456,N_28109,N_25164);
and UO_1457 (O_1457,N_26082,N_25158);
nor UO_1458 (O_1458,N_25210,N_29736);
and UO_1459 (O_1459,N_27127,N_28969);
or UO_1460 (O_1460,N_25444,N_28549);
nor UO_1461 (O_1461,N_28074,N_27140);
xor UO_1462 (O_1462,N_28486,N_28955);
xnor UO_1463 (O_1463,N_28640,N_27802);
and UO_1464 (O_1464,N_27759,N_27420);
or UO_1465 (O_1465,N_26506,N_29701);
and UO_1466 (O_1466,N_25930,N_29132);
nor UO_1467 (O_1467,N_26342,N_25659);
nor UO_1468 (O_1468,N_27575,N_27700);
nand UO_1469 (O_1469,N_26274,N_26346);
nor UO_1470 (O_1470,N_28830,N_26800);
or UO_1471 (O_1471,N_26055,N_29737);
nor UO_1472 (O_1472,N_28247,N_28582);
nand UO_1473 (O_1473,N_26212,N_25046);
nand UO_1474 (O_1474,N_27326,N_27360);
or UO_1475 (O_1475,N_26977,N_29208);
or UO_1476 (O_1476,N_25649,N_29339);
or UO_1477 (O_1477,N_27116,N_28592);
nand UO_1478 (O_1478,N_26567,N_29287);
nor UO_1479 (O_1479,N_27081,N_26190);
nor UO_1480 (O_1480,N_29413,N_29804);
and UO_1481 (O_1481,N_26690,N_29019);
nand UO_1482 (O_1482,N_29336,N_27425);
xor UO_1483 (O_1483,N_25064,N_27125);
xnor UO_1484 (O_1484,N_28332,N_28394);
or UO_1485 (O_1485,N_25500,N_28767);
xor UO_1486 (O_1486,N_27806,N_25940);
and UO_1487 (O_1487,N_27358,N_27380);
nand UO_1488 (O_1488,N_28707,N_28543);
or UO_1489 (O_1489,N_25713,N_25589);
or UO_1490 (O_1490,N_27611,N_25817);
and UO_1491 (O_1491,N_27030,N_27415);
nand UO_1492 (O_1492,N_28968,N_29247);
xnor UO_1493 (O_1493,N_26306,N_25520);
or UO_1494 (O_1494,N_26244,N_28965);
nand UO_1495 (O_1495,N_27029,N_27204);
and UO_1496 (O_1496,N_26930,N_25499);
nand UO_1497 (O_1497,N_28261,N_28489);
or UO_1498 (O_1498,N_26636,N_27040);
xnor UO_1499 (O_1499,N_26673,N_28905);
and UO_1500 (O_1500,N_29572,N_27798);
and UO_1501 (O_1501,N_29149,N_29138);
nand UO_1502 (O_1502,N_26754,N_25162);
nand UO_1503 (O_1503,N_28002,N_27766);
nor UO_1504 (O_1504,N_27119,N_27971);
or UO_1505 (O_1505,N_28913,N_28459);
nand UO_1506 (O_1506,N_28431,N_28028);
nand UO_1507 (O_1507,N_27260,N_25440);
or UO_1508 (O_1508,N_26070,N_28122);
nor UO_1509 (O_1509,N_28478,N_29376);
and UO_1510 (O_1510,N_28573,N_28626);
nand UO_1511 (O_1511,N_25464,N_26988);
and UO_1512 (O_1512,N_27300,N_25950);
nor UO_1513 (O_1513,N_27592,N_28250);
and UO_1514 (O_1514,N_27939,N_26675);
or UO_1515 (O_1515,N_27387,N_29753);
nor UO_1516 (O_1516,N_25456,N_26918);
xor UO_1517 (O_1517,N_26458,N_25860);
xnor UO_1518 (O_1518,N_26247,N_28886);
or UO_1519 (O_1519,N_27259,N_27272);
and UO_1520 (O_1520,N_25362,N_26559);
nor UO_1521 (O_1521,N_28687,N_29690);
and UO_1522 (O_1522,N_28418,N_29654);
nor UO_1523 (O_1523,N_29032,N_26990);
nor UO_1524 (O_1524,N_28363,N_28641);
and UO_1525 (O_1525,N_29883,N_26756);
nand UO_1526 (O_1526,N_29728,N_26275);
or UO_1527 (O_1527,N_29143,N_26702);
nand UO_1528 (O_1528,N_27831,N_29349);
nor UO_1529 (O_1529,N_26224,N_25438);
or UO_1530 (O_1530,N_25850,N_26461);
or UO_1531 (O_1531,N_28613,N_29312);
nand UO_1532 (O_1532,N_28303,N_26710);
nand UO_1533 (O_1533,N_27636,N_27606);
or UO_1534 (O_1534,N_25848,N_29845);
and UO_1535 (O_1535,N_27540,N_25981);
and UO_1536 (O_1536,N_25287,N_28040);
xor UO_1537 (O_1537,N_28078,N_25597);
nor UO_1538 (O_1538,N_26483,N_27527);
and UO_1539 (O_1539,N_25100,N_27123);
xnor UO_1540 (O_1540,N_25693,N_26826);
or UO_1541 (O_1541,N_28879,N_26547);
nor UO_1542 (O_1542,N_25363,N_28115);
nand UO_1543 (O_1543,N_26985,N_27462);
nand UO_1544 (O_1544,N_27245,N_27148);
and UO_1545 (O_1545,N_28237,N_25936);
and UO_1546 (O_1546,N_29382,N_27033);
and UO_1547 (O_1547,N_25184,N_26729);
xor UO_1548 (O_1548,N_27091,N_26404);
nand UO_1549 (O_1549,N_27506,N_28755);
nor UO_1550 (O_1550,N_28888,N_29670);
xnor UO_1551 (O_1551,N_28698,N_29011);
nor UO_1552 (O_1552,N_27825,N_29489);
nand UO_1553 (O_1553,N_25601,N_27344);
or UO_1554 (O_1554,N_27401,N_25878);
xor UO_1555 (O_1555,N_29291,N_29085);
nor UO_1556 (O_1556,N_29289,N_25038);
xnor UO_1557 (O_1557,N_28321,N_26850);
xor UO_1558 (O_1558,N_25315,N_27786);
and UO_1559 (O_1559,N_26889,N_25406);
and UO_1560 (O_1560,N_27676,N_27230);
nand UO_1561 (O_1561,N_28442,N_29416);
or UO_1562 (O_1562,N_29989,N_28308);
and UO_1563 (O_1563,N_25881,N_26472);
and UO_1564 (O_1564,N_27343,N_29609);
xnor UO_1565 (O_1565,N_27201,N_25908);
or UO_1566 (O_1566,N_26065,N_25782);
xor UO_1567 (O_1567,N_28403,N_26330);
xnor UO_1568 (O_1568,N_25146,N_28977);
nor UO_1569 (O_1569,N_27333,N_25921);
or UO_1570 (O_1570,N_26814,N_28947);
nand UO_1571 (O_1571,N_29069,N_28209);
xor UO_1572 (O_1572,N_26637,N_25771);
and UO_1573 (O_1573,N_27981,N_25581);
nor UO_1574 (O_1574,N_25387,N_25424);
nand UO_1575 (O_1575,N_25453,N_25776);
xnor UO_1576 (O_1576,N_25727,N_27439);
and UO_1577 (O_1577,N_26122,N_26862);
or UO_1578 (O_1578,N_27995,N_29448);
nor UO_1579 (O_1579,N_27566,N_27153);
xnor UO_1580 (O_1580,N_26433,N_28228);
xor UO_1581 (O_1581,N_28165,N_29071);
and UO_1582 (O_1582,N_26768,N_25282);
xor UO_1583 (O_1583,N_28335,N_28827);
nand UO_1584 (O_1584,N_25251,N_28134);
or UO_1585 (O_1585,N_25679,N_28733);
and UO_1586 (O_1586,N_25163,N_25984);
and UO_1587 (O_1587,N_27329,N_27408);
nor UO_1588 (O_1588,N_26934,N_27146);
or UO_1589 (O_1589,N_29187,N_29745);
nor UO_1590 (O_1590,N_28736,N_27834);
or UO_1591 (O_1591,N_29344,N_29780);
and UO_1592 (O_1592,N_27613,N_25258);
xor UO_1593 (O_1593,N_26171,N_26528);
and UO_1594 (O_1594,N_27649,N_28944);
and UO_1595 (O_1595,N_29027,N_29854);
nor UO_1596 (O_1596,N_25191,N_29740);
or UO_1597 (O_1597,N_29148,N_28937);
xor UO_1598 (O_1598,N_25052,N_26821);
xnor UO_1599 (O_1599,N_25916,N_26585);
xor UO_1600 (O_1600,N_28572,N_27255);
nor UO_1601 (O_1601,N_29342,N_26961);
or UO_1602 (O_1602,N_25150,N_27475);
nand UO_1603 (O_1603,N_26041,N_25608);
xnor UO_1604 (O_1604,N_26619,N_28068);
xnor UO_1605 (O_1605,N_26494,N_26907);
and UO_1606 (O_1606,N_25410,N_28208);
nand UO_1607 (O_1607,N_29517,N_28021);
xor UO_1608 (O_1608,N_27144,N_29365);
or UO_1609 (O_1609,N_27283,N_26271);
xor UO_1610 (O_1610,N_29625,N_25733);
nor UO_1611 (O_1611,N_29157,N_25266);
xor UO_1612 (O_1612,N_25227,N_27671);
nor UO_1613 (O_1613,N_25995,N_28116);
xnor UO_1614 (O_1614,N_28272,N_29101);
nor UO_1615 (O_1615,N_26440,N_26580);
and UO_1616 (O_1616,N_25480,N_28591);
and UO_1617 (O_1617,N_27719,N_27712);
nand UO_1618 (O_1618,N_29114,N_26935);
nor UO_1619 (O_1619,N_25177,N_25277);
xor UO_1620 (O_1620,N_29345,N_25030);
and UO_1621 (O_1621,N_27994,N_29200);
xor UO_1622 (O_1622,N_26402,N_29269);
nand UO_1623 (O_1623,N_29614,N_29968);
xnor UO_1624 (O_1624,N_28410,N_26419);
nand UO_1625 (O_1625,N_26179,N_26525);
or UO_1626 (O_1626,N_28704,N_26069);
and UO_1627 (O_1627,N_26778,N_29481);
or UO_1628 (O_1628,N_27843,N_29077);
nand UO_1629 (O_1629,N_29543,N_29099);
xor UO_1630 (O_1630,N_25723,N_29328);
and UO_1631 (O_1631,N_27447,N_26144);
xor UO_1632 (O_1632,N_25037,N_27107);
and UO_1633 (O_1633,N_26533,N_27218);
or UO_1634 (O_1634,N_25443,N_25795);
or UO_1635 (O_1635,N_28164,N_27906);
xor UO_1636 (O_1636,N_28302,N_26076);
nand UO_1637 (O_1637,N_28758,N_28665);
or UO_1638 (O_1638,N_27240,N_26663);
nand UO_1639 (O_1639,N_29665,N_28730);
or UO_1640 (O_1640,N_25065,N_25900);
nand UO_1641 (O_1641,N_27414,N_26513);
xor UO_1642 (O_1642,N_28839,N_29380);
and UO_1643 (O_1643,N_25945,N_26912);
and UO_1644 (O_1644,N_28820,N_26687);
or UO_1645 (O_1645,N_27101,N_25120);
xor UO_1646 (O_1646,N_28323,N_25765);
xnor UO_1647 (O_1647,N_25768,N_28392);
nor UO_1648 (O_1648,N_25752,N_27388);
and UO_1649 (O_1649,N_29571,N_29831);
nand UO_1650 (O_1650,N_28889,N_29685);
nor UO_1651 (O_1651,N_26343,N_28542);
nand UO_1652 (O_1652,N_26121,N_27365);
xnor UO_1653 (O_1653,N_28759,N_26874);
nand UO_1654 (O_1654,N_25924,N_26872);
nand UO_1655 (O_1655,N_26784,N_28979);
xor UO_1656 (O_1656,N_25705,N_28873);
nand UO_1657 (O_1657,N_25208,N_29255);
nand UO_1658 (O_1658,N_26392,N_25882);
xor UO_1659 (O_1659,N_29928,N_28366);
nor UO_1660 (O_1660,N_27770,N_27874);
and UO_1661 (O_1661,N_27026,N_29326);
nand UO_1662 (O_1662,N_29404,N_29039);
xnor UO_1663 (O_1663,N_29023,N_27803);
or UO_1664 (O_1664,N_28786,N_29796);
nand UO_1665 (O_1665,N_25944,N_26923);
xnor UO_1666 (O_1666,N_27755,N_28064);
xor UO_1667 (O_1667,N_25617,N_29616);
and UO_1668 (O_1668,N_28373,N_27036);
and UO_1669 (O_1669,N_25033,N_27957);
nand UO_1670 (O_1670,N_28581,N_29992);
xnor UO_1671 (O_1671,N_29351,N_28488);
nor UO_1672 (O_1672,N_28559,N_27624);
nor UO_1673 (O_1673,N_28929,N_26646);
nor UO_1674 (O_1674,N_27419,N_29444);
or UO_1675 (O_1675,N_25031,N_27965);
xor UO_1676 (O_1676,N_28346,N_29364);
nor UO_1677 (O_1677,N_25035,N_26153);
nand UO_1678 (O_1678,N_29700,N_27782);
and UO_1679 (O_1679,N_25171,N_26873);
xor UO_1680 (O_1680,N_28961,N_25190);
or UO_1681 (O_1681,N_26700,N_26880);
and UO_1682 (O_1682,N_26385,N_25799);
xor UO_1683 (O_1683,N_27496,N_26788);
nand UO_1684 (O_1684,N_25622,N_27710);
or UO_1685 (O_1685,N_26123,N_28659);
xor UO_1686 (O_1686,N_27353,N_28829);
xor UO_1687 (O_1687,N_27635,N_27039);
xor UO_1688 (O_1688,N_26164,N_29335);
nand UO_1689 (O_1689,N_28380,N_25722);
or UO_1690 (O_1690,N_29014,N_29990);
and UO_1691 (O_1691,N_28997,N_27381);
nor UO_1692 (O_1692,N_26096,N_26202);
nand UO_1693 (O_1693,N_25276,N_27050);
xnor UO_1694 (O_1694,N_29639,N_27677);
nand UO_1695 (O_1695,N_25346,N_25931);
nand UO_1696 (O_1696,N_27591,N_29230);
or UO_1697 (O_1697,N_28526,N_27749);
nor UO_1698 (O_1698,N_27977,N_26027);
xor UO_1699 (O_1699,N_27077,N_25436);
nor UO_1700 (O_1700,N_26277,N_25784);
nor UO_1701 (O_1701,N_29356,N_29880);
and UO_1702 (O_1702,N_28590,N_25159);
nand UO_1703 (O_1703,N_26017,N_25990);
xor UO_1704 (O_1704,N_27714,N_26314);
xnor UO_1705 (O_1705,N_28254,N_25837);
nand UO_1706 (O_1706,N_28159,N_27431);
nor UO_1707 (O_1707,N_27241,N_27276);
nor UO_1708 (O_1708,N_25117,N_26944);
xnor UO_1709 (O_1709,N_25205,N_29611);
or UO_1710 (O_1710,N_25588,N_25584);
xnor UO_1711 (O_1711,N_27956,N_28256);
and UO_1712 (O_1712,N_28047,N_27219);
or UO_1713 (O_1713,N_25913,N_26143);
nor UO_1714 (O_1714,N_28633,N_26272);
nor UO_1715 (O_1715,N_27368,N_27974);
or UO_1716 (O_1716,N_26925,N_29683);
xor UO_1717 (O_1717,N_27109,N_28378);
nor UO_1718 (O_1718,N_27601,N_26131);
and UO_1719 (O_1719,N_26750,N_28038);
and UO_1720 (O_1720,N_25478,N_26887);
xnor UO_1721 (O_1721,N_29769,N_29043);
or UO_1722 (O_1722,N_25024,N_28460);
xnor UO_1723 (O_1723,N_25643,N_29102);
and UO_1724 (O_1724,N_27363,N_26371);
nor UO_1725 (O_1725,N_26490,N_25076);
nor UO_1726 (O_1726,N_29515,N_26824);
nand UO_1727 (O_1727,N_25974,N_28966);
nand UO_1728 (O_1728,N_26780,N_26060);
nand UO_1729 (O_1729,N_29066,N_25690);
and UO_1730 (O_1730,N_27067,N_29983);
nor UO_1731 (O_1731,N_26858,N_28617);
nand UO_1732 (O_1732,N_28429,N_25070);
nand UO_1733 (O_1733,N_27229,N_26167);
nand UO_1734 (O_1734,N_28854,N_28835);
nand UO_1735 (O_1735,N_29202,N_25122);
or UO_1736 (O_1736,N_29523,N_28841);
nand UO_1737 (O_1737,N_25743,N_25022);
nor UO_1738 (O_1738,N_28023,N_28917);
xor UO_1739 (O_1739,N_29070,N_26305);
and UO_1740 (O_1740,N_29240,N_28602);
nand UO_1741 (O_1741,N_28847,N_27894);
nor UO_1742 (O_1742,N_27082,N_28849);
nand UO_1743 (O_1743,N_26279,N_25983);
nor UO_1744 (O_1744,N_26048,N_26012);
nand UO_1745 (O_1745,N_28390,N_29386);
nor UO_1746 (O_1746,N_28587,N_29218);
and UO_1747 (O_1747,N_26280,N_25103);
nand UO_1748 (O_1748,N_25747,N_29271);
or UO_1749 (O_1749,N_27324,N_25255);
nand UO_1750 (O_1750,N_28695,N_25741);
xnor UO_1751 (O_1751,N_27070,N_26016);
xnor UO_1752 (O_1752,N_27890,N_27281);
and UO_1753 (O_1753,N_27097,N_28596);
xnor UO_1754 (O_1754,N_25764,N_29813);
nor UO_1755 (O_1755,N_29446,N_25963);
nor UO_1756 (O_1756,N_27117,N_27924);
or UO_1757 (O_1757,N_28398,N_26094);
nand UO_1758 (O_1758,N_25364,N_25910);
nand UO_1759 (O_1759,N_29935,N_28018);
nor UO_1760 (O_1760,N_29399,N_28067);
xor UO_1761 (O_1761,N_25791,N_28850);
nand UO_1762 (O_1762,N_29681,N_27446);
nor UO_1763 (O_1763,N_27352,N_28579);
nand UO_1764 (O_1764,N_27052,N_29920);
or UO_1765 (O_1765,N_29710,N_25042);
or UO_1766 (O_1766,N_27561,N_28731);
xor UO_1767 (O_1767,N_27821,N_28760);
nor UO_1768 (O_1768,N_25169,N_25989);
nor UO_1769 (O_1769,N_27143,N_28092);
nand UO_1770 (O_1770,N_27385,N_25054);
or UO_1771 (O_1771,N_25341,N_26564);
or UO_1772 (O_1772,N_29480,N_28477);
xnor UO_1773 (O_1773,N_27093,N_26047);
nand UO_1774 (O_1774,N_29219,N_26273);
nand UO_1775 (O_1775,N_28006,N_26665);
nand UO_1776 (O_1776,N_29073,N_27302);
nor UO_1777 (O_1777,N_25195,N_26762);
nand UO_1778 (O_1778,N_29911,N_25091);
xor UO_1779 (O_1779,N_26287,N_27233);
and UO_1780 (O_1780,N_28932,N_26013);
and UO_1781 (O_1781,N_25053,N_28570);
nor UO_1782 (O_1782,N_28479,N_26595);
nor UO_1783 (O_1783,N_26558,N_27655);
nor UO_1784 (O_1784,N_27590,N_28344);
xnor UO_1785 (O_1785,N_26956,N_29256);
or UO_1786 (O_1786,N_28892,N_27500);
xor UO_1787 (O_1787,N_28071,N_25861);
nand UO_1788 (O_1788,N_28752,N_29548);
and UO_1789 (O_1789,N_28202,N_25824);
nand UO_1790 (O_1790,N_26672,N_25306);
and UO_1791 (O_1791,N_25960,N_25147);
or UO_1792 (O_1792,N_27633,N_27106);
nand UO_1793 (O_1793,N_29829,N_29050);
nor UO_1794 (O_1794,N_29672,N_27943);
nor UO_1795 (O_1795,N_29746,N_27149);
and UO_1796 (O_1796,N_29977,N_26168);
or UO_1797 (O_1797,N_27778,N_29105);
or UO_1798 (O_1798,N_29258,N_26046);
and UO_1799 (O_1799,N_25451,N_28598);
or UO_1800 (O_1800,N_25627,N_28155);
xor UO_1801 (O_1801,N_29885,N_25384);
and UO_1802 (O_1802,N_27809,N_25918);
or UO_1803 (O_1803,N_27417,N_27377);
xnor UO_1804 (O_1804,N_28552,N_27836);
nor UO_1805 (O_1805,N_27441,N_29324);
or UO_1806 (O_1806,N_29874,N_28674);
or UO_1807 (O_1807,N_25724,N_28962);
or UO_1808 (O_1808,N_28564,N_28290);
nor UO_1809 (O_1809,N_26926,N_25545);
or UO_1810 (O_1810,N_29196,N_26393);
nand UO_1811 (O_1811,N_26847,N_26155);
nand UO_1812 (O_1812,N_26942,N_27173);
nand UO_1813 (O_1813,N_29853,N_28295);
nor UO_1814 (O_1814,N_28643,N_27618);
and UO_1815 (O_1815,N_25976,N_26252);
and UO_1816 (O_1816,N_29346,N_26304);
and UO_1817 (O_1817,N_27320,N_28395);
or UO_1818 (O_1818,N_27554,N_28383);
nand UO_1819 (O_1819,N_26536,N_25680);
nor UO_1820 (O_1820,N_26450,N_29348);
xor UO_1821 (O_1821,N_25825,N_28031);
nor UO_1822 (O_1822,N_26549,N_29462);
and UO_1823 (O_1823,N_26162,N_26787);
nor UO_1824 (O_1824,N_28140,N_25338);
nor UO_1825 (O_1825,N_26302,N_27926);
and UO_1826 (O_1826,N_27334,N_27646);
or UO_1827 (O_1827,N_25907,N_27078);
and UO_1828 (O_1828,N_28471,N_25128);
nand UO_1829 (O_1829,N_26596,N_25005);
xor UO_1830 (O_1830,N_27877,N_25668);
nand UO_1831 (O_1831,N_29120,N_25632);
and UO_1832 (O_1832,N_27944,N_28119);
xnor UO_1833 (O_1833,N_29645,N_28817);
nor UO_1834 (O_1834,N_28522,N_26184);
nand UO_1835 (O_1835,N_26615,N_29599);
xnor UO_1836 (O_1836,N_28894,N_27481);
and UO_1837 (O_1837,N_25807,N_26011);
or UO_1838 (O_1838,N_28312,N_29937);
xnor UO_1839 (O_1839,N_28161,N_26652);
and UO_1840 (O_1840,N_27172,N_26101);
xnor UO_1841 (O_1841,N_28318,N_29197);
nand UO_1842 (O_1842,N_28053,N_26709);
nand UO_1843 (O_1843,N_28848,N_25763);
nand UO_1844 (O_1844,N_28327,N_28940);
nor UO_1845 (O_1845,N_26684,N_29922);
xnor UO_1846 (O_1846,N_25957,N_27936);
nand UO_1847 (O_1847,N_27041,N_27095);
and UO_1848 (O_1848,N_28924,N_26865);
xnor UO_1849 (O_1849,N_27856,N_28405);
nand UO_1850 (O_1850,N_26157,N_28551);
or UO_1851 (O_1851,N_29119,N_25885);
xnor UO_1852 (O_1852,N_29037,N_25466);
xor UO_1853 (O_1853,N_25658,N_26482);
xnor UO_1854 (O_1854,N_25620,N_26924);
xnor UO_1855 (O_1855,N_29999,N_25114);
nand UO_1856 (O_1856,N_29475,N_27340);
and UO_1857 (O_1857,N_26759,N_25239);
xor UO_1858 (O_1858,N_27709,N_28123);
nor UO_1859 (O_1859,N_28976,N_27147);
and UO_1860 (O_1860,N_26644,N_27808);
xor UO_1861 (O_1861,N_26656,N_28553);
or UO_1862 (O_1862,N_25203,N_29784);
nor UO_1863 (O_1863,N_26650,N_28282);
or UO_1864 (O_1864,N_27704,N_25377);
nand UO_1865 (O_1865,N_26263,N_28324);
nor UO_1866 (O_1866,N_28216,N_26954);
or UO_1867 (O_1867,N_25993,N_27725);
nand UO_1868 (O_1868,N_29026,N_25891);
xnor UO_1869 (O_1869,N_28287,N_28599);
xnor UO_1870 (O_1870,N_25874,N_28908);
or UO_1871 (O_1871,N_28773,N_27697);
nand UO_1872 (O_1872,N_27310,N_28355);
xnor UO_1873 (O_1873,N_25400,N_29501);
xor UO_1874 (O_1874,N_26996,N_25598);
nand UO_1875 (O_1875,N_25975,N_25709);
nand UO_1876 (O_1876,N_25358,N_25437);
or UO_1877 (O_1877,N_26399,N_29418);
nor UO_1878 (O_1878,N_25672,N_29347);
nor UO_1879 (O_1879,N_29934,N_28162);
nor UO_1880 (O_1880,N_29995,N_29744);
nor UO_1881 (O_1881,N_26947,N_27145);
nand UO_1882 (O_1882,N_28397,N_27285);
and UO_1883 (O_1883,N_25197,N_27378);
xor UO_1884 (O_1884,N_26195,N_27200);
nor UO_1885 (O_1885,N_29261,N_28608);
nor UO_1886 (O_1886,N_29776,N_29858);
and UO_1887 (O_1887,N_27120,N_29139);
nor UO_1888 (O_1888,N_26337,N_28118);
nand UO_1889 (O_1889,N_25295,N_26995);
or UO_1890 (O_1890,N_27314,N_26486);
or UO_1891 (O_1891,N_26220,N_26006);
xor UO_1892 (O_1892,N_27128,N_27322);
or UO_1893 (O_1893,N_28722,N_29169);
xnor UO_1894 (O_1894,N_29165,N_29606);
or UO_1895 (O_1895,N_27607,N_28831);
or UO_1896 (O_1896,N_29891,N_25663);
nand UO_1897 (O_1897,N_29802,N_25193);
nand UO_1898 (O_1898,N_25228,N_26206);
nand UO_1899 (O_1899,N_26207,N_28178);
and UO_1900 (O_1900,N_25987,N_25246);
or UO_1901 (O_1901,N_27653,N_28868);
or UO_1902 (O_1902,N_27785,N_26617);
nor UO_1903 (O_1903,N_25796,N_27126);
xnor UO_1904 (O_1904,N_28627,N_25797);
xnor UO_1905 (O_1905,N_26038,N_29916);
or UO_1906 (O_1906,N_29822,N_29993);
xnor UO_1907 (O_1907,N_25644,N_28644);
or UO_1908 (O_1908,N_27286,N_29361);
or UO_1909 (O_1909,N_26534,N_27290);
and UO_1910 (O_1910,N_26648,N_28655);
nand UO_1911 (O_1911,N_28706,N_27501);
xor UO_1912 (O_1912,N_29500,N_28433);
nor UO_1913 (O_1913,N_26723,N_28331);
xnor UO_1914 (O_1914,N_27409,N_25378);
nand UO_1915 (O_1915,N_29930,N_28938);
or UO_1916 (O_1916,N_26294,N_27861);
nand UO_1917 (O_1917,N_28493,N_28249);
nor UO_1918 (O_1918,N_26291,N_28233);
or UO_1919 (O_1919,N_28371,N_27392);
or UO_1920 (O_1920,N_27311,N_29846);
xor UO_1921 (O_1921,N_28569,N_27312);
xnor UO_1922 (O_1922,N_28154,N_25553);
and UO_1923 (O_1923,N_26653,N_29397);
or UO_1924 (O_1924,N_29721,N_25836);
nor UO_1925 (O_1925,N_27293,N_28796);
or UO_1926 (O_1926,N_26208,N_29815);
and UO_1927 (O_1927,N_26969,N_26050);
nor UO_1928 (O_1928,N_29355,N_26891);
nand UO_1929 (O_1929,N_26898,N_29152);
nand UO_1930 (O_1930,N_25461,N_26080);
or UO_1931 (O_1931,N_27668,N_28089);
and UO_1932 (O_1932,N_25912,N_25133);
or UO_1933 (O_1933,N_26193,N_26515);
nor UO_1934 (O_1934,N_25800,N_29235);
and UO_1935 (O_1935,N_29958,N_26582);
nor UO_1936 (O_1936,N_27764,N_27376);
xnor UO_1937 (O_1937,N_26315,N_27557);
and UO_1938 (O_1938,N_28789,N_26783);
nor UO_1939 (O_1939,N_25223,N_28032);
nand UO_1940 (O_1940,N_29203,N_26386);
nor UO_1941 (O_1941,N_26991,N_25067);
and UO_1942 (O_1942,N_26902,N_26185);
xor UO_1943 (O_1943,N_25801,N_28090);
or UO_1944 (O_1944,N_28107,N_27402);
nor UO_1945 (O_1945,N_27711,N_27357);
nor UO_1946 (O_1946,N_27410,N_29876);
xor UO_1947 (O_1947,N_26074,N_29381);
or UO_1948 (O_1948,N_27202,N_29805);
xnor UO_1949 (O_1949,N_27339,N_28084);
and UO_1950 (O_1950,N_28732,N_29082);
nand UO_1951 (O_1951,N_25818,N_25901);
nor UO_1952 (O_1952,N_29785,N_26158);
nor UO_1953 (O_1953,N_26639,N_29038);
xor UO_1954 (O_1954,N_29167,N_29511);
xnor UO_1955 (O_1955,N_25725,N_25043);
xnor UO_1956 (O_1956,N_25157,N_26284);
or UO_1957 (O_1957,N_27379,N_28837);
or UO_1958 (O_1958,N_25775,N_27641);
nand UO_1959 (O_1959,N_29007,N_25844);
xnor UO_1960 (O_1960,N_29253,N_29061);
or UO_1961 (O_1961,N_26095,N_28197);
nand UO_1962 (O_1962,N_25301,N_25056);
xor UO_1963 (O_1963,N_28753,N_26739);
or UO_1964 (O_1964,N_26602,N_28389);
or UO_1965 (O_1965,N_26692,N_27102);
nor UO_1966 (O_1966,N_28609,N_25248);
or UO_1967 (O_1967,N_26910,N_25564);
and UO_1968 (O_1968,N_27963,N_25962);
xnor UO_1969 (O_1969,N_27242,N_27960);
and UO_1970 (O_1970,N_27562,N_28113);
xnor UO_1971 (O_1971,N_29001,N_25261);
nor UO_1972 (O_1972,N_25636,N_25345);
nor UO_1973 (O_1973,N_25746,N_27435);
and UO_1974 (O_1974,N_27084,N_26381);
nor UO_1975 (O_1975,N_26507,N_26608);
or UO_1976 (O_1976,N_29129,N_25607);
xor UO_1977 (O_1977,N_29373,N_28832);
and UO_1978 (O_1978,N_25317,N_26052);
nor UO_1979 (O_1979,N_28776,N_26383);
nand UO_1980 (O_1980,N_28978,N_28780);
or UO_1981 (O_1981,N_29932,N_27182);
or UO_1982 (O_1982,N_27824,N_28077);
or UO_1983 (O_1983,N_25112,N_26763);
and UO_1984 (O_1984,N_29064,N_26772);
nor UO_1985 (O_1985,N_27413,N_28386);
and UO_1986 (O_1986,N_27342,N_27973);
and UO_1987 (O_1987,N_25490,N_25585);
nor UO_1988 (O_1988,N_28419,N_25847);
or UO_1989 (O_1989,N_29975,N_29875);
nand UO_1990 (O_1990,N_28600,N_27542);
and UO_1991 (O_1991,N_25740,N_27359);
and UO_1992 (O_1992,N_28269,N_28343);
and UO_1993 (O_1993,N_25549,N_26974);
nor UO_1994 (O_1994,N_27005,N_27914);
nand UO_1995 (O_1995,N_25333,N_27003);
and UO_1996 (O_1996,N_28601,N_26015);
xor UO_1997 (O_1997,N_25512,N_26950);
and UO_1998 (O_1998,N_25127,N_27531);
xnor UO_1999 (O_1999,N_25253,N_26782);
or UO_2000 (O_2000,N_29390,N_26634);
and UO_2001 (O_2001,N_25115,N_27865);
and UO_2002 (O_2002,N_26660,N_29761);
nor UO_2003 (O_2003,N_26720,N_27031);
and UO_2004 (O_2004,N_27108,N_29576);
or UO_2005 (O_2005,N_25828,N_28629);
and UO_2006 (O_2006,N_29422,N_27823);
nor UO_2007 (O_2007,N_26398,N_25685);
and UO_2008 (O_2008,N_25667,N_29163);
or UO_2009 (O_2009,N_25126,N_28057);
and UO_2010 (O_2010,N_26929,N_28690);
and UO_2011 (O_2011,N_25753,N_27927);
and UO_2012 (O_2012,N_25467,N_28852);
and UO_2013 (O_2013,N_29330,N_25392);
or UO_2014 (O_2014,N_25555,N_26659);
or UO_2015 (O_2015,N_26697,N_26604);
and UO_2016 (O_2016,N_27581,N_27983);
and UO_2017 (O_2017,N_25474,N_26760);
and UO_2018 (O_2018,N_29234,N_28515);
and UO_2019 (O_2019,N_29659,N_26857);
nand UO_2020 (O_2020,N_27848,N_25829);
nand UO_2021 (O_2021,N_29541,N_27319);
xnor UO_2022 (O_2022,N_28680,N_27657);
nor UO_2023 (O_2023,N_25186,N_27849);
nor UO_2024 (O_2024,N_28434,N_26281);
nor UO_2025 (O_2025,N_28325,N_26307);
or UO_2026 (O_2026,N_28846,N_28636);
nor UO_2027 (O_2027,N_27693,N_29303);
xor UO_2028 (O_2028,N_28699,N_29315);
and UO_2029 (O_2029,N_29180,N_26223);
nand UO_2030 (O_2030,N_27911,N_26916);
xor UO_2031 (O_2031,N_26351,N_29633);
xnor UO_2032 (O_2032,N_27743,N_26825);
nand UO_2033 (O_2033,N_25506,N_27389);
nor UO_2034 (O_2034,N_27552,N_29597);
xor UO_2035 (O_2035,N_27056,N_29223);
xor UO_2036 (O_2036,N_26414,N_25044);
and UO_2037 (O_2037,N_27461,N_27972);
and UO_2038 (O_2038,N_26770,N_26899);
and UO_2039 (O_2039,N_26312,N_26413);
xnor UO_2040 (O_2040,N_29311,N_28379);
nand UO_2041 (O_2041,N_26003,N_25884);
xor UO_2042 (O_2042,N_26566,N_25331);
or UO_2043 (O_2043,N_29729,N_28217);
or UO_2044 (O_2044,N_27814,N_26537);
nand UO_2045 (O_2045,N_27403,N_29350);
nor UO_2046 (O_2046,N_26751,N_27541);
nor UO_2047 (O_2047,N_29532,N_26972);
or UO_2048 (O_2048,N_28823,N_29764);
xnor UO_2049 (O_2049,N_25613,N_29810);
or UO_2050 (O_2050,N_28270,N_29629);
or UO_2051 (O_2051,N_27156,N_27092);
or UO_2052 (O_2052,N_28692,N_25448);
nand UO_2053 (O_2053,N_26372,N_25831);
nor UO_2054 (O_2054,N_25926,N_29204);
xnor UO_2055 (O_2055,N_27799,N_29919);
or UO_2056 (O_2056,N_26747,N_26454);
nor UO_2057 (O_2057,N_29586,N_26909);
nor UO_2058 (O_2058,N_26110,N_25998);
nand UO_2059 (O_2059,N_25641,N_27361);
nand UO_2060 (O_2060,N_28499,N_28145);
or UO_2061 (O_2061,N_28170,N_25051);
xor UO_2062 (O_2062,N_26701,N_28851);
nand UO_2063 (O_2063,N_29048,N_27167);
or UO_2064 (O_2064,N_26408,N_27421);
and UO_2065 (O_2065,N_28798,N_26922);
xnor UO_2066 (O_2066,N_26338,N_27266);
or UO_2067 (O_2067,N_26447,N_29392);
nor UO_2068 (O_2068,N_28062,N_27767);
and UO_2069 (O_2069,N_27583,N_28274);
nor UO_2070 (O_2070,N_29453,N_25580);
and UO_2071 (O_2071,N_28422,N_28326);
or UO_2072 (O_2072,N_27837,N_27812);
nand UO_2073 (O_2073,N_28491,N_26859);
and UO_2074 (O_2074,N_29936,N_28151);
xor UO_2075 (O_2075,N_25846,N_25367);
xnor UO_2076 (O_2076,N_26728,N_28876);
and UO_2077 (O_2077,N_27670,N_25278);
or UO_2078 (O_2078,N_29325,N_27539);
nand UO_2079 (O_2079,N_28035,N_29409);
or UO_2080 (O_2080,N_26234,N_26647);
or UO_2081 (O_2081,N_25339,N_27228);
and UO_2082 (O_2082,N_29965,N_25754);
or UO_2083 (O_2083,N_26467,N_25271);
nor UO_2084 (O_2084,N_29320,N_26009);
nor UO_2085 (O_2085,N_29857,N_26218);
nor UO_2086 (O_2086,N_25573,N_26597);
and UO_2087 (O_2087,N_28294,N_28801);
xnor UO_2088 (O_2088,N_29587,N_26848);
xor UO_2089 (O_2089,N_27997,N_28819);
or UO_2090 (O_2090,N_28382,N_28464);
nor UO_2091 (O_2091,N_25090,N_28281);
nor UO_2092 (O_2092,N_25148,N_25014);
xnor UO_2093 (O_2093,N_29244,N_28063);
and UO_2094 (O_2094,N_25933,N_25342);
nand UO_2095 (O_2095,N_29762,N_25420);
and UO_2096 (O_2096,N_25408,N_26496);
and UO_2097 (O_2097,N_25838,N_27489);
nor UO_2098 (O_2098,N_25956,N_29655);
or UO_2099 (O_2099,N_27001,N_29903);
nor UO_2100 (O_2100,N_29264,N_27787);
or UO_2101 (O_2101,N_29505,N_26588);
nand UO_2102 (O_2102,N_26072,N_29634);
and UO_2103 (O_2103,N_28328,N_29799);
nand UO_2104 (O_2104,N_26831,N_27945);
nor UO_2105 (O_2105,N_26339,N_29140);
nand UO_2106 (O_2106,N_26696,N_25452);
and UO_2107 (O_2107,N_28440,N_25326);
and UO_2108 (O_2108,N_25283,N_25623);
nor UO_2109 (O_2109,N_27051,N_27918);
nand UO_2110 (O_2110,N_25224,N_29438);
nand UO_2111 (O_2111,N_25582,N_27362);
or UO_2112 (O_2112,N_26621,N_27129);
xnor UO_2113 (O_2113,N_27669,N_26364);
or UO_2114 (O_2114,N_25721,N_28286);
xnor UO_2115 (O_2115,N_28330,N_29679);
nand UO_2116 (O_2116,N_26601,N_29584);
or UO_2117 (O_2117,N_25965,N_28610);
and UO_2118 (O_2118,N_25600,N_29445);
or UO_2119 (O_2119,N_28271,N_28443);
or UO_2120 (O_2120,N_27321,N_25118);
and UO_2121 (O_2121,N_25843,N_25353);
nor UO_2122 (O_2122,N_29674,N_27076);
xor UO_2123 (O_2123,N_25482,N_25249);
and UO_2124 (O_2124,N_28577,N_28996);
and UO_2125 (O_2125,N_29695,N_28523);
or UO_2126 (O_2126,N_27243,N_26322);
nand UO_2127 (O_2127,N_25206,N_26903);
nor UO_2128 (O_2128,N_28967,N_26791);
or UO_2129 (O_2129,N_27014,N_27337);
xnor UO_2130 (O_2130,N_27304,N_27318);
nor UO_2131 (O_2131,N_26235,N_25745);
nand UO_2132 (O_2132,N_26115,N_27269);
or UO_2133 (O_2133,N_26463,N_25676);
nor UO_2134 (O_2134,N_29600,N_29188);
nand UO_2135 (O_2135,N_26492,N_28142);
nor UO_2136 (O_2136,N_25089,N_27822);
and UO_2137 (O_2137,N_25917,N_26999);
or UO_2138 (O_2138,N_27951,N_26250);
or UO_2139 (O_2139,N_29507,N_25744);
or UO_2140 (O_2140,N_25786,N_28508);
or UO_2141 (O_2141,N_26051,N_27301);
xnor UO_2142 (O_2142,N_28768,N_27297);
or UO_2143 (O_2143,N_25832,N_29942);
nor UO_2144 (O_2144,N_28186,N_25422);
xnor UO_2145 (O_2145,N_26476,N_25074);
xnor UO_2146 (O_2146,N_28213,N_26460);
or UO_2147 (O_2147,N_26860,N_28015);
nor UO_2148 (O_2148,N_28083,N_25041);
xnor UO_2149 (O_2149,N_28361,N_28757);
or UO_2150 (O_2150,N_29141,N_29452);
xor UO_2151 (O_2151,N_26232,N_26261);
nor UO_2152 (O_2152,N_28547,N_26530);
or UO_2153 (O_2153,N_28914,N_27526);
xnor UO_2154 (O_2154,N_29963,N_26877);
or UO_2155 (O_2155,N_25508,N_26415);
nand UO_2156 (O_2156,N_26410,N_25586);
and UO_2157 (O_2157,N_25369,N_28341);
and UO_2158 (O_2158,N_29028,N_27978);
nor UO_2159 (O_2159,N_27284,N_29703);
and UO_2160 (O_2160,N_26577,N_25397);
xor UO_2161 (O_2161,N_28930,N_27341);
nand UO_2162 (O_2162,N_29951,N_28815);
or UO_2163 (O_2163,N_27390,N_26384);
nand UO_2164 (O_2164,N_28235,N_29299);
nand UO_2165 (O_2165,N_28385,N_29573);
and UO_2166 (O_2166,N_26732,N_25399);
and UO_2167 (O_2167,N_29768,N_29210);
nor UO_2168 (O_2168,N_28806,N_25864);
or UO_2169 (O_2169,N_27728,N_29697);
or UO_2170 (O_2170,N_27330,N_28676);
xnor UO_2171 (O_2171,N_27134,N_28258);
xor UO_2172 (O_2172,N_28487,N_26125);
nor UO_2173 (O_2173,N_26845,N_26512);
nor UO_2174 (O_2174,N_28280,N_25762);
nor UO_2175 (O_2175,N_25412,N_28536);
or UO_2176 (O_2176,N_29305,N_27555);
and UO_2177 (O_2177,N_27317,N_26396);
or UO_2178 (O_2178,N_28878,N_25999);
nor UO_2179 (O_2179,N_29012,N_29454);
nor UO_2180 (O_2180,N_28778,N_25699);
or UO_2181 (O_2181,N_28019,N_26508);
xor UO_2182 (O_2182,N_27909,N_28288);
or UO_2183 (O_2183,N_28951,N_27351);
or UO_2184 (O_2184,N_25937,N_25979);
xor UO_2185 (O_2185,N_28013,N_25314);
or UO_2186 (O_2186,N_28425,N_28374);
nor UO_2187 (O_2187,N_25536,N_29754);
nor UO_2188 (O_2188,N_26655,N_29758);
nand UO_2189 (O_2189,N_29274,N_26678);
nor UO_2190 (O_2190,N_29384,N_25731);
and UO_2191 (O_2191,N_26238,N_29047);
or UO_2192 (O_2192,N_29075,N_27628);
xnor UO_2193 (O_2193,N_28352,N_28480);
or UO_2194 (O_2194,N_25105,N_25025);
and UO_2195 (O_2195,N_26569,N_28278);
nor UO_2196 (O_2196,N_27113,N_25562);
nand UO_2197 (O_2197,N_28939,N_29096);
xor UO_2198 (O_2198,N_29525,N_25405);
and UO_2199 (O_2199,N_25008,N_28921);
nor UO_2200 (O_2200,N_27622,N_27463);
xnor UO_2201 (O_2201,N_28415,N_29147);
and UO_2202 (O_2202,N_28152,N_25435);
nor UO_2203 (O_2203,N_25686,N_28638);
nor UO_2204 (O_2204,N_27295,N_28833);
xnor UO_2205 (O_2205,N_27404,N_25568);
xor UO_2206 (O_2206,N_25321,N_28227);
or UO_2207 (O_2207,N_29029,N_28494);
nand UO_2208 (O_2208,N_26695,N_27867);
or UO_2209 (O_2209,N_25288,N_25160);
nor UO_2210 (O_2210,N_25559,N_26264);
or UO_2211 (O_2211,N_29425,N_27616);
nand UO_2212 (O_2212,N_27872,N_29801);
xor UO_2213 (O_2213,N_29627,N_28370);
nand UO_2214 (O_2214,N_28588,N_27519);
nor UO_2215 (O_2215,N_27087,N_25648);
or UO_2216 (O_2216,N_29786,N_27131);
and UO_2217 (O_2217,N_29160,N_29793);
nor UO_2218 (O_2218,N_26059,N_29495);
xnor UO_2219 (O_2219,N_26920,N_26466);
xor UO_2220 (O_2220,N_27261,N_25374);
nor UO_2221 (O_2221,N_27551,N_29582);
or UO_2222 (O_2222,N_28348,N_28176);
and UO_2223 (O_2223,N_26479,N_28528);
and UO_2224 (O_2224,N_27306,N_28423);
xor UO_2225 (O_2225,N_26058,N_26994);
nor UO_2226 (O_2226,N_28739,N_25488);
and UO_2227 (O_2227,N_29126,N_29275);
nand UO_2228 (O_2228,N_26488,N_27962);
xnor UO_2229 (O_2229,N_27348,N_26864);
nor UO_2230 (O_2230,N_27632,N_26262);
or UO_2231 (O_2231,N_27913,N_26594);
nand UO_2232 (O_2232,N_29093,N_28301);
nor UO_2233 (O_2233,N_26188,N_25029);
or UO_2234 (O_2234,N_26443,N_26546);
nor UO_2235 (O_2235,N_27852,N_28120);
nand UO_2236 (O_2236,N_28683,N_26225);
and UO_2237 (O_2237,N_29213,N_27935);
or UO_2238 (O_2238,N_27667,N_26790);
xor UO_2239 (O_2239,N_28441,N_25502);
or UO_2240 (O_2240,N_25513,N_27630);
nand UO_2241 (O_2241,N_27124,N_26140);
or UO_2242 (O_2242,N_29696,N_25182);
nand UO_2243 (O_2243,N_26139,N_25492);
nor UO_2244 (O_2244,N_28711,N_26635);
nor UO_2245 (O_2245,N_27157,N_27017);
xor UO_2246 (O_2246,N_27434,N_28772);
nor UO_2247 (O_2247,N_29944,N_27733);
or UO_2248 (O_2248,N_27862,N_27405);
nor UO_2249 (O_2249,N_26423,N_28470);
nor UO_2250 (O_2250,N_26610,N_27044);
or UO_2251 (O_2251,N_25245,N_25535);
or UO_2252 (O_2252,N_25875,N_28105);
nor UO_2253 (O_2253,N_25010,N_28056);
nand UO_2254 (O_2254,N_29231,N_25149);
nor UO_2255 (O_2255,N_25903,N_28532);
and UO_2256 (O_2256,N_26445,N_25446);
or UO_2257 (O_2257,N_29383,N_25017);
nor UO_2258 (O_2258,N_27288,N_27038);
or UO_2259 (O_2259,N_27164,N_27870);
and UO_2260 (O_2260,N_29338,N_27079);
or UO_2261 (O_2261,N_28259,N_25080);
nor UO_2262 (O_2262,N_25802,N_27885);
nand UO_2263 (O_2263,N_27863,N_28337);
and UO_2264 (O_2264,N_29791,N_27571);
xnor UO_2265 (O_2265,N_27063,N_27666);
and UO_2266 (O_2266,N_29268,N_25661);
nor UO_2267 (O_2267,N_25525,N_26033);
nor UO_2268 (O_2268,N_29546,N_26029);
nand UO_2269 (O_2269,N_27948,N_25198);
or UO_2270 (O_2270,N_26227,N_26132);
and UO_2271 (O_2271,N_25716,N_26084);
or UO_2272 (O_2272,N_29551,N_28407);
xor UO_2273 (O_2273,N_26259,N_27829);
and UO_2274 (O_2274,N_26380,N_29237);
and UO_2275 (O_2275,N_29982,N_25595);
and UO_2276 (O_2276,N_25948,N_28229);
or UO_2277 (O_2277,N_25865,N_27596);
nand UO_2278 (O_2278,N_28306,N_25141);
xor UO_2279 (O_2279,N_27498,N_29049);
nand UO_2280 (O_2280,N_26109,N_28185);
or UO_2281 (O_2281,N_29923,N_25343);
or UO_2282 (O_2282,N_27103,N_28604);
or UO_2283 (O_2283,N_26389,N_29387);
and UO_2284 (O_2284,N_26138,N_29086);
and UO_2285 (O_2285,N_28264,N_27556);
nor UO_2286 (O_2286,N_29193,N_25552);
xor UO_2287 (O_2287,N_26539,N_25615);
nor UO_2288 (O_2288,N_29925,N_27194);
xor UO_2289 (O_2289,N_29807,N_28180);
and UO_2290 (O_2290,N_26253,N_27841);
and UO_2291 (O_2291,N_25633,N_28181);
or UO_2292 (O_2292,N_26842,N_26278);
xnor UO_2293 (O_2293,N_27642,N_25803);
or UO_2294 (O_2294,N_26489,N_27190);
nand UO_2295 (O_2295,N_27136,N_26666);
or UO_2296 (O_2296,N_27449,N_26744);
nor UO_2297 (O_2297,N_28862,N_25259);
or UO_2298 (O_2298,N_26962,N_26855);
or UO_2299 (O_2299,N_29110,N_27840);
and UO_2300 (O_2300,N_28150,N_26174);
nor UO_2301 (O_2301,N_28444,N_29658);
nand UO_2302 (O_2302,N_27477,N_26693);
xor UO_2303 (O_2303,N_27442,N_25108);
nand UO_2304 (O_2304,N_25959,N_28840);
and UO_2305 (O_2305,N_26662,N_26890);
nand UO_2306 (O_2306,N_26183,N_26349);
xor UO_2307 (O_2307,N_29855,N_29912);
and UO_2308 (O_2308,N_25131,N_25479);
and UO_2309 (O_2309,N_26289,N_28723);
nand UO_2310 (O_2310,N_27024,N_28942);
nand UO_2311 (O_2311,N_28670,N_25423);
xnor UO_2312 (O_2312,N_29808,N_27665);
nand UO_2313 (O_2313,N_26178,N_26194);
nor UO_2314 (O_2314,N_28686,N_26633);
or UO_2315 (O_2315,N_26946,N_27881);
and UO_2316 (O_2316,N_29749,N_28584);
nor UO_2317 (O_2317,N_28548,N_29904);
and UO_2318 (O_2318,N_25123,N_29068);
nor UO_2319 (O_2319,N_27723,N_25703);
nand UO_2320 (O_2320,N_26707,N_28793);
nand UO_2321 (O_2321,N_28476,N_29692);
and UO_2322 (O_2322,N_25083,N_25196);
and UO_2323 (O_2323,N_27751,N_26300);
nor UO_2324 (O_2324,N_27268,N_26452);
xnor UO_2325 (O_2325,N_26730,N_26382);
or UO_2326 (O_2326,N_25394,N_29245);
nor UO_2327 (O_2327,N_28502,N_26026);
xnor UO_2328 (O_2328,N_29457,N_28625);
nand UO_2329 (O_2329,N_27558,N_28874);
and UO_2330 (O_2330,N_27215,N_27000);
or UO_2331 (O_2331,N_25477,N_27754);
nor UO_2332 (O_2332,N_28541,N_27335);
nand UO_2333 (O_2333,N_28309,N_26797);
or UO_2334 (O_2334,N_29565,N_25515);
or UO_2335 (O_2335,N_28427,N_28052);
and UO_2336 (O_2336,N_27869,N_27152);
nand UO_2337 (O_2337,N_28211,N_29121);
xor UO_2338 (O_2338,N_28903,N_25202);
or UO_2339 (O_2339,N_25431,N_25414);
xnor UO_2340 (O_2340,N_27740,N_28642);
and UO_2341 (O_2341,N_28484,N_26426);
xor UO_2342 (O_2342,N_26216,N_29640);
nor UO_2343 (O_2343,N_27085,N_29682);
nand UO_2344 (O_2344,N_25718,N_29839);
or UO_2345 (O_2345,N_28428,N_29374);
or UO_2346 (O_2346,N_25292,N_29567);
or UO_2347 (O_2347,N_25904,N_27347);
and UO_2348 (O_2348,N_26849,N_25385);
and UO_2349 (O_2349,N_26679,N_29419);
nand UO_2350 (O_2350,N_27212,N_26283);
nand UO_2351 (O_2351,N_25689,N_29620);
nor UO_2352 (O_2352,N_28782,N_29803);
and UO_2353 (O_2353,N_25592,N_28184);
or UO_2354 (O_2354,N_25695,N_28075);
xor UO_2355 (O_2355,N_28561,N_28177);
nor UO_2356 (O_2356,N_29527,N_28183);
or UO_2357 (O_2357,N_28748,N_28243);
and UO_2358 (O_2358,N_29730,N_29602);
and UO_2359 (O_2359,N_27457,N_29224);
xor UO_2360 (O_2360,N_29984,N_29331);
nand UO_2361 (O_2361,N_26691,N_27226);
and UO_2362 (O_2362,N_29278,N_28503);
and UO_2363 (O_2363,N_25870,N_26203);
and UO_2364 (O_2364,N_29795,N_26453);
and UO_2365 (O_2365,N_25792,N_28156);
nor UO_2366 (O_2366,N_28970,N_26724);
nor UO_2367 (O_2367,N_27900,N_29476);
or UO_2368 (O_2368,N_26722,N_28016);
nand UO_2369 (O_2369,N_27009,N_25511);
or UO_2370 (O_2370,N_26374,N_28230);
xnor UO_2371 (O_2371,N_29778,N_27793);
xor UO_2372 (O_2372,N_28039,N_25660);
nand UO_2373 (O_2373,N_27930,N_26511);
or UO_2374 (O_2374,N_29123,N_29058);
nand UO_2375 (O_2375,N_25546,N_25368);
and UO_2376 (O_2376,N_26348,N_28960);
nand UO_2377 (O_2377,N_25677,N_29971);
nand UO_2378 (O_2378,N_28721,N_29896);
and UO_2379 (O_2379,N_28501,N_27497);
xnor UO_2380 (O_2380,N_27683,N_27231);
nor UO_2381 (O_2381,N_27650,N_27270);
and UO_2382 (O_2382,N_25006,N_29402);
nor UO_2383 (O_2383,N_25635,N_29298);
nor UO_2384 (O_2384,N_29013,N_26118);
or UO_2385 (O_2385,N_25471,N_27904);
or UO_2386 (O_2386,N_29111,N_26557);
nor UO_2387 (O_2387,N_29252,N_25857);
or UO_2388 (O_2388,N_29106,N_28742);
or UO_2389 (O_2389,N_25473,N_25662);
and UO_2390 (O_2390,N_27781,N_28320);
nand UO_2391 (O_2391,N_28220,N_29375);
nand UO_2392 (O_2392,N_25140,N_28558);
or UO_2393 (O_2393,N_27681,N_28396);
and UO_2394 (O_2394,N_25229,N_27925);
xor UO_2395 (O_2395,N_26980,N_29092);
nor UO_2396 (O_2396,N_27813,N_25526);
or UO_2397 (O_2397,N_27474,N_28000);
nand UO_2398 (O_2398,N_26368,N_28073);
or UO_2399 (O_2399,N_25000,N_28268);
nand UO_2400 (O_2400,N_26911,N_28205);
nand UO_2401 (O_2401,N_25732,N_25165);
or UO_2402 (O_2402,N_29580,N_25531);
nand UO_2403 (O_2403,N_29366,N_29295);
xor UO_2404 (O_2404,N_27371,N_26145);
nand UO_2405 (O_2405,N_28715,N_29420);
or UO_2406 (O_2406,N_25463,N_26888);
and UO_2407 (O_2407,N_29886,N_25943);
nor UO_2408 (O_2408,N_27465,N_28678);
xnor UO_2409 (O_2409,N_26853,N_27570);
and UO_2410 (O_2410,N_25057,N_25935);
or UO_2411 (O_2411,N_27096,N_29403);
nor UO_2412 (O_2412,N_28631,N_27423);
nand UO_2413 (O_2413,N_29502,N_26840);
nor UO_2414 (O_2414,N_27548,N_27221);
nand UO_2415 (O_2415,N_28925,N_27213);
xor UO_2416 (O_2416,N_26504,N_29080);
and UO_2417 (O_2417,N_26045,N_27742);
nor UO_2418 (O_2418,N_28384,N_25066);
xnor UO_2419 (O_2419,N_25569,N_27612);
nand UO_2420 (O_2420,N_27188,N_28651);
nor UO_2421 (O_2421,N_25234,N_25176);
and UO_2422 (O_2422,N_29862,N_25702);
and UO_2423 (O_2423,N_29474,N_28466);
and UO_2424 (O_2424,N_27614,N_25449);
nand UO_2425 (O_2425,N_27752,N_29956);
or UO_2426 (O_2426,N_29003,N_29561);
or UO_2427 (O_2427,N_28729,N_26429);
or UO_2428 (O_2428,N_28128,N_27903);
or UO_2429 (O_2429,N_27058,N_29458);
xnor UO_2430 (O_2430,N_25599,N_25909);
nor UO_2431 (O_2431,N_25356,N_28082);
xor UO_2432 (O_2432,N_25809,N_27992);
or UO_2433 (O_2433,N_25393,N_25481);
xor UO_2434 (O_2434,N_27453,N_29427);
nor UO_2435 (O_2435,N_28810,N_28783);
and UO_2436 (O_2436,N_29466,N_25496);
nor UO_2437 (O_2437,N_27452,N_29128);
xnor UO_2438 (O_2438,N_25804,N_29771);
xor UO_2439 (O_2439,N_28887,N_27133);
and UO_2440 (O_2440,N_26064,N_25093);
nand UO_2441 (O_2441,N_25297,N_28953);
or UO_2442 (O_2442,N_28761,N_27499);
nand UO_2443 (O_2443,N_28709,N_27237);
xor UO_2444 (O_2444,N_26127,N_26979);
nand UO_2445 (O_2445,N_25411,N_27954);
nand UO_2446 (O_2446,N_29884,N_27071);
nor UO_2447 (O_2447,N_28560,N_29217);
or UO_2448 (O_2448,N_27214,N_26951);
or UO_2449 (O_2449,N_28198,N_28372);
nor UO_2450 (O_2450,N_25016,N_25285);
and UO_2451 (O_2451,N_28510,N_29250);
nand UO_2452 (O_2452,N_25366,N_25777);
nand UO_2453 (O_2453,N_25113,N_25107);
or UO_2454 (O_2454,N_27827,N_27198);
xor UO_2455 (O_2455,N_28224,N_27586);
nand UO_2456 (O_2456,N_26459,N_26400);
or UO_2457 (O_2457,N_26254,N_25593);
and UO_2458 (O_2458,N_25966,N_25840);
nor UO_2459 (O_2459,N_25372,N_25863);
nand UO_2460 (O_2460,N_26711,N_27524);
and UO_2461 (O_2461,N_25780,N_26141);
xor UO_2462 (O_2462,N_29800,N_29901);
nand UO_2463 (O_2463,N_27154,N_26598);
and UO_2464 (O_2464,N_27859,N_26161);
nor UO_2465 (O_2465,N_27046,N_26037);
nand UO_2466 (O_2466,N_26435,N_27659);
or UO_2467 (O_2467,N_28037,N_28125);
nor UO_2468 (O_2468,N_26014,N_26093);
xnor UO_2469 (O_2469,N_25867,N_27758);
or UO_2470 (O_2470,N_25772,N_28544);
nand UO_2471 (O_2471,N_25657,N_26777);
or UO_2472 (O_2472,N_28987,N_28045);
nand UO_2473 (O_2473,N_26403,N_28246);
and UO_2474 (O_2474,N_28720,N_25311);
nor UO_2475 (O_2475,N_26943,N_26606);
nand UO_2476 (O_2476,N_29297,N_29554);
nor UO_2477 (O_2477,N_26552,N_28195);
xnor UO_2478 (O_2478,N_28884,N_25336);
nand UO_2479 (O_2479,N_25023,N_28675);
and UO_2480 (O_2480,N_29718,N_26098);
nor UO_2481 (O_2481,N_29538,N_28933);
nand UO_2482 (O_2482,N_27271,N_28192);
or UO_2483 (O_2483,N_25538,N_28922);
xor UO_2484 (O_2484,N_28980,N_26336);
nor UO_2485 (O_2485,N_28273,N_25914);
or UO_2486 (O_2486,N_26233,N_28081);
xor UO_2487 (O_2487,N_28196,N_28895);
nor UO_2488 (O_2488,N_26495,N_25877);
nor UO_2489 (O_2489,N_26915,N_28498);
nor UO_2490 (O_2490,N_28621,N_28029);
and UO_2491 (O_2491,N_29694,N_25068);
or UO_2492 (O_2492,N_25579,N_29724);
and UO_2493 (O_2493,N_25180,N_27523);
nand UO_2494 (O_2494,N_29103,N_27845);
or UO_2495 (O_2495,N_25591,N_28472);
and UO_2496 (O_2496,N_29996,N_26043);
and UO_2497 (O_2497,N_29738,N_25653);
or UO_2498 (O_2498,N_28737,N_28716);
and UO_2499 (O_2499,N_26584,N_28409);
and UO_2500 (O_2500,N_25654,N_27894);
nor UO_2501 (O_2501,N_25337,N_27407);
or UO_2502 (O_2502,N_25561,N_27486);
xnor UO_2503 (O_2503,N_28734,N_27440);
xnor UO_2504 (O_2504,N_25719,N_25846);
xor UO_2505 (O_2505,N_29601,N_27892);
nand UO_2506 (O_2506,N_27497,N_26566);
nand UO_2507 (O_2507,N_27868,N_28830);
xnor UO_2508 (O_2508,N_28757,N_27357);
nand UO_2509 (O_2509,N_28994,N_28923);
and UO_2510 (O_2510,N_29321,N_26485);
or UO_2511 (O_2511,N_26697,N_27177);
and UO_2512 (O_2512,N_28159,N_28848);
and UO_2513 (O_2513,N_29609,N_25351);
nor UO_2514 (O_2514,N_27025,N_27853);
nor UO_2515 (O_2515,N_28316,N_26526);
or UO_2516 (O_2516,N_25418,N_29256);
and UO_2517 (O_2517,N_29092,N_29543);
or UO_2518 (O_2518,N_25245,N_28512);
or UO_2519 (O_2519,N_28299,N_28269);
nor UO_2520 (O_2520,N_28628,N_29299);
xnor UO_2521 (O_2521,N_29679,N_25327);
nor UO_2522 (O_2522,N_26577,N_28843);
or UO_2523 (O_2523,N_29471,N_26671);
xor UO_2524 (O_2524,N_25026,N_27202);
or UO_2525 (O_2525,N_26938,N_27800);
or UO_2526 (O_2526,N_25706,N_28333);
xor UO_2527 (O_2527,N_27758,N_25143);
nand UO_2528 (O_2528,N_29577,N_25740);
xor UO_2529 (O_2529,N_26971,N_26288);
nand UO_2530 (O_2530,N_26750,N_28945);
xnor UO_2531 (O_2531,N_27526,N_27969);
nand UO_2532 (O_2532,N_25336,N_26322);
or UO_2533 (O_2533,N_28429,N_28190);
or UO_2534 (O_2534,N_26320,N_28900);
nand UO_2535 (O_2535,N_29173,N_28290);
nand UO_2536 (O_2536,N_26048,N_28805);
and UO_2537 (O_2537,N_29104,N_27295);
nand UO_2538 (O_2538,N_26811,N_27735);
nand UO_2539 (O_2539,N_25016,N_27929);
and UO_2540 (O_2540,N_25242,N_26934);
or UO_2541 (O_2541,N_27058,N_25254);
xor UO_2542 (O_2542,N_29978,N_28107);
or UO_2543 (O_2543,N_26803,N_25672);
and UO_2544 (O_2544,N_27178,N_27753);
and UO_2545 (O_2545,N_25938,N_27538);
or UO_2546 (O_2546,N_27473,N_25027);
xnor UO_2547 (O_2547,N_28224,N_29163);
nand UO_2548 (O_2548,N_29836,N_25348);
nor UO_2549 (O_2549,N_26781,N_26355);
and UO_2550 (O_2550,N_29770,N_28232);
or UO_2551 (O_2551,N_28117,N_25013);
and UO_2552 (O_2552,N_28914,N_25690);
nor UO_2553 (O_2553,N_28743,N_26975);
and UO_2554 (O_2554,N_26021,N_26856);
xnor UO_2555 (O_2555,N_27431,N_26390);
nand UO_2556 (O_2556,N_26461,N_27834);
xnor UO_2557 (O_2557,N_27940,N_26423);
nor UO_2558 (O_2558,N_26585,N_26299);
or UO_2559 (O_2559,N_27156,N_28697);
nand UO_2560 (O_2560,N_29435,N_25921);
xnor UO_2561 (O_2561,N_26628,N_25515);
nand UO_2562 (O_2562,N_28112,N_29267);
or UO_2563 (O_2563,N_27849,N_29224);
nor UO_2564 (O_2564,N_26397,N_29394);
nor UO_2565 (O_2565,N_28485,N_29544);
or UO_2566 (O_2566,N_29762,N_25383);
nand UO_2567 (O_2567,N_27657,N_25545);
nor UO_2568 (O_2568,N_25307,N_25723);
xor UO_2569 (O_2569,N_29063,N_25487);
and UO_2570 (O_2570,N_26039,N_26124);
and UO_2571 (O_2571,N_26021,N_25105);
xor UO_2572 (O_2572,N_26044,N_29543);
and UO_2573 (O_2573,N_28247,N_29927);
and UO_2574 (O_2574,N_26272,N_27077);
and UO_2575 (O_2575,N_29991,N_27216);
nand UO_2576 (O_2576,N_27510,N_25854);
or UO_2577 (O_2577,N_28632,N_27094);
nor UO_2578 (O_2578,N_25797,N_25812);
and UO_2579 (O_2579,N_27933,N_27856);
nand UO_2580 (O_2580,N_27985,N_25962);
or UO_2581 (O_2581,N_29267,N_26790);
or UO_2582 (O_2582,N_27043,N_25313);
and UO_2583 (O_2583,N_29345,N_25478);
nand UO_2584 (O_2584,N_27015,N_27965);
or UO_2585 (O_2585,N_25536,N_28638);
and UO_2586 (O_2586,N_26242,N_25409);
and UO_2587 (O_2587,N_28410,N_26979);
nand UO_2588 (O_2588,N_29612,N_25568);
nor UO_2589 (O_2589,N_26230,N_27750);
xnor UO_2590 (O_2590,N_26844,N_27666);
xor UO_2591 (O_2591,N_27311,N_25409);
and UO_2592 (O_2592,N_29738,N_26583);
nor UO_2593 (O_2593,N_29062,N_25249);
xor UO_2594 (O_2594,N_29887,N_25978);
nor UO_2595 (O_2595,N_25291,N_26512);
xnor UO_2596 (O_2596,N_29716,N_29208);
and UO_2597 (O_2597,N_25275,N_26453);
nor UO_2598 (O_2598,N_29302,N_28968);
or UO_2599 (O_2599,N_27215,N_25207);
nor UO_2600 (O_2600,N_28948,N_26434);
xnor UO_2601 (O_2601,N_25301,N_28011);
and UO_2602 (O_2602,N_28914,N_25166);
or UO_2603 (O_2603,N_27969,N_29974);
nand UO_2604 (O_2604,N_26038,N_28781);
or UO_2605 (O_2605,N_29397,N_28948);
xnor UO_2606 (O_2606,N_26477,N_29451);
or UO_2607 (O_2607,N_28131,N_27478);
or UO_2608 (O_2608,N_25556,N_29067);
and UO_2609 (O_2609,N_26101,N_25159);
and UO_2610 (O_2610,N_25365,N_26038);
or UO_2611 (O_2611,N_26431,N_27170);
xor UO_2612 (O_2612,N_26967,N_26574);
xnor UO_2613 (O_2613,N_26630,N_28344);
or UO_2614 (O_2614,N_25172,N_27708);
or UO_2615 (O_2615,N_25331,N_28701);
nor UO_2616 (O_2616,N_25108,N_26304);
or UO_2617 (O_2617,N_25110,N_29842);
or UO_2618 (O_2618,N_25764,N_28069);
or UO_2619 (O_2619,N_26479,N_28939);
nor UO_2620 (O_2620,N_25880,N_25225);
and UO_2621 (O_2621,N_26567,N_27373);
nor UO_2622 (O_2622,N_29208,N_25698);
or UO_2623 (O_2623,N_27876,N_25388);
xor UO_2624 (O_2624,N_29355,N_29501);
nand UO_2625 (O_2625,N_27483,N_27728);
nand UO_2626 (O_2626,N_28317,N_29796);
xor UO_2627 (O_2627,N_25669,N_27394);
xor UO_2628 (O_2628,N_29125,N_28642);
xnor UO_2629 (O_2629,N_28852,N_27691);
nor UO_2630 (O_2630,N_28378,N_29071);
nand UO_2631 (O_2631,N_26028,N_27003);
or UO_2632 (O_2632,N_25906,N_27324);
and UO_2633 (O_2633,N_27804,N_29703);
nand UO_2634 (O_2634,N_25371,N_25463);
xnor UO_2635 (O_2635,N_25769,N_29280);
xor UO_2636 (O_2636,N_25888,N_25793);
nand UO_2637 (O_2637,N_27047,N_27381);
nand UO_2638 (O_2638,N_25007,N_27021);
or UO_2639 (O_2639,N_26419,N_25196);
nand UO_2640 (O_2640,N_27940,N_27878);
xnor UO_2641 (O_2641,N_27969,N_25106);
and UO_2642 (O_2642,N_28340,N_27220);
xnor UO_2643 (O_2643,N_25097,N_29722);
nand UO_2644 (O_2644,N_25069,N_29541);
xor UO_2645 (O_2645,N_26398,N_25162);
nor UO_2646 (O_2646,N_26225,N_28655);
or UO_2647 (O_2647,N_29576,N_26184);
and UO_2648 (O_2648,N_27393,N_28177);
xnor UO_2649 (O_2649,N_27317,N_28246);
xnor UO_2650 (O_2650,N_27499,N_25679);
nand UO_2651 (O_2651,N_27516,N_28090);
nand UO_2652 (O_2652,N_29594,N_29509);
nand UO_2653 (O_2653,N_28749,N_26896);
xor UO_2654 (O_2654,N_25227,N_29763);
nand UO_2655 (O_2655,N_25975,N_26708);
and UO_2656 (O_2656,N_26182,N_25108);
and UO_2657 (O_2657,N_27075,N_29156);
nand UO_2658 (O_2658,N_28746,N_29788);
and UO_2659 (O_2659,N_25914,N_26040);
xnor UO_2660 (O_2660,N_27321,N_29958);
xnor UO_2661 (O_2661,N_27573,N_27332);
nand UO_2662 (O_2662,N_26978,N_25040);
and UO_2663 (O_2663,N_27006,N_27306);
and UO_2664 (O_2664,N_28685,N_29146);
xor UO_2665 (O_2665,N_28593,N_28268);
nor UO_2666 (O_2666,N_28535,N_27779);
xnor UO_2667 (O_2667,N_28569,N_29106);
xnor UO_2668 (O_2668,N_25814,N_27922);
nor UO_2669 (O_2669,N_27231,N_26429);
nor UO_2670 (O_2670,N_25243,N_25641);
xor UO_2671 (O_2671,N_29320,N_28748);
nand UO_2672 (O_2672,N_25236,N_26910);
and UO_2673 (O_2673,N_25939,N_27561);
or UO_2674 (O_2674,N_25462,N_28052);
xor UO_2675 (O_2675,N_28970,N_27240);
and UO_2676 (O_2676,N_29964,N_29639);
nand UO_2677 (O_2677,N_29420,N_29943);
nand UO_2678 (O_2678,N_25260,N_27128);
or UO_2679 (O_2679,N_27090,N_26407);
nor UO_2680 (O_2680,N_26006,N_25877);
nor UO_2681 (O_2681,N_26206,N_25621);
nand UO_2682 (O_2682,N_26216,N_25531);
and UO_2683 (O_2683,N_27607,N_25075);
nor UO_2684 (O_2684,N_29671,N_28862);
or UO_2685 (O_2685,N_27004,N_26514);
and UO_2686 (O_2686,N_26699,N_25454);
xor UO_2687 (O_2687,N_28047,N_29988);
and UO_2688 (O_2688,N_26780,N_25878);
or UO_2689 (O_2689,N_27864,N_26768);
and UO_2690 (O_2690,N_27350,N_28903);
or UO_2691 (O_2691,N_29384,N_27716);
and UO_2692 (O_2692,N_25128,N_28073);
and UO_2693 (O_2693,N_28336,N_28268);
nand UO_2694 (O_2694,N_25111,N_29606);
or UO_2695 (O_2695,N_25183,N_25214);
xnor UO_2696 (O_2696,N_25178,N_28356);
and UO_2697 (O_2697,N_25163,N_28958);
nand UO_2698 (O_2698,N_29631,N_29532);
nor UO_2699 (O_2699,N_25961,N_29749);
nor UO_2700 (O_2700,N_26338,N_29198);
and UO_2701 (O_2701,N_25000,N_29381);
or UO_2702 (O_2702,N_25553,N_27771);
or UO_2703 (O_2703,N_27343,N_28595);
xor UO_2704 (O_2704,N_27181,N_29422);
nand UO_2705 (O_2705,N_26046,N_25526);
and UO_2706 (O_2706,N_27654,N_28013);
or UO_2707 (O_2707,N_25642,N_27140);
or UO_2708 (O_2708,N_27688,N_29222);
nand UO_2709 (O_2709,N_28490,N_26470);
nand UO_2710 (O_2710,N_25929,N_25142);
nand UO_2711 (O_2711,N_28720,N_27038);
nor UO_2712 (O_2712,N_26994,N_29057);
or UO_2713 (O_2713,N_25954,N_27233);
nand UO_2714 (O_2714,N_27573,N_29957);
nor UO_2715 (O_2715,N_26042,N_25535);
nand UO_2716 (O_2716,N_25863,N_27607);
nand UO_2717 (O_2717,N_29425,N_27266);
nand UO_2718 (O_2718,N_27747,N_25645);
and UO_2719 (O_2719,N_27724,N_25015);
or UO_2720 (O_2720,N_29213,N_28692);
xor UO_2721 (O_2721,N_28812,N_28958);
nor UO_2722 (O_2722,N_27490,N_28980);
xnor UO_2723 (O_2723,N_26016,N_27009);
or UO_2724 (O_2724,N_26253,N_28577);
nand UO_2725 (O_2725,N_29531,N_27260);
and UO_2726 (O_2726,N_25919,N_29676);
and UO_2727 (O_2727,N_29575,N_25283);
nand UO_2728 (O_2728,N_27473,N_28532);
and UO_2729 (O_2729,N_25701,N_27234);
or UO_2730 (O_2730,N_26663,N_27347);
and UO_2731 (O_2731,N_28303,N_25727);
or UO_2732 (O_2732,N_28168,N_29246);
and UO_2733 (O_2733,N_29117,N_26083);
nand UO_2734 (O_2734,N_25148,N_28825);
nor UO_2735 (O_2735,N_29615,N_25459);
nor UO_2736 (O_2736,N_26889,N_27529);
xor UO_2737 (O_2737,N_29667,N_26111);
and UO_2738 (O_2738,N_28539,N_29217);
or UO_2739 (O_2739,N_29115,N_29539);
xnor UO_2740 (O_2740,N_29118,N_28436);
or UO_2741 (O_2741,N_29579,N_28009);
or UO_2742 (O_2742,N_27745,N_28873);
nand UO_2743 (O_2743,N_27780,N_26582);
xnor UO_2744 (O_2744,N_27975,N_28760);
nand UO_2745 (O_2745,N_28165,N_27517);
and UO_2746 (O_2746,N_27097,N_25599);
or UO_2747 (O_2747,N_27057,N_26026);
xor UO_2748 (O_2748,N_29142,N_27208);
xnor UO_2749 (O_2749,N_25429,N_25827);
xnor UO_2750 (O_2750,N_29283,N_28333);
and UO_2751 (O_2751,N_26259,N_27808);
xor UO_2752 (O_2752,N_28069,N_26595);
nor UO_2753 (O_2753,N_26363,N_26204);
or UO_2754 (O_2754,N_28286,N_27300);
xnor UO_2755 (O_2755,N_27722,N_28365);
nand UO_2756 (O_2756,N_27964,N_27075);
xor UO_2757 (O_2757,N_25873,N_27352);
and UO_2758 (O_2758,N_28107,N_29463);
nor UO_2759 (O_2759,N_29683,N_27058);
or UO_2760 (O_2760,N_26423,N_27832);
or UO_2761 (O_2761,N_29457,N_25788);
and UO_2762 (O_2762,N_29470,N_27057);
and UO_2763 (O_2763,N_29137,N_25253);
nand UO_2764 (O_2764,N_28460,N_26484);
or UO_2765 (O_2765,N_27232,N_26328);
nand UO_2766 (O_2766,N_25560,N_29571);
xnor UO_2767 (O_2767,N_29022,N_25522);
nor UO_2768 (O_2768,N_28959,N_28824);
nor UO_2769 (O_2769,N_27955,N_28996);
xnor UO_2770 (O_2770,N_25303,N_27593);
or UO_2771 (O_2771,N_25805,N_28265);
and UO_2772 (O_2772,N_26171,N_29296);
nor UO_2773 (O_2773,N_28665,N_29732);
or UO_2774 (O_2774,N_29502,N_29916);
nor UO_2775 (O_2775,N_27754,N_27352);
nand UO_2776 (O_2776,N_25278,N_27917);
or UO_2777 (O_2777,N_25218,N_29794);
or UO_2778 (O_2778,N_29784,N_25819);
or UO_2779 (O_2779,N_28699,N_26394);
nand UO_2780 (O_2780,N_25572,N_25937);
xnor UO_2781 (O_2781,N_29448,N_29572);
xnor UO_2782 (O_2782,N_26507,N_28541);
and UO_2783 (O_2783,N_26655,N_29405);
and UO_2784 (O_2784,N_29347,N_26275);
nand UO_2785 (O_2785,N_28318,N_29350);
nor UO_2786 (O_2786,N_27987,N_28248);
or UO_2787 (O_2787,N_26749,N_27566);
or UO_2788 (O_2788,N_27520,N_26537);
or UO_2789 (O_2789,N_29140,N_26381);
nor UO_2790 (O_2790,N_25878,N_27758);
and UO_2791 (O_2791,N_28837,N_29754);
nand UO_2792 (O_2792,N_27199,N_25329);
xor UO_2793 (O_2793,N_26437,N_29438);
nor UO_2794 (O_2794,N_25906,N_29044);
nor UO_2795 (O_2795,N_26904,N_26188);
or UO_2796 (O_2796,N_27585,N_25725);
or UO_2797 (O_2797,N_25770,N_27705);
xor UO_2798 (O_2798,N_29448,N_26943);
or UO_2799 (O_2799,N_28519,N_27426);
nor UO_2800 (O_2800,N_26747,N_26273);
xnor UO_2801 (O_2801,N_28397,N_26731);
nand UO_2802 (O_2802,N_28925,N_26906);
or UO_2803 (O_2803,N_26758,N_25031);
nand UO_2804 (O_2804,N_29810,N_26700);
and UO_2805 (O_2805,N_25525,N_26092);
and UO_2806 (O_2806,N_26506,N_28319);
and UO_2807 (O_2807,N_25056,N_26227);
nand UO_2808 (O_2808,N_25622,N_26108);
and UO_2809 (O_2809,N_29965,N_29348);
nand UO_2810 (O_2810,N_28168,N_26740);
xnor UO_2811 (O_2811,N_26440,N_28196);
nor UO_2812 (O_2812,N_29144,N_26644);
nand UO_2813 (O_2813,N_27715,N_25904);
xor UO_2814 (O_2814,N_28845,N_25959);
or UO_2815 (O_2815,N_25504,N_25948);
xor UO_2816 (O_2816,N_28455,N_25776);
xor UO_2817 (O_2817,N_29581,N_27343);
xnor UO_2818 (O_2818,N_27571,N_25416);
xor UO_2819 (O_2819,N_27871,N_25390);
nor UO_2820 (O_2820,N_27933,N_27307);
or UO_2821 (O_2821,N_25858,N_27328);
and UO_2822 (O_2822,N_28068,N_27464);
or UO_2823 (O_2823,N_28314,N_27555);
and UO_2824 (O_2824,N_26936,N_29691);
and UO_2825 (O_2825,N_25643,N_28363);
xnor UO_2826 (O_2826,N_29296,N_25532);
nand UO_2827 (O_2827,N_28519,N_29106);
xnor UO_2828 (O_2828,N_26001,N_27779);
xor UO_2829 (O_2829,N_26493,N_27077);
nand UO_2830 (O_2830,N_27685,N_27864);
and UO_2831 (O_2831,N_27003,N_28145);
or UO_2832 (O_2832,N_27148,N_29087);
or UO_2833 (O_2833,N_25317,N_25269);
or UO_2834 (O_2834,N_28922,N_28572);
nor UO_2835 (O_2835,N_28461,N_29612);
xor UO_2836 (O_2836,N_27840,N_27192);
nor UO_2837 (O_2837,N_26392,N_25722);
or UO_2838 (O_2838,N_26418,N_27083);
or UO_2839 (O_2839,N_25623,N_26960);
and UO_2840 (O_2840,N_27056,N_26097);
nor UO_2841 (O_2841,N_27154,N_28614);
nand UO_2842 (O_2842,N_26286,N_29061);
nor UO_2843 (O_2843,N_27277,N_25679);
or UO_2844 (O_2844,N_27962,N_27191);
xor UO_2845 (O_2845,N_26455,N_26160);
or UO_2846 (O_2846,N_28655,N_27531);
nor UO_2847 (O_2847,N_25146,N_27598);
xnor UO_2848 (O_2848,N_28013,N_27321);
nand UO_2849 (O_2849,N_27030,N_26012);
xor UO_2850 (O_2850,N_27127,N_25180);
nor UO_2851 (O_2851,N_25040,N_25028);
and UO_2852 (O_2852,N_26436,N_28947);
or UO_2853 (O_2853,N_26213,N_29492);
nor UO_2854 (O_2854,N_28819,N_28797);
nand UO_2855 (O_2855,N_29144,N_25818);
xor UO_2856 (O_2856,N_28502,N_27168);
and UO_2857 (O_2857,N_25350,N_26664);
nor UO_2858 (O_2858,N_28292,N_25497);
xnor UO_2859 (O_2859,N_27879,N_28071);
nand UO_2860 (O_2860,N_25802,N_27729);
and UO_2861 (O_2861,N_29771,N_26950);
or UO_2862 (O_2862,N_27360,N_25072);
nand UO_2863 (O_2863,N_26196,N_26074);
and UO_2864 (O_2864,N_28725,N_26800);
and UO_2865 (O_2865,N_25504,N_27954);
nor UO_2866 (O_2866,N_28050,N_26340);
xor UO_2867 (O_2867,N_26723,N_27599);
xor UO_2868 (O_2868,N_25540,N_27218);
nor UO_2869 (O_2869,N_25801,N_28986);
or UO_2870 (O_2870,N_26595,N_26456);
nand UO_2871 (O_2871,N_28510,N_27764);
nor UO_2872 (O_2872,N_27407,N_26431);
xor UO_2873 (O_2873,N_25658,N_29382);
or UO_2874 (O_2874,N_25435,N_26509);
xor UO_2875 (O_2875,N_27964,N_26732);
xor UO_2876 (O_2876,N_27867,N_27232);
xnor UO_2877 (O_2877,N_25277,N_29009);
xor UO_2878 (O_2878,N_29888,N_28708);
nand UO_2879 (O_2879,N_25230,N_28814);
nor UO_2880 (O_2880,N_28433,N_27686);
and UO_2881 (O_2881,N_25163,N_29976);
nor UO_2882 (O_2882,N_28351,N_26087);
nand UO_2883 (O_2883,N_25541,N_27140);
nand UO_2884 (O_2884,N_25131,N_29201);
or UO_2885 (O_2885,N_29081,N_29336);
or UO_2886 (O_2886,N_27938,N_29707);
nand UO_2887 (O_2887,N_27594,N_27520);
and UO_2888 (O_2888,N_27582,N_28282);
nor UO_2889 (O_2889,N_29198,N_28147);
nor UO_2890 (O_2890,N_27642,N_26035);
or UO_2891 (O_2891,N_27245,N_26445);
xor UO_2892 (O_2892,N_26450,N_27226);
and UO_2893 (O_2893,N_29621,N_28083);
xnor UO_2894 (O_2894,N_27863,N_25149);
and UO_2895 (O_2895,N_25327,N_25407);
xnor UO_2896 (O_2896,N_28548,N_25762);
and UO_2897 (O_2897,N_27224,N_25274);
and UO_2898 (O_2898,N_26824,N_27017);
and UO_2899 (O_2899,N_27621,N_26478);
and UO_2900 (O_2900,N_25485,N_28222);
and UO_2901 (O_2901,N_27365,N_25912);
xnor UO_2902 (O_2902,N_26234,N_29841);
and UO_2903 (O_2903,N_28464,N_29890);
and UO_2904 (O_2904,N_27834,N_25213);
or UO_2905 (O_2905,N_29862,N_29323);
nor UO_2906 (O_2906,N_28242,N_29535);
and UO_2907 (O_2907,N_26321,N_29404);
nand UO_2908 (O_2908,N_29204,N_25338);
xnor UO_2909 (O_2909,N_26813,N_29936);
or UO_2910 (O_2910,N_25602,N_27099);
and UO_2911 (O_2911,N_27574,N_25393);
or UO_2912 (O_2912,N_25354,N_26643);
and UO_2913 (O_2913,N_29602,N_28552);
nand UO_2914 (O_2914,N_28349,N_28948);
or UO_2915 (O_2915,N_29647,N_27123);
nor UO_2916 (O_2916,N_28401,N_26127);
nand UO_2917 (O_2917,N_29356,N_25895);
nor UO_2918 (O_2918,N_25199,N_29765);
or UO_2919 (O_2919,N_28252,N_27034);
xor UO_2920 (O_2920,N_25681,N_28350);
and UO_2921 (O_2921,N_29349,N_29458);
or UO_2922 (O_2922,N_25737,N_25381);
nand UO_2923 (O_2923,N_25516,N_29962);
nand UO_2924 (O_2924,N_26519,N_27485);
xor UO_2925 (O_2925,N_26854,N_26998);
and UO_2926 (O_2926,N_29453,N_27848);
nor UO_2927 (O_2927,N_29354,N_25396);
nor UO_2928 (O_2928,N_29659,N_26723);
or UO_2929 (O_2929,N_29175,N_26407);
and UO_2930 (O_2930,N_25371,N_25158);
and UO_2931 (O_2931,N_25269,N_26856);
nor UO_2932 (O_2932,N_28605,N_28730);
nor UO_2933 (O_2933,N_29302,N_29669);
nor UO_2934 (O_2934,N_29875,N_26453);
xor UO_2935 (O_2935,N_29355,N_27861);
xnor UO_2936 (O_2936,N_26279,N_26802);
nor UO_2937 (O_2937,N_28783,N_28652);
or UO_2938 (O_2938,N_28622,N_27442);
nor UO_2939 (O_2939,N_25888,N_29216);
xor UO_2940 (O_2940,N_29693,N_27390);
nor UO_2941 (O_2941,N_25626,N_28365);
and UO_2942 (O_2942,N_29369,N_26588);
xnor UO_2943 (O_2943,N_28442,N_29736);
and UO_2944 (O_2944,N_25899,N_26027);
xnor UO_2945 (O_2945,N_26288,N_27650);
and UO_2946 (O_2946,N_25024,N_28359);
xnor UO_2947 (O_2947,N_27051,N_29576);
nand UO_2948 (O_2948,N_27673,N_28896);
and UO_2949 (O_2949,N_29538,N_26423);
xnor UO_2950 (O_2950,N_29473,N_28627);
xor UO_2951 (O_2951,N_28742,N_27923);
or UO_2952 (O_2952,N_26315,N_28829);
xor UO_2953 (O_2953,N_28859,N_29204);
or UO_2954 (O_2954,N_26667,N_27189);
or UO_2955 (O_2955,N_29904,N_29713);
xnor UO_2956 (O_2956,N_27769,N_28299);
nand UO_2957 (O_2957,N_26386,N_27292);
nor UO_2958 (O_2958,N_29693,N_25367);
nor UO_2959 (O_2959,N_25328,N_28068);
or UO_2960 (O_2960,N_28086,N_29289);
and UO_2961 (O_2961,N_29676,N_27846);
xnor UO_2962 (O_2962,N_25684,N_29533);
or UO_2963 (O_2963,N_25852,N_29753);
or UO_2964 (O_2964,N_28896,N_26838);
and UO_2965 (O_2965,N_25003,N_28910);
xor UO_2966 (O_2966,N_26024,N_28679);
nor UO_2967 (O_2967,N_27513,N_29544);
or UO_2968 (O_2968,N_27034,N_26272);
and UO_2969 (O_2969,N_28524,N_26844);
xor UO_2970 (O_2970,N_25962,N_26630);
nor UO_2971 (O_2971,N_28482,N_28023);
nor UO_2972 (O_2972,N_28328,N_26129);
nor UO_2973 (O_2973,N_25740,N_26196);
nor UO_2974 (O_2974,N_25684,N_27526);
or UO_2975 (O_2975,N_28447,N_27929);
or UO_2976 (O_2976,N_29438,N_26414);
xnor UO_2977 (O_2977,N_27572,N_28271);
or UO_2978 (O_2978,N_29510,N_27926);
or UO_2979 (O_2979,N_27940,N_25913);
or UO_2980 (O_2980,N_27168,N_27330);
xor UO_2981 (O_2981,N_26400,N_25334);
or UO_2982 (O_2982,N_29700,N_28580);
or UO_2983 (O_2983,N_28726,N_29728);
xor UO_2984 (O_2984,N_29122,N_28935);
nor UO_2985 (O_2985,N_28714,N_29609);
nor UO_2986 (O_2986,N_27803,N_26785);
xnor UO_2987 (O_2987,N_27048,N_27226);
or UO_2988 (O_2988,N_26554,N_25748);
or UO_2989 (O_2989,N_26492,N_25629);
xnor UO_2990 (O_2990,N_28143,N_29295);
or UO_2991 (O_2991,N_25023,N_28516);
nand UO_2992 (O_2992,N_28696,N_28488);
nand UO_2993 (O_2993,N_26005,N_26924);
nor UO_2994 (O_2994,N_28374,N_28940);
or UO_2995 (O_2995,N_28384,N_25202);
or UO_2996 (O_2996,N_26488,N_25289);
nor UO_2997 (O_2997,N_27763,N_26056);
or UO_2998 (O_2998,N_29376,N_29130);
or UO_2999 (O_2999,N_26902,N_27373);
and UO_3000 (O_3000,N_28345,N_25971);
nand UO_3001 (O_3001,N_27973,N_25221);
nor UO_3002 (O_3002,N_29959,N_26212);
and UO_3003 (O_3003,N_25863,N_27484);
or UO_3004 (O_3004,N_29095,N_27126);
nand UO_3005 (O_3005,N_27144,N_26076);
xor UO_3006 (O_3006,N_26682,N_26900);
nand UO_3007 (O_3007,N_27490,N_25550);
and UO_3008 (O_3008,N_26118,N_27804);
and UO_3009 (O_3009,N_27710,N_29682);
nand UO_3010 (O_3010,N_25860,N_26922);
and UO_3011 (O_3011,N_28676,N_25598);
xor UO_3012 (O_3012,N_26028,N_26101);
and UO_3013 (O_3013,N_25032,N_25981);
nand UO_3014 (O_3014,N_25363,N_28328);
and UO_3015 (O_3015,N_25500,N_25781);
nor UO_3016 (O_3016,N_27858,N_25804);
xnor UO_3017 (O_3017,N_29948,N_28578);
nor UO_3018 (O_3018,N_29100,N_28544);
nand UO_3019 (O_3019,N_26136,N_26769);
nor UO_3020 (O_3020,N_28290,N_26491);
or UO_3021 (O_3021,N_26303,N_26829);
or UO_3022 (O_3022,N_29023,N_25653);
nor UO_3023 (O_3023,N_29789,N_25278);
and UO_3024 (O_3024,N_27152,N_26089);
or UO_3025 (O_3025,N_28299,N_29987);
or UO_3026 (O_3026,N_29870,N_27187);
nand UO_3027 (O_3027,N_29294,N_28190);
or UO_3028 (O_3028,N_25372,N_27791);
nand UO_3029 (O_3029,N_25341,N_29595);
xnor UO_3030 (O_3030,N_27998,N_25866);
nor UO_3031 (O_3031,N_25474,N_25034);
nand UO_3032 (O_3032,N_26041,N_25423);
xnor UO_3033 (O_3033,N_25225,N_26034);
nand UO_3034 (O_3034,N_25780,N_29622);
nand UO_3035 (O_3035,N_29226,N_26529);
or UO_3036 (O_3036,N_29609,N_25906);
nor UO_3037 (O_3037,N_26465,N_29368);
nand UO_3038 (O_3038,N_29163,N_27074);
xnor UO_3039 (O_3039,N_25385,N_29276);
or UO_3040 (O_3040,N_28417,N_29158);
or UO_3041 (O_3041,N_29000,N_29644);
or UO_3042 (O_3042,N_25658,N_27816);
xnor UO_3043 (O_3043,N_25984,N_27206);
nor UO_3044 (O_3044,N_29262,N_29504);
or UO_3045 (O_3045,N_25147,N_29676);
nor UO_3046 (O_3046,N_25917,N_26650);
and UO_3047 (O_3047,N_26251,N_28324);
xnor UO_3048 (O_3048,N_25955,N_29204);
nor UO_3049 (O_3049,N_27068,N_26959);
xor UO_3050 (O_3050,N_29071,N_28852);
nand UO_3051 (O_3051,N_27605,N_27326);
nand UO_3052 (O_3052,N_26614,N_27195);
xor UO_3053 (O_3053,N_27396,N_29982);
nor UO_3054 (O_3054,N_25958,N_29039);
nor UO_3055 (O_3055,N_28696,N_29247);
or UO_3056 (O_3056,N_29215,N_25347);
xnor UO_3057 (O_3057,N_27116,N_27227);
nor UO_3058 (O_3058,N_28270,N_29999);
or UO_3059 (O_3059,N_29098,N_26430);
nand UO_3060 (O_3060,N_28308,N_26015);
nand UO_3061 (O_3061,N_28407,N_25780);
xnor UO_3062 (O_3062,N_28096,N_25371);
xnor UO_3063 (O_3063,N_25536,N_29458);
nor UO_3064 (O_3064,N_29877,N_29785);
or UO_3065 (O_3065,N_26306,N_26720);
and UO_3066 (O_3066,N_25817,N_26519);
nand UO_3067 (O_3067,N_27653,N_26258);
or UO_3068 (O_3068,N_26081,N_28426);
nor UO_3069 (O_3069,N_29921,N_28493);
xor UO_3070 (O_3070,N_25086,N_26625);
xor UO_3071 (O_3071,N_25483,N_25154);
nor UO_3072 (O_3072,N_28579,N_26987);
xnor UO_3073 (O_3073,N_25328,N_25109);
and UO_3074 (O_3074,N_29982,N_26317);
nor UO_3075 (O_3075,N_25034,N_27945);
xnor UO_3076 (O_3076,N_26116,N_29227);
nor UO_3077 (O_3077,N_29326,N_27613);
or UO_3078 (O_3078,N_28413,N_28467);
and UO_3079 (O_3079,N_25429,N_25995);
xor UO_3080 (O_3080,N_25957,N_27074);
nand UO_3081 (O_3081,N_29461,N_28619);
and UO_3082 (O_3082,N_28125,N_26152);
nand UO_3083 (O_3083,N_28975,N_25677);
xnor UO_3084 (O_3084,N_25016,N_25125);
nand UO_3085 (O_3085,N_29025,N_25575);
nand UO_3086 (O_3086,N_28785,N_27271);
nor UO_3087 (O_3087,N_25590,N_25420);
xnor UO_3088 (O_3088,N_26322,N_26056);
or UO_3089 (O_3089,N_25361,N_28373);
xnor UO_3090 (O_3090,N_26927,N_28814);
nand UO_3091 (O_3091,N_25251,N_26887);
or UO_3092 (O_3092,N_29653,N_27917);
xnor UO_3093 (O_3093,N_29687,N_26017);
or UO_3094 (O_3094,N_28817,N_25695);
nand UO_3095 (O_3095,N_28350,N_29068);
nor UO_3096 (O_3096,N_28413,N_25096);
xnor UO_3097 (O_3097,N_25645,N_29553);
xor UO_3098 (O_3098,N_25384,N_28032);
xor UO_3099 (O_3099,N_28801,N_27909);
nand UO_3100 (O_3100,N_25298,N_27316);
nor UO_3101 (O_3101,N_26482,N_25463);
and UO_3102 (O_3102,N_29982,N_27206);
or UO_3103 (O_3103,N_29979,N_26569);
and UO_3104 (O_3104,N_27769,N_27893);
and UO_3105 (O_3105,N_29396,N_28429);
and UO_3106 (O_3106,N_26862,N_28301);
nor UO_3107 (O_3107,N_27530,N_27729);
nand UO_3108 (O_3108,N_29567,N_27530);
xor UO_3109 (O_3109,N_27233,N_27105);
xor UO_3110 (O_3110,N_28150,N_25065);
or UO_3111 (O_3111,N_26220,N_25877);
nor UO_3112 (O_3112,N_27335,N_25043);
or UO_3113 (O_3113,N_27678,N_29370);
xor UO_3114 (O_3114,N_26808,N_29189);
nor UO_3115 (O_3115,N_25573,N_27708);
and UO_3116 (O_3116,N_25040,N_27072);
xnor UO_3117 (O_3117,N_27083,N_25616);
xor UO_3118 (O_3118,N_26455,N_27514);
and UO_3119 (O_3119,N_26168,N_28617);
nor UO_3120 (O_3120,N_28955,N_28811);
nor UO_3121 (O_3121,N_29062,N_25805);
or UO_3122 (O_3122,N_28159,N_28892);
and UO_3123 (O_3123,N_27793,N_27678);
and UO_3124 (O_3124,N_26056,N_27314);
xor UO_3125 (O_3125,N_26132,N_29114);
or UO_3126 (O_3126,N_29030,N_28600);
nor UO_3127 (O_3127,N_29336,N_25277);
nand UO_3128 (O_3128,N_27251,N_28124);
nand UO_3129 (O_3129,N_29913,N_27731);
and UO_3130 (O_3130,N_29724,N_26175);
and UO_3131 (O_3131,N_25820,N_26298);
nand UO_3132 (O_3132,N_29385,N_25543);
xor UO_3133 (O_3133,N_29144,N_26173);
and UO_3134 (O_3134,N_27933,N_28205);
and UO_3135 (O_3135,N_28854,N_25076);
nand UO_3136 (O_3136,N_29932,N_27416);
or UO_3137 (O_3137,N_28095,N_28748);
nand UO_3138 (O_3138,N_25599,N_26733);
or UO_3139 (O_3139,N_29092,N_27124);
nor UO_3140 (O_3140,N_27952,N_25197);
xnor UO_3141 (O_3141,N_25747,N_28025);
nor UO_3142 (O_3142,N_27347,N_26399);
xor UO_3143 (O_3143,N_29190,N_27734);
or UO_3144 (O_3144,N_28517,N_26619);
nand UO_3145 (O_3145,N_27167,N_26386);
xnor UO_3146 (O_3146,N_27351,N_29505);
nor UO_3147 (O_3147,N_27193,N_26779);
and UO_3148 (O_3148,N_26287,N_27366);
and UO_3149 (O_3149,N_28697,N_25520);
xor UO_3150 (O_3150,N_27891,N_27555);
xor UO_3151 (O_3151,N_26412,N_26202);
xor UO_3152 (O_3152,N_25510,N_25506);
and UO_3153 (O_3153,N_26344,N_25802);
or UO_3154 (O_3154,N_29849,N_25430);
xor UO_3155 (O_3155,N_28277,N_29460);
or UO_3156 (O_3156,N_25187,N_25122);
nand UO_3157 (O_3157,N_26375,N_25429);
nor UO_3158 (O_3158,N_29071,N_27687);
nand UO_3159 (O_3159,N_27267,N_28537);
nand UO_3160 (O_3160,N_26729,N_29777);
and UO_3161 (O_3161,N_26293,N_28451);
or UO_3162 (O_3162,N_25379,N_27788);
and UO_3163 (O_3163,N_27759,N_26395);
nor UO_3164 (O_3164,N_28764,N_28042);
nor UO_3165 (O_3165,N_27154,N_25506);
and UO_3166 (O_3166,N_26980,N_25562);
nand UO_3167 (O_3167,N_25835,N_28540);
nor UO_3168 (O_3168,N_25890,N_29460);
nor UO_3169 (O_3169,N_26884,N_26614);
nand UO_3170 (O_3170,N_25914,N_27032);
nor UO_3171 (O_3171,N_29667,N_27086);
and UO_3172 (O_3172,N_27913,N_28099);
nor UO_3173 (O_3173,N_25119,N_26680);
nor UO_3174 (O_3174,N_29961,N_29387);
nand UO_3175 (O_3175,N_26997,N_28393);
nor UO_3176 (O_3176,N_28605,N_26134);
xor UO_3177 (O_3177,N_27335,N_28715);
nand UO_3178 (O_3178,N_28630,N_25437);
and UO_3179 (O_3179,N_29054,N_28786);
nor UO_3180 (O_3180,N_29394,N_25652);
xnor UO_3181 (O_3181,N_27780,N_25114);
xnor UO_3182 (O_3182,N_29636,N_26181);
xor UO_3183 (O_3183,N_28652,N_26968);
nand UO_3184 (O_3184,N_25038,N_26226);
nor UO_3185 (O_3185,N_26224,N_27471);
xnor UO_3186 (O_3186,N_25710,N_27124);
or UO_3187 (O_3187,N_29124,N_26387);
and UO_3188 (O_3188,N_27312,N_25322);
nor UO_3189 (O_3189,N_25164,N_25902);
and UO_3190 (O_3190,N_28593,N_26271);
nor UO_3191 (O_3191,N_26845,N_27712);
nor UO_3192 (O_3192,N_28405,N_25323);
nor UO_3193 (O_3193,N_25606,N_26726);
and UO_3194 (O_3194,N_26242,N_25161);
and UO_3195 (O_3195,N_28022,N_27692);
xnor UO_3196 (O_3196,N_27475,N_25075);
and UO_3197 (O_3197,N_26918,N_29496);
xor UO_3198 (O_3198,N_26542,N_26195);
xor UO_3199 (O_3199,N_25565,N_26795);
xnor UO_3200 (O_3200,N_29886,N_28682);
nor UO_3201 (O_3201,N_27486,N_25903);
nand UO_3202 (O_3202,N_28804,N_27897);
nand UO_3203 (O_3203,N_25320,N_27703);
and UO_3204 (O_3204,N_28243,N_26067);
and UO_3205 (O_3205,N_26468,N_29242);
and UO_3206 (O_3206,N_28728,N_27571);
nor UO_3207 (O_3207,N_29741,N_26948);
xnor UO_3208 (O_3208,N_26938,N_29269);
nor UO_3209 (O_3209,N_25443,N_27459);
or UO_3210 (O_3210,N_28123,N_25748);
xnor UO_3211 (O_3211,N_25360,N_26956);
nand UO_3212 (O_3212,N_29879,N_27508);
and UO_3213 (O_3213,N_29849,N_28666);
nand UO_3214 (O_3214,N_28454,N_29272);
and UO_3215 (O_3215,N_25962,N_28512);
or UO_3216 (O_3216,N_27668,N_25603);
nand UO_3217 (O_3217,N_27530,N_29787);
nand UO_3218 (O_3218,N_26542,N_27656);
xnor UO_3219 (O_3219,N_26474,N_29635);
and UO_3220 (O_3220,N_29370,N_28870);
xnor UO_3221 (O_3221,N_27654,N_25718);
or UO_3222 (O_3222,N_25006,N_29983);
nor UO_3223 (O_3223,N_25987,N_28781);
nand UO_3224 (O_3224,N_25099,N_28781);
or UO_3225 (O_3225,N_27751,N_29943);
nor UO_3226 (O_3226,N_27243,N_25645);
nand UO_3227 (O_3227,N_28152,N_27678);
or UO_3228 (O_3228,N_27044,N_28624);
or UO_3229 (O_3229,N_26618,N_27662);
nand UO_3230 (O_3230,N_25886,N_25873);
or UO_3231 (O_3231,N_27533,N_25285);
nor UO_3232 (O_3232,N_29034,N_29874);
xor UO_3233 (O_3233,N_26729,N_26570);
nand UO_3234 (O_3234,N_26522,N_27460);
nand UO_3235 (O_3235,N_27713,N_25640);
xor UO_3236 (O_3236,N_25877,N_25264);
and UO_3237 (O_3237,N_26550,N_25035);
or UO_3238 (O_3238,N_25137,N_27235);
nor UO_3239 (O_3239,N_28603,N_28246);
xor UO_3240 (O_3240,N_26282,N_26605);
and UO_3241 (O_3241,N_27593,N_26020);
or UO_3242 (O_3242,N_25282,N_26990);
xor UO_3243 (O_3243,N_27488,N_29373);
and UO_3244 (O_3244,N_28673,N_26388);
xor UO_3245 (O_3245,N_28562,N_26361);
or UO_3246 (O_3246,N_26602,N_26206);
xnor UO_3247 (O_3247,N_25943,N_25604);
nor UO_3248 (O_3248,N_29433,N_27894);
and UO_3249 (O_3249,N_27492,N_28679);
xor UO_3250 (O_3250,N_27375,N_25815);
xnor UO_3251 (O_3251,N_26100,N_25741);
nand UO_3252 (O_3252,N_29425,N_29142);
nor UO_3253 (O_3253,N_25546,N_28400);
nor UO_3254 (O_3254,N_25470,N_26779);
nand UO_3255 (O_3255,N_28238,N_26592);
nand UO_3256 (O_3256,N_29597,N_25873);
or UO_3257 (O_3257,N_25435,N_25025);
nor UO_3258 (O_3258,N_25874,N_28759);
nor UO_3259 (O_3259,N_25061,N_26531);
or UO_3260 (O_3260,N_28597,N_28435);
nand UO_3261 (O_3261,N_29245,N_26273);
and UO_3262 (O_3262,N_26722,N_27867);
and UO_3263 (O_3263,N_29895,N_25268);
nor UO_3264 (O_3264,N_28325,N_28742);
xor UO_3265 (O_3265,N_27402,N_27403);
xor UO_3266 (O_3266,N_28261,N_27496);
and UO_3267 (O_3267,N_28997,N_25052);
xor UO_3268 (O_3268,N_29378,N_29225);
nor UO_3269 (O_3269,N_28775,N_25889);
nand UO_3270 (O_3270,N_26476,N_27605);
nor UO_3271 (O_3271,N_26245,N_29464);
or UO_3272 (O_3272,N_29395,N_26263);
nand UO_3273 (O_3273,N_26946,N_28687);
nand UO_3274 (O_3274,N_27668,N_28824);
or UO_3275 (O_3275,N_29975,N_29267);
nand UO_3276 (O_3276,N_25823,N_26014);
nor UO_3277 (O_3277,N_27648,N_28749);
xor UO_3278 (O_3278,N_25907,N_25791);
or UO_3279 (O_3279,N_25862,N_27386);
nor UO_3280 (O_3280,N_25580,N_27424);
and UO_3281 (O_3281,N_29308,N_29762);
nand UO_3282 (O_3282,N_27715,N_29974);
and UO_3283 (O_3283,N_26191,N_29905);
nand UO_3284 (O_3284,N_27652,N_27950);
nand UO_3285 (O_3285,N_25176,N_26971);
or UO_3286 (O_3286,N_25795,N_29974);
xor UO_3287 (O_3287,N_26075,N_29062);
or UO_3288 (O_3288,N_28061,N_26286);
or UO_3289 (O_3289,N_26770,N_26441);
nor UO_3290 (O_3290,N_25113,N_28838);
or UO_3291 (O_3291,N_28473,N_25474);
or UO_3292 (O_3292,N_26385,N_29882);
xnor UO_3293 (O_3293,N_25396,N_25429);
nand UO_3294 (O_3294,N_27879,N_25768);
or UO_3295 (O_3295,N_27262,N_26788);
and UO_3296 (O_3296,N_26767,N_29737);
nand UO_3297 (O_3297,N_29988,N_29797);
or UO_3298 (O_3298,N_25919,N_25671);
nand UO_3299 (O_3299,N_28282,N_28219);
and UO_3300 (O_3300,N_26501,N_29206);
and UO_3301 (O_3301,N_25750,N_28815);
xnor UO_3302 (O_3302,N_26646,N_28338);
nor UO_3303 (O_3303,N_29302,N_28830);
nand UO_3304 (O_3304,N_27375,N_29090);
and UO_3305 (O_3305,N_26418,N_25116);
xor UO_3306 (O_3306,N_29269,N_27989);
nand UO_3307 (O_3307,N_27991,N_25906);
and UO_3308 (O_3308,N_29627,N_28900);
and UO_3309 (O_3309,N_29238,N_27591);
and UO_3310 (O_3310,N_26487,N_29754);
xor UO_3311 (O_3311,N_27989,N_29472);
or UO_3312 (O_3312,N_28982,N_29974);
nand UO_3313 (O_3313,N_28214,N_27731);
nand UO_3314 (O_3314,N_25269,N_27782);
or UO_3315 (O_3315,N_28986,N_26338);
nand UO_3316 (O_3316,N_28107,N_29854);
xnor UO_3317 (O_3317,N_27135,N_26552);
xnor UO_3318 (O_3318,N_25023,N_27116);
nor UO_3319 (O_3319,N_26883,N_25703);
nand UO_3320 (O_3320,N_29524,N_28056);
and UO_3321 (O_3321,N_26956,N_28888);
nand UO_3322 (O_3322,N_27279,N_28883);
xor UO_3323 (O_3323,N_26691,N_25769);
or UO_3324 (O_3324,N_29921,N_25897);
and UO_3325 (O_3325,N_25989,N_25420);
or UO_3326 (O_3326,N_29450,N_25045);
and UO_3327 (O_3327,N_27126,N_28595);
nand UO_3328 (O_3328,N_26009,N_29299);
or UO_3329 (O_3329,N_29367,N_28060);
nor UO_3330 (O_3330,N_29262,N_28056);
nand UO_3331 (O_3331,N_27391,N_29995);
nor UO_3332 (O_3332,N_27693,N_27257);
and UO_3333 (O_3333,N_29027,N_27916);
and UO_3334 (O_3334,N_29124,N_27070);
or UO_3335 (O_3335,N_26049,N_28508);
nor UO_3336 (O_3336,N_28063,N_26485);
xor UO_3337 (O_3337,N_26233,N_27663);
nand UO_3338 (O_3338,N_27685,N_26495);
nor UO_3339 (O_3339,N_28790,N_26036);
xnor UO_3340 (O_3340,N_26782,N_29485);
xor UO_3341 (O_3341,N_27979,N_26310);
xor UO_3342 (O_3342,N_25899,N_26737);
nor UO_3343 (O_3343,N_27714,N_25675);
nand UO_3344 (O_3344,N_26752,N_28494);
or UO_3345 (O_3345,N_27899,N_27802);
or UO_3346 (O_3346,N_27947,N_26468);
nor UO_3347 (O_3347,N_27524,N_29292);
or UO_3348 (O_3348,N_26670,N_29684);
and UO_3349 (O_3349,N_27758,N_26279);
or UO_3350 (O_3350,N_27442,N_28350);
nand UO_3351 (O_3351,N_26580,N_25123);
xor UO_3352 (O_3352,N_29073,N_28386);
nand UO_3353 (O_3353,N_28093,N_28150);
xnor UO_3354 (O_3354,N_27602,N_28592);
nor UO_3355 (O_3355,N_26361,N_25860);
or UO_3356 (O_3356,N_29507,N_28898);
nand UO_3357 (O_3357,N_27240,N_25358);
and UO_3358 (O_3358,N_27503,N_28210);
and UO_3359 (O_3359,N_28144,N_27768);
xor UO_3360 (O_3360,N_28379,N_27774);
xnor UO_3361 (O_3361,N_26379,N_27470);
nor UO_3362 (O_3362,N_28390,N_27651);
xnor UO_3363 (O_3363,N_27620,N_25358);
or UO_3364 (O_3364,N_25687,N_28029);
nand UO_3365 (O_3365,N_27008,N_26928);
xor UO_3366 (O_3366,N_29264,N_27212);
nand UO_3367 (O_3367,N_29420,N_25692);
and UO_3368 (O_3368,N_29985,N_27881);
xor UO_3369 (O_3369,N_28781,N_28710);
nor UO_3370 (O_3370,N_25075,N_25115);
nor UO_3371 (O_3371,N_26486,N_27048);
nand UO_3372 (O_3372,N_27414,N_26694);
nand UO_3373 (O_3373,N_27274,N_26283);
nor UO_3374 (O_3374,N_25934,N_28721);
nand UO_3375 (O_3375,N_29556,N_26266);
xnor UO_3376 (O_3376,N_26547,N_27898);
nor UO_3377 (O_3377,N_25428,N_28202);
nand UO_3378 (O_3378,N_29336,N_25221);
xnor UO_3379 (O_3379,N_25041,N_26730);
nand UO_3380 (O_3380,N_27514,N_25993);
or UO_3381 (O_3381,N_25809,N_29764);
and UO_3382 (O_3382,N_28849,N_27262);
and UO_3383 (O_3383,N_27850,N_29427);
or UO_3384 (O_3384,N_28244,N_25965);
and UO_3385 (O_3385,N_27155,N_26985);
xnor UO_3386 (O_3386,N_25153,N_28709);
nor UO_3387 (O_3387,N_25764,N_26382);
or UO_3388 (O_3388,N_26862,N_29864);
and UO_3389 (O_3389,N_29230,N_26499);
or UO_3390 (O_3390,N_29978,N_28072);
or UO_3391 (O_3391,N_26253,N_25363);
nand UO_3392 (O_3392,N_28509,N_26108);
xor UO_3393 (O_3393,N_25570,N_25787);
and UO_3394 (O_3394,N_27126,N_26652);
nand UO_3395 (O_3395,N_26579,N_29871);
nor UO_3396 (O_3396,N_29801,N_29206);
xnor UO_3397 (O_3397,N_27687,N_26407);
nand UO_3398 (O_3398,N_29372,N_25032);
nand UO_3399 (O_3399,N_28278,N_29204);
or UO_3400 (O_3400,N_28812,N_28772);
or UO_3401 (O_3401,N_28860,N_29081);
xnor UO_3402 (O_3402,N_25485,N_29706);
xnor UO_3403 (O_3403,N_29199,N_25451);
nor UO_3404 (O_3404,N_26004,N_29026);
and UO_3405 (O_3405,N_28158,N_29866);
xnor UO_3406 (O_3406,N_26952,N_28371);
or UO_3407 (O_3407,N_26055,N_27256);
nor UO_3408 (O_3408,N_27457,N_26167);
nand UO_3409 (O_3409,N_26222,N_25574);
or UO_3410 (O_3410,N_27493,N_25127);
or UO_3411 (O_3411,N_25384,N_29400);
and UO_3412 (O_3412,N_25210,N_28144);
nor UO_3413 (O_3413,N_28153,N_27568);
xor UO_3414 (O_3414,N_29071,N_28250);
nor UO_3415 (O_3415,N_28457,N_29272);
or UO_3416 (O_3416,N_29341,N_29739);
and UO_3417 (O_3417,N_28091,N_25232);
nand UO_3418 (O_3418,N_27117,N_29891);
and UO_3419 (O_3419,N_28284,N_27534);
and UO_3420 (O_3420,N_28858,N_26872);
xor UO_3421 (O_3421,N_25632,N_26821);
and UO_3422 (O_3422,N_27534,N_26592);
xnor UO_3423 (O_3423,N_28133,N_27869);
or UO_3424 (O_3424,N_27688,N_25904);
xor UO_3425 (O_3425,N_26385,N_27267);
and UO_3426 (O_3426,N_29337,N_25375);
xnor UO_3427 (O_3427,N_29445,N_25712);
or UO_3428 (O_3428,N_29160,N_29968);
nand UO_3429 (O_3429,N_27531,N_28593);
or UO_3430 (O_3430,N_26280,N_26516);
or UO_3431 (O_3431,N_27514,N_27294);
and UO_3432 (O_3432,N_29393,N_27114);
or UO_3433 (O_3433,N_26133,N_25876);
or UO_3434 (O_3434,N_27971,N_25504);
nand UO_3435 (O_3435,N_29306,N_27327);
or UO_3436 (O_3436,N_27696,N_28920);
xnor UO_3437 (O_3437,N_25106,N_28066);
nor UO_3438 (O_3438,N_25787,N_26011);
nor UO_3439 (O_3439,N_26575,N_26449);
nor UO_3440 (O_3440,N_25280,N_28659);
or UO_3441 (O_3441,N_28880,N_29673);
nor UO_3442 (O_3442,N_25832,N_27371);
and UO_3443 (O_3443,N_25254,N_27360);
and UO_3444 (O_3444,N_26289,N_27337);
xor UO_3445 (O_3445,N_26100,N_26645);
nor UO_3446 (O_3446,N_29944,N_29319);
or UO_3447 (O_3447,N_25337,N_29627);
and UO_3448 (O_3448,N_29120,N_29863);
nor UO_3449 (O_3449,N_27208,N_28952);
xor UO_3450 (O_3450,N_29913,N_26936);
or UO_3451 (O_3451,N_27408,N_28931);
nand UO_3452 (O_3452,N_28973,N_29699);
and UO_3453 (O_3453,N_27259,N_28119);
nand UO_3454 (O_3454,N_28078,N_29564);
or UO_3455 (O_3455,N_26478,N_29846);
nor UO_3456 (O_3456,N_29131,N_27447);
and UO_3457 (O_3457,N_26274,N_25778);
nand UO_3458 (O_3458,N_25710,N_28604);
xor UO_3459 (O_3459,N_27143,N_28103);
nor UO_3460 (O_3460,N_25838,N_26065);
or UO_3461 (O_3461,N_28099,N_26408);
or UO_3462 (O_3462,N_25751,N_29510);
nand UO_3463 (O_3463,N_28872,N_28300);
nor UO_3464 (O_3464,N_29042,N_29903);
xnor UO_3465 (O_3465,N_29269,N_29201);
nor UO_3466 (O_3466,N_26882,N_25670);
nor UO_3467 (O_3467,N_28275,N_27716);
nand UO_3468 (O_3468,N_29487,N_28308);
nor UO_3469 (O_3469,N_25171,N_25821);
xnor UO_3470 (O_3470,N_25361,N_28645);
nand UO_3471 (O_3471,N_28801,N_29524);
and UO_3472 (O_3472,N_28497,N_28890);
and UO_3473 (O_3473,N_27538,N_25651);
nor UO_3474 (O_3474,N_28029,N_26013);
or UO_3475 (O_3475,N_28711,N_26489);
xnor UO_3476 (O_3476,N_29447,N_29767);
or UO_3477 (O_3477,N_27427,N_27838);
nor UO_3478 (O_3478,N_28328,N_26325);
nor UO_3479 (O_3479,N_25216,N_29585);
or UO_3480 (O_3480,N_26902,N_29035);
nand UO_3481 (O_3481,N_26110,N_25347);
and UO_3482 (O_3482,N_26327,N_27388);
xor UO_3483 (O_3483,N_27226,N_25535);
or UO_3484 (O_3484,N_28690,N_25768);
nor UO_3485 (O_3485,N_28533,N_29523);
xor UO_3486 (O_3486,N_25882,N_25462);
and UO_3487 (O_3487,N_27332,N_27374);
or UO_3488 (O_3488,N_28311,N_28697);
or UO_3489 (O_3489,N_26925,N_26087);
nand UO_3490 (O_3490,N_28218,N_29551);
nand UO_3491 (O_3491,N_29862,N_28840);
xor UO_3492 (O_3492,N_28450,N_26333);
xor UO_3493 (O_3493,N_25050,N_28986);
or UO_3494 (O_3494,N_27247,N_26394);
xnor UO_3495 (O_3495,N_28270,N_29045);
and UO_3496 (O_3496,N_26255,N_28692);
and UO_3497 (O_3497,N_27293,N_29918);
xnor UO_3498 (O_3498,N_27892,N_25498);
nand UO_3499 (O_3499,N_27731,N_29243);
endmodule