module basic_500_3000_500_4_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_100,In_387);
nor U1 (N_1,In_168,In_282);
nand U2 (N_2,In_226,In_225);
xor U3 (N_3,In_390,In_362);
nor U4 (N_4,In_359,In_244);
nand U5 (N_5,In_140,In_292);
nor U6 (N_6,In_323,In_399);
nand U7 (N_7,In_178,In_305);
xor U8 (N_8,In_254,In_435);
nor U9 (N_9,In_147,In_122);
or U10 (N_10,In_21,In_398);
or U11 (N_11,In_407,In_162);
nor U12 (N_12,In_106,In_396);
and U13 (N_13,In_316,In_330);
and U14 (N_14,In_159,In_291);
xnor U15 (N_15,In_319,In_146);
or U16 (N_16,In_44,In_329);
nand U17 (N_17,In_496,In_184);
xor U18 (N_18,In_246,In_462);
and U19 (N_19,In_322,In_203);
nor U20 (N_20,In_361,In_43);
and U21 (N_21,In_190,In_348);
xor U22 (N_22,In_149,In_321);
nand U23 (N_23,In_125,In_6);
xor U24 (N_24,In_448,In_80);
and U25 (N_25,In_13,In_299);
and U26 (N_26,In_290,In_74);
and U27 (N_27,In_369,In_341);
nand U28 (N_28,In_377,In_9);
nor U29 (N_29,In_12,In_55);
nand U30 (N_30,In_423,In_453);
nand U31 (N_31,In_183,In_495);
and U32 (N_32,In_429,In_351);
nor U33 (N_33,In_481,In_5);
nand U34 (N_34,In_438,In_163);
xnor U35 (N_35,In_179,In_175);
nor U36 (N_36,In_67,In_284);
xor U37 (N_37,In_86,In_275);
or U38 (N_38,In_54,In_93);
and U39 (N_39,In_451,In_214);
nor U40 (N_40,In_280,In_199);
or U41 (N_41,In_486,In_216);
nor U42 (N_42,In_132,In_70);
nand U43 (N_43,In_16,In_381);
nand U44 (N_44,In_27,In_219);
xor U45 (N_45,In_334,In_490);
or U46 (N_46,In_176,In_118);
and U47 (N_47,In_213,In_402);
or U48 (N_48,In_157,In_430);
xnor U49 (N_49,In_343,In_456);
nand U50 (N_50,In_392,In_302);
nor U51 (N_51,In_131,In_272);
or U52 (N_52,In_289,In_10);
or U53 (N_53,In_364,In_459);
nor U54 (N_54,In_307,In_276);
xnor U55 (N_55,In_57,In_136);
xor U56 (N_56,In_35,In_463);
or U57 (N_57,In_354,In_95);
nor U58 (N_58,In_77,In_360);
and U59 (N_59,In_473,In_248);
or U60 (N_60,In_38,In_241);
xor U61 (N_61,In_417,In_26);
nor U62 (N_62,In_471,In_220);
or U63 (N_63,In_209,In_313);
nand U64 (N_64,In_328,In_293);
xnor U65 (N_65,In_224,In_439);
nor U66 (N_66,In_105,In_151);
or U67 (N_67,In_294,In_240);
xor U68 (N_68,In_156,In_185);
xnor U69 (N_69,In_180,In_452);
or U70 (N_70,In_267,In_342);
and U71 (N_71,In_412,In_22);
nand U72 (N_72,In_484,In_123);
xor U73 (N_73,In_62,In_20);
xnor U74 (N_74,In_424,In_194);
xor U75 (N_75,In_264,In_266);
and U76 (N_76,In_251,In_90);
nor U77 (N_77,In_455,In_346);
xnor U78 (N_78,In_450,In_25);
or U79 (N_79,In_464,In_60);
and U80 (N_80,In_207,In_262);
nand U81 (N_81,In_11,In_258);
or U82 (N_82,In_8,In_18);
xnor U83 (N_83,In_245,In_212);
and U84 (N_84,In_4,In_477);
xor U85 (N_85,In_375,In_337);
and U86 (N_86,In_152,In_68);
or U87 (N_87,In_7,In_204);
nand U88 (N_88,In_483,In_432);
xor U89 (N_89,In_431,In_201);
nand U90 (N_90,In_187,In_482);
and U91 (N_91,In_99,In_130);
xor U92 (N_92,In_139,In_102);
or U93 (N_93,In_253,In_72);
nor U94 (N_94,In_470,In_278);
and U95 (N_95,In_161,In_263);
nor U96 (N_96,In_103,In_104);
nor U97 (N_97,In_303,In_332);
or U98 (N_98,In_457,In_494);
xnor U99 (N_99,In_380,In_306);
nand U100 (N_100,In_206,In_368);
nor U101 (N_101,In_189,In_311);
or U102 (N_102,In_465,In_41);
xor U103 (N_103,In_52,In_120);
nand U104 (N_104,In_79,In_59);
or U105 (N_105,In_141,In_37);
xnor U106 (N_106,In_223,In_304);
or U107 (N_107,In_405,In_480);
nor U108 (N_108,In_394,In_409);
xnor U109 (N_109,In_325,In_217);
or U110 (N_110,In_138,In_458);
or U111 (N_111,In_443,In_107);
nand U112 (N_112,In_49,In_478);
or U113 (N_113,In_447,In_273);
and U114 (N_114,In_286,In_234);
nor U115 (N_115,In_476,In_376);
and U116 (N_116,In_42,In_265);
and U117 (N_117,In_47,In_356);
nor U118 (N_118,In_296,In_411);
nor U119 (N_119,In_171,In_421);
and U120 (N_120,In_249,In_188);
nor U121 (N_121,In_378,In_488);
xor U122 (N_122,In_434,In_413);
nand U123 (N_123,In_472,In_349);
xnor U124 (N_124,In_418,In_269);
or U125 (N_125,In_479,In_250);
nand U126 (N_126,In_193,In_256);
nor U127 (N_127,In_14,In_98);
xnor U128 (N_128,In_24,In_338);
and U129 (N_129,In_200,In_40);
xor U130 (N_130,In_371,In_144);
xor U131 (N_131,In_285,In_358);
and U132 (N_132,In_333,In_404);
nor U133 (N_133,In_135,In_196);
xor U134 (N_134,In_255,In_382);
nand U135 (N_135,In_274,In_56);
nor U136 (N_136,In_485,In_314);
xor U137 (N_137,In_31,In_46);
or U138 (N_138,In_350,In_487);
or U139 (N_139,In_133,In_383);
and U140 (N_140,In_208,In_395);
or U141 (N_141,In_230,In_89);
or U142 (N_142,In_239,In_119);
nor U143 (N_143,In_357,In_397);
xnor U144 (N_144,In_23,In_379);
nor U145 (N_145,In_493,In_1);
or U146 (N_146,In_489,In_422);
nor U147 (N_147,In_372,In_83);
and U148 (N_148,In_327,In_344);
and U149 (N_149,In_50,In_96);
nor U150 (N_150,In_449,In_320);
nand U151 (N_151,In_66,In_0);
or U152 (N_152,In_425,In_177);
xor U153 (N_153,In_416,In_326);
or U154 (N_154,In_15,In_352);
or U155 (N_155,In_36,In_270);
and U156 (N_156,In_17,In_331);
nand U157 (N_157,In_384,In_69);
nor U158 (N_158,In_257,In_137);
or U159 (N_159,In_259,In_353);
xor U160 (N_160,In_437,In_169);
xor U161 (N_161,In_410,In_153);
xnor U162 (N_162,In_128,In_82);
nor U163 (N_163,In_114,In_115);
xor U164 (N_164,In_288,In_497);
and U165 (N_165,In_295,In_433);
or U166 (N_166,In_242,In_324);
nand U167 (N_167,In_406,In_181);
nor U168 (N_168,In_460,In_142);
or U169 (N_169,In_155,In_88);
nor U170 (N_170,In_94,In_475);
nand U171 (N_171,In_440,In_143);
nor U172 (N_172,In_76,In_312);
nand U173 (N_173,In_126,In_309);
nand U174 (N_174,In_491,In_370);
nand U175 (N_175,In_414,In_283);
or U176 (N_176,In_391,In_297);
and U177 (N_177,In_197,In_363);
xor U178 (N_178,In_347,In_393);
and U179 (N_179,In_243,In_191);
and U180 (N_180,In_237,In_474);
nor U181 (N_181,In_173,In_164);
nand U182 (N_182,In_277,In_221);
nand U183 (N_183,In_29,In_335);
xor U184 (N_184,In_172,In_415);
nor U185 (N_185,In_174,In_45);
nand U186 (N_186,In_75,In_150);
nand U187 (N_187,In_64,In_444);
and U188 (N_188,In_218,In_63);
and U189 (N_189,In_116,In_428);
nor U190 (N_190,In_365,In_236);
nand U191 (N_191,In_461,In_2);
nand U192 (N_192,In_227,In_260);
nor U193 (N_193,In_233,In_110);
and U194 (N_194,In_252,In_81);
and U195 (N_195,In_192,In_71);
nand U196 (N_196,In_318,In_401);
nand U197 (N_197,In_310,In_367);
and U198 (N_198,In_129,In_202);
nand U199 (N_199,In_33,In_373);
nand U200 (N_200,In_385,In_400);
xnor U201 (N_201,In_108,In_408);
nor U202 (N_202,In_61,In_420);
or U203 (N_203,In_232,In_186);
or U204 (N_204,In_134,In_281);
xor U205 (N_205,In_84,In_469);
or U206 (N_206,In_298,In_231);
xnor U207 (N_207,In_468,In_148);
nand U208 (N_208,In_235,In_182);
and U209 (N_209,In_101,In_467);
nand U210 (N_210,In_34,In_211);
and U211 (N_211,In_78,In_441);
xor U212 (N_212,In_336,In_73);
xor U213 (N_213,In_268,In_121);
and U214 (N_214,In_85,In_386);
and U215 (N_215,In_345,In_53);
xor U216 (N_216,In_160,In_97);
xor U217 (N_217,In_222,In_51);
and U218 (N_218,In_158,In_127);
nand U219 (N_219,In_58,In_446);
or U220 (N_220,In_32,In_205);
xnor U221 (N_221,In_109,In_166);
nor U222 (N_222,In_198,In_287);
and U223 (N_223,In_145,In_65);
and U224 (N_224,In_403,In_315);
nor U225 (N_225,In_374,In_492);
and U226 (N_226,In_339,In_317);
nand U227 (N_227,In_426,In_301);
or U228 (N_228,In_48,In_366);
and U229 (N_229,In_39,In_113);
nor U230 (N_230,In_229,In_340);
or U231 (N_231,In_195,In_466);
nor U232 (N_232,In_442,In_427);
nand U233 (N_233,In_300,In_308);
nand U234 (N_234,In_92,In_170);
nand U235 (N_235,In_261,In_124);
or U236 (N_236,In_210,In_117);
nand U237 (N_237,In_498,In_271);
and U238 (N_238,In_499,In_279);
xor U239 (N_239,In_228,In_215);
or U240 (N_240,In_419,In_247);
and U241 (N_241,In_454,In_112);
or U242 (N_242,In_445,In_111);
and U243 (N_243,In_436,In_165);
or U244 (N_244,In_388,In_167);
or U245 (N_245,In_19,In_355);
nor U246 (N_246,In_3,In_91);
or U247 (N_247,In_30,In_87);
xor U248 (N_248,In_238,In_28);
xnor U249 (N_249,In_389,In_154);
or U250 (N_250,In_171,In_466);
xnor U251 (N_251,In_389,In_443);
nand U252 (N_252,In_300,In_165);
or U253 (N_253,In_184,In_190);
and U254 (N_254,In_269,In_298);
and U255 (N_255,In_37,In_348);
nand U256 (N_256,In_399,In_85);
nand U257 (N_257,In_311,In_162);
nor U258 (N_258,In_103,In_383);
and U259 (N_259,In_53,In_136);
nor U260 (N_260,In_31,In_405);
nand U261 (N_261,In_111,In_363);
or U262 (N_262,In_228,In_410);
nand U263 (N_263,In_288,In_379);
nor U264 (N_264,In_221,In_79);
nor U265 (N_265,In_32,In_2);
xnor U266 (N_266,In_406,In_237);
xor U267 (N_267,In_206,In_418);
nand U268 (N_268,In_433,In_363);
or U269 (N_269,In_381,In_193);
nor U270 (N_270,In_371,In_117);
nor U271 (N_271,In_72,In_170);
or U272 (N_272,In_320,In_299);
xnor U273 (N_273,In_486,In_458);
nor U274 (N_274,In_332,In_451);
xor U275 (N_275,In_310,In_249);
and U276 (N_276,In_70,In_84);
nand U277 (N_277,In_125,In_111);
nor U278 (N_278,In_178,In_279);
nand U279 (N_279,In_82,In_9);
xnor U280 (N_280,In_87,In_316);
nor U281 (N_281,In_201,In_35);
nor U282 (N_282,In_364,In_387);
or U283 (N_283,In_358,In_425);
nor U284 (N_284,In_111,In_309);
or U285 (N_285,In_75,In_338);
nor U286 (N_286,In_107,In_54);
and U287 (N_287,In_355,In_431);
or U288 (N_288,In_144,In_393);
xnor U289 (N_289,In_208,In_162);
or U290 (N_290,In_265,In_121);
nand U291 (N_291,In_198,In_211);
nor U292 (N_292,In_56,In_425);
nand U293 (N_293,In_226,In_148);
and U294 (N_294,In_394,In_219);
and U295 (N_295,In_312,In_127);
or U296 (N_296,In_298,In_189);
xnor U297 (N_297,In_457,In_220);
or U298 (N_298,In_111,In_489);
nor U299 (N_299,In_167,In_275);
nand U300 (N_300,In_283,In_114);
nor U301 (N_301,In_87,In_109);
nor U302 (N_302,In_474,In_185);
xor U303 (N_303,In_373,In_356);
xor U304 (N_304,In_251,In_81);
nor U305 (N_305,In_373,In_371);
and U306 (N_306,In_79,In_310);
xor U307 (N_307,In_220,In_344);
nand U308 (N_308,In_451,In_43);
nor U309 (N_309,In_299,In_445);
or U310 (N_310,In_238,In_416);
nand U311 (N_311,In_37,In_214);
or U312 (N_312,In_109,In_55);
or U313 (N_313,In_452,In_321);
or U314 (N_314,In_256,In_105);
xor U315 (N_315,In_431,In_169);
nand U316 (N_316,In_57,In_458);
nand U317 (N_317,In_250,In_367);
nand U318 (N_318,In_361,In_436);
or U319 (N_319,In_170,In_468);
or U320 (N_320,In_285,In_444);
nor U321 (N_321,In_324,In_464);
xor U322 (N_322,In_444,In_113);
xor U323 (N_323,In_395,In_433);
xnor U324 (N_324,In_328,In_348);
or U325 (N_325,In_355,In_60);
nor U326 (N_326,In_177,In_223);
xnor U327 (N_327,In_125,In_445);
nor U328 (N_328,In_314,In_482);
xor U329 (N_329,In_151,In_462);
or U330 (N_330,In_203,In_310);
xor U331 (N_331,In_258,In_57);
nor U332 (N_332,In_120,In_437);
and U333 (N_333,In_266,In_179);
or U334 (N_334,In_453,In_360);
xnor U335 (N_335,In_286,In_495);
nor U336 (N_336,In_28,In_366);
or U337 (N_337,In_86,In_254);
nand U338 (N_338,In_45,In_359);
and U339 (N_339,In_120,In_66);
and U340 (N_340,In_472,In_150);
or U341 (N_341,In_14,In_408);
nand U342 (N_342,In_6,In_207);
and U343 (N_343,In_410,In_450);
xor U344 (N_344,In_58,In_461);
xnor U345 (N_345,In_50,In_36);
or U346 (N_346,In_222,In_260);
or U347 (N_347,In_492,In_133);
xnor U348 (N_348,In_454,In_188);
and U349 (N_349,In_215,In_72);
nor U350 (N_350,In_252,In_288);
and U351 (N_351,In_55,In_16);
nor U352 (N_352,In_106,In_22);
nand U353 (N_353,In_274,In_345);
and U354 (N_354,In_203,In_426);
and U355 (N_355,In_261,In_240);
nand U356 (N_356,In_298,In_15);
and U357 (N_357,In_279,In_436);
or U358 (N_358,In_421,In_451);
nor U359 (N_359,In_313,In_72);
xor U360 (N_360,In_30,In_60);
or U361 (N_361,In_235,In_92);
and U362 (N_362,In_234,In_4);
nor U363 (N_363,In_156,In_250);
and U364 (N_364,In_284,In_443);
or U365 (N_365,In_496,In_181);
and U366 (N_366,In_315,In_455);
and U367 (N_367,In_485,In_126);
and U368 (N_368,In_358,In_112);
nand U369 (N_369,In_492,In_92);
nor U370 (N_370,In_335,In_350);
or U371 (N_371,In_497,In_118);
xnor U372 (N_372,In_16,In_289);
nor U373 (N_373,In_400,In_162);
or U374 (N_374,In_241,In_271);
or U375 (N_375,In_339,In_120);
and U376 (N_376,In_46,In_194);
and U377 (N_377,In_281,In_18);
xor U378 (N_378,In_47,In_12);
and U379 (N_379,In_314,In_379);
nor U380 (N_380,In_321,In_488);
nand U381 (N_381,In_266,In_359);
xnor U382 (N_382,In_244,In_420);
nor U383 (N_383,In_441,In_229);
nand U384 (N_384,In_30,In_280);
xor U385 (N_385,In_254,In_79);
or U386 (N_386,In_151,In_160);
or U387 (N_387,In_52,In_299);
xnor U388 (N_388,In_93,In_389);
and U389 (N_389,In_203,In_419);
nand U390 (N_390,In_74,In_252);
or U391 (N_391,In_484,In_165);
or U392 (N_392,In_348,In_383);
xor U393 (N_393,In_304,In_192);
and U394 (N_394,In_57,In_248);
nand U395 (N_395,In_114,In_128);
nand U396 (N_396,In_146,In_7);
nand U397 (N_397,In_477,In_405);
and U398 (N_398,In_329,In_235);
and U399 (N_399,In_116,In_425);
nand U400 (N_400,In_166,In_201);
and U401 (N_401,In_87,In_428);
xor U402 (N_402,In_147,In_38);
xnor U403 (N_403,In_411,In_238);
and U404 (N_404,In_34,In_149);
and U405 (N_405,In_282,In_374);
nand U406 (N_406,In_118,In_172);
xor U407 (N_407,In_438,In_450);
or U408 (N_408,In_211,In_425);
nor U409 (N_409,In_451,In_277);
or U410 (N_410,In_157,In_213);
and U411 (N_411,In_250,In_119);
nand U412 (N_412,In_27,In_41);
or U413 (N_413,In_137,In_139);
or U414 (N_414,In_67,In_339);
nor U415 (N_415,In_31,In_142);
and U416 (N_416,In_251,In_89);
and U417 (N_417,In_91,In_403);
or U418 (N_418,In_476,In_364);
and U419 (N_419,In_287,In_136);
nor U420 (N_420,In_261,In_17);
nand U421 (N_421,In_433,In_159);
xor U422 (N_422,In_449,In_292);
xnor U423 (N_423,In_181,In_43);
or U424 (N_424,In_75,In_394);
nand U425 (N_425,In_313,In_238);
xor U426 (N_426,In_342,In_325);
or U427 (N_427,In_69,In_479);
nand U428 (N_428,In_414,In_174);
nand U429 (N_429,In_197,In_253);
nand U430 (N_430,In_117,In_431);
and U431 (N_431,In_356,In_393);
nor U432 (N_432,In_307,In_271);
and U433 (N_433,In_85,In_165);
nor U434 (N_434,In_387,In_418);
nand U435 (N_435,In_370,In_136);
nor U436 (N_436,In_466,In_410);
or U437 (N_437,In_278,In_499);
nand U438 (N_438,In_28,In_202);
nand U439 (N_439,In_324,In_195);
or U440 (N_440,In_87,In_96);
xnor U441 (N_441,In_170,In_336);
and U442 (N_442,In_458,In_106);
nor U443 (N_443,In_182,In_76);
or U444 (N_444,In_385,In_15);
or U445 (N_445,In_494,In_332);
nor U446 (N_446,In_337,In_220);
and U447 (N_447,In_115,In_428);
nor U448 (N_448,In_401,In_290);
nand U449 (N_449,In_399,In_367);
nand U450 (N_450,In_26,In_471);
nor U451 (N_451,In_52,In_192);
nand U452 (N_452,In_62,In_369);
xnor U453 (N_453,In_261,In_181);
nor U454 (N_454,In_117,In_357);
and U455 (N_455,In_472,In_385);
nor U456 (N_456,In_237,In_380);
nand U457 (N_457,In_350,In_266);
nor U458 (N_458,In_136,In_225);
nand U459 (N_459,In_224,In_5);
xor U460 (N_460,In_286,In_161);
nor U461 (N_461,In_143,In_316);
or U462 (N_462,In_64,In_252);
nor U463 (N_463,In_59,In_399);
nand U464 (N_464,In_448,In_88);
nor U465 (N_465,In_162,In_55);
and U466 (N_466,In_326,In_437);
nand U467 (N_467,In_163,In_48);
or U468 (N_468,In_383,In_293);
nand U469 (N_469,In_285,In_164);
xor U470 (N_470,In_204,In_123);
nor U471 (N_471,In_171,In_266);
nor U472 (N_472,In_222,In_364);
nand U473 (N_473,In_315,In_338);
or U474 (N_474,In_346,In_360);
nor U475 (N_475,In_242,In_292);
nand U476 (N_476,In_53,In_362);
xor U477 (N_477,In_425,In_73);
nor U478 (N_478,In_46,In_92);
nor U479 (N_479,In_272,In_480);
or U480 (N_480,In_423,In_257);
or U481 (N_481,In_400,In_113);
and U482 (N_482,In_50,In_161);
and U483 (N_483,In_290,In_321);
xnor U484 (N_484,In_201,In_105);
nor U485 (N_485,In_422,In_378);
and U486 (N_486,In_453,In_45);
or U487 (N_487,In_459,In_499);
and U488 (N_488,In_199,In_343);
nand U489 (N_489,In_257,In_487);
or U490 (N_490,In_113,In_384);
and U491 (N_491,In_487,In_162);
nor U492 (N_492,In_160,In_57);
nand U493 (N_493,In_354,In_61);
or U494 (N_494,In_225,In_480);
nand U495 (N_495,In_350,In_24);
and U496 (N_496,In_144,In_455);
and U497 (N_497,In_382,In_355);
or U498 (N_498,In_413,In_266);
nor U499 (N_499,In_228,In_61);
or U500 (N_500,In_374,In_168);
or U501 (N_501,In_229,In_475);
nand U502 (N_502,In_312,In_372);
xor U503 (N_503,In_441,In_80);
and U504 (N_504,In_108,In_420);
and U505 (N_505,In_328,In_337);
and U506 (N_506,In_110,In_362);
nand U507 (N_507,In_39,In_131);
or U508 (N_508,In_173,In_28);
or U509 (N_509,In_225,In_187);
or U510 (N_510,In_462,In_41);
or U511 (N_511,In_474,In_24);
nor U512 (N_512,In_288,In_476);
or U513 (N_513,In_132,In_197);
nor U514 (N_514,In_128,In_47);
and U515 (N_515,In_98,In_435);
nor U516 (N_516,In_185,In_47);
xor U517 (N_517,In_298,In_314);
nor U518 (N_518,In_415,In_395);
nor U519 (N_519,In_406,In_102);
and U520 (N_520,In_286,In_28);
nand U521 (N_521,In_272,In_204);
or U522 (N_522,In_387,In_94);
nor U523 (N_523,In_272,In_395);
and U524 (N_524,In_451,In_285);
and U525 (N_525,In_168,In_152);
and U526 (N_526,In_284,In_337);
or U527 (N_527,In_272,In_439);
and U528 (N_528,In_442,In_87);
nor U529 (N_529,In_158,In_172);
or U530 (N_530,In_60,In_73);
nor U531 (N_531,In_124,In_115);
nor U532 (N_532,In_206,In_431);
nor U533 (N_533,In_441,In_346);
or U534 (N_534,In_193,In_89);
nand U535 (N_535,In_328,In_53);
or U536 (N_536,In_180,In_86);
nand U537 (N_537,In_296,In_91);
and U538 (N_538,In_210,In_389);
xnor U539 (N_539,In_344,In_246);
and U540 (N_540,In_396,In_156);
nand U541 (N_541,In_338,In_325);
nand U542 (N_542,In_387,In_45);
nor U543 (N_543,In_148,In_326);
and U544 (N_544,In_458,In_351);
and U545 (N_545,In_22,In_323);
and U546 (N_546,In_26,In_260);
and U547 (N_547,In_201,In_383);
and U548 (N_548,In_310,In_294);
xor U549 (N_549,In_291,In_287);
nand U550 (N_550,In_102,In_138);
nor U551 (N_551,In_393,In_412);
nand U552 (N_552,In_385,In_268);
nand U553 (N_553,In_479,In_307);
and U554 (N_554,In_17,In_408);
nand U555 (N_555,In_429,In_90);
nor U556 (N_556,In_314,In_448);
nand U557 (N_557,In_279,In_51);
nand U558 (N_558,In_267,In_281);
and U559 (N_559,In_71,In_483);
nand U560 (N_560,In_405,In_226);
xnor U561 (N_561,In_32,In_121);
nor U562 (N_562,In_172,In_198);
xor U563 (N_563,In_189,In_153);
xnor U564 (N_564,In_272,In_489);
or U565 (N_565,In_63,In_490);
or U566 (N_566,In_243,In_370);
or U567 (N_567,In_184,In_366);
and U568 (N_568,In_411,In_208);
xnor U569 (N_569,In_42,In_463);
nand U570 (N_570,In_468,In_283);
nor U571 (N_571,In_266,In_24);
nor U572 (N_572,In_410,In_235);
and U573 (N_573,In_399,In_474);
and U574 (N_574,In_154,In_338);
or U575 (N_575,In_138,In_438);
nand U576 (N_576,In_312,In_205);
or U577 (N_577,In_39,In_198);
nand U578 (N_578,In_88,In_134);
or U579 (N_579,In_315,In_105);
nor U580 (N_580,In_377,In_119);
or U581 (N_581,In_184,In_106);
xnor U582 (N_582,In_472,In_201);
or U583 (N_583,In_83,In_485);
xor U584 (N_584,In_48,In_57);
or U585 (N_585,In_198,In_297);
xnor U586 (N_586,In_68,In_197);
nand U587 (N_587,In_432,In_46);
and U588 (N_588,In_443,In_124);
nand U589 (N_589,In_16,In_258);
xnor U590 (N_590,In_34,In_75);
xor U591 (N_591,In_91,In_351);
and U592 (N_592,In_262,In_461);
nand U593 (N_593,In_216,In_56);
and U594 (N_594,In_73,In_38);
nor U595 (N_595,In_56,In_80);
nor U596 (N_596,In_309,In_453);
nand U597 (N_597,In_0,In_265);
and U598 (N_598,In_228,In_123);
nor U599 (N_599,In_63,In_387);
xor U600 (N_600,In_247,In_243);
xnor U601 (N_601,In_394,In_428);
nor U602 (N_602,In_40,In_37);
xor U603 (N_603,In_142,In_322);
or U604 (N_604,In_91,In_486);
and U605 (N_605,In_53,In_51);
or U606 (N_606,In_284,In_9);
and U607 (N_607,In_453,In_153);
nor U608 (N_608,In_146,In_89);
or U609 (N_609,In_222,In_219);
xnor U610 (N_610,In_396,In_395);
nand U611 (N_611,In_414,In_81);
nand U612 (N_612,In_338,In_226);
or U613 (N_613,In_156,In_337);
nor U614 (N_614,In_384,In_63);
nand U615 (N_615,In_318,In_406);
xnor U616 (N_616,In_272,In_457);
and U617 (N_617,In_429,In_360);
nand U618 (N_618,In_10,In_376);
or U619 (N_619,In_230,In_109);
xor U620 (N_620,In_371,In_309);
nor U621 (N_621,In_412,In_277);
and U622 (N_622,In_29,In_367);
or U623 (N_623,In_375,In_410);
nand U624 (N_624,In_174,In_125);
nand U625 (N_625,In_250,In_208);
nand U626 (N_626,In_368,In_140);
and U627 (N_627,In_241,In_368);
or U628 (N_628,In_450,In_7);
nor U629 (N_629,In_325,In_319);
nand U630 (N_630,In_455,In_140);
xor U631 (N_631,In_216,In_28);
nand U632 (N_632,In_27,In_449);
or U633 (N_633,In_225,In_172);
and U634 (N_634,In_361,In_117);
nor U635 (N_635,In_13,In_219);
xnor U636 (N_636,In_57,In_8);
nor U637 (N_637,In_269,In_106);
nor U638 (N_638,In_56,In_51);
or U639 (N_639,In_299,In_461);
nand U640 (N_640,In_292,In_15);
nand U641 (N_641,In_375,In_33);
xnor U642 (N_642,In_325,In_369);
and U643 (N_643,In_237,In_278);
and U644 (N_644,In_450,In_375);
or U645 (N_645,In_418,In_331);
or U646 (N_646,In_447,In_379);
or U647 (N_647,In_365,In_2);
nor U648 (N_648,In_209,In_169);
or U649 (N_649,In_436,In_211);
xnor U650 (N_650,In_155,In_398);
nor U651 (N_651,In_353,In_408);
and U652 (N_652,In_65,In_180);
nand U653 (N_653,In_409,In_76);
xnor U654 (N_654,In_419,In_322);
nand U655 (N_655,In_425,In_411);
nand U656 (N_656,In_344,In_398);
xnor U657 (N_657,In_52,In_479);
and U658 (N_658,In_137,In_458);
nand U659 (N_659,In_332,In_12);
or U660 (N_660,In_140,In_363);
and U661 (N_661,In_12,In_351);
nand U662 (N_662,In_138,In_72);
nor U663 (N_663,In_247,In_190);
xnor U664 (N_664,In_78,In_295);
or U665 (N_665,In_187,In_183);
xnor U666 (N_666,In_428,In_456);
xnor U667 (N_667,In_47,In_59);
nand U668 (N_668,In_426,In_334);
or U669 (N_669,In_236,In_329);
and U670 (N_670,In_379,In_389);
nand U671 (N_671,In_400,In_187);
and U672 (N_672,In_154,In_351);
nor U673 (N_673,In_313,In_79);
nor U674 (N_674,In_498,In_327);
or U675 (N_675,In_43,In_486);
and U676 (N_676,In_370,In_80);
nor U677 (N_677,In_185,In_237);
or U678 (N_678,In_216,In_434);
nor U679 (N_679,In_196,In_167);
and U680 (N_680,In_34,In_128);
or U681 (N_681,In_447,In_134);
nor U682 (N_682,In_89,In_64);
and U683 (N_683,In_366,In_51);
xnor U684 (N_684,In_366,In_193);
nand U685 (N_685,In_404,In_337);
nand U686 (N_686,In_488,In_305);
nor U687 (N_687,In_35,In_308);
xnor U688 (N_688,In_62,In_131);
and U689 (N_689,In_187,In_442);
nand U690 (N_690,In_190,In_89);
and U691 (N_691,In_86,In_370);
or U692 (N_692,In_212,In_167);
xnor U693 (N_693,In_261,In_350);
nand U694 (N_694,In_170,In_445);
xor U695 (N_695,In_432,In_29);
xnor U696 (N_696,In_144,In_243);
nand U697 (N_697,In_284,In_356);
and U698 (N_698,In_244,In_72);
nor U699 (N_699,In_346,In_211);
xnor U700 (N_700,In_388,In_328);
and U701 (N_701,In_207,In_92);
and U702 (N_702,In_69,In_408);
nor U703 (N_703,In_165,In_260);
and U704 (N_704,In_400,In_305);
or U705 (N_705,In_115,In_148);
and U706 (N_706,In_263,In_297);
nand U707 (N_707,In_465,In_369);
and U708 (N_708,In_197,In_327);
and U709 (N_709,In_437,In_199);
xnor U710 (N_710,In_183,In_385);
nand U711 (N_711,In_476,In_205);
nand U712 (N_712,In_205,In_202);
and U713 (N_713,In_454,In_298);
nand U714 (N_714,In_139,In_340);
nand U715 (N_715,In_477,In_173);
xor U716 (N_716,In_426,In_162);
xor U717 (N_717,In_334,In_72);
nor U718 (N_718,In_142,In_239);
and U719 (N_719,In_236,In_204);
nor U720 (N_720,In_320,In_417);
or U721 (N_721,In_414,In_342);
xnor U722 (N_722,In_302,In_121);
xor U723 (N_723,In_282,In_25);
nand U724 (N_724,In_499,In_267);
nand U725 (N_725,In_171,In_275);
xor U726 (N_726,In_476,In_93);
and U727 (N_727,In_352,In_461);
nor U728 (N_728,In_228,In_211);
or U729 (N_729,In_486,In_168);
and U730 (N_730,In_101,In_48);
or U731 (N_731,In_283,In_324);
xnor U732 (N_732,In_319,In_135);
nor U733 (N_733,In_428,In_279);
nand U734 (N_734,In_396,In_132);
nand U735 (N_735,In_300,In_253);
xnor U736 (N_736,In_140,In_149);
or U737 (N_737,In_271,In_145);
nand U738 (N_738,In_307,In_411);
or U739 (N_739,In_262,In_283);
and U740 (N_740,In_331,In_221);
xnor U741 (N_741,In_185,In_426);
nor U742 (N_742,In_150,In_381);
xnor U743 (N_743,In_380,In_276);
nor U744 (N_744,In_398,In_234);
nor U745 (N_745,In_420,In_194);
nand U746 (N_746,In_202,In_306);
nor U747 (N_747,In_295,In_281);
nor U748 (N_748,In_135,In_494);
and U749 (N_749,In_122,In_342);
and U750 (N_750,N_665,N_472);
and U751 (N_751,N_163,N_549);
nand U752 (N_752,N_183,N_365);
and U753 (N_753,N_193,N_146);
and U754 (N_754,N_309,N_172);
nand U755 (N_755,N_112,N_496);
and U756 (N_756,N_134,N_581);
and U757 (N_757,N_250,N_529);
and U758 (N_758,N_741,N_44);
nor U759 (N_759,N_318,N_248);
xnor U760 (N_760,N_370,N_206);
xnor U761 (N_761,N_368,N_634);
and U762 (N_762,N_594,N_585);
nand U763 (N_763,N_60,N_438);
xnor U764 (N_764,N_568,N_666);
or U765 (N_765,N_316,N_562);
nand U766 (N_766,N_537,N_314);
nor U767 (N_767,N_119,N_552);
and U768 (N_768,N_45,N_371);
nand U769 (N_769,N_258,N_38);
or U770 (N_770,N_343,N_694);
nor U771 (N_771,N_720,N_280);
or U772 (N_772,N_490,N_432);
nand U773 (N_773,N_593,N_136);
nor U774 (N_774,N_405,N_703);
or U775 (N_775,N_685,N_51);
nor U776 (N_776,N_200,N_20);
nand U777 (N_777,N_606,N_94);
and U778 (N_778,N_174,N_623);
xnor U779 (N_779,N_11,N_246);
and U780 (N_780,N_379,N_538);
and U781 (N_781,N_313,N_483);
xor U782 (N_782,N_58,N_546);
and U783 (N_783,N_710,N_672);
nor U784 (N_784,N_281,N_444);
xor U785 (N_785,N_213,N_503);
xnor U786 (N_786,N_353,N_168);
xor U787 (N_787,N_460,N_505);
nand U788 (N_788,N_180,N_488);
xor U789 (N_789,N_56,N_140);
xor U790 (N_790,N_400,N_252);
and U791 (N_791,N_143,N_609);
nor U792 (N_792,N_473,N_127);
and U793 (N_793,N_514,N_648);
xor U794 (N_794,N_734,N_73);
nor U795 (N_795,N_475,N_737);
or U796 (N_796,N_504,N_743);
or U797 (N_797,N_435,N_676);
nand U798 (N_798,N_169,N_285);
or U799 (N_799,N_6,N_21);
or U800 (N_800,N_103,N_108);
nor U801 (N_801,N_532,N_417);
and U802 (N_802,N_42,N_71);
or U803 (N_803,N_566,N_544);
or U804 (N_804,N_380,N_458);
nor U805 (N_805,N_339,N_523);
nand U806 (N_806,N_461,N_224);
or U807 (N_807,N_231,N_525);
nand U808 (N_808,N_567,N_306);
and U809 (N_809,N_357,N_730);
and U810 (N_810,N_154,N_557);
nor U811 (N_811,N_684,N_257);
or U812 (N_812,N_31,N_499);
nor U813 (N_813,N_77,N_713);
xnor U814 (N_814,N_479,N_465);
nor U815 (N_815,N_655,N_5);
and U816 (N_816,N_745,N_81);
or U817 (N_817,N_447,N_282);
nand U818 (N_818,N_57,N_419);
xnor U819 (N_819,N_642,N_327);
and U820 (N_820,N_412,N_205);
xnor U821 (N_821,N_251,N_645);
or U822 (N_822,N_320,N_506);
nand U823 (N_823,N_203,N_521);
and U824 (N_824,N_291,N_346);
xnor U825 (N_825,N_748,N_111);
and U826 (N_826,N_364,N_36);
or U827 (N_827,N_548,N_559);
nor U828 (N_828,N_9,N_293);
and U829 (N_829,N_484,N_86);
and U830 (N_830,N_120,N_126);
and U831 (N_831,N_109,N_363);
and U832 (N_832,N_321,N_675);
nor U833 (N_833,N_133,N_325);
or U834 (N_834,N_330,N_345);
nand U835 (N_835,N_302,N_234);
or U836 (N_836,N_115,N_312);
and U837 (N_837,N_425,N_512);
nor U838 (N_838,N_278,N_605);
or U839 (N_839,N_614,N_697);
and U840 (N_840,N_22,N_65);
nor U841 (N_841,N_630,N_137);
nand U842 (N_842,N_607,N_121);
or U843 (N_843,N_715,N_315);
nand U844 (N_844,N_68,N_263);
and U845 (N_845,N_449,N_49);
or U846 (N_846,N_553,N_156);
and U847 (N_847,N_101,N_84);
xor U848 (N_848,N_667,N_261);
or U849 (N_849,N_30,N_153);
xor U850 (N_850,N_377,N_705);
nand U851 (N_851,N_192,N_236);
nor U852 (N_852,N_210,N_196);
nand U853 (N_853,N_443,N_732);
and U854 (N_854,N_673,N_360);
and U855 (N_855,N_212,N_125);
or U856 (N_856,N_721,N_481);
nand U857 (N_857,N_67,N_608);
and U858 (N_858,N_445,N_437);
or U859 (N_859,N_116,N_396);
and U860 (N_860,N_588,N_641);
nand U861 (N_861,N_452,N_480);
or U862 (N_862,N_90,N_34);
xnor U863 (N_863,N_340,N_170);
nor U864 (N_864,N_467,N_502);
or U865 (N_865,N_24,N_424);
nand U866 (N_866,N_324,N_696);
and U867 (N_867,N_262,N_157);
or U868 (N_868,N_601,N_47);
or U869 (N_869,N_564,N_178);
nand U870 (N_870,N_249,N_563);
nand U871 (N_871,N_188,N_66);
or U872 (N_872,N_15,N_344);
or U873 (N_873,N_332,N_747);
or U874 (N_874,N_139,N_241);
xor U875 (N_875,N_573,N_375);
or U876 (N_876,N_430,N_79);
nand U877 (N_877,N_464,N_387);
and U878 (N_878,N_207,N_88);
xnor U879 (N_879,N_495,N_16);
or U880 (N_880,N_201,N_602);
nor U881 (N_881,N_590,N_215);
xor U882 (N_882,N_184,N_310);
xnor U883 (N_883,N_268,N_305);
nor U884 (N_884,N_735,N_516);
nand U885 (N_885,N_358,N_238);
nor U886 (N_886,N_1,N_338);
nand U887 (N_887,N_329,N_220);
nand U888 (N_888,N_352,N_227);
nand U889 (N_889,N_547,N_422);
xor U890 (N_890,N_295,N_385);
nand U891 (N_891,N_415,N_738);
nand U892 (N_892,N_378,N_289);
and U893 (N_893,N_431,N_40);
or U894 (N_894,N_52,N_674);
nor U895 (N_895,N_511,N_359);
xor U896 (N_896,N_2,N_202);
or U897 (N_897,N_644,N_383);
and U898 (N_898,N_621,N_190);
nor U899 (N_899,N_414,N_12);
nor U900 (N_900,N_639,N_704);
xor U901 (N_901,N_519,N_392);
nand U902 (N_902,N_749,N_124);
xor U903 (N_903,N_105,N_668);
or U904 (N_904,N_98,N_144);
and U905 (N_905,N_501,N_149);
and U906 (N_906,N_23,N_613);
and U907 (N_907,N_554,N_135);
nand U908 (N_908,N_384,N_612);
xor U909 (N_909,N_189,N_221);
and U910 (N_910,N_17,N_647);
xor U911 (N_911,N_104,N_270);
nor U912 (N_912,N_80,N_398);
or U913 (N_913,N_381,N_93);
nor U914 (N_914,N_530,N_349);
or U915 (N_915,N_633,N_274);
nand U916 (N_916,N_436,N_264);
nor U917 (N_917,N_138,N_287);
and U918 (N_918,N_265,N_151);
xnor U919 (N_919,N_520,N_651);
xnor U920 (N_920,N_493,N_322);
nand U921 (N_921,N_652,N_256);
nor U922 (N_922,N_600,N_545);
nand U923 (N_923,N_725,N_575);
nor U924 (N_924,N_117,N_500);
and U925 (N_925,N_14,N_217);
nand U926 (N_926,N_240,N_509);
nand U927 (N_927,N_173,N_448);
xnor U928 (N_928,N_555,N_524);
and U929 (N_929,N_197,N_631);
xnor U930 (N_930,N_147,N_617);
xnor U931 (N_931,N_198,N_239);
xor U932 (N_932,N_334,N_54);
or U933 (N_933,N_476,N_474);
nor U934 (N_934,N_686,N_536);
nand U935 (N_935,N_401,N_578);
xor U936 (N_936,N_700,N_211);
nor U937 (N_937,N_660,N_37);
xnor U938 (N_938,N_102,N_551);
xor U939 (N_939,N_319,N_307);
nor U940 (N_940,N_328,N_724);
xor U941 (N_941,N_335,N_507);
nor U942 (N_942,N_470,N_457);
nand U943 (N_943,N_418,N_742);
nor U944 (N_944,N_204,N_373);
nand U945 (N_945,N_254,N_403);
nand U946 (N_946,N_455,N_97);
and U947 (N_947,N_550,N_679);
nor U948 (N_948,N_191,N_326);
nor U949 (N_949,N_699,N_277);
xnor U950 (N_950,N_497,N_736);
and U951 (N_951,N_229,N_517);
and U952 (N_952,N_454,N_311);
and U953 (N_953,N_331,N_463);
nand U954 (N_954,N_283,N_267);
and U955 (N_955,N_466,N_43);
and U956 (N_956,N_59,N_450);
xnor U957 (N_957,N_150,N_531);
nor U958 (N_958,N_235,N_708);
and U959 (N_959,N_656,N_245);
xor U960 (N_960,N_462,N_572);
xor U961 (N_961,N_19,N_626);
and U962 (N_962,N_485,N_355);
nor U963 (N_963,N_471,N_255);
xor U964 (N_964,N_680,N_8);
xor U965 (N_965,N_688,N_629);
nor U966 (N_966,N_587,N_657);
nor U967 (N_967,N_266,N_690);
nor U968 (N_968,N_649,N_214);
and U969 (N_969,N_286,N_627);
or U970 (N_970,N_440,N_638);
nor U971 (N_971,N_62,N_195);
nor U972 (N_972,N_176,N_25);
nor U973 (N_973,N_386,N_692);
nand U974 (N_974,N_388,N_162);
nor U975 (N_975,N_498,N_661);
and U976 (N_976,N_625,N_701);
or U977 (N_977,N_671,N_740);
xor U978 (N_978,N_0,N_230);
xor U979 (N_979,N_323,N_716);
nand U980 (N_980,N_618,N_522);
xnor U981 (N_981,N_635,N_271);
xor U982 (N_982,N_64,N_603);
nand U983 (N_983,N_32,N_539);
and U984 (N_984,N_29,N_534);
or U985 (N_985,N_372,N_711);
and U986 (N_986,N_413,N_518);
xor U987 (N_987,N_244,N_159);
nand U988 (N_988,N_7,N_693);
xor U989 (N_989,N_269,N_468);
or U990 (N_990,N_604,N_46);
and U991 (N_991,N_82,N_728);
or U992 (N_992,N_114,N_243);
nand U993 (N_993,N_279,N_175);
nand U994 (N_994,N_561,N_397);
xnor U995 (N_995,N_194,N_222);
or U996 (N_996,N_446,N_399);
nor U997 (N_997,N_533,N_160);
or U998 (N_998,N_219,N_208);
nor U999 (N_999,N_275,N_515);
or U1000 (N_1000,N_719,N_589);
xnor U1001 (N_1001,N_181,N_376);
nor U1002 (N_1002,N_273,N_167);
nor U1003 (N_1003,N_717,N_408);
xnor U1004 (N_1004,N_658,N_714);
or U1005 (N_1005,N_106,N_420);
nand U1006 (N_1006,N_145,N_259);
xor U1007 (N_1007,N_27,N_663);
and U1008 (N_1008,N_75,N_570);
xor U1009 (N_1009,N_723,N_610);
and U1010 (N_1010,N_620,N_712);
nand U1011 (N_1011,N_491,N_574);
xor U1012 (N_1012,N_225,N_599);
nand U1013 (N_1013,N_689,N_682);
nor U1014 (N_1014,N_739,N_237);
nand U1015 (N_1015,N_233,N_50);
nand U1016 (N_1016,N_39,N_441);
nand U1017 (N_1017,N_10,N_317);
nor U1018 (N_1018,N_336,N_28);
nand U1019 (N_1019,N_583,N_702);
or U1020 (N_1020,N_337,N_669);
nand U1021 (N_1021,N_678,N_95);
xnor U1022 (N_1022,N_406,N_643);
nor U1023 (N_1023,N_107,N_410);
and U1024 (N_1024,N_69,N_70);
and U1025 (N_1025,N_299,N_100);
and U1026 (N_1026,N_456,N_622);
xnor U1027 (N_1027,N_292,N_87);
xor U1028 (N_1028,N_152,N_584);
nand U1029 (N_1029,N_628,N_63);
nor U1030 (N_1030,N_571,N_284);
nand U1031 (N_1031,N_421,N_513);
or U1032 (N_1032,N_131,N_367);
and U1033 (N_1033,N_288,N_654);
or U1034 (N_1034,N_394,N_55);
or U1035 (N_1035,N_722,N_541);
xnor U1036 (N_1036,N_492,N_596);
nor U1037 (N_1037,N_158,N_580);
xnor U1038 (N_1038,N_186,N_26);
and U1039 (N_1039,N_347,N_303);
nand U1040 (N_1040,N_402,N_391);
or U1041 (N_1041,N_253,N_487);
or U1042 (N_1042,N_89,N_565);
nor U1043 (N_1043,N_369,N_129);
nand U1044 (N_1044,N_232,N_92);
and U1045 (N_1045,N_577,N_659);
and U1046 (N_1046,N_74,N_560);
xor U1047 (N_1047,N_304,N_171);
and U1048 (N_1048,N_218,N_395);
nor U1049 (N_1049,N_640,N_187);
and U1050 (N_1050,N_427,N_698);
and U1051 (N_1051,N_113,N_664);
or U1052 (N_1052,N_416,N_290);
nand U1053 (N_1053,N_374,N_662);
or U1054 (N_1054,N_61,N_744);
xor U1055 (N_1055,N_18,N_4);
and U1056 (N_1056,N_366,N_351);
or U1057 (N_1057,N_733,N_110);
xor U1058 (N_1058,N_382,N_122);
nor U1059 (N_1059,N_508,N_362);
xnor U1060 (N_1060,N_434,N_482);
or U1061 (N_1061,N_569,N_439);
nor U1062 (N_1062,N_165,N_540);
and U1063 (N_1063,N_615,N_228);
or U1064 (N_1064,N_216,N_528);
or U1065 (N_1065,N_718,N_478);
nand U1066 (N_1066,N_428,N_132);
nor U1067 (N_1067,N_469,N_650);
and U1068 (N_1068,N_709,N_526);
xnor U1069 (N_1069,N_543,N_260);
and U1070 (N_1070,N_3,N_726);
xor U1071 (N_1071,N_33,N_85);
or U1072 (N_1072,N_247,N_161);
nor U1073 (N_1073,N_677,N_276);
or U1074 (N_1074,N_209,N_598);
and U1075 (N_1075,N_272,N_558);
xor U1076 (N_1076,N_308,N_142);
and U1077 (N_1077,N_459,N_342);
nor U1078 (N_1078,N_595,N_99);
xor U1079 (N_1079,N_582,N_148);
nand U1080 (N_1080,N_48,N_477);
xor U1081 (N_1081,N_242,N_494);
xnor U1082 (N_1082,N_389,N_729);
nor U1083 (N_1083,N_489,N_354);
xnor U1084 (N_1084,N_350,N_96);
xnor U1085 (N_1085,N_141,N_576);
nor U1086 (N_1086,N_393,N_527);
and U1087 (N_1087,N_155,N_35);
or U1088 (N_1088,N_199,N_636);
nand U1089 (N_1089,N_185,N_619);
nor U1090 (N_1090,N_423,N_226);
or U1091 (N_1091,N_687,N_300);
and U1092 (N_1092,N_53,N_653);
xnor U1093 (N_1093,N_510,N_691);
xor U1094 (N_1094,N_632,N_333);
xnor U1095 (N_1095,N_646,N_182);
nor U1096 (N_1096,N_13,N_341);
and U1097 (N_1097,N_616,N_223);
nor U1098 (N_1098,N_586,N_404);
nor U1099 (N_1099,N_177,N_611);
and U1100 (N_1100,N_297,N_356);
or U1101 (N_1101,N_429,N_411);
or U1102 (N_1102,N_637,N_592);
and U1103 (N_1103,N_486,N_597);
xnor U1104 (N_1104,N_542,N_731);
or U1105 (N_1105,N_451,N_118);
xor U1106 (N_1106,N_556,N_409);
and U1107 (N_1107,N_301,N_76);
nor U1108 (N_1108,N_130,N_361);
nand U1109 (N_1109,N_166,N_683);
xor U1110 (N_1110,N_348,N_579);
nor U1111 (N_1111,N_298,N_681);
and U1112 (N_1112,N_179,N_296);
or U1113 (N_1113,N_707,N_695);
and U1114 (N_1114,N_41,N_591);
nand U1115 (N_1115,N_294,N_433);
xnor U1116 (N_1116,N_91,N_78);
nand U1117 (N_1117,N_128,N_706);
or U1118 (N_1118,N_390,N_727);
and U1119 (N_1119,N_123,N_442);
and U1120 (N_1120,N_426,N_670);
nand U1121 (N_1121,N_407,N_453);
and U1122 (N_1122,N_72,N_164);
and U1123 (N_1123,N_624,N_535);
nand U1124 (N_1124,N_746,N_83);
xnor U1125 (N_1125,N_631,N_604);
and U1126 (N_1126,N_294,N_503);
nand U1127 (N_1127,N_688,N_656);
or U1128 (N_1128,N_706,N_188);
and U1129 (N_1129,N_135,N_65);
nor U1130 (N_1130,N_745,N_443);
nor U1131 (N_1131,N_645,N_537);
xnor U1132 (N_1132,N_140,N_497);
nand U1133 (N_1133,N_467,N_478);
or U1134 (N_1134,N_547,N_288);
nand U1135 (N_1135,N_147,N_384);
xor U1136 (N_1136,N_390,N_393);
or U1137 (N_1137,N_600,N_447);
nand U1138 (N_1138,N_101,N_134);
or U1139 (N_1139,N_660,N_202);
nand U1140 (N_1140,N_179,N_636);
and U1141 (N_1141,N_420,N_311);
or U1142 (N_1142,N_663,N_318);
nor U1143 (N_1143,N_218,N_417);
or U1144 (N_1144,N_700,N_646);
xor U1145 (N_1145,N_729,N_439);
and U1146 (N_1146,N_473,N_164);
xnor U1147 (N_1147,N_154,N_680);
xor U1148 (N_1148,N_490,N_713);
and U1149 (N_1149,N_358,N_422);
nand U1150 (N_1150,N_105,N_249);
nor U1151 (N_1151,N_88,N_281);
and U1152 (N_1152,N_439,N_508);
and U1153 (N_1153,N_572,N_42);
nand U1154 (N_1154,N_9,N_166);
or U1155 (N_1155,N_118,N_73);
or U1156 (N_1156,N_69,N_536);
nand U1157 (N_1157,N_73,N_665);
xnor U1158 (N_1158,N_121,N_167);
or U1159 (N_1159,N_566,N_95);
and U1160 (N_1160,N_660,N_170);
nor U1161 (N_1161,N_509,N_335);
nor U1162 (N_1162,N_681,N_667);
and U1163 (N_1163,N_617,N_218);
nand U1164 (N_1164,N_723,N_675);
xnor U1165 (N_1165,N_376,N_145);
nand U1166 (N_1166,N_504,N_388);
nand U1167 (N_1167,N_447,N_320);
and U1168 (N_1168,N_385,N_234);
xnor U1169 (N_1169,N_502,N_83);
nor U1170 (N_1170,N_712,N_263);
nor U1171 (N_1171,N_570,N_350);
or U1172 (N_1172,N_26,N_553);
and U1173 (N_1173,N_339,N_410);
and U1174 (N_1174,N_518,N_735);
and U1175 (N_1175,N_492,N_424);
nand U1176 (N_1176,N_409,N_115);
nor U1177 (N_1177,N_476,N_322);
or U1178 (N_1178,N_361,N_737);
or U1179 (N_1179,N_309,N_465);
xor U1180 (N_1180,N_28,N_215);
nor U1181 (N_1181,N_190,N_25);
xnor U1182 (N_1182,N_710,N_321);
xnor U1183 (N_1183,N_64,N_634);
and U1184 (N_1184,N_91,N_668);
or U1185 (N_1185,N_162,N_511);
nor U1186 (N_1186,N_6,N_152);
nor U1187 (N_1187,N_583,N_438);
nand U1188 (N_1188,N_21,N_317);
or U1189 (N_1189,N_53,N_720);
nor U1190 (N_1190,N_307,N_368);
or U1191 (N_1191,N_123,N_398);
nor U1192 (N_1192,N_115,N_579);
xor U1193 (N_1193,N_254,N_115);
or U1194 (N_1194,N_377,N_329);
or U1195 (N_1195,N_458,N_27);
nand U1196 (N_1196,N_320,N_691);
xor U1197 (N_1197,N_728,N_671);
nor U1198 (N_1198,N_412,N_443);
or U1199 (N_1199,N_37,N_420);
or U1200 (N_1200,N_146,N_636);
nand U1201 (N_1201,N_185,N_600);
nand U1202 (N_1202,N_335,N_84);
and U1203 (N_1203,N_360,N_399);
nor U1204 (N_1204,N_350,N_600);
nor U1205 (N_1205,N_628,N_259);
nor U1206 (N_1206,N_122,N_25);
and U1207 (N_1207,N_426,N_326);
and U1208 (N_1208,N_154,N_152);
or U1209 (N_1209,N_431,N_715);
nor U1210 (N_1210,N_106,N_42);
nor U1211 (N_1211,N_640,N_685);
nor U1212 (N_1212,N_748,N_607);
xor U1213 (N_1213,N_229,N_349);
xnor U1214 (N_1214,N_0,N_236);
and U1215 (N_1215,N_749,N_633);
and U1216 (N_1216,N_29,N_264);
xor U1217 (N_1217,N_340,N_690);
nand U1218 (N_1218,N_722,N_323);
nand U1219 (N_1219,N_352,N_525);
or U1220 (N_1220,N_481,N_189);
xnor U1221 (N_1221,N_163,N_605);
or U1222 (N_1222,N_396,N_689);
or U1223 (N_1223,N_464,N_233);
nor U1224 (N_1224,N_29,N_687);
nand U1225 (N_1225,N_206,N_76);
and U1226 (N_1226,N_250,N_504);
nor U1227 (N_1227,N_321,N_347);
and U1228 (N_1228,N_514,N_191);
nor U1229 (N_1229,N_530,N_124);
nor U1230 (N_1230,N_438,N_154);
or U1231 (N_1231,N_669,N_54);
nand U1232 (N_1232,N_741,N_393);
or U1233 (N_1233,N_129,N_535);
xor U1234 (N_1234,N_14,N_302);
and U1235 (N_1235,N_659,N_622);
or U1236 (N_1236,N_251,N_266);
and U1237 (N_1237,N_639,N_50);
nor U1238 (N_1238,N_145,N_222);
nor U1239 (N_1239,N_612,N_665);
nor U1240 (N_1240,N_527,N_384);
and U1241 (N_1241,N_372,N_487);
and U1242 (N_1242,N_231,N_538);
xnor U1243 (N_1243,N_565,N_305);
xor U1244 (N_1244,N_465,N_704);
xor U1245 (N_1245,N_37,N_263);
nand U1246 (N_1246,N_528,N_157);
and U1247 (N_1247,N_514,N_138);
xnor U1248 (N_1248,N_361,N_693);
and U1249 (N_1249,N_636,N_598);
nor U1250 (N_1250,N_301,N_536);
xnor U1251 (N_1251,N_745,N_701);
xor U1252 (N_1252,N_112,N_250);
or U1253 (N_1253,N_478,N_440);
and U1254 (N_1254,N_727,N_453);
xor U1255 (N_1255,N_541,N_484);
xnor U1256 (N_1256,N_627,N_410);
or U1257 (N_1257,N_139,N_290);
nor U1258 (N_1258,N_613,N_8);
xor U1259 (N_1259,N_255,N_104);
xor U1260 (N_1260,N_257,N_310);
and U1261 (N_1261,N_86,N_356);
or U1262 (N_1262,N_64,N_487);
and U1263 (N_1263,N_199,N_608);
nor U1264 (N_1264,N_277,N_133);
nand U1265 (N_1265,N_596,N_591);
nor U1266 (N_1266,N_8,N_0);
or U1267 (N_1267,N_489,N_180);
nand U1268 (N_1268,N_83,N_3);
xnor U1269 (N_1269,N_233,N_363);
and U1270 (N_1270,N_292,N_29);
nor U1271 (N_1271,N_9,N_673);
nand U1272 (N_1272,N_607,N_485);
xnor U1273 (N_1273,N_485,N_134);
nor U1274 (N_1274,N_180,N_609);
or U1275 (N_1275,N_549,N_339);
nor U1276 (N_1276,N_205,N_663);
nor U1277 (N_1277,N_327,N_602);
nor U1278 (N_1278,N_214,N_585);
xnor U1279 (N_1279,N_686,N_390);
nor U1280 (N_1280,N_205,N_294);
xor U1281 (N_1281,N_32,N_344);
nor U1282 (N_1282,N_200,N_749);
and U1283 (N_1283,N_691,N_116);
xor U1284 (N_1284,N_449,N_342);
and U1285 (N_1285,N_55,N_657);
nor U1286 (N_1286,N_399,N_341);
and U1287 (N_1287,N_412,N_234);
or U1288 (N_1288,N_411,N_616);
and U1289 (N_1289,N_721,N_606);
or U1290 (N_1290,N_26,N_717);
nor U1291 (N_1291,N_664,N_443);
nand U1292 (N_1292,N_141,N_359);
xor U1293 (N_1293,N_567,N_376);
or U1294 (N_1294,N_710,N_448);
nand U1295 (N_1295,N_140,N_1);
or U1296 (N_1296,N_348,N_312);
nand U1297 (N_1297,N_593,N_34);
and U1298 (N_1298,N_177,N_219);
xnor U1299 (N_1299,N_220,N_695);
nor U1300 (N_1300,N_592,N_621);
or U1301 (N_1301,N_533,N_738);
nand U1302 (N_1302,N_24,N_468);
nor U1303 (N_1303,N_220,N_655);
nand U1304 (N_1304,N_39,N_166);
xnor U1305 (N_1305,N_288,N_404);
xor U1306 (N_1306,N_742,N_194);
or U1307 (N_1307,N_211,N_408);
nand U1308 (N_1308,N_239,N_405);
and U1309 (N_1309,N_692,N_430);
xor U1310 (N_1310,N_614,N_341);
and U1311 (N_1311,N_690,N_673);
or U1312 (N_1312,N_284,N_698);
nor U1313 (N_1313,N_595,N_231);
nor U1314 (N_1314,N_586,N_65);
nor U1315 (N_1315,N_95,N_354);
xnor U1316 (N_1316,N_542,N_67);
nor U1317 (N_1317,N_273,N_338);
xor U1318 (N_1318,N_32,N_621);
and U1319 (N_1319,N_118,N_156);
nand U1320 (N_1320,N_545,N_294);
nand U1321 (N_1321,N_73,N_574);
nand U1322 (N_1322,N_495,N_639);
xnor U1323 (N_1323,N_94,N_132);
nor U1324 (N_1324,N_281,N_503);
and U1325 (N_1325,N_274,N_394);
nand U1326 (N_1326,N_271,N_470);
xnor U1327 (N_1327,N_476,N_601);
or U1328 (N_1328,N_3,N_502);
nor U1329 (N_1329,N_653,N_10);
xor U1330 (N_1330,N_410,N_289);
and U1331 (N_1331,N_692,N_476);
nor U1332 (N_1332,N_369,N_501);
nand U1333 (N_1333,N_303,N_665);
nor U1334 (N_1334,N_274,N_382);
nor U1335 (N_1335,N_154,N_6);
nor U1336 (N_1336,N_54,N_682);
nor U1337 (N_1337,N_587,N_542);
xor U1338 (N_1338,N_665,N_337);
and U1339 (N_1339,N_411,N_634);
nor U1340 (N_1340,N_289,N_443);
nor U1341 (N_1341,N_485,N_455);
or U1342 (N_1342,N_180,N_550);
nor U1343 (N_1343,N_128,N_458);
xnor U1344 (N_1344,N_659,N_713);
nand U1345 (N_1345,N_447,N_109);
nor U1346 (N_1346,N_462,N_114);
nor U1347 (N_1347,N_591,N_411);
xnor U1348 (N_1348,N_737,N_519);
nor U1349 (N_1349,N_9,N_251);
nand U1350 (N_1350,N_721,N_442);
xor U1351 (N_1351,N_15,N_343);
nor U1352 (N_1352,N_492,N_233);
nand U1353 (N_1353,N_500,N_243);
or U1354 (N_1354,N_602,N_497);
xor U1355 (N_1355,N_66,N_685);
nor U1356 (N_1356,N_303,N_295);
nor U1357 (N_1357,N_581,N_347);
nor U1358 (N_1358,N_680,N_460);
and U1359 (N_1359,N_349,N_699);
nor U1360 (N_1360,N_248,N_16);
xnor U1361 (N_1361,N_147,N_544);
nor U1362 (N_1362,N_265,N_735);
nor U1363 (N_1363,N_504,N_132);
xnor U1364 (N_1364,N_301,N_540);
and U1365 (N_1365,N_422,N_741);
nor U1366 (N_1366,N_364,N_277);
nand U1367 (N_1367,N_129,N_542);
or U1368 (N_1368,N_680,N_524);
and U1369 (N_1369,N_392,N_543);
or U1370 (N_1370,N_282,N_183);
xnor U1371 (N_1371,N_376,N_355);
xnor U1372 (N_1372,N_696,N_170);
nor U1373 (N_1373,N_715,N_330);
and U1374 (N_1374,N_68,N_465);
and U1375 (N_1375,N_149,N_58);
nand U1376 (N_1376,N_397,N_595);
and U1377 (N_1377,N_296,N_131);
or U1378 (N_1378,N_143,N_352);
and U1379 (N_1379,N_479,N_188);
xnor U1380 (N_1380,N_660,N_658);
nand U1381 (N_1381,N_300,N_730);
and U1382 (N_1382,N_408,N_382);
nor U1383 (N_1383,N_637,N_572);
nor U1384 (N_1384,N_11,N_137);
xnor U1385 (N_1385,N_712,N_189);
or U1386 (N_1386,N_375,N_246);
nand U1387 (N_1387,N_738,N_559);
nand U1388 (N_1388,N_620,N_242);
nor U1389 (N_1389,N_519,N_564);
nor U1390 (N_1390,N_633,N_132);
and U1391 (N_1391,N_74,N_716);
and U1392 (N_1392,N_659,N_339);
nand U1393 (N_1393,N_50,N_14);
xor U1394 (N_1394,N_88,N_526);
nor U1395 (N_1395,N_124,N_535);
xor U1396 (N_1396,N_227,N_370);
nand U1397 (N_1397,N_618,N_396);
xor U1398 (N_1398,N_624,N_607);
and U1399 (N_1399,N_175,N_307);
nor U1400 (N_1400,N_351,N_308);
nand U1401 (N_1401,N_3,N_77);
nor U1402 (N_1402,N_36,N_399);
nor U1403 (N_1403,N_709,N_555);
and U1404 (N_1404,N_30,N_446);
and U1405 (N_1405,N_186,N_52);
xor U1406 (N_1406,N_64,N_678);
nor U1407 (N_1407,N_21,N_742);
nor U1408 (N_1408,N_122,N_185);
and U1409 (N_1409,N_95,N_293);
xor U1410 (N_1410,N_381,N_192);
xnor U1411 (N_1411,N_299,N_254);
nand U1412 (N_1412,N_1,N_389);
nor U1413 (N_1413,N_278,N_573);
nand U1414 (N_1414,N_697,N_218);
and U1415 (N_1415,N_316,N_18);
or U1416 (N_1416,N_557,N_41);
and U1417 (N_1417,N_315,N_419);
xor U1418 (N_1418,N_167,N_105);
xnor U1419 (N_1419,N_664,N_171);
xor U1420 (N_1420,N_165,N_159);
xnor U1421 (N_1421,N_540,N_150);
nand U1422 (N_1422,N_656,N_253);
or U1423 (N_1423,N_10,N_22);
nor U1424 (N_1424,N_56,N_623);
and U1425 (N_1425,N_377,N_599);
nand U1426 (N_1426,N_501,N_7);
nor U1427 (N_1427,N_347,N_509);
and U1428 (N_1428,N_577,N_158);
nor U1429 (N_1429,N_744,N_197);
nor U1430 (N_1430,N_338,N_720);
nand U1431 (N_1431,N_339,N_739);
nor U1432 (N_1432,N_129,N_228);
and U1433 (N_1433,N_626,N_110);
xnor U1434 (N_1434,N_117,N_163);
xor U1435 (N_1435,N_425,N_268);
xor U1436 (N_1436,N_416,N_455);
and U1437 (N_1437,N_456,N_385);
xnor U1438 (N_1438,N_435,N_678);
and U1439 (N_1439,N_664,N_136);
nor U1440 (N_1440,N_403,N_108);
nand U1441 (N_1441,N_45,N_534);
or U1442 (N_1442,N_58,N_634);
or U1443 (N_1443,N_99,N_385);
xnor U1444 (N_1444,N_451,N_182);
and U1445 (N_1445,N_126,N_235);
or U1446 (N_1446,N_532,N_560);
nor U1447 (N_1447,N_82,N_656);
xnor U1448 (N_1448,N_172,N_701);
nor U1449 (N_1449,N_157,N_12);
and U1450 (N_1450,N_317,N_113);
or U1451 (N_1451,N_468,N_747);
nor U1452 (N_1452,N_174,N_661);
and U1453 (N_1453,N_25,N_569);
and U1454 (N_1454,N_666,N_693);
nand U1455 (N_1455,N_404,N_740);
nand U1456 (N_1456,N_131,N_459);
and U1457 (N_1457,N_467,N_574);
or U1458 (N_1458,N_597,N_519);
xnor U1459 (N_1459,N_60,N_266);
or U1460 (N_1460,N_189,N_135);
nand U1461 (N_1461,N_439,N_600);
and U1462 (N_1462,N_3,N_649);
or U1463 (N_1463,N_413,N_29);
nor U1464 (N_1464,N_396,N_507);
xnor U1465 (N_1465,N_451,N_426);
xnor U1466 (N_1466,N_471,N_115);
or U1467 (N_1467,N_698,N_108);
nand U1468 (N_1468,N_34,N_546);
nand U1469 (N_1469,N_538,N_501);
nor U1470 (N_1470,N_695,N_185);
xnor U1471 (N_1471,N_345,N_290);
xnor U1472 (N_1472,N_126,N_222);
nor U1473 (N_1473,N_75,N_543);
nand U1474 (N_1474,N_203,N_470);
and U1475 (N_1475,N_442,N_404);
xnor U1476 (N_1476,N_442,N_61);
or U1477 (N_1477,N_666,N_504);
nand U1478 (N_1478,N_611,N_585);
or U1479 (N_1479,N_652,N_200);
or U1480 (N_1480,N_674,N_458);
or U1481 (N_1481,N_539,N_445);
nand U1482 (N_1482,N_701,N_668);
nor U1483 (N_1483,N_95,N_389);
and U1484 (N_1484,N_545,N_280);
xor U1485 (N_1485,N_215,N_672);
nor U1486 (N_1486,N_204,N_742);
nor U1487 (N_1487,N_369,N_238);
nand U1488 (N_1488,N_712,N_217);
or U1489 (N_1489,N_150,N_323);
or U1490 (N_1490,N_10,N_701);
nor U1491 (N_1491,N_71,N_462);
xnor U1492 (N_1492,N_57,N_427);
nor U1493 (N_1493,N_709,N_560);
and U1494 (N_1494,N_539,N_529);
or U1495 (N_1495,N_231,N_553);
and U1496 (N_1496,N_325,N_683);
or U1497 (N_1497,N_604,N_317);
nor U1498 (N_1498,N_113,N_264);
and U1499 (N_1499,N_53,N_404);
nand U1500 (N_1500,N_1338,N_873);
or U1501 (N_1501,N_895,N_1446);
nor U1502 (N_1502,N_1371,N_831);
xnor U1503 (N_1503,N_1306,N_1158);
and U1504 (N_1504,N_968,N_1349);
nor U1505 (N_1505,N_1055,N_1029);
nor U1506 (N_1506,N_1324,N_1017);
xnor U1507 (N_1507,N_893,N_1109);
or U1508 (N_1508,N_1107,N_931);
and U1509 (N_1509,N_942,N_1414);
xor U1510 (N_1510,N_1042,N_1229);
and U1511 (N_1511,N_861,N_1407);
and U1512 (N_1512,N_818,N_1309);
xnor U1513 (N_1513,N_1332,N_838);
and U1514 (N_1514,N_1365,N_1149);
nor U1515 (N_1515,N_1172,N_1215);
nor U1516 (N_1516,N_1007,N_1199);
xnor U1517 (N_1517,N_1067,N_1277);
nor U1518 (N_1518,N_975,N_1232);
or U1519 (N_1519,N_820,N_1267);
nor U1520 (N_1520,N_965,N_917);
nand U1521 (N_1521,N_1266,N_835);
and U1522 (N_1522,N_1219,N_1207);
and U1523 (N_1523,N_1111,N_933);
xor U1524 (N_1524,N_1481,N_1316);
nand U1525 (N_1525,N_1386,N_1060);
nand U1526 (N_1526,N_1099,N_1401);
or U1527 (N_1527,N_1133,N_1265);
or U1528 (N_1528,N_765,N_1186);
nor U1529 (N_1529,N_757,N_1453);
nand U1530 (N_1530,N_991,N_981);
or U1531 (N_1531,N_887,N_1305);
and U1532 (N_1532,N_1369,N_1169);
or U1533 (N_1533,N_1159,N_1122);
or U1534 (N_1534,N_868,N_1069);
and U1535 (N_1535,N_901,N_786);
xor U1536 (N_1536,N_1478,N_1283);
nor U1537 (N_1537,N_1014,N_1114);
nand U1538 (N_1538,N_852,N_1058);
nor U1539 (N_1539,N_879,N_1342);
or U1540 (N_1540,N_1239,N_1056);
or U1541 (N_1541,N_994,N_836);
nand U1542 (N_1542,N_1004,N_945);
nand U1543 (N_1543,N_1032,N_771);
or U1544 (N_1544,N_1320,N_1418);
nand U1545 (N_1545,N_1065,N_1070);
nand U1546 (N_1546,N_956,N_1209);
and U1547 (N_1547,N_793,N_1436);
xor U1548 (N_1548,N_1413,N_905);
xnor U1549 (N_1549,N_927,N_1043);
nand U1550 (N_1550,N_1328,N_819);
nor U1551 (N_1551,N_1129,N_1459);
and U1552 (N_1552,N_928,N_1078);
or U1553 (N_1553,N_1173,N_1441);
xor U1554 (N_1554,N_1221,N_1467);
and U1555 (N_1555,N_1088,N_809);
and U1556 (N_1556,N_1304,N_1112);
nor U1557 (N_1557,N_1497,N_1091);
nor U1558 (N_1558,N_1167,N_1053);
nor U1559 (N_1559,N_805,N_896);
xor U1560 (N_1560,N_1174,N_1351);
nand U1561 (N_1561,N_1260,N_1347);
xor U1562 (N_1562,N_1404,N_1483);
xor U1563 (N_1563,N_1355,N_824);
or U1564 (N_1564,N_932,N_1329);
or U1565 (N_1565,N_1137,N_1457);
nor U1566 (N_1566,N_1333,N_1061);
nor U1567 (N_1567,N_1302,N_1241);
nand U1568 (N_1568,N_1444,N_1432);
nand U1569 (N_1569,N_783,N_1144);
xor U1570 (N_1570,N_972,N_1339);
nand U1571 (N_1571,N_890,N_1242);
nor U1572 (N_1572,N_1045,N_1185);
nor U1573 (N_1573,N_792,N_814);
and U1574 (N_1574,N_912,N_1374);
xnor U1575 (N_1575,N_1227,N_1311);
xnor U1576 (N_1576,N_1202,N_1212);
xnor U1577 (N_1577,N_1276,N_1358);
xnor U1578 (N_1578,N_1104,N_878);
nor U1579 (N_1579,N_1254,N_1188);
nor U1580 (N_1580,N_758,N_1279);
nor U1581 (N_1581,N_1100,N_1068);
nor U1582 (N_1582,N_1161,N_1147);
xnor U1583 (N_1583,N_813,N_1142);
xor U1584 (N_1584,N_902,N_1354);
nand U1585 (N_1585,N_839,N_1390);
or U1586 (N_1586,N_955,N_1325);
nand U1587 (N_1587,N_1257,N_997);
nand U1588 (N_1588,N_894,N_1310);
nor U1589 (N_1589,N_1396,N_1127);
xnor U1590 (N_1590,N_1164,N_1005);
nand U1591 (N_1591,N_1288,N_1015);
nor U1592 (N_1592,N_1486,N_781);
and U1593 (N_1593,N_1204,N_1422);
nor U1594 (N_1594,N_1250,N_801);
xnor U1595 (N_1595,N_1222,N_907);
nor U1596 (N_1596,N_987,N_1256);
nor U1597 (N_1597,N_1334,N_1367);
and U1598 (N_1598,N_1116,N_1024);
nor U1599 (N_1599,N_1300,N_990);
xnor U1600 (N_1600,N_970,N_1203);
xnor U1601 (N_1601,N_1409,N_1124);
xor U1602 (N_1602,N_1195,N_1400);
nand U1603 (N_1603,N_791,N_840);
or U1604 (N_1604,N_941,N_1388);
nand U1605 (N_1605,N_1106,N_867);
nor U1606 (N_1606,N_1220,N_1489);
xor U1607 (N_1607,N_830,N_1020);
nor U1608 (N_1608,N_989,N_984);
or U1609 (N_1609,N_1314,N_1179);
xnor U1610 (N_1610,N_1170,N_1073);
xor U1611 (N_1611,N_1191,N_1050);
or U1612 (N_1612,N_983,N_1000);
nor U1613 (N_1613,N_949,N_1447);
or U1614 (N_1614,N_1148,N_954);
nand U1615 (N_1615,N_1139,N_935);
xnor U1616 (N_1616,N_1378,N_947);
nor U1617 (N_1617,N_1255,N_769);
xnor U1618 (N_1618,N_859,N_936);
nand U1619 (N_1619,N_1008,N_986);
xor U1620 (N_1620,N_1284,N_1468);
and U1621 (N_1621,N_1397,N_799);
nand U1622 (N_1622,N_1151,N_1079);
xnor U1623 (N_1623,N_1370,N_1214);
nand U1624 (N_1624,N_763,N_844);
xnor U1625 (N_1625,N_1016,N_1103);
xnor U1626 (N_1626,N_1415,N_1076);
nand U1627 (N_1627,N_1477,N_1417);
nand U1628 (N_1628,N_1443,N_1197);
or U1629 (N_1629,N_1132,N_1383);
xnor U1630 (N_1630,N_755,N_1101);
nand U1631 (N_1631,N_1348,N_1335);
xor U1632 (N_1632,N_770,N_1162);
or U1633 (N_1633,N_800,N_1271);
nor U1634 (N_1634,N_898,N_953);
nor U1635 (N_1635,N_1461,N_885);
xor U1636 (N_1636,N_909,N_1323);
or U1637 (N_1637,N_976,N_1321);
nand U1638 (N_1638,N_1428,N_1449);
or U1639 (N_1639,N_1228,N_871);
nor U1640 (N_1640,N_1084,N_1287);
or U1641 (N_1641,N_1140,N_1072);
and U1642 (N_1642,N_1393,N_1036);
nor U1643 (N_1643,N_863,N_969);
nor U1644 (N_1644,N_1463,N_1493);
and U1645 (N_1645,N_759,N_1094);
and U1646 (N_1646,N_1379,N_1048);
or U1647 (N_1647,N_1405,N_1187);
or U1648 (N_1648,N_1165,N_939);
and U1649 (N_1649,N_1431,N_1089);
xor U1650 (N_1650,N_1308,N_1160);
xnor U1651 (N_1651,N_1336,N_1495);
nor U1652 (N_1652,N_1006,N_866);
nor U1653 (N_1653,N_1264,N_850);
xnor U1654 (N_1654,N_847,N_1201);
and U1655 (N_1655,N_1190,N_916);
nor U1656 (N_1656,N_827,N_1157);
xor U1657 (N_1657,N_1085,N_921);
xnor U1658 (N_1658,N_1387,N_764);
nor U1659 (N_1659,N_1097,N_903);
nor U1660 (N_1660,N_767,N_1438);
or U1661 (N_1661,N_846,N_1297);
xnor U1662 (N_1662,N_1426,N_978);
or U1663 (N_1663,N_858,N_1131);
or U1664 (N_1664,N_1217,N_752);
nand U1665 (N_1665,N_948,N_1293);
nor U1666 (N_1666,N_1052,N_982);
nand U1667 (N_1667,N_1128,N_1208);
and U1668 (N_1668,N_1291,N_1350);
nand U1669 (N_1669,N_1421,N_998);
xor U1670 (N_1670,N_1166,N_1152);
xor U1671 (N_1671,N_964,N_1259);
or U1672 (N_1672,N_929,N_795);
nor U1673 (N_1673,N_1253,N_845);
nand U1674 (N_1674,N_973,N_1391);
nand U1675 (N_1675,N_807,N_779);
nand U1676 (N_1676,N_1275,N_922);
nor U1677 (N_1677,N_751,N_869);
xor U1678 (N_1678,N_784,N_1019);
nor U1679 (N_1679,N_1230,N_1030);
nand U1680 (N_1680,N_1315,N_906);
nor U1681 (N_1681,N_1134,N_1427);
and U1682 (N_1682,N_993,N_911);
or U1683 (N_1683,N_1218,N_1246);
nand U1684 (N_1684,N_967,N_1041);
or U1685 (N_1685,N_923,N_1281);
and U1686 (N_1686,N_1086,N_860);
and U1687 (N_1687,N_1343,N_1364);
or U1688 (N_1688,N_1237,N_750);
nand U1689 (N_1689,N_1098,N_1345);
and U1690 (N_1690,N_798,N_1492);
or U1691 (N_1691,N_856,N_1485);
nand U1692 (N_1692,N_1423,N_806);
nand U1693 (N_1693,N_1143,N_1194);
nand U1694 (N_1694,N_1245,N_1464);
or U1695 (N_1695,N_1233,N_963);
nor U1696 (N_1696,N_768,N_1487);
and U1697 (N_1697,N_1049,N_940);
nor U1698 (N_1698,N_1223,N_1382);
xor U1699 (N_1699,N_995,N_1327);
or U1700 (N_1700,N_958,N_1080);
xor U1701 (N_1701,N_1211,N_1482);
or U1702 (N_1702,N_1352,N_919);
nand U1703 (N_1703,N_812,N_1296);
xnor U1704 (N_1704,N_1150,N_1430);
nand U1705 (N_1705,N_1282,N_1154);
xnor U1706 (N_1706,N_920,N_1040);
or U1707 (N_1707,N_1225,N_1126);
nor U1708 (N_1708,N_1025,N_1480);
or U1709 (N_1709,N_1460,N_837);
nand U1710 (N_1710,N_1189,N_1398);
and U1711 (N_1711,N_1499,N_817);
nand U1712 (N_1712,N_971,N_1363);
nor U1713 (N_1713,N_864,N_899);
nor U1714 (N_1714,N_1322,N_1471);
xor U1715 (N_1715,N_849,N_1361);
nand U1716 (N_1716,N_1317,N_1385);
and U1717 (N_1717,N_774,N_1394);
or U1718 (N_1718,N_900,N_1263);
and U1719 (N_1719,N_1392,N_1135);
nand U1720 (N_1720,N_1096,N_1377);
nor U1721 (N_1721,N_1424,N_914);
nand U1722 (N_1722,N_1003,N_1023);
and U1723 (N_1723,N_1366,N_1163);
nand U1724 (N_1724,N_1047,N_1054);
nor U1725 (N_1725,N_1033,N_1251);
nor U1726 (N_1726,N_1285,N_1341);
xor U1727 (N_1727,N_1469,N_1071);
nand U1728 (N_1728,N_1018,N_1092);
xnor U1729 (N_1729,N_756,N_1198);
nor U1730 (N_1730,N_1380,N_1268);
nor U1731 (N_1731,N_874,N_1434);
or U1732 (N_1732,N_1235,N_1435);
nor U1733 (N_1733,N_1236,N_1344);
xnor U1734 (N_1734,N_1238,N_1326);
nand U1735 (N_1735,N_1368,N_1410);
or U1736 (N_1736,N_1295,N_1240);
and U1737 (N_1737,N_1445,N_1090);
nor U1738 (N_1738,N_999,N_862);
nor U1739 (N_1739,N_1110,N_1027);
xor U1740 (N_1740,N_1066,N_1115);
xnor U1741 (N_1741,N_754,N_943);
nand U1742 (N_1742,N_946,N_1184);
and U1743 (N_1743,N_773,N_1470);
nand U1744 (N_1744,N_1412,N_760);
nor U1745 (N_1745,N_1454,N_1113);
or U1746 (N_1746,N_1474,N_1416);
or U1747 (N_1747,N_889,N_886);
xnor U1748 (N_1748,N_832,N_1330);
nand U1749 (N_1749,N_1360,N_855);
nor U1750 (N_1750,N_790,N_753);
and U1751 (N_1751,N_1168,N_944);
nor U1752 (N_1752,N_957,N_1269);
nand U1753 (N_1753,N_1312,N_794);
nor U1754 (N_1754,N_1439,N_1231);
nor U1755 (N_1755,N_1138,N_962);
or U1756 (N_1756,N_1181,N_1034);
nand U1757 (N_1757,N_851,N_1337);
and U1758 (N_1758,N_1272,N_1491);
and U1759 (N_1759,N_1108,N_1062);
xor U1760 (N_1760,N_1498,N_816);
nor U1761 (N_1761,N_918,N_1301);
xnor U1762 (N_1762,N_1216,N_833);
xor U1763 (N_1763,N_1087,N_1026);
xor U1764 (N_1764,N_823,N_1121);
nor U1765 (N_1765,N_865,N_1118);
nand U1766 (N_1766,N_1299,N_1130);
or U1767 (N_1767,N_788,N_1175);
or U1768 (N_1768,N_1145,N_853);
nand U1769 (N_1769,N_848,N_1331);
or U1770 (N_1770,N_1433,N_804);
or U1771 (N_1771,N_891,N_1357);
xnor U1772 (N_1772,N_1009,N_1248);
nor U1773 (N_1773,N_880,N_934);
and U1774 (N_1774,N_766,N_1440);
and U1775 (N_1775,N_1346,N_937);
and U1776 (N_1776,N_826,N_780);
and U1777 (N_1777,N_1125,N_1252);
nor U1778 (N_1778,N_1156,N_1200);
nand U1779 (N_1779,N_1451,N_1462);
nor U1780 (N_1780,N_1153,N_1313);
nor U1781 (N_1781,N_882,N_1002);
nand U1782 (N_1782,N_884,N_1117);
nand U1783 (N_1783,N_821,N_857);
and U1784 (N_1784,N_1082,N_1213);
xor U1785 (N_1785,N_1473,N_1183);
and U1786 (N_1786,N_1455,N_782);
or U1787 (N_1787,N_1384,N_1408);
xnor U1788 (N_1788,N_1081,N_1146);
nor U1789 (N_1789,N_881,N_777);
and U1790 (N_1790,N_1075,N_1362);
nor U1791 (N_1791,N_1001,N_854);
xor U1792 (N_1792,N_1206,N_876);
or U1793 (N_1793,N_1083,N_1051);
nor U1794 (N_1794,N_1286,N_959);
xor U1795 (N_1795,N_1476,N_1171);
nand U1796 (N_1796,N_1466,N_1064);
and U1797 (N_1797,N_803,N_952);
nor U1798 (N_1798,N_1465,N_966);
or U1799 (N_1799,N_761,N_1307);
and U1800 (N_1800,N_1450,N_1381);
or U1801 (N_1801,N_1210,N_1294);
xnor U1802 (N_1802,N_796,N_1290);
and U1803 (N_1803,N_951,N_1249);
nor U1804 (N_1804,N_950,N_870);
and U1805 (N_1805,N_1429,N_842);
and U1806 (N_1806,N_1359,N_1488);
or U1807 (N_1807,N_1292,N_1105);
or U1808 (N_1808,N_789,N_1012);
nand U1809 (N_1809,N_875,N_961);
nor U1810 (N_1810,N_1031,N_1120);
nor U1811 (N_1811,N_1472,N_841);
xnor U1812 (N_1812,N_1261,N_1419);
and U1813 (N_1813,N_1475,N_1298);
xnor U1814 (N_1814,N_1376,N_1057);
or U1815 (N_1815,N_1077,N_1319);
and U1816 (N_1816,N_926,N_1234);
nand U1817 (N_1817,N_930,N_1403);
nor U1818 (N_1818,N_1028,N_810);
nor U1819 (N_1819,N_1278,N_1356);
xor U1820 (N_1820,N_1102,N_1420);
nand U1821 (N_1821,N_1496,N_1093);
or U1822 (N_1822,N_1013,N_988);
nor U1823 (N_1823,N_1375,N_808);
nand U1824 (N_1824,N_822,N_1373);
nor U1825 (N_1825,N_1141,N_1010);
or U1826 (N_1826,N_1479,N_892);
xor U1827 (N_1827,N_1452,N_778);
and U1828 (N_1828,N_1484,N_1258);
nor U1829 (N_1829,N_1046,N_785);
nor U1830 (N_1830,N_1243,N_980);
or U1831 (N_1831,N_1456,N_1244);
nand U1832 (N_1832,N_904,N_1289);
and U1833 (N_1833,N_925,N_1192);
xnor U1834 (N_1834,N_787,N_1011);
and U1835 (N_1835,N_883,N_762);
or U1836 (N_1836,N_992,N_1063);
nor U1837 (N_1837,N_1038,N_1193);
nand U1838 (N_1838,N_1411,N_1395);
and U1839 (N_1839,N_772,N_1205);
xnor U1840 (N_1840,N_1425,N_1178);
nor U1841 (N_1841,N_802,N_811);
xor U1842 (N_1842,N_979,N_815);
nor U1843 (N_1843,N_1402,N_915);
nand U1844 (N_1844,N_1494,N_1176);
xnor U1845 (N_1845,N_1442,N_1155);
nor U1846 (N_1846,N_1274,N_828);
nor U1847 (N_1847,N_775,N_1177);
nor U1848 (N_1848,N_877,N_913);
nand U1849 (N_1849,N_1372,N_1021);
nand U1850 (N_1850,N_996,N_1224);
or U1851 (N_1851,N_960,N_1037);
nor U1852 (N_1852,N_1273,N_924);
or U1853 (N_1853,N_1270,N_888);
xnor U1854 (N_1854,N_1318,N_825);
and U1855 (N_1855,N_1123,N_938);
xnor U1856 (N_1856,N_834,N_985);
xor U1857 (N_1857,N_1247,N_1119);
or U1858 (N_1858,N_1182,N_1022);
and U1859 (N_1859,N_1074,N_1262);
xor U1860 (N_1860,N_910,N_908);
xor U1861 (N_1861,N_1448,N_1389);
nor U1862 (N_1862,N_1039,N_1044);
nand U1863 (N_1863,N_1353,N_1399);
nand U1864 (N_1864,N_897,N_1303);
nor U1865 (N_1865,N_1035,N_977);
or U1866 (N_1866,N_1458,N_1406);
xor U1867 (N_1867,N_1059,N_1437);
nand U1868 (N_1868,N_1280,N_1095);
nor U1869 (N_1869,N_872,N_1340);
and U1870 (N_1870,N_843,N_974);
or U1871 (N_1871,N_797,N_1226);
xor U1872 (N_1872,N_1136,N_829);
or U1873 (N_1873,N_1490,N_1196);
xor U1874 (N_1874,N_776,N_1180);
or U1875 (N_1875,N_1229,N_979);
or U1876 (N_1876,N_1194,N_1476);
xnor U1877 (N_1877,N_1495,N_864);
nand U1878 (N_1878,N_935,N_996);
nand U1879 (N_1879,N_829,N_1389);
nand U1880 (N_1880,N_1413,N_1445);
or U1881 (N_1881,N_1026,N_1271);
or U1882 (N_1882,N_1440,N_1290);
or U1883 (N_1883,N_1303,N_976);
and U1884 (N_1884,N_1274,N_864);
nor U1885 (N_1885,N_1311,N_1055);
nand U1886 (N_1886,N_831,N_791);
nor U1887 (N_1887,N_774,N_1164);
xnor U1888 (N_1888,N_1427,N_785);
and U1889 (N_1889,N_1099,N_1117);
nand U1890 (N_1890,N_850,N_924);
nor U1891 (N_1891,N_815,N_991);
nor U1892 (N_1892,N_1457,N_908);
or U1893 (N_1893,N_1296,N_1341);
nor U1894 (N_1894,N_1216,N_1051);
nor U1895 (N_1895,N_788,N_1070);
nand U1896 (N_1896,N_1289,N_1205);
nor U1897 (N_1897,N_1231,N_1045);
xnor U1898 (N_1898,N_951,N_764);
nand U1899 (N_1899,N_1353,N_1147);
and U1900 (N_1900,N_878,N_1024);
nor U1901 (N_1901,N_951,N_1212);
nand U1902 (N_1902,N_770,N_857);
or U1903 (N_1903,N_1487,N_1150);
nor U1904 (N_1904,N_1151,N_933);
or U1905 (N_1905,N_913,N_1044);
nor U1906 (N_1906,N_808,N_1492);
xnor U1907 (N_1907,N_811,N_1164);
or U1908 (N_1908,N_847,N_1163);
and U1909 (N_1909,N_1385,N_1354);
nand U1910 (N_1910,N_758,N_1429);
nand U1911 (N_1911,N_1024,N_939);
xnor U1912 (N_1912,N_1070,N_1245);
nand U1913 (N_1913,N_1097,N_1079);
nor U1914 (N_1914,N_1151,N_1063);
nor U1915 (N_1915,N_1029,N_978);
and U1916 (N_1916,N_1380,N_1343);
or U1917 (N_1917,N_1107,N_966);
nor U1918 (N_1918,N_1073,N_1093);
nand U1919 (N_1919,N_1222,N_847);
xnor U1920 (N_1920,N_1425,N_1109);
nor U1921 (N_1921,N_1124,N_1153);
nand U1922 (N_1922,N_1400,N_1299);
xor U1923 (N_1923,N_1190,N_1479);
or U1924 (N_1924,N_867,N_1476);
nand U1925 (N_1925,N_1219,N_845);
or U1926 (N_1926,N_861,N_978);
xor U1927 (N_1927,N_913,N_1100);
nand U1928 (N_1928,N_1023,N_1138);
nand U1929 (N_1929,N_1497,N_796);
and U1930 (N_1930,N_922,N_1288);
xnor U1931 (N_1931,N_1111,N_1179);
and U1932 (N_1932,N_1269,N_1174);
nand U1933 (N_1933,N_1110,N_878);
or U1934 (N_1934,N_1444,N_847);
nor U1935 (N_1935,N_1476,N_1415);
nor U1936 (N_1936,N_1318,N_948);
nor U1937 (N_1937,N_1181,N_872);
nand U1938 (N_1938,N_886,N_1310);
or U1939 (N_1939,N_1345,N_1125);
nor U1940 (N_1940,N_1489,N_1102);
nor U1941 (N_1941,N_976,N_1270);
xor U1942 (N_1942,N_1344,N_1442);
nand U1943 (N_1943,N_1473,N_1455);
nand U1944 (N_1944,N_849,N_1119);
nor U1945 (N_1945,N_1476,N_1297);
nand U1946 (N_1946,N_1270,N_1440);
nor U1947 (N_1947,N_1385,N_1242);
nor U1948 (N_1948,N_798,N_881);
and U1949 (N_1949,N_808,N_1015);
nor U1950 (N_1950,N_1248,N_1163);
and U1951 (N_1951,N_1025,N_858);
or U1952 (N_1952,N_1099,N_1171);
and U1953 (N_1953,N_1190,N_955);
xor U1954 (N_1954,N_1407,N_1281);
xor U1955 (N_1955,N_1104,N_1459);
and U1956 (N_1956,N_1496,N_1187);
and U1957 (N_1957,N_1135,N_1090);
or U1958 (N_1958,N_909,N_966);
xnor U1959 (N_1959,N_1270,N_1351);
and U1960 (N_1960,N_947,N_1434);
or U1961 (N_1961,N_1409,N_1198);
and U1962 (N_1962,N_1337,N_783);
nor U1963 (N_1963,N_1485,N_819);
nand U1964 (N_1964,N_1466,N_1401);
or U1965 (N_1965,N_1325,N_985);
and U1966 (N_1966,N_1401,N_1179);
xor U1967 (N_1967,N_1281,N_752);
nand U1968 (N_1968,N_1147,N_962);
or U1969 (N_1969,N_1377,N_1355);
nor U1970 (N_1970,N_1213,N_1027);
nand U1971 (N_1971,N_1497,N_795);
xnor U1972 (N_1972,N_922,N_1145);
or U1973 (N_1973,N_975,N_1302);
or U1974 (N_1974,N_760,N_961);
and U1975 (N_1975,N_1278,N_862);
or U1976 (N_1976,N_823,N_1149);
xor U1977 (N_1977,N_1068,N_807);
or U1978 (N_1978,N_1340,N_1346);
nor U1979 (N_1979,N_1334,N_1064);
nor U1980 (N_1980,N_1412,N_1338);
nor U1981 (N_1981,N_953,N_813);
nand U1982 (N_1982,N_763,N_909);
and U1983 (N_1983,N_1294,N_1089);
nand U1984 (N_1984,N_811,N_988);
xnor U1985 (N_1985,N_1031,N_1132);
xor U1986 (N_1986,N_1373,N_1323);
nor U1987 (N_1987,N_888,N_1289);
xnor U1988 (N_1988,N_762,N_767);
nor U1989 (N_1989,N_1203,N_897);
and U1990 (N_1990,N_1349,N_1461);
or U1991 (N_1991,N_1121,N_953);
xnor U1992 (N_1992,N_1112,N_1287);
and U1993 (N_1993,N_1140,N_1160);
xor U1994 (N_1994,N_1123,N_1205);
nand U1995 (N_1995,N_1111,N_1258);
nor U1996 (N_1996,N_1153,N_1005);
xor U1997 (N_1997,N_999,N_1233);
nand U1998 (N_1998,N_1290,N_1111);
or U1999 (N_1999,N_1002,N_977);
nor U2000 (N_2000,N_1301,N_975);
xor U2001 (N_2001,N_1357,N_939);
or U2002 (N_2002,N_1189,N_981);
nor U2003 (N_2003,N_1423,N_1331);
or U2004 (N_2004,N_1468,N_1273);
and U2005 (N_2005,N_950,N_1000);
xor U2006 (N_2006,N_830,N_944);
nor U2007 (N_2007,N_1106,N_1278);
and U2008 (N_2008,N_987,N_1078);
and U2009 (N_2009,N_1140,N_1173);
nand U2010 (N_2010,N_1010,N_911);
nand U2011 (N_2011,N_1265,N_817);
or U2012 (N_2012,N_1321,N_1079);
or U2013 (N_2013,N_1316,N_1462);
and U2014 (N_2014,N_1155,N_1118);
nand U2015 (N_2015,N_1061,N_820);
and U2016 (N_2016,N_1184,N_1400);
nor U2017 (N_2017,N_1072,N_963);
xnor U2018 (N_2018,N_992,N_1442);
nor U2019 (N_2019,N_1306,N_1440);
nand U2020 (N_2020,N_1242,N_980);
nand U2021 (N_2021,N_1324,N_1091);
or U2022 (N_2022,N_948,N_1423);
and U2023 (N_2023,N_1166,N_1011);
or U2024 (N_2024,N_777,N_1317);
and U2025 (N_2025,N_996,N_783);
nand U2026 (N_2026,N_1454,N_1067);
or U2027 (N_2027,N_1171,N_1130);
nor U2028 (N_2028,N_1429,N_1284);
and U2029 (N_2029,N_1237,N_1018);
nand U2030 (N_2030,N_805,N_962);
xor U2031 (N_2031,N_1043,N_1499);
xnor U2032 (N_2032,N_1307,N_1472);
nor U2033 (N_2033,N_1383,N_1246);
or U2034 (N_2034,N_1158,N_756);
nor U2035 (N_2035,N_911,N_1121);
nor U2036 (N_2036,N_1447,N_890);
nor U2037 (N_2037,N_1278,N_1413);
nand U2038 (N_2038,N_922,N_762);
xnor U2039 (N_2039,N_933,N_1167);
nand U2040 (N_2040,N_1495,N_1390);
or U2041 (N_2041,N_911,N_1072);
nor U2042 (N_2042,N_771,N_1485);
nand U2043 (N_2043,N_1316,N_1273);
xnor U2044 (N_2044,N_874,N_807);
nand U2045 (N_2045,N_771,N_858);
nor U2046 (N_2046,N_881,N_1172);
xor U2047 (N_2047,N_1010,N_1140);
nor U2048 (N_2048,N_1070,N_1098);
nor U2049 (N_2049,N_1004,N_1318);
nor U2050 (N_2050,N_1265,N_807);
and U2051 (N_2051,N_1475,N_1483);
nor U2052 (N_2052,N_1469,N_812);
and U2053 (N_2053,N_758,N_1060);
or U2054 (N_2054,N_1366,N_1114);
and U2055 (N_2055,N_1288,N_1345);
xnor U2056 (N_2056,N_1230,N_1294);
xor U2057 (N_2057,N_880,N_810);
and U2058 (N_2058,N_812,N_1120);
or U2059 (N_2059,N_827,N_1178);
and U2060 (N_2060,N_1260,N_1479);
nor U2061 (N_2061,N_1341,N_1307);
or U2062 (N_2062,N_991,N_1315);
or U2063 (N_2063,N_1254,N_1351);
or U2064 (N_2064,N_842,N_846);
or U2065 (N_2065,N_1251,N_1013);
xor U2066 (N_2066,N_1039,N_1174);
nand U2067 (N_2067,N_803,N_1469);
nor U2068 (N_2068,N_1158,N_848);
nand U2069 (N_2069,N_872,N_945);
nor U2070 (N_2070,N_1463,N_1160);
and U2071 (N_2071,N_1458,N_1043);
or U2072 (N_2072,N_1184,N_902);
nand U2073 (N_2073,N_796,N_1304);
xnor U2074 (N_2074,N_1031,N_1258);
and U2075 (N_2075,N_1142,N_1288);
xor U2076 (N_2076,N_1246,N_1247);
xnor U2077 (N_2077,N_1375,N_1105);
and U2078 (N_2078,N_947,N_869);
or U2079 (N_2079,N_1221,N_1100);
xnor U2080 (N_2080,N_1172,N_842);
or U2081 (N_2081,N_783,N_895);
or U2082 (N_2082,N_1360,N_1165);
and U2083 (N_2083,N_1050,N_1178);
nor U2084 (N_2084,N_1288,N_1164);
nand U2085 (N_2085,N_1313,N_1273);
or U2086 (N_2086,N_934,N_1254);
nand U2087 (N_2087,N_1455,N_1407);
nand U2088 (N_2088,N_1401,N_897);
nand U2089 (N_2089,N_1269,N_1362);
nand U2090 (N_2090,N_1406,N_1207);
nor U2091 (N_2091,N_948,N_1358);
and U2092 (N_2092,N_1190,N_1075);
nor U2093 (N_2093,N_1049,N_924);
nand U2094 (N_2094,N_834,N_1326);
nor U2095 (N_2095,N_1119,N_1495);
and U2096 (N_2096,N_1127,N_1343);
nand U2097 (N_2097,N_1367,N_1294);
nand U2098 (N_2098,N_1076,N_1077);
nor U2099 (N_2099,N_1412,N_766);
xor U2100 (N_2100,N_1257,N_1195);
xnor U2101 (N_2101,N_1429,N_1384);
nor U2102 (N_2102,N_1495,N_1299);
and U2103 (N_2103,N_956,N_1462);
nor U2104 (N_2104,N_791,N_1354);
nor U2105 (N_2105,N_897,N_1160);
and U2106 (N_2106,N_786,N_1494);
or U2107 (N_2107,N_1189,N_1254);
nor U2108 (N_2108,N_989,N_1402);
and U2109 (N_2109,N_1468,N_1386);
or U2110 (N_2110,N_1129,N_1400);
nor U2111 (N_2111,N_1220,N_821);
nor U2112 (N_2112,N_1104,N_1075);
nand U2113 (N_2113,N_778,N_1425);
and U2114 (N_2114,N_921,N_1204);
nand U2115 (N_2115,N_1005,N_865);
nand U2116 (N_2116,N_1202,N_1130);
nand U2117 (N_2117,N_986,N_1054);
nand U2118 (N_2118,N_899,N_800);
or U2119 (N_2119,N_1456,N_818);
nor U2120 (N_2120,N_830,N_778);
and U2121 (N_2121,N_1183,N_1078);
and U2122 (N_2122,N_1496,N_813);
or U2123 (N_2123,N_1138,N_851);
xor U2124 (N_2124,N_822,N_1188);
or U2125 (N_2125,N_1103,N_1425);
nor U2126 (N_2126,N_764,N_1038);
and U2127 (N_2127,N_1304,N_1290);
nand U2128 (N_2128,N_768,N_942);
nor U2129 (N_2129,N_799,N_1277);
xor U2130 (N_2130,N_1192,N_1095);
or U2131 (N_2131,N_1438,N_1276);
and U2132 (N_2132,N_966,N_1137);
xor U2133 (N_2133,N_1281,N_1050);
nor U2134 (N_2134,N_798,N_1002);
xor U2135 (N_2135,N_976,N_1026);
xnor U2136 (N_2136,N_938,N_1456);
nor U2137 (N_2137,N_1248,N_1164);
xnor U2138 (N_2138,N_1012,N_1225);
or U2139 (N_2139,N_1184,N_1417);
nor U2140 (N_2140,N_1336,N_1056);
or U2141 (N_2141,N_1322,N_1203);
nor U2142 (N_2142,N_902,N_1365);
nand U2143 (N_2143,N_899,N_995);
or U2144 (N_2144,N_1153,N_822);
or U2145 (N_2145,N_989,N_1080);
or U2146 (N_2146,N_1297,N_1017);
and U2147 (N_2147,N_1478,N_1133);
and U2148 (N_2148,N_1450,N_1371);
and U2149 (N_2149,N_1048,N_1360);
and U2150 (N_2150,N_1375,N_1301);
xnor U2151 (N_2151,N_1410,N_1242);
xnor U2152 (N_2152,N_1367,N_988);
or U2153 (N_2153,N_761,N_917);
xnor U2154 (N_2154,N_1161,N_954);
nand U2155 (N_2155,N_1223,N_968);
nand U2156 (N_2156,N_1332,N_1252);
nand U2157 (N_2157,N_1101,N_1454);
nand U2158 (N_2158,N_1487,N_1215);
or U2159 (N_2159,N_788,N_945);
and U2160 (N_2160,N_907,N_1122);
nor U2161 (N_2161,N_868,N_1151);
or U2162 (N_2162,N_1346,N_1364);
nor U2163 (N_2163,N_1007,N_1213);
xor U2164 (N_2164,N_955,N_1327);
nor U2165 (N_2165,N_963,N_1241);
nand U2166 (N_2166,N_778,N_1265);
and U2167 (N_2167,N_1217,N_1278);
xor U2168 (N_2168,N_1120,N_1393);
xnor U2169 (N_2169,N_1108,N_1364);
nand U2170 (N_2170,N_1264,N_1439);
and U2171 (N_2171,N_886,N_1470);
xnor U2172 (N_2172,N_839,N_1149);
or U2173 (N_2173,N_752,N_1481);
nor U2174 (N_2174,N_1488,N_1484);
nand U2175 (N_2175,N_1293,N_1439);
nand U2176 (N_2176,N_994,N_1169);
nand U2177 (N_2177,N_1248,N_1497);
nor U2178 (N_2178,N_834,N_1236);
nor U2179 (N_2179,N_1109,N_1455);
nor U2180 (N_2180,N_1435,N_1328);
and U2181 (N_2181,N_1182,N_1114);
xnor U2182 (N_2182,N_1136,N_1429);
nand U2183 (N_2183,N_1476,N_1059);
xnor U2184 (N_2184,N_997,N_839);
nand U2185 (N_2185,N_1467,N_1099);
nor U2186 (N_2186,N_822,N_857);
or U2187 (N_2187,N_1035,N_1393);
xor U2188 (N_2188,N_771,N_914);
and U2189 (N_2189,N_827,N_1375);
nor U2190 (N_2190,N_955,N_1470);
nor U2191 (N_2191,N_809,N_1256);
xnor U2192 (N_2192,N_839,N_1266);
nand U2193 (N_2193,N_1402,N_781);
nand U2194 (N_2194,N_1375,N_754);
or U2195 (N_2195,N_1290,N_923);
and U2196 (N_2196,N_1330,N_819);
nor U2197 (N_2197,N_1334,N_1128);
and U2198 (N_2198,N_760,N_994);
or U2199 (N_2199,N_1175,N_1274);
nand U2200 (N_2200,N_1265,N_1270);
nand U2201 (N_2201,N_1120,N_1410);
or U2202 (N_2202,N_1155,N_1334);
nand U2203 (N_2203,N_1304,N_860);
xnor U2204 (N_2204,N_928,N_1359);
nor U2205 (N_2205,N_1099,N_1487);
or U2206 (N_2206,N_1442,N_1397);
or U2207 (N_2207,N_999,N_1437);
or U2208 (N_2208,N_1423,N_1405);
nor U2209 (N_2209,N_818,N_860);
or U2210 (N_2210,N_1055,N_763);
or U2211 (N_2211,N_781,N_917);
xor U2212 (N_2212,N_1152,N_1178);
or U2213 (N_2213,N_1392,N_1440);
or U2214 (N_2214,N_1063,N_1407);
xor U2215 (N_2215,N_844,N_1494);
or U2216 (N_2216,N_1328,N_1152);
or U2217 (N_2217,N_920,N_1187);
nor U2218 (N_2218,N_1307,N_1063);
and U2219 (N_2219,N_756,N_1306);
nor U2220 (N_2220,N_1332,N_1027);
or U2221 (N_2221,N_1211,N_994);
xor U2222 (N_2222,N_1045,N_1496);
or U2223 (N_2223,N_850,N_965);
or U2224 (N_2224,N_1304,N_1127);
xnor U2225 (N_2225,N_838,N_1076);
xnor U2226 (N_2226,N_844,N_1242);
nor U2227 (N_2227,N_1381,N_1296);
or U2228 (N_2228,N_1380,N_1172);
xor U2229 (N_2229,N_758,N_1327);
or U2230 (N_2230,N_873,N_870);
nand U2231 (N_2231,N_1396,N_1178);
or U2232 (N_2232,N_1157,N_1127);
or U2233 (N_2233,N_1305,N_1162);
nor U2234 (N_2234,N_1475,N_1146);
and U2235 (N_2235,N_1110,N_1156);
and U2236 (N_2236,N_1425,N_1443);
and U2237 (N_2237,N_1213,N_1196);
nand U2238 (N_2238,N_1254,N_1071);
nor U2239 (N_2239,N_1291,N_1273);
or U2240 (N_2240,N_1133,N_1225);
or U2241 (N_2241,N_1285,N_1051);
nand U2242 (N_2242,N_1368,N_875);
nand U2243 (N_2243,N_1008,N_1184);
nor U2244 (N_2244,N_1291,N_856);
or U2245 (N_2245,N_1332,N_855);
nor U2246 (N_2246,N_1256,N_1149);
nor U2247 (N_2247,N_791,N_1187);
nor U2248 (N_2248,N_910,N_1252);
nor U2249 (N_2249,N_1116,N_1461);
nor U2250 (N_2250,N_1706,N_2041);
xnor U2251 (N_2251,N_2089,N_2155);
and U2252 (N_2252,N_1523,N_2006);
or U2253 (N_2253,N_1661,N_1692);
and U2254 (N_2254,N_1936,N_1537);
or U2255 (N_2255,N_1805,N_1818);
nand U2256 (N_2256,N_1753,N_1509);
nand U2257 (N_2257,N_1823,N_1865);
nand U2258 (N_2258,N_1882,N_1991);
nand U2259 (N_2259,N_1717,N_1644);
or U2260 (N_2260,N_2170,N_1867);
nand U2261 (N_2261,N_2037,N_1983);
and U2262 (N_2262,N_1530,N_1840);
or U2263 (N_2263,N_2192,N_2118);
nor U2264 (N_2264,N_1768,N_1819);
xnor U2265 (N_2265,N_2227,N_2177);
xor U2266 (N_2266,N_1709,N_1951);
or U2267 (N_2267,N_1757,N_2003);
xor U2268 (N_2268,N_1653,N_2033);
nor U2269 (N_2269,N_1816,N_2190);
nand U2270 (N_2270,N_1890,N_2233);
xnor U2271 (N_2271,N_1993,N_2107);
nor U2272 (N_2272,N_1813,N_1538);
nor U2273 (N_2273,N_1939,N_1617);
or U2274 (N_2274,N_2034,N_2103);
nand U2275 (N_2275,N_1596,N_2054);
xnor U2276 (N_2276,N_1919,N_2012);
and U2277 (N_2277,N_1806,N_1884);
and U2278 (N_2278,N_2130,N_2174);
and U2279 (N_2279,N_2182,N_2204);
or U2280 (N_2280,N_1728,N_2042);
nand U2281 (N_2281,N_2168,N_1896);
or U2282 (N_2282,N_1933,N_1871);
xnor U2283 (N_2283,N_2196,N_1658);
nor U2284 (N_2284,N_2163,N_2117);
nor U2285 (N_2285,N_1914,N_1662);
xnor U2286 (N_2286,N_2028,N_1995);
nor U2287 (N_2287,N_2077,N_1925);
nor U2288 (N_2288,N_1718,N_2005);
nor U2289 (N_2289,N_1854,N_2022);
or U2290 (N_2290,N_1513,N_1756);
or U2291 (N_2291,N_1879,N_1640);
nor U2292 (N_2292,N_1698,N_2166);
or U2293 (N_2293,N_1752,N_1830);
and U2294 (N_2294,N_2154,N_1949);
and U2295 (N_2295,N_2181,N_1808);
or U2296 (N_2296,N_2193,N_1671);
or U2297 (N_2297,N_1916,N_1541);
or U2298 (N_2298,N_1815,N_1520);
xnor U2299 (N_2299,N_1736,N_1976);
and U2300 (N_2300,N_1587,N_1743);
nor U2301 (N_2301,N_2208,N_1650);
xor U2302 (N_2302,N_1906,N_1584);
or U2303 (N_2303,N_2020,N_2113);
nand U2304 (N_2304,N_2071,N_1901);
xnor U2305 (N_2305,N_1900,N_1626);
nor U2306 (N_2306,N_1895,N_1997);
nand U2307 (N_2307,N_1804,N_1544);
or U2308 (N_2308,N_2026,N_1668);
or U2309 (N_2309,N_1712,N_2156);
and U2310 (N_2310,N_1777,N_1585);
nor U2311 (N_2311,N_2220,N_1690);
nor U2312 (N_2312,N_1562,N_1855);
nand U2313 (N_2313,N_1631,N_2091);
nand U2314 (N_2314,N_1968,N_2235);
nand U2315 (N_2315,N_1826,N_1674);
or U2316 (N_2316,N_1892,N_2200);
and U2317 (N_2317,N_1829,N_1904);
and U2318 (N_2318,N_1985,N_1528);
nand U2319 (N_2319,N_2141,N_1740);
and U2320 (N_2320,N_1580,N_1902);
xor U2321 (N_2321,N_1858,N_2145);
nand U2322 (N_2322,N_1911,N_1570);
xnor U2323 (N_2323,N_1921,N_2068);
or U2324 (N_2324,N_1682,N_2194);
xor U2325 (N_2325,N_2223,N_2218);
and U2326 (N_2326,N_1848,N_2161);
and U2327 (N_2327,N_2102,N_1885);
nand U2328 (N_2328,N_1694,N_2053);
or U2329 (N_2329,N_1713,N_1772);
and U2330 (N_2330,N_1611,N_1665);
xnor U2331 (N_2331,N_1536,N_2189);
xor U2332 (N_2332,N_1844,N_1605);
nor U2333 (N_2333,N_2184,N_1504);
or U2334 (N_2334,N_1832,N_1930);
nand U2335 (N_2335,N_1500,N_1646);
or U2336 (N_2336,N_1586,N_1681);
or U2337 (N_2337,N_1648,N_1917);
xor U2338 (N_2338,N_1510,N_1572);
nor U2339 (N_2339,N_1573,N_1702);
xor U2340 (N_2340,N_1783,N_1856);
xor U2341 (N_2341,N_1851,N_2008);
and U2342 (N_2342,N_2221,N_2225);
xnor U2343 (N_2343,N_2086,N_1569);
nand U2344 (N_2344,N_1566,N_1834);
and U2345 (N_2345,N_1872,N_2110);
or U2346 (N_2346,N_1874,N_1628);
nand U2347 (N_2347,N_1934,N_1532);
nor U2348 (N_2348,N_1618,N_2224);
or U2349 (N_2349,N_1591,N_2176);
and U2350 (N_2350,N_1685,N_1927);
or U2351 (N_2351,N_1535,N_2134);
nor U2352 (N_2352,N_1669,N_1620);
xnor U2353 (N_2353,N_1947,N_1994);
xor U2354 (N_2354,N_1775,N_2180);
or U2355 (N_2355,N_2125,N_1634);
xor U2356 (N_2356,N_1602,N_1898);
nor U2357 (N_2357,N_1771,N_2013);
nor U2358 (N_2358,N_1866,N_1747);
or U2359 (N_2359,N_1864,N_1937);
nand U2360 (N_2360,N_2032,N_2081);
nand U2361 (N_2361,N_1543,N_1796);
or U2362 (N_2362,N_1691,N_2001);
nor U2363 (N_2363,N_2052,N_1522);
or U2364 (N_2364,N_1999,N_2245);
nor U2365 (N_2365,N_1836,N_1894);
nor U2366 (N_2366,N_2215,N_1781);
nand U2367 (N_2367,N_2136,N_1652);
or U2368 (N_2368,N_2098,N_2138);
or U2369 (N_2369,N_1589,N_2109);
nand U2370 (N_2370,N_2160,N_1920);
nand U2371 (N_2371,N_1732,N_2228);
and U2372 (N_2372,N_1735,N_2165);
nor U2373 (N_2373,N_1956,N_1784);
xor U2374 (N_2374,N_1779,N_1827);
or U2375 (N_2375,N_1553,N_1770);
nor U2376 (N_2376,N_1769,N_2124);
and U2377 (N_2377,N_1825,N_1643);
and U2378 (N_2378,N_1579,N_2039);
xor U2379 (N_2379,N_1765,N_1737);
nand U2380 (N_2380,N_1787,N_2007);
nor U2381 (N_2381,N_2048,N_2159);
nand U2382 (N_2382,N_2179,N_2056);
and U2383 (N_2383,N_2019,N_1555);
nor U2384 (N_2384,N_1824,N_1660);
xor U2385 (N_2385,N_1869,N_1636);
nand U2386 (N_2386,N_1593,N_2164);
and U2387 (N_2387,N_2199,N_2188);
nand U2388 (N_2388,N_2072,N_2214);
xor U2389 (N_2389,N_1946,N_1749);
nor U2390 (N_2390,N_1567,N_2011);
xnor U2391 (N_2391,N_1963,N_1820);
and U2392 (N_2392,N_2240,N_1727);
and U2393 (N_2393,N_1683,N_1563);
or U2394 (N_2394,N_1533,N_1501);
and U2395 (N_2395,N_1529,N_1928);
and U2396 (N_2396,N_1881,N_2187);
or U2397 (N_2397,N_1809,N_1801);
xor U2398 (N_2398,N_1974,N_2079);
xor U2399 (N_2399,N_1812,N_1868);
nor U2400 (N_2400,N_2151,N_1721);
or U2401 (N_2401,N_1785,N_2016);
nand U2402 (N_2402,N_1739,N_1597);
xnor U2403 (N_2403,N_1959,N_2060);
xnor U2404 (N_2404,N_1613,N_1512);
nor U2405 (N_2405,N_2206,N_1641);
xnor U2406 (N_2406,N_1670,N_1950);
and U2407 (N_2407,N_2241,N_1745);
or U2408 (N_2408,N_1595,N_1847);
nor U2409 (N_2409,N_1942,N_2062);
and U2410 (N_2410,N_2146,N_2015);
and U2411 (N_2411,N_1841,N_1688);
xor U2412 (N_2412,N_1516,N_1755);
nor U2413 (N_2413,N_1701,N_1657);
or U2414 (N_2414,N_2096,N_1507);
or U2415 (N_2415,N_1984,N_2036);
nand U2416 (N_2416,N_2129,N_1664);
and U2417 (N_2417,N_1792,N_2158);
xor U2418 (N_2418,N_1857,N_1799);
xnor U2419 (N_2419,N_1515,N_2122);
nor U2420 (N_2420,N_2067,N_1511);
nor U2421 (N_2421,N_1789,N_2152);
xnor U2422 (N_2422,N_1738,N_2093);
nand U2423 (N_2423,N_1838,N_1565);
xnor U2424 (N_2424,N_1550,N_2197);
and U2425 (N_2425,N_2069,N_1655);
or U2426 (N_2426,N_2135,N_1932);
nand U2427 (N_2427,N_2234,N_1955);
or U2428 (N_2428,N_2116,N_2104);
nor U2429 (N_2429,N_2078,N_1810);
nor U2430 (N_2430,N_2148,N_1659);
xnor U2431 (N_2431,N_2216,N_2131);
nand U2432 (N_2432,N_1996,N_2202);
or U2433 (N_2433,N_2066,N_1548);
nor U2434 (N_2434,N_1645,N_1619);
xnor U2435 (N_2435,N_1758,N_1850);
and U2436 (N_2436,N_2178,N_1908);
nand U2437 (N_2437,N_1680,N_1803);
and U2438 (N_2438,N_1534,N_1577);
and U2439 (N_2439,N_1606,N_1891);
nand U2440 (N_2440,N_1524,N_1609);
nand U2441 (N_2441,N_1922,N_1977);
nor U2442 (N_2442,N_2108,N_1964);
and U2443 (N_2443,N_2211,N_2140);
and U2444 (N_2444,N_1817,N_2043);
and U2445 (N_2445,N_2201,N_1807);
and U2446 (N_2446,N_2172,N_1731);
or U2447 (N_2447,N_1849,N_1910);
nor U2448 (N_2448,N_1859,N_1853);
or U2449 (N_2449,N_1907,N_1663);
nand U2450 (N_2450,N_1845,N_1887);
or U2451 (N_2451,N_2099,N_1633);
and U2452 (N_2452,N_2047,N_2112);
or U2453 (N_2453,N_1554,N_2120);
nor U2454 (N_2454,N_1893,N_1592);
and U2455 (N_2455,N_1734,N_1981);
nand U2456 (N_2456,N_1635,N_2065);
or U2457 (N_2457,N_1962,N_2186);
nor U2458 (N_2458,N_1998,N_2213);
xor U2459 (N_2459,N_2173,N_1839);
and U2460 (N_2460,N_1912,N_1647);
nand U2461 (N_2461,N_1821,N_1940);
nand U2462 (N_2462,N_1601,N_1831);
or U2463 (N_2463,N_2029,N_1835);
xor U2464 (N_2464,N_2243,N_1899);
and U2465 (N_2465,N_1935,N_1542);
nor U2466 (N_2466,N_1989,N_1588);
nand U2467 (N_2467,N_1707,N_1627);
nand U2468 (N_2468,N_1654,N_1873);
or U2469 (N_2469,N_1557,N_1514);
xnor U2470 (N_2470,N_1766,N_1764);
and U2471 (N_2471,N_2080,N_1651);
xor U2472 (N_2472,N_1625,N_1623);
or U2473 (N_2473,N_1878,N_1795);
xnor U2474 (N_2474,N_1979,N_1941);
nand U2475 (N_2475,N_1750,N_1571);
nor U2476 (N_2476,N_1621,N_2239);
nor U2477 (N_2477,N_1666,N_2046);
or U2478 (N_2478,N_1726,N_1742);
or U2479 (N_2479,N_1695,N_2030);
nor U2480 (N_2480,N_2142,N_2105);
nand U2481 (N_2481,N_1614,N_1677);
and U2482 (N_2482,N_1583,N_2111);
or U2483 (N_2483,N_1748,N_2126);
nand U2484 (N_2484,N_2021,N_1797);
nor U2485 (N_2485,N_2205,N_1700);
nor U2486 (N_2486,N_2088,N_1988);
xnor U2487 (N_2487,N_1679,N_1773);
or U2488 (N_2488,N_1790,N_1699);
nor U2489 (N_2489,N_1967,N_2232);
nor U2490 (N_2490,N_1876,N_1926);
nor U2491 (N_2491,N_1886,N_2024);
or U2492 (N_2492,N_1696,N_1719);
or U2493 (N_2493,N_2010,N_1561);
and U2494 (N_2494,N_1776,N_1880);
xnor U2495 (N_2495,N_1610,N_1877);
nor U2496 (N_2496,N_1608,N_1576);
nand U2497 (N_2497,N_1972,N_1547);
xor U2498 (N_2498,N_2175,N_2242);
nand U2499 (N_2499,N_1637,N_1704);
or U2500 (N_2500,N_1990,N_2229);
nand U2501 (N_2501,N_1708,N_1929);
nor U2502 (N_2502,N_1710,N_1822);
nand U2503 (N_2503,N_1711,N_1889);
nor U2504 (N_2504,N_2185,N_2035);
nand U2505 (N_2505,N_1924,N_1656);
nand U2506 (N_2506,N_2219,N_2094);
nand U2507 (N_2507,N_1675,N_2040);
nor U2508 (N_2508,N_1842,N_2147);
nor U2509 (N_2509,N_2133,N_1551);
nand U2510 (N_2510,N_2017,N_1630);
and U2511 (N_2511,N_2023,N_2127);
xor U2512 (N_2512,N_1600,N_1705);
and U2513 (N_2513,N_1870,N_1986);
xnor U2514 (N_2514,N_1545,N_1761);
xor U2515 (N_2515,N_2203,N_1837);
xnor U2516 (N_2516,N_1556,N_2100);
or U2517 (N_2517,N_1746,N_2123);
nand U2518 (N_2518,N_2082,N_1560);
or U2519 (N_2519,N_1508,N_2097);
and U2520 (N_2520,N_1791,N_1574);
nand U2521 (N_2521,N_2244,N_1686);
or U2522 (N_2522,N_1843,N_2195);
or U2523 (N_2523,N_2132,N_1754);
and U2524 (N_2524,N_1794,N_1763);
xnor U2525 (N_2525,N_2045,N_2063);
or U2526 (N_2526,N_1525,N_1527);
or U2527 (N_2527,N_1505,N_1943);
or U2528 (N_2528,N_1923,N_1944);
and U2529 (N_2529,N_1578,N_1519);
nor U2530 (N_2530,N_1875,N_1622);
xnor U2531 (N_2531,N_2231,N_1774);
nand U2532 (N_2532,N_1506,N_2064);
xor U2533 (N_2533,N_1552,N_1862);
nor U2534 (N_2534,N_1715,N_1684);
and U2535 (N_2535,N_2237,N_1639);
nand U2536 (N_2536,N_1828,N_1973);
and U2537 (N_2537,N_1975,N_1960);
and U2538 (N_2538,N_1649,N_2238);
and U2539 (N_2539,N_2115,N_2198);
and U2540 (N_2540,N_1594,N_2018);
or U2541 (N_2541,N_1539,N_2246);
xnor U2542 (N_2542,N_2002,N_1833);
or U2543 (N_2543,N_1720,N_1852);
and U2544 (N_2544,N_1948,N_1678);
nand U2545 (N_2545,N_2055,N_1980);
xor U2546 (N_2546,N_2143,N_1915);
or U2547 (N_2547,N_2084,N_1759);
nand U2548 (N_2548,N_1978,N_2038);
xor U2549 (N_2549,N_1612,N_2073);
nor U2550 (N_2550,N_1966,N_1970);
xor U2551 (N_2551,N_2004,N_2247);
and U2552 (N_2552,N_1760,N_2083);
nor U2553 (N_2553,N_1800,N_1793);
and U2554 (N_2554,N_2114,N_1909);
xnor U2555 (N_2555,N_1778,N_2087);
or U2556 (N_2556,N_1992,N_1938);
nor U2557 (N_2557,N_2000,N_1861);
and U2558 (N_2558,N_1863,N_1559);
or U2559 (N_2559,N_1518,N_2058);
nor U2560 (N_2560,N_1604,N_2049);
xor U2561 (N_2561,N_1786,N_1897);
or U2562 (N_2562,N_1762,N_2144);
or U2563 (N_2563,N_1582,N_1540);
nor U2564 (N_2564,N_2076,N_1767);
or U2565 (N_2565,N_2169,N_2217);
xnor U2566 (N_2566,N_1521,N_1811);
xor U2567 (N_2567,N_1733,N_2230);
or U2568 (N_2568,N_1971,N_2207);
nor U2569 (N_2569,N_1603,N_1503);
and U2570 (N_2570,N_2150,N_1599);
or U2571 (N_2571,N_2014,N_1846);
xnor U2572 (N_2572,N_1958,N_1729);
nand U2573 (N_2573,N_2248,N_2212);
xnor U2574 (N_2574,N_1689,N_1517);
or U2575 (N_2575,N_1741,N_1730);
nor U2576 (N_2576,N_2209,N_1632);
nor U2577 (N_2577,N_2075,N_1502);
nor U2578 (N_2578,N_1982,N_2121);
nand U2579 (N_2579,N_1575,N_1624);
xor U2580 (N_2580,N_1581,N_2171);
nand U2581 (N_2581,N_1987,N_2095);
xor U2582 (N_2582,N_1802,N_1903);
nor U2583 (N_2583,N_1905,N_2050);
or U2584 (N_2584,N_2092,N_1782);
xnor U2585 (N_2585,N_1931,N_2070);
nand U2586 (N_2586,N_2149,N_2157);
nor U2587 (N_2587,N_1744,N_2074);
nand U2588 (N_2588,N_2101,N_1615);
or U2589 (N_2589,N_1888,N_1883);
nor U2590 (N_2590,N_1952,N_1687);
nand U2591 (N_2591,N_1969,N_1714);
or U2592 (N_2592,N_2137,N_1629);
nand U2593 (N_2593,N_2222,N_1798);
nand U2594 (N_2594,N_1780,N_1672);
nor U2595 (N_2595,N_1693,N_1546);
nor U2596 (N_2596,N_2153,N_1526);
nor U2597 (N_2597,N_1642,N_2119);
xnor U2598 (N_2598,N_2139,N_1722);
nand U2599 (N_2599,N_2090,N_1616);
nor U2600 (N_2600,N_2009,N_2061);
xor U2601 (N_2601,N_1957,N_1697);
and U2602 (N_2602,N_1568,N_2236);
nor U2603 (N_2603,N_1751,N_2057);
nand U2604 (N_2604,N_2027,N_1590);
or U2605 (N_2605,N_1598,N_2106);
xor U2606 (N_2606,N_1945,N_1531);
xnor U2607 (N_2607,N_1965,N_2051);
or U2608 (N_2608,N_1814,N_2226);
or U2609 (N_2609,N_1724,N_1961);
xnor U2610 (N_2610,N_1673,N_1918);
xor U2611 (N_2611,N_1860,N_1716);
xor U2612 (N_2612,N_1564,N_2128);
and U2613 (N_2613,N_2059,N_2085);
xnor U2614 (N_2614,N_1607,N_2191);
or U2615 (N_2615,N_1723,N_1953);
nor U2616 (N_2616,N_2044,N_2167);
or U2617 (N_2617,N_2031,N_1549);
and U2618 (N_2618,N_1667,N_2025);
nand U2619 (N_2619,N_1954,N_1788);
or U2620 (N_2620,N_1725,N_1676);
nand U2621 (N_2621,N_2183,N_1703);
and U2622 (N_2622,N_1913,N_1558);
or U2623 (N_2623,N_2210,N_2249);
xor U2624 (N_2624,N_1638,N_2162);
and U2625 (N_2625,N_1704,N_1549);
or U2626 (N_2626,N_1660,N_1585);
nand U2627 (N_2627,N_1798,N_1556);
or U2628 (N_2628,N_1889,N_1631);
xnor U2629 (N_2629,N_2193,N_2151);
and U2630 (N_2630,N_1998,N_1742);
xnor U2631 (N_2631,N_1975,N_1950);
or U2632 (N_2632,N_1674,N_2157);
or U2633 (N_2633,N_1954,N_2157);
xnor U2634 (N_2634,N_1656,N_1847);
nand U2635 (N_2635,N_2245,N_1812);
or U2636 (N_2636,N_1710,N_2166);
xnor U2637 (N_2637,N_2118,N_1790);
nor U2638 (N_2638,N_2085,N_2241);
xor U2639 (N_2639,N_1896,N_2117);
xor U2640 (N_2640,N_2008,N_2247);
or U2641 (N_2641,N_1677,N_1860);
or U2642 (N_2642,N_2074,N_1997);
and U2643 (N_2643,N_2198,N_1926);
nor U2644 (N_2644,N_1532,N_1686);
nand U2645 (N_2645,N_1540,N_1799);
nor U2646 (N_2646,N_2012,N_1846);
or U2647 (N_2647,N_2102,N_1603);
or U2648 (N_2648,N_1764,N_1583);
nand U2649 (N_2649,N_1758,N_1514);
nand U2650 (N_2650,N_1508,N_1763);
xor U2651 (N_2651,N_2079,N_2238);
xor U2652 (N_2652,N_1603,N_1740);
nor U2653 (N_2653,N_2044,N_1739);
nor U2654 (N_2654,N_2103,N_2177);
xor U2655 (N_2655,N_2188,N_1813);
xnor U2656 (N_2656,N_1816,N_1632);
nor U2657 (N_2657,N_1600,N_1613);
or U2658 (N_2658,N_2032,N_1737);
nor U2659 (N_2659,N_2217,N_2092);
and U2660 (N_2660,N_1752,N_1614);
nand U2661 (N_2661,N_1638,N_1728);
or U2662 (N_2662,N_2138,N_1617);
nor U2663 (N_2663,N_1696,N_1670);
nor U2664 (N_2664,N_1985,N_1723);
nand U2665 (N_2665,N_2031,N_1543);
nor U2666 (N_2666,N_1672,N_1598);
nor U2667 (N_2667,N_1883,N_1920);
or U2668 (N_2668,N_1627,N_1827);
or U2669 (N_2669,N_1699,N_2033);
nand U2670 (N_2670,N_1723,N_2061);
xor U2671 (N_2671,N_1758,N_1555);
or U2672 (N_2672,N_1927,N_1578);
or U2673 (N_2673,N_2026,N_1698);
and U2674 (N_2674,N_2090,N_1893);
nor U2675 (N_2675,N_1856,N_2015);
nand U2676 (N_2676,N_1767,N_1793);
or U2677 (N_2677,N_1828,N_2103);
or U2678 (N_2678,N_1976,N_1856);
or U2679 (N_2679,N_1920,N_1696);
or U2680 (N_2680,N_1643,N_2043);
nor U2681 (N_2681,N_1752,N_1713);
nor U2682 (N_2682,N_2071,N_1897);
or U2683 (N_2683,N_2127,N_1701);
and U2684 (N_2684,N_1735,N_2005);
or U2685 (N_2685,N_2228,N_1597);
nand U2686 (N_2686,N_2218,N_1569);
or U2687 (N_2687,N_2148,N_1558);
xnor U2688 (N_2688,N_2228,N_1514);
nor U2689 (N_2689,N_2136,N_2181);
and U2690 (N_2690,N_1729,N_2094);
nand U2691 (N_2691,N_1744,N_1706);
or U2692 (N_2692,N_1728,N_2232);
nand U2693 (N_2693,N_1869,N_1942);
xor U2694 (N_2694,N_1681,N_2145);
and U2695 (N_2695,N_1802,N_2180);
or U2696 (N_2696,N_2005,N_2028);
nand U2697 (N_2697,N_1944,N_2179);
or U2698 (N_2698,N_2229,N_1885);
and U2699 (N_2699,N_2187,N_1887);
nor U2700 (N_2700,N_2078,N_1805);
and U2701 (N_2701,N_1508,N_1949);
xnor U2702 (N_2702,N_1763,N_2004);
nor U2703 (N_2703,N_2016,N_1525);
and U2704 (N_2704,N_2224,N_2212);
and U2705 (N_2705,N_1933,N_2104);
xor U2706 (N_2706,N_1753,N_1823);
nor U2707 (N_2707,N_2166,N_1723);
nor U2708 (N_2708,N_1989,N_2194);
nand U2709 (N_2709,N_1981,N_1951);
nor U2710 (N_2710,N_1512,N_1941);
nand U2711 (N_2711,N_2164,N_1636);
xnor U2712 (N_2712,N_1705,N_2056);
nor U2713 (N_2713,N_1639,N_1901);
or U2714 (N_2714,N_1985,N_1565);
and U2715 (N_2715,N_2035,N_2173);
nor U2716 (N_2716,N_1711,N_1905);
or U2717 (N_2717,N_1754,N_2235);
xnor U2718 (N_2718,N_2220,N_1697);
xnor U2719 (N_2719,N_2052,N_1974);
xor U2720 (N_2720,N_1941,N_2047);
xor U2721 (N_2721,N_1825,N_1949);
and U2722 (N_2722,N_1863,N_2060);
and U2723 (N_2723,N_2006,N_1933);
nor U2724 (N_2724,N_2076,N_1940);
nand U2725 (N_2725,N_2188,N_1728);
nand U2726 (N_2726,N_1906,N_1973);
nand U2727 (N_2727,N_1594,N_2102);
xnor U2728 (N_2728,N_1794,N_1813);
xor U2729 (N_2729,N_1874,N_1746);
and U2730 (N_2730,N_2169,N_1935);
nand U2731 (N_2731,N_1656,N_2201);
nor U2732 (N_2732,N_1861,N_1828);
nor U2733 (N_2733,N_1706,N_1636);
nor U2734 (N_2734,N_1546,N_1647);
nand U2735 (N_2735,N_1654,N_2209);
nand U2736 (N_2736,N_2216,N_2199);
or U2737 (N_2737,N_1962,N_1521);
nand U2738 (N_2738,N_1588,N_1705);
nand U2739 (N_2739,N_2215,N_2082);
xor U2740 (N_2740,N_1631,N_1718);
nand U2741 (N_2741,N_2142,N_2129);
nor U2742 (N_2742,N_1621,N_1586);
or U2743 (N_2743,N_2236,N_1850);
nand U2744 (N_2744,N_2092,N_1879);
xor U2745 (N_2745,N_1814,N_1966);
nor U2746 (N_2746,N_1571,N_1908);
and U2747 (N_2747,N_1941,N_2148);
or U2748 (N_2748,N_1861,N_1673);
nor U2749 (N_2749,N_2073,N_2215);
nand U2750 (N_2750,N_1931,N_1781);
xor U2751 (N_2751,N_2222,N_1586);
xor U2752 (N_2752,N_1779,N_1581);
nor U2753 (N_2753,N_1774,N_2114);
nor U2754 (N_2754,N_1693,N_2156);
or U2755 (N_2755,N_1954,N_1851);
nor U2756 (N_2756,N_2188,N_2142);
nand U2757 (N_2757,N_2025,N_1780);
xor U2758 (N_2758,N_2032,N_1796);
xor U2759 (N_2759,N_2015,N_2007);
or U2760 (N_2760,N_1511,N_1811);
and U2761 (N_2761,N_1829,N_2096);
or U2762 (N_2762,N_1725,N_1818);
nor U2763 (N_2763,N_2229,N_2047);
or U2764 (N_2764,N_2021,N_1783);
nand U2765 (N_2765,N_1908,N_2221);
nor U2766 (N_2766,N_1903,N_1881);
or U2767 (N_2767,N_1646,N_1819);
xnor U2768 (N_2768,N_1633,N_2051);
xor U2769 (N_2769,N_1623,N_1591);
and U2770 (N_2770,N_1688,N_1886);
nor U2771 (N_2771,N_2067,N_2043);
nor U2772 (N_2772,N_1683,N_1603);
nor U2773 (N_2773,N_1640,N_1662);
xnor U2774 (N_2774,N_2173,N_2107);
or U2775 (N_2775,N_1936,N_1607);
xor U2776 (N_2776,N_1529,N_1678);
nor U2777 (N_2777,N_1754,N_2041);
xor U2778 (N_2778,N_1978,N_1961);
and U2779 (N_2779,N_1864,N_2227);
and U2780 (N_2780,N_1615,N_2020);
and U2781 (N_2781,N_1825,N_1508);
or U2782 (N_2782,N_1727,N_1526);
nor U2783 (N_2783,N_1761,N_1778);
xor U2784 (N_2784,N_1698,N_1971);
or U2785 (N_2785,N_1833,N_2040);
and U2786 (N_2786,N_1802,N_2167);
nor U2787 (N_2787,N_2175,N_1874);
nand U2788 (N_2788,N_1835,N_2117);
nor U2789 (N_2789,N_1846,N_1619);
or U2790 (N_2790,N_2015,N_1723);
nand U2791 (N_2791,N_2083,N_1833);
xor U2792 (N_2792,N_2179,N_2197);
nor U2793 (N_2793,N_1533,N_2073);
or U2794 (N_2794,N_1909,N_1512);
and U2795 (N_2795,N_1887,N_1506);
nand U2796 (N_2796,N_1661,N_1961);
or U2797 (N_2797,N_2109,N_1533);
nand U2798 (N_2798,N_2149,N_1807);
or U2799 (N_2799,N_1907,N_1593);
nor U2800 (N_2800,N_2163,N_1775);
and U2801 (N_2801,N_1792,N_2033);
nand U2802 (N_2802,N_1671,N_1607);
or U2803 (N_2803,N_1688,N_1917);
and U2804 (N_2804,N_2016,N_2065);
nand U2805 (N_2805,N_1726,N_1912);
nand U2806 (N_2806,N_2200,N_1868);
and U2807 (N_2807,N_1986,N_1533);
and U2808 (N_2808,N_2037,N_2186);
or U2809 (N_2809,N_2004,N_1989);
xor U2810 (N_2810,N_2032,N_1847);
or U2811 (N_2811,N_2051,N_1827);
nand U2812 (N_2812,N_2136,N_1749);
nor U2813 (N_2813,N_1805,N_2114);
nand U2814 (N_2814,N_1954,N_2112);
xor U2815 (N_2815,N_1583,N_1816);
and U2816 (N_2816,N_2056,N_1589);
nor U2817 (N_2817,N_2170,N_1968);
and U2818 (N_2818,N_1844,N_2216);
or U2819 (N_2819,N_1574,N_1889);
nand U2820 (N_2820,N_1945,N_2156);
nand U2821 (N_2821,N_1528,N_1562);
and U2822 (N_2822,N_2126,N_1724);
nand U2823 (N_2823,N_1688,N_1540);
xor U2824 (N_2824,N_2236,N_1754);
nand U2825 (N_2825,N_2221,N_2212);
nor U2826 (N_2826,N_2031,N_1858);
and U2827 (N_2827,N_1871,N_1600);
nor U2828 (N_2828,N_2029,N_1726);
and U2829 (N_2829,N_1532,N_1799);
xnor U2830 (N_2830,N_2066,N_2205);
nor U2831 (N_2831,N_1987,N_1617);
nor U2832 (N_2832,N_1979,N_1531);
xor U2833 (N_2833,N_1724,N_1593);
and U2834 (N_2834,N_1662,N_1630);
xor U2835 (N_2835,N_1560,N_2170);
and U2836 (N_2836,N_1610,N_1917);
xor U2837 (N_2837,N_2024,N_2190);
xnor U2838 (N_2838,N_2071,N_1730);
nand U2839 (N_2839,N_2069,N_1539);
nand U2840 (N_2840,N_1575,N_2231);
xnor U2841 (N_2841,N_1824,N_2036);
nor U2842 (N_2842,N_1534,N_1592);
nand U2843 (N_2843,N_2158,N_1529);
nor U2844 (N_2844,N_2123,N_1799);
xnor U2845 (N_2845,N_1757,N_1877);
and U2846 (N_2846,N_2141,N_2191);
and U2847 (N_2847,N_1518,N_1771);
nand U2848 (N_2848,N_2171,N_1598);
or U2849 (N_2849,N_2129,N_1703);
xnor U2850 (N_2850,N_2207,N_2113);
or U2851 (N_2851,N_1789,N_2249);
or U2852 (N_2852,N_1810,N_1691);
nor U2853 (N_2853,N_1736,N_1601);
nand U2854 (N_2854,N_1808,N_1754);
or U2855 (N_2855,N_1774,N_2087);
or U2856 (N_2856,N_1987,N_1609);
xnor U2857 (N_2857,N_1959,N_1837);
nor U2858 (N_2858,N_1669,N_2090);
or U2859 (N_2859,N_2159,N_1549);
and U2860 (N_2860,N_1502,N_1625);
nor U2861 (N_2861,N_1737,N_1893);
and U2862 (N_2862,N_1725,N_2096);
nand U2863 (N_2863,N_1712,N_1702);
and U2864 (N_2864,N_1841,N_1741);
and U2865 (N_2865,N_1582,N_2100);
and U2866 (N_2866,N_1528,N_2197);
xor U2867 (N_2867,N_2231,N_2002);
nor U2868 (N_2868,N_1539,N_1579);
and U2869 (N_2869,N_1539,N_1506);
nand U2870 (N_2870,N_1503,N_1695);
nand U2871 (N_2871,N_2011,N_2133);
nor U2872 (N_2872,N_1851,N_1762);
or U2873 (N_2873,N_1794,N_1921);
or U2874 (N_2874,N_1633,N_2169);
xor U2875 (N_2875,N_1612,N_2224);
xor U2876 (N_2876,N_2077,N_1756);
nor U2877 (N_2877,N_1997,N_1662);
or U2878 (N_2878,N_1712,N_1625);
and U2879 (N_2879,N_2134,N_1507);
nor U2880 (N_2880,N_2014,N_1558);
nor U2881 (N_2881,N_1816,N_1621);
or U2882 (N_2882,N_1856,N_2009);
or U2883 (N_2883,N_1991,N_1659);
nor U2884 (N_2884,N_2227,N_2100);
xor U2885 (N_2885,N_2074,N_2240);
or U2886 (N_2886,N_2054,N_1721);
xor U2887 (N_2887,N_1997,N_1633);
and U2888 (N_2888,N_2056,N_2136);
xnor U2889 (N_2889,N_1700,N_2104);
or U2890 (N_2890,N_1909,N_1508);
xor U2891 (N_2891,N_1669,N_2199);
nor U2892 (N_2892,N_1682,N_1690);
xor U2893 (N_2893,N_1866,N_2102);
xor U2894 (N_2894,N_2188,N_1641);
and U2895 (N_2895,N_2048,N_1615);
or U2896 (N_2896,N_1899,N_1962);
nand U2897 (N_2897,N_2238,N_1565);
xnor U2898 (N_2898,N_1603,N_1838);
nand U2899 (N_2899,N_1595,N_2144);
nand U2900 (N_2900,N_2031,N_1854);
and U2901 (N_2901,N_2206,N_1912);
nor U2902 (N_2902,N_2068,N_1536);
xnor U2903 (N_2903,N_2000,N_1945);
nand U2904 (N_2904,N_2023,N_1853);
xnor U2905 (N_2905,N_1863,N_1560);
nor U2906 (N_2906,N_1982,N_1926);
nor U2907 (N_2907,N_1794,N_2148);
and U2908 (N_2908,N_1567,N_1603);
xor U2909 (N_2909,N_1987,N_1611);
nand U2910 (N_2910,N_1660,N_1694);
nand U2911 (N_2911,N_1702,N_1733);
or U2912 (N_2912,N_1992,N_1830);
or U2913 (N_2913,N_1552,N_2012);
xnor U2914 (N_2914,N_2145,N_2032);
nand U2915 (N_2915,N_1631,N_1705);
and U2916 (N_2916,N_1607,N_1834);
or U2917 (N_2917,N_1712,N_2157);
and U2918 (N_2918,N_1826,N_1815);
and U2919 (N_2919,N_1728,N_1795);
xor U2920 (N_2920,N_2072,N_1837);
and U2921 (N_2921,N_1856,N_1612);
xor U2922 (N_2922,N_1512,N_2111);
nor U2923 (N_2923,N_1576,N_1806);
xor U2924 (N_2924,N_1976,N_1743);
and U2925 (N_2925,N_1979,N_2003);
xnor U2926 (N_2926,N_2109,N_2093);
and U2927 (N_2927,N_1588,N_1824);
and U2928 (N_2928,N_1952,N_1702);
nand U2929 (N_2929,N_1907,N_2010);
xor U2930 (N_2930,N_2052,N_2187);
nor U2931 (N_2931,N_1761,N_2210);
nand U2932 (N_2932,N_2063,N_2025);
or U2933 (N_2933,N_1908,N_2004);
nor U2934 (N_2934,N_2144,N_2094);
and U2935 (N_2935,N_1545,N_1982);
or U2936 (N_2936,N_1981,N_1651);
nor U2937 (N_2937,N_2103,N_2015);
nand U2938 (N_2938,N_2144,N_1702);
nor U2939 (N_2939,N_1536,N_1988);
or U2940 (N_2940,N_2214,N_2249);
xor U2941 (N_2941,N_1909,N_2177);
or U2942 (N_2942,N_2165,N_1675);
xor U2943 (N_2943,N_1711,N_2127);
and U2944 (N_2944,N_2128,N_1705);
nand U2945 (N_2945,N_1832,N_1928);
or U2946 (N_2946,N_1574,N_1648);
xnor U2947 (N_2947,N_2118,N_1770);
and U2948 (N_2948,N_1592,N_1823);
and U2949 (N_2949,N_1826,N_1693);
or U2950 (N_2950,N_2189,N_1857);
xor U2951 (N_2951,N_1643,N_1743);
and U2952 (N_2952,N_1518,N_2210);
or U2953 (N_2953,N_1529,N_2143);
and U2954 (N_2954,N_2118,N_1798);
xnor U2955 (N_2955,N_1502,N_1980);
and U2956 (N_2956,N_2068,N_2054);
xor U2957 (N_2957,N_1627,N_1901);
xnor U2958 (N_2958,N_1908,N_1560);
nor U2959 (N_2959,N_1855,N_1572);
nand U2960 (N_2960,N_1650,N_1867);
and U2961 (N_2961,N_2167,N_1989);
nand U2962 (N_2962,N_1781,N_2056);
and U2963 (N_2963,N_2167,N_2173);
nor U2964 (N_2964,N_1807,N_1895);
or U2965 (N_2965,N_1837,N_1868);
nand U2966 (N_2966,N_1568,N_1861);
or U2967 (N_2967,N_1714,N_1569);
or U2968 (N_2968,N_1639,N_2077);
and U2969 (N_2969,N_2190,N_2091);
and U2970 (N_2970,N_2135,N_2136);
or U2971 (N_2971,N_1623,N_1707);
or U2972 (N_2972,N_2075,N_1851);
xor U2973 (N_2973,N_1806,N_1902);
xnor U2974 (N_2974,N_2170,N_2136);
xnor U2975 (N_2975,N_2152,N_1722);
xor U2976 (N_2976,N_2204,N_2169);
nor U2977 (N_2977,N_2215,N_1925);
or U2978 (N_2978,N_1756,N_2062);
xor U2979 (N_2979,N_1653,N_1878);
xor U2980 (N_2980,N_2003,N_2123);
nand U2981 (N_2981,N_2231,N_2220);
nor U2982 (N_2982,N_2114,N_1589);
nand U2983 (N_2983,N_2248,N_2134);
nand U2984 (N_2984,N_1628,N_1936);
nand U2985 (N_2985,N_1919,N_1585);
or U2986 (N_2986,N_2059,N_1746);
nand U2987 (N_2987,N_1884,N_2058);
nor U2988 (N_2988,N_1635,N_1613);
xor U2989 (N_2989,N_1514,N_1964);
nor U2990 (N_2990,N_2101,N_1770);
nor U2991 (N_2991,N_2203,N_1946);
xor U2992 (N_2992,N_2021,N_1752);
nand U2993 (N_2993,N_2197,N_2171);
nand U2994 (N_2994,N_2017,N_1838);
nor U2995 (N_2995,N_1831,N_1813);
nor U2996 (N_2996,N_1515,N_1916);
and U2997 (N_2997,N_1774,N_2012);
xor U2998 (N_2998,N_1585,N_1730);
xnor U2999 (N_2999,N_1858,N_2105);
nor UO_0 (O_0,N_2685,N_2809);
xor UO_1 (O_1,N_2480,N_2855);
and UO_2 (O_2,N_2278,N_2386);
nor UO_3 (O_3,N_2727,N_2394);
or UO_4 (O_4,N_2811,N_2526);
nor UO_5 (O_5,N_2385,N_2790);
xnor UO_6 (O_6,N_2307,N_2618);
or UO_7 (O_7,N_2766,N_2761);
nor UO_8 (O_8,N_2688,N_2428);
xor UO_9 (O_9,N_2446,N_2515);
and UO_10 (O_10,N_2641,N_2689);
or UO_11 (O_11,N_2315,N_2771);
xor UO_12 (O_12,N_2499,N_2258);
and UO_13 (O_13,N_2910,N_2354);
nand UO_14 (O_14,N_2457,N_2464);
or UO_15 (O_15,N_2624,N_2617);
and UO_16 (O_16,N_2778,N_2709);
xor UO_17 (O_17,N_2593,N_2942);
and UO_18 (O_18,N_2266,N_2741);
nand UO_19 (O_19,N_2305,N_2352);
nand UO_20 (O_20,N_2740,N_2976);
nand UO_21 (O_21,N_2667,N_2532);
or UO_22 (O_22,N_2605,N_2523);
or UO_23 (O_23,N_2857,N_2481);
and UO_24 (O_24,N_2886,N_2812);
xnor UO_25 (O_25,N_2989,N_2412);
nor UO_26 (O_26,N_2748,N_2531);
nor UO_27 (O_27,N_2253,N_2670);
nor UO_28 (O_28,N_2834,N_2721);
nand UO_29 (O_29,N_2953,N_2729);
nand UO_30 (O_30,N_2340,N_2776);
xor UO_31 (O_31,N_2427,N_2666);
and UO_32 (O_32,N_2567,N_2978);
and UO_33 (O_33,N_2357,N_2272);
xor UO_34 (O_34,N_2369,N_2918);
nand UO_35 (O_35,N_2580,N_2676);
and UO_36 (O_36,N_2877,N_2609);
xor UO_37 (O_37,N_2908,N_2804);
nor UO_38 (O_38,N_2629,N_2512);
or UO_39 (O_39,N_2549,N_2797);
xor UO_40 (O_40,N_2536,N_2979);
xnor UO_41 (O_41,N_2551,N_2830);
xnor UO_42 (O_42,N_2682,N_2255);
or UO_43 (O_43,N_2880,N_2840);
and UO_44 (O_44,N_2905,N_2632);
or UO_45 (O_45,N_2575,N_2296);
nor UO_46 (O_46,N_2756,N_2985);
nand UO_47 (O_47,N_2610,N_2252);
nand UO_48 (O_48,N_2450,N_2290);
nor UO_49 (O_49,N_2644,N_2510);
or UO_50 (O_50,N_2966,N_2940);
or UO_51 (O_51,N_2430,N_2681);
or UO_52 (O_52,N_2795,N_2260);
xor UO_53 (O_53,N_2562,N_2263);
nor UO_54 (O_54,N_2365,N_2922);
or UO_55 (O_55,N_2954,N_2298);
or UO_56 (O_56,N_2683,N_2715);
xnor UO_57 (O_57,N_2926,N_2406);
nor UO_58 (O_58,N_2498,N_2946);
or UO_59 (O_59,N_2903,N_2917);
xor UO_60 (O_60,N_2588,N_2483);
xnor UO_61 (O_61,N_2441,N_2547);
or UO_62 (O_62,N_2702,N_2294);
and UO_63 (O_63,N_2583,N_2770);
nand UO_64 (O_64,N_2813,N_2881);
xor UO_65 (O_65,N_2915,N_2935);
and UO_66 (O_66,N_2755,N_2521);
or UO_67 (O_67,N_2322,N_2858);
nand UO_68 (O_68,N_2424,N_2691);
nor UO_69 (O_69,N_2321,N_2820);
nor UO_70 (O_70,N_2458,N_2661);
nand UO_71 (O_71,N_2492,N_2387);
and UO_72 (O_72,N_2995,N_2724);
or UO_73 (O_73,N_2972,N_2791);
or UO_74 (O_74,N_2655,N_2752);
xor UO_75 (O_75,N_2494,N_2675);
and UO_76 (O_76,N_2569,N_2348);
nand UO_77 (O_77,N_2587,N_2389);
and UO_78 (O_78,N_2726,N_2653);
or UO_79 (O_79,N_2529,N_2448);
or UO_80 (O_80,N_2873,N_2939);
or UO_81 (O_81,N_2723,N_2975);
nor UO_82 (O_82,N_2714,N_2734);
or UO_83 (O_83,N_2274,N_2982);
nand UO_84 (O_84,N_2410,N_2535);
nand UO_85 (O_85,N_2534,N_2784);
xor UO_86 (O_86,N_2713,N_2779);
xor UO_87 (O_87,N_2454,N_2506);
nor UO_88 (O_88,N_2563,N_2422);
and UO_89 (O_89,N_2388,N_2974);
or UO_90 (O_90,N_2678,N_2810);
and UO_91 (O_91,N_2692,N_2868);
nor UO_92 (O_92,N_2434,N_2620);
or UO_93 (O_93,N_2671,N_2827);
xnor UO_94 (O_94,N_2656,N_2347);
xnor UO_95 (O_95,N_2329,N_2901);
xnor UO_96 (O_96,N_2833,N_2559);
xor UO_97 (O_97,N_2735,N_2798);
and UO_98 (O_98,N_2495,N_2436);
xnor UO_99 (O_99,N_2651,N_2311);
and UO_100 (O_100,N_2851,N_2381);
nor UO_101 (O_101,N_2493,N_2867);
nand UO_102 (O_102,N_2687,N_2951);
xnor UO_103 (O_103,N_2716,N_2533);
nor UO_104 (O_104,N_2647,N_2376);
nor UO_105 (O_105,N_2906,N_2317);
nand UO_106 (O_106,N_2279,N_2608);
nor UO_107 (O_107,N_2442,N_2539);
or UO_108 (O_108,N_2413,N_2701);
or UO_109 (O_109,N_2527,N_2557);
nand UO_110 (O_110,N_2635,N_2368);
xor UO_111 (O_111,N_2850,N_2631);
or UO_112 (O_112,N_2358,N_2423);
xor UO_113 (O_113,N_2911,N_2316);
xor UO_114 (O_114,N_2808,N_2821);
and UO_115 (O_115,N_2379,N_2262);
and UO_116 (O_116,N_2383,N_2849);
xor UO_117 (O_117,N_2257,N_2875);
nand UO_118 (O_118,N_2265,N_2615);
and UO_119 (O_119,N_2775,N_2805);
nand UO_120 (O_120,N_2513,N_2612);
or UO_121 (O_121,N_2957,N_2479);
nor UO_122 (O_122,N_2576,N_2505);
nand UO_123 (O_123,N_2443,N_2623);
nor UO_124 (O_124,N_2919,N_2544);
nand UO_125 (O_125,N_2967,N_2891);
nor UO_126 (O_126,N_2718,N_2930);
nand UO_127 (O_127,N_2362,N_2611);
nand UO_128 (O_128,N_2301,N_2327);
nand UO_129 (O_129,N_2338,N_2598);
nor UO_130 (O_130,N_2658,N_2283);
xnor UO_131 (O_131,N_2669,N_2330);
or UO_132 (O_132,N_2254,N_2486);
or UO_133 (O_133,N_2607,N_2997);
nor UO_134 (O_134,N_2275,N_2318);
nand UO_135 (O_135,N_2261,N_2816);
nand UO_136 (O_136,N_2990,N_2277);
nor UO_137 (O_137,N_2405,N_2497);
nor UO_138 (O_138,N_2916,N_2956);
and UO_139 (O_139,N_2984,N_2633);
nor UO_140 (O_140,N_2509,N_2473);
or UO_141 (O_141,N_2859,N_2308);
or UO_142 (O_142,N_2794,N_2627);
nor UO_143 (O_143,N_2304,N_2963);
xor UO_144 (O_144,N_2426,N_2626);
nor UO_145 (O_145,N_2991,N_2973);
nand UO_146 (O_146,N_2416,N_2664);
xor UO_147 (O_147,N_2927,N_2898);
or UO_148 (O_148,N_2584,N_2904);
nand UO_149 (O_149,N_2342,N_2380);
nor UO_150 (O_150,N_2907,N_2392);
xor UO_151 (O_151,N_2297,N_2802);
nor UO_152 (O_152,N_2838,N_2731);
xor UO_153 (O_153,N_2414,N_2391);
nand UO_154 (O_154,N_2780,N_2879);
or UO_155 (O_155,N_2920,N_2993);
and UO_156 (O_156,N_2981,N_2478);
or UO_157 (O_157,N_2417,N_2606);
and UO_158 (O_158,N_2467,N_2654);
or UO_159 (O_159,N_2351,N_2518);
nand UO_160 (O_160,N_2968,N_2408);
nor UO_161 (O_161,N_2648,N_2936);
or UO_162 (O_162,N_2396,N_2461);
nor UO_163 (O_163,N_2789,N_2807);
and UO_164 (O_164,N_2883,N_2597);
and UO_165 (O_165,N_2772,N_2370);
nand UO_166 (O_166,N_2395,N_2604);
or UO_167 (O_167,N_2839,N_2335);
xnor UO_168 (O_168,N_2703,N_2896);
xor UO_169 (O_169,N_2646,N_2568);
nand UO_170 (O_170,N_2961,N_2738);
nor UO_171 (O_171,N_2359,N_2679);
or UO_172 (O_172,N_2720,N_2519);
nand UO_173 (O_173,N_2814,N_2705);
xnor UO_174 (O_174,N_2281,N_2842);
and UO_175 (O_175,N_2996,N_2466);
or UO_176 (O_176,N_2508,N_2432);
and UO_177 (O_177,N_2783,N_2323);
xor UO_178 (O_178,N_2398,N_2694);
or UO_179 (O_179,N_2642,N_2640);
and UO_180 (O_180,N_2937,N_2476);
xor UO_181 (O_181,N_2962,N_2882);
xnor UO_182 (O_182,N_2938,N_2751);
or UO_183 (O_183,N_2449,N_2540);
nor UO_184 (O_184,N_2339,N_2300);
xor UO_185 (O_185,N_2952,N_2522);
and UO_186 (O_186,N_2295,N_2420);
xor UO_187 (O_187,N_2969,N_2933);
nor UO_188 (O_188,N_2674,N_2332);
nor UO_189 (O_189,N_2582,N_2276);
xor UO_190 (O_190,N_2453,N_2970);
nand UO_191 (O_191,N_2268,N_2749);
xor UO_192 (O_192,N_2292,N_2707);
xnor UO_193 (O_193,N_2825,N_2831);
nor UO_194 (O_194,N_2538,N_2367);
and UO_195 (O_195,N_2556,N_2287);
and UO_196 (O_196,N_2586,N_2421);
nor UO_197 (O_197,N_2866,N_2595);
xor UO_198 (O_198,N_2754,N_2841);
nor UO_199 (O_199,N_2484,N_2665);
xor UO_200 (O_200,N_2913,N_2774);
nand UO_201 (O_201,N_2474,N_2490);
nand UO_202 (O_202,N_2662,N_2353);
and UO_203 (O_203,N_2429,N_2819);
nor UO_204 (O_204,N_2284,N_2697);
xor UO_205 (O_205,N_2573,N_2343);
nor UO_206 (O_206,N_2485,N_2334);
nor UO_207 (O_207,N_2561,N_2302);
or UO_208 (O_208,N_2267,N_2328);
or UO_209 (O_209,N_2832,N_2259);
xor UO_210 (O_210,N_2264,N_2433);
nor UO_211 (O_211,N_2570,N_2344);
and UO_212 (O_212,N_2826,N_2759);
xnor UO_213 (O_213,N_2899,N_2271);
or UO_214 (O_214,N_2585,N_2852);
xnor UO_215 (O_215,N_2792,N_2680);
nand UO_216 (O_216,N_2693,N_2829);
and UO_217 (O_217,N_2520,N_2965);
or UO_218 (O_218,N_2350,N_2463);
xor UO_219 (O_219,N_2372,N_2553);
nor UO_220 (O_220,N_2845,N_2313);
and UO_221 (O_221,N_2944,N_2730);
nand UO_222 (O_222,N_2541,N_2945);
or UO_223 (O_223,N_2710,N_2923);
xor UO_224 (O_224,N_2530,N_2711);
and UO_225 (O_225,N_2411,N_2765);
or UO_226 (O_226,N_2864,N_2601);
nand UO_227 (O_227,N_2803,N_2817);
or UO_228 (O_228,N_2337,N_2579);
nand UO_229 (O_229,N_2487,N_2760);
nor UO_230 (O_230,N_2890,N_2309);
nor UO_231 (O_231,N_2793,N_2986);
nor UO_232 (O_232,N_2998,N_2762);
and UO_233 (O_233,N_2571,N_2844);
xnor UO_234 (O_234,N_2614,N_2737);
nor UO_235 (O_235,N_2673,N_2282);
nor UO_236 (O_236,N_2708,N_2404);
or UO_237 (O_237,N_2577,N_2397);
nor UO_238 (O_238,N_2941,N_2346);
nor UO_239 (O_239,N_2451,N_2955);
and UO_240 (O_240,N_2949,N_2796);
xor UO_241 (O_241,N_2336,N_2285);
or UO_242 (O_242,N_2932,N_2743);
xor UO_243 (O_243,N_2786,N_2848);
xnor UO_244 (O_244,N_2983,N_2399);
or UO_245 (O_245,N_2602,N_2757);
nor UO_246 (O_246,N_2482,N_2739);
nand UO_247 (O_247,N_2860,N_2865);
xnor UO_248 (O_248,N_2668,N_2725);
nand UO_249 (O_249,N_2660,N_2489);
nand UO_250 (O_250,N_2280,N_2550);
xnor UO_251 (O_251,N_2528,N_2500);
or UO_252 (O_252,N_2468,N_2377);
nand UO_253 (O_253,N_2785,N_2672);
nor UO_254 (O_254,N_2872,N_2360);
nor UO_255 (O_255,N_2431,N_2843);
or UO_256 (O_256,N_2750,N_2987);
nand UO_257 (O_257,N_2341,N_2948);
nand UO_258 (O_258,N_2472,N_2909);
or UO_259 (O_259,N_2289,N_2924);
or UO_260 (O_260,N_2603,N_2856);
nor UO_261 (O_261,N_2270,N_2502);
xnor UO_262 (O_262,N_2578,N_2470);
nand UO_263 (O_263,N_2677,N_2628);
nor UO_264 (O_264,N_2950,N_2592);
nand UO_265 (O_265,N_2828,N_2299);
or UO_266 (O_266,N_2921,N_2686);
or UO_267 (O_267,N_2732,N_2992);
xor UO_268 (O_268,N_2884,N_2736);
and UO_269 (O_269,N_2496,N_2545);
and UO_270 (O_270,N_2980,N_2320);
or UO_271 (O_271,N_2349,N_2787);
xnor UO_272 (O_272,N_2554,N_2616);
and UO_273 (O_273,N_2768,N_2524);
nand UO_274 (O_274,N_2690,N_2929);
xor UO_275 (O_275,N_2488,N_2581);
xnor UO_276 (O_276,N_2650,N_2250);
nor UO_277 (O_277,N_2501,N_2684);
or UO_278 (O_278,N_2878,N_2897);
nor UO_279 (O_279,N_2887,N_2543);
nor UO_280 (O_280,N_2902,N_2471);
or UO_281 (O_281,N_2364,N_2425);
and UO_282 (O_282,N_2799,N_2815);
or UO_283 (O_283,N_2574,N_2621);
and UO_284 (O_284,N_2636,N_2712);
xnor UO_285 (O_285,N_2767,N_2822);
nor UO_286 (O_286,N_2371,N_2645);
xnor UO_287 (O_287,N_2455,N_2537);
xor UO_288 (O_288,N_2800,N_2475);
xor UO_289 (O_289,N_2853,N_2409);
xnor UO_290 (O_290,N_2744,N_2477);
or UO_291 (O_291,N_2900,N_2415);
and UO_292 (O_292,N_2630,N_2312);
or UO_293 (O_293,N_2456,N_2333);
and UO_294 (O_294,N_2638,N_2491);
nand UO_295 (O_295,N_2959,N_2625);
xor UO_296 (O_296,N_2912,N_2600);
or UO_297 (O_297,N_2773,N_2303);
and UO_298 (O_298,N_2781,N_2874);
nor UO_299 (O_299,N_2373,N_2728);
and UO_300 (O_300,N_2407,N_2733);
nand UO_301 (O_301,N_2764,N_2704);
and UO_302 (O_302,N_2291,N_2862);
and UO_303 (O_303,N_2637,N_2652);
nor UO_304 (O_304,N_2552,N_2861);
nand UO_305 (O_305,N_2403,N_2769);
or UO_306 (O_306,N_2892,N_2869);
or UO_307 (O_307,N_2746,N_2445);
or UO_308 (O_308,N_2657,N_2871);
and UO_309 (O_309,N_2719,N_2314);
nor UO_310 (O_310,N_2435,N_2469);
or UO_311 (O_311,N_2440,N_2504);
xnor UO_312 (O_312,N_2639,N_2696);
nand UO_313 (O_313,N_2459,N_2251);
nor UO_314 (O_314,N_2854,N_2273);
nand UO_315 (O_315,N_2465,N_2971);
xnor UO_316 (O_316,N_2402,N_2400);
xnor UO_317 (O_317,N_2511,N_2447);
nand UO_318 (O_318,N_2836,N_2777);
nand UO_319 (O_319,N_2462,N_2325);
nor UO_320 (O_320,N_2516,N_2698);
nand UO_321 (O_321,N_2823,N_2566);
or UO_322 (O_322,N_2548,N_2288);
nor UO_323 (O_323,N_2999,N_2460);
xnor UO_324 (O_324,N_2925,N_2564);
nand UO_325 (O_325,N_2885,N_2594);
nor UO_326 (O_326,N_2835,N_2356);
nand UO_327 (O_327,N_2437,N_2525);
nor UO_328 (O_328,N_2914,N_2782);
or UO_329 (O_329,N_2401,N_2363);
xor UO_330 (O_330,N_2293,N_2977);
or UO_331 (O_331,N_2390,N_2355);
and UO_332 (O_332,N_2634,N_2560);
nand UO_333 (O_333,N_2326,N_2555);
xor UO_334 (O_334,N_2507,N_2452);
xnor UO_335 (O_335,N_2663,N_2888);
and UO_336 (O_336,N_2366,N_2958);
and UO_337 (O_337,N_2310,N_2863);
or UO_338 (O_338,N_2806,N_2947);
nor UO_339 (O_339,N_2894,N_2444);
xnor UO_340 (O_340,N_2438,N_2895);
xor UO_341 (O_341,N_2382,N_2599);
xor UO_342 (O_342,N_2384,N_2643);
xnor UO_343 (O_343,N_2622,N_2818);
xor UO_344 (O_344,N_2876,N_2659);
or UO_345 (O_345,N_2619,N_2590);
and UO_346 (O_346,N_2717,N_2994);
and UO_347 (O_347,N_2589,N_2699);
nor UO_348 (O_348,N_2591,N_2801);
or UO_349 (O_349,N_2565,N_2546);
or UO_350 (O_350,N_2722,N_2747);
or UO_351 (O_351,N_2256,N_2788);
and UO_352 (O_352,N_2988,N_2331);
xor UO_353 (O_353,N_2753,N_2319);
nand UO_354 (O_354,N_2378,N_2286);
xnor UO_355 (O_355,N_2763,N_2613);
xnor UO_356 (O_356,N_2419,N_2517);
nand UO_357 (O_357,N_2306,N_2893);
xnor UO_358 (O_358,N_2846,N_2324);
and UO_359 (O_359,N_2745,N_2928);
xor UO_360 (O_360,N_2960,N_2649);
xnor UO_361 (O_361,N_2542,N_2572);
nor UO_362 (O_362,N_2758,N_2889);
and UO_363 (O_363,N_2931,N_2706);
and UO_364 (O_364,N_2700,N_2374);
nor UO_365 (O_365,N_2514,N_2361);
or UO_366 (O_366,N_2964,N_2269);
nor UO_367 (O_367,N_2870,N_2393);
and UO_368 (O_368,N_2558,N_2439);
nand UO_369 (O_369,N_2742,N_2837);
xnor UO_370 (O_370,N_2847,N_2824);
and UO_371 (O_371,N_2345,N_2418);
nand UO_372 (O_372,N_2503,N_2934);
and UO_373 (O_373,N_2596,N_2943);
nand UO_374 (O_374,N_2375,N_2695);
or UO_375 (O_375,N_2727,N_2640);
xnor UO_376 (O_376,N_2913,N_2402);
nand UO_377 (O_377,N_2533,N_2467);
or UO_378 (O_378,N_2437,N_2516);
nor UO_379 (O_379,N_2551,N_2363);
nor UO_380 (O_380,N_2298,N_2308);
nor UO_381 (O_381,N_2732,N_2565);
nor UO_382 (O_382,N_2463,N_2959);
nand UO_383 (O_383,N_2594,N_2973);
xnor UO_384 (O_384,N_2564,N_2549);
nor UO_385 (O_385,N_2755,N_2931);
nor UO_386 (O_386,N_2783,N_2276);
xnor UO_387 (O_387,N_2832,N_2348);
xor UO_388 (O_388,N_2960,N_2271);
nor UO_389 (O_389,N_2667,N_2824);
nand UO_390 (O_390,N_2478,N_2665);
or UO_391 (O_391,N_2342,N_2385);
xor UO_392 (O_392,N_2642,N_2289);
xnor UO_393 (O_393,N_2713,N_2325);
xor UO_394 (O_394,N_2568,N_2578);
and UO_395 (O_395,N_2965,N_2275);
xnor UO_396 (O_396,N_2701,N_2615);
nor UO_397 (O_397,N_2868,N_2650);
nor UO_398 (O_398,N_2949,N_2543);
or UO_399 (O_399,N_2775,N_2984);
nand UO_400 (O_400,N_2425,N_2591);
xor UO_401 (O_401,N_2730,N_2258);
nor UO_402 (O_402,N_2844,N_2523);
and UO_403 (O_403,N_2582,N_2318);
or UO_404 (O_404,N_2550,N_2797);
nand UO_405 (O_405,N_2929,N_2977);
nand UO_406 (O_406,N_2450,N_2272);
xor UO_407 (O_407,N_2643,N_2650);
xor UO_408 (O_408,N_2893,N_2770);
and UO_409 (O_409,N_2507,N_2839);
nor UO_410 (O_410,N_2745,N_2897);
nand UO_411 (O_411,N_2283,N_2264);
or UO_412 (O_412,N_2335,N_2334);
xor UO_413 (O_413,N_2260,N_2882);
nor UO_414 (O_414,N_2638,N_2844);
nand UO_415 (O_415,N_2281,N_2445);
or UO_416 (O_416,N_2924,N_2379);
xnor UO_417 (O_417,N_2315,N_2775);
and UO_418 (O_418,N_2327,N_2755);
or UO_419 (O_419,N_2949,N_2995);
or UO_420 (O_420,N_2350,N_2582);
nand UO_421 (O_421,N_2665,N_2992);
or UO_422 (O_422,N_2965,N_2287);
nor UO_423 (O_423,N_2961,N_2623);
and UO_424 (O_424,N_2391,N_2369);
xor UO_425 (O_425,N_2822,N_2546);
xor UO_426 (O_426,N_2814,N_2260);
nand UO_427 (O_427,N_2885,N_2434);
and UO_428 (O_428,N_2661,N_2654);
and UO_429 (O_429,N_2981,N_2377);
nand UO_430 (O_430,N_2962,N_2281);
and UO_431 (O_431,N_2794,N_2743);
and UO_432 (O_432,N_2726,N_2612);
xor UO_433 (O_433,N_2541,N_2581);
and UO_434 (O_434,N_2466,N_2503);
or UO_435 (O_435,N_2978,N_2702);
xor UO_436 (O_436,N_2361,N_2430);
nor UO_437 (O_437,N_2901,N_2502);
nand UO_438 (O_438,N_2959,N_2594);
and UO_439 (O_439,N_2693,N_2404);
or UO_440 (O_440,N_2370,N_2341);
or UO_441 (O_441,N_2925,N_2700);
and UO_442 (O_442,N_2845,N_2659);
nor UO_443 (O_443,N_2465,N_2816);
or UO_444 (O_444,N_2870,N_2850);
or UO_445 (O_445,N_2809,N_2936);
or UO_446 (O_446,N_2371,N_2980);
nor UO_447 (O_447,N_2313,N_2314);
or UO_448 (O_448,N_2594,N_2500);
xnor UO_449 (O_449,N_2580,N_2648);
nor UO_450 (O_450,N_2797,N_2773);
nand UO_451 (O_451,N_2627,N_2251);
nor UO_452 (O_452,N_2708,N_2552);
and UO_453 (O_453,N_2545,N_2692);
or UO_454 (O_454,N_2981,N_2551);
and UO_455 (O_455,N_2705,N_2658);
nand UO_456 (O_456,N_2321,N_2477);
nand UO_457 (O_457,N_2915,N_2270);
nor UO_458 (O_458,N_2760,N_2684);
nor UO_459 (O_459,N_2790,N_2477);
nor UO_460 (O_460,N_2642,N_2379);
nor UO_461 (O_461,N_2444,N_2880);
nand UO_462 (O_462,N_2494,N_2391);
and UO_463 (O_463,N_2874,N_2379);
xnor UO_464 (O_464,N_2868,N_2309);
and UO_465 (O_465,N_2275,N_2401);
xnor UO_466 (O_466,N_2946,N_2780);
xnor UO_467 (O_467,N_2746,N_2971);
or UO_468 (O_468,N_2334,N_2250);
and UO_469 (O_469,N_2612,N_2540);
nor UO_470 (O_470,N_2440,N_2953);
nor UO_471 (O_471,N_2496,N_2267);
and UO_472 (O_472,N_2513,N_2369);
nand UO_473 (O_473,N_2969,N_2876);
nor UO_474 (O_474,N_2442,N_2944);
or UO_475 (O_475,N_2805,N_2364);
or UO_476 (O_476,N_2864,N_2296);
nor UO_477 (O_477,N_2830,N_2268);
nor UO_478 (O_478,N_2675,N_2746);
nor UO_479 (O_479,N_2553,N_2810);
xor UO_480 (O_480,N_2299,N_2790);
xor UO_481 (O_481,N_2704,N_2998);
nor UO_482 (O_482,N_2602,N_2305);
xor UO_483 (O_483,N_2397,N_2398);
nor UO_484 (O_484,N_2520,N_2952);
and UO_485 (O_485,N_2500,N_2619);
xnor UO_486 (O_486,N_2974,N_2419);
or UO_487 (O_487,N_2398,N_2305);
nor UO_488 (O_488,N_2824,N_2991);
xor UO_489 (O_489,N_2485,N_2898);
nand UO_490 (O_490,N_2799,N_2402);
and UO_491 (O_491,N_2590,N_2366);
nand UO_492 (O_492,N_2373,N_2470);
or UO_493 (O_493,N_2933,N_2774);
or UO_494 (O_494,N_2349,N_2713);
nand UO_495 (O_495,N_2834,N_2475);
nand UO_496 (O_496,N_2445,N_2976);
and UO_497 (O_497,N_2411,N_2390);
nor UO_498 (O_498,N_2288,N_2316);
nand UO_499 (O_499,N_2773,N_2832);
endmodule