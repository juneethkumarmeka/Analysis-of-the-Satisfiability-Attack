module basic_1500_15000_2000_20_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_1327,In_502);
xor U1 (N_1,In_89,In_772);
and U2 (N_2,In_514,In_1320);
nand U3 (N_3,In_1368,In_1393);
nand U4 (N_4,In_983,In_474);
nor U5 (N_5,In_520,In_367);
nor U6 (N_6,In_62,In_789);
nand U7 (N_7,In_820,In_534);
or U8 (N_8,In_700,In_477);
nor U9 (N_9,In_480,In_1353);
and U10 (N_10,In_1418,In_1406);
nand U11 (N_11,In_3,In_855);
nand U12 (N_12,In_1111,In_766);
and U13 (N_13,In_1232,In_1275);
or U14 (N_14,In_90,In_1147);
or U15 (N_15,In_1400,In_59);
or U16 (N_16,In_438,In_719);
and U17 (N_17,In_954,In_452);
or U18 (N_18,In_408,In_93);
nand U19 (N_19,In_291,In_1105);
or U20 (N_20,In_1284,In_724);
nand U21 (N_21,In_1499,In_49);
and U22 (N_22,In_875,In_821);
nor U23 (N_23,In_1397,In_911);
nand U24 (N_24,In_336,In_196);
xor U25 (N_25,In_453,In_808);
nor U26 (N_26,In_481,In_551);
nor U27 (N_27,In_380,In_276);
and U28 (N_28,In_646,In_638);
or U29 (N_29,In_1340,In_1045);
xor U30 (N_30,In_223,In_629);
and U31 (N_31,In_245,In_234);
nand U32 (N_32,In_591,In_91);
nand U33 (N_33,In_240,In_1040);
or U34 (N_34,In_1480,In_1276);
xor U35 (N_35,In_1092,In_1435);
or U36 (N_36,In_197,In_1362);
nor U37 (N_37,In_280,In_423);
or U38 (N_38,In_1159,In_1234);
and U39 (N_39,In_1237,In_230);
xnor U40 (N_40,In_921,In_1321);
nand U41 (N_41,In_256,In_834);
and U42 (N_42,In_773,In_347);
or U43 (N_43,In_258,In_1027);
nor U44 (N_44,In_787,In_1255);
nand U45 (N_45,In_856,In_265);
nand U46 (N_46,In_546,In_560);
or U47 (N_47,In_684,In_1077);
or U48 (N_48,In_139,In_137);
xnor U49 (N_49,In_956,In_450);
xor U50 (N_50,In_315,In_1174);
nor U51 (N_51,In_266,In_1495);
and U52 (N_52,In_774,In_1460);
or U53 (N_53,In_1361,In_1223);
nand U54 (N_54,In_1248,In_470);
xnor U55 (N_55,In_817,In_704);
nand U56 (N_56,In_55,In_1145);
or U57 (N_57,In_729,In_15);
or U58 (N_58,In_640,In_1048);
nand U59 (N_59,In_394,In_30);
or U60 (N_60,In_877,In_779);
nand U61 (N_61,In_1380,In_199);
or U62 (N_62,In_525,In_594);
or U63 (N_63,In_34,In_878);
nand U64 (N_64,In_516,In_239);
or U65 (N_65,In_1347,In_379);
or U66 (N_66,In_861,In_651);
or U67 (N_67,In_893,In_695);
nand U68 (N_68,In_166,In_575);
nand U69 (N_69,In_1462,In_402);
xor U70 (N_70,In_513,In_28);
nand U71 (N_71,In_974,In_1150);
xor U72 (N_72,In_688,In_1099);
and U73 (N_73,In_332,In_792);
nand U74 (N_74,In_709,In_717);
or U75 (N_75,In_851,In_167);
nor U76 (N_76,In_1337,In_102);
nor U77 (N_77,In_1496,In_707);
or U78 (N_78,In_1371,In_896);
nand U79 (N_79,In_866,In_1485);
and U80 (N_80,In_88,In_1124);
and U81 (N_81,In_1262,In_469);
nand U82 (N_82,In_232,In_178);
nor U83 (N_83,In_1486,In_1442);
or U84 (N_84,In_1475,In_115);
nand U85 (N_85,In_107,In_917);
or U86 (N_86,In_720,In_894);
and U87 (N_87,In_1446,In_565);
nor U88 (N_88,In_1383,In_271);
and U89 (N_89,In_282,In_1333);
nand U90 (N_90,In_791,In_955);
nand U91 (N_91,In_657,In_543);
or U92 (N_92,In_1372,In_82);
nor U93 (N_93,In_1043,In_1144);
or U94 (N_94,In_136,In_716);
or U95 (N_95,In_171,In_811);
or U96 (N_96,In_235,In_564);
nand U97 (N_97,In_1296,In_1018);
nor U98 (N_98,In_882,In_1363);
nor U99 (N_99,In_128,In_73);
or U100 (N_100,In_1443,In_975);
nand U101 (N_101,In_1113,In_242);
nand U102 (N_102,In_970,In_1295);
nor U103 (N_103,In_1009,In_562);
nor U104 (N_104,In_1025,In_1414);
nand U105 (N_105,In_506,In_1019);
or U106 (N_106,In_297,In_1430);
nor U107 (N_107,In_530,In_623);
and U108 (N_108,In_1004,In_1120);
or U109 (N_109,In_494,In_505);
nand U110 (N_110,In_53,In_1434);
nand U111 (N_111,In_935,In_1230);
nor U112 (N_112,In_1125,In_961);
xor U113 (N_113,In_1089,In_846);
or U114 (N_114,In_85,In_1313);
and U115 (N_115,In_289,In_236);
and U116 (N_116,In_883,In_781);
nor U117 (N_117,In_827,In_1044);
nor U118 (N_118,In_805,In_76);
xor U119 (N_119,In_363,In_205);
nand U120 (N_120,In_31,In_517);
nor U121 (N_121,In_1464,In_1267);
and U122 (N_122,In_960,In_905);
nor U123 (N_123,In_400,In_884);
nand U124 (N_124,In_133,In_927);
and U125 (N_125,In_1408,In_995);
or U126 (N_126,In_913,In_841);
or U127 (N_127,In_1242,In_1104);
nor U128 (N_128,In_1058,In_752);
or U129 (N_129,In_10,In_1229);
and U130 (N_130,In_1236,In_725);
xor U131 (N_131,In_260,In_687);
and U132 (N_132,In_938,In_1195);
or U133 (N_133,In_1038,In_831);
nor U134 (N_134,In_484,In_346);
and U135 (N_135,In_949,In_1076);
and U136 (N_136,In_341,In_570);
and U137 (N_137,In_1492,In_359);
nor U138 (N_138,In_616,In_1222);
and U139 (N_139,In_1239,In_391);
nand U140 (N_140,In_1289,In_918);
and U141 (N_141,In_300,In_407);
xnor U142 (N_142,In_1404,In_1218);
nand U143 (N_143,In_1140,In_1473);
nor U144 (N_144,In_1398,In_309);
and U145 (N_145,In_593,In_561);
nor U146 (N_146,In_1319,In_432);
nor U147 (N_147,In_410,In_1101);
xor U148 (N_148,In_212,In_1220);
nor U149 (N_149,In_814,In_1279);
or U150 (N_150,In_253,In_768);
or U151 (N_151,In_930,In_372);
or U152 (N_152,In_1471,In_165);
nor U153 (N_153,In_1031,In_1359);
and U154 (N_154,In_1117,In_1155);
nor U155 (N_155,In_1254,In_192);
and U156 (N_156,In_1423,In_1128);
and U157 (N_157,In_340,In_891);
and U158 (N_158,In_966,In_1421);
nand U159 (N_159,In_1345,In_1198);
nand U160 (N_160,In_1299,In_277);
nand U161 (N_161,In_1169,In_225);
and U162 (N_162,In_1263,In_1268);
and U163 (N_163,In_965,In_68);
or U164 (N_164,In_830,In_442);
nor U165 (N_165,In_1352,In_943);
nor U166 (N_166,In_1122,In_174);
nand U167 (N_167,In_74,In_1415);
or U168 (N_168,In_540,In_144);
nor U169 (N_169,In_1357,In_1209);
or U170 (N_170,In_678,In_1420);
nand U171 (N_171,In_135,In_741);
nand U172 (N_172,In_153,In_1015);
and U173 (N_173,In_971,In_1342);
nor U174 (N_174,In_409,In_463);
or U175 (N_175,In_1312,In_378);
nand U176 (N_176,In_320,In_881);
nand U177 (N_177,In_1334,In_843);
or U178 (N_178,In_1167,In_116);
or U179 (N_179,In_1463,In_1324);
nand U180 (N_180,In_193,In_306);
nor U181 (N_181,In_1252,In_840);
and U182 (N_182,In_365,In_11);
and U183 (N_183,In_1098,In_357);
nor U184 (N_184,In_285,In_800);
or U185 (N_185,In_1211,In_78);
nand U186 (N_186,In_749,In_238);
or U187 (N_187,In_269,In_1068);
or U188 (N_188,In_335,In_334);
and U189 (N_189,In_1282,In_179);
nand U190 (N_190,In_736,In_414);
and U191 (N_191,In_764,In_886);
and U192 (N_192,In_1301,In_198);
nor U193 (N_193,In_1186,In_595);
and U194 (N_194,In_1216,In_1095);
or U195 (N_195,In_1032,In_1494);
nor U196 (N_196,In_899,In_682);
xnor U197 (N_197,In_1188,In_1037);
nand U198 (N_198,In_1257,In_156);
and U199 (N_199,In_888,In_748);
nor U200 (N_200,In_0,In_1343);
or U201 (N_201,In_201,In_1082);
xor U202 (N_202,In_84,In_337);
or U203 (N_203,In_1164,In_216);
and U204 (N_204,In_588,In_157);
or U205 (N_205,In_399,In_487);
and U206 (N_206,In_864,In_951);
nor U207 (N_207,In_801,In_1086);
xnor U208 (N_208,In_512,In_544);
nor U209 (N_209,In_1062,In_962);
nand U210 (N_210,In_658,In_865);
xor U211 (N_211,In_1235,In_576);
xor U212 (N_212,In_301,In_532);
nor U213 (N_213,In_241,In_40);
and U214 (N_214,In_1308,In_702);
nand U215 (N_215,In_1154,In_1226);
nor U216 (N_216,In_308,In_1179);
and U217 (N_217,In_1029,In_1253);
or U218 (N_218,In_1190,In_906);
or U219 (N_219,In_425,In_415);
and U220 (N_220,In_635,In_994);
and U221 (N_221,In_858,In_413);
and U222 (N_222,In_1273,In_257);
nand U223 (N_223,In_243,In_1160);
nor U224 (N_224,In_942,In_224);
and U225 (N_225,In_454,In_914);
or U226 (N_226,In_20,In_1016);
nor U227 (N_227,In_1452,In_339);
nand U228 (N_228,In_1061,In_889);
and U229 (N_229,In_1083,In_1156);
nand U230 (N_230,In_1157,In_778);
or U231 (N_231,In_1131,In_118);
and U232 (N_232,In_1067,In_677);
and U233 (N_233,In_526,In_1379);
nor U234 (N_234,In_529,In_690);
and U235 (N_235,In_501,In_554);
nand U236 (N_236,In_839,In_210);
nand U237 (N_237,In_92,In_247);
or U238 (N_238,In_1141,In_319);
nor U239 (N_239,In_1259,In_1412);
nor U240 (N_240,In_1401,In_1331);
and U241 (N_241,In_1208,In_1056);
or U242 (N_242,In_175,In_521);
nand U243 (N_243,In_842,In_950);
or U244 (N_244,In_605,In_292);
and U245 (N_245,In_987,In_1042);
or U246 (N_246,In_1134,In_1472);
and U247 (N_247,In_322,In_1005);
and U248 (N_248,In_348,In_87);
nor U249 (N_249,In_472,In_1395);
nor U250 (N_250,In_1265,In_204);
nand U251 (N_251,In_184,In_1286);
and U252 (N_252,In_944,In_761);
nor U253 (N_253,In_1310,In_14);
nand U254 (N_254,In_898,In_283);
nor U255 (N_255,In_86,In_1030);
xnor U256 (N_256,In_1024,In_1488);
nor U257 (N_257,In_731,In_1079);
and U258 (N_258,In_1036,In_744);
and U259 (N_259,In_373,In_665);
or U260 (N_260,In_737,In_388);
or U261 (N_261,In_1476,In_1376);
nor U262 (N_262,In_868,In_967);
and U263 (N_263,In_1054,In_619);
xor U264 (N_264,In_1467,In_1449);
nor U265 (N_265,In_132,In_125);
xnor U266 (N_266,In_539,In_104);
xor U267 (N_267,In_27,In_747);
xor U268 (N_268,In_1228,In_762);
and U269 (N_269,In_989,In_1007);
and U270 (N_270,In_75,In_1162);
and U271 (N_271,In_797,In_859);
or U272 (N_272,In_77,In_427);
xnor U273 (N_273,In_1152,In_627);
nor U274 (N_274,In_1350,In_1137);
nor U275 (N_275,In_1478,In_323);
xor U276 (N_276,In_1138,In_1484);
and U277 (N_277,In_486,In_1087);
xor U278 (N_278,In_895,In_710);
and U279 (N_279,In_900,In_1123);
nor U280 (N_280,In_255,In_114);
or U281 (N_281,In_1440,In_360);
nand U282 (N_282,In_1246,In_485);
and U283 (N_283,In_172,In_755);
xnor U284 (N_284,In_429,In_447);
nor U285 (N_285,In_639,In_1006);
nor U286 (N_286,In_305,In_1240);
nor U287 (N_287,In_941,In_1028);
or U288 (N_288,In_609,In_1481);
xor U289 (N_289,In_849,In_173);
nand U290 (N_290,In_1204,In_314);
or U291 (N_291,In_1171,In_1102);
and U292 (N_292,In_1142,In_503);
nor U293 (N_293,In_522,In_42);
xnor U294 (N_294,In_1338,In_351);
xor U295 (N_295,In_195,In_287);
nor U296 (N_296,In_67,In_786);
nand U297 (N_297,In_798,In_765);
nor U298 (N_298,In_614,In_54);
nor U299 (N_299,In_1097,In_141);
nand U300 (N_300,In_310,In_160);
nor U301 (N_301,In_631,In_739);
or U302 (N_302,In_862,In_1210);
or U303 (N_303,In_304,In_608);
nor U304 (N_304,In_644,In_355);
or U305 (N_305,In_549,In_9);
xor U306 (N_306,In_1251,In_655);
nand U307 (N_307,In_1135,In_1163);
or U308 (N_308,In_169,In_1205);
or U309 (N_309,In_272,In_1292);
and U310 (N_310,In_1184,In_937);
and U311 (N_311,In_1072,In_1173);
and U312 (N_312,In_154,In_142);
and U313 (N_313,In_823,In_180);
xnor U314 (N_314,In_2,In_892);
and U315 (N_315,In_1139,In_857);
and U316 (N_316,In_1489,In_316);
and U317 (N_317,In_663,In_499);
nor U318 (N_318,In_455,In_1118);
nand U319 (N_319,In_1304,In_969);
xnor U320 (N_320,In_1182,In_395);
nand U321 (N_321,In_286,In_213);
and U322 (N_322,In_145,In_71);
and U323 (N_323,In_1483,In_466);
or U324 (N_324,In_1444,In_799);
nand U325 (N_325,In_251,In_29);
nor U326 (N_326,In_1305,In_215);
nor U327 (N_327,In_233,In_401);
nand U328 (N_328,In_620,In_1022);
or U329 (N_329,In_330,In_103);
nor U330 (N_330,In_1431,In_978);
and U331 (N_331,In_1318,In_1168);
nor U332 (N_332,In_767,In_815);
and U333 (N_333,In_933,In_37);
nand U334 (N_334,In_100,In_745);
nand U335 (N_335,In_325,In_686);
nor U336 (N_336,In_1017,In_844);
nor U337 (N_337,In_728,In_541);
nand U338 (N_338,In_863,In_812);
and U339 (N_339,In_1046,In_527);
nand U340 (N_340,In_458,In_838);
or U341 (N_341,In_428,In_1189);
nand U342 (N_342,In_1197,In_723);
and U343 (N_343,In_254,In_1426);
nand U344 (N_344,In_699,In_1110);
nand U345 (N_345,In_785,In_390);
or U346 (N_346,In_267,In_16);
or U347 (N_347,In_1245,In_488);
nor U348 (N_348,In_352,In_919);
nor U349 (N_349,In_207,In_735);
and U350 (N_350,In_845,In_268);
and U351 (N_351,In_1356,In_420);
nand U352 (N_352,In_81,In_1093);
xor U353 (N_353,In_504,In_1403);
or U354 (N_354,In_349,In_5);
or U355 (N_355,In_621,In_385);
and U356 (N_356,In_531,In_1219);
or U357 (N_357,In_569,In_794);
nand U358 (N_358,In_191,In_558);
nor U359 (N_359,In_998,In_934);
nand U360 (N_360,In_1344,In_1377);
nor U361 (N_361,In_43,In_1391);
xor U362 (N_362,In_23,In_370);
nor U363 (N_363,In_12,In_498);
nand U364 (N_364,In_177,In_7);
xor U365 (N_365,In_1477,In_35);
or U366 (N_366,In_1425,In_1130);
nand U367 (N_367,In_57,In_417);
nand U368 (N_368,In_51,In_17);
and U369 (N_369,In_1090,In_860);
nor U370 (N_370,In_353,In_1461);
nor U371 (N_371,In_929,In_947);
nand U372 (N_372,In_915,In_262);
nand U373 (N_373,In_124,In_580);
and U374 (N_374,In_158,In_1041);
xnor U375 (N_375,In_317,In_1317);
nand U376 (N_376,In_1121,In_916);
or U377 (N_377,In_907,In_742);
and U378 (N_378,In_18,In_396);
or U379 (N_379,In_219,In_1063);
or U380 (N_380,In_109,In_607);
nand U381 (N_381,In_997,In_1241);
and U382 (N_382,In_284,In_273);
and U383 (N_383,In_1326,In_1281);
and U384 (N_384,In_1196,In_804);
or U385 (N_385,In_362,In_1419);
nand U386 (N_386,In_1238,In_294);
nand U387 (N_387,In_632,In_307);
or U388 (N_388,In_925,In_510);
and U389 (N_389,In_659,In_1256);
nand U390 (N_390,In_1055,In_190);
nand U391 (N_391,In_416,In_419);
nor U392 (N_392,In_1386,In_1176);
or U393 (N_393,In_819,In_464);
nor U394 (N_394,In_164,In_1033);
nand U395 (N_395,In_1405,In_430);
nor U396 (N_396,In_775,In_1422);
nand U397 (N_397,In_1491,In_1428);
and U398 (N_398,In_1224,In_1207);
nor U399 (N_399,In_555,In_13);
nand U400 (N_400,In_1010,In_39);
or U401 (N_401,In_1382,In_1348);
nor U402 (N_402,In_1081,In_1271);
and U403 (N_403,In_386,In_1065);
nor U404 (N_404,In_500,In_666);
nand U405 (N_405,In_1451,In_19);
xor U406 (N_406,In_945,In_1192);
nor U407 (N_407,In_475,In_1064);
and U408 (N_408,In_1433,In_1250);
and U409 (N_409,In_1341,In_829);
nor U410 (N_410,In_1258,In_296);
or U411 (N_411,In_331,In_6);
nand U412 (N_412,In_1206,In_572);
and U413 (N_413,In_446,In_471);
nand U414 (N_414,In_751,In_290);
nor U415 (N_415,In_313,In_398);
or U416 (N_416,In_999,In_924);
or U417 (N_417,In_1441,In_1374);
xnor U418 (N_418,In_1244,In_733);
nor U419 (N_419,In_972,In_818);
nand U420 (N_420,In_563,In_926);
or U421 (N_421,In_381,In_976);
nor U422 (N_422,In_596,In_1158);
nand U423 (N_423,In_887,In_211);
and U424 (N_424,In_1214,In_489);
and U425 (N_425,In_753,In_991);
nor U426 (N_426,In_161,In_209);
nor U427 (N_427,In_1482,In_403);
nand U428 (N_428,In_777,In_451);
xor U429 (N_429,In_518,In_63);
nand U430 (N_430,In_1177,In_1322);
or U431 (N_431,In_382,In_24);
or U432 (N_432,In_1119,In_264);
xor U433 (N_433,In_389,In_1215);
nand U434 (N_434,In_1456,In_1103);
and U435 (N_435,In_782,In_832);
nand U436 (N_436,In_788,In_170);
nor U437 (N_437,In_189,In_870);
and U438 (N_438,In_795,In_387);
and U439 (N_439,In_1358,In_143);
and U440 (N_440,In_664,In_1183);
and U441 (N_441,In_459,In_1285);
or U442 (N_442,In_208,In_902);
nand U443 (N_443,In_750,In_1243);
nand U444 (N_444,In_96,In_112);
and U445 (N_445,In_1287,In_1088);
nor U446 (N_446,In_1302,In_97);
or U447 (N_447,In_681,In_566);
nor U448 (N_448,In_244,In_985);
or U449 (N_449,In_181,In_1384);
or U450 (N_450,In_1012,In_483);
or U451 (N_451,In_873,In_783);
nor U452 (N_452,In_222,In_123);
nand U453 (N_453,In_1127,In_1008);
or U454 (N_454,In_507,In_448);
xnor U455 (N_455,In_1278,In_1115);
nand U456 (N_456,In_1497,In_126);
nand U457 (N_457,In_374,In_1490);
and U458 (N_458,In_228,In_1096);
and U459 (N_459,In_746,In_1165);
or U460 (N_460,In_436,In_1366);
nor U461 (N_461,In_642,In_108);
nand U462 (N_462,In_931,In_1306);
nor U463 (N_463,In_393,In_1070);
and U464 (N_464,In_584,In_397);
and U465 (N_465,In_369,In_760);
nand U466 (N_466,In_248,In_26);
and U467 (N_467,In_1293,In_550);
or U468 (N_468,In_1225,In_923);
nor U469 (N_469,In_901,In_1448);
nor U470 (N_470,In_1272,In_647);
nand U471 (N_471,In_650,In_1199);
nor U472 (N_472,In_4,In_8);
nand U473 (N_473,In_662,In_679);
or U474 (N_474,In_652,In_854);
or U475 (N_475,In_1399,In_1203);
xor U476 (N_476,In_1277,In_1021);
nand U477 (N_477,In_482,In_672);
or U478 (N_478,In_64,In_1290);
or U479 (N_479,In_50,In_816);
xnor U480 (N_480,In_803,In_162);
and U481 (N_481,In_508,In_705);
and U482 (N_482,In_643,In_127);
xnor U483 (N_483,In_261,In_111);
nor U484 (N_484,In_922,In_876);
and U485 (N_485,In_249,In_72);
nor U486 (N_486,In_150,In_33);
xor U487 (N_487,In_1487,In_1339);
or U488 (N_488,In_155,In_617);
xor U489 (N_489,In_524,In_567);
or U490 (N_490,In_708,In_437);
nor U491 (N_491,In_721,In_611);
nor U492 (N_492,In_443,In_1075);
or U493 (N_493,In_1360,In_404);
nor U494 (N_494,In_920,In_984);
nor U495 (N_495,In_1438,In_796);
or U496 (N_496,In_1170,In_1002);
nor U497 (N_497,In_117,In_730);
or U498 (N_498,In_288,In_809);
xnor U499 (N_499,In_669,In_250);
or U500 (N_500,In_467,In_790);
and U501 (N_501,In_758,In_909);
or U502 (N_502,In_147,In_1417);
or U503 (N_503,In_129,In_58);
and U504 (N_504,In_1074,In_345);
nand U505 (N_505,In_1330,In_979);
nor U506 (N_506,In_491,In_633);
or U507 (N_507,In_1416,In_368);
or U508 (N_508,In_824,In_461);
nand U509 (N_509,In_689,In_959);
or U510 (N_510,In_671,In_1274);
nand U511 (N_511,In_932,In_904);
and U512 (N_512,In_557,In_439);
or U513 (N_513,In_612,In_714);
nor U514 (N_514,In_578,In_186);
nor U515 (N_515,In_618,In_698);
nand U516 (N_516,In_465,In_46);
or U517 (N_517,In_270,In_802);
nor U518 (N_518,In_433,In_1364);
or U519 (N_519,In_113,In_613);
and U520 (N_520,In_21,In_1023);
nand U521 (N_521,In_624,In_992);
or U522 (N_522,In_542,In_847);
or U523 (N_523,In_606,In_106);
or U524 (N_524,In_333,In_1411);
nor U525 (N_525,In_1402,In_47);
or U526 (N_526,In_1283,In_715);
nand U527 (N_527,In_1231,In_445);
nand U528 (N_528,In_431,In_1409);
xnor U529 (N_529,In_449,In_214);
nand U530 (N_530,In_110,In_1071);
or U531 (N_531,In_1453,In_121);
nand U532 (N_532,In_732,In_1291);
nor U533 (N_533,In_754,In_1309);
nor U534 (N_534,In_600,In_1212);
nand U535 (N_535,In_371,In_602);
nand U536 (N_536,In_422,In_908);
and U537 (N_537,In_328,In_476);
and U538 (N_538,In_1247,In_869);
nor U539 (N_539,In_329,In_1185);
nor U540 (N_540,In_1470,In_311);
or U541 (N_541,In_836,In_693);
and U542 (N_542,In_685,In_654);
nor U543 (N_543,In_1498,In_1161);
nand U544 (N_544,In_1109,In_776);
nand U545 (N_545,In_303,In_694);
nand U546 (N_546,In_1059,In_615);
and U547 (N_547,In_361,In_628);
nand U548 (N_548,In_1047,In_1387);
or U549 (N_549,In_1108,In_726);
or U550 (N_550,In_119,In_1148);
nand U551 (N_551,In_848,In_852);
and U552 (N_552,In_188,In_1388);
xor U553 (N_553,In_590,In_637);
or U554 (N_554,In_528,In_825);
or U555 (N_555,In_1085,In_692);
nand U556 (N_556,In_780,In_1260);
or U557 (N_557,In_598,In_871);
xnor U558 (N_558,In_281,In_1073);
or U559 (N_559,In_496,In_218);
or U560 (N_560,In_1003,In_1175);
and U561 (N_561,In_95,In_828);
xnor U562 (N_562,In_793,In_1458);
or U563 (N_563,In_1227,In_1328);
or U564 (N_564,In_478,In_1413);
nand U565 (N_565,In_1136,In_630);
nand U566 (N_566,In_1249,In_1354);
nor U567 (N_567,In_610,In_185);
nor U568 (N_568,In_1266,In_743);
or U569 (N_569,In_1389,In_1202);
nand U570 (N_570,In_101,In_1132);
and U571 (N_571,In_536,In_722);
xor U572 (N_572,In_149,In_939);
nor U573 (N_573,In_1213,In_1378);
nor U574 (N_574,In_1126,In_771);
nand U575 (N_575,In_1133,In_718);
nand U576 (N_576,In_298,In_1264);
nand U577 (N_577,In_727,In_1373);
nor U578 (N_578,In_105,In_1026);
nand U579 (N_579,In_936,In_151);
nand U580 (N_580,In_1447,In_41);
or U581 (N_581,In_1396,In_1445);
and U582 (N_582,In_599,In_581);
nor U583 (N_583,In_973,In_252);
or U584 (N_584,In_200,In_535);
or U585 (N_585,In_299,In_187);
nand U586 (N_586,In_556,In_131);
nand U587 (N_587,In_740,In_1013);
nor U588 (N_588,In_1457,In_675);
nor U589 (N_589,In_910,In_1049);
and U590 (N_590,In_1166,In_411);
and U591 (N_591,In_1107,In_479);
nor U592 (N_592,In_1261,In_203);
and U593 (N_593,In_293,In_1427);
nand U594 (N_594,In_1493,In_1436);
and U595 (N_595,In_1011,In_533);
or U596 (N_596,In_579,In_495);
nand U597 (N_597,In_1355,In_1069);
or U598 (N_598,In_1297,In_1051);
and U599 (N_599,In_1392,In_988);
xnor U600 (N_600,In_1335,In_1311);
and U601 (N_601,In_1437,In_130);
nor U602 (N_602,In_473,In_712);
nor U603 (N_603,In_952,In_1060);
and U604 (N_604,In_835,In_734);
and U605 (N_605,In_426,In_661);
nor U606 (N_606,In_826,In_1294);
or U607 (N_607,In_1314,In_986);
and U608 (N_608,In_582,In_176);
nor U609 (N_609,In_327,In_993);
and U610 (N_610,In_574,In_32);
and U611 (N_611,In_667,In_691);
and U612 (N_612,In_412,In_1315);
nor U613 (N_613,In_653,In_1390);
and U614 (N_614,In_622,In_996);
nand U615 (N_615,In_377,In_405);
or U616 (N_616,In_1080,In_897);
nand U617 (N_617,In_1050,In_589);
nor U618 (N_618,In_1336,In_221);
nor U619 (N_619,In_641,In_1084);
and U620 (N_620,In_376,In_440);
nor U621 (N_621,In_48,In_981);
or U622 (N_622,In_1300,In_1370);
and U623 (N_623,In_1349,In_738);
xor U624 (N_624,In_953,In_990);
and U625 (N_625,In_1474,In_434);
and U626 (N_626,In_538,In_1351);
or U627 (N_627,In_853,In_879);
and U628 (N_628,In_1180,In_1187);
or U629 (N_629,In_25,In_964);
and U630 (N_630,In_706,In_60);
and U631 (N_631,In_770,In_680);
xnor U632 (N_632,In_146,In_1178);
or U633 (N_633,In_457,In_1375);
nor U634 (N_634,In_318,In_649);
or U635 (N_635,In_676,In_278);
and U636 (N_636,In_375,In_1323);
xor U637 (N_637,In_1114,In_1221);
or U638 (N_638,In_321,In_577);
nand U639 (N_639,In_231,In_963);
nand U640 (N_640,In_79,In_492);
nor U641 (N_641,In_1369,In_1066);
nor U642 (N_642,In_1385,In_807);
nor U643 (N_643,In_1052,In_1143);
nand U644 (N_644,In_648,In_537);
nor U645 (N_645,In_406,In_354);
nand U646 (N_646,In_1078,In_65);
or U647 (N_647,In_634,In_573);
nand U648 (N_648,In_237,In_45);
or U649 (N_649,In_134,In_44);
xor U650 (N_650,In_490,In_592);
or U651 (N_651,In_302,In_1465);
or U652 (N_652,In_52,In_148);
xor U653 (N_653,In_94,In_342);
nand U654 (N_654,In_1094,In_1394);
or U655 (N_655,In_1307,In_547);
nor U656 (N_656,In_497,In_227);
and U657 (N_657,In_152,In_226);
nor U658 (N_658,In_366,In_636);
nand U659 (N_659,In_421,In_384);
nor U660 (N_660,In_1429,In_880);
nand U661 (N_661,In_312,In_1365);
and U662 (N_662,In_597,In_660);
and U663 (N_663,In_460,In_757);
nand U664 (N_664,In_601,In_217);
xnor U665 (N_665,In_645,In_1057);
nor U666 (N_666,In_202,In_1112);
nand U667 (N_667,In_22,In_1450);
nor U668 (N_668,In_1479,In_568);
and U669 (N_669,In_1149,In_545);
nor U670 (N_670,In_1459,In_38);
nor U671 (N_671,In_603,In_697);
nor U672 (N_672,In_295,In_822);
xor U673 (N_673,In_958,In_872);
xor U674 (N_674,In_696,In_946);
and U675 (N_675,In_1000,In_1129);
and U676 (N_676,In_813,In_559);
nor U677 (N_677,In_99,In_1280);
and U678 (N_678,In_1288,In_344);
xnor U679 (N_679,In_1381,In_66);
nor U680 (N_680,In_220,In_1346);
and U681 (N_681,In_553,In_668);
and U682 (N_682,In_552,In_683);
xor U683 (N_683,In_523,In_229);
or U684 (N_684,In_246,In_625);
nand U685 (N_685,In_274,In_279);
or U686 (N_686,In_890,In_364);
nand U687 (N_687,In_850,In_468);
and U688 (N_688,In_159,In_183);
or U689 (N_689,In_120,In_70);
nand U690 (N_690,In_1367,In_586);
nor U691 (N_691,In_1,In_759);
nor U692 (N_692,In_585,In_1193);
xnor U693 (N_693,In_56,In_1466);
nor U694 (N_694,In_1191,In_940);
nor U695 (N_695,In_968,In_1298);
or U696 (N_696,In_1039,In_1454);
nor U697 (N_697,In_275,In_324);
or U698 (N_698,In_1432,In_874);
or U699 (N_699,In_1014,In_1469);
xor U700 (N_700,In_509,In_571);
nor U701 (N_701,In_263,In_674);
and U702 (N_702,In_1455,In_810);
nor U703 (N_703,In_837,In_1269);
xnor U704 (N_704,In_61,In_350);
or U705 (N_705,In_515,In_626);
and U706 (N_706,In_326,In_784);
nand U707 (N_707,In_356,In_1332);
xnor U708 (N_708,In_583,In_1194);
and U709 (N_709,In_83,In_912);
or U710 (N_710,In_493,In_867);
nor U711 (N_711,In_138,In_462);
xnor U712 (N_712,In_670,In_1001);
and U713 (N_713,In_957,In_656);
nor U714 (N_714,In_182,In_982);
and U715 (N_715,In_587,In_338);
and U716 (N_716,In_1329,In_1303);
or U717 (N_717,In_1172,In_519);
nand U718 (N_718,In_548,In_1153);
or U719 (N_719,In_703,In_140);
and U720 (N_720,In_435,In_1053);
or U721 (N_721,In_977,In_1410);
nand U722 (N_722,In_1201,In_441);
nor U723 (N_723,In_1325,In_259);
nor U724 (N_724,In_1233,In_763);
or U725 (N_725,In_1316,In_1116);
nand U726 (N_726,In_1468,In_1020);
nor U727 (N_727,In_1439,In_383);
xor U728 (N_728,In_1146,In_1106);
nor U729 (N_729,In_948,In_1151);
or U730 (N_730,In_168,In_713);
and U731 (N_731,In_806,In_1091);
or U732 (N_732,In_604,In_701);
and U733 (N_733,In_1100,In_928);
or U734 (N_734,In_1035,In_1181);
nand U735 (N_735,In_673,In_980);
or U736 (N_736,In_343,In_833);
nand U737 (N_737,In_511,In_1200);
or U738 (N_738,In_358,In_36);
xnor U739 (N_739,In_885,In_1407);
or U740 (N_740,In_98,In_711);
or U741 (N_741,In_769,In_756);
and U742 (N_742,In_163,In_194);
and U743 (N_743,In_424,In_903);
nand U744 (N_744,In_1217,In_418);
or U745 (N_745,In_206,In_444);
nand U746 (N_746,In_392,In_80);
nor U747 (N_747,In_1034,In_1424);
nand U748 (N_748,In_456,In_69);
xnor U749 (N_749,In_1270,In_122);
xor U750 (N_750,N_127,N_563);
or U751 (N_751,N_485,N_110);
nor U752 (N_752,N_575,N_94);
and U753 (N_753,N_505,N_84);
nand U754 (N_754,N_689,N_481);
xnor U755 (N_755,N_403,N_239);
nor U756 (N_756,N_363,N_638);
nand U757 (N_757,N_2,N_371);
and U758 (N_758,N_188,N_649);
or U759 (N_759,N_144,N_646);
or U760 (N_760,N_426,N_396);
or U761 (N_761,N_669,N_738);
xnor U762 (N_762,N_235,N_639);
nand U763 (N_763,N_693,N_514);
and U764 (N_764,N_676,N_620);
or U765 (N_765,N_37,N_550);
nor U766 (N_766,N_245,N_421);
nand U767 (N_767,N_709,N_40);
nor U768 (N_768,N_310,N_398);
nor U769 (N_769,N_629,N_648);
nand U770 (N_770,N_488,N_197);
nand U771 (N_771,N_609,N_109);
nand U772 (N_772,N_584,N_7);
nand U773 (N_773,N_597,N_280);
xor U774 (N_774,N_46,N_315);
or U775 (N_775,N_636,N_521);
and U776 (N_776,N_680,N_251);
xnor U777 (N_777,N_591,N_205);
nand U778 (N_778,N_335,N_414);
nand U779 (N_779,N_287,N_356);
or U780 (N_780,N_65,N_719);
nor U781 (N_781,N_552,N_555);
nand U782 (N_782,N_498,N_723);
nor U783 (N_783,N_464,N_511);
nand U784 (N_784,N_444,N_373);
or U785 (N_785,N_473,N_141);
xor U786 (N_786,N_523,N_455);
nand U787 (N_787,N_282,N_492);
and U788 (N_788,N_657,N_89);
xnor U789 (N_789,N_705,N_580);
nand U790 (N_790,N_391,N_49);
or U791 (N_791,N_469,N_601);
nand U792 (N_792,N_194,N_710);
or U793 (N_793,N_113,N_634);
or U794 (N_794,N_377,N_101);
nor U795 (N_795,N_17,N_168);
xnor U796 (N_796,N_351,N_302);
nor U797 (N_797,N_131,N_456);
and U798 (N_798,N_29,N_367);
nor U799 (N_799,N_295,N_428);
nand U800 (N_800,N_561,N_123);
nor U801 (N_801,N_327,N_354);
nand U802 (N_802,N_407,N_355);
nand U803 (N_803,N_610,N_106);
and U804 (N_804,N_714,N_677);
nand U805 (N_805,N_218,N_128);
or U806 (N_806,N_497,N_577);
nor U807 (N_807,N_735,N_688);
or U808 (N_808,N_173,N_733);
nor U809 (N_809,N_328,N_274);
and U810 (N_810,N_27,N_85);
or U811 (N_811,N_558,N_269);
nor U812 (N_812,N_527,N_411);
nor U813 (N_813,N_494,N_319);
and U814 (N_814,N_368,N_486);
nand U815 (N_815,N_534,N_423);
nor U816 (N_816,N_145,N_210);
xor U817 (N_817,N_654,N_734);
xor U818 (N_818,N_692,N_663);
nand U819 (N_819,N_618,N_31);
and U820 (N_820,N_358,N_78);
nand U821 (N_821,N_572,N_275);
and U822 (N_822,N_71,N_250);
or U823 (N_823,N_38,N_139);
nor U824 (N_824,N_415,N_519);
or U825 (N_825,N_294,N_124);
or U826 (N_826,N_542,N_196);
nor U827 (N_827,N_360,N_329);
and U828 (N_828,N_81,N_731);
nor U829 (N_829,N_721,N_320);
xnor U830 (N_830,N_62,N_349);
nor U831 (N_831,N_400,N_202);
and U832 (N_832,N_626,N_437);
nand U833 (N_833,N_612,N_209);
nor U834 (N_834,N_248,N_331);
nand U835 (N_835,N_633,N_568);
nor U836 (N_836,N_416,N_249);
nand U837 (N_837,N_233,N_503);
nand U838 (N_838,N_531,N_678);
and U839 (N_839,N_402,N_201);
nand U840 (N_840,N_291,N_425);
nand U841 (N_841,N_451,N_67);
nor U842 (N_842,N_348,N_450);
nand U843 (N_843,N_615,N_696);
and U844 (N_844,N_433,N_230);
xnor U845 (N_845,N_495,N_125);
xor U846 (N_846,N_658,N_284);
nor U847 (N_847,N_301,N_483);
and U848 (N_848,N_379,N_224);
nand U849 (N_849,N_409,N_478);
nand U850 (N_850,N_161,N_446);
or U851 (N_851,N_720,N_30);
or U852 (N_852,N_55,N_187);
nand U853 (N_853,N_326,N_616);
or U854 (N_854,N_745,N_666);
and U855 (N_855,N_436,N_134);
and U856 (N_856,N_340,N_59);
xor U857 (N_857,N_376,N_681);
nor U858 (N_858,N_530,N_401);
and U859 (N_859,N_637,N_178);
or U860 (N_860,N_660,N_748);
nand U861 (N_861,N_405,N_307);
nor U862 (N_862,N_431,N_42);
xnor U863 (N_863,N_271,N_581);
nor U864 (N_864,N_189,N_621);
nand U865 (N_865,N_70,N_547);
nor U866 (N_866,N_607,N_746);
or U867 (N_867,N_664,N_64);
nor U868 (N_868,N_41,N_66);
or U869 (N_869,N_448,N_83);
nor U870 (N_870,N_685,N_317);
and U871 (N_871,N_278,N_247);
and U872 (N_872,N_728,N_491);
or U873 (N_873,N_632,N_102);
nor U874 (N_874,N_182,N_430);
nand U875 (N_875,N_704,N_252);
or U876 (N_876,N_6,N_179);
nand U877 (N_877,N_347,N_242);
and U878 (N_878,N_261,N_465);
and U879 (N_879,N_397,N_309);
xnor U880 (N_880,N_72,N_87);
nand U881 (N_881,N_298,N_36);
nor U882 (N_882,N_590,N_333);
or U883 (N_883,N_622,N_132);
nand U884 (N_884,N_671,N_191);
and U885 (N_885,N_549,N_545);
nor U886 (N_886,N_60,N_346);
nor U887 (N_887,N_662,N_493);
or U888 (N_888,N_596,N_404);
and U889 (N_889,N_151,N_244);
nor U890 (N_890,N_741,N_470);
or U891 (N_891,N_33,N_263);
and U892 (N_892,N_541,N_19);
xnor U893 (N_893,N_175,N_611);
xor U894 (N_894,N_744,N_14);
xnor U895 (N_895,N_392,N_177);
nand U896 (N_896,N_500,N_595);
xnor U897 (N_897,N_86,N_198);
nor U898 (N_898,N_655,N_343);
nand U899 (N_899,N_708,N_359);
or U900 (N_900,N_344,N_484);
nor U901 (N_901,N_332,N_614);
xnor U902 (N_902,N_142,N_449);
nor U903 (N_903,N_199,N_155);
and U904 (N_904,N_119,N_135);
nand U905 (N_905,N_221,N_675);
or U906 (N_906,N_700,N_672);
nor U907 (N_907,N_538,N_297);
nand U908 (N_908,N_279,N_435);
and U909 (N_909,N_747,N_10);
or U910 (N_910,N_441,N_389);
or U911 (N_911,N_432,N_73);
and U912 (N_912,N_157,N_589);
and U913 (N_913,N_195,N_463);
nand U914 (N_914,N_540,N_160);
nor U915 (N_915,N_467,N_385);
nor U916 (N_916,N_183,N_28);
or U917 (N_917,N_159,N_129);
xor U918 (N_918,N_91,N_418);
nor U919 (N_919,N_115,N_559);
nor U920 (N_920,N_314,N_554);
and U921 (N_921,N_578,N_476);
or U922 (N_922,N_305,N_624);
nor U923 (N_923,N_39,N_643);
nand U924 (N_924,N_501,N_118);
nor U925 (N_925,N_154,N_608);
nand U926 (N_926,N_574,N_277);
nor U927 (N_927,N_691,N_477);
and U928 (N_928,N_682,N_535);
and U929 (N_929,N_587,N_509);
or U930 (N_930,N_176,N_651);
nor U931 (N_931,N_592,N_18);
or U932 (N_932,N_267,N_0);
and U933 (N_933,N_701,N_726);
or U934 (N_934,N_730,N_338);
or U935 (N_935,N_516,N_126);
nor U936 (N_936,N_512,N_466);
nand U937 (N_937,N_241,N_47);
nand U938 (N_938,N_650,N_95);
nor U939 (N_939,N_399,N_357);
xor U940 (N_940,N_236,N_57);
nor U941 (N_941,N_533,N_253);
nor U942 (N_942,N_163,N_231);
nand U943 (N_943,N_1,N_300);
and U944 (N_944,N_15,N_353);
nor U945 (N_945,N_164,N_312);
and U946 (N_946,N_684,N_717);
and U947 (N_947,N_321,N_487);
nand U948 (N_948,N_56,N_200);
or U949 (N_949,N_507,N_63);
xnor U950 (N_950,N_690,N_311);
xor U951 (N_951,N_293,N_105);
nor U952 (N_952,N_656,N_214);
or U953 (N_953,N_289,N_556);
nor U954 (N_954,N_417,N_537);
and U955 (N_955,N_204,N_228);
nand U956 (N_956,N_502,N_605);
nor U957 (N_957,N_130,N_61);
or U958 (N_958,N_50,N_171);
xnor U959 (N_959,N_193,N_292);
xnor U960 (N_960,N_564,N_165);
and U961 (N_961,N_153,N_69);
nor U962 (N_962,N_108,N_75);
nor U963 (N_963,N_736,N_186);
or U964 (N_964,N_255,N_270);
and U965 (N_965,N_223,N_243);
xor U966 (N_966,N_361,N_58);
nand U967 (N_967,N_48,N_35);
nand U968 (N_968,N_99,N_652);
nand U969 (N_969,N_699,N_352);
nor U970 (N_970,N_316,N_372);
nor U971 (N_971,N_583,N_336);
xnor U972 (N_972,N_96,N_222);
nor U973 (N_973,N_16,N_167);
nor U974 (N_974,N_419,N_604);
nand U975 (N_975,N_11,N_54);
xnor U976 (N_976,N_140,N_136);
and U977 (N_977,N_475,N_266);
or U978 (N_978,N_232,N_458);
nand U979 (N_979,N_718,N_613);
xnor U980 (N_980,N_603,N_472);
and U981 (N_981,N_378,N_260);
and U982 (N_982,N_529,N_74);
or U983 (N_983,N_90,N_532);
and U984 (N_984,N_713,N_100);
nand U985 (N_985,N_536,N_229);
and U986 (N_986,N_468,N_264);
or U987 (N_987,N_619,N_286);
and U988 (N_988,N_308,N_749);
or U989 (N_989,N_370,N_114);
and U990 (N_990,N_546,N_234);
nand U991 (N_991,N_518,N_240);
xnor U992 (N_992,N_219,N_121);
nand U993 (N_993,N_422,N_285);
nor U994 (N_994,N_77,N_427);
nor U995 (N_995,N_686,N_12);
nor U996 (N_996,N_52,N_438);
nor U997 (N_997,N_299,N_152);
and U998 (N_998,N_216,N_715);
or U999 (N_999,N_350,N_306);
xnor U1000 (N_1000,N_26,N_3);
and U1001 (N_1001,N_585,N_169);
xor U1002 (N_1002,N_23,N_103);
and U1003 (N_1003,N_600,N_215);
or U1004 (N_1004,N_362,N_288);
or U1005 (N_1005,N_45,N_474);
nand U1006 (N_1006,N_325,N_625);
nor U1007 (N_1007,N_694,N_174);
and U1008 (N_1008,N_462,N_387);
or U1009 (N_1009,N_192,N_138);
or U1010 (N_1010,N_586,N_739);
or U1011 (N_1011,N_670,N_318);
nand U1012 (N_1012,N_383,N_479);
xnor U1013 (N_1013,N_573,N_567);
nand U1014 (N_1014,N_97,N_457);
nor U1015 (N_1015,N_459,N_21);
or U1016 (N_1016,N_642,N_185);
nand U1017 (N_1017,N_420,N_122);
or U1018 (N_1018,N_665,N_434);
nand U1019 (N_1019,N_339,N_345);
nand U1020 (N_1020,N_543,N_548);
nand U1021 (N_1021,N_562,N_172);
nand U1022 (N_1022,N_8,N_668);
and U1023 (N_1023,N_220,N_257);
nor U1024 (N_1024,N_226,N_147);
nand U1025 (N_1025,N_445,N_645);
nor U1026 (N_1026,N_259,N_588);
and U1027 (N_1027,N_313,N_203);
nand U1028 (N_1028,N_208,N_544);
nor U1029 (N_1029,N_517,N_729);
nand U1030 (N_1030,N_528,N_149);
nor U1031 (N_1031,N_722,N_212);
nand U1032 (N_1032,N_5,N_453);
nand U1033 (N_1033,N_594,N_213);
or U1034 (N_1034,N_256,N_447);
and U1035 (N_1035,N_93,N_323);
nand U1036 (N_1036,N_217,N_413);
nand U1037 (N_1037,N_570,N_272);
nor U1038 (N_1038,N_166,N_439);
nor U1039 (N_1039,N_80,N_206);
or U1040 (N_1040,N_265,N_667);
xor U1041 (N_1041,N_566,N_262);
and U1042 (N_1042,N_742,N_246);
nand U1043 (N_1043,N_82,N_565);
or U1044 (N_1044,N_724,N_111);
nand U1045 (N_1045,N_579,N_380);
or U1046 (N_1046,N_706,N_725);
or U1047 (N_1047,N_366,N_471);
nor U1048 (N_1048,N_640,N_375);
nor U1049 (N_1049,N_679,N_582);
or U1050 (N_1050,N_390,N_381);
nand U1051 (N_1051,N_190,N_184);
or U1052 (N_1052,N_254,N_51);
nand U1053 (N_1053,N_628,N_330);
and U1054 (N_1054,N_79,N_238);
nand U1055 (N_1055,N_489,N_661);
xor U1056 (N_1056,N_551,N_698);
nand U1057 (N_1057,N_408,N_395);
or U1058 (N_1058,N_225,N_296);
nor U1059 (N_1059,N_697,N_211);
xor U1060 (N_1060,N_88,N_647);
and U1061 (N_1061,N_342,N_20);
nor U1062 (N_1062,N_364,N_557);
nor U1063 (N_1063,N_442,N_24);
and U1064 (N_1064,N_635,N_560);
nor U1065 (N_1065,N_496,N_281);
nor U1066 (N_1066,N_273,N_116);
nand U1067 (N_1067,N_695,N_606);
or U1068 (N_1068,N_461,N_424);
nor U1069 (N_1069,N_452,N_599);
nand U1070 (N_1070,N_460,N_480);
and U1071 (N_1071,N_290,N_34);
nor U1072 (N_1072,N_576,N_386);
nor U1073 (N_1073,N_388,N_410);
nand U1074 (N_1074,N_513,N_227);
and U1075 (N_1075,N_641,N_683);
nand U1076 (N_1076,N_148,N_393);
nand U1077 (N_1077,N_727,N_22);
or U1078 (N_1078,N_394,N_9);
nor U1079 (N_1079,N_4,N_482);
or U1080 (N_1080,N_207,N_68);
and U1081 (N_1081,N_508,N_593);
nand U1082 (N_1082,N_539,N_743);
nand U1083 (N_1083,N_598,N_630);
or U1084 (N_1084,N_737,N_571);
xor U1085 (N_1085,N_53,N_740);
nand U1086 (N_1086,N_631,N_156);
and U1087 (N_1087,N_158,N_687);
nand U1088 (N_1088,N_412,N_443);
and U1089 (N_1089,N_322,N_520);
and U1090 (N_1090,N_644,N_341);
and U1091 (N_1091,N_524,N_525);
and U1092 (N_1092,N_659,N_499);
and U1093 (N_1093,N_107,N_334);
or U1094 (N_1094,N_133,N_653);
nor U1095 (N_1095,N_711,N_440);
nand U1096 (N_1096,N_374,N_703);
and U1097 (N_1097,N_522,N_98);
nand U1098 (N_1098,N_707,N_429);
xor U1099 (N_1099,N_673,N_569);
or U1100 (N_1100,N_143,N_120);
or U1101 (N_1101,N_162,N_490);
or U1102 (N_1102,N_702,N_369);
and U1103 (N_1103,N_732,N_76);
xnor U1104 (N_1104,N_43,N_454);
nand U1105 (N_1105,N_674,N_170);
nor U1106 (N_1106,N_627,N_506);
and U1107 (N_1107,N_515,N_268);
or U1108 (N_1108,N_324,N_180);
xor U1109 (N_1109,N_276,N_716);
or U1110 (N_1110,N_92,N_623);
or U1111 (N_1111,N_137,N_553);
nor U1112 (N_1112,N_365,N_25);
nand U1113 (N_1113,N_617,N_504);
nor U1114 (N_1114,N_510,N_337);
xor U1115 (N_1115,N_303,N_712);
nand U1116 (N_1116,N_258,N_112);
and U1117 (N_1117,N_104,N_382);
nor U1118 (N_1118,N_237,N_384);
and U1119 (N_1119,N_526,N_283);
or U1120 (N_1120,N_304,N_13);
and U1121 (N_1121,N_117,N_32);
xor U1122 (N_1122,N_150,N_146);
nor U1123 (N_1123,N_44,N_406);
nand U1124 (N_1124,N_181,N_602);
and U1125 (N_1125,N_649,N_541);
nor U1126 (N_1126,N_496,N_602);
nor U1127 (N_1127,N_150,N_254);
or U1128 (N_1128,N_565,N_201);
or U1129 (N_1129,N_393,N_109);
nor U1130 (N_1130,N_11,N_310);
nand U1131 (N_1131,N_590,N_574);
nor U1132 (N_1132,N_46,N_342);
and U1133 (N_1133,N_315,N_692);
nand U1134 (N_1134,N_166,N_241);
xor U1135 (N_1135,N_277,N_111);
nor U1136 (N_1136,N_668,N_83);
nand U1137 (N_1137,N_626,N_130);
and U1138 (N_1138,N_227,N_194);
nor U1139 (N_1139,N_568,N_183);
nor U1140 (N_1140,N_635,N_436);
or U1141 (N_1141,N_422,N_641);
or U1142 (N_1142,N_694,N_517);
nand U1143 (N_1143,N_250,N_604);
or U1144 (N_1144,N_573,N_586);
and U1145 (N_1145,N_617,N_712);
nor U1146 (N_1146,N_72,N_301);
nor U1147 (N_1147,N_331,N_237);
nor U1148 (N_1148,N_121,N_577);
nor U1149 (N_1149,N_742,N_269);
and U1150 (N_1150,N_619,N_575);
and U1151 (N_1151,N_392,N_246);
nor U1152 (N_1152,N_673,N_537);
nor U1153 (N_1153,N_310,N_541);
or U1154 (N_1154,N_548,N_560);
or U1155 (N_1155,N_137,N_292);
or U1156 (N_1156,N_299,N_404);
nand U1157 (N_1157,N_685,N_318);
and U1158 (N_1158,N_340,N_563);
or U1159 (N_1159,N_150,N_319);
nor U1160 (N_1160,N_56,N_308);
nor U1161 (N_1161,N_549,N_394);
nand U1162 (N_1162,N_11,N_569);
nor U1163 (N_1163,N_86,N_713);
nor U1164 (N_1164,N_55,N_275);
or U1165 (N_1165,N_684,N_164);
nor U1166 (N_1166,N_716,N_299);
or U1167 (N_1167,N_343,N_476);
nand U1168 (N_1168,N_304,N_366);
and U1169 (N_1169,N_347,N_245);
or U1170 (N_1170,N_323,N_598);
nand U1171 (N_1171,N_231,N_352);
nand U1172 (N_1172,N_121,N_130);
nand U1173 (N_1173,N_525,N_277);
and U1174 (N_1174,N_12,N_730);
nor U1175 (N_1175,N_357,N_212);
or U1176 (N_1176,N_368,N_674);
nor U1177 (N_1177,N_718,N_689);
nand U1178 (N_1178,N_212,N_22);
nor U1179 (N_1179,N_428,N_252);
nand U1180 (N_1180,N_389,N_293);
nor U1181 (N_1181,N_209,N_485);
or U1182 (N_1182,N_207,N_160);
nand U1183 (N_1183,N_188,N_339);
or U1184 (N_1184,N_33,N_469);
and U1185 (N_1185,N_324,N_686);
nor U1186 (N_1186,N_52,N_295);
and U1187 (N_1187,N_472,N_425);
or U1188 (N_1188,N_452,N_720);
xor U1189 (N_1189,N_498,N_525);
or U1190 (N_1190,N_277,N_174);
nor U1191 (N_1191,N_452,N_346);
or U1192 (N_1192,N_550,N_499);
nor U1193 (N_1193,N_337,N_708);
nor U1194 (N_1194,N_614,N_423);
and U1195 (N_1195,N_209,N_382);
xnor U1196 (N_1196,N_731,N_639);
xor U1197 (N_1197,N_462,N_689);
nand U1198 (N_1198,N_278,N_210);
and U1199 (N_1199,N_86,N_29);
nor U1200 (N_1200,N_355,N_9);
nor U1201 (N_1201,N_727,N_682);
nor U1202 (N_1202,N_135,N_375);
nor U1203 (N_1203,N_438,N_230);
nor U1204 (N_1204,N_429,N_14);
and U1205 (N_1205,N_291,N_253);
nor U1206 (N_1206,N_434,N_613);
and U1207 (N_1207,N_486,N_225);
nand U1208 (N_1208,N_233,N_418);
nand U1209 (N_1209,N_372,N_654);
nor U1210 (N_1210,N_306,N_65);
or U1211 (N_1211,N_81,N_732);
and U1212 (N_1212,N_267,N_17);
or U1213 (N_1213,N_542,N_497);
and U1214 (N_1214,N_679,N_512);
and U1215 (N_1215,N_591,N_53);
and U1216 (N_1216,N_457,N_269);
or U1217 (N_1217,N_730,N_175);
or U1218 (N_1218,N_235,N_279);
and U1219 (N_1219,N_171,N_642);
nand U1220 (N_1220,N_206,N_545);
or U1221 (N_1221,N_400,N_121);
and U1222 (N_1222,N_395,N_609);
nand U1223 (N_1223,N_712,N_545);
and U1224 (N_1224,N_109,N_140);
nor U1225 (N_1225,N_268,N_128);
and U1226 (N_1226,N_667,N_80);
nand U1227 (N_1227,N_340,N_305);
and U1228 (N_1228,N_608,N_491);
or U1229 (N_1229,N_681,N_84);
or U1230 (N_1230,N_361,N_319);
xnor U1231 (N_1231,N_706,N_404);
nand U1232 (N_1232,N_147,N_722);
and U1233 (N_1233,N_287,N_33);
nand U1234 (N_1234,N_403,N_545);
and U1235 (N_1235,N_396,N_257);
nor U1236 (N_1236,N_153,N_653);
nor U1237 (N_1237,N_579,N_433);
nand U1238 (N_1238,N_518,N_604);
and U1239 (N_1239,N_694,N_237);
nand U1240 (N_1240,N_443,N_269);
and U1241 (N_1241,N_719,N_732);
nand U1242 (N_1242,N_414,N_144);
nor U1243 (N_1243,N_661,N_208);
nand U1244 (N_1244,N_60,N_264);
nand U1245 (N_1245,N_185,N_245);
or U1246 (N_1246,N_318,N_483);
nand U1247 (N_1247,N_36,N_321);
nand U1248 (N_1248,N_625,N_666);
nand U1249 (N_1249,N_208,N_466);
or U1250 (N_1250,N_314,N_464);
nor U1251 (N_1251,N_511,N_339);
nor U1252 (N_1252,N_406,N_212);
and U1253 (N_1253,N_4,N_498);
nor U1254 (N_1254,N_577,N_166);
and U1255 (N_1255,N_281,N_493);
nor U1256 (N_1256,N_141,N_26);
and U1257 (N_1257,N_88,N_213);
and U1258 (N_1258,N_617,N_336);
and U1259 (N_1259,N_561,N_251);
or U1260 (N_1260,N_634,N_101);
nor U1261 (N_1261,N_180,N_161);
nand U1262 (N_1262,N_358,N_277);
and U1263 (N_1263,N_576,N_642);
nand U1264 (N_1264,N_50,N_183);
nor U1265 (N_1265,N_587,N_308);
nor U1266 (N_1266,N_724,N_438);
nand U1267 (N_1267,N_589,N_34);
or U1268 (N_1268,N_85,N_735);
xnor U1269 (N_1269,N_372,N_107);
nor U1270 (N_1270,N_245,N_215);
or U1271 (N_1271,N_196,N_33);
nand U1272 (N_1272,N_411,N_627);
nand U1273 (N_1273,N_667,N_204);
nand U1274 (N_1274,N_189,N_239);
nor U1275 (N_1275,N_61,N_340);
and U1276 (N_1276,N_712,N_742);
nand U1277 (N_1277,N_308,N_28);
nand U1278 (N_1278,N_731,N_192);
or U1279 (N_1279,N_63,N_590);
and U1280 (N_1280,N_587,N_571);
and U1281 (N_1281,N_165,N_299);
nor U1282 (N_1282,N_394,N_60);
and U1283 (N_1283,N_402,N_133);
and U1284 (N_1284,N_234,N_491);
xnor U1285 (N_1285,N_588,N_518);
nor U1286 (N_1286,N_8,N_193);
nor U1287 (N_1287,N_222,N_635);
and U1288 (N_1288,N_709,N_611);
or U1289 (N_1289,N_6,N_14);
or U1290 (N_1290,N_539,N_738);
and U1291 (N_1291,N_228,N_169);
nor U1292 (N_1292,N_423,N_216);
and U1293 (N_1293,N_539,N_721);
and U1294 (N_1294,N_738,N_137);
xnor U1295 (N_1295,N_467,N_14);
nor U1296 (N_1296,N_343,N_23);
and U1297 (N_1297,N_677,N_267);
nor U1298 (N_1298,N_405,N_711);
xnor U1299 (N_1299,N_52,N_313);
nor U1300 (N_1300,N_722,N_222);
nand U1301 (N_1301,N_238,N_59);
nor U1302 (N_1302,N_456,N_342);
and U1303 (N_1303,N_486,N_223);
and U1304 (N_1304,N_193,N_580);
or U1305 (N_1305,N_59,N_186);
or U1306 (N_1306,N_229,N_518);
or U1307 (N_1307,N_577,N_186);
xnor U1308 (N_1308,N_699,N_647);
nand U1309 (N_1309,N_232,N_724);
and U1310 (N_1310,N_366,N_359);
nor U1311 (N_1311,N_558,N_286);
or U1312 (N_1312,N_145,N_466);
nor U1313 (N_1313,N_252,N_123);
nand U1314 (N_1314,N_593,N_63);
nand U1315 (N_1315,N_44,N_634);
nor U1316 (N_1316,N_270,N_358);
and U1317 (N_1317,N_167,N_725);
nor U1318 (N_1318,N_353,N_687);
nand U1319 (N_1319,N_64,N_647);
xor U1320 (N_1320,N_37,N_545);
xnor U1321 (N_1321,N_51,N_91);
xor U1322 (N_1322,N_391,N_67);
and U1323 (N_1323,N_746,N_423);
or U1324 (N_1324,N_14,N_650);
and U1325 (N_1325,N_488,N_149);
nor U1326 (N_1326,N_685,N_416);
or U1327 (N_1327,N_116,N_733);
and U1328 (N_1328,N_456,N_78);
xnor U1329 (N_1329,N_233,N_353);
and U1330 (N_1330,N_311,N_551);
and U1331 (N_1331,N_5,N_386);
nand U1332 (N_1332,N_462,N_478);
or U1333 (N_1333,N_653,N_635);
nor U1334 (N_1334,N_425,N_345);
and U1335 (N_1335,N_681,N_8);
nand U1336 (N_1336,N_424,N_613);
nand U1337 (N_1337,N_632,N_701);
nand U1338 (N_1338,N_280,N_577);
nand U1339 (N_1339,N_351,N_651);
nor U1340 (N_1340,N_380,N_114);
and U1341 (N_1341,N_255,N_72);
and U1342 (N_1342,N_50,N_277);
nand U1343 (N_1343,N_621,N_427);
xnor U1344 (N_1344,N_273,N_420);
and U1345 (N_1345,N_4,N_474);
nor U1346 (N_1346,N_288,N_571);
nor U1347 (N_1347,N_260,N_371);
or U1348 (N_1348,N_199,N_590);
and U1349 (N_1349,N_539,N_231);
nor U1350 (N_1350,N_174,N_644);
nand U1351 (N_1351,N_520,N_539);
nor U1352 (N_1352,N_59,N_231);
or U1353 (N_1353,N_270,N_16);
and U1354 (N_1354,N_147,N_76);
and U1355 (N_1355,N_337,N_212);
nor U1356 (N_1356,N_459,N_391);
nand U1357 (N_1357,N_195,N_731);
or U1358 (N_1358,N_232,N_648);
nand U1359 (N_1359,N_343,N_623);
and U1360 (N_1360,N_749,N_618);
or U1361 (N_1361,N_408,N_310);
xnor U1362 (N_1362,N_326,N_514);
xor U1363 (N_1363,N_595,N_129);
nor U1364 (N_1364,N_128,N_584);
or U1365 (N_1365,N_128,N_706);
nand U1366 (N_1366,N_405,N_146);
nand U1367 (N_1367,N_440,N_408);
and U1368 (N_1368,N_636,N_247);
nor U1369 (N_1369,N_216,N_552);
nor U1370 (N_1370,N_45,N_294);
and U1371 (N_1371,N_193,N_10);
and U1372 (N_1372,N_502,N_40);
and U1373 (N_1373,N_69,N_167);
and U1374 (N_1374,N_242,N_587);
nor U1375 (N_1375,N_701,N_602);
nor U1376 (N_1376,N_464,N_130);
nand U1377 (N_1377,N_647,N_235);
nand U1378 (N_1378,N_152,N_326);
nor U1379 (N_1379,N_358,N_544);
nand U1380 (N_1380,N_568,N_36);
or U1381 (N_1381,N_404,N_123);
and U1382 (N_1382,N_103,N_217);
or U1383 (N_1383,N_725,N_583);
and U1384 (N_1384,N_585,N_253);
and U1385 (N_1385,N_639,N_674);
and U1386 (N_1386,N_264,N_48);
and U1387 (N_1387,N_342,N_742);
or U1388 (N_1388,N_109,N_195);
nor U1389 (N_1389,N_28,N_26);
nand U1390 (N_1390,N_576,N_267);
nand U1391 (N_1391,N_396,N_587);
nor U1392 (N_1392,N_275,N_219);
nand U1393 (N_1393,N_408,N_716);
or U1394 (N_1394,N_47,N_637);
and U1395 (N_1395,N_295,N_495);
nor U1396 (N_1396,N_322,N_7);
nor U1397 (N_1397,N_449,N_151);
nor U1398 (N_1398,N_329,N_262);
xor U1399 (N_1399,N_410,N_733);
nand U1400 (N_1400,N_439,N_535);
or U1401 (N_1401,N_667,N_649);
and U1402 (N_1402,N_708,N_620);
or U1403 (N_1403,N_399,N_248);
or U1404 (N_1404,N_70,N_505);
or U1405 (N_1405,N_641,N_179);
and U1406 (N_1406,N_268,N_53);
and U1407 (N_1407,N_303,N_144);
and U1408 (N_1408,N_270,N_693);
or U1409 (N_1409,N_705,N_153);
or U1410 (N_1410,N_243,N_392);
nand U1411 (N_1411,N_204,N_164);
or U1412 (N_1412,N_390,N_334);
nor U1413 (N_1413,N_695,N_549);
nand U1414 (N_1414,N_655,N_232);
and U1415 (N_1415,N_8,N_263);
and U1416 (N_1416,N_471,N_266);
xor U1417 (N_1417,N_295,N_38);
and U1418 (N_1418,N_129,N_93);
nor U1419 (N_1419,N_81,N_166);
and U1420 (N_1420,N_532,N_414);
xor U1421 (N_1421,N_122,N_376);
or U1422 (N_1422,N_693,N_547);
or U1423 (N_1423,N_596,N_511);
nand U1424 (N_1424,N_243,N_95);
and U1425 (N_1425,N_648,N_694);
nor U1426 (N_1426,N_167,N_235);
and U1427 (N_1427,N_208,N_726);
and U1428 (N_1428,N_289,N_67);
nand U1429 (N_1429,N_423,N_690);
nor U1430 (N_1430,N_571,N_539);
nor U1431 (N_1431,N_407,N_404);
nand U1432 (N_1432,N_212,N_427);
nor U1433 (N_1433,N_279,N_277);
and U1434 (N_1434,N_636,N_696);
nand U1435 (N_1435,N_330,N_460);
nor U1436 (N_1436,N_506,N_249);
and U1437 (N_1437,N_199,N_44);
or U1438 (N_1438,N_544,N_231);
xnor U1439 (N_1439,N_376,N_584);
and U1440 (N_1440,N_171,N_127);
and U1441 (N_1441,N_282,N_399);
nor U1442 (N_1442,N_540,N_560);
and U1443 (N_1443,N_717,N_705);
nand U1444 (N_1444,N_488,N_414);
and U1445 (N_1445,N_676,N_470);
or U1446 (N_1446,N_696,N_31);
or U1447 (N_1447,N_468,N_151);
nand U1448 (N_1448,N_606,N_116);
xnor U1449 (N_1449,N_326,N_273);
nor U1450 (N_1450,N_623,N_598);
nand U1451 (N_1451,N_162,N_377);
nand U1452 (N_1452,N_240,N_624);
and U1453 (N_1453,N_378,N_246);
nor U1454 (N_1454,N_91,N_426);
nand U1455 (N_1455,N_204,N_281);
nor U1456 (N_1456,N_109,N_560);
or U1457 (N_1457,N_728,N_522);
xor U1458 (N_1458,N_172,N_589);
nor U1459 (N_1459,N_50,N_661);
and U1460 (N_1460,N_144,N_682);
nor U1461 (N_1461,N_197,N_156);
and U1462 (N_1462,N_56,N_41);
nand U1463 (N_1463,N_612,N_279);
nand U1464 (N_1464,N_336,N_555);
and U1465 (N_1465,N_650,N_175);
and U1466 (N_1466,N_446,N_593);
nand U1467 (N_1467,N_687,N_606);
xor U1468 (N_1468,N_162,N_630);
nor U1469 (N_1469,N_471,N_650);
or U1470 (N_1470,N_222,N_620);
or U1471 (N_1471,N_510,N_304);
nor U1472 (N_1472,N_631,N_173);
and U1473 (N_1473,N_109,N_491);
nand U1474 (N_1474,N_573,N_125);
or U1475 (N_1475,N_356,N_621);
nand U1476 (N_1476,N_146,N_216);
or U1477 (N_1477,N_548,N_262);
nor U1478 (N_1478,N_382,N_126);
xor U1479 (N_1479,N_618,N_400);
nor U1480 (N_1480,N_356,N_354);
nor U1481 (N_1481,N_635,N_251);
nand U1482 (N_1482,N_497,N_387);
and U1483 (N_1483,N_83,N_314);
and U1484 (N_1484,N_517,N_117);
nand U1485 (N_1485,N_175,N_376);
nor U1486 (N_1486,N_722,N_160);
xor U1487 (N_1487,N_728,N_89);
nor U1488 (N_1488,N_241,N_306);
nand U1489 (N_1489,N_412,N_497);
or U1490 (N_1490,N_590,N_563);
xnor U1491 (N_1491,N_185,N_405);
and U1492 (N_1492,N_624,N_142);
or U1493 (N_1493,N_142,N_78);
or U1494 (N_1494,N_432,N_348);
nand U1495 (N_1495,N_735,N_253);
nand U1496 (N_1496,N_291,N_749);
and U1497 (N_1497,N_245,N_371);
nand U1498 (N_1498,N_560,N_305);
nor U1499 (N_1499,N_341,N_173);
and U1500 (N_1500,N_991,N_1308);
nand U1501 (N_1501,N_1330,N_926);
or U1502 (N_1502,N_984,N_1039);
xor U1503 (N_1503,N_888,N_1398);
or U1504 (N_1504,N_1034,N_1225);
or U1505 (N_1505,N_760,N_869);
and U1506 (N_1506,N_1060,N_1223);
nor U1507 (N_1507,N_1464,N_1085);
xor U1508 (N_1508,N_1078,N_1089);
or U1509 (N_1509,N_1116,N_1099);
nand U1510 (N_1510,N_1117,N_1327);
and U1511 (N_1511,N_1028,N_1322);
and U1512 (N_1512,N_1363,N_1016);
and U1513 (N_1513,N_824,N_961);
and U1514 (N_1514,N_898,N_1254);
and U1515 (N_1515,N_1093,N_765);
xor U1516 (N_1516,N_1177,N_921);
nand U1517 (N_1517,N_822,N_1451);
nand U1518 (N_1518,N_1165,N_1010);
nor U1519 (N_1519,N_1154,N_1475);
or U1520 (N_1520,N_1247,N_1120);
and U1521 (N_1521,N_1394,N_838);
nor U1522 (N_1522,N_856,N_1113);
and U1523 (N_1523,N_1101,N_1454);
nor U1524 (N_1524,N_1468,N_1022);
nor U1525 (N_1525,N_1407,N_1395);
or U1526 (N_1526,N_1412,N_771);
nand U1527 (N_1527,N_1420,N_863);
nor U1528 (N_1528,N_1459,N_1440);
and U1529 (N_1529,N_1405,N_1448);
xor U1530 (N_1530,N_1240,N_879);
nor U1531 (N_1531,N_1059,N_1343);
nand U1532 (N_1532,N_1350,N_1422);
nand U1533 (N_1533,N_1178,N_1014);
nand U1534 (N_1534,N_1311,N_1300);
and U1535 (N_1535,N_1435,N_1095);
and U1536 (N_1536,N_1072,N_1157);
nand U1537 (N_1537,N_759,N_1358);
or U1538 (N_1538,N_1334,N_828);
and U1539 (N_1539,N_1442,N_779);
nand U1540 (N_1540,N_1069,N_1482);
nand U1541 (N_1541,N_1104,N_1004);
or U1542 (N_1542,N_1032,N_797);
and U1543 (N_1543,N_900,N_975);
nand U1544 (N_1544,N_1195,N_945);
nand U1545 (N_1545,N_761,N_1337);
xor U1546 (N_1546,N_1091,N_1074);
nor U1547 (N_1547,N_1159,N_920);
nor U1548 (N_1548,N_1299,N_1233);
or U1549 (N_1549,N_1105,N_978);
nor U1550 (N_1550,N_1203,N_1474);
and U1551 (N_1551,N_1441,N_1268);
or U1552 (N_1552,N_1281,N_820);
nand U1553 (N_1553,N_1346,N_783);
and U1554 (N_1554,N_874,N_878);
or U1555 (N_1555,N_834,N_1221);
and U1556 (N_1556,N_1293,N_1287);
nand U1557 (N_1557,N_1055,N_1109);
nand U1558 (N_1558,N_1415,N_1166);
nand U1559 (N_1559,N_854,N_1296);
and U1560 (N_1560,N_1145,N_1298);
xor U1561 (N_1561,N_1027,N_876);
and U1562 (N_1562,N_1487,N_1385);
or U1563 (N_1563,N_968,N_950);
or U1564 (N_1564,N_793,N_1042);
and U1565 (N_1565,N_754,N_864);
nor U1566 (N_1566,N_826,N_1488);
and U1567 (N_1567,N_1272,N_1494);
or U1568 (N_1568,N_1457,N_1273);
or U1569 (N_1569,N_1124,N_1387);
and U1570 (N_1570,N_932,N_1163);
nand U1571 (N_1571,N_1244,N_847);
or U1572 (N_1572,N_1253,N_1108);
or U1573 (N_1573,N_1131,N_1406);
xnor U1574 (N_1574,N_1278,N_1252);
xor U1575 (N_1575,N_1054,N_1066);
nand U1576 (N_1576,N_1188,N_1368);
nand U1577 (N_1577,N_887,N_1047);
or U1578 (N_1578,N_767,N_1257);
nand U1579 (N_1579,N_936,N_1173);
and U1580 (N_1580,N_948,N_852);
nor U1581 (N_1581,N_1447,N_1477);
and U1582 (N_1582,N_867,N_1226);
and U1583 (N_1583,N_1331,N_1160);
nand U1584 (N_1584,N_1062,N_1276);
or U1585 (N_1585,N_832,N_1456);
or U1586 (N_1586,N_938,N_962);
xnor U1587 (N_1587,N_997,N_1029);
xnor U1588 (N_1588,N_1156,N_1248);
or U1589 (N_1589,N_877,N_1017);
xnor U1590 (N_1590,N_897,N_1121);
or U1591 (N_1591,N_947,N_1008);
and U1592 (N_1592,N_1191,N_934);
nor U1593 (N_1593,N_1262,N_1251);
nor U1594 (N_1594,N_976,N_1397);
and U1595 (N_1595,N_843,N_780);
nor U1596 (N_1596,N_808,N_971);
nor U1597 (N_1597,N_1041,N_1045);
and U1598 (N_1598,N_811,N_1158);
and U1599 (N_1599,N_1270,N_1123);
xor U1600 (N_1600,N_794,N_1438);
and U1601 (N_1601,N_953,N_775);
or U1602 (N_1602,N_1470,N_1354);
nor U1603 (N_1603,N_1367,N_1023);
nor U1604 (N_1604,N_1351,N_1231);
or U1605 (N_1605,N_883,N_972);
and U1606 (N_1606,N_1100,N_1467);
and U1607 (N_1607,N_1134,N_836);
nand U1608 (N_1608,N_770,N_1349);
and U1609 (N_1609,N_1288,N_1384);
nand U1610 (N_1610,N_1185,N_807);
nor U1611 (N_1611,N_1238,N_1040);
and U1612 (N_1612,N_848,N_930);
nor U1613 (N_1613,N_1208,N_1266);
nand U1614 (N_1614,N_1135,N_1212);
or U1615 (N_1615,N_964,N_1321);
xnor U1616 (N_1616,N_777,N_1403);
nor U1617 (N_1617,N_985,N_1046);
nand U1618 (N_1618,N_1162,N_1480);
nand U1619 (N_1619,N_1472,N_1357);
or U1620 (N_1620,N_1033,N_855);
nand U1621 (N_1621,N_1437,N_899);
nor U1622 (N_1622,N_1003,N_1416);
nand U1623 (N_1623,N_1277,N_1176);
xor U1624 (N_1624,N_1137,N_1168);
nor U1625 (N_1625,N_1218,N_784);
or U1626 (N_1626,N_1199,N_1297);
nand U1627 (N_1627,N_861,N_918);
xor U1628 (N_1628,N_1414,N_1289);
nor U1629 (N_1629,N_816,N_1138);
nand U1630 (N_1630,N_1064,N_798);
nand U1631 (N_1631,N_1020,N_1361);
or U1632 (N_1632,N_1452,N_1431);
or U1633 (N_1633,N_1471,N_805);
nor U1634 (N_1634,N_1317,N_1386);
nor U1635 (N_1635,N_956,N_1312);
nand U1636 (N_1636,N_1473,N_1338);
and U1637 (N_1637,N_789,N_1460);
and U1638 (N_1638,N_873,N_1360);
or U1639 (N_1639,N_1082,N_1413);
nand U1640 (N_1640,N_1325,N_1110);
nor U1641 (N_1641,N_967,N_1285);
or U1642 (N_1642,N_882,N_939);
nand U1643 (N_1643,N_1161,N_815);
xnor U1644 (N_1644,N_1106,N_1002);
xnor U1645 (N_1645,N_1122,N_1115);
or U1646 (N_1646,N_1245,N_829);
and U1647 (N_1647,N_1219,N_924);
or U1648 (N_1648,N_1282,N_868);
nor U1649 (N_1649,N_951,N_1453);
nor U1650 (N_1650,N_943,N_1377);
and U1651 (N_1651,N_1205,N_764);
and U1652 (N_1652,N_954,N_1497);
xor U1653 (N_1653,N_1392,N_766);
nor U1654 (N_1654,N_1376,N_1190);
nand U1655 (N_1655,N_941,N_1126);
or U1656 (N_1656,N_916,N_1409);
or U1657 (N_1657,N_1379,N_965);
xnor U1658 (N_1658,N_1133,N_917);
or U1659 (N_1659,N_757,N_1043);
or U1660 (N_1660,N_772,N_1426);
nand U1661 (N_1661,N_823,N_1214);
nand U1662 (N_1662,N_1466,N_751);
nor U1663 (N_1663,N_1209,N_1217);
nand U1664 (N_1664,N_1388,N_1275);
nand U1665 (N_1665,N_933,N_1345);
nand U1666 (N_1666,N_911,N_1206);
and U1667 (N_1667,N_1381,N_1071);
nor U1668 (N_1668,N_804,N_1329);
nor U1669 (N_1669,N_1044,N_1035);
xor U1670 (N_1670,N_1344,N_1210);
or U1671 (N_1671,N_1433,N_891);
nor U1672 (N_1672,N_1179,N_859);
nor U1673 (N_1673,N_974,N_1012);
or U1674 (N_1674,N_831,N_788);
nor U1675 (N_1675,N_884,N_1286);
and U1676 (N_1676,N_1372,N_889);
nor U1677 (N_1677,N_1320,N_803);
xnor U1678 (N_1678,N_922,N_1485);
xor U1679 (N_1679,N_928,N_1242);
nor U1680 (N_1680,N_1196,N_1142);
and U1681 (N_1681,N_1170,N_1256);
xor U1682 (N_1682,N_1332,N_1025);
or U1683 (N_1683,N_850,N_980);
and U1684 (N_1684,N_791,N_774);
and U1685 (N_1685,N_833,N_1063);
and U1686 (N_1686,N_769,N_1175);
xnor U1687 (N_1687,N_894,N_1213);
nor U1688 (N_1688,N_1495,N_1197);
and U1689 (N_1689,N_905,N_1303);
and U1690 (N_1690,N_909,N_1198);
nor U1691 (N_1691,N_1237,N_1476);
and U1692 (N_1692,N_973,N_1427);
nand U1693 (N_1693,N_1499,N_778);
or U1694 (N_1694,N_758,N_1302);
xnor U1695 (N_1695,N_993,N_812);
xor U1696 (N_1696,N_750,N_1061);
and U1697 (N_1697,N_762,N_810);
and U1698 (N_1698,N_1235,N_969);
nand U1699 (N_1699,N_935,N_994);
or U1700 (N_1700,N_1411,N_1114);
and U1701 (N_1701,N_1193,N_1383);
and U1702 (N_1702,N_919,N_957);
and U1703 (N_1703,N_1141,N_1481);
xnor U1704 (N_1704,N_1182,N_1271);
or U1705 (N_1705,N_1184,N_801);
nand U1706 (N_1706,N_1153,N_1150);
nand U1707 (N_1707,N_1366,N_987);
nor U1708 (N_1708,N_837,N_1132);
or U1709 (N_1709,N_1102,N_1006);
xnor U1710 (N_1710,N_1484,N_785);
and U1711 (N_1711,N_1018,N_875);
or U1712 (N_1712,N_809,N_1201);
and U1713 (N_1713,N_1274,N_979);
and U1714 (N_1714,N_1015,N_1423);
nand U1715 (N_1715,N_782,N_763);
or U1716 (N_1716,N_914,N_1469);
nand U1717 (N_1717,N_1463,N_1404);
nand U1718 (N_1718,N_1450,N_1342);
nand U1719 (N_1719,N_990,N_942);
and U1720 (N_1720,N_1211,N_1465);
and U1721 (N_1721,N_1417,N_923);
or U1722 (N_1722,N_960,N_1369);
nand U1723 (N_1723,N_1455,N_1491);
or U1724 (N_1724,N_1310,N_1019);
and U1725 (N_1725,N_1048,N_892);
or U1726 (N_1726,N_1283,N_1186);
xnor U1727 (N_1727,N_1216,N_1077);
nand U1728 (N_1728,N_949,N_1147);
and U1729 (N_1729,N_1348,N_1097);
nand U1730 (N_1730,N_1373,N_860);
xor U1731 (N_1731,N_1391,N_1424);
or U1732 (N_1732,N_806,N_925);
nor U1733 (N_1733,N_1462,N_1228);
and U1734 (N_1734,N_1084,N_1478);
and U1735 (N_1735,N_1449,N_1169);
nand U1736 (N_1736,N_1425,N_871);
nand U1737 (N_1737,N_1492,N_1396);
nor U1738 (N_1738,N_1430,N_865);
nand U1739 (N_1739,N_986,N_776);
or U1740 (N_1740,N_1222,N_1443);
or U1741 (N_1741,N_1336,N_958);
xnor U1742 (N_1742,N_1374,N_1259);
nor U1743 (N_1743,N_1439,N_952);
and U1744 (N_1744,N_1079,N_1056);
and U1745 (N_1745,N_1402,N_1068);
and U1746 (N_1746,N_931,N_1075);
xor U1747 (N_1747,N_1207,N_818);
nand U1748 (N_1748,N_1243,N_1128);
or U1749 (N_1749,N_1227,N_1365);
nor U1750 (N_1750,N_1410,N_1378);
or U1751 (N_1751,N_800,N_1189);
xnor U1752 (N_1752,N_1496,N_1419);
or U1753 (N_1753,N_1340,N_827);
xnor U1754 (N_1754,N_1498,N_1401);
nor U1755 (N_1755,N_1052,N_795);
nand U1756 (N_1756,N_1341,N_857);
and U1757 (N_1757,N_1000,N_752);
nand U1758 (N_1758,N_907,N_1295);
nor U1759 (N_1759,N_1230,N_940);
nor U1760 (N_1760,N_981,N_1202);
or U1761 (N_1761,N_1316,N_1284);
and U1762 (N_1762,N_813,N_1364);
nor U1763 (N_1763,N_1051,N_893);
nand U1764 (N_1764,N_1490,N_1021);
and U1765 (N_1765,N_1380,N_1130);
and U1766 (N_1766,N_1359,N_1418);
and U1767 (N_1767,N_1118,N_1294);
and U1768 (N_1768,N_1049,N_1053);
nand U1769 (N_1769,N_839,N_1306);
xor U1770 (N_1770,N_1011,N_1445);
nor U1771 (N_1771,N_1493,N_904);
and U1772 (N_1772,N_1323,N_858);
or U1773 (N_1773,N_1009,N_781);
nor U1774 (N_1774,N_1146,N_1333);
and U1775 (N_1775,N_1382,N_1239);
nor U1776 (N_1776,N_885,N_870);
nand U1777 (N_1777,N_1094,N_1088);
nand U1778 (N_1778,N_1024,N_906);
nor U1779 (N_1779,N_1241,N_872);
nand U1780 (N_1780,N_773,N_846);
nand U1781 (N_1781,N_1080,N_1328);
nand U1782 (N_1782,N_1220,N_1136);
or U1783 (N_1783,N_1172,N_1255);
nand U1784 (N_1784,N_853,N_880);
nand U1785 (N_1785,N_1057,N_1371);
or U1786 (N_1786,N_866,N_851);
and U1787 (N_1787,N_1070,N_1090);
nand U1788 (N_1788,N_1125,N_903);
nand U1789 (N_1789,N_1249,N_1280);
and U1790 (N_1790,N_825,N_1107);
and U1791 (N_1791,N_1180,N_1187);
nand U1792 (N_1792,N_996,N_1319);
nand U1793 (N_1793,N_1355,N_1483);
or U1794 (N_1794,N_929,N_1432);
xor U1795 (N_1795,N_1013,N_1204);
and U1796 (N_1796,N_1461,N_1353);
and U1797 (N_1797,N_1087,N_1339);
and U1798 (N_1798,N_937,N_1007);
nand U1799 (N_1799,N_844,N_799);
and U1800 (N_1800,N_1489,N_1076);
or U1801 (N_1801,N_1215,N_1446);
xnor U1802 (N_1802,N_1098,N_988);
or U1803 (N_1803,N_755,N_1326);
and U1804 (N_1804,N_1267,N_1479);
and U1805 (N_1805,N_1264,N_802);
nand U1806 (N_1806,N_1183,N_1092);
or U1807 (N_1807,N_966,N_1192);
and U1808 (N_1808,N_908,N_1307);
nand U1809 (N_1809,N_1375,N_1026);
and U1810 (N_1810,N_1038,N_983);
nand U1811 (N_1811,N_1001,N_1164);
or U1812 (N_1812,N_1086,N_970);
and U1813 (N_1813,N_1291,N_756);
nand U1814 (N_1814,N_1246,N_1143);
xor U1815 (N_1815,N_1167,N_841);
nand U1816 (N_1816,N_946,N_1436);
and U1817 (N_1817,N_901,N_1428);
or U1818 (N_1818,N_1305,N_896);
nand U1819 (N_1819,N_787,N_1096);
nand U1820 (N_1820,N_790,N_1058);
and U1821 (N_1821,N_1065,N_963);
xnor U1822 (N_1822,N_1356,N_1194);
nand U1823 (N_1823,N_1149,N_1083);
nand U1824 (N_1824,N_998,N_1393);
nor U1825 (N_1825,N_1151,N_1486);
and U1826 (N_1826,N_817,N_1031);
nand U1827 (N_1827,N_1434,N_1144);
and U1828 (N_1828,N_1429,N_1313);
nor U1829 (N_1829,N_910,N_1352);
and U1830 (N_1830,N_913,N_1234);
and U1831 (N_1831,N_1155,N_992);
or U1832 (N_1832,N_1250,N_1260);
and U1833 (N_1833,N_1309,N_753);
nand U1834 (N_1834,N_1389,N_1301);
or U1835 (N_1835,N_1129,N_995);
nand U1836 (N_1836,N_1458,N_1390);
or U1837 (N_1837,N_1236,N_982);
and U1838 (N_1838,N_999,N_1111);
nor U1839 (N_1839,N_1112,N_1036);
or U1840 (N_1840,N_835,N_1152);
or U1841 (N_1841,N_845,N_1050);
nor U1842 (N_1842,N_840,N_1258);
and U1843 (N_1843,N_1139,N_1370);
nand U1844 (N_1844,N_1400,N_1399);
nor U1845 (N_1845,N_902,N_895);
nand U1846 (N_1846,N_1229,N_881);
nand U1847 (N_1847,N_786,N_890);
and U1848 (N_1848,N_944,N_1261);
or U1849 (N_1849,N_819,N_1103);
and U1850 (N_1850,N_955,N_1140);
xor U1851 (N_1851,N_1269,N_792);
xnor U1852 (N_1852,N_912,N_1119);
xor U1853 (N_1853,N_886,N_927);
and U1854 (N_1854,N_1315,N_1037);
and U1855 (N_1855,N_862,N_821);
xor U1856 (N_1856,N_1318,N_1127);
and U1857 (N_1857,N_1174,N_977);
or U1858 (N_1858,N_1314,N_1005);
nand U1859 (N_1859,N_1408,N_1324);
or U1860 (N_1860,N_1073,N_1224);
or U1861 (N_1861,N_989,N_842);
and U1862 (N_1862,N_830,N_1279);
nor U1863 (N_1863,N_796,N_1335);
or U1864 (N_1864,N_1148,N_1265);
xor U1865 (N_1865,N_1292,N_959);
nor U1866 (N_1866,N_1421,N_1362);
or U1867 (N_1867,N_1200,N_814);
xnor U1868 (N_1868,N_915,N_1290);
nand U1869 (N_1869,N_1263,N_1081);
and U1870 (N_1870,N_1171,N_768);
or U1871 (N_1871,N_1181,N_1347);
or U1872 (N_1872,N_1067,N_849);
nor U1873 (N_1873,N_1444,N_1304);
and U1874 (N_1874,N_1030,N_1232);
nor U1875 (N_1875,N_1238,N_1384);
nor U1876 (N_1876,N_1242,N_1437);
or U1877 (N_1877,N_1136,N_1241);
or U1878 (N_1878,N_812,N_1275);
nand U1879 (N_1879,N_1110,N_1375);
xor U1880 (N_1880,N_1080,N_1250);
and U1881 (N_1881,N_1106,N_1380);
nor U1882 (N_1882,N_1080,N_893);
nor U1883 (N_1883,N_1243,N_1026);
nor U1884 (N_1884,N_1090,N_781);
nor U1885 (N_1885,N_948,N_1096);
nor U1886 (N_1886,N_999,N_992);
and U1887 (N_1887,N_971,N_1048);
nand U1888 (N_1888,N_1245,N_1483);
and U1889 (N_1889,N_779,N_1356);
nor U1890 (N_1890,N_834,N_812);
or U1891 (N_1891,N_867,N_1387);
nor U1892 (N_1892,N_1484,N_1276);
nor U1893 (N_1893,N_1341,N_902);
or U1894 (N_1894,N_881,N_758);
and U1895 (N_1895,N_888,N_753);
and U1896 (N_1896,N_1072,N_907);
nor U1897 (N_1897,N_1122,N_958);
nand U1898 (N_1898,N_1394,N_892);
nand U1899 (N_1899,N_1175,N_1466);
and U1900 (N_1900,N_1097,N_1027);
and U1901 (N_1901,N_1038,N_946);
or U1902 (N_1902,N_822,N_781);
and U1903 (N_1903,N_786,N_753);
nand U1904 (N_1904,N_1371,N_1049);
and U1905 (N_1905,N_1110,N_1062);
or U1906 (N_1906,N_937,N_958);
nand U1907 (N_1907,N_1464,N_1149);
or U1908 (N_1908,N_963,N_844);
and U1909 (N_1909,N_929,N_837);
or U1910 (N_1910,N_1209,N_1011);
nor U1911 (N_1911,N_827,N_753);
xor U1912 (N_1912,N_983,N_825);
nand U1913 (N_1913,N_950,N_1441);
or U1914 (N_1914,N_1291,N_1181);
or U1915 (N_1915,N_904,N_967);
and U1916 (N_1916,N_1144,N_868);
nor U1917 (N_1917,N_1442,N_1187);
nand U1918 (N_1918,N_1074,N_1171);
nand U1919 (N_1919,N_841,N_1362);
xor U1920 (N_1920,N_1251,N_1357);
and U1921 (N_1921,N_1373,N_1419);
xnor U1922 (N_1922,N_999,N_1367);
or U1923 (N_1923,N_1468,N_1099);
nor U1924 (N_1924,N_1172,N_989);
nand U1925 (N_1925,N_896,N_1074);
and U1926 (N_1926,N_1069,N_1000);
and U1927 (N_1927,N_1373,N_785);
nand U1928 (N_1928,N_762,N_764);
nand U1929 (N_1929,N_1021,N_1062);
nor U1930 (N_1930,N_1390,N_1284);
nor U1931 (N_1931,N_1207,N_826);
or U1932 (N_1932,N_1209,N_1095);
nor U1933 (N_1933,N_1432,N_1257);
nor U1934 (N_1934,N_1173,N_1168);
nor U1935 (N_1935,N_1293,N_1441);
xor U1936 (N_1936,N_1230,N_1472);
and U1937 (N_1937,N_968,N_1190);
or U1938 (N_1938,N_1138,N_1085);
nand U1939 (N_1939,N_1293,N_1124);
and U1940 (N_1940,N_1397,N_986);
nor U1941 (N_1941,N_1443,N_1036);
nor U1942 (N_1942,N_1375,N_1228);
and U1943 (N_1943,N_1460,N_1453);
and U1944 (N_1944,N_1023,N_1346);
and U1945 (N_1945,N_912,N_887);
and U1946 (N_1946,N_1361,N_1113);
nand U1947 (N_1947,N_1202,N_1335);
nand U1948 (N_1948,N_1183,N_1220);
nor U1949 (N_1949,N_1476,N_1367);
or U1950 (N_1950,N_1305,N_879);
nor U1951 (N_1951,N_1007,N_903);
or U1952 (N_1952,N_971,N_904);
xor U1953 (N_1953,N_910,N_1019);
nand U1954 (N_1954,N_818,N_1431);
or U1955 (N_1955,N_930,N_1425);
xnor U1956 (N_1956,N_1319,N_780);
and U1957 (N_1957,N_1231,N_806);
xor U1958 (N_1958,N_1422,N_956);
nand U1959 (N_1959,N_1490,N_968);
and U1960 (N_1960,N_1334,N_1038);
and U1961 (N_1961,N_970,N_1043);
nand U1962 (N_1962,N_1153,N_1259);
or U1963 (N_1963,N_1156,N_1254);
or U1964 (N_1964,N_1057,N_1027);
and U1965 (N_1965,N_1335,N_1331);
or U1966 (N_1966,N_1467,N_1265);
and U1967 (N_1967,N_1430,N_1388);
xnor U1968 (N_1968,N_1237,N_829);
xor U1969 (N_1969,N_1404,N_1279);
nor U1970 (N_1970,N_1023,N_920);
or U1971 (N_1971,N_953,N_1266);
or U1972 (N_1972,N_1032,N_1219);
nand U1973 (N_1973,N_935,N_1283);
or U1974 (N_1974,N_800,N_1293);
nand U1975 (N_1975,N_1301,N_1247);
nand U1976 (N_1976,N_1411,N_1245);
nor U1977 (N_1977,N_790,N_1259);
nand U1978 (N_1978,N_1467,N_1001);
nand U1979 (N_1979,N_1177,N_1202);
or U1980 (N_1980,N_938,N_966);
and U1981 (N_1981,N_1254,N_974);
and U1982 (N_1982,N_967,N_766);
or U1983 (N_1983,N_1081,N_1000);
or U1984 (N_1984,N_1410,N_806);
and U1985 (N_1985,N_1331,N_1393);
or U1986 (N_1986,N_1040,N_1086);
or U1987 (N_1987,N_1225,N_1261);
nand U1988 (N_1988,N_985,N_1244);
or U1989 (N_1989,N_808,N_810);
nor U1990 (N_1990,N_1496,N_1392);
or U1991 (N_1991,N_1003,N_1152);
or U1992 (N_1992,N_997,N_1435);
nand U1993 (N_1993,N_1355,N_1225);
nand U1994 (N_1994,N_1495,N_1160);
or U1995 (N_1995,N_1148,N_1154);
and U1996 (N_1996,N_1417,N_833);
and U1997 (N_1997,N_926,N_775);
and U1998 (N_1998,N_903,N_1264);
and U1999 (N_1999,N_1439,N_937);
nand U2000 (N_2000,N_1144,N_943);
and U2001 (N_2001,N_1197,N_1133);
and U2002 (N_2002,N_1451,N_1360);
nand U2003 (N_2003,N_1308,N_1332);
nor U2004 (N_2004,N_896,N_1399);
xnor U2005 (N_2005,N_753,N_957);
xnor U2006 (N_2006,N_757,N_819);
xor U2007 (N_2007,N_1328,N_1403);
nand U2008 (N_2008,N_989,N_1039);
or U2009 (N_2009,N_1421,N_1451);
and U2010 (N_2010,N_1205,N_987);
nor U2011 (N_2011,N_803,N_796);
nand U2012 (N_2012,N_758,N_1252);
nand U2013 (N_2013,N_779,N_1012);
nand U2014 (N_2014,N_1228,N_1125);
and U2015 (N_2015,N_987,N_1184);
or U2016 (N_2016,N_1443,N_1339);
and U2017 (N_2017,N_1345,N_1384);
and U2018 (N_2018,N_1403,N_1072);
and U2019 (N_2019,N_1429,N_1195);
or U2020 (N_2020,N_1218,N_1407);
xnor U2021 (N_2021,N_1099,N_755);
and U2022 (N_2022,N_1367,N_1020);
xnor U2023 (N_2023,N_1440,N_939);
nand U2024 (N_2024,N_1379,N_1014);
and U2025 (N_2025,N_1306,N_1467);
xor U2026 (N_2026,N_850,N_1416);
nor U2027 (N_2027,N_903,N_967);
nand U2028 (N_2028,N_861,N_1017);
nor U2029 (N_2029,N_1269,N_1046);
or U2030 (N_2030,N_1199,N_961);
and U2031 (N_2031,N_966,N_774);
nor U2032 (N_2032,N_1297,N_1060);
and U2033 (N_2033,N_1456,N_1065);
nand U2034 (N_2034,N_1164,N_928);
and U2035 (N_2035,N_839,N_772);
nand U2036 (N_2036,N_758,N_1427);
or U2037 (N_2037,N_1165,N_1394);
or U2038 (N_2038,N_797,N_800);
and U2039 (N_2039,N_1273,N_1153);
nand U2040 (N_2040,N_1374,N_982);
nor U2041 (N_2041,N_1474,N_1062);
nor U2042 (N_2042,N_1192,N_986);
and U2043 (N_2043,N_777,N_1347);
nor U2044 (N_2044,N_936,N_819);
or U2045 (N_2045,N_1225,N_869);
nor U2046 (N_2046,N_1203,N_775);
nor U2047 (N_2047,N_1461,N_1331);
and U2048 (N_2048,N_1321,N_860);
nor U2049 (N_2049,N_839,N_943);
or U2050 (N_2050,N_1036,N_794);
and U2051 (N_2051,N_855,N_790);
nand U2052 (N_2052,N_1184,N_832);
and U2053 (N_2053,N_982,N_1382);
xnor U2054 (N_2054,N_1464,N_1347);
nor U2055 (N_2055,N_1497,N_1380);
or U2056 (N_2056,N_1368,N_1124);
nand U2057 (N_2057,N_775,N_1408);
xor U2058 (N_2058,N_804,N_962);
nand U2059 (N_2059,N_1032,N_1495);
or U2060 (N_2060,N_985,N_984);
nor U2061 (N_2061,N_1395,N_1460);
or U2062 (N_2062,N_1109,N_1280);
nand U2063 (N_2063,N_991,N_884);
and U2064 (N_2064,N_1341,N_1489);
nand U2065 (N_2065,N_1051,N_916);
nor U2066 (N_2066,N_1166,N_808);
or U2067 (N_2067,N_1325,N_955);
nand U2068 (N_2068,N_842,N_1053);
nor U2069 (N_2069,N_755,N_1162);
nand U2070 (N_2070,N_875,N_1446);
nand U2071 (N_2071,N_1128,N_1357);
xor U2072 (N_2072,N_1140,N_1399);
nand U2073 (N_2073,N_886,N_1388);
xor U2074 (N_2074,N_1274,N_1414);
and U2075 (N_2075,N_844,N_835);
and U2076 (N_2076,N_803,N_1400);
nor U2077 (N_2077,N_1021,N_751);
nor U2078 (N_2078,N_1192,N_814);
nor U2079 (N_2079,N_1256,N_1367);
nand U2080 (N_2080,N_1384,N_1148);
or U2081 (N_2081,N_789,N_1239);
nand U2082 (N_2082,N_1442,N_828);
nand U2083 (N_2083,N_803,N_1385);
and U2084 (N_2084,N_1037,N_1471);
and U2085 (N_2085,N_1275,N_1155);
nand U2086 (N_2086,N_1403,N_891);
or U2087 (N_2087,N_924,N_847);
or U2088 (N_2088,N_844,N_1053);
nor U2089 (N_2089,N_1371,N_1292);
or U2090 (N_2090,N_1128,N_955);
nand U2091 (N_2091,N_1406,N_785);
or U2092 (N_2092,N_1150,N_1167);
or U2093 (N_2093,N_1017,N_905);
nand U2094 (N_2094,N_1152,N_837);
nand U2095 (N_2095,N_1116,N_1403);
nor U2096 (N_2096,N_1251,N_936);
nand U2097 (N_2097,N_896,N_1057);
xor U2098 (N_2098,N_1320,N_965);
nand U2099 (N_2099,N_1011,N_1435);
or U2100 (N_2100,N_1433,N_1229);
nand U2101 (N_2101,N_1153,N_1282);
and U2102 (N_2102,N_799,N_1148);
xnor U2103 (N_2103,N_1358,N_1109);
or U2104 (N_2104,N_994,N_931);
or U2105 (N_2105,N_1091,N_1023);
nand U2106 (N_2106,N_1196,N_1152);
nor U2107 (N_2107,N_960,N_1289);
or U2108 (N_2108,N_827,N_1464);
and U2109 (N_2109,N_1221,N_1246);
nor U2110 (N_2110,N_985,N_936);
nor U2111 (N_2111,N_1420,N_809);
nand U2112 (N_2112,N_1300,N_777);
nor U2113 (N_2113,N_1320,N_754);
xnor U2114 (N_2114,N_773,N_1047);
nand U2115 (N_2115,N_1277,N_879);
or U2116 (N_2116,N_1170,N_1352);
nand U2117 (N_2117,N_1136,N_1316);
nand U2118 (N_2118,N_940,N_929);
nand U2119 (N_2119,N_1048,N_1388);
nor U2120 (N_2120,N_754,N_786);
nand U2121 (N_2121,N_867,N_1369);
nand U2122 (N_2122,N_1196,N_955);
nor U2123 (N_2123,N_1061,N_1290);
nand U2124 (N_2124,N_1140,N_992);
nand U2125 (N_2125,N_1099,N_817);
and U2126 (N_2126,N_1408,N_955);
xor U2127 (N_2127,N_1089,N_1179);
or U2128 (N_2128,N_1383,N_1405);
nor U2129 (N_2129,N_1019,N_1199);
or U2130 (N_2130,N_1441,N_943);
nor U2131 (N_2131,N_1152,N_887);
nor U2132 (N_2132,N_1446,N_1491);
nand U2133 (N_2133,N_1429,N_1406);
or U2134 (N_2134,N_1265,N_1212);
or U2135 (N_2135,N_863,N_847);
xor U2136 (N_2136,N_787,N_896);
nor U2137 (N_2137,N_1412,N_1461);
nor U2138 (N_2138,N_1326,N_1201);
and U2139 (N_2139,N_1311,N_1332);
nor U2140 (N_2140,N_1180,N_768);
nand U2141 (N_2141,N_1075,N_1230);
and U2142 (N_2142,N_1204,N_1109);
nor U2143 (N_2143,N_1029,N_1269);
nor U2144 (N_2144,N_970,N_1390);
or U2145 (N_2145,N_1488,N_856);
or U2146 (N_2146,N_1155,N_1165);
nor U2147 (N_2147,N_1283,N_1037);
and U2148 (N_2148,N_1490,N_1124);
nor U2149 (N_2149,N_1499,N_1367);
nand U2150 (N_2150,N_764,N_1113);
and U2151 (N_2151,N_1153,N_1454);
or U2152 (N_2152,N_1494,N_1379);
xnor U2153 (N_2153,N_1323,N_1387);
and U2154 (N_2154,N_1015,N_1183);
or U2155 (N_2155,N_863,N_800);
nor U2156 (N_2156,N_784,N_1095);
xnor U2157 (N_2157,N_974,N_1092);
and U2158 (N_2158,N_1150,N_1105);
and U2159 (N_2159,N_1116,N_1359);
nand U2160 (N_2160,N_1254,N_986);
and U2161 (N_2161,N_1338,N_1314);
xnor U2162 (N_2162,N_806,N_1439);
or U2163 (N_2163,N_1086,N_974);
nand U2164 (N_2164,N_1145,N_926);
or U2165 (N_2165,N_939,N_903);
and U2166 (N_2166,N_1327,N_941);
or U2167 (N_2167,N_1015,N_1056);
nand U2168 (N_2168,N_1294,N_931);
or U2169 (N_2169,N_1198,N_1395);
nor U2170 (N_2170,N_1042,N_1137);
and U2171 (N_2171,N_1337,N_1433);
and U2172 (N_2172,N_846,N_1434);
nand U2173 (N_2173,N_1356,N_1130);
and U2174 (N_2174,N_818,N_1097);
nor U2175 (N_2175,N_905,N_1496);
xnor U2176 (N_2176,N_1054,N_1239);
or U2177 (N_2177,N_1407,N_1498);
nand U2178 (N_2178,N_1436,N_1388);
and U2179 (N_2179,N_1236,N_905);
nand U2180 (N_2180,N_863,N_1157);
and U2181 (N_2181,N_1338,N_1405);
nor U2182 (N_2182,N_1030,N_1159);
or U2183 (N_2183,N_778,N_1300);
and U2184 (N_2184,N_914,N_1218);
and U2185 (N_2185,N_1396,N_1240);
and U2186 (N_2186,N_1242,N_1003);
and U2187 (N_2187,N_1228,N_1062);
and U2188 (N_2188,N_750,N_1240);
nand U2189 (N_2189,N_1400,N_945);
and U2190 (N_2190,N_903,N_1140);
and U2191 (N_2191,N_1137,N_891);
and U2192 (N_2192,N_1493,N_775);
nand U2193 (N_2193,N_1036,N_1139);
or U2194 (N_2194,N_990,N_1298);
nand U2195 (N_2195,N_1037,N_1495);
or U2196 (N_2196,N_1216,N_1382);
or U2197 (N_2197,N_1241,N_982);
nand U2198 (N_2198,N_1163,N_879);
and U2199 (N_2199,N_1407,N_978);
nor U2200 (N_2200,N_1286,N_1322);
nor U2201 (N_2201,N_1173,N_1304);
and U2202 (N_2202,N_943,N_829);
xor U2203 (N_2203,N_773,N_809);
nand U2204 (N_2204,N_782,N_1447);
nor U2205 (N_2205,N_1320,N_1339);
or U2206 (N_2206,N_932,N_1330);
or U2207 (N_2207,N_1169,N_981);
nor U2208 (N_2208,N_983,N_1175);
and U2209 (N_2209,N_856,N_1082);
and U2210 (N_2210,N_880,N_885);
nor U2211 (N_2211,N_1396,N_860);
nor U2212 (N_2212,N_1368,N_979);
nor U2213 (N_2213,N_779,N_1289);
or U2214 (N_2214,N_1233,N_1070);
or U2215 (N_2215,N_1350,N_852);
or U2216 (N_2216,N_1281,N_828);
nor U2217 (N_2217,N_1320,N_1396);
and U2218 (N_2218,N_1198,N_1314);
xor U2219 (N_2219,N_770,N_1344);
nand U2220 (N_2220,N_1014,N_949);
xnor U2221 (N_2221,N_1447,N_961);
and U2222 (N_2222,N_1321,N_1151);
xnor U2223 (N_2223,N_910,N_791);
and U2224 (N_2224,N_929,N_993);
nand U2225 (N_2225,N_793,N_1194);
xnor U2226 (N_2226,N_962,N_1367);
and U2227 (N_2227,N_789,N_1311);
nor U2228 (N_2228,N_1279,N_914);
nor U2229 (N_2229,N_869,N_1167);
nand U2230 (N_2230,N_1485,N_840);
nor U2231 (N_2231,N_1194,N_1240);
nor U2232 (N_2232,N_1185,N_1040);
nor U2233 (N_2233,N_997,N_1109);
and U2234 (N_2234,N_1313,N_1297);
or U2235 (N_2235,N_1113,N_1181);
xnor U2236 (N_2236,N_852,N_1088);
or U2237 (N_2237,N_882,N_762);
and U2238 (N_2238,N_975,N_784);
or U2239 (N_2239,N_1443,N_1042);
nor U2240 (N_2240,N_760,N_928);
nor U2241 (N_2241,N_1074,N_1484);
nor U2242 (N_2242,N_910,N_901);
and U2243 (N_2243,N_1119,N_1063);
xnor U2244 (N_2244,N_1296,N_856);
or U2245 (N_2245,N_1093,N_1068);
nor U2246 (N_2246,N_934,N_1176);
nand U2247 (N_2247,N_970,N_1406);
or U2248 (N_2248,N_951,N_1091);
nand U2249 (N_2249,N_844,N_814);
and U2250 (N_2250,N_1955,N_1899);
nand U2251 (N_2251,N_2220,N_1858);
or U2252 (N_2252,N_1882,N_1799);
or U2253 (N_2253,N_1838,N_2125);
nand U2254 (N_2254,N_1522,N_2203);
nor U2255 (N_2255,N_2093,N_1632);
nand U2256 (N_2256,N_1631,N_1897);
xor U2257 (N_2257,N_1728,N_1788);
nor U2258 (N_2258,N_1571,N_2242);
nor U2259 (N_2259,N_1677,N_2191);
xnor U2260 (N_2260,N_1873,N_1576);
nand U2261 (N_2261,N_2235,N_1626);
nor U2262 (N_2262,N_1640,N_2034);
or U2263 (N_2263,N_1768,N_1989);
nand U2264 (N_2264,N_1525,N_1773);
or U2265 (N_2265,N_1692,N_1660);
nor U2266 (N_2266,N_1560,N_2150);
or U2267 (N_2267,N_2067,N_1961);
nand U2268 (N_2268,N_2101,N_1974);
nor U2269 (N_2269,N_1709,N_2082);
or U2270 (N_2270,N_2192,N_1988);
and U2271 (N_2271,N_1934,N_2176);
or U2272 (N_2272,N_1745,N_1545);
or U2273 (N_2273,N_2048,N_1703);
and U2274 (N_2274,N_1654,N_2142);
nand U2275 (N_2275,N_2092,N_1732);
nor U2276 (N_2276,N_2062,N_2043);
nor U2277 (N_2277,N_1714,N_1985);
nand U2278 (N_2278,N_1859,N_1887);
or U2279 (N_2279,N_1509,N_1785);
nand U2280 (N_2280,N_2061,N_1845);
nor U2281 (N_2281,N_2181,N_1592);
nand U2282 (N_2282,N_2066,N_1796);
nor U2283 (N_2283,N_1972,N_1963);
or U2284 (N_2284,N_1754,N_1682);
and U2285 (N_2285,N_1551,N_2204);
nand U2286 (N_2286,N_1952,N_1621);
and U2287 (N_2287,N_2124,N_1673);
and U2288 (N_2288,N_2033,N_1958);
nor U2289 (N_2289,N_1968,N_1615);
nor U2290 (N_2290,N_1751,N_1526);
xor U2291 (N_2291,N_1618,N_1720);
and U2292 (N_2292,N_1800,N_1775);
or U2293 (N_2293,N_1715,N_2106);
or U2294 (N_2294,N_2017,N_2076);
nor U2295 (N_2295,N_2073,N_1794);
and U2296 (N_2296,N_1717,N_1835);
xor U2297 (N_2297,N_1512,N_2196);
and U2298 (N_2298,N_1916,N_1574);
nor U2299 (N_2299,N_1726,N_1550);
nand U2300 (N_2300,N_1605,N_1774);
or U2301 (N_2301,N_2223,N_1687);
nand U2302 (N_2302,N_2138,N_1929);
nand U2303 (N_2303,N_1661,N_2208);
or U2304 (N_2304,N_1757,N_2098);
nand U2305 (N_2305,N_1834,N_1538);
nand U2306 (N_2306,N_2039,N_1824);
xor U2307 (N_2307,N_1601,N_2221);
nor U2308 (N_2308,N_1613,N_1639);
or U2309 (N_2309,N_1847,N_1894);
nand U2310 (N_2310,N_2108,N_1623);
and U2311 (N_2311,N_2209,N_1539);
and U2312 (N_2312,N_2162,N_1875);
or U2313 (N_2313,N_1888,N_1826);
or U2314 (N_2314,N_1884,N_1575);
or U2315 (N_2315,N_1561,N_1619);
nand U2316 (N_2316,N_1765,N_1832);
xnor U2317 (N_2317,N_1595,N_1827);
nand U2318 (N_2318,N_2238,N_1579);
and U2319 (N_2319,N_1914,N_2128);
or U2320 (N_2320,N_1542,N_1516);
or U2321 (N_2321,N_2083,N_1635);
nor U2322 (N_2322,N_1904,N_1982);
or U2323 (N_2323,N_1948,N_1992);
and U2324 (N_2324,N_2074,N_2240);
and U2325 (N_2325,N_1998,N_1655);
and U2326 (N_2326,N_1762,N_1685);
nand U2327 (N_2327,N_2031,N_2040);
nand U2328 (N_2328,N_1636,N_1730);
or U2329 (N_2329,N_1721,N_2207);
or U2330 (N_2330,N_2236,N_1851);
nand U2331 (N_2331,N_1840,N_1764);
or U2332 (N_2332,N_1846,N_2072);
nor U2333 (N_2333,N_2079,N_2111);
nor U2334 (N_2334,N_1849,N_1686);
and U2335 (N_2335,N_1528,N_1920);
nand U2336 (N_2336,N_2174,N_1722);
or U2337 (N_2337,N_1783,N_1602);
and U2338 (N_2338,N_2117,N_2152);
nor U2339 (N_2339,N_1710,N_1776);
xnor U2340 (N_2340,N_1706,N_1587);
and U2341 (N_2341,N_1688,N_2244);
xor U2342 (N_2342,N_1848,N_1557);
and U2343 (N_2343,N_1928,N_1629);
nand U2344 (N_2344,N_1801,N_1986);
and U2345 (N_2345,N_2112,N_1809);
or U2346 (N_2346,N_1637,N_1674);
xor U2347 (N_2347,N_1867,N_2032);
nand U2348 (N_2348,N_1570,N_2064);
nor U2349 (N_2349,N_1535,N_1970);
nand U2350 (N_2350,N_1918,N_2171);
and U2351 (N_2351,N_1877,N_1964);
and U2352 (N_2352,N_1907,N_1939);
nand U2353 (N_2353,N_1979,N_2219);
or U2354 (N_2354,N_2087,N_1584);
nand U2355 (N_2355,N_1962,N_2179);
nand U2356 (N_2356,N_2049,N_2089);
nor U2357 (N_2357,N_1508,N_2164);
nand U2358 (N_2358,N_1777,N_1871);
nor U2359 (N_2359,N_2183,N_1506);
or U2360 (N_2360,N_1811,N_2206);
nor U2361 (N_2361,N_2055,N_1523);
or U2362 (N_2362,N_1944,N_1564);
nor U2363 (N_2363,N_1905,N_1500);
nand U2364 (N_2364,N_1903,N_1759);
nor U2365 (N_2365,N_1747,N_1781);
and U2366 (N_2366,N_2218,N_2188);
or U2367 (N_2367,N_1742,N_2044);
nor U2368 (N_2368,N_1924,N_1643);
or U2369 (N_2369,N_1900,N_1828);
nor U2370 (N_2370,N_1702,N_1942);
nand U2371 (N_2371,N_1633,N_2146);
nor U2372 (N_2372,N_1779,N_2160);
and U2373 (N_2373,N_2140,N_1855);
nand U2374 (N_2374,N_1530,N_1559);
and U2375 (N_2375,N_1960,N_2195);
nand U2376 (N_2376,N_1701,N_1541);
and U2377 (N_2377,N_2145,N_2038);
nand U2378 (N_2378,N_2161,N_1567);
nand U2379 (N_2379,N_1980,N_2009);
nand U2380 (N_2380,N_1863,N_2025);
xor U2381 (N_2381,N_2151,N_1708);
or U2382 (N_2382,N_1868,N_1667);
nand U2383 (N_2383,N_1969,N_1983);
nand U2384 (N_2384,N_1933,N_2080);
nand U2385 (N_2385,N_2222,N_1610);
nand U2386 (N_2386,N_2132,N_2027);
nor U2387 (N_2387,N_1735,N_1596);
nand U2388 (N_2388,N_1698,N_1756);
or U2389 (N_2389,N_1861,N_1895);
nand U2390 (N_2390,N_1505,N_1566);
or U2391 (N_2391,N_1893,N_1598);
and U2392 (N_2392,N_1513,N_1681);
and U2393 (N_2393,N_1780,N_1693);
or U2394 (N_2394,N_2156,N_1825);
nor U2395 (N_2395,N_2109,N_1733);
or U2396 (N_2396,N_1691,N_2028);
nand U2397 (N_2397,N_1731,N_1938);
and U2398 (N_2398,N_1634,N_1556);
nand U2399 (N_2399,N_1608,N_1786);
and U2400 (N_2400,N_1886,N_1880);
nor U2401 (N_2401,N_1600,N_1977);
and U2402 (N_2402,N_1750,N_1752);
or U2403 (N_2403,N_1727,N_1614);
and U2404 (N_2404,N_2078,N_2126);
or U2405 (N_2405,N_1519,N_1588);
or U2406 (N_2406,N_1529,N_2154);
nand U2407 (N_2407,N_1946,N_2190);
xnor U2408 (N_2408,N_1767,N_2201);
nand U2409 (N_2409,N_2029,N_1669);
xor U2410 (N_2410,N_2205,N_1902);
nor U2411 (N_2411,N_1625,N_1548);
and U2412 (N_2412,N_1737,N_1606);
and U2413 (N_2413,N_2100,N_2229);
nand U2414 (N_2414,N_1864,N_1740);
or U2415 (N_2415,N_2001,N_2070);
or U2416 (N_2416,N_1707,N_2051);
nor U2417 (N_2417,N_2042,N_1844);
or U2418 (N_2418,N_1736,N_1531);
and U2419 (N_2419,N_2099,N_1911);
nor U2420 (N_2420,N_1947,N_1568);
nand U2421 (N_2421,N_2011,N_2130);
and U2422 (N_2422,N_1760,N_1990);
nor U2423 (N_2423,N_2157,N_1791);
nand U2424 (N_2424,N_1951,N_1976);
nand U2425 (N_2425,N_1872,N_1883);
nand U2426 (N_2426,N_1697,N_1926);
nor U2427 (N_2427,N_2135,N_2212);
or U2428 (N_2428,N_1581,N_2050);
nand U2429 (N_2429,N_1815,N_1547);
nor U2430 (N_2430,N_1622,N_1569);
and U2431 (N_2431,N_1603,N_1890);
and U2432 (N_2432,N_2008,N_2063);
nand U2433 (N_2433,N_2088,N_1803);
nor U2434 (N_2434,N_1975,N_2006);
nand U2435 (N_2435,N_1954,N_1843);
nor U2436 (N_2436,N_1790,N_1689);
nand U2437 (N_2437,N_1941,N_1554);
or U2438 (N_2438,N_2184,N_1818);
nand U2439 (N_2439,N_1782,N_1544);
nand U2440 (N_2440,N_1819,N_1758);
nor U2441 (N_2441,N_2210,N_1833);
and U2442 (N_2442,N_2081,N_1922);
xor U2443 (N_2443,N_1578,N_2211);
and U2444 (N_2444,N_1841,N_1789);
nor U2445 (N_2445,N_2185,N_2041);
and U2446 (N_2446,N_2000,N_1562);
nor U2447 (N_2447,N_2148,N_1769);
nor U2448 (N_2448,N_1668,N_1604);
or U2449 (N_2449,N_2246,N_1919);
or U2450 (N_2450,N_2169,N_2232);
nor U2451 (N_2451,N_2247,N_1766);
nor U2452 (N_2452,N_1662,N_1869);
nor U2453 (N_2453,N_2077,N_1741);
or U2454 (N_2454,N_1593,N_1937);
nand U2455 (N_2455,N_1532,N_2086);
and U2456 (N_2456,N_1599,N_1684);
xor U2457 (N_2457,N_1949,N_1664);
or U2458 (N_2458,N_2075,N_1549);
xnor U2459 (N_2459,N_1704,N_1837);
nand U2460 (N_2460,N_2186,N_2180);
nor U2461 (N_2461,N_1514,N_1906);
nor U2462 (N_2462,N_2230,N_1797);
nor U2463 (N_2463,N_1573,N_2141);
and U2464 (N_2464,N_1738,N_1582);
nand U2465 (N_2465,N_2239,N_1812);
or U2466 (N_2466,N_2199,N_2052);
nand U2467 (N_2467,N_2013,N_1945);
nand U2468 (N_2468,N_1817,N_1744);
nor U2469 (N_2469,N_2143,N_2133);
xor U2470 (N_2470,N_1795,N_1925);
nor U2471 (N_2471,N_1718,N_1950);
nand U2472 (N_2472,N_1874,N_1694);
or U2473 (N_2473,N_1908,N_2022);
or U2474 (N_2474,N_1829,N_2007);
or U2475 (N_2475,N_1679,N_1555);
nand U2476 (N_2476,N_2163,N_1638);
or U2477 (N_2477,N_1746,N_2026);
nand U2478 (N_2478,N_1690,N_1839);
xor U2479 (N_2479,N_1870,N_2149);
and U2480 (N_2480,N_1991,N_1713);
or U2481 (N_2481,N_2134,N_1889);
or U2482 (N_2482,N_1763,N_2095);
and U2483 (N_2483,N_2037,N_1719);
nor U2484 (N_2484,N_1808,N_2019);
and U2485 (N_2485,N_1898,N_1771);
nor U2486 (N_2486,N_1778,N_2094);
and U2487 (N_2487,N_1927,N_1973);
nor U2488 (N_2488,N_1607,N_2147);
nand U2489 (N_2489,N_1611,N_1915);
xnor U2490 (N_2490,N_1725,N_1862);
xnor U2491 (N_2491,N_1540,N_1501);
nor U2492 (N_2492,N_1616,N_1770);
xor U2493 (N_2493,N_1802,N_2241);
xnor U2494 (N_2494,N_1642,N_1935);
and U2495 (N_2495,N_1565,N_2053);
or U2496 (N_2496,N_1987,N_2137);
nand U2497 (N_2497,N_2036,N_1931);
nand U2498 (N_2498,N_2168,N_1749);
nor U2499 (N_2499,N_1936,N_1683);
and U2500 (N_2500,N_1813,N_1806);
nand U2501 (N_2501,N_1617,N_1881);
nand U2502 (N_2502,N_2194,N_2096);
and U2503 (N_2503,N_1537,N_2198);
xor U2504 (N_2504,N_2228,N_1892);
or U2505 (N_2505,N_1511,N_2159);
nor U2506 (N_2506,N_1836,N_1663);
nor U2507 (N_2507,N_1820,N_1504);
nor U2508 (N_2508,N_2123,N_2131);
or U2509 (N_2509,N_1711,N_2003);
and U2510 (N_2510,N_1739,N_1930);
nand U2511 (N_2511,N_1517,N_2226);
nor U2512 (N_2512,N_1648,N_1659);
nand U2513 (N_2513,N_2177,N_1885);
or U2514 (N_2514,N_1995,N_1502);
and U2515 (N_2515,N_1999,N_1705);
and U2516 (N_2516,N_1628,N_2097);
nand U2517 (N_2517,N_2237,N_2139);
and U2518 (N_2518,N_1563,N_1695);
or U2519 (N_2519,N_2016,N_1657);
nand U2520 (N_2520,N_2107,N_2213);
or U2521 (N_2521,N_1647,N_1901);
or U2522 (N_2522,N_1856,N_2058);
nor U2523 (N_2523,N_2113,N_1981);
and U2524 (N_2524,N_1850,N_1804);
and U2525 (N_2525,N_2021,N_1787);
nor U2526 (N_2526,N_1723,N_1965);
xnor U2527 (N_2527,N_2002,N_1696);
nor U2528 (N_2528,N_1743,N_1585);
or U2529 (N_2529,N_1821,N_2224);
or U2530 (N_2530,N_1503,N_2122);
or U2531 (N_2531,N_1921,N_2071);
nor U2532 (N_2532,N_1580,N_2182);
and U2533 (N_2533,N_1993,N_1597);
nand U2534 (N_2534,N_2090,N_1822);
or U2535 (N_2535,N_1755,N_1645);
and U2536 (N_2536,N_2172,N_2118);
nor U2537 (N_2537,N_1805,N_2010);
nor U2538 (N_2538,N_1997,N_1807);
and U2539 (N_2539,N_2018,N_1671);
and U2540 (N_2540,N_1876,N_2173);
xor U2541 (N_2541,N_1543,N_2069);
and U2542 (N_2542,N_1665,N_1798);
or U2543 (N_2543,N_1641,N_1957);
and U2544 (N_2544,N_2103,N_1854);
and U2545 (N_2545,N_1609,N_2120);
xor U2546 (N_2546,N_1912,N_1699);
and U2547 (N_2547,N_2119,N_1831);
and U2548 (N_2548,N_1510,N_1910);
nand U2549 (N_2549,N_1956,N_1646);
or U2550 (N_2550,N_1761,N_1984);
nor U2551 (N_2551,N_1577,N_2158);
nand U2552 (N_2552,N_1594,N_2065);
or U2553 (N_2553,N_1830,N_2248);
nor U2554 (N_2554,N_2155,N_1524);
and U2555 (N_2555,N_2129,N_2054);
or U2556 (N_2556,N_2202,N_1670);
nand U2557 (N_2557,N_1913,N_1966);
nor U2558 (N_2558,N_2102,N_1729);
xnor U2559 (N_2559,N_1612,N_1959);
and U2560 (N_2560,N_1515,N_1932);
and U2561 (N_2561,N_2170,N_1656);
nand U2562 (N_2562,N_2193,N_1630);
nor U2563 (N_2563,N_1590,N_1649);
nand U2564 (N_2564,N_1734,N_1680);
and U2565 (N_2565,N_1852,N_2200);
nor U2566 (N_2566,N_2047,N_1586);
and U2567 (N_2567,N_1534,N_1784);
nand U2568 (N_2568,N_1520,N_2127);
nand U2569 (N_2569,N_2114,N_1996);
nand U2570 (N_2570,N_1521,N_2175);
or U2571 (N_2571,N_1823,N_2023);
and U2572 (N_2572,N_2187,N_2216);
xnor U2573 (N_2573,N_2215,N_2105);
nand U2574 (N_2574,N_2046,N_1940);
or U2575 (N_2575,N_1971,N_1572);
nor U2576 (N_2576,N_2012,N_1792);
nor U2577 (N_2577,N_1917,N_1860);
nand U2578 (N_2578,N_2243,N_1878);
nand U2579 (N_2579,N_1658,N_2004);
or U2580 (N_2580,N_1943,N_1712);
xor U2581 (N_2581,N_2136,N_1650);
and U2582 (N_2582,N_2110,N_1978);
xnor U2583 (N_2583,N_1624,N_2189);
or U2584 (N_2584,N_1953,N_2085);
or U2585 (N_2585,N_2104,N_2056);
nor U2586 (N_2586,N_2144,N_2153);
and U2587 (N_2587,N_1552,N_2084);
nand U2588 (N_2588,N_2015,N_1967);
and U2589 (N_2589,N_1810,N_2059);
and U2590 (N_2590,N_1536,N_1620);
nand U2591 (N_2591,N_1652,N_1627);
or U2592 (N_2592,N_1546,N_1842);
or U2593 (N_2593,N_1866,N_1716);
nand U2594 (N_2594,N_1644,N_1676);
xor U2595 (N_2595,N_2057,N_1651);
and U2596 (N_2596,N_2167,N_1558);
nor U2597 (N_2597,N_2245,N_1753);
nand U2598 (N_2598,N_2014,N_1793);
nand U2599 (N_2599,N_1816,N_1748);
and U2600 (N_2600,N_2024,N_1923);
nand U2601 (N_2601,N_1675,N_2116);
nand U2602 (N_2602,N_2234,N_1583);
and U2603 (N_2603,N_1896,N_1994);
or U2604 (N_2604,N_1533,N_1589);
nand U2605 (N_2605,N_2227,N_1591);
and U2606 (N_2606,N_2233,N_1879);
nor U2607 (N_2607,N_1853,N_1909);
nor U2608 (N_2608,N_2060,N_2091);
and U2609 (N_2609,N_1891,N_1865);
or U2610 (N_2610,N_2068,N_2249);
and U2611 (N_2611,N_2231,N_1772);
nand U2612 (N_2612,N_2020,N_1653);
nand U2613 (N_2613,N_2121,N_2214);
and U2614 (N_2614,N_2197,N_2166);
and U2615 (N_2615,N_2178,N_2225);
nand U2616 (N_2616,N_2005,N_1724);
nor U2617 (N_2617,N_1857,N_1553);
nand U2618 (N_2618,N_1678,N_2030);
nand U2619 (N_2619,N_2217,N_1666);
nand U2620 (N_2620,N_1527,N_1814);
xor U2621 (N_2621,N_1700,N_1672);
nor U2622 (N_2622,N_2115,N_1507);
and U2623 (N_2623,N_2165,N_2045);
and U2624 (N_2624,N_1518,N_2035);
nor U2625 (N_2625,N_1524,N_1963);
nand U2626 (N_2626,N_2238,N_1614);
nand U2627 (N_2627,N_2054,N_2052);
nand U2628 (N_2628,N_2097,N_2079);
nor U2629 (N_2629,N_1901,N_1891);
nor U2630 (N_2630,N_1747,N_1877);
xnor U2631 (N_2631,N_2195,N_2095);
nor U2632 (N_2632,N_1895,N_2088);
nand U2633 (N_2633,N_1649,N_1739);
or U2634 (N_2634,N_1504,N_1996);
xnor U2635 (N_2635,N_1806,N_1767);
nand U2636 (N_2636,N_1903,N_2130);
and U2637 (N_2637,N_2226,N_2036);
nor U2638 (N_2638,N_1737,N_1563);
and U2639 (N_2639,N_2177,N_1609);
nand U2640 (N_2640,N_2229,N_1793);
or U2641 (N_2641,N_2157,N_1760);
xor U2642 (N_2642,N_1644,N_1646);
or U2643 (N_2643,N_2128,N_1765);
nor U2644 (N_2644,N_1781,N_1725);
nor U2645 (N_2645,N_1717,N_1971);
or U2646 (N_2646,N_1880,N_1916);
or U2647 (N_2647,N_1578,N_1513);
nand U2648 (N_2648,N_1974,N_2212);
nor U2649 (N_2649,N_1573,N_1604);
nand U2650 (N_2650,N_1909,N_2083);
xor U2651 (N_2651,N_2202,N_2179);
and U2652 (N_2652,N_1877,N_1633);
or U2653 (N_2653,N_2099,N_1591);
and U2654 (N_2654,N_1532,N_2045);
nor U2655 (N_2655,N_2059,N_1508);
and U2656 (N_2656,N_1578,N_1958);
or U2657 (N_2657,N_1886,N_1769);
nor U2658 (N_2658,N_1938,N_1935);
or U2659 (N_2659,N_1657,N_2212);
nor U2660 (N_2660,N_1772,N_1630);
and U2661 (N_2661,N_1624,N_1866);
and U2662 (N_2662,N_1562,N_1633);
nor U2663 (N_2663,N_2185,N_1666);
and U2664 (N_2664,N_2155,N_1723);
nor U2665 (N_2665,N_1632,N_1908);
xor U2666 (N_2666,N_1736,N_2246);
or U2667 (N_2667,N_2053,N_2092);
nor U2668 (N_2668,N_1723,N_2039);
or U2669 (N_2669,N_2126,N_1656);
or U2670 (N_2670,N_2048,N_2003);
xor U2671 (N_2671,N_2177,N_1863);
xnor U2672 (N_2672,N_1681,N_2071);
nor U2673 (N_2673,N_1860,N_2213);
and U2674 (N_2674,N_2190,N_1610);
and U2675 (N_2675,N_1891,N_1944);
and U2676 (N_2676,N_2245,N_2198);
and U2677 (N_2677,N_1539,N_2230);
nor U2678 (N_2678,N_1540,N_1842);
xor U2679 (N_2679,N_2189,N_1759);
nand U2680 (N_2680,N_1694,N_1617);
nand U2681 (N_2681,N_1731,N_2160);
nor U2682 (N_2682,N_2175,N_1523);
xor U2683 (N_2683,N_2189,N_1645);
and U2684 (N_2684,N_2150,N_2144);
xnor U2685 (N_2685,N_1860,N_1626);
or U2686 (N_2686,N_2231,N_2136);
nor U2687 (N_2687,N_2173,N_1689);
and U2688 (N_2688,N_2076,N_2152);
or U2689 (N_2689,N_1944,N_2184);
nand U2690 (N_2690,N_1517,N_1535);
nand U2691 (N_2691,N_2127,N_2210);
or U2692 (N_2692,N_2148,N_1961);
or U2693 (N_2693,N_1724,N_1840);
nand U2694 (N_2694,N_2012,N_1835);
xor U2695 (N_2695,N_1663,N_1970);
nand U2696 (N_2696,N_1634,N_1506);
nand U2697 (N_2697,N_1949,N_2183);
or U2698 (N_2698,N_1981,N_1651);
or U2699 (N_2699,N_1805,N_1560);
and U2700 (N_2700,N_2019,N_2066);
nor U2701 (N_2701,N_2190,N_1666);
and U2702 (N_2702,N_1918,N_1856);
nor U2703 (N_2703,N_1583,N_1951);
or U2704 (N_2704,N_1620,N_1957);
nand U2705 (N_2705,N_2083,N_2068);
or U2706 (N_2706,N_1756,N_2206);
and U2707 (N_2707,N_1623,N_2123);
nand U2708 (N_2708,N_2094,N_1537);
nor U2709 (N_2709,N_1654,N_1544);
nand U2710 (N_2710,N_2062,N_1645);
nor U2711 (N_2711,N_2016,N_1734);
or U2712 (N_2712,N_1847,N_1709);
nor U2713 (N_2713,N_1996,N_1818);
nand U2714 (N_2714,N_1713,N_1893);
or U2715 (N_2715,N_1916,N_1509);
xnor U2716 (N_2716,N_1588,N_1942);
and U2717 (N_2717,N_1807,N_1752);
and U2718 (N_2718,N_2085,N_1921);
nand U2719 (N_2719,N_1870,N_2052);
nor U2720 (N_2720,N_1842,N_1704);
xor U2721 (N_2721,N_2210,N_1834);
or U2722 (N_2722,N_1696,N_1799);
and U2723 (N_2723,N_1947,N_1859);
nand U2724 (N_2724,N_1613,N_1857);
nand U2725 (N_2725,N_1701,N_1579);
xor U2726 (N_2726,N_1785,N_1877);
nand U2727 (N_2727,N_1923,N_1592);
and U2728 (N_2728,N_1928,N_1661);
nand U2729 (N_2729,N_1573,N_2057);
and U2730 (N_2730,N_1531,N_2137);
or U2731 (N_2731,N_1612,N_1685);
nand U2732 (N_2732,N_1904,N_1763);
xnor U2733 (N_2733,N_1833,N_2104);
and U2734 (N_2734,N_1575,N_2154);
nor U2735 (N_2735,N_1652,N_2023);
or U2736 (N_2736,N_2148,N_1798);
nor U2737 (N_2737,N_2071,N_2143);
nor U2738 (N_2738,N_1982,N_1906);
nor U2739 (N_2739,N_1656,N_2222);
xor U2740 (N_2740,N_1993,N_2125);
and U2741 (N_2741,N_2136,N_1636);
and U2742 (N_2742,N_2069,N_1824);
and U2743 (N_2743,N_1544,N_1846);
nor U2744 (N_2744,N_1931,N_2233);
nor U2745 (N_2745,N_2180,N_2082);
or U2746 (N_2746,N_1738,N_1592);
and U2747 (N_2747,N_2227,N_1884);
nand U2748 (N_2748,N_1614,N_1658);
xor U2749 (N_2749,N_2009,N_1527);
nor U2750 (N_2750,N_1903,N_1533);
nor U2751 (N_2751,N_1948,N_2104);
nand U2752 (N_2752,N_2203,N_1959);
nand U2753 (N_2753,N_1829,N_2008);
nor U2754 (N_2754,N_2231,N_2076);
nor U2755 (N_2755,N_1949,N_2223);
nand U2756 (N_2756,N_2244,N_1866);
or U2757 (N_2757,N_2047,N_1581);
and U2758 (N_2758,N_1809,N_2048);
nor U2759 (N_2759,N_1960,N_2111);
nor U2760 (N_2760,N_1714,N_2166);
and U2761 (N_2761,N_1847,N_2137);
nand U2762 (N_2762,N_1601,N_1594);
and U2763 (N_2763,N_2098,N_1567);
or U2764 (N_2764,N_2016,N_1868);
and U2765 (N_2765,N_2024,N_1696);
or U2766 (N_2766,N_1857,N_1513);
xor U2767 (N_2767,N_2195,N_2242);
or U2768 (N_2768,N_2029,N_1653);
nand U2769 (N_2769,N_1809,N_2210);
nand U2770 (N_2770,N_1751,N_1659);
or U2771 (N_2771,N_1531,N_2145);
and U2772 (N_2772,N_2156,N_2199);
or U2773 (N_2773,N_1914,N_2215);
nor U2774 (N_2774,N_1565,N_1868);
and U2775 (N_2775,N_2062,N_1937);
and U2776 (N_2776,N_1609,N_2195);
or U2777 (N_2777,N_1711,N_1685);
or U2778 (N_2778,N_1550,N_2122);
nor U2779 (N_2779,N_1569,N_1555);
and U2780 (N_2780,N_1907,N_1937);
or U2781 (N_2781,N_1965,N_2182);
nor U2782 (N_2782,N_1596,N_2048);
nor U2783 (N_2783,N_1893,N_1906);
nor U2784 (N_2784,N_1655,N_1741);
nand U2785 (N_2785,N_2206,N_2095);
nor U2786 (N_2786,N_2058,N_1589);
nand U2787 (N_2787,N_1977,N_1896);
nor U2788 (N_2788,N_2138,N_1615);
nor U2789 (N_2789,N_2011,N_1788);
nand U2790 (N_2790,N_1820,N_1718);
nand U2791 (N_2791,N_1775,N_1557);
and U2792 (N_2792,N_1754,N_1529);
xnor U2793 (N_2793,N_1767,N_1916);
nand U2794 (N_2794,N_1721,N_1650);
xnor U2795 (N_2795,N_2127,N_2173);
and U2796 (N_2796,N_2099,N_1784);
nand U2797 (N_2797,N_1767,N_1773);
and U2798 (N_2798,N_2095,N_2166);
nor U2799 (N_2799,N_1935,N_1553);
or U2800 (N_2800,N_2121,N_1640);
and U2801 (N_2801,N_2119,N_1824);
or U2802 (N_2802,N_2037,N_1511);
nor U2803 (N_2803,N_1617,N_2179);
nor U2804 (N_2804,N_1587,N_2030);
or U2805 (N_2805,N_1878,N_2148);
nand U2806 (N_2806,N_1954,N_1691);
nand U2807 (N_2807,N_1978,N_1772);
and U2808 (N_2808,N_1573,N_1820);
or U2809 (N_2809,N_1589,N_2094);
and U2810 (N_2810,N_2221,N_1593);
and U2811 (N_2811,N_1667,N_1550);
nor U2812 (N_2812,N_1612,N_1806);
and U2813 (N_2813,N_1781,N_2103);
nor U2814 (N_2814,N_1826,N_1563);
nor U2815 (N_2815,N_1540,N_1746);
or U2816 (N_2816,N_2136,N_1707);
nand U2817 (N_2817,N_1892,N_1978);
or U2818 (N_2818,N_2217,N_1713);
and U2819 (N_2819,N_1640,N_1876);
nand U2820 (N_2820,N_2118,N_1648);
and U2821 (N_2821,N_2137,N_2100);
or U2822 (N_2822,N_2197,N_1620);
nand U2823 (N_2823,N_1634,N_2059);
nand U2824 (N_2824,N_2185,N_1500);
nor U2825 (N_2825,N_1506,N_2039);
xor U2826 (N_2826,N_1903,N_1785);
nor U2827 (N_2827,N_1696,N_1987);
nand U2828 (N_2828,N_1997,N_2120);
or U2829 (N_2829,N_2086,N_2039);
nor U2830 (N_2830,N_1625,N_1951);
xnor U2831 (N_2831,N_1748,N_2240);
or U2832 (N_2832,N_1771,N_1894);
or U2833 (N_2833,N_2163,N_1813);
nand U2834 (N_2834,N_2006,N_1735);
nor U2835 (N_2835,N_1592,N_1931);
nor U2836 (N_2836,N_1768,N_2117);
and U2837 (N_2837,N_1960,N_1535);
xnor U2838 (N_2838,N_2038,N_2028);
xor U2839 (N_2839,N_2082,N_1603);
nand U2840 (N_2840,N_1607,N_2098);
and U2841 (N_2841,N_2211,N_1971);
or U2842 (N_2842,N_2244,N_1663);
nor U2843 (N_2843,N_1729,N_1892);
or U2844 (N_2844,N_1813,N_1546);
nor U2845 (N_2845,N_1541,N_1625);
nor U2846 (N_2846,N_1758,N_1860);
nand U2847 (N_2847,N_2199,N_2176);
or U2848 (N_2848,N_1641,N_2213);
and U2849 (N_2849,N_1587,N_1692);
nor U2850 (N_2850,N_1573,N_1920);
and U2851 (N_2851,N_1845,N_1516);
and U2852 (N_2852,N_1570,N_2137);
xor U2853 (N_2853,N_2173,N_2009);
nor U2854 (N_2854,N_1523,N_1825);
or U2855 (N_2855,N_1612,N_2107);
or U2856 (N_2856,N_1991,N_1869);
and U2857 (N_2857,N_2244,N_1660);
or U2858 (N_2858,N_1896,N_1851);
or U2859 (N_2859,N_1634,N_2162);
nand U2860 (N_2860,N_1860,N_2050);
and U2861 (N_2861,N_2222,N_1502);
and U2862 (N_2862,N_1554,N_2126);
xor U2863 (N_2863,N_1829,N_1827);
or U2864 (N_2864,N_1949,N_2061);
and U2865 (N_2865,N_2061,N_1977);
or U2866 (N_2866,N_2057,N_1967);
and U2867 (N_2867,N_1970,N_2005);
xnor U2868 (N_2868,N_1796,N_1800);
nand U2869 (N_2869,N_1695,N_2057);
nor U2870 (N_2870,N_1871,N_2221);
and U2871 (N_2871,N_1584,N_2121);
nor U2872 (N_2872,N_1863,N_1963);
xor U2873 (N_2873,N_1806,N_1617);
nand U2874 (N_2874,N_2171,N_2233);
nand U2875 (N_2875,N_1919,N_1850);
and U2876 (N_2876,N_1858,N_1604);
and U2877 (N_2877,N_1645,N_2190);
or U2878 (N_2878,N_1570,N_1549);
or U2879 (N_2879,N_1969,N_1654);
and U2880 (N_2880,N_1621,N_1563);
xor U2881 (N_2881,N_1921,N_2110);
nor U2882 (N_2882,N_2234,N_1797);
or U2883 (N_2883,N_2104,N_1597);
nor U2884 (N_2884,N_2049,N_1628);
nand U2885 (N_2885,N_2152,N_2103);
nand U2886 (N_2886,N_1939,N_1861);
nand U2887 (N_2887,N_1753,N_1571);
nand U2888 (N_2888,N_2195,N_2191);
nand U2889 (N_2889,N_1818,N_1763);
nor U2890 (N_2890,N_1624,N_1917);
and U2891 (N_2891,N_1661,N_1889);
or U2892 (N_2892,N_1923,N_1577);
or U2893 (N_2893,N_1897,N_1660);
nor U2894 (N_2894,N_1977,N_1811);
nand U2895 (N_2895,N_1567,N_2143);
nand U2896 (N_2896,N_1806,N_1771);
xnor U2897 (N_2897,N_1808,N_1539);
nor U2898 (N_2898,N_1807,N_2053);
and U2899 (N_2899,N_1936,N_1867);
and U2900 (N_2900,N_2157,N_1739);
and U2901 (N_2901,N_1788,N_1515);
and U2902 (N_2902,N_2025,N_1620);
and U2903 (N_2903,N_1992,N_1821);
or U2904 (N_2904,N_2084,N_1839);
nand U2905 (N_2905,N_1666,N_1928);
nand U2906 (N_2906,N_1650,N_1837);
and U2907 (N_2907,N_2094,N_1629);
or U2908 (N_2908,N_1777,N_1566);
nand U2909 (N_2909,N_2074,N_1750);
xnor U2910 (N_2910,N_2215,N_1536);
and U2911 (N_2911,N_1520,N_2178);
or U2912 (N_2912,N_2215,N_2054);
xnor U2913 (N_2913,N_2168,N_1670);
and U2914 (N_2914,N_1862,N_1686);
nand U2915 (N_2915,N_1768,N_1899);
nand U2916 (N_2916,N_1862,N_1677);
or U2917 (N_2917,N_1842,N_1863);
nor U2918 (N_2918,N_1889,N_1913);
or U2919 (N_2919,N_2151,N_1871);
nor U2920 (N_2920,N_1987,N_1899);
and U2921 (N_2921,N_1924,N_2062);
nand U2922 (N_2922,N_2181,N_1879);
nor U2923 (N_2923,N_1606,N_1607);
xor U2924 (N_2924,N_1796,N_1906);
nor U2925 (N_2925,N_1958,N_1662);
nor U2926 (N_2926,N_2093,N_2014);
nor U2927 (N_2927,N_1944,N_2147);
nor U2928 (N_2928,N_2132,N_1975);
or U2929 (N_2929,N_2180,N_1687);
nor U2930 (N_2930,N_1896,N_2019);
or U2931 (N_2931,N_2121,N_2060);
and U2932 (N_2932,N_1970,N_1506);
and U2933 (N_2933,N_1593,N_1599);
nand U2934 (N_2934,N_1681,N_2103);
nor U2935 (N_2935,N_1689,N_1624);
xor U2936 (N_2936,N_2018,N_1888);
nand U2937 (N_2937,N_1632,N_1896);
and U2938 (N_2938,N_1620,N_1692);
or U2939 (N_2939,N_1529,N_1549);
or U2940 (N_2940,N_1926,N_2178);
xnor U2941 (N_2941,N_1741,N_1679);
nor U2942 (N_2942,N_1630,N_2063);
nor U2943 (N_2943,N_1934,N_1997);
xnor U2944 (N_2944,N_1814,N_1575);
nor U2945 (N_2945,N_1909,N_1810);
and U2946 (N_2946,N_2105,N_2043);
and U2947 (N_2947,N_1742,N_1807);
or U2948 (N_2948,N_2110,N_1576);
nor U2949 (N_2949,N_2070,N_2221);
nand U2950 (N_2950,N_1645,N_1756);
nor U2951 (N_2951,N_1530,N_2078);
nor U2952 (N_2952,N_1748,N_1526);
xnor U2953 (N_2953,N_1516,N_1770);
nand U2954 (N_2954,N_1736,N_2147);
nand U2955 (N_2955,N_2245,N_2163);
nand U2956 (N_2956,N_1617,N_2039);
xor U2957 (N_2957,N_2168,N_1728);
xnor U2958 (N_2958,N_1652,N_1614);
and U2959 (N_2959,N_1911,N_2111);
and U2960 (N_2960,N_1548,N_1866);
nor U2961 (N_2961,N_2091,N_2075);
nor U2962 (N_2962,N_1721,N_2214);
nand U2963 (N_2963,N_1836,N_2248);
xnor U2964 (N_2964,N_1997,N_1795);
and U2965 (N_2965,N_1643,N_1883);
or U2966 (N_2966,N_1752,N_1683);
nand U2967 (N_2967,N_1723,N_1771);
nand U2968 (N_2968,N_1579,N_1577);
nand U2969 (N_2969,N_2237,N_2018);
xor U2970 (N_2970,N_1502,N_1696);
xnor U2971 (N_2971,N_1624,N_2206);
nor U2972 (N_2972,N_1588,N_1961);
nor U2973 (N_2973,N_1786,N_1679);
nor U2974 (N_2974,N_1817,N_1595);
or U2975 (N_2975,N_1695,N_1684);
xor U2976 (N_2976,N_1816,N_1769);
nand U2977 (N_2977,N_2105,N_1968);
xnor U2978 (N_2978,N_1813,N_1615);
nand U2979 (N_2979,N_2221,N_2018);
xor U2980 (N_2980,N_1745,N_1893);
or U2981 (N_2981,N_1878,N_2180);
xnor U2982 (N_2982,N_1560,N_1700);
or U2983 (N_2983,N_1742,N_2185);
or U2984 (N_2984,N_1520,N_2035);
and U2985 (N_2985,N_1612,N_2113);
nor U2986 (N_2986,N_1853,N_1924);
xor U2987 (N_2987,N_2181,N_1990);
or U2988 (N_2988,N_2186,N_1617);
or U2989 (N_2989,N_1632,N_1627);
and U2990 (N_2990,N_1545,N_1727);
nor U2991 (N_2991,N_1937,N_1622);
or U2992 (N_2992,N_1670,N_2165);
xor U2993 (N_2993,N_1650,N_1514);
xor U2994 (N_2994,N_1941,N_2109);
or U2995 (N_2995,N_1728,N_1875);
nand U2996 (N_2996,N_2096,N_1606);
xnor U2997 (N_2997,N_1510,N_1676);
xnor U2998 (N_2998,N_1746,N_1744);
and U2999 (N_2999,N_1755,N_1694);
nor U3000 (N_3000,N_2413,N_2758);
or U3001 (N_3001,N_2660,N_2869);
nor U3002 (N_3002,N_2584,N_2813);
nand U3003 (N_3003,N_2770,N_2775);
nand U3004 (N_3004,N_2401,N_2490);
xor U3005 (N_3005,N_2583,N_2495);
or U3006 (N_3006,N_2559,N_2663);
or U3007 (N_3007,N_2965,N_2313);
and U3008 (N_3008,N_2947,N_2318);
nor U3009 (N_3009,N_2473,N_2738);
or U3010 (N_3010,N_2784,N_2375);
and U3011 (N_3011,N_2740,N_2968);
nor U3012 (N_3012,N_2700,N_2661);
nand U3013 (N_3013,N_2930,N_2695);
and U3014 (N_3014,N_2647,N_2529);
nor U3015 (N_3015,N_2315,N_2847);
nor U3016 (N_3016,N_2260,N_2448);
nor U3017 (N_3017,N_2861,N_2333);
nor U3018 (N_3018,N_2891,N_2256);
nor U3019 (N_3019,N_2677,N_2554);
and U3020 (N_3020,N_2602,N_2270);
nand U3021 (N_3021,N_2701,N_2696);
nand U3022 (N_3022,N_2773,N_2644);
nand U3023 (N_3023,N_2766,N_2938);
and U3024 (N_3024,N_2340,N_2295);
and U3025 (N_3025,N_2625,N_2634);
or U3026 (N_3026,N_2522,N_2285);
or U3027 (N_3027,N_2936,N_2655);
nand U3028 (N_3028,N_2859,N_2386);
or U3029 (N_3029,N_2452,N_2320);
xor U3030 (N_3030,N_2842,N_2935);
and U3031 (N_3031,N_2761,N_2835);
nor U3032 (N_3032,N_2369,N_2988);
and U3033 (N_3033,N_2540,N_2789);
or U3034 (N_3034,N_2864,N_2404);
and U3035 (N_3035,N_2759,N_2253);
nand U3036 (N_3036,N_2564,N_2389);
nor U3037 (N_3037,N_2361,N_2860);
nand U3038 (N_3038,N_2347,N_2402);
nand U3039 (N_3039,N_2580,N_2458);
and U3040 (N_3040,N_2420,N_2801);
and U3041 (N_3041,N_2905,N_2697);
nand U3042 (N_3042,N_2341,N_2378);
and U3043 (N_3043,N_2960,N_2379);
xor U3044 (N_3044,N_2376,N_2870);
and U3045 (N_3045,N_2373,N_2337);
nor U3046 (N_3046,N_2676,N_2531);
nor U3047 (N_3047,N_2631,N_2913);
or U3048 (N_3048,N_2539,N_2585);
xnor U3049 (N_3049,N_2727,N_2591);
xor U3050 (N_3050,N_2872,N_2547);
and U3051 (N_3051,N_2818,N_2915);
or U3052 (N_3052,N_2920,N_2501);
nand U3053 (N_3053,N_2298,N_2506);
nand U3054 (N_3054,N_2508,N_2480);
and U3055 (N_3055,N_2488,N_2868);
or U3056 (N_3056,N_2551,N_2550);
and U3057 (N_3057,N_2989,N_2571);
and U3058 (N_3058,N_2787,N_2314);
and U3059 (N_3059,N_2967,N_2768);
or U3060 (N_3060,N_2713,N_2962);
nand U3061 (N_3061,N_2980,N_2577);
and U3062 (N_3062,N_2502,N_2291);
nand U3063 (N_3063,N_2678,N_2690);
and U3064 (N_3064,N_2549,N_2335);
or U3065 (N_3065,N_2463,N_2416);
or U3066 (N_3066,N_2892,N_2259);
nand U3067 (N_3067,N_2900,N_2805);
or U3068 (N_3068,N_2767,N_2772);
nand U3069 (N_3069,N_2654,N_2664);
nand U3070 (N_3070,N_2865,N_2675);
and U3071 (N_3071,N_2693,N_2412);
and U3072 (N_3072,N_2945,N_2477);
nor U3073 (N_3073,N_2894,N_2575);
nand U3074 (N_3074,N_2565,N_2781);
nor U3075 (N_3075,N_2994,N_2466);
and U3076 (N_3076,N_2293,N_2266);
nor U3077 (N_3077,N_2574,N_2380);
and U3078 (N_3078,N_2395,N_2685);
nor U3079 (N_3079,N_2494,N_2358);
or U3080 (N_3080,N_2757,N_2810);
nor U3081 (N_3081,N_2826,N_2966);
xnor U3082 (N_3082,N_2512,N_2568);
and U3083 (N_3083,N_2462,N_2306);
and U3084 (N_3084,N_2741,N_2521);
or U3085 (N_3085,N_2925,N_2852);
nor U3086 (N_3086,N_2409,N_2288);
or U3087 (N_3087,N_2804,N_2706);
and U3088 (N_3088,N_2519,N_2455);
and U3089 (N_3089,N_2659,N_2997);
or U3090 (N_3090,N_2652,N_2476);
and U3091 (N_3091,N_2811,N_2536);
nand U3092 (N_3092,N_2623,N_2453);
nor U3093 (N_3093,N_2504,N_2895);
nand U3094 (N_3094,N_2702,N_2717);
and U3095 (N_3095,N_2614,N_2914);
xnor U3096 (N_3096,N_2489,N_2934);
nand U3097 (N_3097,N_2563,N_2820);
or U3098 (N_3098,N_2721,N_2704);
or U3099 (N_3099,N_2326,N_2941);
nor U3100 (N_3100,N_2526,N_2986);
xor U3101 (N_3101,N_2507,N_2523);
nand U3102 (N_3102,N_2626,N_2586);
nor U3103 (N_3103,N_2977,N_2332);
or U3104 (N_3104,N_2751,N_2567);
and U3105 (N_3105,N_2394,N_2884);
and U3106 (N_3106,N_2898,N_2427);
xor U3107 (N_3107,N_2274,N_2569);
nor U3108 (N_3108,N_2893,N_2537);
or U3109 (N_3109,N_2595,N_2518);
nor U3110 (N_3110,N_2349,N_2527);
nand U3111 (N_3111,N_2771,N_2525);
or U3112 (N_3112,N_2733,N_2434);
nand U3113 (N_3113,N_2823,N_2750);
or U3114 (N_3114,N_2788,N_2710);
and U3115 (N_3115,N_2352,N_2929);
nor U3116 (N_3116,N_2981,N_2628);
or U3117 (N_3117,N_2292,N_2827);
nand U3118 (N_3118,N_2845,N_2742);
nand U3119 (N_3119,N_2610,N_2912);
nand U3120 (N_3120,N_2774,N_2449);
and U3121 (N_3121,N_2728,N_2809);
nand U3122 (N_3122,N_2570,N_2290);
or U3123 (N_3123,N_2438,N_2381);
nand U3124 (N_3124,N_2323,N_2346);
nand U3125 (N_3125,N_2712,N_2856);
nand U3126 (N_3126,N_2698,N_2599);
nand U3127 (N_3127,N_2843,N_2533);
and U3128 (N_3128,N_2776,N_2368);
xor U3129 (N_3129,N_2933,N_2437);
and U3130 (N_3130,N_2408,N_2642);
and U3131 (N_3131,N_2435,N_2328);
and U3132 (N_3132,N_2544,N_2909);
and U3133 (N_3133,N_2545,N_2271);
nor U3134 (N_3134,N_2275,N_2593);
xor U3135 (N_3135,N_2737,N_2907);
nand U3136 (N_3136,N_2483,N_2803);
or U3137 (N_3137,N_2307,N_2429);
and U3138 (N_3138,N_2921,N_2639);
and U3139 (N_3139,N_2558,N_2719);
and U3140 (N_3140,N_2978,N_2500);
or U3141 (N_3141,N_2927,N_2633);
and U3142 (N_3142,N_2680,N_2431);
nor U3143 (N_3143,N_2786,N_2976);
nor U3144 (N_3144,N_2468,N_2880);
xor U3145 (N_3145,N_2798,N_2783);
nor U3146 (N_3146,N_2854,N_2688);
nand U3147 (N_3147,N_2613,N_2645);
nor U3148 (N_3148,N_2792,N_2396);
nor U3149 (N_3149,N_2419,N_2871);
xor U3150 (N_3150,N_2600,N_2257);
or U3151 (N_3151,N_2808,N_2836);
and U3152 (N_3152,N_2604,N_2724);
nand U3153 (N_3153,N_2999,N_2755);
nand U3154 (N_3154,N_2284,N_2879);
or U3155 (N_3155,N_2418,N_2590);
nor U3156 (N_3156,N_2345,N_2902);
or U3157 (N_3157,N_2481,N_2354);
and U3158 (N_3158,N_2447,N_2594);
nor U3159 (N_3159,N_2319,N_2904);
nand U3160 (N_3160,N_2387,N_2867);
nand U3161 (N_3161,N_2683,N_2679);
nor U3162 (N_3162,N_2262,N_2487);
or U3163 (N_3163,N_2436,N_2943);
or U3164 (N_3164,N_2428,N_2838);
and U3165 (N_3165,N_2374,N_2325);
and U3166 (N_3166,N_2991,N_2731);
and U3167 (N_3167,N_2362,N_2658);
or U3168 (N_3168,N_2874,N_2649);
or U3169 (N_3169,N_2573,N_2530);
nand U3170 (N_3170,N_2255,N_2665);
nand U3171 (N_3171,N_2953,N_2806);
or U3172 (N_3172,N_2674,N_2524);
xnor U3173 (N_3173,N_2417,N_2839);
and U3174 (N_3174,N_2819,N_2311);
and U3175 (N_3175,N_2283,N_2336);
nor U3176 (N_3176,N_2310,N_2250);
and U3177 (N_3177,N_2881,N_2763);
and U3178 (N_3178,N_2754,N_2372);
or U3179 (N_3179,N_2735,N_2825);
and U3180 (N_3180,N_2397,N_2391);
and U3181 (N_3181,N_2736,N_2334);
and U3182 (N_3182,N_2265,N_2648);
and U3183 (N_3183,N_2300,N_2460);
or U3184 (N_3184,N_2961,N_2356);
nand U3185 (N_3185,N_2272,N_2327);
nand U3186 (N_3186,N_2425,N_2432);
and U3187 (N_3187,N_2998,N_2329);
or U3188 (N_3188,N_2446,N_2456);
or U3189 (N_3189,N_2777,N_2622);
and U3190 (N_3190,N_2305,N_2399);
nor U3191 (N_3191,N_2392,N_2261);
or U3192 (N_3192,N_2692,N_2297);
nor U3193 (N_3193,N_2765,N_2673);
nor U3194 (N_3194,N_2791,N_2670);
nand U3195 (N_3195,N_2922,N_2830);
nor U3196 (N_3196,N_2753,N_2520);
nor U3197 (N_3197,N_2667,N_2946);
and U3198 (N_3198,N_2450,N_2708);
or U3199 (N_3199,N_2707,N_2889);
and U3200 (N_3200,N_2739,N_2878);
nor U3201 (N_3201,N_2899,N_2726);
nor U3202 (N_3202,N_2903,N_2722);
nor U3203 (N_3203,N_2883,N_2479);
or U3204 (N_3204,N_2385,N_2546);
nor U3205 (N_3205,N_2343,N_2672);
nand U3206 (N_3206,N_2982,N_2411);
nand U3207 (N_3207,N_2364,N_2850);
nand U3208 (N_3208,N_2862,N_2355);
nor U3209 (N_3209,N_2687,N_2752);
and U3210 (N_3210,N_2897,N_2485);
or U3211 (N_3211,N_2282,N_2331);
nor U3212 (N_3212,N_2746,N_2919);
or U3213 (N_3213,N_2555,N_2597);
and U3214 (N_3214,N_2908,N_2312);
nor U3215 (N_3215,N_2668,N_2430);
nand U3216 (N_3216,N_2681,N_2360);
or U3217 (N_3217,N_2576,N_2730);
nor U3218 (N_3218,N_2640,N_2882);
or U3219 (N_3219,N_2484,N_2492);
nand U3220 (N_3220,N_2511,N_2371);
or U3221 (N_3221,N_2280,N_2344);
and U3222 (N_3222,N_2444,N_2918);
and U3223 (N_3223,N_2756,N_2888);
nand U3224 (N_3224,N_2800,N_2302);
or U3225 (N_3225,N_2607,N_2421);
nand U3226 (N_3226,N_2954,N_2932);
nor U3227 (N_3227,N_2415,N_2618);
or U3228 (N_3228,N_2393,N_2617);
and U3229 (N_3229,N_2612,N_2951);
or U3230 (N_3230,N_2834,N_2684);
and U3231 (N_3231,N_2699,N_2384);
nor U3232 (N_3232,N_2797,N_2829);
xor U3233 (N_3233,N_2474,N_2917);
nor U3234 (N_3234,N_2445,N_2470);
nor U3235 (N_3235,N_2273,N_2632);
and U3236 (N_3236,N_2475,N_2461);
nand U3237 (N_3237,N_2985,N_2407);
and U3238 (N_3238,N_2970,N_2923);
or U3239 (N_3239,N_2471,N_2308);
nor U3240 (N_3240,N_2482,N_2541);
nand U3241 (N_3241,N_2983,N_2296);
or U3242 (N_3242,N_2560,N_2718);
nand U3243 (N_3243,N_2831,N_2636);
or U3244 (N_3244,N_2464,N_2542);
and U3245 (N_3245,N_2388,N_2469);
xor U3246 (N_3246,N_2581,N_2566);
nand U3247 (N_3247,N_2348,N_2299);
or U3248 (N_3248,N_2548,N_2359);
and U3249 (N_3249,N_2269,N_2732);
nand U3250 (N_3250,N_2646,N_2322);
nand U3251 (N_3251,N_2656,N_2383);
nor U3252 (N_3252,N_2258,N_2303);
nor U3253 (N_3253,N_2799,N_2924);
or U3254 (N_3254,N_2254,N_2782);
xor U3255 (N_3255,N_2744,N_2630);
or U3256 (N_3256,N_2916,N_2451);
or U3257 (N_3257,N_2992,N_2802);
xor U3258 (N_3258,N_2264,N_2886);
and U3259 (N_3259,N_2906,N_2844);
and U3260 (N_3260,N_2794,N_2592);
or U3261 (N_3261,N_2263,N_2338);
nand U3262 (N_3262,N_2390,N_2588);
and U3263 (N_3263,N_2509,N_2779);
and U3264 (N_3264,N_2911,N_2817);
and U3265 (N_3265,N_2846,N_2734);
and U3266 (N_3266,N_2764,N_2339);
nand U3267 (N_3267,N_2534,N_2552);
nand U3268 (N_3268,N_2638,N_2609);
nor U3269 (N_3269,N_2964,N_2366);
nand U3270 (N_3270,N_2400,N_2990);
nor U3271 (N_3271,N_2637,N_2828);
xor U3272 (N_3272,N_2330,N_2928);
and U3273 (N_3273,N_2824,N_2324);
nand U3274 (N_3274,N_2745,N_2793);
nand U3275 (N_3275,N_2532,N_2875);
nor U3276 (N_3276,N_2422,N_2984);
nor U3277 (N_3277,N_2457,N_2975);
xnor U3278 (N_3278,N_2365,N_2505);
xor U3279 (N_3279,N_2866,N_2406);
nand U3280 (N_3280,N_2851,N_2309);
or U3281 (N_3281,N_2948,N_2703);
nand U3282 (N_3282,N_2493,N_2952);
nor U3283 (N_3283,N_2287,N_2276);
or U3284 (N_3284,N_2651,N_2382);
nand U3285 (N_3285,N_2840,N_2926);
and U3286 (N_3286,N_2478,N_2440);
or U3287 (N_3287,N_2849,N_2725);
or U3288 (N_3288,N_2553,N_2949);
and U3289 (N_3289,N_2942,N_2812);
and U3290 (N_3290,N_2301,N_2723);
or U3291 (N_3291,N_2979,N_2627);
and U3292 (N_3292,N_2398,N_2514);
or U3293 (N_3293,N_2465,N_2510);
nand U3294 (N_3294,N_2277,N_2956);
or U3295 (N_3295,N_2317,N_2996);
nand U3296 (N_3296,N_2971,N_2589);
or U3297 (N_3297,N_2987,N_2972);
xor U3298 (N_3298,N_2749,N_2937);
nand U3299 (N_3299,N_2837,N_2497);
or U3300 (N_3300,N_2426,N_2855);
nand U3301 (N_3301,N_2896,N_2433);
or U3302 (N_3302,N_2498,N_2516);
nor U3303 (N_3303,N_2821,N_2528);
nand U3304 (N_3304,N_2621,N_2885);
and U3305 (N_3305,N_2579,N_2790);
and U3306 (N_3306,N_2857,N_2833);
nor U3307 (N_3307,N_2769,N_2944);
or U3308 (N_3308,N_2410,N_2795);
and U3309 (N_3309,N_2289,N_2760);
nand U3310 (N_3310,N_2321,N_2641);
nand U3311 (N_3311,N_2294,N_2281);
nand U3312 (N_3312,N_2691,N_2729);
xor U3313 (N_3313,N_2832,N_2743);
nor U3314 (N_3314,N_2513,N_2268);
or U3315 (N_3315,N_2686,N_2762);
or U3316 (N_3316,N_2496,N_2543);
and U3317 (N_3317,N_2278,N_2562);
and U3318 (N_3318,N_2403,N_2424);
nor U3319 (N_3319,N_2414,N_2304);
nand U3320 (N_3320,N_2596,N_2657);
nor U3321 (N_3321,N_2608,N_2814);
nand U3322 (N_3322,N_2443,N_2561);
nand U3323 (N_3323,N_2705,N_2969);
and U3324 (N_3324,N_2711,N_2643);
or U3325 (N_3325,N_2557,N_2682);
nand U3326 (N_3326,N_2252,N_2377);
and U3327 (N_3327,N_2910,N_2459);
and U3328 (N_3328,N_2503,N_2615);
and U3329 (N_3329,N_2650,N_2538);
or U3330 (N_3330,N_2901,N_2535);
or U3331 (N_3331,N_2620,N_2587);
and U3332 (N_3332,N_2286,N_2689);
and U3333 (N_3333,N_2370,N_2715);
or U3334 (N_3334,N_2876,N_2441);
nand U3335 (N_3335,N_2841,N_2556);
xnor U3336 (N_3336,N_2350,N_2662);
and U3337 (N_3337,N_2363,N_2694);
and U3338 (N_3338,N_2472,N_2666);
and U3339 (N_3339,N_2423,N_2367);
and U3340 (N_3340,N_2796,N_2351);
nor U3341 (N_3341,N_2963,N_2747);
and U3342 (N_3342,N_2822,N_2486);
nand U3343 (N_3343,N_2957,N_2454);
or U3344 (N_3344,N_2491,N_2606);
and U3345 (N_3345,N_2955,N_2353);
nor U3346 (N_3346,N_2578,N_2785);
and U3347 (N_3347,N_2974,N_2950);
xnor U3348 (N_3348,N_2635,N_2671);
nand U3349 (N_3349,N_2887,N_2939);
and U3350 (N_3350,N_2442,N_2439);
nand U3351 (N_3351,N_2959,N_2624);
or U3352 (N_3352,N_2720,N_2467);
nand U3353 (N_3353,N_2877,N_2931);
nor U3354 (N_3354,N_2582,N_2815);
or U3355 (N_3355,N_2993,N_2778);
xor U3356 (N_3356,N_2995,N_2714);
or U3357 (N_3357,N_2499,N_2853);
nor U3358 (N_3358,N_2848,N_2405);
nor U3359 (N_3359,N_2342,N_2748);
nand U3360 (N_3360,N_2598,N_2807);
and U3361 (N_3361,N_2611,N_2669);
nor U3362 (N_3362,N_2316,N_2940);
and U3363 (N_3363,N_2780,N_2619);
or U3364 (N_3364,N_2709,N_2716);
xnor U3365 (N_3365,N_2858,N_2605);
nor U3366 (N_3366,N_2616,N_2515);
and U3367 (N_3367,N_2601,N_2816);
nor U3368 (N_3368,N_2279,N_2958);
nand U3369 (N_3369,N_2890,N_2603);
and U3370 (N_3370,N_2873,N_2251);
nand U3371 (N_3371,N_2517,N_2653);
or U3372 (N_3372,N_2357,N_2629);
xor U3373 (N_3373,N_2973,N_2267);
and U3374 (N_3374,N_2863,N_2572);
or U3375 (N_3375,N_2802,N_2401);
and U3376 (N_3376,N_2527,N_2717);
or U3377 (N_3377,N_2555,N_2468);
and U3378 (N_3378,N_2447,N_2922);
xor U3379 (N_3379,N_2674,N_2287);
nor U3380 (N_3380,N_2869,N_2626);
and U3381 (N_3381,N_2866,N_2520);
and U3382 (N_3382,N_2386,N_2713);
and U3383 (N_3383,N_2292,N_2645);
nand U3384 (N_3384,N_2352,N_2428);
nand U3385 (N_3385,N_2416,N_2999);
nand U3386 (N_3386,N_2792,N_2855);
and U3387 (N_3387,N_2547,N_2410);
nor U3388 (N_3388,N_2490,N_2314);
or U3389 (N_3389,N_2730,N_2806);
nor U3390 (N_3390,N_2686,N_2257);
and U3391 (N_3391,N_2862,N_2938);
and U3392 (N_3392,N_2408,N_2915);
nor U3393 (N_3393,N_2341,N_2728);
xor U3394 (N_3394,N_2813,N_2715);
nand U3395 (N_3395,N_2350,N_2782);
nand U3396 (N_3396,N_2711,N_2563);
nand U3397 (N_3397,N_2575,N_2852);
or U3398 (N_3398,N_2956,N_2575);
nor U3399 (N_3399,N_2393,N_2621);
or U3400 (N_3400,N_2719,N_2924);
or U3401 (N_3401,N_2675,N_2807);
and U3402 (N_3402,N_2872,N_2341);
and U3403 (N_3403,N_2888,N_2949);
and U3404 (N_3404,N_2522,N_2512);
xor U3405 (N_3405,N_2333,N_2604);
or U3406 (N_3406,N_2320,N_2635);
nor U3407 (N_3407,N_2942,N_2596);
nor U3408 (N_3408,N_2689,N_2520);
nand U3409 (N_3409,N_2666,N_2599);
nand U3410 (N_3410,N_2755,N_2454);
nor U3411 (N_3411,N_2661,N_2816);
xnor U3412 (N_3412,N_2915,N_2395);
and U3413 (N_3413,N_2696,N_2561);
nor U3414 (N_3414,N_2646,N_2756);
and U3415 (N_3415,N_2274,N_2743);
or U3416 (N_3416,N_2279,N_2738);
nand U3417 (N_3417,N_2755,N_2607);
and U3418 (N_3418,N_2630,N_2977);
nand U3419 (N_3419,N_2377,N_2405);
nand U3420 (N_3420,N_2678,N_2778);
and U3421 (N_3421,N_2560,N_2434);
or U3422 (N_3422,N_2552,N_2798);
nor U3423 (N_3423,N_2269,N_2929);
and U3424 (N_3424,N_2403,N_2585);
xor U3425 (N_3425,N_2637,N_2337);
xnor U3426 (N_3426,N_2911,N_2297);
nand U3427 (N_3427,N_2374,N_2535);
xor U3428 (N_3428,N_2960,N_2814);
nor U3429 (N_3429,N_2922,N_2884);
nand U3430 (N_3430,N_2521,N_2933);
or U3431 (N_3431,N_2976,N_2863);
nor U3432 (N_3432,N_2299,N_2559);
xnor U3433 (N_3433,N_2305,N_2410);
nand U3434 (N_3434,N_2446,N_2873);
or U3435 (N_3435,N_2266,N_2868);
xnor U3436 (N_3436,N_2740,N_2287);
nand U3437 (N_3437,N_2331,N_2337);
and U3438 (N_3438,N_2941,N_2823);
nor U3439 (N_3439,N_2418,N_2654);
and U3440 (N_3440,N_2748,N_2855);
or U3441 (N_3441,N_2644,N_2712);
nand U3442 (N_3442,N_2800,N_2742);
xnor U3443 (N_3443,N_2935,N_2659);
nor U3444 (N_3444,N_2933,N_2585);
and U3445 (N_3445,N_2607,N_2790);
or U3446 (N_3446,N_2608,N_2972);
or U3447 (N_3447,N_2357,N_2660);
nand U3448 (N_3448,N_2475,N_2295);
xor U3449 (N_3449,N_2893,N_2660);
nand U3450 (N_3450,N_2738,N_2808);
nand U3451 (N_3451,N_2357,N_2639);
or U3452 (N_3452,N_2673,N_2703);
nor U3453 (N_3453,N_2647,N_2585);
xor U3454 (N_3454,N_2891,N_2715);
or U3455 (N_3455,N_2505,N_2815);
nor U3456 (N_3456,N_2808,N_2356);
nand U3457 (N_3457,N_2764,N_2594);
or U3458 (N_3458,N_2294,N_2881);
or U3459 (N_3459,N_2773,N_2661);
and U3460 (N_3460,N_2751,N_2324);
and U3461 (N_3461,N_2925,N_2924);
and U3462 (N_3462,N_2473,N_2501);
or U3463 (N_3463,N_2775,N_2454);
nor U3464 (N_3464,N_2730,N_2280);
nand U3465 (N_3465,N_2800,N_2372);
or U3466 (N_3466,N_2944,N_2440);
or U3467 (N_3467,N_2561,N_2545);
xor U3468 (N_3468,N_2721,N_2646);
nor U3469 (N_3469,N_2270,N_2916);
nand U3470 (N_3470,N_2454,N_2591);
and U3471 (N_3471,N_2470,N_2973);
or U3472 (N_3472,N_2425,N_2858);
nor U3473 (N_3473,N_2286,N_2419);
and U3474 (N_3474,N_2343,N_2321);
or U3475 (N_3475,N_2859,N_2860);
xor U3476 (N_3476,N_2802,N_2756);
nand U3477 (N_3477,N_2598,N_2620);
and U3478 (N_3478,N_2838,N_2423);
nor U3479 (N_3479,N_2563,N_2968);
nor U3480 (N_3480,N_2287,N_2742);
and U3481 (N_3481,N_2689,N_2714);
nor U3482 (N_3482,N_2544,N_2348);
or U3483 (N_3483,N_2658,N_2938);
nand U3484 (N_3484,N_2448,N_2532);
nor U3485 (N_3485,N_2734,N_2843);
or U3486 (N_3486,N_2296,N_2969);
nor U3487 (N_3487,N_2649,N_2943);
nor U3488 (N_3488,N_2942,N_2568);
xor U3489 (N_3489,N_2887,N_2902);
or U3490 (N_3490,N_2532,N_2464);
or U3491 (N_3491,N_2583,N_2852);
or U3492 (N_3492,N_2686,N_2379);
or U3493 (N_3493,N_2630,N_2860);
xor U3494 (N_3494,N_2811,N_2266);
or U3495 (N_3495,N_2287,N_2881);
or U3496 (N_3496,N_2422,N_2735);
nand U3497 (N_3497,N_2368,N_2991);
and U3498 (N_3498,N_2288,N_2271);
and U3499 (N_3499,N_2777,N_2281);
and U3500 (N_3500,N_2798,N_2373);
and U3501 (N_3501,N_2509,N_2526);
or U3502 (N_3502,N_2631,N_2354);
nor U3503 (N_3503,N_2266,N_2657);
or U3504 (N_3504,N_2306,N_2630);
nand U3505 (N_3505,N_2427,N_2482);
or U3506 (N_3506,N_2884,N_2807);
and U3507 (N_3507,N_2925,N_2263);
and U3508 (N_3508,N_2322,N_2356);
nor U3509 (N_3509,N_2796,N_2835);
nor U3510 (N_3510,N_2738,N_2377);
nor U3511 (N_3511,N_2458,N_2870);
or U3512 (N_3512,N_2953,N_2741);
nor U3513 (N_3513,N_2476,N_2636);
and U3514 (N_3514,N_2650,N_2419);
or U3515 (N_3515,N_2487,N_2804);
or U3516 (N_3516,N_2575,N_2538);
nor U3517 (N_3517,N_2978,N_2470);
nand U3518 (N_3518,N_2961,N_2483);
or U3519 (N_3519,N_2896,N_2365);
nand U3520 (N_3520,N_2540,N_2544);
nor U3521 (N_3521,N_2923,N_2483);
or U3522 (N_3522,N_2960,N_2609);
nor U3523 (N_3523,N_2717,N_2819);
nor U3524 (N_3524,N_2678,N_2869);
or U3525 (N_3525,N_2614,N_2790);
xnor U3526 (N_3526,N_2755,N_2265);
nor U3527 (N_3527,N_2259,N_2774);
nand U3528 (N_3528,N_2813,N_2662);
nand U3529 (N_3529,N_2848,N_2891);
and U3530 (N_3530,N_2822,N_2839);
nor U3531 (N_3531,N_2998,N_2844);
nand U3532 (N_3532,N_2671,N_2795);
or U3533 (N_3533,N_2698,N_2656);
or U3534 (N_3534,N_2591,N_2477);
and U3535 (N_3535,N_2493,N_2739);
or U3536 (N_3536,N_2483,N_2270);
xnor U3537 (N_3537,N_2685,N_2977);
xor U3538 (N_3538,N_2382,N_2729);
xor U3539 (N_3539,N_2313,N_2614);
nor U3540 (N_3540,N_2974,N_2307);
or U3541 (N_3541,N_2830,N_2626);
and U3542 (N_3542,N_2602,N_2442);
nor U3543 (N_3543,N_2383,N_2534);
and U3544 (N_3544,N_2727,N_2379);
nand U3545 (N_3545,N_2707,N_2969);
and U3546 (N_3546,N_2738,N_2280);
nand U3547 (N_3547,N_2511,N_2470);
and U3548 (N_3548,N_2917,N_2886);
and U3549 (N_3549,N_2861,N_2975);
nor U3550 (N_3550,N_2373,N_2473);
and U3551 (N_3551,N_2823,N_2901);
and U3552 (N_3552,N_2633,N_2299);
nor U3553 (N_3553,N_2621,N_2607);
or U3554 (N_3554,N_2772,N_2710);
or U3555 (N_3555,N_2851,N_2770);
nor U3556 (N_3556,N_2539,N_2564);
nor U3557 (N_3557,N_2732,N_2309);
nor U3558 (N_3558,N_2323,N_2528);
or U3559 (N_3559,N_2470,N_2261);
nand U3560 (N_3560,N_2866,N_2460);
nand U3561 (N_3561,N_2674,N_2884);
xnor U3562 (N_3562,N_2527,N_2391);
xnor U3563 (N_3563,N_2393,N_2883);
and U3564 (N_3564,N_2390,N_2846);
or U3565 (N_3565,N_2478,N_2753);
and U3566 (N_3566,N_2855,N_2992);
nor U3567 (N_3567,N_2752,N_2361);
or U3568 (N_3568,N_2782,N_2744);
nand U3569 (N_3569,N_2750,N_2920);
nand U3570 (N_3570,N_2415,N_2910);
nand U3571 (N_3571,N_2780,N_2638);
or U3572 (N_3572,N_2260,N_2859);
xnor U3573 (N_3573,N_2738,N_2576);
nor U3574 (N_3574,N_2987,N_2307);
or U3575 (N_3575,N_2259,N_2927);
and U3576 (N_3576,N_2488,N_2578);
and U3577 (N_3577,N_2297,N_2964);
xnor U3578 (N_3578,N_2754,N_2676);
xor U3579 (N_3579,N_2500,N_2603);
nand U3580 (N_3580,N_2611,N_2873);
or U3581 (N_3581,N_2400,N_2575);
nor U3582 (N_3582,N_2730,N_2273);
xnor U3583 (N_3583,N_2398,N_2277);
nor U3584 (N_3584,N_2417,N_2535);
nand U3585 (N_3585,N_2536,N_2766);
and U3586 (N_3586,N_2272,N_2282);
or U3587 (N_3587,N_2512,N_2575);
nor U3588 (N_3588,N_2517,N_2556);
or U3589 (N_3589,N_2362,N_2509);
nor U3590 (N_3590,N_2690,N_2938);
or U3591 (N_3591,N_2587,N_2322);
and U3592 (N_3592,N_2356,N_2998);
nor U3593 (N_3593,N_2636,N_2781);
or U3594 (N_3594,N_2664,N_2335);
nand U3595 (N_3595,N_2325,N_2974);
nor U3596 (N_3596,N_2790,N_2717);
and U3597 (N_3597,N_2833,N_2283);
nand U3598 (N_3598,N_2554,N_2669);
or U3599 (N_3599,N_2769,N_2977);
xnor U3600 (N_3600,N_2967,N_2353);
xnor U3601 (N_3601,N_2541,N_2470);
xnor U3602 (N_3602,N_2578,N_2457);
nor U3603 (N_3603,N_2730,N_2315);
nor U3604 (N_3604,N_2934,N_2715);
nand U3605 (N_3605,N_2953,N_2536);
xor U3606 (N_3606,N_2287,N_2286);
and U3607 (N_3607,N_2606,N_2553);
and U3608 (N_3608,N_2550,N_2491);
nand U3609 (N_3609,N_2359,N_2537);
or U3610 (N_3610,N_2711,N_2705);
and U3611 (N_3611,N_2717,N_2333);
nand U3612 (N_3612,N_2255,N_2853);
nor U3613 (N_3613,N_2900,N_2841);
nor U3614 (N_3614,N_2644,N_2523);
or U3615 (N_3615,N_2847,N_2819);
and U3616 (N_3616,N_2404,N_2347);
nand U3617 (N_3617,N_2597,N_2825);
nor U3618 (N_3618,N_2446,N_2407);
nor U3619 (N_3619,N_2771,N_2519);
nand U3620 (N_3620,N_2731,N_2946);
nand U3621 (N_3621,N_2873,N_2759);
nor U3622 (N_3622,N_2708,N_2585);
or U3623 (N_3623,N_2722,N_2752);
nor U3624 (N_3624,N_2821,N_2737);
nand U3625 (N_3625,N_2262,N_2381);
and U3626 (N_3626,N_2950,N_2401);
nand U3627 (N_3627,N_2651,N_2408);
nor U3628 (N_3628,N_2992,N_2292);
nor U3629 (N_3629,N_2748,N_2794);
or U3630 (N_3630,N_2497,N_2409);
and U3631 (N_3631,N_2329,N_2704);
nand U3632 (N_3632,N_2554,N_2732);
nor U3633 (N_3633,N_2749,N_2783);
or U3634 (N_3634,N_2306,N_2618);
nor U3635 (N_3635,N_2281,N_2874);
nor U3636 (N_3636,N_2297,N_2536);
xor U3637 (N_3637,N_2329,N_2741);
nor U3638 (N_3638,N_2815,N_2679);
nor U3639 (N_3639,N_2435,N_2899);
nand U3640 (N_3640,N_2633,N_2336);
nand U3641 (N_3641,N_2758,N_2876);
nand U3642 (N_3642,N_2843,N_2956);
or U3643 (N_3643,N_2865,N_2795);
or U3644 (N_3644,N_2560,N_2913);
and U3645 (N_3645,N_2736,N_2406);
nor U3646 (N_3646,N_2972,N_2865);
and U3647 (N_3647,N_2843,N_2690);
and U3648 (N_3648,N_2313,N_2952);
nor U3649 (N_3649,N_2970,N_2855);
or U3650 (N_3650,N_2886,N_2471);
nor U3651 (N_3651,N_2712,N_2514);
nand U3652 (N_3652,N_2469,N_2344);
or U3653 (N_3653,N_2694,N_2498);
xor U3654 (N_3654,N_2307,N_2750);
and U3655 (N_3655,N_2905,N_2877);
and U3656 (N_3656,N_2628,N_2391);
nand U3657 (N_3657,N_2344,N_2686);
nand U3658 (N_3658,N_2724,N_2753);
and U3659 (N_3659,N_2378,N_2779);
nor U3660 (N_3660,N_2665,N_2298);
nor U3661 (N_3661,N_2831,N_2404);
xnor U3662 (N_3662,N_2539,N_2656);
nand U3663 (N_3663,N_2745,N_2645);
and U3664 (N_3664,N_2830,N_2320);
and U3665 (N_3665,N_2387,N_2270);
nor U3666 (N_3666,N_2899,N_2584);
and U3667 (N_3667,N_2992,N_2402);
nor U3668 (N_3668,N_2268,N_2588);
nand U3669 (N_3669,N_2599,N_2583);
xor U3670 (N_3670,N_2547,N_2727);
nand U3671 (N_3671,N_2736,N_2254);
nor U3672 (N_3672,N_2682,N_2818);
xor U3673 (N_3673,N_2663,N_2599);
nor U3674 (N_3674,N_2651,N_2854);
and U3675 (N_3675,N_2482,N_2298);
nor U3676 (N_3676,N_2456,N_2498);
or U3677 (N_3677,N_2683,N_2367);
and U3678 (N_3678,N_2341,N_2952);
or U3679 (N_3679,N_2253,N_2595);
xor U3680 (N_3680,N_2933,N_2390);
and U3681 (N_3681,N_2639,N_2618);
or U3682 (N_3682,N_2500,N_2365);
and U3683 (N_3683,N_2856,N_2277);
nor U3684 (N_3684,N_2609,N_2801);
or U3685 (N_3685,N_2698,N_2526);
nor U3686 (N_3686,N_2890,N_2530);
nand U3687 (N_3687,N_2296,N_2795);
nand U3688 (N_3688,N_2320,N_2418);
nor U3689 (N_3689,N_2421,N_2535);
and U3690 (N_3690,N_2724,N_2429);
or U3691 (N_3691,N_2564,N_2546);
xor U3692 (N_3692,N_2887,N_2522);
nand U3693 (N_3693,N_2809,N_2326);
or U3694 (N_3694,N_2956,N_2690);
nor U3695 (N_3695,N_2764,N_2251);
nor U3696 (N_3696,N_2850,N_2929);
or U3697 (N_3697,N_2918,N_2817);
or U3698 (N_3698,N_2259,N_2754);
nand U3699 (N_3699,N_2290,N_2495);
or U3700 (N_3700,N_2631,N_2785);
nand U3701 (N_3701,N_2343,N_2826);
or U3702 (N_3702,N_2481,N_2427);
nor U3703 (N_3703,N_2892,N_2535);
nor U3704 (N_3704,N_2820,N_2791);
nor U3705 (N_3705,N_2783,N_2753);
nor U3706 (N_3706,N_2420,N_2306);
and U3707 (N_3707,N_2514,N_2799);
nand U3708 (N_3708,N_2513,N_2536);
nor U3709 (N_3709,N_2470,N_2469);
nand U3710 (N_3710,N_2956,N_2538);
nand U3711 (N_3711,N_2345,N_2508);
and U3712 (N_3712,N_2774,N_2827);
and U3713 (N_3713,N_2323,N_2328);
nor U3714 (N_3714,N_2623,N_2378);
or U3715 (N_3715,N_2960,N_2325);
or U3716 (N_3716,N_2756,N_2918);
nand U3717 (N_3717,N_2805,N_2843);
or U3718 (N_3718,N_2899,N_2594);
and U3719 (N_3719,N_2870,N_2294);
nor U3720 (N_3720,N_2937,N_2469);
xor U3721 (N_3721,N_2957,N_2532);
and U3722 (N_3722,N_2974,N_2965);
or U3723 (N_3723,N_2796,N_2984);
nand U3724 (N_3724,N_2642,N_2509);
nand U3725 (N_3725,N_2720,N_2824);
nand U3726 (N_3726,N_2934,N_2327);
and U3727 (N_3727,N_2930,N_2929);
and U3728 (N_3728,N_2534,N_2794);
and U3729 (N_3729,N_2941,N_2451);
or U3730 (N_3730,N_2864,N_2434);
xor U3731 (N_3731,N_2295,N_2554);
and U3732 (N_3732,N_2643,N_2912);
or U3733 (N_3733,N_2919,N_2894);
nand U3734 (N_3734,N_2840,N_2361);
nor U3735 (N_3735,N_2519,N_2395);
nor U3736 (N_3736,N_2446,N_2677);
nand U3737 (N_3737,N_2800,N_2938);
nand U3738 (N_3738,N_2677,N_2692);
nor U3739 (N_3739,N_2832,N_2924);
nand U3740 (N_3740,N_2538,N_2944);
nand U3741 (N_3741,N_2686,N_2704);
and U3742 (N_3742,N_2824,N_2996);
nor U3743 (N_3743,N_2475,N_2722);
and U3744 (N_3744,N_2641,N_2524);
and U3745 (N_3745,N_2523,N_2516);
nand U3746 (N_3746,N_2596,N_2288);
and U3747 (N_3747,N_2816,N_2683);
or U3748 (N_3748,N_2308,N_2551);
and U3749 (N_3749,N_2540,N_2487);
and U3750 (N_3750,N_3172,N_3079);
or U3751 (N_3751,N_3053,N_3303);
nor U3752 (N_3752,N_3205,N_3318);
nand U3753 (N_3753,N_3319,N_3094);
or U3754 (N_3754,N_3480,N_3173);
and U3755 (N_3755,N_3555,N_3314);
or U3756 (N_3756,N_3166,N_3552);
and U3757 (N_3757,N_3670,N_3295);
nand U3758 (N_3758,N_3710,N_3320);
nand U3759 (N_3759,N_3143,N_3284);
xor U3760 (N_3760,N_3547,N_3666);
xnor U3761 (N_3761,N_3663,N_3713);
xnor U3762 (N_3762,N_3431,N_3656);
nand U3763 (N_3763,N_3133,N_3048);
xor U3764 (N_3764,N_3603,N_3429);
or U3765 (N_3765,N_3466,N_3139);
nor U3766 (N_3766,N_3434,N_3088);
nor U3767 (N_3767,N_3129,N_3646);
and U3768 (N_3768,N_3719,N_3605);
and U3769 (N_3769,N_3575,N_3261);
nor U3770 (N_3770,N_3685,N_3438);
and U3771 (N_3771,N_3359,N_3019);
and U3772 (N_3772,N_3649,N_3706);
nor U3773 (N_3773,N_3563,N_3032);
or U3774 (N_3774,N_3356,N_3215);
and U3775 (N_3775,N_3285,N_3223);
or U3776 (N_3776,N_3152,N_3185);
nor U3777 (N_3777,N_3615,N_3136);
or U3778 (N_3778,N_3745,N_3541);
nor U3779 (N_3779,N_3699,N_3083);
xor U3780 (N_3780,N_3684,N_3391);
nor U3781 (N_3781,N_3569,N_3148);
nand U3782 (N_3782,N_3055,N_3735);
nor U3783 (N_3783,N_3170,N_3457);
and U3784 (N_3784,N_3386,N_3325);
and U3785 (N_3785,N_3105,N_3749);
and U3786 (N_3786,N_3622,N_3114);
and U3787 (N_3787,N_3609,N_3479);
or U3788 (N_3788,N_3729,N_3062);
nand U3789 (N_3789,N_3151,N_3401);
nand U3790 (N_3790,N_3167,N_3257);
nand U3791 (N_3791,N_3056,N_3351);
nor U3792 (N_3792,N_3385,N_3580);
nor U3793 (N_3793,N_3592,N_3157);
and U3794 (N_3794,N_3201,N_3168);
xnor U3795 (N_3795,N_3447,N_3623);
xor U3796 (N_3796,N_3349,N_3428);
or U3797 (N_3797,N_3190,N_3442);
and U3798 (N_3798,N_3472,N_3544);
nand U3799 (N_3799,N_3436,N_3244);
nor U3800 (N_3800,N_3113,N_3263);
and U3801 (N_3801,N_3535,N_3739);
nor U3802 (N_3802,N_3276,N_3637);
nand U3803 (N_3803,N_3695,N_3110);
or U3804 (N_3804,N_3095,N_3581);
nand U3805 (N_3805,N_3724,N_3744);
or U3806 (N_3806,N_3494,N_3577);
nand U3807 (N_3807,N_3028,N_3260);
nor U3808 (N_3808,N_3194,N_3039);
and U3809 (N_3809,N_3002,N_3636);
nand U3810 (N_3810,N_3630,N_3455);
xnor U3811 (N_3811,N_3548,N_3456);
xnor U3812 (N_3812,N_3131,N_3097);
and U3813 (N_3813,N_3366,N_3415);
or U3814 (N_3814,N_3186,N_3049);
and U3815 (N_3815,N_3126,N_3253);
and U3816 (N_3816,N_3045,N_3551);
and U3817 (N_3817,N_3337,N_3362);
nor U3818 (N_3818,N_3732,N_3515);
xnor U3819 (N_3819,N_3388,N_3449);
or U3820 (N_3820,N_3726,N_3367);
or U3821 (N_3821,N_3546,N_3200);
and U3822 (N_3822,N_3071,N_3489);
nand U3823 (N_3823,N_3315,N_3336);
and U3824 (N_3824,N_3274,N_3738);
or U3825 (N_3825,N_3708,N_3321);
nand U3826 (N_3826,N_3207,N_3024);
nand U3827 (N_3827,N_3631,N_3183);
and U3828 (N_3828,N_3254,N_3165);
xor U3829 (N_3829,N_3498,N_3427);
nand U3830 (N_3830,N_3523,N_3397);
nand U3831 (N_3831,N_3103,N_3027);
and U3832 (N_3832,N_3030,N_3217);
and U3833 (N_3833,N_3288,N_3502);
nand U3834 (N_3834,N_3317,N_3237);
and U3835 (N_3835,N_3363,N_3638);
or U3836 (N_3836,N_3218,N_3299);
or U3837 (N_3837,N_3291,N_3704);
or U3838 (N_3838,N_3070,N_3443);
or U3839 (N_3839,N_3490,N_3013);
nand U3840 (N_3840,N_3524,N_3180);
nor U3841 (N_3841,N_3398,N_3270);
nor U3842 (N_3842,N_3379,N_3432);
and U3843 (N_3843,N_3387,N_3423);
nand U3844 (N_3844,N_3350,N_3286);
or U3845 (N_3845,N_3231,N_3554);
or U3846 (N_3846,N_3671,N_3411);
nor U3847 (N_3847,N_3068,N_3216);
and U3848 (N_3848,N_3347,N_3195);
and U3849 (N_3849,N_3196,N_3664);
or U3850 (N_3850,N_3247,N_3723);
nor U3851 (N_3851,N_3702,N_3747);
and U3852 (N_3852,N_3301,N_3677);
nand U3853 (N_3853,N_3283,N_3520);
nand U3854 (N_3854,N_3582,N_3383);
and U3855 (N_3855,N_3694,N_3517);
nand U3856 (N_3856,N_3252,N_3178);
or U3857 (N_3857,N_3731,N_3674);
and U3858 (N_3858,N_3426,N_3175);
nand U3859 (N_3859,N_3403,N_3132);
and U3860 (N_3860,N_3042,N_3437);
nor U3861 (N_3861,N_3146,N_3184);
and U3862 (N_3862,N_3203,N_3565);
nand U3863 (N_3863,N_3331,N_3080);
and U3864 (N_3864,N_3294,N_3102);
nor U3865 (N_3865,N_3163,N_3007);
nand U3866 (N_3866,N_3737,N_3330);
and U3867 (N_3867,N_3158,N_3249);
nand U3868 (N_3868,N_3335,N_3448);
or U3869 (N_3869,N_3292,N_3073);
nor U3870 (N_3870,N_3599,N_3138);
xnor U3871 (N_3871,N_3240,N_3516);
nand U3872 (N_3872,N_3420,N_3134);
and U3873 (N_3873,N_3323,N_3100);
nand U3874 (N_3874,N_3093,N_3632);
nand U3875 (N_3875,N_3643,N_3038);
or U3876 (N_3876,N_3251,N_3587);
nand U3877 (N_3877,N_3115,N_3500);
nor U3878 (N_3878,N_3271,N_3471);
and U3879 (N_3879,N_3589,N_3108);
or U3880 (N_3880,N_3003,N_3698);
or U3881 (N_3881,N_3553,N_3345);
and U3882 (N_3882,N_3084,N_3267);
nor U3883 (N_3883,N_3090,N_3673);
and U3884 (N_3884,N_3235,N_3230);
nand U3885 (N_3885,N_3462,N_3122);
nor U3886 (N_3886,N_3691,N_3504);
nand U3887 (N_3887,N_3680,N_3051);
nor U3888 (N_3888,N_3475,N_3004);
and U3889 (N_3889,N_3338,N_3117);
nand U3890 (N_3890,N_3255,N_3091);
nor U3891 (N_3891,N_3688,N_3141);
or U3892 (N_3892,N_3730,N_3016);
nand U3893 (N_3893,N_3054,N_3177);
or U3894 (N_3894,N_3741,N_3645);
nand U3895 (N_3895,N_3487,N_3574);
or U3896 (N_3896,N_3204,N_3058);
nor U3897 (N_3897,N_3078,N_3302);
nand U3898 (N_3898,N_3140,N_3096);
or U3899 (N_3899,N_3689,N_3369);
and U3900 (N_3900,N_3562,N_3043);
nor U3901 (N_3901,N_3652,N_3259);
nand U3902 (N_3902,N_3705,N_3557);
nand U3903 (N_3903,N_3258,N_3144);
nor U3904 (N_3904,N_3406,N_3586);
or U3905 (N_3905,N_3594,N_3486);
xnor U3906 (N_3906,N_3539,N_3389);
nand U3907 (N_3907,N_3616,N_3282);
nor U3908 (N_3908,N_3300,N_3613);
and U3909 (N_3909,N_3496,N_3460);
and U3910 (N_3910,N_3101,N_3005);
or U3911 (N_3911,N_3085,N_3193);
or U3912 (N_3912,N_3459,N_3568);
nand U3913 (N_3913,N_3069,N_3425);
and U3914 (N_3914,N_3307,N_3125);
nand U3915 (N_3915,N_3561,N_3036);
xnor U3916 (N_3916,N_3346,N_3044);
nand U3917 (N_3917,N_3440,N_3407);
and U3918 (N_3918,N_3208,N_3210);
nor U3919 (N_3919,N_3556,N_3246);
and U3920 (N_3920,N_3275,N_3109);
nor U3921 (N_3921,N_3721,N_3501);
and U3922 (N_3922,N_3000,N_3474);
xnor U3923 (N_3923,N_3687,N_3659);
and U3924 (N_3924,N_3202,N_3463);
and U3925 (N_3925,N_3416,N_3518);
and U3926 (N_3926,N_3527,N_3625);
nor U3927 (N_3927,N_3660,N_3588);
nand U3928 (N_3928,N_3748,N_3430);
or U3929 (N_3929,N_3405,N_3221);
and U3930 (N_3930,N_3650,N_3720);
and U3931 (N_3931,N_3313,N_3099);
and U3932 (N_3932,N_3339,N_3224);
nor U3933 (N_3933,N_3476,N_3644);
or U3934 (N_3934,N_3075,N_3162);
nor U3935 (N_3935,N_3679,N_3392);
or U3936 (N_3936,N_3662,N_3227);
or U3937 (N_3937,N_3268,N_3607);
or U3938 (N_3938,N_3453,N_3365);
and U3939 (N_3939,N_3106,N_3717);
xor U3940 (N_3940,N_3654,N_3454);
nor U3941 (N_3941,N_3278,N_3011);
nor U3942 (N_3942,N_3293,N_3001);
nor U3943 (N_3943,N_3250,N_3226);
and U3944 (N_3944,N_3233,N_3364);
or U3945 (N_3945,N_3701,N_3505);
nand U3946 (N_3946,N_3040,N_3238);
or U3947 (N_3947,N_3481,N_3528);
and U3948 (N_3948,N_3025,N_3409);
or U3949 (N_3949,N_3082,N_3611);
nor U3950 (N_3950,N_3222,N_3718);
and U3951 (N_3951,N_3606,N_3209);
nand U3952 (N_3952,N_3050,N_3711);
nor U3953 (N_3953,N_3290,N_3642);
nand U3954 (N_3954,N_3281,N_3120);
nand U3955 (N_3955,N_3709,N_3297);
and U3956 (N_3956,N_3191,N_3627);
or U3957 (N_3957,N_3121,N_3273);
or U3958 (N_3958,N_3234,N_3412);
or U3959 (N_3959,N_3511,N_3329);
nand U3960 (N_3960,N_3262,N_3006);
nand U3961 (N_3961,N_3452,N_3444);
and U3962 (N_3962,N_3550,N_3031);
nor U3963 (N_3963,N_3700,N_3635);
and U3964 (N_3964,N_3560,N_3107);
and U3965 (N_3965,N_3326,N_3219);
or U3966 (N_3966,N_3488,N_3311);
nor U3967 (N_3967,N_3341,N_3074);
nor U3968 (N_3968,N_3525,N_3641);
or U3969 (N_3969,N_3390,N_3353);
and U3970 (N_3970,N_3026,N_3465);
and U3971 (N_3971,N_3441,N_3161);
nand U3972 (N_3972,N_3601,N_3225);
nor U3973 (N_3973,N_3682,N_3450);
or U3974 (N_3974,N_3057,N_3188);
nor U3975 (N_3975,N_3506,N_3150);
nor U3976 (N_3976,N_3018,N_3265);
or U3977 (N_3977,N_3340,N_3232);
and U3978 (N_3978,N_3707,N_3657);
or U3979 (N_3979,N_3399,N_3012);
nand U3980 (N_3980,N_3064,N_3736);
nand U3981 (N_3981,N_3473,N_3182);
nor U3982 (N_3982,N_3360,N_3316);
xnor U3983 (N_3983,N_3445,N_3681);
nor U3984 (N_3984,N_3600,N_3715);
xor U3985 (N_3985,N_3740,N_3571);
nor U3986 (N_3986,N_3047,N_3352);
nand U3987 (N_3987,N_3692,N_3703);
nor U3988 (N_3988,N_3618,N_3743);
xor U3989 (N_3989,N_3570,N_3483);
or U3990 (N_3990,N_3065,N_3344);
or U3991 (N_3991,N_3154,N_3081);
and U3992 (N_3992,N_3619,N_3361);
or U3993 (N_3993,N_3725,N_3728);
nand U3994 (N_3994,N_3628,N_3417);
nor U3995 (N_3995,N_3066,N_3526);
xnor U3996 (N_3996,N_3010,N_3022);
nand U3997 (N_3997,N_3128,N_3593);
or U3998 (N_3998,N_3742,N_3298);
nand U3999 (N_3999,N_3578,N_3639);
nand U4000 (N_4000,N_3127,N_3585);
or U4001 (N_4001,N_3328,N_3634);
nor U4002 (N_4002,N_3591,N_3212);
and U4003 (N_4003,N_3089,N_3280);
nor U4004 (N_4004,N_3513,N_3176);
xnor U4005 (N_4005,N_3722,N_3327);
nor U4006 (N_4006,N_3029,N_3422);
or U4007 (N_4007,N_3598,N_3714);
and U4008 (N_4008,N_3484,N_3245);
xnor U4009 (N_4009,N_3400,N_3469);
nand U4010 (N_4010,N_3633,N_3312);
and U4011 (N_4011,N_3059,N_3477);
nor U4012 (N_4012,N_3590,N_3495);
nand U4013 (N_4013,N_3533,N_3137);
xnor U4014 (N_4014,N_3375,N_3530);
or U4015 (N_4015,N_3368,N_3174);
nor U4016 (N_4016,N_3531,N_3355);
nor U4017 (N_4017,N_3604,N_3716);
and U4018 (N_4018,N_3264,N_3468);
nor U4019 (N_4019,N_3035,N_3510);
and U4020 (N_4020,N_3072,N_3414);
nand U4021 (N_4021,N_3658,N_3061);
nor U4022 (N_4022,N_3023,N_3086);
nand U4023 (N_4023,N_3690,N_3354);
and U4024 (N_4024,N_3564,N_3380);
nand U4025 (N_4025,N_3647,N_3077);
nor U4026 (N_4026,N_3147,N_3461);
and U4027 (N_4027,N_3624,N_3478);
nor U4028 (N_4028,N_3395,N_3037);
nand U4029 (N_4029,N_3534,N_3197);
nand U4030 (N_4030,N_3381,N_3169);
nand U4031 (N_4031,N_3467,N_3522);
nand U4032 (N_4032,N_3171,N_3651);
or U4033 (N_4033,N_3111,N_3377);
or U4034 (N_4034,N_3015,N_3669);
nand U4035 (N_4035,N_3214,N_3746);
nor U4036 (N_4036,N_3529,N_3503);
or U4037 (N_4037,N_3211,N_3402);
and U4038 (N_4038,N_3597,N_3532);
or U4039 (N_4039,N_3579,N_3334);
and U4040 (N_4040,N_3421,N_3418);
and U4041 (N_4041,N_3566,N_3187);
and U4042 (N_4042,N_3092,N_3009);
nor U4043 (N_4043,N_3608,N_3734);
and U4044 (N_4044,N_3145,N_3493);
or U4045 (N_4045,N_3155,N_3119);
and U4046 (N_4046,N_3378,N_3602);
nand U4047 (N_4047,N_3614,N_3192);
or U4048 (N_4048,N_3371,N_3538);
nor U4049 (N_4049,N_3665,N_3576);
or U4050 (N_4050,N_3289,N_3492);
nand U4051 (N_4051,N_3324,N_3583);
or U4052 (N_4052,N_3159,N_3491);
nor U4053 (N_4053,N_3304,N_3393);
nand U4054 (N_4054,N_3149,N_3676);
nand U4055 (N_4055,N_3668,N_3104);
nand U4056 (N_4056,N_3277,N_3220);
nand U4057 (N_4057,N_3512,N_3266);
nand U4058 (N_4058,N_3308,N_3499);
or U4059 (N_4059,N_3382,N_3439);
nand U4060 (N_4060,N_3686,N_3451);
nor U4061 (N_4061,N_3620,N_3241);
or U4062 (N_4062,N_3584,N_3370);
nor U4063 (N_4063,N_3497,N_3123);
nand U4064 (N_4064,N_3508,N_3228);
and U4065 (N_4065,N_3567,N_3020);
nand U4066 (N_4066,N_3063,N_3612);
or U4067 (N_4067,N_3135,N_3675);
and U4068 (N_4068,N_3348,N_3198);
xnor U4069 (N_4069,N_3482,N_3626);
nand U4070 (N_4070,N_3408,N_3098);
and U4071 (N_4071,N_3446,N_3067);
nand U4072 (N_4072,N_3130,N_3629);
and U4073 (N_4073,N_3309,N_3610);
nand U4074 (N_4074,N_3310,N_3021);
and U4075 (N_4075,N_3655,N_3322);
or U4076 (N_4076,N_3118,N_3573);
and U4077 (N_4077,N_3404,N_3470);
or U4078 (N_4078,N_3374,N_3256);
nand U4079 (N_4079,N_3543,N_3596);
nor U4080 (N_4080,N_3236,N_3521);
nor U4081 (N_4081,N_3153,N_3542);
nor U4082 (N_4082,N_3433,N_3733);
nand U4083 (N_4083,N_3558,N_3199);
xor U4084 (N_4084,N_3559,N_3621);
and U4085 (N_4085,N_3358,N_3424);
nand U4086 (N_4086,N_3343,N_3572);
nand U4087 (N_4087,N_3046,N_3419);
or U4088 (N_4088,N_3357,N_3536);
nor U4089 (N_4089,N_3124,N_3164);
or U4090 (N_4090,N_3248,N_3008);
and U4091 (N_4091,N_3617,N_3667);
and U4092 (N_4092,N_3017,N_3697);
or U4093 (N_4093,N_3239,N_3332);
or U4094 (N_4094,N_3342,N_3076);
or U4095 (N_4095,N_3272,N_3229);
nand U4096 (N_4096,N_3333,N_3060);
nor U4097 (N_4097,N_3384,N_3160);
xnor U4098 (N_4098,N_3112,N_3242);
or U4099 (N_4099,N_3712,N_3519);
nand U4100 (N_4100,N_3435,N_3413);
nor U4101 (N_4101,N_3410,N_3052);
nand U4102 (N_4102,N_3640,N_3116);
nand U4103 (N_4103,N_3464,N_3279);
nor U4104 (N_4104,N_3727,N_3296);
nor U4105 (N_4105,N_3372,N_3033);
or U4106 (N_4106,N_3305,N_3287);
or U4107 (N_4107,N_3509,N_3213);
nor U4108 (N_4108,N_3034,N_3179);
nand U4109 (N_4109,N_3545,N_3014);
xor U4110 (N_4110,N_3206,N_3373);
nor U4111 (N_4111,N_3507,N_3678);
nor U4112 (N_4112,N_3672,N_3661);
nand U4113 (N_4113,N_3142,N_3595);
nand U4114 (N_4114,N_3189,N_3181);
or U4115 (N_4115,N_3394,N_3540);
or U4116 (N_4116,N_3514,N_3041);
nor U4117 (N_4117,N_3396,N_3243);
xnor U4118 (N_4118,N_3653,N_3376);
and U4119 (N_4119,N_3458,N_3537);
nand U4120 (N_4120,N_3648,N_3269);
nand U4121 (N_4121,N_3549,N_3693);
nor U4122 (N_4122,N_3087,N_3696);
nand U4123 (N_4123,N_3683,N_3485);
or U4124 (N_4124,N_3156,N_3306);
nand U4125 (N_4125,N_3563,N_3050);
nand U4126 (N_4126,N_3256,N_3003);
nor U4127 (N_4127,N_3415,N_3074);
and U4128 (N_4128,N_3721,N_3222);
nor U4129 (N_4129,N_3133,N_3619);
nand U4130 (N_4130,N_3265,N_3311);
or U4131 (N_4131,N_3577,N_3665);
nor U4132 (N_4132,N_3526,N_3739);
nor U4133 (N_4133,N_3439,N_3369);
nor U4134 (N_4134,N_3527,N_3605);
nor U4135 (N_4135,N_3012,N_3676);
nor U4136 (N_4136,N_3429,N_3736);
nand U4137 (N_4137,N_3685,N_3688);
and U4138 (N_4138,N_3403,N_3259);
nor U4139 (N_4139,N_3283,N_3685);
or U4140 (N_4140,N_3699,N_3644);
and U4141 (N_4141,N_3498,N_3078);
or U4142 (N_4142,N_3009,N_3206);
or U4143 (N_4143,N_3114,N_3073);
and U4144 (N_4144,N_3226,N_3285);
and U4145 (N_4145,N_3655,N_3278);
nor U4146 (N_4146,N_3437,N_3278);
and U4147 (N_4147,N_3472,N_3470);
or U4148 (N_4148,N_3256,N_3159);
xnor U4149 (N_4149,N_3328,N_3149);
or U4150 (N_4150,N_3363,N_3442);
and U4151 (N_4151,N_3165,N_3613);
and U4152 (N_4152,N_3687,N_3653);
or U4153 (N_4153,N_3628,N_3129);
or U4154 (N_4154,N_3541,N_3383);
nor U4155 (N_4155,N_3312,N_3020);
nand U4156 (N_4156,N_3089,N_3500);
or U4157 (N_4157,N_3464,N_3551);
nor U4158 (N_4158,N_3046,N_3578);
and U4159 (N_4159,N_3628,N_3159);
nor U4160 (N_4160,N_3093,N_3285);
and U4161 (N_4161,N_3321,N_3560);
xor U4162 (N_4162,N_3380,N_3432);
nand U4163 (N_4163,N_3057,N_3609);
and U4164 (N_4164,N_3115,N_3280);
nand U4165 (N_4165,N_3243,N_3177);
nand U4166 (N_4166,N_3514,N_3728);
or U4167 (N_4167,N_3434,N_3297);
and U4168 (N_4168,N_3004,N_3119);
nand U4169 (N_4169,N_3325,N_3257);
or U4170 (N_4170,N_3619,N_3031);
nor U4171 (N_4171,N_3562,N_3299);
nand U4172 (N_4172,N_3059,N_3273);
or U4173 (N_4173,N_3548,N_3296);
and U4174 (N_4174,N_3581,N_3025);
and U4175 (N_4175,N_3661,N_3523);
nand U4176 (N_4176,N_3517,N_3680);
xnor U4177 (N_4177,N_3091,N_3533);
nand U4178 (N_4178,N_3692,N_3715);
xnor U4179 (N_4179,N_3088,N_3107);
xor U4180 (N_4180,N_3223,N_3365);
xnor U4181 (N_4181,N_3735,N_3041);
and U4182 (N_4182,N_3703,N_3165);
nand U4183 (N_4183,N_3487,N_3520);
xnor U4184 (N_4184,N_3042,N_3510);
nor U4185 (N_4185,N_3265,N_3617);
nand U4186 (N_4186,N_3082,N_3740);
and U4187 (N_4187,N_3525,N_3556);
and U4188 (N_4188,N_3731,N_3086);
nor U4189 (N_4189,N_3276,N_3518);
and U4190 (N_4190,N_3048,N_3201);
or U4191 (N_4191,N_3713,N_3307);
nor U4192 (N_4192,N_3440,N_3082);
nand U4193 (N_4193,N_3235,N_3214);
nor U4194 (N_4194,N_3732,N_3502);
nor U4195 (N_4195,N_3347,N_3636);
or U4196 (N_4196,N_3644,N_3241);
and U4197 (N_4197,N_3592,N_3509);
nor U4198 (N_4198,N_3456,N_3260);
or U4199 (N_4199,N_3024,N_3097);
xor U4200 (N_4200,N_3610,N_3662);
and U4201 (N_4201,N_3485,N_3592);
and U4202 (N_4202,N_3714,N_3686);
and U4203 (N_4203,N_3217,N_3615);
nand U4204 (N_4204,N_3465,N_3239);
or U4205 (N_4205,N_3599,N_3548);
and U4206 (N_4206,N_3440,N_3732);
xor U4207 (N_4207,N_3315,N_3093);
nand U4208 (N_4208,N_3669,N_3069);
xor U4209 (N_4209,N_3522,N_3353);
and U4210 (N_4210,N_3162,N_3295);
nand U4211 (N_4211,N_3544,N_3047);
or U4212 (N_4212,N_3386,N_3211);
nand U4213 (N_4213,N_3550,N_3609);
nor U4214 (N_4214,N_3694,N_3447);
nor U4215 (N_4215,N_3613,N_3215);
nor U4216 (N_4216,N_3320,N_3463);
and U4217 (N_4217,N_3520,N_3033);
nand U4218 (N_4218,N_3494,N_3061);
or U4219 (N_4219,N_3468,N_3391);
or U4220 (N_4220,N_3432,N_3505);
or U4221 (N_4221,N_3699,N_3745);
nand U4222 (N_4222,N_3492,N_3440);
nand U4223 (N_4223,N_3276,N_3554);
or U4224 (N_4224,N_3649,N_3594);
and U4225 (N_4225,N_3011,N_3212);
and U4226 (N_4226,N_3441,N_3658);
nor U4227 (N_4227,N_3697,N_3587);
or U4228 (N_4228,N_3142,N_3571);
nor U4229 (N_4229,N_3378,N_3647);
or U4230 (N_4230,N_3160,N_3151);
or U4231 (N_4231,N_3422,N_3078);
and U4232 (N_4232,N_3581,N_3268);
nor U4233 (N_4233,N_3322,N_3425);
nor U4234 (N_4234,N_3051,N_3130);
or U4235 (N_4235,N_3238,N_3490);
xnor U4236 (N_4236,N_3266,N_3595);
and U4237 (N_4237,N_3379,N_3229);
xnor U4238 (N_4238,N_3556,N_3414);
xor U4239 (N_4239,N_3715,N_3531);
nor U4240 (N_4240,N_3336,N_3114);
nand U4241 (N_4241,N_3389,N_3254);
or U4242 (N_4242,N_3705,N_3388);
nand U4243 (N_4243,N_3372,N_3480);
or U4244 (N_4244,N_3218,N_3399);
nor U4245 (N_4245,N_3099,N_3069);
or U4246 (N_4246,N_3494,N_3202);
or U4247 (N_4247,N_3681,N_3074);
nand U4248 (N_4248,N_3134,N_3514);
or U4249 (N_4249,N_3419,N_3054);
or U4250 (N_4250,N_3084,N_3041);
nor U4251 (N_4251,N_3109,N_3564);
nand U4252 (N_4252,N_3503,N_3460);
and U4253 (N_4253,N_3106,N_3095);
or U4254 (N_4254,N_3489,N_3604);
nor U4255 (N_4255,N_3089,N_3583);
or U4256 (N_4256,N_3087,N_3092);
nand U4257 (N_4257,N_3235,N_3019);
nand U4258 (N_4258,N_3286,N_3407);
and U4259 (N_4259,N_3523,N_3368);
xor U4260 (N_4260,N_3609,N_3398);
nor U4261 (N_4261,N_3084,N_3023);
or U4262 (N_4262,N_3451,N_3709);
nor U4263 (N_4263,N_3651,N_3710);
xor U4264 (N_4264,N_3610,N_3248);
nand U4265 (N_4265,N_3605,N_3364);
nand U4266 (N_4266,N_3722,N_3418);
nand U4267 (N_4267,N_3186,N_3207);
nand U4268 (N_4268,N_3643,N_3277);
or U4269 (N_4269,N_3606,N_3225);
and U4270 (N_4270,N_3016,N_3560);
nand U4271 (N_4271,N_3737,N_3345);
nand U4272 (N_4272,N_3215,N_3341);
or U4273 (N_4273,N_3511,N_3328);
and U4274 (N_4274,N_3204,N_3490);
xnor U4275 (N_4275,N_3313,N_3216);
or U4276 (N_4276,N_3435,N_3142);
or U4277 (N_4277,N_3239,N_3389);
nand U4278 (N_4278,N_3213,N_3070);
and U4279 (N_4279,N_3634,N_3290);
and U4280 (N_4280,N_3431,N_3325);
nor U4281 (N_4281,N_3219,N_3593);
and U4282 (N_4282,N_3730,N_3061);
and U4283 (N_4283,N_3154,N_3552);
or U4284 (N_4284,N_3545,N_3425);
nor U4285 (N_4285,N_3599,N_3390);
or U4286 (N_4286,N_3244,N_3565);
or U4287 (N_4287,N_3363,N_3236);
nand U4288 (N_4288,N_3652,N_3478);
and U4289 (N_4289,N_3266,N_3682);
or U4290 (N_4290,N_3411,N_3712);
nand U4291 (N_4291,N_3074,N_3609);
xor U4292 (N_4292,N_3617,N_3582);
nor U4293 (N_4293,N_3660,N_3671);
nor U4294 (N_4294,N_3220,N_3319);
nand U4295 (N_4295,N_3209,N_3111);
nor U4296 (N_4296,N_3609,N_3404);
and U4297 (N_4297,N_3026,N_3643);
and U4298 (N_4298,N_3624,N_3548);
and U4299 (N_4299,N_3329,N_3326);
nand U4300 (N_4300,N_3094,N_3385);
nor U4301 (N_4301,N_3539,N_3034);
nand U4302 (N_4302,N_3313,N_3208);
nor U4303 (N_4303,N_3338,N_3475);
or U4304 (N_4304,N_3593,N_3362);
nor U4305 (N_4305,N_3212,N_3370);
nand U4306 (N_4306,N_3132,N_3404);
and U4307 (N_4307,N_3246,N_3149);
xor U4308 (N_4308,N_3382,N_3228);
nor U4309 (N_4309,N_3452,N_3730);
nand U4310 (N_4310,N_3176,N_3511);
and U4311 (N_4311,N_3223,N_3362);
nor U4312 (N_4312,N_3730,N_3629);
nand U4313 (N_4313,N_3085,N_3215);
nor U4314 (N_4314,N_3317,N_3221);
and U4315 (N_4315,N_3641,N_3034);
or U4316 (N_4316,N_3502,N_3118);
xor U4317 (N_4317,N_3499,N_3733);
or U4318 (N_4318,N_3295,N_3490);
nor U4319 (N_4319,N_3139,N_3701);
nand U4320 (N_4320,N_3227,N_3630);
and U4321 (N_4321,N_3107,N_3042);
and U4322 (N_4322,N_3523,N_3641);
xnor U4323 (N_4323,N_3631,N_3323);
or U4324 (N_4324,N_3225,N_3623);
nor U4325 (N_4325,N_3656,N_3274);
xnor U4326 (N_4326,N_3605,N_3413);
nor U4327 (N_4327,N_3338,N_3711);
nor U4328 (N_4328,N_3309,N_3505);
or U4329 (N_4329,N_3016,N_3024);
nor U4330 (N_4330,N_3619,N_3179);
and U4331 (N_4331,N_3153,N_3522);
nor U4332 (N_4332,N_3730,N_3359);
nor U4333 (N_4333,N_3336,N_3127);
nor U4334 (N_4334,N_3639,N_3443);
or U4335 (N_4335,N_3396,N_3467);
nor U4336 (N_4336,N_3171,N_3527);
nand U4337 (N_4337,N_3095,N_3734);
xnor U4338 (N_4338,N_3156,N_3639);
or U4339 (N_4339,N_3440,N_3141);
nand U4340 (N_4340,N_3153,N_3540);
nor U4341 (N_4341,N_3099,N_3296);
xnor U4342 (N_4342,N_3587,N_3052);
or U4343 (N_4343,N_3577,N_3556);
and U4344 (N_4344,N_3383,N_3722);
nor U4345 (N_4345,N_3347,N_3043);
and U4346 (N_4346,N_3676,N_3048);
nor U4347 (N_4347,N_3558,N_3399);
or U4348 (N_4348,N_3677,N_3144);
nor U4349 (N_4349,N_3239,N_3011);
and U4350 (N_4350,N_3014,N_3343);
or U4351 (N_4351,N_3173,N_3592);
nand U4352 (N_4352,N_3448,N_3635);
nor U4353 (N_4353,N_3290,N_3725);
nor U4354 (N_4354,N_3199,N_3734);
nor U4355 (N_4355,N_3599,N_3160);
or U4356 (N_4356,N_3013,N_3439);
and U4357 (N_4357,N_3415,N_3503);
and U4358 (N_4358,N_3398,N_3339);
nor U4359 (N_4359,N_3633,N_3322);
nand U4360 (N_4360,N_3402,N_3135);
nand U4361 (N_4361,N_3315,N_3281);
and U4362 (N_4362,N_3093,N_3378);
and U4363 (N_4363,N_3370,N_3437);
nor U4364 (N_4364,N_3212,N_3548);
or U4365 (N_4365,N_3068,N_3222);
xnor U4366 (N_4366,N_3098,N_3222);
nor U4367 (N_4367,N_3527,N_3720);
or U4368 (N_4368,N_3143,N_3381);
and U4369 (N_4369,N_3252,N_3053);
and U4370 (N_4370,N_3345,N_3336);
nor U4371 (N_4371,N_3736,N_3639);
or U4372 (N_4372,N_3517,N_3525);
nand U4373 (N_4373,N_3298,N_3673);
nand U4374 (N_4374,N_3323,N_3497);
nand U4375 (N_4375,N_3149,N_3099);
or U4376 (N_4376,N_3326,N_3191);
or U4377 (N_4377,N_3331,N_3460);
nor U4378 (N_4378,N_3095,N_3298);
xor U4379 (N_4379,N_3666,N_3324);
or U4380 (N_4380,N_3360,N_3259);
and U4381 (N_4381,N_3482,N_3363);
or U4382 (N_4382,N_3016,N_3667);
and U4383 (N_4383,N_3094,N_3170);
or U4384 (N_4384,N_3408,N_3687);
or U4385 (N_4385,N_3116,N_3338);
or U4386 (N_4386,N_3369,N_3457);
and U4387 (N_4387,N_3311,N_3282);
nand U4388 (N_4388,N_3284,N_3174);
nand U4389 (N_4389,N_3534,N_3725);
nand U4390 (N_4390,N_3502,N_3623);
and U4391 (N_4391,N_3416,N_3460);
or U4392 (N_4392,N_3244,N_3320);
nor U4393 (N_4393,N_3097,N_3353);
and U4394 (N_4394,N_3513,N_3642);
and U4395 (N_4395,N_3693,N_3662);
nor U4396 (N_4396,N_3549,N_3586);
nand U4397 (N_4397,N_3459,N_3461);
or U4398 (N_4398,N_3362,N_3399);
and U4399 (N_4399,N_3414,N_3082);
and U4400 (N_4400,N_3650,N_3463);
nor U4401 (N_4401,N_3118,N_3112);
nor U4402 (N_4402,N_3379,N_3354);
and U4403 (N_4403,N_3091,N_3127);
and U4404 (N_4404,N_3439,N_3637);
nand U4405 (N_4405,N_3660,N_3112);
or U4406 (N_4406,N_3029,N_3156);
and U4407 (N_4407,N_3127,N_3459);
nand U4408 (N_4408,N_3007,N_3016);
xor U4409 (N_4409,N_3301,N_3355);
nor U4410 (N_4410,N_3113,N_3480);
nand U4411 (N_4411,N_3478,N_3062);
nor U4412 (N_4412,N_3589,N_3442);
nand U4413 (N_4413,N_3014,N_3413);
and U4414 (N_4414,N_3612,N_3460);
nor U4415 (N_4415,N_3344,N_3505);
and U4416 (N_4416,N_3074,N_3498);
and U4417 (N_4417,N_3546,N_3064);
nand U4418 (N_4418,N_3435,N_3536);
and U4419 (N_4419,N_3364,N_3511);
xnor U4420 (N_4420,N_3286,N_3137);
xnor U4421 (N_4421,N_3149,N_3384);
nand U4422 (N_4422,N_3747,N_3363);
or U4423 (N_4423,N_3103,N_3276);
nor U4424 (N_4424,N_3629,N_3128);
nor U4425 (N_4425,N_3625,N_3566);
nand U4426 (N_4426,N_3608,N_3596);
xor U4427 (N_4427,N_3336,N_3676);
or U4428 (N_4428,N_3021,N_3174);
or U4429 (N_4429,N_3083,N_3030);
and U4430 (N_4430,N_3453,N_3039);
and U4431 (N_4431,N_3079,N_3315);
or U4432 (N_4432,N_3673,N_3354);
or U4433 (N_4433,N_3191,N_3230);
nor U4434 (N_4434,N_3104,N_3463);
xor U4435 (N_4435,N_3318,N_3651);
xor U4436 (N_4436,N_3726,N_3747);
or U4437 (N_4437,N_3735,N_3595);
and U4438 (N_4438,N_3086,N_3104);
nand U4439 (N_4439,N_3253,N_3497);
and U4440 (N_4440,N_3289,N_3490);
xor U4441 (N_4441,N_3515,N_3312);
or U4442 (N_4442,N_3197,N_3681);
nor U4443 (N_4443,N_3568,N_3163);
nand U4444 (N_4444,N_3080,N_3733);
nand U4445 (N_4445,N_3291,N_3277);
nor U4446 (N_4446,N_3739,N_3028);
xor U4447 (N_4447,N_3033,N_3086);
xnor U4448 (N_4448,N_3246,N_3513);
or U4449 (N_4449,N_3182,N_3534);
or U4450 (N_4450,N_3621,N_3335);
nand U4451 (N_4451,N_3329,N_3421);
nand U4452 (N_4452,N_3682,N_3551);
nand U4453 (N_4453,N_3121,N_3559);
nor U4454 (N_4454,N_3185,N_3620);
xor U4455 (N_4455,N_3457,N_3648);
and U4456 (N_4456,N_3556,N_3096);
nand U4457 (N_4457,N_3388,N_3163);
and U4458 (N_4458,N_3026,N_3077);
nand U4459 (N_4459,N_3045,N_3424);
nor U4460 (N_4460,N_3078,N_3547);
nor U4461 (N_4461,N_3041,N_3444);
and U4462 (N_4462,N_3053,N_3619);
nor U4463 (N_4463,N_3567,N_3534);
nor U4464 (N_4464,N_3249,N_3167);
nor U4465 (N_4465,N_3239,N_3302);
nor U4466 (N_4466,N_3351,N_3128);
xnor U4467 (N_4467,N_3498,N_3028);
and U4468 (N_4468,N_3201,N_3280);
xor U4469 (N_4469,N_3739,N_3748);
nor U4470 (N_4470,N_3245,N_3362);
nor U4471 (N_4471,N_3556,N_3477);
and U4472 (N_4472,N_3442,N_3551);
or U4473 (N_4473,N_3684,N_3697);
and U4474 (N_4474,N_3617,N_3559);
or U4475 (N_4475,N_3268,N_3587);
or U4476 (N_4476,N_3134,N_3392);
and U4477 (N_4477,N_3513,N_3492);
and U4478 (N_4478,N_3286,N_3686);
nand U4479 (N_4479,N_3087,N_3523);
nand U4480 (N_4480,N_3077,N_3275);
or U4481 (N_4481,N_3066,N_3263);
or U4482 (N_4482,N_3010,N_3737);
xnor U4483 (N_4483,N_3248,N_3692);
or U4484 (N_4484,N_3376,N_3138);
or U4485 (N_4485,N_3592,N_3318);
xnor U4486 (N_4486,N_3360,N_3653);
or U4487 (N_4487,N_3357,N_3499);
xor U4488 (N_4488,N_3668,N_3053);
or U4489 (N_4489,N_3413,N_3609);
nor U4490 (N_4490,N_3028,N_3503);
or U4491 (N_4491,N_3490,N_3300);
or U4492 (N_4492,N_3164,N_3062);
and U4493 (N_4493,N_3035,N_3066);
nand U4494 (N_4494,N_3486,N_3298);
and U4495 (N_4495,N_3071,N_3524);
nor U4496 (N_4496,N_3337,N_3389);
and U4497 (N_4497,N_3629,N_3628);
or U4498 (N_4498,N_3110,N_3369);
nand U4499 (N_4499,N_3671,N_3000);
and U4500 (N_4500,N_4492,N_4242);
or U4501 (N_4501,N_4418,N_4357);
nand U4502 (N_4502,N_3825,N_4459);
and U4503 (N_4503,N_3764,N_4140);
nand U4504 (N_4504,N_3941,N_4384);
and U4505 (N_4505,N_3810,N_3828);
nand U4506 (N_4506,N_4283,N_4158);
xnor U4507 (N_4507,N_4008,N_4135);
and U4508 (N_4508,N_4007,N_4347);
or U4509 (N_4509,N_4106,N_4236);
or U4510 (N_4510,N_4373,N_4289);
and U4511 (N_4511,N_4467,N_4068);
or U4512 (N_4512,N_4063,N_4225);
nand U4513 (N_4513,N_3847,N_4235);
or U4514 (N_4514,N_4443,N_4109);
nand U4515 (N_4515,N_4339,N_4138);
and U4516 (N_4516,N_4082,N_4209);
nor U4517 (N_4517,N_3814,N_3800);
and U4518 (N_4518,N_4487,N_3774);
nor U4519 (N_4519,N_4496,N_4305);
and U4520 (N_4520,N_3874,N_4057);
and U4521 (N_4521,N_4491,N_4108);
xnor U4522 (N_4522,N_4254,N_4243);
or U4523 (N_4523,N_4200,N_4121);
and U4524 (N_4524,N_3899,N_3805);
and U4525 (N_4525,N_3753,N_4388);
nor U4526 (N_4526,N_4086,N_3757);
xnor U4527 (N_4527,N_3913,N_4326);
xnor U4528 (N_4528,N_3851,N_4398);
nand U4529 (N_4529,N_4294,N_4119);
or U4530 (N_4530,N_4032,N_3832);
nor U4531 (N_4531,N_3750,N_3813);
nand U4532 (N_4532,N_3924,N_4221);
nor U4533 (N_4533,N_3815,N_4027);
nor U4534 (N_4534,N_4197,N_4075);
nor U4535 (N_4535,N_4081,N_3817);
nand U4536 (N_4536,N_4462,N_4178);
or U4537 (N_4537,N_3868,N_4447);
nand U4538 (N_4538,N_4295,N_4296);
nor U4539 (N_4539,N_3793,N_4275);
nand U4540 (N_4540,N_4441,N_4228);
xnor U4541 (N_4541,N_4037,N_4132);
and U4542 (N_4542,N_4021,N_3752);
and U4543 (N_4543,N_4160,N_4202);
or U4544 (N_4544,N_4499,N_4133);
nor U4545 (N_4545,N_4488,N_4372);
nor U4546 (N_4546,N_4024,N_4039);
or U4547 (N_4547,N_4371,N_4205);
and U4548 (N_4548,N_3782,N_3838);
nor U4549 (N_4549,N_4169,N_3910);
nor U4550 (N_4550,N_4185,N_4028);
or U4551 (N_4551,N_3806,N_4446);
nand U4552 (N_4552,N_4153,N_3863);
or U4553 (N_4553,N_4097,N_4286);
or U4554 (N_4554,N_3783,N_3890);
nand U4555 (N_4555,N_4117,N_3820);
nor U4556 (N_4556,N_3798,N_4461);
nand U4557 (N_4557,N_4203,N_4112);
and U4558 (N_4558,N_3875,N_4310);
and U4559 (N_4559,N_4293,N_4183);
or U4560 (N_4560,N_3984,N_3835);
and U4561 (N_4561,N_3902,N_4216);
nand U4562 (N_4562,N_4247,N_4069);
nand U4563 (N_4563,N_4052,N_3988);
nand U4564 (N_4564,N_3892,N_4155);
nand U4565 (N_4565,N_4479,N_4448);
and U4566 (N_4566,N_4046,N_4167);
nand U4567 (N_4567,N_4374,N_4012);
xor U4568 (N_4568,N_3856,N_4055);
nand U4569 (N_4569,N_4300,N_3778);
nand U4570 (N_4570,N_4279,N_4166);
or U4571 (N_4571,N_4278,N_3865);
nand U4572 (N_4572,N_4192,N_4437);
nor U4573 (N_4573,N_4299,N_3836);
nor U4574 (N_4574,N_3975,N_4190);
nor U4575 (N_4575,N_4451,N_4490);
nand U4576 (N_4576,N_4266,N_3969);
and U4577 (N_4577,N_4274,N_3982);
or U4578 (N_4578,N_3827,N_4114);
nor U4579 (N_4579,N_4429,N_4474);
and U4580 (N_4580,N_3760,N_3853);
and U4581 (N_4581,N_4250,N_4379);
nand U4582 (N_4582,N_3769,N_4297);
xnor U4583 (N_4583,N_3844,N_4292);
nand U4584 (N_4584,N_3862,N_4449);
and U4585 (N_4585,N_4147,N_3861);
nor U4586 (N_4586,N_3966,N_3879);
nand U4587 (N_4587,N_4195,N_4395);
nand U4588 (N_4588,N_3873,N_3963);
xor U4589 (N_4589,N_3822,N_4409);
and U4590 (N_4590,N_4270,N_3766);
nand U4591 (N_4591,N_3979,N_4025);
nand U4592 (N_4592,N_4497,N_3953);
or U4593 (N_4593,N_3944,N_4005);
and U4594 (N_4594,N_4423,N_4337);
and U4595 (N_4595,N_3762,N_4103);
and U4596 (N_4596,N_3765,N_4466);
nand U4597 (N_4597,N_4102,N_4092);
and U4598 (N_4598,N_3903,N_4416);
and U4599 (N_4599,N_4201,N_3916);
nor U4600 (N_4600,N_4218,N_4468);
and U4601 (N_4601,N_3780,N_4498);
nand U4602 (N_4602,N_4356,N_3809);
and U4603 (N_4603,N_3895,N_4420);
and U4604 (N_4604,N_4071,N_4436);
nand U4605 (N_4605,N_4177,N_4208);
xnor U4606 (N_4606,N_4115,N_4353);
and U4607 (N_4607,N_4091,N_3768);
and U4608 (N_4608,N_4306,N_4058);
xnor U4609 (N_4609,N_3877,N_4127);
or U4610 (N_4610,N_4062,N_4471);
nand U4611 (N_4611,N_4405,N_3808);
nor U4612 (N_4612,N_3907,N_4431);
and U4613 (N_4613,N_4029,N_3787);
nor U4614 (N_4614,N_4036,N_4085);
xnor U4615 (N_4615,N_3839,N_3962);
and U4616 (N_4616,N_4181,N_4164);
nand U4617 (N_4617,N_4146,N_4249);
and U4618 (N_4618,N_3818,N_4302);
and U4619 (N_4619,N_3990,N_4013);
nand U4620 (N_4620,N_4060,N_4154);
xor U4621 (N_4621,N_3830,N_3755);
nor U4622 (N_4622,N_4308,N_4022);
nor U4623 (N_4623,N_4330,N_4126);
xor U4624 (N_4624,N_4172,N_3926);
and U4625 (N_4625,N_3860,N_3758);
and U4626 (N_4626,N_3970,N_3871);
nor U4627 (N_4627,N_4244,N_4457);
nand U4628 (N_4628,N_4311,N_4199);
and U4629 (N_4629,N_4397,N_4137);
and U4630 (N_4630,N_4333,N_3850);
or U4631 (N_4631,N_4174,N_4282);
or U4632 (N_4632,N_3854,N_4232);
or U4633 (N_4633,N_4433,N_4262);
or U4634 (N_4634,N_4042,N_4000);
nand U4635 (N_4635,N_4322,N_3837);
or U4636 (N_4636,N_4442,N_4224);
or U4637 (N_4637,N_3812,N_3884);
nand U4638 (N_4638,N_3952,N_4239);
or U4639 (N_4639,N_4298,N_4041);
and U4640 (N_4640,N_3869,N_4168);
and U4641 (N_4641,N_4328,N_4156);
nor U4642 (N_4642,N_4151,N_4145);
nand U4643 (N_4643,N_3824,N_4482);
and U4644 (N_4644,N_3949,N_4403);
xor U4645 (N_4645,N_3876,N_3788);
nor U4646 (N_4646,N_4040,N_4413);
nor U4647 (N_4647,N_3819,N_4453);
nand U4648 (N_4648,N_3936,N_3846);
xor U4649 (N_4649,N_4125,N_4348);
nor U4650 (N_4650,N_4455,N_4342);
and U4651 (N_4651,N_3789,N_4354);
xor U4652 (N_4652,N_4495,N_4408);
xnor U4653 (N_4653,N_4309,N_4229);
or U4654 (N_4654,N_3772,N_4401);
nor U4655 (N_4655,N_4314,N_3909);
nor U4656 (N_4656,N_4268,N_3914);
nor U4657 (N_4657,N_4385,N_3870);
and U4658 (N_4658,N_3954,N_3786);
nand U4659 (N_4659,N_3947,N_4198);
and U4660 (N_4660,N_4271,N_4179);
nor U4661 (N_4661,N_4051,N_4233);
xnor U4662 (N_4662,N_3843,N_3840);
and U4663 (N_4663,N_4020,N_4157);
nor U4664 (N_4664,N_4325,N_3826);
or U4665 (N_4665,N_3905,N_4445);
nand U4666 (N_4666,N_4226,N_4427);
nand U4667 (N_4667,N_4281,N_4318);
or U4668 (N_4668,N_4422,N_4350);
or U4669 (N_4669,N_3933,N_4186);
nor U4670 (N_4670,N_3833,N_4044);
xnor U4671 (N_4671,N_4316,N_4359);
xnor U4672 (N_4672,N_4470,N_3849);
or U4673 (N_4673,N_4362,N_4483);
nand U4674 (N_4674,N_3938,N_3911);
nand U4675 (N_4675,N_4360,N_4273);
nand U4676 (N_4676,N_4258,N_3790);
xor U4677 (N_4677,N_4463,N_4452);
nand U4678 (N_4678,N_4473,N_4241);
xnor U4679 (N_4679,N_4043,N_3930);
nor U4680 (N_4680,N_4159,N_3928);
nor U4681 (N_4681,N_4180,N_4149);
or U4682 (N_4682,N_4187,N_4381);
nand U4683 (N_4683,N_3784,N_4368);
nand U4684 (N_4684,N_4079,N_3891);
nand U4685 (N_4685,N_3794,N_4400);
and U4686 (N_4686,N_4004,N_4340);
nand U4687 (N_4687,N_4345,N_4240);
nor U4688 (N_4688,N_4313,N_4394);
nand U4689 (N_4689,N_3959,N_4072);
or U4690 (N_4690,N_3823,N_4475);
nand U4691 (N_4691,N_4128,N_4001);
or U4692 (N_4692,N_4033,N_3932);
nor U4693 (N_4693,N_4349,N_4494);
or U4694 (N_4694,N_4280,N_4095);
and U4695 (N_4695,N_3881,N_3977);
or U4696 (N_4696,N_3857,N_4404);
xor U4697 (N_4697,N_3864,N_4272);
nor U4698 (N_4698,N_4321,N_4438);
or U4699 (N_4699,N_4018,N_4257);
nand U4700 (N_4700,N_4396,N_3971);
and U4701 (N_4701,N_3915,N_3796);
nand U4702 (N_4702,N_4113,N_4074);
or U4703 (N_4703,N_4392,N_3751);
xor U4704 (N_4704,N_3931,N_4426);
nor U4705 (N_4705,N_4141,N_4087);
nor U4706 (N_4706,N_4261,N_3978);
nor U4707 (N_4707,N_4331,N_3807);
or U4708 (N_4708,N_4458,N_4231);
and U4709 (N_4709,N_4376,N_4263);
nor U4710 (N_4710,N_4152,N_4324);
and U4711 (N_4711,N_4084,N_4425);
nor U4712 (N_4712,N_4026,N_4134);
nor U4713 (N_4713,N_4323,N_3991);
and U4714 (N_4714,N_3995,N_4377);
nor U4715 (N_4715,N_4104,N_4329);
or U4716 (N_4716,N_4212,N_4450);
nand U4717 (N_4717,N_3945,N_3918);
nor U4718 (N_4718,N_4089,N_3779);
or U4719 (N_4719,N_4485,N_3872);
nor U4720 (N_4720,N_4142,N_3802);
or U4721 (N_4721,N_4378,N_4415);
and U4722 (N_4722,N_4288,N_4066);
nand U4723 (N_4723,N_3785,N_4122);
nand U4724 (N_4724,N_4213,N_4383);
nand U4725 (N_4725,N_3948,N_4162);
or U4726 (N_4726,N_3957,N_4171);
or U4727 (N_4727,N_3898,N_3883);
and U4728 (N_4728,N_4129,N_3934);
nor U4729 (N_4729,N_4204,N_3972);
nor U4730 (N_4730,N_4364,N_3770);
or U4731 (N_4731,N_3773,N_4456);
or U4732 (N_4732,N_3956,N_3834);
xnor U4733 (N_4733,N_4303,N_4386);
nand U4734 (N_4734,N_4493,N_3893);
nand U4735 (N_4735,N_4019,N_4419);
nor U4736 (N_4736,N_3803,N_4207);
and U4737 (N_4737,N_3763,N_3937);
nand U4738 (N_4738,N_4034,N_4284);
or U4739 (N_4739,N_4355,N_4143);
nor U4740 (N_4740,N_4038,N_4375);
nand U4741 (N_4741,N_4111,N_3940);
nand U4742 (N_4742,N_3888,N_4173);
and U4743 (N_4743,N_4070,N_3961);
xnor U4744 (N_4744,N_4315,N_4237);
nand U4745 (N_4745,N_3831,N_4469);
or U4746 (N_4746,N_4460,N_3885);
xnor U4747 (N_4747,N_4105,N_3829);
and U4748 (N_4748,N_3999,N_4214);
or U4749 (N_4749,N_3929,N_3998);
xor U4750 (N_4750,N_4402,N_3922);
and U4751 (N_4751,N_4002,N_4163);
and U4752 (N_4752,N_3882,N_4053);
and U4753 (N_4753,N_4399,N_4370);
and U4754 (N_4754,N_4107,N_3921);
nand U4755 (N_4755,N_3965,N_4206);
nand U4756 (N_4756,N_3908,N_3775);
or U4757 (N_4757,N_4477,N_4428);
nand U4758 (N_4758,N_4454,N_4480);
nand U4759 (N_4759,N_4335,N_4389);
xnor U4760 (N_4760,N_4253,N_4170);
and U4761 (N_4761,N_3901,N_4031);
nand U4762 (N_4762,N_4077,N_3951);
nand U4763 (N_4763,N_3950,N_4245);
or U4764 (N_4764,N_4338,N_4083);
nor U4765 (N_4765,N_4116,N_4352);
and U4766 (N_4766,N_4098,N_4317);
and U4767 (N_4767,N_4435,N_4176);
or U4768 (N_4768,N_4035,N_4045);
nand U4769 (N_4769,N_3811,N_4067);
and U4770 (N_4770,N_3859,N_3958);
xnor U4771 (N_4771,N_4100,N_4434);
and U4772 (N_4772,N_3912,N_4161);
nor U4773 (N_4773,N_3904,N_4217);
and U4774 (N_4774,N_4439,N_4367);
xnor U4775 (N_4775,N_4489,N_3985);
and U4776 (N_4776,N_4227,N_4124);
and U4777 (N_4777,N_3993,N_4059);
nor U4778 (N_4778,N_3974,N_4090);
nor U4779 (N_4779,N_3842,N_4110);
or U4780 (N_4780,N_4312,N_3935);
nor U4781 (N_4781,N_3976,N_4332);
nand U4782 (N_4782,N_4363,N_4136);
and U4783 (N_4783,N_3756,N_3797);
nor U4784 (N_4784,N_4030,N_3989);
nand U4785 (N_4785,N_4343,N_4391);
nor U4786 (N_4786,N_4088,N_4073);
or U4787 (N_4787,N_4476,N_4011);
nor U4788 (N_4788,N_3767,N_4016);
or U4789 (N_4789,N_4341,N_4056);
or U4790 (N_4790,N_3858,N_4320);
nor U4791 (N_4791,N_3896,N_3841);
nor U4792 (N_4792,N_4064,N_4050);
and U4793 (N_4793,N_4220,N_4382);
xor U4794 (N_4794,N_3761,N_4259);
nand U4795 (N_4795,N_3927,N_4023);
or U4796 (N_4796,N_4246,N_4410);
or U4797 (N_4797,N_4265,N_4150);
nand U4798 (N_4798,N_4078,N_3816);
and U4799 (N_4799,N_3923,N_4215);
or U4800 (N_4800,N_3759,N_4211);
nor U4801 (N_4801,N_4234,N_3946);
and U4802 (N_4802,N_3799,N_4061);
nor U4803 (N_4803,N_3925,N_3866);
or U4804 (N_4804,N_4290,N_3821);
xor U4805 (N_4805,N_3801,N_4464);
or U4806 (N_4806,N_3996,N_3771);
nor U4807 (N_4807,N_4365,N_4264);
xnor U4808 (N_4808,N_3889,N_3777);
nand U4809 (N_4809,N_4049,N_4344);
and U4810 (N_4810,N_4120,N_3973);
nand U4811 (N_4811,N_4047,N_3919);
nor U4812 (N_4812,N_4484,N_4380);
nand U4813 (N_4813,N_4118,N_3994);
nand U4814 (N_4814,N_4387,N_4346);
nand U4815 (N_4815,N_4248,N_4251);
nor U4816 (N_4816,N_3880,N_4131);
nand U4817 (N_4817,N_4424,N_4210);
and U4818 (N_4818,N_4196,N_4193);
and U4819 (N_4819,N_4076,N_4319);
nor U4820 (N_4820,N_3983,N_4444);
nor U4821 (N_4821,N_4017,N_4014);
and U4822 (N_4822,N_4123,N_3845);
and U4823 (N_4823,N_4361,N_3867);
and U4824 (N_4824,N_4291,N_4407);
nor U4825 (N_4825,N_3920,N_4358);
nor U4826 (N_4826,N_3900,N_4276);
or U4827 (N_4827,N_4277,N_3968);
nor U4828 (N_4828,N_4430,N_4465);
nor U4829 (N_4829,N_4165,N_4189);
nor U4830 (N_4830,N_4238,N_3776);
nor U4831 (N_4831,N_4182,N_4094);
or U4832 (N_4832,N_3997,N_4412);
nand U4833 (N_4833,N_4054,N_4010);
nor U4834 (N_4834,N_4369,N_3886);
and U4835 (N_4835,N_3781,N_3791);
and U4836 (N_4836,N_4003,N_4406);
xnor U4837 (N_4837,N_4015,N_4336);
nor U4838 (N_4838,N_3878,N_4269);
nand U4839 (N_4839,N_4006,N_4256);
nand U4840 (N_4840,N_3967,N_4219);
nand U4841 (N_4841,N_4194,N_4304);
or U4842 (N_4842,N_4417,N_4301);
nor U4843 (N_4843,N_3897,N_4260);
and U4844 (N_4844,N_3955,N_3906);
xor U4845 (N_4845,N_4080,N_4223);
and U4846 (N_4846,N_4101,N_4188);
nor U4847 (N_4847,N_4139,N_3754);
nand U4848 (N_4848,N_4307,N_3804);
nor U4849 (N_4849,N_4093,N_4065);
xor U4850 (N_4850,N_3942,N_3917);
xor U4851 (N_4851,N_3792,N_4148);
or U4852 (N_4852,N_3964,N_4414);
and U4853 (N_4853,N_4287,N_4130);
nor U4854 (N_4854,N_4144,N_4440);
nand U4855 (N_4855,N_4481,N_4421);
nor U4856 (N_4856,N_3848,N_3981);
and U4857 (N_4857,N_3855,N_4486);
or U4858 (N_4858,N_4175,N_3943);
and U4859 (N_4859,N_3992,N_4184);
nor U4860 (N_4860,N_3894,N_3795);
nor U4861 (N_4861,N_4366,N_4267);
or U4862 (N_4862,N_4252,N_3987);
and U4863 (N_4863,N_4009,N_3960);
nand U4864 (N_4864,N_4327,N_4048);
or U4865 (N_4865,N_4334,N_3986);
and U4866 (N_4866,N_4096,N_4411);
xnor U4867 (N_4867,N_4099,N_4191);
nand U4868 (N_4868,N_4285,N_4222);
or U4869 (N_4869,N_3852,N_4390);
or U4870 (N_4870,N_4472,N_3887);
nor U4871 (N_4871,N_4230,N_4255);
and U4872 (N_4872,N_4478,N_4351);
or U4873 (N_4873,N_4393,N_4432);
nand U4874 (N_4874,N_3939,N_3980);
xor U4875 (N_4875,N_4061,N_3806);
or U4876 (N_4876,N_3921,N_4096);
or U4877 (N_4877,N_4202,N_4376);
nor U4878 (N_4878,N_4069,N_4243);
nor U4879 (N_4879,N_4262,N_3760);
or U4880 (N_4880,N_3912,N_3772);
nor U4881 (N_4881,N_4474,N_4144);
xor U4882 (N_4882,N_4239,N_4194);
nand U4883 (N_4883,N_4361,N_3798);
nor U4884 (N_4884,N_4127,N_4213);
nor U4885 (N_4885,N_4286,N_3988);
nor U4886 (N_4886,N_4225,N_4275);
or U4887 (N_4887,N_3992,N_3939);
and U4888 (N_4888,N_3993,N_4405);
nor U4889 (N_4889,N_4367,N_4148);
xor U4890 (N_4890,N_4179,N_3813);
nor U4891 (N_4891,N_4310,N_3806);
or U4892 (N_4892,N_3931,N_4210);
nor U4893 (N_4893,N_4220,N_4014);
nor U4894 (N_4894,N_4189,N_3911);
nor U4895 (N_4895,N_4402,N_4457);
nor U4896 (N_4896,N_3802,N_3936);
and U4897 (N_4897,N_3800,N_3829);
nand U4898 (N_4898,N_4050,N_4156);
and U4899 (N_4899,N_4404,N_3828);
nor U4900 (N_4900,N_3857,N_4200);
nor U4901 (N_4901,N_4325,N_3938);
nand U4902 (N_4902,N_3866,N_4477);
or U4903 (N_4903,N_4351,N_4401);
and U4904 (N_4904,N_3769,N_4379);
or U4905 (N_4905,N_3898,N_4187);
nor U4906 (N_4906,N_4101,N_4044);
xnor U4907 (N_4907,N_4099,N_3879);
nor U4908 (N_4908,N_4413,N_4316);
and U4909 (N_4909,N_3894,N_3862);
and U4910 (N_4910,N_4333,N_4435);
xnor U4911 (N_4911,N_3858,N_4463);
and U4912 (N_4912,N_4020,N_4430);
nor U4913 (N_4913,N_4147,N_4235);
nor U4914 (N_4914,N_4126,N_3923);
and U4915 (N_4915,N_3983,N_4463);
nor U4916 (N_4916,N_4445,N_4372);
nor U4917 (N_4917,N_4242,N_4063);
xnor U4918 (N_4918,N_4461,N_4425);
nand U4919 (N_4919,N_4159,N_3770);
and U4920 (N_4920,N_4095,N_4265);
and U4921 (N_4921,N_4353,N_4167);
nand U4922 (N_4922,N_3949,N_3885);
nor U4923 (N_4923,N_4258,N_3952);
xor U4924 (N_4924,N_3834,N_3948);
nand U4925 (N_4925,N_4026,N_4428);
and U4926 (N_4926,N_4378,N_3919);
nor U4927 (N_4927,N_4034,N_4401);
xnor U4928 (N_4928,N_3803,N_3759);
or U4929 (N_4929,N_3883,N_4071);
and U4930 (N_4930,N_3823,N_4004);
and U4931 (N_4931,N_4497,N_3780);
and U4932 (N_4932,N_3846,N_4354);
nand U4933 (N_4933,N_4106,N_4287);
or U4934 (N_4934,N_4129,N_4111);
or U4935 (N_4935,N_3887,N_4205);
and U4936 (N_4936,N_4457,N_4025);
xor U4937 (N_4937,N_4194,N_4489);
or U4938 (N_4938,N_4232,N_4375);
or U4939 (N_4939,N_4221,N_4025);
nor U4940 (N_4940,N_3870,N_3932);
or U4941 (N_4941,N_4378,N_4212);
nor U4942 (N_4942,N_4359,N_4252);
nor U4943 (N_4943,N_3821,N_3867);
xor U4944 (N_4944,N_3912,N_4255);
and U4945 (N_4945,N_4298,N_3856);
nand U4946 (N_4946,N_4096,N_3752);
or U4947 (N_4947,N_4408,N_4064);
or U4948 (N_4948,N_4091,N_4135);
nor U4949 (N_4949,N_4297,N_4241);
and U4950 (N_4950,N_4379,N_4118);
nor U4951 (N_4951,N_4398,N_3786);
nand U4952 (N_4952,N_4202,N_4059);
or U4953 (N_4953,N_4405,N_4175);
xnor U4954 (N_4954,N_4230,N_4415);
or U4955 (N_4955,N_4484,N_3907);
or U4956 (N_4956,N_4451,N_4252);
nand U4957 (N_4957,N_4000,N_4482);
xor U4958 (N_4958,N_4073,N_4148);
nand U4959 (N_4959,N_4070,N_3871);
xnor U4960 (N_4960,N_4309,N_4366);
xor U4961 (N_4961,N_4083,N_4298);
and U4962 (N_4962,N_4419,N_3878);
or U4963 (N_4963,N_3838,N_4331);
nand U4964 (N_4964,N_3876,N_4282);
nand U4965 (N_4965,N_4433,N_4475);
or U4966 (N_4966,N_3858,N_4315);
or U4967 (N_4967,N_4388,N_4468);
and U4968 (N_4968,N_4173,N_4276);
and U4969 (N_4969,N_3775,N_4494);
nor U4970 (N_4970,N_4025,N_3764);
nand U4971 (N_4971,N_4025,N_3958);
xor U4972 (N_4972,N_4270,N_4245);
nor U4973 (N_4973,N_3869,N_3757);
nand U4974 (N_4974,N_3855,N_4091);
xnor U4975 (N_4975,N_4049,N_4295);
and U4976 (N_4976,N_4033,N_4326);
and U4977 (N_4977,N_4077,N_3961);
or U4978 (N_4978,N_3867,N_3761);
nand U4979 (N_4979,N_4352,N_4296);
nor U4980 (N_4980,N_4107,N_4458);
or U4981 (N_4981,N_4132,N_4074);
nor U4982 (N_4982,N_4324,N_3872);
and U4983 (N_4983,N_3799,N_4474);
or U4984 (N_4984,N_4484,N_3753);
or U4985 (N_4985,N_4345,N_4178);
and U4986 (N_4986,N_4333,N_4398);
or U4987 (N_4987,N_4075,N_4315);
nor U4988 (N_4988,N_3835,N_4045);
and U4989 (N_4989,N_3957,N_4183);
nand U4990 (N_4990,N_4295,N_4055);
nor U4991 (N_4991,N_3835,N_4455);
and U4992 (N_4992,N_3796,N_3955);
nor U4993 (N_4993,N_4408,N_4146);
and U4994 (N_4994,N_4210,N_4132);
nor U4995 (N_4995,N_3872,N_4368);
nand U4996 (N_4996,N_3807,N_4359);
nor U4997 (N_4997,N_3989,N_4295);
nor U4998 (N_4998,N_3917,N_3930);
nor U4999 (N_4999,N_4420,N_4147);
nor U5000 (N_5000,N_3760,N_4268);
nand U5001 (N_5001,N_4341,N_4475);
and U5002 (N_5002,N_4133,N_3797);
nand U5003 (N_5003,N_4149,N_4278);
nand U5004 (N_5004,N_4477,N_4310);
nor U5005 (N_5005,N_4148,N_4210);
nand U5006 (N_5006,N_3858,N_4233);
nand U5007 (N_5007,N_4187,N_3897);
xor U5008 (N_5008,N_4043,N_4298);
nor U5009 (N_5009,N_4195,N_3942);
and U5010 (N_5010,N_4277,N_4322);
nor U5011 (N_5011,N_4057,N_3955);
nor U5012 (N_5012,N_3903,N_4257);
and U5013 (N_5013,N_4175,N_4304);
and U5014 (N_5014,N_4390,N_4452);
nor U5015 (N_5015,N_4029,N_4254);
or U5016 (N_5016,N_4146,N_3988);
nand U5017 (N_5017,N_3769,N_4357);
or U5018 (N_5018,N_4469,N_4280);
or U5019 (N_5019,N_4180,N_3766);
or U5020 (N_5020,N_4023,N_4380);
and U5021 (N_5021,N_4143,N_4105);
and U5022 (N_5022,N_4410,N_3823);
nand U5023 (N_5023,N_4432,N_4076);
nor U5024 (N_5024,N_3851,N_4201);
nor U5025 (N_5025,N_4326,N_4027);
nand U5026 (N_5026,N_3957,N_4076);
xnor U5027 (N_5027,N_3991,N_4043);
nor U5028 (N_5028,N_4428,N_4175);
nand U5029 (N_5029,N_4376,N_3931);
and U5030 (N_5030,N_4324,N_3986);
or U5031 (N_5031,N_4266,N_4450);
or U5032 (N_5032,N_4349,N_4027);
xor U5033 (N_5033,N_3750,N_4247);
or U5034 (N_5034,N_4171,N_3886);
xor U5035 (N_5035,N_3990,N_4298);
or U5036 (N_5036,N_4237,N_4246);
nand U5037 (N_5037,N_4447,N_3850);
and U5038 (N_5038,N_3966,N_4059);
xnor U5039 (N_5039,N_4333,N_4068);
or U5040 (N_5040,N_3896,N_4149);
or U5041 (N_5041,N_3978,N_4471);
or U5042 (N_5042,N_4207,N_4116);
nand U5043 (N_5043,N_3960,N_3862);
nand U5044 (N_5044,N_3906,N_4489);
or U5045 (N_5045,N_3809,N_3867);
and U5046 (N_5046,N_3861,N_4255);
nand U5047 (N_5047,N_3986,N_3991);
nor U5048 (N_5048,N_3974,N_4448);
or U5049 (N_5049,N_3949,N_4009);
nand U5050 (N_5050,N_4141,N_4494);
xor U5051 (N_5051,N_4226,N_4014);
xnor U5052 (N_5052,N_4136,N_4344);
and U5053 (N_5053,N_3758,N_4022);
nor U5054 (N_5054,N_4271,N_4456);
nand U5055 (N_5055,N_4295,N_3786);
or U5056 (N_5056,N_3887,N_4336);
nand U5057 (N_5057,N_4061,N_3934);
nand U5058 (N_5058,N_4012,N_4089);
xor U5059 (N_5059,N_4142,N_4460);
or U5060 (N_5060,N_4304,N_4159);
or U5061 (N_5061,N_4364,N_4315);
or U5062 (N_5062,N_4487,N_4231);
and U5063 (N_5063,N_3793,N_3967);
nor U5064 (N_5064,N_3806,N_4032);
nor U5065 (N_5065,N_4066,N_4393);
xnor U5066 (N_5066,N_4390,N_3938);
nand U5067 (N_5067,N_3772,N_3853);
or U5068 (N_5068,N_4147,N_4221);
nand U5069 (N_5069,N_3813,N_3987);
nand U5070 (N_5070,N_4411,N_3935);
and U5071 (N_5071,N_4366,N_4417);
or U5072 (N_5072,N_3904,N_4073);
nand U5073 (N_5073,N_4434,N_4420);
or U5074 (N_5074,N_4077,N_3920);
nand U5075 (N_5075,N_3870,N_4127);
or U5076 (N_5076,N_3870,N_4174);
nand U5077 (N_5077,N_4205,N_4007);
nor U5078 (N_5078,N_3934,N_4195);
and U5079 (N_5079,N_3939,N_4477);
nor U5080 (N_5080,N_4109,N_4284);
xor U5081 (N_5081,N_4225,N_4229);
xor U5082 (N_5082,N_3843,N_3966);
nor U5083 (N_5083,N_4423,N_4124);
nand U5084 (N_5084,N_4110,N_3759);
nor U5085 (N_5085,N_3995,N_3796);
nor U5086 (N_5086,N_4116,N_4239);
nor U5087 (N_5087,N_4294,N_4067);
nand U5088 (N_5088,N_4324,N_4419);
xnor U5089 (N_5089,N_4267,N_3870);
or U5090 (N_5090,N_4131,N_4006);
or U5091 (N_5091,N_3984,N_3847);
xnor U5092 (N_5092,N_3923,N_4371);
xnor U5093 (N_5093,N_4461,N_4295);
nor U5094 (N_5094,N_4496,N_4312);
nand U5095 (N_5095,N_3824,N_4265);
nand U5096 (N_5096,N_4191,N_3974);
nand U5097 (N_5097,N_4273,N_3840);
or U5098 (N_5098,N_4475,N_4376);
and U5099 (N_5099,N_4427,N_4308);
and U5100 (N_5100,N_4174,N_4150);
and U5101 (N_5101,N_4237,N_4404);
nor U5102 (N_5102,N_4361,N_4204);
nand U5103 (N_5103,N_4249,N_3765);
xor U5104 (N_5104,N_4152,N_4260);
and U5105 (N_5105,N_3892,N_4202);
nor U5106 (N_5106,N_4421,N_4196);
and U5107 (N_5107,N_4115,N_3942);
nor U5108 (N_5108,N_3940,N_4233);
nor U5109 (N_5109,N_3815,N_4384);
or U5110 (N_5110,N_4301,N_4002);
nand U5111 (N_5111,N_4223,N_3941);
or U5112 (N_5112,N_4174,N_3829);
and U5113 (N_5113,N_4067,N_3835);
or U5114 (N_5114,N_4475,N_3846);
nand U5115 (N_5115,N_4078,N_4085);
or U5116 (N_5116,N_4099,N_4212);
nor U5117 (N_5117,N_3828,N_4444);
and U5118 (N_5118,N_4033,N_4295);
nor U5119 (N_5119,N_3792,N_3785);
or U5120 (N_5120,N_4000,N_4209);
nor U5121 (N_5121,N_4073,N_3790);
or U5122 (N_5122,N_4159,N_3885);
nor U5123 (N_5123,N_4007,N_3985);
nand U5124 (N_5124,N_4304,N_4366);
nand U5125 (N_5125,N_3763,N_4447);
nor U5126 (N_5126,N_4432,N_4281);
and U5127 (N_5127,N_4008,N_4043);
nor U5128 (N_5128,N_4285,N_4484);
nor U5129 (N_5129,N_4409,N_3986);
and U5130 (N_5130,N_4145,N_4401);
and U5131 (N_5131,N_4248,N_3963);
nor U5132 (N_5132,N_3851,N_3906);
nor U5133 (N_5133,N_4046,N_3905);
nand U5134 (N_5134,N_3818,N_4169);
nand U5135 (N_5135,N_3820,N_4491);
or U5136 (N_5136,N_4158,N_3788);
and U5137 (N_5137,N_4116,N_4168);
and U5138 (N_5138,N_3885,N_4020);
nor U5139 (N_5139,N_4018,N_4422);
or U5140 (N_5140,N_4357,N_4449);
or U5141 (N_5141,N_4236,N_4151);
nor U5142 (N_5142,N_4473,N_4329);
and U5143 (N_5143,N_4032,N_4414);
and U5144 (N_5144,N_4259,N_3850);
or U5145 (N_5145,N_3873,N_4094);
nor U5146 (N_5146,N_4009,N_4305);
and U5147 (N_5147,N_4288,N_4304);
nor U5148 (N_5148,N_4034,N_4301);
and U5149 (N_5149,N_4172,N_4367);
or U5150 (N_5150,N_4193,N_4329);
or U5151 (N_5151,N_3846,N_4022);
and U5152 (N_5152,N_4085,N_4160);
or U5153 (N_5153,N_3764,N_4434);
nor U5154 (N_5154,N_4348,N_3781);
nor U5155 (N_5155,N_4011,N_4082);
and U5156 (N_5156,N_3755,N_4160);
xnor U5157 (N_5157,N_3884,N_4424);
nor U5158 (N_5158,N_3807,N_3828);
xor U5159 (N_5159,N_4158,N_3954);
xnor U5160 (N_5160,N_3754,N_4035);
nor U5161 (N_5161,N_4250,N_4474);
nand U5162 (N_5162,N_3990,N_4253);
and U5163 (N_5163,N_4349,N_4326);
xnor U5164 (N_5164,N_4274,N_4391);
or U5165 (N_5165,N_4014,N_4310);
nor U5166 (N_5166,N_3939,N_3782);
nor U5167 (N_5167,N_4315,N_4463);
nand U5168 (N_5168,N_4335,N_4068);
nor U5169 (N_5169,N_4101,N_4168);
xor U5170 (N_5170,N_4192,N_4206);
nand U5171 (N_5171,N_3960,N_4146);
nor U5172 (N_5172,N_4057,N_3892);
nor U5173 (N_5173,N_4077,N_3801);
nor U5174 (N_5174,N_4324,N_4364);
nor U5175 (N_5175,N_4319,N_4167);
or U5176 (N_5176,N_4165,N_3980);
xor U5177 (N_5177,N_3847,N_4254);
and U5178 (N_5178,N_3981,N_4416);
or U5179 (N_5179,N_3907,N_4012);
nor U5180 (N_5180,N_4245,N_3845);
and U5181 (N_5181,N_3979,N_3923);
nand U5182 (N_5182,N_3914,N_4112);
nor U5183 (N_5183,N_4027,N_3784);
nand U5184 (N_5184,N_3862,N_4259);
nor U5185 (N_5185,N_3906,N_4284);
nor U5186 (N_5186,N_3990,N_4182);
xnor U5187 (N_5187,N_4212,N_4002);
nand U5188 (N_5188,N_4270,N_4320);
nand U5189 (N_5189,N_4152,N_3942);
nand U5190 (N_5190,N_3989,N_4163);
nor U5191 (N_5191,N_4434,N_4157);
nand U5192 (N_5192,N_4161,N_4463);
and U5193 (N_5193,N_4108,N_4296);
or U5194 (N_5194,N_4343,N_4024);
nand U5195 (N_5195,N_3893,N_4285);
xnor U5196 (N_5196,N_3930,N_4090);
nand U5197 (N_5197,N_3976,N_4393);
and U5198 (N_5198,N_3884,N_4107);
nor U5199 (N_5199,N_3853,N_4008);
nand U5200 (N_5200,N_4232,N_3800);
or U5201 (N_5201,N_4186,N_3799);
or U5202 (N_5202,N_4154,N_4158);
or U5203 (N_5203,N_3933,N_4198);
nor U5204 (N_5204,N_4083,N_4166);
and U5205 (N_5205,N_3939,N_4327);
and U5206 (N_5206,N_4360,N_4067);
nand U5207 (N_5207,N_3782,N_4430);
nor U5208 (N_5208,N_3907,N_3755);
or U5209 (N_5209,N_4358,N_3843);
nand U5210 (N_5210,N_4283,N_4444);
nand U5211 (N_5211,N_4184,N_4326);
nor U5212 (N_5212,N_3825,N_4201);
and U5213 (N_5213,N_4081,N_4186);
or U5214 (N_5214,N_3893,N_3846);
and U5215 (N_5215,N_4282,N_4442);
nor U5216 (N_5216,N_4161,N_3941);
and U5217 (N_5217,N_4100,N_4326);
xor U5218 (N_5218,N_4338,N_4428);
or U5219 (N_5219,N_4063,N_4217);
nor U5220 (N_5220,N_4159,N_4418);
nor U5221 (N_5221,N_3763,N_4025);
xnor U5222 (N_5222,N_4161,N_3994);
and U5223 (N_5223,N_4465,N_4062);
nand U5224 (N_5224,N_4472,N_4244);
nand U5225 (N_5225,N_4053,N_4006);
nor U5226 (N_5226,N_4398,N_4052);
nor U5227 (N_5227,N_3913,N_3809);
or U5228 (N_5228,N_4100,N_4486);
and U5229 (N_5229,N_4069,N_4038);
or U5230 (N_5230,N_4007,N_4432);
and U5231 (N_5231,N_4021,N_4019);
or U5232 (N_5232,N_3822,N_3944);
and U5233 (N_5233,N_4466,N_4301);
or U5234 (N_5234,N_4335,N_4166);
nor U5235 (N_5235,N_3799,N_4101);
and U5236 (N_5236,N_4150,N_4033);
and U5237 (N_5237,N_4061,N_4450);
nand U5238 (N_5238,N_4078,N_4491);
and U5239 (N_5239,N_3768,N_4120);
or U5240 (N_5240,N_3908,N_4385);
nor U5241 (N_5241,N_4018,N_4250);
and U5242 (N_5242,N_4264,N_4012);
or U5243 (N_5243,N_4202,N_4398);
nor U5244 (N_5244,N_4367,N_3900);
and U5245 (N_5245,N_3845,N_4209);
and U5246 (N_5246,N_3986,N_3825);
xor U5247 (N_5247,N_4169,N_4204);
or U5248 (N_5248,N_3800,N_3853);
nand U5249 (N_5249,N_4106,N_3879);
nand U5250 (N_5250,N_5057,N_4971);
and U5251 (N_5251,N_4522,N_4761);
nor U5252 (N_5252,N_4632,N_4717);
or U5253 (N_5253,N_4669,N_4558);
nand U5254 (N_5254,N_4885,N_5220);
nand U5255 (N_5255,N_4663,N_5092);
or U5256 (N_5256,N_4561,N_4641);
or U5257 (N_5257,N_4538,N_4700);
nand U5258 (N_5258,N_4913,N_4598);
nor U5259 (N_5259,N_4869,N_4588);
xnor U5260 (N_5260,N_4575,N_5178);
nor U5261 (N_5261,N_4515,N_5051);
or U5262 (N_5262,N_4978,N_5099);
nand U5263 (N_5263,N_4672,N_4698);
nand U5264 (N_5264,N_4639,N_4676);
nor U5265 (N_5265,N_4610,N_4963);
and U5266 (N_5266,N_5015,N_5088);
or U5267 (N_5267,N_4535,N_4827);
and U5268 (N_5268,N_5127,N_4715);
or U5269 (N_5269,N_4880,N_4748);
xor U5270 (N_5270,N_5226,N_4998);
or U5271 (N_5271,N_4769,N_5045);
or U5272 (N_5272,N_5222,N_4525);
or U5273 (N_5273,N_5221,N_5105);
nand U5274 (N_5274,N_5113,N_4886);
nor U5275 (N_5275,N_5235,N_4648);
or U5276 (N_5276,N_4810,N_4758);
and U5277 (N_5277,N_4803,N_5173);
nand U5278 (N_5278,N_4794,N_4988);
nand U5279 (N_5279,N_4787,N_4604);
nor U5280 (N_5280,N_5144,N_5076);
and U5281 (N_5281,N_5019,N_5209);
xor U5282 (N_5282,N_5208,N_4824);
or U5283 (N_5283,N_4741,N_4569);
nand U5284 (N_5284,N_4937,N_5174);
nand U5285 (N_5285,N_5093,N_4829);
and U5286 (N_5286,N_4613,N_4601);
or U5287 (N_5287,N_4776,N_4782);
nor U5288 (N_5288,N_4714,N_4750);
and U5289 (N_5289,N_4557,N_4883);
nor U5290 (N_5290,N_4625,N_4730);
and U5291 (N_5291,N_4990,N_4865);
nor U5292 (N_5292,N_4950,N_4821);
and U5293 (N_5293,N_5110,N_4868);
or U5294 (N_5294,N_4529,N_5103);
and U5295 (N_5295,N_4766,N_5137);
xor U5296 (N_5296,N_4927,N_4890);
and U5297 (N_5297,N_4960,N_4893);
nor U5298 (N_5298,N_4790,N_4853);
nand U5299 (N_5299,N_4981,N_5072);
nor U5300 (N_5300,N_4837,N_5042);
nand U5301 (N_5301,N_4905,N_5095);
nand U5302 (N_5302,N_5081,N_4563);
xor U5303 (N_5303,N_4986,N_4595);
xor U5304 (N_5304,N_4550,N_4689);
nor U5305 (N_5305,N_5115,N_4933);
and U5306 (N_5306,N_4656,N_4936);
or U5307 (N_5307,N_4926,N_5244);
or U5308 (N_5308,N_4809,N_4819);
nand U5309 (N_5309,N_4932,N_5247);
nand U5310 (N_5310,N_4875,N_5071);
and U5311 (N_5311,N_5217,N_4553);
or U5312 (N_5312,N_5213,N_4593);
nor U5313 (N_5313,N_4954,N_4832);
or U5314 (N_5314,N_4582,N_4543);
xor U5315 (N_5315,N_5024,N_5248);
nand U5316 (N_5316,N_5100,N_4697);
nand U5317 (N_5317,N_4939,N_5000);
and U5318 (N_5318,N_4737,N_4762);
nand U5319 (N_5319,N_5167,N_4953);
and U5320 (N_5320,N_4531,N_5157);
nor U5321 (N_5321,N_4540,N_4802);
or U5322 (N_5322,N_4681,N_5234);
and U5323 (N_5323,N_4728,N_4644);
nor U5324 (N_5324,N_5188,N_4510);
nor U5325 (N_5325,N_4683,N_4620);
or U5326 (N_5326,N_4940,N_4823);
nand U5327 (N_5327,N_4907,N_5169);
nand U5328 (N_5328,N_4814,N_5021);
nor U5329 (N_5329,N_4660,N_4835);
nand U5330 (N_5330,N_4655,N_5034);
and U5331 (N_5331,N_4645,N_4712);
xor U5332 (N_5332,N_4735,N_5008);
xor U5333 (N_5333,N_4901,N_4921);
nand U5334 (N_5334,N_4898,N_4584);
nor U5335 (N_5335,N_4920,N_4984);
nor U5336 (N_5336,N_5053,N_4688);
nand U5337 (N_5337,N_4874,N_4753);
nor U5338 (N_5338,N_5128,N_5163);
nand U5339 (N_5339,N_4675,N_4581);
xor U5340 (N_5340,N_4616,N_5049);
xnor U5341 (N_5341,N_4851,N_4845);
or U5342 (N_5342,N_4935,N_5196);
or U5343 (N_5343,N_4554,N_4710);
nor U5344 (N_5344,N_5148,N_4979);
and U5345 (N_5345,N_4873,N_5218);
xor U5346 (N_5346,N_4603,N_4774);
and U5347 (N_5347,N_4820,N_4552);
nor U5348 (N_5348,N_4701,N_4590);
or U5349 (N_5349,N_4505,N_4864);
nand U5350 (N_5350,N_4638,N_5048);
nor U5351 (N_5351,N_4565,N_4560);
nor U5352 (N_5352,N_4574,N_4580);
or U5353 (N_5353,N_4773,N_4770);
nor U5354 (N_5354,N_4825,N_4928);
nand U5355 (N_5355,N_5140,N_4941);
and U5356 (N_5356,N_4679,N_4629);
or U5357 (N_5357,N_4972,N_4951);
nor U5358 (N_5358,N_4678,N_4804);
nor U5359 (N_5359,N_4997,N_5199);
nor U5360 (N_5360,N_5175,N_4577);
nand U5361 (N_5361,N_4504,N_4796);
nand U5362 (N_5362,N_4884,N_4947);
or U5363 (N_5363,N_4547,N_5031);
xnor U5364 (N_5364,N_4703,N_5176);
and U5365 (N_5365,N_4597,N_4686);
xor U5366 (N_5366,N_5044,N_4844);
nand U5367 (N_5367,N_4786,N_5134);
nor U5368 (N_5368,N_4843,N_4571);
nand U5369 (N_5369,N_4667,N_4812);
xor U5370 (N_5370,N_5006,N_4536);
and U5371 (N_5371,N_5060,N_4608);
and U5372 (N_5372,N_4549,N_4514);
or U5373 (N_5373,N_4719,N_4716);
and U5374 (N_5374,N_4799,N_4720);
and U5375 (N_5375,N_4793,N_5201);
and U5376 (N_5376,N_5181,N_4702);
or U5377 (N_5377,N_4973,N_4925);
or U5378 (N_5378,N_4520,N_5022);
and U5379 (N_5379,N_4602,N_4779);
and U5380 (N_5380,N_4573,N_5186);
nor U5381 (N_5381,N_4713,N_4975);
nand U5382 (N_5382,N_4881,N_4709);
or U5383 (N_5383,N_4706,N_4636);
nor U5384 (N_5384,N_4976,N_4503);
nand U5385 (N_5385,N_5180,N_4815);
and U5386 (N_5386,N_4768,N_5183);
and U5387 (N_5387,N_4548,N_4949);
nand U5388 (N_5388,N_5078,N_4858);
nand U5389 (N_5389,N_4662,N_4765);
nor U5390 (N_5390,N_5032,N_4665);
nor U5391 (N_5391,N_4943,N_4551);
nand U5392 (N_5392,N_5224,N_5237);
or U5393 (N_5393,N_4740,N_4980);
and U5394 (N_5394,N_4628,N_5233);
nor U5395 (N_5395,N_4867,N_4957);
nand U5396 (N_5396,N_4738,N_5239);
and U5397 (N_5397,N_5086,N_4879);
nand U5398 (N_5398,N_4922,N_4870);
nand U5399 (N_5399,N_5067,N_5164);
nand U5400 (N_5400,N_4784,N_4674);
xor U5401 (N_5401,N_5056,N_4813);
and U5402 (N_5402,N_4594,N_4859);
nor U5403 (N_5403,N_5055,N_5106);
or U5404 (N_5404,N_4760,N_4643);
nand U5405 (N_5405,N_5166,N_4772);
nand U5406 (N_5406,N_5131,N_4734);
nand U5407 (N_5407,N_4912,N_4904);
nand U5408 (N_5408,N_4727,N_4591);
and U5409 (N_5409,N_4704,N_4631);
or U5410 (N_5410,N_5107,N_4742);
and U5411 (N_5411,N_5133,N_5039);
and U5412 (N_5412,N_5108,N_5033);
nor U5413 (N_5413,N_4541,N_4956);
or U5414 (N_5414,N_4527,N_5138);
nor U5415 (N_5415,N_5159,N_5013);
nand U5416 (N_5416,N_5118,N_4725);
or U5417 (N_5417,N_4944,N_4755);
and U5418 (N_5418,N_4559,N_4839);
nand U5419 (N_5419,N_4897,N_5069);
nand U5420 (N_5420,N_4994,N_4671);
nor U5421 (N_5421,N_5195,N_4684);
nor U5422 (N_5422,N_5065,N_4707);
or U5423 (N_5423,N_4847,N_4838);
nor U5424 (N_5424,N_4860,N_5066);
nor U5425 (N_5425,N_5091,N_4854);
nor U5426 (N_5426,N_4614,N_5179);
xor U5427 (N_5427,N_4955,N_5172);
or U5428 (N_5428,N_5132,N_5171);
nand U5429 (N_5429,N_4919,N_4917);
nor U5430 (N_5430,N_5047,N_5227);
xnor U5431 (N_5431,N_4830,N_4649);
nand U5432 (N_5432,N_4544,N_5121);
nor U5433 (N_5433,N_4892,N_4948);
and U5434 (N_5434,N_4661,N_4857);
nor U5435 (N_5435,N_4789,N_5097);
nand U5436 (N_5436,N_5194,N_4846);
or U5437 (N_5437,N_4539,N_4657);
and U5438 (N_5438,N_4938,N_5136);
nand U5439 (N_5439,N_4617,N_4658);
nor U5440 (N_5440,N_4775,N_5184);
nand U5441 (N_5441,N_5187,N_4958);
nand U5442 (N_5442,N_5029,N_4506);
or U5443 (N_5443,N_4991,N_4512);
nor U5444 (N_5444,N_4586,N_4836);
nor U5445 (N_5445,N_5109,N_4583);
and U5446 (N_5446,N_4805,N_5154);
or U5447 (N_5447,N_4611,N_5145);
nor U5448 (N_5448,N_4524,N_5007);
nand U5449 (N_5449,N_5116,N_4771);
or U5450 (N_5450,N_5153,N_5002);
and U5451 (N_5451,N_4627,N_4866);
nand U5452 (N_5452,N_5059,N_4841);
and U5453 (N_5453,N_4599,N_4916);
or U5454 (N_5454,N_5054,N_4721);
xor U5455 (N_5455,N_4695,N_4791);
and U5456 (N_5456,N_4545,N_5241);
nor U5457 (N_5457,N_5214,N_4600);
and U5458 (N_5458,N_4877,N_4596);
nand U5459 (N_5459,N_4747,N_4767);
nand U5460 (N_5460,N_5098,N_4806);
nand U5461 (N_5461,N_4763,N_4511);
and U5462 (N_5462,N_5094,N_5219);
xnor U5463 (N_5463,N_4739,N_4816);
or U5464 (N_5464,N_5165,N_5011);
xor U5465 (N_5465,N_4895,N_4612);
nand U5466 (N_5466,N_4903,N_5185);
and U5467 (N_5467,N_4526,N_5156);
nand U5468 (N_5468,N_4607,N_5070);
or U5469 (N_5469,N_5182,N_4743);
and U5470 (N_5470,N_4637,N_4855);
or U5471 (N_5471,N_4652,N_4899);
and U5472 (N_5472,N_4621,N_5158);
nand U5473 (N_5473,N_5096,N_5212);
nand U5474 (N_5474,N_4871,N_5077);
nor U5475 (N_5475,N_4718,N_4894);
and U5476 (N_5476,N_5130,N_4729);
xnor U5477 (N_5477,N_5014,N_5223);
nor U5478 (N_5478,N_4754,N_5228);
nand U5479 (N_5479,N_5139,N_4723);
nor U5480 (N_5480,N_5177,N_5023);
and U5481 (N_5481,N_4831,N_5168);
nor U5482 (N_5482,N_4568,N_4646);
nor U5483 (N_5483,N_4930,N_5225);
nand U5484 (N_5484,N_4587,N_4759);
and U5485 (N_5485,N_4934,N_4882);
nand U5486 (N_5486,N_4680,N_5193);
nand U5487 (N_5487,N_5210,N_5117);
or U5488 (N_5488,N_4731,N_4502);
nand U5489 (N_5489,N_5090,N_4959);
and U5490 (N_5490,N_4924,N_4992);
or U5491 (N_5491,N_4798,N_5020);
nor U5492 (N_5492,N_4834,N_5012);
or U5493 (N_5493,N_4630,N_4746);
nor U5494 (N_5494,N_4682,N_4744);
and U5495 (N_5495,N_5245,N_4668);
or U5496 (N_5496,N_4908,N_4605);
nor U5497 (N_5497,N_4906,N_4696);
nand U5498 (N_5498,N_5030,N_5206);
and U5499 (N_5499,N_4902,N_5240);
nand U5500 (N_5500,N_5135,N_4778);
or U5501 (N_5501,N_5005,N_5238);
or U5502 (N_5502,N_5063,N_4777);
nand U5503 (N_5503,N_5232,N_4840);
or U5504 (N_5504,N_4626,N_4530);
nor U5505 (N_5505,N_4781,N_5120);
nand U5506 (N_5506,N_4732,N_4622);
and U5507 (N_5507,N_5203,N_5200);
and U5508 (N_5508,N_5236,N_4914);
xnor U5509 (N_5509,N_5204,N_4619);
and U5510 (N_5510,N_4592,N_5089);
or U5511 (N_5511,N_4647,N_4915);
or U5512 (N_5512,N_5150,N_4523);
and U5513 (N_5513,N_4785,N_4516);
xnor U5514 (N_5514,N_5162,N_5104);
xor U5515 (N_5515,N_4736,N_5202);
and U5516 (N_5516,N_4962,N_4685);
nand U5517 (N_5517,N_4896,N_5124);
and U5518 (N_5518,N_4751,N_4861);
nand U5519 (N_5519,N_5027,N_4811);
xor U5520 (N_5520,N_4817,N_4993);
or U5521 (N_5521,N_5038,N_4666);
or U5522 (N_5522,N_4711,N_5192);
xor U5523 (N_5523,N_5035,N_4966);
nand U5524 (N_5524,N_4964,N_4764);
nor U5525 (N_5525,N_4757,N_5125);
or U5526 (N_5526,N_4609,N_5040);
or U5527 (N_5527,N_5061,N_4989);
nor U5528 (N_5528,N_4642,N_4722);
or U5529 (N_5529,N_4889,N_4519);
or U5530 (N_5530,N_4677,N_5142);
nor U5531 (N_5531,N_4995,N_4640);
and U5532 (N_5532,N_4537,N_4850);
and U5533 (N_5533,N_5074,N_4826);
nor U5534 (N_5534,N_4726,N_4876);
or U5535 (N_5535,N_5025,N_4566);
nor U5536 (N_5536,N_5143,N_5149);
and U5537 (N_5537,N_4942,N_4961);
or U5538 (N_5538,N_4733,N_4507);
or U5539 (N_5539,N_5198,N_4659);
nand U5540 (N_5540,N_5191,N_4833);
or U5541 (N_5541,N_4570,N_4752);
and U5542 (N_5542,N_4635,N_5052);
or U5543 (N_5543,N_4694,N_4572);
or U5544 (N_5544,N_4518,N_5009);
nor U5545 (N_5545,N_5036,N_4862);
or U5546 (N_5546,N_4923,N_4900);
and U5547 (N_5547,N_5190,N_5147);
or U5548 (N_5548,N_5111,N_4521);
and U5549 (N_5549,N_4969,N_4567);
nand U5550 (N_5550,N_5058,N_5155);
nor U5551 (N_5551,N_4578,N_5126);
or U5552 (N_5552,N_4965,N_5119);
and U5553 (N_5553,N_4690,N_4780);
xnor U5554 (N_5554,N_4872,N_5216);
or U5555 (N_5555,N_4999,N_5112);
nand U5556 (N_5556,N_5085,N_5151);
or U5557 (N_5557,N_5001,N_5064);
or U5558 (N_5558,N_4888,N_4977);
or U5559 (N_5559,N_4807,N_4887);
or U5560 (N_5560,N_4756,N_4650);
nand U5561 (N_5561,N_4500,N_5211);
or U5562 (N_5562,N_5073,N_5189);
or U5563 (N_5563,N_5062,N_4606);
nand U5564 (N_5564,N_5084,N_4705);
xor U5565 (N_5565,N_5080,N_4970);
or U5566 (N_5566,N_4693,N_5004);
nor U5567 (N_5567,N_5050,N_5231);
and U5568 (N_5568,N_4983,N_5123);
nand U5569 (N_5569,N_4653,N_4967);
and U5570 (N_5570,N_5122,N_4501);
xor U5571 (N_5571,N_4533,N_4546);
nor U5572 (N_5572,N_4910,N_5215);
nand U5573 (N_5573,N_4795,N_5037);
and U5574 (N_5574,N_5230,N_4863);
or U5575 (N_5575,N_4664,N_4985);
nor U5576 (N_5576,N_4974,N_5017);
nor U5577 (N_5577,N_5026,N_4788);
or U5578 (N_5578,N_4542,N_5043);
xor U5579 (N_5579,N_4848,N_4708);
nand U5580 (N_5580,N_5003,N_4918);
or U5581 (N_5581,N_4534,N_4856);
or U5582 (N_5582,N_4909,N_5101);
nor U5583 (N_5583,N_5152,N_4987);
nor U5584 (N_5584,N_4946,N_5079);
or U5585 (N_5585,N_4528,N_4842);
nor U5586 (N_5586,N_4692,N_5205);
nand U5587 (N_5587,N_4509,N_4745);
nor U5588 (N_5588,N_4783,N_4911);
nor U5589 (N_5589,N_5129,N_4508);
and U5590 (N_5590,N_5197,N_4797);
nor U5591 (N_5591,N_4699,N_4564);
nand U5592 (N_5592,N_4800,N_5041);
nand U5593 (N_5593,N_4691,N_4852);
nor U5594 (N_5594,N_4687,N_4532);
nor U5595 (N_5595,N_4849,N_4555);
and U5596 (N_5596,N_4945,N_4952);
nand U5597 (N_5597,N_4562,N_5028);
or U5598 (N_5598,N_4968,N_4792);
nor U5599 (N_5599,N_4517,N_4615);
nand U5600 (N_5600,N_5242,N_4579);
nor U5601 (N_5601,N_4624,N_5018);
xor U5602 (N_5602,N_5146,N_4891);
nor U5603 (N_5603,N_4749,N_5161);
and U5604 (N_5604,N_4801,N_5082);
nand U5605 (N_5605,N_5016,N_5243);
nor U5606 (N_5606,N_5075,N_5114);
nor U5607 (N_5607,N_5046,N_5087);
and U5608 (N_5608,N_4982,N_4618);
or U5609 (N_5609,N_5249,N_4929);
nor U5610 (N_5610,N_4634,N_4654);
nor U5611 (N_5611,N_4996,N_4670);
nor U5612 (N_5612,N_5229,N_4822);
nand U5613 (N_5613,N_5102,N_5170);
nand U5614 (N_5614,N_4808,N_4724);
xnor U5615 (N_5615,N_5083,N_5207);
or U5616 (N_5616,N_4828,N_5068);
and U5617 (N_5617,N_4673,N_4513);
nor U5618 (N_5618,N_4576,N_4623);
xor U5619 (N_5619,N_4585,N_5246);
nor U5620 (N_5620,N_5010,N_4651);
nand U5621 (N_5621,N_5141,N_5160);
nand U5622 (N_5622,N_4589,N_4556);
nor U5623 (N_5623,N_4931,N_4818);
xnor U5624 (N_5624,N_4633,N_4878);
and U5625 (N_5625,N_4770,N_5097);
and U5626 (N_5626,N_4890,N_4836);
and U5627 (N_5627,N_4719,N_5230);
nand U5628 (N_5628,N_4943,N_4871);
nand U5629 (N_5629,N_5169,N_4508);
or U5630 (N_5630,N_4833,N_4609);
nand U5631 (N_5631,N_4974,N_4571);
xor U5632 (N_5632,N_5058,N_4786);
and U5633 (N_5633,N_4956,N_4965);
or U5634 (N_5634,N_4863,N_4787);
nor U5635 (N_5635,N_5192,N_4792);
nand U5636 (N_5636,N_4683,N_4817);
and U5637 (N_5637,N_5041,N_5237);
or U5638 (N_5638,N_4934,N_4621);
and U5639 (N_5639,N_4550,N_4544);
nand U5640 (N_5640,N_4583,N_4540);
and U5641 (N_5641,N_4920,N_5048);
nand U5642 (N_5642,N_4561,N_4816);
and U5643 (N_5643,N_5077,N_4625);
nand U5644 (N_5644,N_5006,N_4598);
and U5645 (N_5645,N_4952,N_5155);
or U5646 (N_5646,N_5055,N_4806);
nand U5647 (N_5647,N_4718,N_4616);
nor U5648 (N_5648,N_5022,N_5123);
and U5649 (N_5649,N_4994,N_5216);
nand U5650 (N_5650,N_4768,N_5210);
or U5651 (N_5651,N_4599,N_4504);
and U5652 (N_5652,N_4541,N_4769);
nor U5653 (N_5653,N_4581,N_4734);
or U5654 (N_5654,N_4697,N_5121);
and U5655 (N_5655,N_5233,N_4760);
or U5656 (N_5656,N_4514,N_4949);
and U5657 (N_5657,N_4687,N_4993);
nor U5658 (N_5658,N_4980,N_4671);
xor U5659 (N_5659,N_5074,N_4660);
nor U5660 (N_5660,N_4684,N_5080);
xor U5661 (N_5661,N_4543,N_5008);
and U5662 (N_5662,N_4613,N_4774);
xor U5663 (N_5663,N_4864,N_5112);
and U5664 (N_5664,N_4708,N_4574);
and U5665 (N_5665,N_4956,N_4775);
or U5666 (N_5666,N_4754,N_4722);
nor U5667 (N_5667,N_5034,N_4981);
or U5668 (N_5668,N_5162,N_5215);
or U5669 (N_5669,N_4965,N_4848);
nand U5670 (N_5670,N_4604,N_4925);
nor U5671 (N_5671,N_4896,N_4768);
nor U5672 (N_5672,N_4939,N_5190);
or U5673 (N_5673,N_4646,N_4791);
and U5674 (N_5674,N_5013,N_4721);
nor U5675 (N_5675,N_5180,N_4773);
nor U5676 (N_5676,N_5053,N_4858);
nor U5677 (N_5677,N_4618,N_4611);
nand U5678 (N_5678,N_4658,N_4542);
and U5679 (N_5679,N_4840,N_4912);
nor U5680 (N_5680,N_4756,N_4933);
nor U5681 (N_5681,N_4971,N_5034);
and U5682 (N_5682,N_5179,N_4808);
xnor U5683 (N_5683,N_5165,N_4585);
or U5684 (N_5684,N_4943,N_5149);
nor U5685 (N_5685,N_5036,N_4892);
nor U5686 (N_5686,N_4742,N_4538);
nor U5687 (N_5687,N_4502,N_5245);
and U5688 (N_5688,N_4836,N_4687);
or U5689 (N_5689,N_4898,N_4710);
nand U5690 (N_5690,N_4647,N_4521);
nor U5691 (N_5691,N_4564,N_4607);
nor U5692 (N_5692,N_4511,N_5098);
nand U5693 (N_5693,N_4918,N_4963);
nand U5694 (N_5694,N_4718,N_4855);
and U5695 (N_5695,N_4976,N_5165);
and U5696 (N_5696,N_5101,N_5190);
or U5697 (N_5697,N_5163,N_5082);
and U5698 (N_5698,N_4692,N_5140);
nand U5699 (N_5699,N_4704,N_5008);
nand U5700 (N_5700,N_4669,N_4589);
nand U5701 (N_5701,N_4630,N_4839);
xnor U5702 (N_5702,N_5043,N_4516);
nor U5703 (N_5703,N_4882,N_5129);
nand U5704 (N_5704,N_5245,N_4982);
and U5705 (N_5705,N_4989,N_5010);
and U5706 (N_5706,N_4594,N_4678);
nor U5707 (N_5707,N_4702,N_4927);
nand U5708 (N_5708,N_5035,N_5015);
nor U5709 (N_5709,N_4554,N_5018);
or U5710 (N_5710,N_4801,N_4899);
nor U5711 (N_5711,N_5173,N_4670);
and U5712 (N_5712,N_5025,N_4846);
and U5713 (N_5713,N_4761,N_5021);
or U5714 (N_5714,N_5123,N_4689);
or U5715 (N_5715,N_4541,N_5183);
and U5716 (N_5716,N_4960,N_4711);
xor U5717 (N_5717,N_4875,N_5243);
nor U5718 (N_5718,N_5005,N_4786);
nand U5719 (N_5719,N_5158,N_4925);
or U5720 (N_5720,N_4764,N_5244);
and U5721 (N_5721,N_4970,N_4793);
and U5722 (N_5722,N_5090,N_5116);
and U5723 (N_5723,N_4739,N_4806);
or U5724 (N_5724,N_4639,N_4622);
nand U5725 (N_5725,N_5091,N_4704);
nor U5726 (N_5726,N_5214,N_4948);
nand U5727 (N_5727,N_4584,N_4871);
nand U5728 (N_5728,N_5062,N_4670);
nor U5729 (N_5729,N_4729,N_5207);
and U5730 (N_5730,N_4931,N_5184);
and U5731 (N_5731,N_4798,N_4528);
and U5732 (N_5732,N_4516,N_5193);
nand U5733 (N_5733,N_5241,N_5210);
xnor U5734 (N_5734,N_4816,N_4737);
nor U5735 (N_5735,N_4946,N_4540);
nor U5736 (N_5736,N_4675,N_4818);
or U5737 (N_5737,N_4757,N_5063);
nand U5738 (N_5738,N_4969,N_4513);
nor U5739 (N_5739,N_5171,N_5161);
nor U5740 (N_5740,N_5222,N_4784);
nand U5741 (N_5741,N_4943,N_5010);
nor U5742 (N_5742,N_4637,N_4837);
or U5743 (N_5743,N_4619,N_5105);
nand U5744 (N_5744,N_4718,N_5160);
nand U5745 (N_5745,N_4766,N_4891);
or U5746 (N_5746,N_4955,N_4736);
nand U5747 (N_5747,N_4969,N_4957);
and U5748 (N_5748,N_4612,N_4992);
or U5749 (N_5749,N_4711,N_5207);
nand U5750 (N_5750,N_5222,N_5212);
or U5751 (N_5751,N_4542,N_4673);
nand U5752 (N_5752,N_5220,N_5049);
xnor U5753 (N_5753,N_4523,N_4735);
nand U5754 (N_5754,N_5020,N_4997);
xnor U5755 (N_5755,N_4958,N_5068);
and U5756 (N_5756,N_4835,N_4552);
nand U5757 (N_5757,N_4824,N_4536);
or U5758 (N_5758,N_4736,N_4537);
nand U5759 (N_5759,N_5049,N_4644);
xnor U5760 (N_5760,N_4923,N_4835);
nor U5761 (N_5761,N_4822,N_4563);
nand U5762 (N_5762,N_4624,N_4598);
nor U5763 (N_5763,N_4981,N_4608);
or U5764 (N_5764,N_5099,N_5184);
or U5765 (N_5765,N_5011,N_5218);
xor U5766 (N_5766,N_4576,N_5136);
or U5767 (N_5767,N_4996,N_4560);
or U5768 (N_5768,N_4533,N_4627);
xnor U5769 (N_5769,N_4992,N_5067);
nand U5770 (N_5770,N_4730,N_4627);
nor U5771 (N_5771,N_4716,N_4760);
nand U5772 (N_5772,N_5018,N_4948);
nor U5773 (N_5773,N_4823,N_5022);
nand U5774 (N_5774,N_4966,N_5062);
nor U5775 (N_5775,N_4911,N_5116);
nand U5776 (N_5776,N_4898,N_4843);
xnor U5777 (N_5777,N_5120,N_4690);
nand U5778 (N_5778,N_4605,N_4892);
or U5779 (N_5779,N_4908,N_5192);
nor U5780 (N_5780,N_4543,N_4576);
nor U5781 (N_5781,N_4624,N_4636);
nor U5782 (N_5782,N_5079,N_4563);
nand U5783 (N_5783,N_5189,N_4851);
xor U5784 (N_5784,N_5150,N_4832);
nor U5785 (N_5785,N_5203,N_4891);
or U5786 (N_5786,N_4523,N_4739);
or U5787 (N_5787,N_4955,N_5059);
and U5788 (N_5788,N_4536,N_5228);
nor U5789 (N_5789,N_4723,N_4696);
nor U5790 (N_5790,N_4578,N_4616);
or U5791 (N_5791,N_4939,N_5009);
or U5792 (N_5792,N_4786,N_5236);
nand U5793 (N_5793,N_4979,N_4655);
or U5794 (N_5794,N_4614,N_4598);
nor U5795 (N_5795,N_5063,N_4742);
xnor U5796 (N_5796,N_4878,N_4539);
nand U5797 (N_5797,N_4536,N_5029);
or U5798 (N_5798,N_4837,N_5179);
xor U5799 (N_5799,N_5095,N_4725);
nor U5800 (N_5800,N_5146,N_4571);
nand U5801 (N_5801,N_4822,N_5195);
xnor U5802 (N_5802,N_5059,N_5043);
or U5803 (N_5803,N_4767,N_4803);
and U5804 (N_5804,N_4571,N_4904);
nand U5805 (N_5805,N_4940,N_5175);
nand U5806 (N_5806,N_5206,N_4595);
and U5807 (N_5807,N_5207,N_4618);
nor U5808 (N_5808,N_5227,N_4800);
nand U5809 (N_5809,N_5154,N_5142);
or U5810 (N_5810,N_4918,N_4581);
or U5811 (N_5811,N_4804,N_4886);
nand U5812 (N_5812,N_4865,N_4722);
xor U5813 (N_5813,N_4583,N_4707);
nand U5814 (N_5814,N_4910,N_5240);
nor U5815 (N_5815,N_4980,N_5122);
nor U5816 (N_5816,N_4789,N_5053);
nor U5817 (N_5817,N_5081,N_5233);
nand U5818 (N_5818,N_4640,N_4922);
or U5819 (N_5819,N_4644,N_5036);
nor U5820 (N_5820,N_5076,N_4683);
nor U5821 (N_5821,N_4659,N_4503);
nor U5822 (N_5822,N_5025,N_5240);
and U5823 (N_5823,N_4616,N_4795);
nand U5824 (N_5824,N_4747,N_4971);
and U5825 (N_5825,N_4501,N_4776);
and U5826 (N_5826,N_4588,N_5171);
nand U5827 (N_5827,N_4858,N_4760);
or U5828 (N_5828,N_4886,N_4688);
or U5829 (N_5829,N_5045,N_4522);
xor U5830 (N_5830,N_4999,N_4748);
nor U5831 (N_5831,N_4789,N_4855);
and U5832 (N_5832,N_4679,N_5011);
nand U5833 (N_5833,N_4961,N_5244);
and U5834 (N_5834,N_4912,N_4817);
or U5835 (N_5835,N_4794,N_4505);
nand U5836 (N_5836,N_4686,N_4738);
xor U5837 (N_5837,N_4718,N_4770);
nand U5838 (N_5838,N_4501,N_5001);
xnor U5839 (N_5839,N_4962,N_4708);
nand U5840 (N_5840,N_4718,N_4658);
nand U5841 (N_5841,N_4755,N_5158);
nand U5842 (N_5842,N_4785,N_4589);
nand U5843 (N_5843,N_5060,N_4657);
and U5844 (N_5844,N_5121,N_4554);
xnor U5845 (N_5845,N_5139,N_5244);
nand U5846 (N_5846,N_4706,N_4593);
and U5847 (N_5847,N_4576,N_4925);
nor U5848 (N_5848,N_4879,N_4671);
nor U5849 (N_5849,N_4644,N_4899);
nor U5850 (N_5850,N_5186,N_5153);
nor U5851 (N_5851,N_5007,N_4984);
or U5852 (N_5852,N_4902,N_4881);
and U5853 (N_5853,N_4773,N_4656);
nor U5854 (N_5854,N_4650,N_4943);
or U5855 (N_5855,N_5083,N_4730);
or U5856 (N_5856,N_4820,N_4706);
nor U5857 (N_5857,N_5197,N_4506);
nand U5858 (N_5858,N_4569,N_5150);
or U5859 (N_5859,N_5202,N_4533);
or U5860 (N_5860,N_4615,N_4541);
nor U5861 (N_5861,N_4741,N_4619);
nand U5862 (N_5862,N_4925,N_4572);
or U5863 (N_5863,N_4799,N_5149);
nand U5864 (N_5864,N_4710,N_4915);
or U5865 (N_5865,N_4701,N_5206);
nand U5866 (N_5866,N_4588,N_4712);
nand U5867 (N_5867,N_4987,N_4821);
nand U5868 (N_5868,N_4984,N_4643);
or U5869 (N_5869,N_4561,N_5019);
nor U5870 (N_5870,N_4829,N_4922);
or U5871 (N_5871,N_4629,N_5217);
nand U5872 (N_5872,N_4526,N_5249);
nand U5873 (N_5873,N_4907,N_4941);
nand U5874 (N_5874,N_5068,N_5205);
and U5875 (N_5875,N_5068,N_4883);
or U5876 (N_5876,N_4846,N_4800);
or U5877 (N_5877,N_5077,N_4960);
or U5878 (N_5878,N_4920,N_4505);
nand U5879 (N_5879,N_5128,N_4517);
nand U5880 (N_5880,N_4928,N_4954);
xnor U5881 (N_5881,N_4573,N_5006);
nor U5882 (N_5882,N_4945,N_5005);
and U5883 (N_5883,N_4814,N_5063);
and U5884 (N_5884,N_5245,N_5196);
nand U5885 (N_5885,N_4604,N_4608);
nand U5886 (N_5886,N_4819,N_5016);
nand U5887 (N_5887,N_4921,N_4947);
and U5888 (N_5888,N_4693,N_4879);
or U5889 (N_5889,N_5146,N_5130);
nand U5890 (N_5890,N_4933,N_5114);
or U5891 (N_5891,N_5128,N_5021);
or U5892 (N_5892,N_5115,N_4701);
or U5893 (N_5893,N_4995,N_4702);
nor U5894 (N_5894,N_4628,N_4714);
or U5895 (N_5895,N_4522,N_4847);
and U5896 (N_5896,N_4999,N_4773);
or U5897 (N_5897,N_4821,N_4735);
or U5898 (N_5898,N_4819,N_4985);
nor U5899 (N_5899,N_5148,N_5113);
nor U5900 (N_5900,N_5103,N_5131);
nor U5901 (N_5901,N_5210,N_4788);
and U5902 (N_5902,N_4681,N_4931);
and U5903 (N_5903,N_5075,N_4689);
nand U5904 (N_5904,N_4659,N_4819);
nor U5905 (N_5905,N_4734,N_4531);
or U5906 (N_5906,N_4654,N_4823);
nand U5907 (N_5907,N_4812,N_5112);
nand U5908 (N_5908,N_5238,N_4826);
nand U5909 (N_5909,N_5185,N_4630);
nor U5910 (N_5910,N_4659,N_4998);
xor U5911 (N_5911,N_4968,N_4847);
xnor U5912 (N_5912,N_4673,N_5231);
nand U5913 (N_5913,N_5048,N_4833);
nand U5914 (N_5914,N_4540,N_4858);
and U5915 (N_5915,N_5125,N_5140);
and U5916 (N_5916,N_4670,N_4568);
and U5917 (N_5917,N_4686,N_5219);
nand U5918 (N_5918,N_4593,N_5102);
or U5919 (N_5919,N_4630,N_5028);
nor U5920 (N_5920,N_4578,N_5090);
or U5921 (N_5921,N_5023,N_5067);
nand U5922 (N_5922,N_4673,N_4921);
nand U5923 (N_5923,N_4866,N_4774);
nor U5924 (N_5924,N_4646,N_5246);
xnor U5925 (N_5925,N_5023,N_4784);
nor U5926 (N_5926,N_4637,N_4500);
and U5927 (N_5927,N_5135,N_4503);
nor U5928 (N_5928,N_4865,N_5174);
and U5929 (N_5929,N_4896,N_4529);
or U5930 (N_5930,N_4738,N_4855);
nand U5931 (N_5931,N_4747,N_5143);
xnor U5932 (N_5932,N_5162,N_5066);
and U5933 (N_5933,N_4953,N_5155);
or U5934 (N_5934,N_5174,N_5057);
and U5935 (N_5935,N_4650,N_5062);
nor U5936 (N_5936,N_5183,N_4639);
nor U5937 (N_5937,N_4748,N_4513);
or U5938 (N_5938,N_5103,N_4546);
nor U5939 (N_5939,N_4601,N_5089);
and U5940 (N_5940,N_5121,N_4560);
nand U5941 (N_5941,N_4872,N_4566);
nor U5942 (N_5942,N_4723,N_4994);
or U5943 (N_5943,N_4971,N_5074);
or U5944 (N_5944,N_5099,N_5068);
nor U5945 (N_5945,N_4790,N_5154);
or U5946 (N_5946,N_4714,N_4823);
and U5947 (N_5947,N_4869,N_4548);
nand U5948 (N_5948,N_4963,N_5011);
nor U5949 (N_5949,N_4765,N_5096);
nand U5950 (N_5950,N_5029,N_5010);
nor U5951 (N_5951,N_5056,N_5203);
or U5952 (N_5952,N_4600,N_5079);
nor U5953 (N_5953,N_5188,N_4545);
or U5954 (N_5954,N_4533,N_4935);
or U5955 (N_5955,N_5100,N_4705);
nand U5956 (N_5956,N_5150,N_4565);
nor U5957 (N_5957,N_4982,N_4964);
nand U5958 (N_5958,N_4700,N_4871);
nand U5959 (N_5959,N_5064,N_4627);
xor U5960 (N_5960,N_4511,N_4547);
xor U5961 (N_5961,N_5115,N_4703);
and U5962 (N_5962,N_5149,N_4848);
and U5963 (N_5963,N_4667,N_5057);
and U5964 (N_5964,N_4909,N_5008);
or U5965 (N_5965,N_5146,N_5227);
nand U5966 (N_5966,N_4828,N_5235);
nor U5967 (N_5967,N_4925,N_4599);
or U5968 (N_5968,N_4896,N_4948);
or U5969 (N_5969,N_4504,N_4952);
or U5970 (N_5970,N_4829,N_4979);
or U5971 (N_5971,N_4605,N_4581);
xnor U5972 (N_5972,N_5240,N_4916);
or U5973 (N_5973,N_4933,N_5071);
nor U5974 (N_5974,N_4654,N_5091);
nand U5975 (N_5975,N_4841,N_5175);
nor U5976 (N_5976,N_5009,N_5093);
and U5977 (N_5977,N_5238,N_4633);
or U5978 (N_5978,N_4897,N_4946);
xor U5979 (N_5979,N_4583,N_5217);
and U5980 (N_5980,N_4682,N_5160);
or U5981 (N_5981,N_4623,N_5088);
and U5982 (N_5982,N_5080,N_5161);
and U5983 (N_5983,N_4938,N_5000);
nor U5984 (N_5984,N_4819,N_5185);
and U5985 (N_5985,N_5099,N_4836);
and U5986 (N_5986,N_4772,N_4784);
or U5987 (N_5987,N_4690,N_4884);
or U5988 (N_5988,N_4815,N_4607);
nor U5989 (N_5989,N_4947,N_4539);
xor U5990 (N_5990,N_4915,N_4658);
and U5991 (N_5991,N_4735,N_5146);
nand U5992 (N_5992,N_4957,N_5068);
and U5993 (N_5993,N_5190,N_4593);
nand U5994 (N_5994,N_4668,N_5059);
nand U5995 (N_5995,N_5104,N_4539);
or U5996 (N_5996,N_5009,N_4728);
or U5997 (N_5997,N_4805,N_4831);
nand U5998 (N_5998,N_5029,N_4614);
and U5999 (N_5999,N_4908,N_4817);
or U6000 (N_6000,N_5676,N_5269);
and U6001 (N_6001,N_5838,N_5482);
nand U6002 (N_6002,N_5680,N_5588);
xnor U6003 (N_6003,N_5740,N_5871);
and U6004 (N_6004,N_5793,N_5656);
and U6005 (N_6005,N_5526,N_5732);
nor U6006 (N_6006,N_5825,N_5869);
nand U6007 (N_6007,N_5916,N_5924);
or U6008 (N_6008,N_5909,N_5747);
nand U6009 (N_6009,N_5559,N_5964);
xor U6010 (N_6010,N_5847,N_5873);
and U6011 (N_6011,N_5726,N_5690);
xnor U6012 (N_6012,N_5837,N_5563);
nor U6013 (N_6013,N_5552,N_5452);
and U6014 (N_6014,N_5432,N_5763);
nand U6015 (N_6015,N_5928,N_5442);
and U6016 (N_6016,N_5765,N_5301);
nor U6017 (N_6017,N_5570,N_5906);
or U6018 (N_6018,N_5773,N_5807);
nor U6019 (N_6019,N_5817,N_5384);
and U6020 (N_6020,N_5761,N_5927);
or U6021 (N_6021,N_5772,N_5706);
or U6022 (N_6022,N_5589,N_5451);
and U6023 (N_6023,N_5988,N_5984);
and U6024 (N_6024,N_5974,N_5897);
or U6025 (N_6025,N_5294,N_5677);
nor U6026 (N_6026,N_5686,N_5290);
nand U6027 (N_6027,N_5867,N_5416);
nand U6028 (N_6028,N_5769,N_5542);
nor U6029 (N_6029,N_5839,N_5537);
nand U6030 (N_6030,N_5692,N_5320);
nor U6031 (N_6031,N_5657,N_5612);
nand U6032 (N_6032,N_5377,N_5637);
and U6033 (N_6033,N_5860,N_5957);
xnor U6034 (N_6034,N_5539,N_5633);
or U6035 (N_6035,N_5971,N_5786);
nand U6036 (N_6036,N_5393,N_5700);
nand U6037 (N_6037,N_5823,N_5851);
nor U6038 (N_6038,N_5444,N_5864);
or U6039 (N_6039,N_5836,N_5749);
and U6040 (N_6040,N_5310,N_5647);
and U6041 (N_6041,N_5306,N_5579);
and U6042 (N_6042,N_5565,N_5337);
and U6043 (N_6043,N_5913,N_5423);
nor U6044 (N_6044,N_5911,N_5620);
nand U6045 (N_6045,N_5986,N_5936);
nand U6046 (N_6046,N_5636,N_5833);
or U6047 (N_6047,N_5580,N_5991);
and U6048 (N_6048,N_5492,N_5983);
and U6049 (N_6049,N_5696,N_5488);
or U6050 (N_6050,N_5336,N_5783);
or U6051 (N_6051,N_5642,N_5972);
nand U6052 (N_6052,N_5907,N_5877);
nor U6053 (N_6053,N_5711,N_5495);
or U6054 (N_6054,N_5595,N_5281);
nor U6055 (N_6055,N_5976,N_5937);
and U6056 (N_6056,N_5594,N_5311);
nand U6057 (N_6057,N_5961,N_5456);
nor U6058 (N_6058,N_5593,N_5804);
nor U6059 (N_6059,N_5938,N_5862);
or U6060 (N_6060,N_5904,N_5868);
and U6061 (N_6061,N_5486,N_5926);
xnor U6062 (N_6062,N_5949,N_5496);
or U6063 (N_6063,N_5331,N_5756);
and U6064 (N_6064,N_5943,N_5303);
nor U6065 (N_6065,N_5410,N_5323);
or U6066 (N_6066,N_5666,N_5601);
nand U6067 (N_6067,N_5374,N_5951);
nand U6068 (N_6068,N_5380,N_5292);
or U6069 (N_6069,N_5822,N_5446);
nand U6070 (N_6070,N_5501,N_5569);
or U6071 (N_6071,N_5679,N_5250);
nor U6072 (N_6072,N_5577,N_5762);
and U6073 (N_6073,N_5436,N_5866);
and U6074 (N_6074,N_5853,N_5895);
nand U6075 (N_6075,N_5258,N_5812);
nor U6076 (N_6076,N_5330,N_5611);
nand U6077 (N_6077,N_5638,N_5314);
nor U6078 (N_6078,N_5992,N_5634);
nor U6079 (N_6079,N_5865,N_5363);
and U6080 (N_6080,N_5473,N_5405);
nor U6081 (N_6081,N_5267,N_5344);
and U6082 (N_6082,N_5465,N_5532);
nand U6083 (N_6083,N_5785,N_5555);
nand U6084 (N_6084,N_5575,N_5746);
or U6085 (N_6085,N_5418,N_5391);
nand U6086 (N_6086,N_5720,N_5343);
nand U6087 (N_6087,N_5508,N_5764);
nand U6088 (N_6088,N_5963,N_5420);
and U6089 (N_6089,N_5382,N_5341);
or U6090 (N_6090,N_5848,N_5828);
or U6091 (N_6091,N_5962,N_5479);
nand U6092 (N_6092,N_5484,N_5313);
xor U6093 (N_6093,N_5574,N_5730);
nor U6094 (N_6094,N_5470,N_5273);
and U6095 (N_6095,N_5725,N_5535);
nor U6096 (N_6096,N_5684,N_5941);
and U6097 (N_6097,N_5315,N_5286);
nor U6098 (N_6098,N_5489,N_5852);
nor U6099 (N_6099,N_5381,N_5931);
and U6100 (N_6100,N_5297,N_5878);
or U6101 (N_6101,N_5985,N_5613);
and U6102 (N_6102,N_5805,N_5285);
nand U6103 (N_6103,N_5854,N_5795);
and U6104 (N_6104,N_5345,N_5792);
nand U6105 (N_6105,N_5824,N_5364);
and U6106 (N_6106,N_5434,N_5815);
or U6107 (N_6107,N_5843,N_5276);
nand U6108 (N_6108,N_5467,N_5806);
and U6109 (N_6109,N_5304,N_5850);
or U6110 (N_6110,N_5955,N_5392);
xor U6111 (N_6111,N_5333,N_5813);
or U6112 (N_6112,N_5958,N_5386);
or U6113 (N_6113,N_5270,N_5447);
nand U6114 (N_6114,N_5426,N_5998);
and U6115 (N_6115,N_5438,N_5491);
or U6116 (N_6116,N_5284,N_5332);
or U6117 (N_6117,N_5758,N_5462);
nand U6118 (N_6118,N_5359,N_5959);
nand U6119 (N_6119,N_5500,N_5728);
and U6120 (N_6120,N_5329,N_5973);
nand U6121 (N_6121,N_5790,N_5340);
nand U6122 (N_6122,N_5404,N_5655);
nand U6123 (N_6123,N_5631,N_5841);
or U6124 (N_6124,N_5327,N_5530);
nor U6125 (N_6125,N_5994,N_5480);
and U6126 (N_6126,N_5752,N_5626);
xor U6127 (N_6127,N_5401,N_5885);
nor U6128 (N_6128,N_5437,N_5770);
and U6129 (N_6129,N_5794,N_5693);
or U6130 (N_6130,N_5921,N_5261);
nor U6131 (N_6131,N_5845,N_5378);
xor U6132 (N_6132,N_5997,N_5506);
nand U6133 (N_6133,N_5471,N_5798);
and U6134 (N_6134,N_5365,N_5578);
or U6135 (N_6135,N_5271,N_5754);
or U6136 (N_6136,N_5424,N_5520);
nand U6137 (N_6137,N_5902,N_5682);
xor U6138 (N_6138,N_5767,N_5400);
nor U6139 (N_6139,N_5893,N_5670);
nand U6140 (N_6140,N_5969,N_5298);
and U6141 (N_6141,N_5940,N_5945);
nand U6142 (N_6142,N_5373,N_5737);
and U6143 (N_6143,N_5981,N_5891);
or U6144 (N_6144,N_5801,N_5347);
and U6145 (N_6145,N_5741,N_5675);
and U6146 (N_6146,N_5319,N_5641);
and U6147 (N_6147,N_5624,N_5414);
and U6148 (N_6148,N_5557,N_5523);
nand U6149 (N_6149,N_5738,N_5629);
and U6150 (N_6150,N_5605,N_5430);
and U6151 (N_6151,N_5650,N_5497);
or U6152 (N_6152,N_5603,N_5614);
and U6153 (N_6153,N_5733,N_5731);
and U6154 (N_6154,N_5457,N_5870);
nand U6155 (N_6155,N_5576,N_5996);
or U6156 (N_6156,N_5439,N_5989);
or U6157 (N_6157,N_5879,N_5361);
or U6158 (N_6158,N_5810,N_5954);
and U6159 (N_6159,N_5698,N_5324);
or U6160 (N_6160,N_5787,N_5277);
and U6161 (N_6161,N_5543,N_5394);
and U6162 (N_6162,N_5397,N_5896);
nor U6163 (N_6163,N_5979,N_5709);
or U6164 (N_6164,N_5428,N_5517);
nor U6165 (N_6165,N_5702,N_5745);
or U6166 (N_6166,N_5604,N_5504);
or U6167 (N_6167,N_5915,N_5369);
nand U6168 (N_6168,N_5708,N_5503);
or U6169 (N_6169,N_5651,N_5948);
or U6170 (N_6170,N_5774,N_5275);
nor U6171 (N_6171,N_5445,N_5606);
and U6172 (N_6172,N_5929,N_5661);
and U6173 (N_6173,N_5944,N_5376);
and U6174 (N_6174,N_5930,N_5912);
nor U6175 (N_6175,N_5265,N_5280);
and U6176 (N_6176,N_5779,N_5540);
nor U6177 (N_6177,N_5339,N_5309);
nand U6178 (N_6178,N_5257,N_5383);
and U6179 (N_6179,N_5547,N_5960);
and U6180 (N_6180,N_5408,N_5987);
nand U6181 (N_6181,N_5548,N_5710);
and U6182 (N_6182,N_5412,N_5308);
and U6183 (N_6183,N_5584,N_5375);
nand U6184 (N_6184,N_5553,N_5556);
or U6185 (N_6185,N_5662,N_5326);
nand U6186 (N_6186,N_5742,N_5653);
nor U6187 (N_6187,N_5466,N_5932);
nor U6188 (N_6188,N_5784,N_5875);
nand U6189 (N_6189,N_5759,N_5478);
or U6190 (N_6190,N_5721,N_5302);
nor U6191 (N_6191,N_5640,N_5328);
or U6192 (N_6192,N_5385,N_5622);
nor U6193 (N_6193,N_5490,N_5671);
nor U6194 (N_6194,N_5321,N_5417);
nand U6195 (N_6195,N_5667,N_5818);
and U6196 (N_6196,N_5287,N_5597);
and U6197 (N_6197,N_5715,N_5609);
or U6198 (N_6198,N_5512,N_5826);
and U6199 (N_6199,N_5534,N_5820);
and U6200 (N_6200,N_5399,N_5630);
nand U6201 (N_6201,N_5712,N_5840);
nor U6202 (N_6202,N_5372,N_5704);
and U6203 (N_6203,N_5914,N_5727);
nand U6204 (N_6204,N_5652,N_5305);
or U6205 (N_6205,N_5683,N_5886);
nor U6206 (N_6206,N_5789,N_5846);
nand U6207 (N_6207,N_5735,N_5856);
or U6208 (N_6208,N_5882,N_5751);
nand U6209 (N_6209,N_5724,N_5977);
nor U6210 (N_6210,N_5799,N_5529);
or U6211 (N_6211,N_5797,N_5664);
nor U6212 (N_6212,N_5599,N_5816);
or U6213 (N_6213,N_5694,N_5645);
nand U6214 (N_6214,N_5362,N_5487);
or U6215 (N_6215,N_5901,N_5583);
nor U6216 (N_6216,N_5649,N_5254);
xnor U6217 (N_6217,N_5561,N_5691);
and U6218 (N_6218,N_5757,N_5398);
and U6219 (N_6219,N_5858,N_5884);
and U6220 (N_6220,N_5502,N_5295);
or U6221 (N_6221,N_5755,N_5481);
nand U6222 (N_6222,N_5252,N_5390);
nor U6223 (N_6223,N_5722,N_5367);
nand U6224 (N_6224,N_5872,N_5768);
nor U6225 (N_6225,N_5293,N_5448);
nor U6226 (N_6226,N_5278,N_5525);
and U6227 (N_6227,N_5995,N_5519);
nand U6228 (N_6228,N_5409,N_5716);
nor U6229 (N_6229,N_5834,N_5253);
and U6230 (N_6230,N_5952,N_5659);
and U6231 (N_6231,N_5739,N_5685);
and U6232 (N_6232,N_5585,N_5499);
nand U6233 (N_6233,N_5978,N_5616);
xor U6234 (N_6234,N_5288,N_5464);
or U6235 (N_6235,N_5353,N_5748);
xnor U6236 (N_6236,N_5586,N_5596);
or U6237 (N_6237,N_5965,N_5348);
and U6238 (N_6238,N_5821,N_5990);
nand U6239 (N_6239,N_5493,N_5279);
nor U6240 (N_6240,N_5617,N_5509);
nor U6241 (N_6241,N_5510,N_5956);
nor U6242 (N_6242,N_5317,N_5713);
xnor U6243 (N_6243,N_5300,N_5842);
or U6244 (N_6244,N_5673,N_5717);
nor U6245 (N_6245,N_5402,N_5411);
nor U6246 (N_6246,N_5366,N_5459);
nand U6247 (N_6247,N_5908,N_5600);
and U6248 (N_6248,N_5474,N_5890);
and U6249 (N_6249,N_5791,N_5455);
or U6250 (N_6250,N_5346,N_5777);
or U6251 (N_6251,N_5796,N_5678);
xnor U6252 (N_6252,N_5263,N_5554);
nand U6253 (N_6253,N_5460,N_5883);
nor U6254 (N_6254,N_5966,N_5358);
or U6255 (N_6255,N_5920,N_5541);
nand U6256 (N_6256,N_5528,N_5546);
and U6257 (N_6257,N_5619,N_5514);
nor U6258 (N_6258,N_5602,N_5674);
nand U6259 (N_6259,N_5814,N_5819);
nand U6260 (N_6260,N_5950,N_5356);
nand U6261 (N_6261,N_5421,N_5888);
or U6262 (N_6262,N_5407,N_5780);
nor U6263 (N_6263,N_5703,N_5933);
or U6264 (N_6264,N_5567,N_5635);
nor U6265 (N_6265,N_5355,N_5894);
and U6266 (N_6266,N_5803,N_5396);
and U6267 (N_6267,N_5458,N_5830);
or U6268 (N_6268,N_5469,N_5935);
and U6269 (N_6269,N_5663,N_5590);
nand U6270 (N_6270,N_5750,N_5370);
or U6271 (N_6271,N_5766,N_5831);
and U6272 (N_6272,N_5349,N_5531);
nor U6273 (N_6273,N_5802,N_5660);
nand U6274 (N_6274,N_5776,N_5403);
and U6275 (N_6275,N_5413,N_5934);
or U6276 (N_6276,N_5621,N_5415);
or U6277 (N_6277,N_5628,N_5863);
nand U6278 (N_6278,N_5454,N_5753);
xor U6279 (N_6279,N_5527,N_5639);
nand U6280 (N_6280,N_5431,N_5476);
nor U6281 (N_6281,N_5551,N_5665);
xor U6282 (N_6282,N_5654,N_5607);
nor U6283 (N_6283,N_5681,N_5699);
nand U6284 (N_6284,N_5433,N_5475);
nor U6285 (N_6285,N_5775,N_5544);
or U6286 (N_6286,N_5472,N_5387);
and U6287 (N_6287,N_5334,N_5573);
or U6288 (N_6288,N_5485,N_5760);
xnor U6289 (N_6289,N_5827,N_5581);
nor U6290 (N_6290,N_5461,N_5782);
or U6291 (N_6291,N_5498,N_5395);
and U6292 (N_6292,N_5264,N_5351);
or U6293 (N_6293,N_5549,N_5947);
nor U6294 (N_6294,N_5919,N_5880);
xor U6295 (N_6295,N_5259,N_5942);
and U6296 (N_6296,N_5272,N_5771);
nor U6297 (N_6297,N_5322,N_5887);
or U6298 (N_6298,N_5483,N_5524);
xnor U6299 (N_6299,N_5505,N_5422);
xor U6300 (N_6300,N_5388,N_5435);
nand U6301 (N_6301,N_5855,N_5354);
nand U6302 (N_6302,N_5350,N_5892);
nor U6303 (N_6303,N_5811,N_5729);
nor U6304 (N_6304,N_5618,N_5695);
nand U6305 (N_6305,N_5256,N_5658);
nor U6306 (N_6306,N_5953,N_5389);
nand U6307 (N_6307,N_5564,N_5874);
nand U6308 (N_6308,N_5342,N_5371);
or U6309 (N_6309,N_5296,N_5861);
nand U6310 (N_6310,N_5781,N_5463);
nand U6311 (N_6311,N_5379,N_5571);
nor U6312 (N_6312,N_5644,N_5357);
and U6313 (N_6313,N_5829,N_5849);
and U6314 (N_6314,N_5723,N_5939);
nor U6315 (N_6315,N_5274,N_5283);
xor U6316 (N_6316,N_5560,N_5844);
nand U6317 (N_6317,N_5477,N_5859);
nor U6318 (N_6318,N_5903,N_5516);
nor U6319 (N_6319,N_5610,N_5587);
nor U6320 (N_6320,N_5425,N_5568);
xnor U6321 (N_6321,N_5689,N_5923);
or U6322 (N_6322,N_5632,N_5441);
nand U6323 (N_6323,N_5307,N_5687);
and U6324 (N_6324,N_5889,N_5905);
and U6325 (N_6325,N_5352,N_5453);
nor U6326 (N_6326,N_5910,N_5545);
nor U6327 (N_6327,N_5688,N_5970);
nor U6328 (N_6328,N_5566,N_5719);
and U6329 (N_6329,N_5513,N_5967);
xnor U6330 (N_6330,N_5917,N_5325);
nor U6331 (N_6331,N_5623,N_5443);
and U6332 (N_6332,N_5668,N_5980);
or U6333 (N_6333,N_5898,N_5922);
or U6334 (N_6334,N_5260,N_5450);
nor U6335 (N_6335,N_5582,N_5521);
or U6336 (N_6336,N_5625,N_5515);
or U6337 (N_6337,N_5946,N_5507);
and U6338 (N_6338,N_5511,N_5429);
xor U6339 (N_6339,N_5266,N_5736);
and U6340 (N_6340,N_5881,N_5262);
and U6341 (N_6341,N_5312,N_5809);
nor U6342 (N_6342,N_5550,N_5646);
or U6343 (N_6343,N_5982,N_5299);
xnor U6344 (N_6344,N_5925,N_5419);
nor U6345 (N_6345,N_5360,N_5562);
and U6346 (N_6346,N_5558,N_5999);
nand U6347 (N_6347,N_5835,N_5316);
nand U6348 (N_6348,N_5572,N_5268);
and U6349 (N_6349,N_5368,N_5788);
nor U6350 (N_6350,N_5282,N_5899);
xnor U6351 (N_6351,N_5251,N_5672);
nand U6352 (N_6352,N_5800,N_5406);
or U6353 (N_6353,N_5522,N_5744);
nand U6354 (N_6354,N_5718,N_5714);
nor U6355 (N_6355,N_5591,N_5968);
and U6356 (N_6356,N_5643,N_5707);
and U6357 (N_6357,N_5518,N_5427);
or U6358 (N_6358,N_5291,N_5975);
xnor U6359 (N_6359,N_5832,N_5705);
nor U6360 (N_6360,N_5449,N_5648);
nor U6361 (N_6361,N_5627,N_5808);
xnor U6362 (N_6362,N_5615,N_5743);
nand U6363 (N_6363,N_5536,N_5669);
or U6364 (N_6364,N_5533,N_5335);
and U6365 (N_6365,N_5494,N_5598);
xnor U6366 (N_6366,N_5338,N_5440);
and U6367 (N_6367,N_5697,N_5918);
or U6368 (N_6368,N_5255,N_5592);
nand U6369 (N_6369,N_5468,N_5734);
nor U6370 (N_6370,N_5538,N_5857);
xor U6371 (N_6371,N_5778,N_5993);
nor U6372 (N_6372,N_5318,N_5876);
nor U6373 (N_6373,N_5701,N_5900);
nor U6374 (N_6374,N_5289,N_5608);
nor U6375 (N_6375,N_5254,N_5341);
nand U6376 (N_6376,N_5719,N_5965);
nand U6377 (N_6377,N_5863,N_5681);
or U6378 (N_6378,N_5473,N_5671);
xnor U6379 (N_6379,N_5675,N_5281);
nor U6380 (N_6380,N_5981,N_5965);
nand U6381 (N_6381,N_5266,N_5293);
nand U6382 (N_6382,N_5613,N_5374);
or U6383 (N_6383,N_5731,N_5830);
or U6384 (N_6384,N_5727,N_5411);
nand U6385 (N_6385,N_5715,N_5991);
or U6386 (N_6386,N_5817,N_5720);
or U6387 (N_6387,N_5429,N_5730);
and U6388 (N_6388,N_5658,N_5697);
nand U6389 (N_6389,N_5310,N_5571);
and U6390 (N_6390,N_5443,N_5972);
nor U6391 (N_6391,N_5614,N_5824);
nor U6392 (N_6392,N_5885,N_5465);
and U6393 (N_6393,N_5872,N_5612);
or U6394 (N_6394,N_5426,N_5936);
or U6395 (N_6395,N_5439,N_5374);
or U6396 (N_6396,N_5295,N_5834);
or U6397 (N_6397,N_5760,N_5767);
nand U6398 (N_6398,N_5291,N_5926);
xor U6399 (N_6399,N_5421,N_5727);
xnor U6400 (N_6400,N_5522,N_5439);
and U6401 (N_6401,N_5656,N_5706);
xor U6402 (N_6402,N_5292,N_5984);
or U6403 (N_6403,N_5432,N_5858);
and U6404 (N_6404,N_5573,N_5765);
xor U6405 (N_6405,N_5943,N_5553);
nor U6406 (N_6406,N_5991,N_5552);
nand U6407 (N_6407,N_5953,N_5739);
and U6408 (N_6408,N_5667,N_5947);
or U6409 (N_6409,N_5280,N_5311);
and U6410 (N_6410,N_5986,N_5533);
or U6411 (N_6411,N_5830,N_5996);
nor U6412 (N_6412,N_5999,N_5626);
nor U6413 (N_6413,N_5915,N_5679);
nor U6414 (N_6414,N_5507,N_5303);
and U6415 (N_6415,N_5573,N_5436);
nor U6416 (N_6416,N_5922,N_5340);
and U6417 (N_6417,N_5607,N_5595);
nor U6418 (N_6418,N_5650,N_5968);
nand U6419 (N_6419,N_5376,N_5965);
and U6420 (N_6420,N_5564,N_5301);
and U6421 (N_6421,N_5281,N_5926);
or U6422 (N_6422,N_5777,N_5592);
nand U6423 (N_6423,N_5493,N_5988);
nand U6424 (N_6424,N_5410,N_5561);
nor U6425 (N_6425,N_5874,N_5882);
nor U6426 (N_6426,N_5524,N_5823);
and U6427 (N_6427,N_5744,N_5597);
nand U6428 (N_6428,N_5278,N_5460);
nor U6429 (N_6429,N_5567,N_5506);
xor U6430 (N_6430,N_5914,N_5510);
xnor U6431 (N_6431,N_5754,N_5317);
nor U6432 (N_6432,N_5312,N_5732);
or U6433 (N_6433,N_5756,N_5530);
nand U6434 (N_6434,N_5836,N_5408);
or U6435 (N_6435,N_5751,N_5417);
or U6436 (N_6436,N_5819,N_5383);
xor U6437 (N_6437,N_5967,N_5990);
nor U6438 (N_6438,N_5581,N_5442);
nand U6439 (N_6439,N_5903,N_5838);
xnor U6440 (N_6440,N_5755,N_5855);
nor U6441 (N_6441,N_5992,N_5443);
or U6442 (N_6442,N_5641,N_5510);
nand U6443 (N_6443,N_5959,N_5256);
xor U6444 (N_6444,N_5593,N_5705);
nand U6445 (N_6445,N_5358,N_5521);
and U6446 (N_6446,N_5585,N_5709);
nor U6447 (N_6447,N_5835,N_5909);
nand U6448 (N_6448,N_5945,N_5459);
nand U6449 (N_6449,N_5571,N_5536);
and U6450 (N_6450,N_5701,N_5883);
and U6451 (N_6451,N_5961,N_5646);
nand U6452 (N_6452,N_5434,N_5795);
xnor U6453 (N_6453,N_5536,N_5711);
nand U6454 (N_6454,N_5809,N_5678);
nand U6455 (N_6455,N_5615,N_5846);
and U6456 (N_6456,N_5507,N_5769);
xor U6457 (N_6457,N_5421,N_5447);
nand U6458 (N_6458,N_5933,N_5300);
nand U6459 (N_6459,N_5628,N_5487);
nor U6460 (N_6460,N_5290,N_5927);
nand U6461 (N_6461,N_5318,N_5347);
and U6462 (N_6462,N_5472,N_5654);
nand U6463 (N_6463,N_5902,N_5366);
nand U6464 (N_6464,N_5284,N_5499);
and U6465 (N_6465,N_5877,N_5333);
or U6466 (N_6466,N_5476,N_5673);
or U6467 (N_6467,N_5755,N_5621);
nor U6468 (N_6468,N_5521,N_5400);
nor U6469 (N_6469,N_5780,N_5319);
nand U6470 (N_6470,N_5395,N_5952);
nor U6471 (N_6471,N_5895,N_5435);
and U6472 (N_6472,N_5657,N_5480);
and U6473 (N_6473,N_5253,N_5451);
or U6474 (N_6474,N_5572,N_5520);
nor U6475 (N_6475,N_5255,N_5369);
or U6476 (N_6476,N_5845,N_5463);
xnor U6477 (N_6477,N_5423,N_5997);
or U6478 (N_6478,N_5880,N_5347);
and U6479 (N_6479,N_5330,N_5735);
or U6480 (N_6480,N_5785,N_5442);
or U6481 (N_6481,N_5558,N_5753);
or U6482 (N_6482,N_5803,N_5872);
nor U6483 (N_6483,N_5610,N_5913);
or U6484 (N_6484,N_5806,N_5775);
and U6485 (N_6485,N_5553,N_5357);
nor U6486 (N_6486,N_5277,N_5568);
nor U6487 (N_6487,N_5740,N_5483);
or U6488 (N_6488,N_5900,N_5620);
and U6489 (N_6489,N_5814,N_5560);
or U6490 (N_6490,N_5591,N_5746);
nor U6491 (N_6491,N_5918,N_5968);
or U6492 (N_6492,N_5689,N_5618);
and U6493 (N_6493,N_5966,N_5732);
nor U6494 (N_6494,N_5358,N_5332);
nand U6495 (N_6495,N_5858,N_5385);
and U6496 (N_6496,N_5386,N_5448);
nand U6497 (N_6497,N_5454,N_5519);
and U6498 (N_6498,N_5620,N_5765);
or U6499 (N_6499,N_5912,N_5390);
nor U6500 (N_6500,N_5355,N_5676);
nand U6501 (N_6501,N_5316,N_5751);
and U6502 (N_6502,N_5862,N_5500);
nor U6503 (N_6503,N_5612,N_5873);
or U6504 (N_6504,N_5933,N_5672);
nand U6505 (N_6505,N_5741,N_5548);
nor U6506 (N_6506,N_5605,N_5575);
xor U6507 (N_6507,N_5813,N_5654);
and U6508 (N_6508,N_5811,N_5935);
nand U6509 (N_6509,N_5398,N_5460);
or U6510 (N_6510,N_5783,N_5908);
or U6511 (N_6511,N_5329,N_5470);
and U6512 (N_6512,N_5653,N_5254);
nand U6513 (N_6513,N_5954,N_5532);
and U6514 (N_6514,N_5917,N_5314);
and U6515 (N_6515,N_5698,N_5761);
nor U6516 (N_6516,N_5293,N_5354);
nand U6517 (N_6517,N_5286,N_5629);
nand U6518 (N_6518,N_5720,N_5257);
or U6519 (N_6519,N_5581,N_5460);
nor U6520 (N_6520,N_5359,N_5679);
nand U6521 (N_6521,N_5393,N_5661);
xnor U6522 (N_6522,N_5717,N_5499);
nand U6523 (N_6523,N_5332,N_5849);
xnor U6524 (N_6524,N_5800,N_5323);
nor U6525 (N_6525,N_5688,N_5943);
and U6526 (N_6526,N_5372,N_5342);
nand U6527 (N_6527,N_5515,N_5385);
or U6528 (N_6528,N_5907,N_5687);
nand U6529 (N_6529,N_5438,N_5475);
or U6530 (N_6530,N_5711,N_5621);
nor U6531 (N_6531,N_5710,N_5330);
and U6532 (N_6532,N_5713,N_5890);
or U6533 (N_6533,N_5825,N_5914);
and U6534 (N_6534,N_5913,N_5727);
nor U6535 (N_6535,N_5315,N_5570);
nor U6536 (N_6536,N_5857,N_5893);
nand U6537 (N_6537,N_5965,N_5461);
and U6538 (N_6538,N_5428,N_5731);
or U6539 (N_6539,N_5322,N_5898);
and U6540 (N_6540,N_5665,N_5583);
or U6541 (N_6541,N_5570,N_5734);
xor U6542 (N_6542,N_5788,N_5782);
and U6543 (N_6543,N_5454,N_5382);
and U6544 (N_6544,N_5310,N_5579);
nand U6545 (N_6545,N_5433,N_5771);
nand U6546 (N_6546,N_5674,N_5941);
and U6547 (N_6547,N_5922,N_5943);
nor U6548 (N_6548,N_5643,N_5285);
nor U6549 (N_6549,N_5577,N_5319);
nand U6550 (N_6550,N_5440,N_5768);
and U6551 (N_6551,N_5310,N_5654);
or U6552 (N_6552,N_5862,N_5978);
or U6553 (N_6553,N_5828,N_5965);
nor U6554 (N_6554,N_5703,N_5806);
nand U6555 (N_6555,N_5787,N_5636);
or U6556 (N_6556,N_5642,N_5377);
nand U6557 (N_6557,N_5658,N_5608);
or U6558 (N_6558,N_5660,N_5671);
nand U6559 (N_6559,N_5963,N_5419);
and U6560 (N_6560,N_5361,N_5917);
nor U6561 (N_6561,N_5539,N_5670);
nor U6562 (N_6562,N_5358,N_5705);
and U6563 (N_6563,N_5565,N_5559);
nand U6564 (N_6564,N_5415,N_5427);
xnor U6565 (N_6565,N_5913,N_5713);
nand U6566 (N_6566,N_5378,N_5784);
nor U6567 (N_6567,N_5822,N_5667);
and U6568 (N_6568,N_5840,N_5666);
nand U6569 (N_6569,N_5329,N_5942);
or U6570 (N_6570,N_5469,N_5539);
nand U6571 (N_6571,N_5319,N_5666);
nor U6572 (N_6572,N_5949,N_5900);
or U6573 (N_6573,N_5651,N_5454);
nor U6574 (N_6574,N_5927,N_5977);
nor U6575 (N_6575,N_5559,N_5444);
and U6576 (N_6576,N_5391,N_5771);
nand U6577 (N_6577,N_5485,N_5822);
and U6578 (N_6578,N_5597,N_5465);
or U6579 (N_6579,N_5562,N_5564);
or U6580 (N_6580,N_5940,N_5859);
and U6581 (N_6581,N_5533,N_5363);
and U6582 (N_6582,N_5378,N_5367);
nor U6583 (N_6583,N_5990,N_5343);
and U6584 (N_6584,N_5510,N_5871);
and U6585 (N_6585,N_5326,N_5657);
nor U6586 (N_6586,N_5393,N_5629);
nor U6587 (N_6587,N_5388,N_5587);
or U6588 (N_6588,N_5264,N_5723);
and U6589 (N_6589,N_5501,N_5545);
nand U6590 (N_6590,N_5369,N_5693);
and U6591 (N_6591,N_5736,N_5800);
and U6592 (N_6592,N_5712,N_5281);
and U6593 (N_6593,N_5400,N_5621);
and U6594 (N_6594,N_5690,N_5587);
or U6595 (N_6595,N_5499,N_5371);
or U6596 (N_6596,N_5885,N_5805);
nor U6597 (N_6597,N_5608,N_5640);
and U6598 (N_6598,N_5844,N_5556);
and U6599 (N_6599,N_5347,N_5963);
nand U6600 (N_6600,N_5423,N_5445);
and U6601 (N_6601,N_5735,N_5987);
nand U6602 (N_6602,N_5814,N_5888);
nor U6603 (N_6603,N_5423,N_5564);
and U6604 (N_6604,N_5256,N_5807);
xor U6605 (N_6605,N_5558,N_5505);
nor U6606 (N_6606,N_5645,N_5396);
nand U6607 (N_6607,N_5490,N_5929);
nor U6608 (N_6608,N_5901,N_5651);
and U6609 (N_6609,N_5331,N_5503);
nor U6610 (N_6610,N_5280,N_5498);
nand U6611 (N_6611,N_5441,N_5933);
xnor U6612 (N_6612,N_5350,N_5391);
or U6613 (N_6613,N_5689,N_5702);
nor U6614 (N_6614,N_5612,N_5685);
or U6615 (N_6615,N_5657,N_5857);
or U6616 (N_6616,N_5363,N_5709);
and U6617 (N_6617,N_5552,N_5671);
or U6618 (N_6618,N_5917,N_5449);
nor U6619 (N_6619,N_5345,N_5462);
nand U6620 (N_6620,N_5880,N_5257);
nor U6621 (N_6621,N_5610,N_5346);
nand U6622 (N_6622,N_5647,N_5689);
and U6623 (N_6623,N_5981,N_5493);
nor U6624 (N_6624,N_5349,N_5264);
and U6625 (N_6625,N_5411,N_5601);
and U6626 (N_6626,N_5883,N_5293);
and U6627 (N_6627,N_5323,N_5862);
nand U6628 (N_6628,N_5575,N_5437);
nand U6629 (N_6629,N_5610,N_5926);
nor U6630 (N_6630,N_5923,N_5264);
or U6631 (N_6631,N_5525,N_5962);
and U6632 (N_6632,N_5733,N_5765);
nand U6633 (N_6633,N_5990,N_5290);
and U6634 (N_6634,N_5437,N_5440);
nand U6635 (N_6635,N_5287,N_5299);
nor U6636 (N_6636,N_5925,N_5322);
and U6637 (N_6637,N_5837,N_5592);
nor U6638 (N_6638,N_5690,N_5317);
nand U6639 (N_6639,N_5652,N_5992);
nand U6640 (N_6640,N_5586,N_5957);
and U6641 (N_6641,N_5592,N_5441);
nor U6642 (N_6642,N_5733,N_5522);
nand U6643 (N_6643,N_5768,N_5711);
nand U6644 (N_6644,N_5880,N_5826);
and U6645 (N_6645,N_5520,N_5558);
xor U6646 (N_6646,N_5462,N_5750);
nor U6647 (N_6647,N_5727,N_5564);
nand U6648 (N_6648,N_5729,N_5456);
and U6649 (N_6649,N_5401,N_5886);
nor U6650 (N_6650,N_5943,N_5378);
nor U6651 (N_6651,N_5550,N_5863);
and U6652 (N_6652,N_5915,N_5758);
nand U6653 (N_6653,N_5302,N_5720);
nand U6654 (N_6654,N_5285,N_5555);
nor U6655 (N_6655,N_5637,N_5299);
nand U6656 (N_6656,N_5861,N_5689);
or U6657 (N_6657,N_5354,N_5689);
nand U6658 (N_6658,N_5509,N_5364);
nor U6659 (N_6659,N_5559,N_5711);
nand U6660 (N_6660,N_5343,N_5759);
nand U6661 (N_6661,N_5514,N_5476);
or U6662 (N_6662,N_5259,N_5505);
and U6663 (N_6663,N_5413,N_5270);
nand U6664 (N_6664,N_5739,N_5603);
xor U6665 (N_6665,N_5508,N_5596);
and U6666 (N_6666,N_5434,N_5587);
xnor U6667 (N_6667,N_5588,N_5730);
and U6668 (N_6668,N_5255,N_5821);
or U6669 (N_6669,N_5443,N_5622);
and U6670 (N_6670,N_5865,N_5783);
xor U6671 (N_6671,N_5923,N_5403);
and U6672 (N_6672,N_5883,N_5485);
xor U6673 (N_6673,N_5446,N_5992);
and U6674 (N_6674,N_5479,N_5427);
or U6675 (N_6675,N_5907,N_5853);
or U6676 (N_6676,N_5413,N_5935);
nand U6677 (N_6677,N_5628,N_5873);
xnor U6678 (N_6678,N_5904,N_5622);
nor U6679 (N_6679,N_5513,N_5400);
or U6680 (N_6680,N_5258,N_5262);
and U6681 (N_6681,N_5715,N_5505);
nand U6682 (N_6682,N_5390,N_5486);
or U6683 (N_6683,N_5393,N_5327);
or U6684 (N_6684,N_5883,N_5591);
and U6685 (N_6685,N_5544,N_5971);
nor U6686 (N_6686,N_5467,N_5699);
or U6687 (N_6687,N_5986,N_5383);
nor U6688 (N_6688,N_5724,N_5531);
and U6689 (N_6689,N_5837,N_5580);
or U6690 (N_6690,N_5817,N_5568);
nor U6691 (N_6691,N_5629,N_5911);
or U6692 (N_6692,N_5436,N_5704);
and U6693 (N_6693,N_5999,N_5986);
nor U6694 (N_6694,N_5761,N_5639);
nor U6695 (N_6695,N_5732,N_5980);
xnor U6696 (N_6696,N_5650,N_5591);
and U6697 (N_6697,N_5894,N_5943);
nor U6698 (N_6698,N_5615,N_5574);
nor U6699 (N_6699,N_5535,N_5660);
and U6700 (N_6700,N_5740,N_5922);
nand U6701 (N_6701,N_5895,N_5627);
nor U6702 (N_6702,N_5727,N_5472);
nor U6703 (N_6703,N_5707,N_5798);
xor U6704 (N_6704,N_5260,N_5451);
nand U6705 (N_6705,N_5833,N_5840);
and U6706 (N_6706,N_5547,N_5711);
xnor U6707 (N_6707,N_5300,N_5869);
nand U6708 (N_6708,N_5914,N_5648);
or U6709 (N_6709,N_5274,N_5659);
nand U6710 (N_6710,N_5916,N_5732);
or U6711 (N_6711,N_5428,N_5943);
nand U6712 (N_6712,N_5736,N_5400);
nand U6713 (N_6713,N_5629,N_5470);
or U6714 (N_6714,N_5380,N_5675);
or U6715 (N_6715,N_5600,N_5441);
or U6716 (N_6716,N_5376,N_5728);
and U6717 (N_6717,N_5317,N_5703);
or U6718 (N_6718,N_5465,N_5602);
and U6719 (N_6719,N_5431,N_5652);
nand U6720 (N_6720,N_5751,N_5987);
nand U6721 (N_6721,N_5333,N_5888);
nand U6722 (N_6722,N_5875,N_5596);
or U6723 (N_6723,N_5727,N_5600);
nand U6724 (N_6724,N_5297,N_5414);
nor U6725 (N_6725,N_5913,N_5936);
nand U6726 (N_6726,N_5498,N_5791);
nand U6727 (N_6727,N_5660,N_5350);
nor U6728 (N_6728,N_5876,N_5940);
or U6729 (N_6729,N_5851,N_5414);
nor U6730 (N_6730,N_5975,N_5311);
nand U6731 (N_6731,N_5847,N_5970);
nand U6732 (N_6732,N_5543,N_5825);
xnor U6733 (N_6733,N_5794,N_5810);
nand U6734 (N_6734,N_5653,N_5783);
or U6735 (N_6735,N_5889,N_5608);
nor U6736 (N_6736,N_5390,N_5382);
nor U6737 (N_6737,N_5730,N_5871);
xor U6738 (N_6738,N_5342,N_5990);
and U6739 (N_6739,N_5954,N_5331);
nand U6740 (N_6740,N_5602,N_5489);
and U6741 (N_6741,N_5534,N_5619);
and U6742 (N_6742,N_5515,N_5495);
nor U6743 (N_6743,N_5643,N_5350);
nand U6744 (N_6744,N_5846,N_5362);
xor U6745 (N_6745,N_5903,N_5555);
and U6746 (N_6746,N_5600,N_5400);
nand U6747 (N_6747,N_5485,N_5817);
nand U6748 (N_6748,N_5686,N_5306);
and U6749 (N_6749,N_5788,N_5522);
or U6750 (N_6750,N_6379,N_6620);
and U6751 (N_6751,N_6673,N_6577);
nor U6752 (N_6752,N_6713,N_6259);
and U6753 (N_6753,N_6035,N_6427);
nand U6754 (N_6754,N_6685,N_6342);
or U6755 (N_6755,N_6677,N_6429);
nor U6756 (N_6756,N_6221,N_6012);
nor U6757 (N_6757,N_6595,N_6572);
nor U6758 (N_6758,N_6301,N_6591);
nand U6759 (N_6759,N_6013,N_6528);
nand U6760 (N_6760,N_6005,N_6455);
nor U6761 (N_6761,N_6740,N_6331);
nor U6762 (N_6762,N_6149,N_6442);
and U6763 (N_6763,N_6090,N_6313);
and U6764 (N_6764,N_6254,N_6169);
nor U6765 (N_6765,N_6218,N_6171);
nand U6766 (N_6766,N_6375,N_6520);
nand U6767 (N_6767,N_6410,N_6075);
or U6768 (N_6768,N_6586,N_6434);
nor U6769 (N_6769,N_6204,N_6100);
or U6770 (N_6770,N_6240,N_6073);
or U6771 (N_6771,N_6199,N_6398);
and U6772 (N_6772,N_6142,N_6278);
and U6773 (N_6773,N_6209,N_6452);
and U6774 (N_6774,N_6648,N_6729);
nor U6775 (N_6775,N_6393,N_6088);
nand U6776 (N_6776,N_6628,N_6409);
nand U6777 (N_6777,N_6462,N_6296);
nand U6778 (N_6778,N_6625,N_6018);
and U6779 (N_6779,N_6086,N_6433);
nand U6780 (N_6780,N_6316,N_6015);
nand U6781 (N_6781,N_6621,N_6505);
nand U6782 (N_6782,N_6089,N_6523);
or U6783 (N_6783,N_6734,N_6573);
nand U6784 (N_6784,N_6238,N_6288);
nor U6785 (N_6785,N_6021,N_6163);
and U6786 (N_6786,N_6704,N_6182);
or U6787 (N_6787,N_6408,N_6599);
nand U6788 (N_6788,N_6168,N_6356);
and U6789 (N_6789,N_6643,N_6099);
or U6790 (N_6790,N_6692,N_6715);
and U6791 (N_6791,N_6242,N_6574);
nor U6792 (N_6792,N_6158,N_6570);
and U6793 (N_6793,N_6435,N_6113);
or U6794 (N_6794,N_6694,N_6051);
nor U6795 (N_6795,N_6110,N_6074);
and U6796 (N_6796,N_6016,N_6691);
nor U6797 (N_6797,N_6693,N_6287);
or U6798 (N_6798,N_6730,N_6217);
or U6799 (N_6799,N_6098,N_6283);
nor U6800 (N_6800,N_6411,N_6629);
and U6801 (N_6801,N_6078,N_6604);
nand U6802 (N_6802,N_6504,N_6450);
nand U6803 (N_6803,N_6426,N_6102);
and U6804 (N_6804,N_6499,N_6206);
and U6805 (N_6805,N_6050,N_6267);
nand U6806 (N_6806,N_6372,N_6070);
nor U6807 (N_6807,N_6183,N_6318);
nand U6808 (N_6808,N_6653,N_6579);
and U6809 (N_6809,N_6525,N_6039);
and U6810 (N_6810,N_6321,N_6065);
and U6811 (N_6811,N_6509,N_6024);
or U6812 (N_6812,N_6323,N_6485);
or U6813 (N_6813,N_6723,N_6087);
or U6814 (N_6814,N_6617,N_6155);
or U6815 (N_6815,N_6063,N_6655);
and U6816 (N_6816,N_6095,N_6170);
or U6817 (N_6817,N_6307,N_6403);
or U6818 (N_6818,N_6735,N_6661);
xor U6819 (N_6819,N_6748,N_6708);
nand U6820 (N_6820,N_6271,N_6080);
nand U6821 (N_6821,N_6680,N_6076);
and U6822 (N_6822,N_6040,N_6608);
nand U6823 (N_6823,N_6516,N_6640);
and U6824 (N_6824,N_6420,N_6417);
and U6825 (N_6825,N_6556,N_6422);
nor U6826 (N_6826,N_6493,N_6732);
nand U6827 (N_6827,N_6418,N_6042);
xor U6828 (N_6828,N_6017,N_6690);
nand U6829 (N_6829,N_6544,N_6044);
nand U6830 (N_6830,N_6533,N_6116);
nor U6831 (N_6831,N_6471,N_6518);
nand U6832 (N_6832,N_6252,N_6214);
nand U6833 (N_6833,N_6592,N_6501);
nor U6834 (N_6834,N_6028,N_6107);
and U6835 (N_6835,N_6285,N_6531);
nand U6836 (N_6836,N_6297,N_6133);
nor U6837 (N_6837,N_6343,N_6233);
and U6838 (N_6838,N_6115,N_6551);
xnor U6839 (N_6839,N_6390,N_6553);
or U6840 (N_6840,N_6440,N_6469);
and U6841 (N_6841,N_6746,N_6624);
and U6842 (N_6842,N_6706,N_6197);
nand U6843 (N_6843,N_6108,N_6695);
or U6844 (N_6844,N_6317,N_6646);
nand U6845 (N_6845,N_6378,N_6507);
and U6846 (N_6846,N_6495,N_6066);
and U6847 (N_6847,N_6446,N_6014);
or U6848 (N_6848,N_6335,N_6344);
nor U6849 (N_6849,N_6645,N_6423);
nor U6850 (N_6850,N_6649,N_6162);
nand U6851 (N_6851,N_6602,N_6008);
xnor U6852 (N_6852,N_6616,N_6487);
or U6853 (N_6853,N_6172,N_6049);
or U6854 (N_6854,N_6451,N_6400);
xor U6855 (N_6855,N_6571,N_6606);
xnor U6856 (N_6856,N_6593,N_6194);
nor U6857 (N_6857,N_6632,N_6043);
and U6858 (N_6858,N_6678,N_6545);
or U6859 (N_6859,N_6581,N_6449);
and U6860 (N_6860,N_6402,N_6031);
nand U6861 (N_6861,N_6486,N_6298);
and U6862 (N_6862,N_6437,N_6262);
nor U6863 (N_6863,N_6697,N_6096);
nand U6864 (N_6864,N_6641,N_6521);
nand U6865 (N_6865,N_6496,N_6213);
or U6866 (N_6866,N_6705,N_6192);
and U6867 (N_6867,N_6510,N_6361);
xnor U6868 (N_6868,N_6247,N_6338);
nand U6869 (N_6869,N_6327,N_6304);
nand U6870 (N_6870,N_6160,N_6707);
or U6871 (N_6871,N_6464,N_6048);
and U6872 (N_6872,N_6167,N_6482);
nand U6873 (N_6873,N_6120,N_6139);
xnor U6874 (N_6874,N_6727,N_6324);
or U6875 (N_6875,N_6749,N_6682);
or U6876 (N_6876,N_6709,N_6532);
xnor U6877 (N_6877,N_6491,N_6166);
or U6878 (N_6878,N_6474,N_6072);
xnor U6879 (N_6879,N_6191,N_6272);
nor U6880 (N_6880,N_6207,N_6293);
nand U6881 (N_6881,N_6414,N_6250);
nand U6882 (N_6882,N_6467,N_6702);
nand U6883 (N_6883,N_6362,N_6527);
nor U6884 (N_6884,N_6371,N_6105);
nand U6885 (N_6885,N_6396,N_6447);
and U6886 (N_6886,N_6263,N_6401);
nand U6887 (N_6887,N_6266,N_6607);
or U6888 (N_6888,N_6558,N_6494);
nor U6889 (N_6889,N_6387,N_6580);
nor U6890 (N_6890,N_6436,N_6244);
xor U6891 (N_6891,N_6226,N_6399);
or U6892 (N_6892,N_6308,N_6281);
nand U6893 (N_6893,N_6610,N_6118);
or U6894 (N_6894,N_6235,N_6314);
nor U6895 (N_6895,N_6548,N_6668);
nor U6896 (N_6896,N_6424,N_6034);
xnor U6897 (N_6897,N_6585,N_6679);
or U6898 (N_6898,N_6141,N_6448);
or U6899 (N_6899,N_6009,N_6228);
nor U6900 (N_6900,N_6148,N_6292);
nand U6901 (N_6901,N_6154,N_6444);
nand U6902 (N_6902,N_6722,N_6660);
nand U6903 (N_6903,N_6475,N_6425);
nand U6904 (N_6904,N_6524,N_6478);
nand U6905 (N_6905,N_6055,N_6470);
or U6906 (N_6906,N_6350,N_6212);
or U6907 (N_6907,N_6377,N_6175);
xnor U6908 (N_6908,N_6612,N_6369);
nand U6909 (N_6909,N_6537,N_6125);
or U6910 (N_6910,N_6582,N_6058);
nor U6911 (N_6911,N_6386,N_6736);
and U6912 (N_6912,N_6472,N_6405);
or U6913 (N_6913,N_6615,N_6060);
nand U6914 (N_6914,N_6686,N_6079);
xor U6915 (N_6915,N_6503,N_6282);
xor U6916 (N_6916,N_6365,N_6502);
and U6917 (N_6917,N_6068,N_6367);
or U6918 (N_6918,N_6306,N_6232);
or U6919 (N_6919,N_6397,N_6134);
and U6920 (N_6920,N_6542,N_6483);
nor U6921 (N_6921,N_6603,N_6032);
or U6922 (N_6922,N_6512,N_6644);
and U6923 (N_6923,N_6081,N_6159);
or U6924 (N_6924,N_6535,N_6563);
and U6925 (N_6925,N_6273,N_6312);
and U6926 (N_6926,N_6636,N_6114);
nand U6927 (N_6927,N_6688,N_6380);
and U6928 (N_6928,N_6560,N_6355);
nand U6929 (N_6929,N_6117,N_6239);
xor U6930 (N_6930,N_6216,N_6284);
and U6931 (N_6931,N_6245,N_6084);
nor U6932 (N_6932,N_6299,N_6453);
xor U6933 (N_6933,N_6265,N_6721);
nand U6934 (N_6934,N_6022,N_6395);
and U6935 (N_6935,N_6174,N_6601);
nand U6936 (N_6936,N_6671,N_6696);
or U6937 (N_6937,N_6569,N_6490);
nor U6938 (N_6938,N_6224,N_6130);
and U6939 (N_6939,N_6187,N_6152);
nand U6940 (N_6940,N_6719,N_6121);
and U6941 (N_6941,N_6623,N_6041);
or U6942 (N_6942,N_6584,N_6295);
nand U6943 (N_6943,N_6202,N_6500);
or U6944 (N_6944,N_6458,N_6346);
xnor U6945 (N_6945,N_6001,N_6161);
and U6946 (N_6946,N_6257,N_6663);
or U6947 (N_6947,N_6007,N_6061);
nand U6948 (N_6948,N_6747,N_6067);
or U6949 (N_6949,N_6492,N_6613);
nand U6950 (N_6950,N_6703,N_6550);
and U6951 (N_6951,N_6020,N_6270);
nor U6952 (N_6952,N_6412,N_6082);
xor U6953 (N_6953,N_6658,N_6195);
or U6954 (N_6954,N_6071,N_6251);
or U6955 (N_6955,N_6374,N_6059);
or U6956 (N_6956,N_6260,N_6203);
nand U6957 (N_6957,N_6700,N_6103);
and U6958 (N_6958,N_6674,N_6030);
nand U6959 (N_6959,N_6559,N_6534);
xnor U6960 (N_6960,N_6315,N_6459);
or U6961 (N_6961,N_6201,N_6083);
nand U6962 (N_6962,N_6258,N_6143);
and U6963 (N_6963,N_6515,N_6328);
or U6964 (N_6964,N_6294,N_6439);
and U6965 (N_6965,N_6611,N_6349);
xnor U6966 (N_6966,N_6476,N_6465);
or U6967 (N_6967,N_6153,N_6618);
nor U6968 (N_6968,N_6320,N_6341);
xnor U6969 (N_6969,N_6144,N_6137);
and U6970 (N_6970,N_6488,N_6670);
and U6971 (N_6971,N_6484,N_6127);
xor U6972 (N_6972,N_6376,N_6246);
or U6973 (N_6973,N_6370,N_6421);
or U6974 (N_6974,N_6151,N_6329);
nor U6975 (N_6975,N_6554,N_6185);
or U6976 (N_6976,N_6650,N_6180);
nand U6977 (N_6977,N_6146,N_6205);
and U6978 (N_6978,N_6305,N_6011);
nor U6979 (N_6979,N_6698,N_6744);
nor U6980 (N_6980,N_6354,N_6481);
or U6981 (N_6981,N_6179,N_6683);
nor U6982 (N_6982,N_6334,N_6119);
nor U6983 (N_6983,N_6046,N_6506);
and U6984 (N_6984,N_6264,N_6633);
nor U6985 (N_6985,N_6236,N_6097);
and U6986 (N_6986,N_6189,N_6069);
nand U6987 (N_6987,N_6415,N_6340);
or U6988 (N_6988,N_6652,N_6373);
and U6989 (N_6989,N_6473,N_6319);
xor U6990 (N_6990,N_6385,N_6587);
nor U6991 (N_6991,N_6546,N_6576);
nand U6992 (N_6992,N_6106,N_6675);
nand U6993 (N_6993,N_6443,N_6511);
nand U6994 (N_6994,N_6064,N_6657);
or U6995 (N_6995,N_6173,N_6345);
and U6996 (N_6996,N_6302,N_6724);
nand U6997 (N_6997,N_6522,N_6025);
nor U6998 (N_6998,N_6131,N_6566);
or U6999 (N_6999,N_6178,N_6513);
or U7000 (N_7000,N_6165,N_6630);
nand U7001 (N_7001,N_6541,N_6358);
nand U7002 (N_7002,N_6164,N_6659);
and U7003 (N_7003,N_6184,N_6508);
nor U7004 (N_7004,N_6589,N_6033);
or U7005 (N_7005,N_6330,N_6514);
nor U7006 (N_7006,N_6177,N_6037);
or U7007 (N_7007,N_6656,N_6394);
and U7008 (N_7008,N_6198,N_6381);
nor U7009 (N_7009,N_6463,N_6456);
and U7010 (N_7010,N_6300,N_6193);
or U7011 (N_7011,N_6441,N_6219);
and U7012 (N_7012,N_6322,N_6145);
and U7013 (N_7013,N_6303,N_6676);
or U7014 (N_7014,N_6222,N_6667);
and U7015 (N_7015,N_6188,N_6339);
xor U7016 (N_7016,N_6045,N_6540);
nand U7017 (N_7017,N_6392,N_6138);
nand U7018 (N_7018,N_6275,N_6109);
or U7019 (N_7019,N_6547,N_6575);
nand U7020 (N_7020,N_6498,N_6052);
nor U7021 (N_7021,N_6594,N_6056);
and U7022 (N_7022,N_6647,N_6227);
or U7023 (N_7023,N_6466,N_6622);
nand U7024 (N_7024,N_6578,N_6389);
or U7025 (N_7025,N_6745,N_6085);
and U7026 (N_7026,N_6225,N_6230);
or U7027 (N_7027,N_6404,N_6363);
nand U7028 (N_7028,N_6104,N_6237);
nor U7029 (N_7029,N_6742,N_6468);
xor U7030 (N_7030,N_6598,N_6712);
or U7031 (N_7031,N_6002,N_6561);
nor U7032 (N_7032,N_6634,N_6062);
and U7033 (N_7033,N_6701,N_6000);
or U7034 (N_7034,N_6639,N_6549);
and U7035 (N_7035,N_6638,N_6432);
nand U7036 (N_7036,N_6132,N_6276);
nor U7037 (N_7037,N_6004,N_6234);
nand U7038 (N_7038,N_6461,N_6190);
xnor U7039 (N_7039,N_6348,N_6687);
nor U7040 (N_7040,N_6325,N_6186);
nor U7041 (N_7041,N_6428,N_6241);
nor U7042 (N_7042,N_6565,N_6057);
and U7043 (N_7043,N_6519,N_6223);
or U7044 (N_7044,N_6023,N_6291);
or U7045 (N_7045,N_6626,N_6637);
xor U7046 (N_7046,N_6564,N_6208);
or U7047 (N_7047,N_6368,N_6631);
or U7048 (N_7048,N_6357,N_6010);
and U7049 (N_7049,N_6047,N_6457);
nor U7050 (N_7050,N_6003,N_6711);
nand U7051 (N_7051,N_6289,N_6269);
or U7052 (N_7052,N_6596,N_6136);
nand U7053 (N_7053,N_6384,N_6477);
nand U7054 (N_7054,N_6360,N_6036);
or U7055 (N_7055,N_6619,N_6200);
and U7056 (N_7056,N_6382,N_6249);
nor U7057 (N_7057,N_6741,N_6430);
or U7058 (N_7058,N_6147,N_6268);
or U7059 (N_7059,N_6718,N_6255);
nor U7060 (N_7060,N_6699,N_6122);
nand U7061 (N_7061,N_6383,N_6347);
or U7062 (N_7062,N_6489,N_6627);
nand U7063 (N_7063,N_6128,N_6157);
and U7064 (N_7064,N_6538,N_6614);
nor U7065 (N_7065,N_6279,N_6651);
xnor U7066 (N_7066,N_6029,N_6609);
and U7067 (N_7067,N_6539,N_6407);
and U7068 (N_7068,N_6027,N_6391);
and U7069 (N_7069,N_6124,N_6311);
xor U7070 (N_7070,N_6526,N_6388);
or U7071 (N_7071,N_6438,N_6353);
and U7072 (N_7072,N_6123,N_6019);
and U7073 (N_7073,N_6588,N_6743);
nor U7074 (N_7074,N_6077,N_6684);
nor U7075 (N_7075,N_6243,N_6597);
and U7076 (N_7076,N_6196,N_6728);
or U7077 (N_7077,N_6738,N_6352);
nand U7078 (N_7078,N_6543,N_6092);
nor U7079 (N_7079,N_6053,N_6445);
and U7080 (N_7080,N_6336,N_6681);
or U7081 (N_7081,N_6366,N_6310);
nor U7082 (N_7082,N_6126,N_6664);
nand U7083 (N_7083,N_6150,N_6256);
nand U7084 (N_7084,N_6156,N_6497);
nor U7085 (N_7085,N_6726,N_6717);
xor U7086 (N_7086,N_6605,N_6006);
or U7087 (N_7087,N_6364,N_6480);
and U7088 (N_7088,N_6220,N_6642);
nor U7089 (N_7089,N_6280,N_6026);
or U7090 (N_7090,N_6529,N_6739);
or U7091 (N_7091,N_6737,N_6454);
nand U7092 (N_7092,N_6666,N_6112);
nand U7093 (N_7093,N_6536,N_6351);
nor U7094 (N_7094,N_6054,N_6714);
nor U7095 (N_7095,N_6211,N_6460);
or U7096 (N_7096,N_6333,N_6662);
and U7097 (N_7097,N_6111,N_6672);
xnor U7098 (N_7098,N_6479,N_6555);
nor U7099 (N_7099,N_6716,N_6731);
and U7100 (N_7100,N_6359,N_6406);
and U7101 (N_7101,N_6665,N_6140);
xor U7102 (N_7102,N_6274,N_6229);
or U7103 (N_7103,N_6261,N_6567);
nor U7104 (N_7104,N_6568,N_6093);
nand U7105 (N_7105,N_6710,N_6530);
nand U7106 (N_7106,N_6253,N_6309);
and U7107 (N_7107,N_6101,N_6654);
nand U7108 (N_7108,N_6215,N_6094);
nor U7109 (N_7109,N_6669,N_6135);
nand U7110 (N_7110,N_6231,N_6635);
nand U7111 (N_7111,N_6332,N_6210);
nand U7112 (N_7112,N_6517,N_6038);
and U7113 (N_7113,N_6590,N_6562);
nor U7114 (N_7114,N_6419,N_6181);
and U7115 (N_7115,N_6557,N_6290);
xnor U7116 (N_7116,N_6413,N_6129);
nand U7117 (N_7117,N_6277,N_6720);
nand U7118 (N_7118,N_6176,N_6337);
and U7119 (N_7119,N_6583,N_6286);
or U7120 (N_7120,N_6600,N_6689);
and U7121 (N_7121,N_6552,N_6733);
nor U7122 (N_7122,N_6431,N_6725);
nand U7123 (N_7123,N_6248,N_6326);
nor U7124 (N_7124,N_6416,N_6091);
nor U7125 (N_7125,N_6465,N_6510);
or U7126 (N_7126,N_6195,N_6191);
xnor U7127 (N_7127,N_6631,N_6714);
and U7128 (N_7128,N_6256,N_6562);
and U7129 (N_7129,N_6517,N_6590);
or U7130 (N_7130,N_6680,N_6459);
and U7131 (N_7131,N_6607,N_6175);
nor U7132 (N_7132,N_6650,N_6646);
and U7133 (N_7133,N_6646,N_6173);
xnor U7134 (N_7134,N_6433,N_6667);
nand U7135 (N_7135,N_6400,N_6643);
and U7136 (N_7136,N_6029,N_6202);
or U7137 (N_7137,N_6079,N_6200);
nor U7138 (N_7138,N_6105,N_6066);
nand U7139 (N_7139,N_6315,N_6100);
or U7140 (N_7140,N_6463,N_6481);
nor U7141 (N_7141,N_6737,N_6148);
nor U7142 (N_7142,N_6503,N_6534);
nand U7143 (N_7143,N_6706,N_6418);
or U7144 (N_7144,N_6640,N_6634);
or U7145 (N_7145,N_6689,N_6642);
xnor U7146 (N_7146,N_6651,N_6329);
nand U7147 (N_7147,N_6136,N_6472);
nand U7148 (N_7148,N_6712,N_6528);
xor U7149 (N_7149,N_6361,N_6661);
nor U7150 (N_7150,N_6252,N_6407);
or U7151 (N_7151,N_6006,N_6528);
nor U7152 (N_7152,N_6614,N_6732);
or U7153 (N_7153,N_6340,N_6360);
and U7154 (N_7154,N_6354,N_6335);
and U7155 (N_7155,N_6087,N_6093);
or U7156 (N_7156,N_6249,N_6092);
xor U7157 (N_7157,N_6109,N_6159);
nand U7158 (N_7158,N_6476,N_6002);
and U7159 (N_7159,N_6666,N_6294);
or U7160 (N_7160,N_6110,N_6318);
nor U7161 (N_7161,N_6034,N_6199);
nor U7162 (N_7162,N_6050,N_6730);
or U7163 (N_7163,N_6359,N_6120);
and U7164 (N_7164,N_6503,N_6002);
and U7165 (N_7165,N_6054,N_6647);
nor U7166 (N_7166,N_6188,N_6209);
or U7167 (N_7167,N_6440,N_6238);
nand U7168 (N_7168,N_6037,N_6062);
and U7169 (N_7169,N_6443,N_6426);
nand U7170 (N_7170,N_6054,N_6157);
or U7171 (N_7171,N_6109,N_6477);
or U7172 (N_7172,N_6656,N_6711);
nor U7173 (N_7173,N_6635,N_6666);
nand U7174 (N_7174,N_6256,N_6326);
or U7175 (N_7175,N_6012,N_6220);
nor U7176 (N_7176,N_6271,N_6619);
or U7177 (N_7177,N_6375,N_6569);
or U7178 (N_7178,N_6196,N_6130);
xnor U7179 (N_7179,N_6144,N_6614);
and U7180 (N_7180,N_6654,N_6042);
or U7181 (N_7181,N_6162,N_6197);
nor U7182 (N_7182,N_6426,N_6604);
and U7183 (N_7183,N_6487,N_6497);
nand U7184 (N_7184,N_6399,N_6322);
or U7185 (N_7185,N_6601,N_6356);
nand U7186 (N_7186,N_6535,N_6092);
and U7187 (N_7187,N_6438,N_6171);
nand U7188 (N_7188,N_6735,N_6745);
nand U7189 (N_7189,N_6606,N_6081);
nor U7190 (N_7190,N_6078,N_6645);
or U7191 (N_7191,N_6444,N_6096);
nand U7192 (N_7192,N_6452,N_6546);
nor U7193 (N_7193,N_6119,N_6235);
and U7194 (N_7194,N_6659,N_6447);
nor U7195 (N_7195,N_6514,N_6648);
nand U7196 (N_7196,N_6352,N_6495);
or U7197 (N_7197,N_6188,N_6740);
xor U7198 (N_7198,N_6618,N_6156);
and U7199 (N_7199,N_6621,N_6272);
and U7200 (N_7200,N_6342,N_6310);
nor U7201 (N_7201,N_6469,N_6360);
nand U7202 (N_7202,N_6004,N_6647);
and U7203 (N_7203,N_6749,N_6642);
nor U7204 (N_7204,N_6327,N_6320);
and U7205 (N_7205,N_6567,N_6161);
and U7206 (N_7206,N_6303,N_6672);
or U7207 (N_7207,N_6320,N_6133);
or U7208 (N_7208,N_6365,N_6636);
nor U7209 (N_7209,N_6357,N_6271);
nand U7210 (N_7210,N_6003,N_6703);
or U7211 (N_7211,N_6634,N_6397);
and U7212 (N_7212,N_6705,N_6534);
or U7213 (N_7213,N_6674,N_6286);
nor U7214 (N_7214,N_6558,N_6161);
nand U7215 (N_7215,N_6047,N_6141);
nor U7216 (N_7216,N_6525,N_6419);
or U7217 (N_7217,N_6598,N_6025);
xor U7218 (N_7218,N_6687,N_6377);
nor U7219 (N_7219,N_6383,N_6540);
or U7220 (N_7220,N_6050,N_6387);
nor U7221 (N_7221,N_6088,N_6074);
or U7222 (N_7222,N_6357,N_6296);
nand U7223 (N_7223,N_6030,N_6377);
or U7224 (N_7224,N_6652,N_6045);
nor U7225 (N_7225,N_6494,N_6485);
or U7226 (N_7226,N_6163,N_6705);
nor U7227 (N_7227,N_6597,N_6139);
or U7228 (N_7228,N_6692,N_6140);
or U7229 (N_7229,N_6627,N_6434);
nand U7230 (N_7230,N_6217,N_6578);
nand U7231 (N_7231,N_6327,N_6330);
nor U7232 (N_7232,N_6645,N_6113);
nand U7233 (N_7233,N_6380,N_6276);
nand U7234 (N_7234,N_6167,N_6420);
xnor U7235 (N_7235,N_6508,N_6226);
nor U7236 (N_7236,N_6494,N_6295);
nand U7237 (N_7237,N_6682,N_6195);
xnor U7238 (N_7238,N_6389,N_6698);
nor U7239 (N_7239,N_6586,N_6556);
xnor U7240 (N_7240,N_6037,N_6204);
nor U7241 (N_7241,N_6300,N_6430);
nand U7242 (N_7242,N_6319,N_6135);
nand U7243 (N_7243,N_6340,N_6272);
nor U7244 (N_7244,N_6679,N_6343);
xor U7245 (N_7245,N_6221,N_6622);
nand U7246 (N_7246,N_6226,N_6001);
and U7247 (N_7247,N_6104,N_6044);
nand U7248 (N_7248,N_6713,N_6239);
or U7249 (N_7249,N_6211,N_6616);
nand U7250 (N_7250,N_6319,N_6468);
nand U7251 (N_7251,N_6524,N_6592);
and U7252 (N_7252,N_6389,N_6714);
or U7253 (N_7253,N_6100,N_6559);
xor U7254 (N_7254,N_6538,N_6128);
nor U7255 (N_7255,N_6438,N_6455);
or U7256 (N_7256,N_6259,N_6227);
nand U7257 (N_7257,N_6748,N_6029);
nor U7258 (N_7258,N_6269,N_6170);
or U7259 (N_7259,N_6618,N_6604);
nand U7260 (N_7260,N_6422,N_6307);
and U7261 (N_7261,N_6672,N_6525);
xor U7262 (N_7262,N_6705,N_6357);
nand U7263 (N_7263,N_6644,N_6556);
nand U7264 (N_7264,N_6449,N_6712);
and U7265 (N_7265,N_6355,N_6198);
and U7266 (N_7266,N_6170,N_6134);
or U7267 (N_7267,N_6091,N_6542);
xnor U7268 (N_7268,N_6238,N_6010);
or U7269 (N_7269,N_6046,N_6726);
nand U7270 (N_7270,N_6622,N_6049);
and U7271 (N_7271,N_6471,N_6407);
and U7272 (N_7272,N_6447,N_6090);
nor U7273 (N_7273,N_6428,N_6180);
or U7274 (N_7274,N_6355,N_6344);
nand U7275 (N_7275,N_6179,N_6656);
nand U7276 (N_7276,N_6054,N_6600);
nand U7277 (N_7277,N_6436,N_6349);
or U7278 (N_7278,N_6578,N_6019);
nor U7279 (N_7279,N_6711,N_6508);
nand U7280 (N_7280,N_6640,N_6531);
or U7281 (N_7281,N_6566,N_6534);
nand U7282 (N_7282,N_6565,N_6207);
nor U7283 (N_7283,N_6591,N_6535);
xnor U7284 (N_7284,N_6329,N_6548);
nand U7285 (N_7285,N_6149,N_6083);
xnor U7286 (N_7286,N_6713,N_6356);
and U7287 (N_7287,N_6194,N_6238);
xor U7288 (N_7288,N_6336,N_6731);
nand U7289 (N_7289,N_6508,N_6018);
or U7290 (N_7290,N_6182,N_6419);
or U7291 (N_7291,N_6625,N_6381);
nand U7292 (N_7292,N_6387,N_6261);
nor U7293 (N_7293,N_6530,N_6226);
nor U7294 (N_7294,N_6174,N_6749);
nor U7295 (N_7295,N_6553,N_6655);
and U7296 (N_7296,N_6693,N_6253);
nor U7297 (N_7297,N_6448,N_6153);
or U7298 (N_7298,N_6618,N_6209);
and U7299 (N_7299,N_6342,N_6641);
nand U7300 (N_7300,N_6441,N_6068);
or U7301 (N_7301,N_6171,N_6656);
nor U7302 (N_7302,N_6059,N_6443);
xnor U7303 (N_7303,N_6181,N_6627);
nand U7304 (N_7304,N_6040,N_6408);
and U7305 (N_7305,N_6680,N_6239);
nor U7306 (N_7306,N_6404,N_6004);
nor U7307 (N_7307,N_6028,N_6141);
or U7308 (N_7308,N_6552,N_6581);
xnor U7309 (N_7309,N_6326,N_6288);
or U7310 (N_7310,N_6161,N_6687);
xor U7311 (N_7311,N_6456,N_6378);
and U7312 (N_7312,N_6352,N_6156);
nor U7313 (N_7313,N_6120,N_6718);
nand U7314 (N_7314,N_6387,N_6708);
nor U7315 (N_7315,N_6670,N_6126);
or U7316 (N_7316,N_6500,N_6643);
and U7317 (N_7317,N_6078,N_6308);
or U7318 (N_7318,N_6130,N_6077);
and U7319 (N_7319,N_6088,N_6570);
nor U7320 (N_7320,N_6443,N_6673);
and U7321 (N_7321,N_6543,N_6211);
and U7322 (N_7322,N_6571,N_6227);
and U7323 (N_7323,N_6570,N_6299);
and U7324 (N_7324,N_6660,N_6344);
and U7325 (N_7325,N_6262,N_6205);
nor U7326 (N_7326,N_6062,N_6563);
nand U7327 (N_7327,N_6162,N_6722);
nand U7328 (N_7328,N_6464,N_6528);
nand U7329 (N_7329,N_6178,N_6080);
or U7330 (N_7330,N_6571,N_6143);
and U7331 (N_7331,N_6095,N_6602);
and U7332 (N_7332,N_6314,N_6553);
xnor U7333 (N_7333,N_6044,N_6186);
nor U7334 (N_7334,N_6454,N_6196);
and U7335 (N_7335,N_6001,N_6187);
nor U7336 (N_7336,N_6355,N_6345);
or U7337 (N_7337,N_6307,N_6626);
nor U7338 (N_7338,N_6449,N_6575);
nor U7339 (N_7339,N_6434,N_6567);
nor U7340 (N_7340,N_6256,N_6009);
nor U7341 (N_7341,N_6043,N_6484);
or U7342 (N_7342,N_6708,N_6619);
or U7343 (N_7343,N_6300,N_6221);
and U7344 (N_7344,N_6599,N_6092);
or U7345 (N_7345,N_6241,N_6022);
xor U7346 (N_7346,N_6176,N_6693);
and U7347 (N_7347,N_6329,N_6019);
nand U7348 (N_7348,N_6080,N_6700);
or U7349 (N_7349,N_6201,N_6410);
and U7350 (N_7350,N_6329,N_6054);
nor U7351 (N_7351,N_6664,N_6322);
or U7352 (N_7352,N_6015,N_6448);
nand U7353 (N_7353,N_6608,N_6249);
xor U7354 (N_7354,N_6688,N_6226);
xnor U7355 (N_7355,N_6042,N_6415);
nand U7356 (N_7356,N_6559,N_6273);
nor U7357 (N_7357,N_6077,N_6033);
and U7358 (N_7358,N_6122,N_6097);
and U7359 (N_7359,N_6198,N_6591);
nand U7360 (N_7360,N_6661,N_6684);
nand U7361 (N_7361,N_6420,N_6475);
xor U7362 (N_7362,N_6020,N_6314);
nor U7363 (N_7363,N_6651,N_6536);
or U7364 (N_7364,N_6029,N_6624);
or U7365 (N_7365,N_6067,N_6579);
and U7366 (N_7366,N_6423,N_6138);
xor U7367 (N_7367,N_6098,N_6612);
nand U7368 (N_7368,N_6365,N_6057);
or U7369 (N_7369,N_6462,N_6346);
or U7370 (N_7370,N_6294,N_6694);
and U7371 (N_7371,N_6526,N_6168);
or U7372 (N_7372,N_6334,N_6715);
nor U7373 (N_7373,N_6519,N_6375);
and U7374 (N_7374,N_6096,N_6274);
and U7375 (N_7375,N_6406,N_6576);
nor U7376 (N_7376,N_6153,N_6140);
or U7377 (N_7377,N_6602,N_6229);
nand U7378 (N_7378,N_6732,N_6686);
nand U7379 (N_7379,N_6631,N_6311);
and U7380 (N_7380,N_6061,N_6580);
nand U7381 (N_7381,N_6608,N_6020);
and U7382 (N_7382,N_6334,N_6090);
nand U7383 (N_7383,N_6715,N_6457);
or U7384 (N_7384,N_6703,N_6086);
and U7385 (N_7385,N_6661,N_6104);
and U7386 (N_7386,N_6128,N_6202);
and U7387 (N_7387,N_6118,N_6373);
or U7388 (N_7388,N_6326,N_6514);
and U7389 (N_7389,N_6591,N_6416);
nor U7390 (N_7390,N_6191,N_6113);
and U7391 (N_7391,N_6482,N_6156);
and U7392 (N_7392,N_6047,N_6348);
or U7393 (N_7393,N_6287,N_6597);
and U7394 (N_7394,N_6685,N_6677);
and U7395 (N_7395,N_6098,N_6108);
or U7396 (N_7396,N_6062,N_6170);
xnor U7397 (N_7397,N_6734,N_6128);
and U7398 (N_7398,N_6067,N_6607);
nor U7399 (N_7399,N_6177,N_6201);
or U7400 (N_7400,N_6162,N_6083);
and U7401 (N_7401,N_6008,N_6182);
nand U7402 (N_7402,N_6257,N_6066);
nor U7403 (N_7403,N_6655,N_6404);
nand U7404 (N_7404,N_6193,N_6421);
nor U7405 (N_7405,N_6167,N_6062);
nand U7406 (N_7406,N_6416,N_6624);
and U7407 (N_7407,N_6034,N_6319);
and U7408 (N_7408,N_6176,N_6212);
or U7409 (N_7409,N_6221,N_6608);
xnor U7410 (N_7410,N_6647,N_6147);
nor U7411 (N_7411,N_6440,N_6073);
or U7412 (N_7412,N_6358,N_6317);
and U7413 (N_7413,N_6479,N_6292);
and U7414 (N_7414,N_6115,N_6613);
or U7415 (N_7415,N_6314,N_6617);
and U7416 (N_7416,N_6378,N_6721);
nand U7417 (N_7417,N_6127,N_6364);
nor U7418 (N_7418,N_6180,N_6381);
and U7419 (N_7419,N_6724,N_6151);
and U7420 (N_7420,N_6722,N_6454);
and U7421 (N_7421,N_6254,N_6640);
nand U7422 (N_7422,N_6562,N_6282);
or U7423 (N_7423,N_6608,N_6247);
nor U7424 (N_7424,N_6571,N_6433);
xor U7425 (N_7425,N_6028,N_6097);
nor U7426 (N_7426,N_6747,N_6457);
and U7427 (N_7427,N_6160,N_6640);
and U7428 (N_7428,N_6364,N_6169);
nor U7429 (N_7429,N_6315,N_6609);
or U7430 (N_7430,N_6416,N_6575);
and U7431 (N_7431,N_6042,N_6729);
and U7432 (N_7432,N_6559,N_6555);
nor U7433 (N_7433,N_6559,N_6405);
and U7434 (N_7434,N_6739,N_6034);
xor U7435 (N_7435,N_6087,N_6383);
xnor U7436 (N_7436,N_6360,N_6364);
nand U7437 (N_7437,N_6465,N_6121);
and U7438 (N_7438,N_6292,N_6074);
nand U7439 (N_7439,N_6292,N_6573);
nor U7440 (N_7440,N_6342,N_6492);
and U7441 (N_7441,N_6472,N_6434);
nand U7442 (N_7442,N_6611,N_6186);
and U7443 (N_7443,N_6016,N_6521);
and U7444 (N_7444,N_6296,N_6420);
and U7445 (N_7445,N_6019,N_6157);
or U7446 (N_7446,N_6728,N_6044);
nand U7447 (N_7447,N_6012,N_6175);
or U7448 (N_7448,N_6024,N_6307);
nand U7449 (N_7449,N_6231,N_6058);
and U7450 (N_7450,N_6142,N_6647);
nand U7451 (N_7451,N_6018,N_6484);
nand U7452 (N_7452,N_6538,N_6372);
or U7453 (N_7453,N_6274,N_6243);
or U7454 (N_7454,N_6278,N_6443);
xor U7455 (N_7455,N_6433,N_6604);
nor U7456 (N_7456,N_6410,N_6129);
nand U7457 (N_7457,N_6148,N_6334);
xnor U7458 (N_7458,N_6443,N_6587);
nand U7459 (N_7459,N_6575,N_6476);
nand U7460 (N_7460,N_6478,N_6438);
or U7461 (N_7461,N_6550,N_6142);
and U7462 (N_7462,N_6207,N_6503);
and U7463 (N_7463,N_6426,N_6289);
or U7464 (N_7464,N_6726,N_6357);
nor U7465 (N_7465,N_6078,N_6036);
or U7466 (N_7466,N_6328,N_6700);
nor U7467 (N_7467,N_6523,N_6303);
and U7468 (N_7468,N_6201,N_6441);
or U7469 (N_7469,N_6250,N_6438);
or U7470 (N_7470,N_6641,N_6231);
and U7471 (N_7471,N_6050,N_6644);
nor U7472 (N_7472,N_6302,N_6330);
nand U7473 (N_7473,N_6233,N_6727);
nand U7474 (N_7474,N_6295,N_6134);
or U7475 (N_7475,N_6149,N_6199);
nand U7476 (N_7476,N_6441,N_6184);
and U7477 (N_7477,N_6554,N_6050);
or U7478 (N_7478,N_6507,N_6742);
nor U7479 (N_7479,N_6200,N_6616);
nor U7480 (N_7480,N_6597,N_6331);
nor U7481 (N_7481,N_6717,N_6432);
or U7482 (N_7482,N_6224,N_6135);
nor U7483 (N_7483,N_6442,N_6502);
nor U7484 (N_7484,N_6715,N_6367);
nand U7485 (N_7485,N_6254,N_6069);
nand U7486 (N_7486,N_6115,N_6686);
and U7487 (N_7487,N_6733,N_6162);
nor U7488 (N_7488,N_6032,N_6639);
nor U7489 (N_7489,N_6127,N_6450);
and U7490 (N_7490,N_6535,N_6215);
nor U7491 (N_7491,N_6604,N_6637);
nand U7492 (N_7492,N_6568,N_6383);
and U7493 (N_7493,N_6128,N_6124);
and U7494 (N_7494,N_6520,N_6087);
nor U7495 (N_7495,N_6742,N_6658);
nor U7496 (N_7496,N_6268,N_6674);
and U7497 (N_7497,N_6132,N_6274);
xnor U7498 (N_7498,N_6096,N_6021);
and U7499 (N_7499,N_6066,N_6696);
or U7500 (N_7500,N_7143,N_6964);
nor U7501 (N_7501,N_7271,N_7374);
and U7502 (N_7502,N_7326,N_7097);
nor U7503 (N_7503,N_7327,N_7165);
xor U7504 (N_7504,N_6854,N_7109);
nor U7505 (N_7505,N_7098,N_7016);
nor U7506 (N_7506,N_6929,N_7434);
nor U7507 (N_7507,N_6855,N_7406);
nor U7508 (N_7508,N_6985,N_7333);
nor U7509 (N_7509,N_6901,N_6918);
xor U7510 (N_7510,N_7226,N_6882);
and U7511 (N_7511,N_6891,N_7268);
and U7512 (N_7512,N_6879,N_6923);
and U7513 (N_7513,N_7070,N_6813);
and U7514 (N_7514,N_7186,N_7026);
nor U7515 (N_7515,N_7207,N_6916);
or U7516 (N_7516,N_6755,N_6806);
nor U7517 (N_7517,N_7339,N_7276);
nor U7518 (N_7518,N_6759,N_7291);
and U7519 (N_7519,N_7308,N_6839);
and U7520 (N_7520,N_7346,N_7388);
and U7521 (N_7521,N_6761,N_7487);
nor U7522 (N_7522,N_7477,N_7221);
and U7523 (N_7523,N_7118,N_7203);
xnor U7524 (N_7524,N_6953,N_6778);
nand U7525 (N_7525,N_7068,N_7037);
nor U7526 (N_7526,N_7412,N_7454);
nand U7527 (N_7527,N_7114,N_7058);
and U7528 (N_7528,N_6851,N_7435);
nor U7529 (N_7529,N_7019,N_7088);
or U7530 (N_7530,N_6814,N_6750);
or U7531 (N_7531,N_6857,N_6769);
or U7532 (N_7532,N_7463,N_7174);
or U7533 (N_7533,N_6856,N_7311);
or U7534 (N_7534,N_7345,N_6842);
nand U7535 (N_7535,N_6995,N_7023);
or U7536 (N_7536,N_6804,N_6858);
nor U7537 (N_7537,N_7307,N_6908);
or U7538 (N_7538,N_7177,N_7219);
nor U7539 (N_7539,N_6961,N_7001);
or U7540 (N_7540,N_6897,N_7384);
or U7541 (N_7541,N_6878,N_7036);
and U7542 (N_7542,N_7314,N_7084);
and U7543 (N_7543,N_7257,N_6817);
or U7544 (N_7544,N_7113,N_7061);
and U7545 (N_7545,N_7330,N_7139);
nand U7546 (N_7546,N_6773,N_7282);
nand U7547 (N_7547,N_6792,N_6799);
and U7548 (N_7548,N_6890,N_6903);
or U7549 (N_7549,N_7022,N_7238);
nor U7550 (N_7550,N_7076,N_6788);
nand U7551 (N_7551,N_6990,N_6979);
or U7552 (N_7552,N_7293,N_7250);
nor U7553 (N_7553,N_7364,N_6829);
and U7554 (N_7554,N_7427,N_7089);
or U7555 (N_7555,N_7342,N_7285);
nand U7556 (N_7556,N_7156,N_6906);
xor U7557 (N_7557,N_6777,N_7056);
or U7558 (N_7558,N_7103,N_7242);
nor U7559 (N_7559,N_6866,N_7252);
nand U7560 (N_7560,N_7087,N_6950);
and U7561 (N_7561,N_7481,N_7366);
nand U7562 (N_7562,N_6970,N_7063);
or U7563 (N_7563,N_7440,N_6904);
xor U7564 (N_7564,N_6931,N_7132);
or U7565 (N_7565,N_7377,N_6927);
or U7566 (N_7566,N_6789,N_7264);
and U7567 (N_7567,N_6768,N_7353);
and U7568 (N_7568,N_7310,N_7192);
or U7569 (N_7569,N_7158,N_7073);
nor U7570 (N_7570,N_7079,N_7419);
nand U7571 (N_7571,N_6946,N_7338);
or U7572 (N_7572,N_7413,N_7441);
and U7573 (N_7573,N_7255,N_6939);
nor U7574 (N_7574,N_6885,N_7205);
nor U7575 (N_7575,N_7395,N_7197);
nor U7576 (N_7576,N_7298,N_6887);
nand U7577 (N_7577,N_6977,N_7410);
nor U7578 (N_7578,N_7288,N_7270);
nor U7579 (N_7579,N_7379,N_7489);
nor U7580 (N_7580,N_6902,N_7124);
nand U7581 (N_7581,N_7052,N_6998);
xor U7582 (N_7582,N_7086,N_7332);
nor U7583 (N_7583,N_7455,N_7072);
nand U7584 (N_7584,N_6968,N_7240);
nand U7585 (N_7585,N_7361,N_7290);
or U7586 (N_7586,N_6880,N_7040);
nor U7587 (N_7587,N_7018,N_7220);
xnor U7588 (N_7588,N_6756,N_7466);
nand U7589 (N_7589,N_7015,N_6774);
and U7590 (N_7590,N_6986,N_6965);
and U7591 (N_7591,N_7033,N_7230);
and U7592 (N_7592,N_7488,N_7247);
or U7593 (N_7593,N_6760,N_7204);
xor U7594 (N_7594,N_7127,N_6919);
or U7595 (N_7595,N_7005,N_7337);
nor U7596 (N_7596,N_6925,N_6809);
or U7597 (N_7597,N_7336,N_7301);
and U7598 (N_7598,N_7246,N_7415);
nand U7599 (N_7599,N_7281,N_7065);
or U7600 (N_7600,N_6975,N_6996);
and U7601 (N_7601,N_7299,N_7212);
nor U7602 (N_7602,N_7468,N_6871);
nand U7603 (N_7603,N_6987,N_7224);
nor U7604 (N_7604,N_7323,N_7331);
nand U7605 (N_7605,N_7400,N_7106);
or U7606 (N_7606,N_6958,N_7320);
nand U7607 (N_7607,N_7296,N_7119);
nand U7608 (N_7608,N_6971,N_7344);
nand U7609 (N_7609,N_7453,N_7451);
nand U7610 (N_7610,N_7375,N_7425);
and U7611 (N_7611,N_7049,N_7222);
xnor U7612 (N_7612,N_7272,N_7141);
nand U7613 (N_7613,N_7128,N_6909);
nor U7614 (N_7614,N_7032,N_7117);
xor U7615 (N_7615,N_7152,N_7029);
nor U7616 (N_7616,N_6988,N_7162);
nor U7617 (N_7617,N_7396,N_7316);
xor U7618 (N_7618,N_7008,N_7045);
nor U7619 (N_7619,N_6831,N_7459);
or U7620 (N_7620,N_7209,N_6811);
nor U7621 (N_7621,N_7229,N_7160);
nor U7622 (N_7622,N_6973,N_7107);
or U7623 (N_7623,N_6924,N_6934);
or U7624 (N_7624,N_6841,N_7499);
nor U7625 (N_7625,N_6893,N_7325);
nand U7626 (N_7626,N_6805,N_7074);
or U7627 (N_7627,N_7357,N_7433);
nor U7628 (N_7628,N_7467,N_7329);
nor U7629 (N_7629,N_6981,N_7170);
and U7630 (N_7630,N_6932,N_7075);
or U7631 (N_7631,N_6818,N_7389);
nor U7632 (N_7632,N_7414,N_6933);
and U7633 (N_7633,N_6948,N_6942);
and U7634 (N_7634,N_6960,N_7085);
nor U7635 (N_7635,N_7111,N_7398);
or U7636 (N_7636,N_6894,N_7360);
or U7637 (N_7637,N_7334,N_7393);
and U7638 (N_7638,N_6983,N_7025);
nor U7639 (N_7639,N_6785,N_7475);
nor U7640 (N_7640,N_6848,N_7173);
nand U7641 (N_7641,N_7116,N_6819);
or U7642 (N_7642,N_6928,N_6826);
nor U7643 (N_7643,N_7274,N_7178);
or U7644 (N_7644,N_6993,N_7135);
xnor U7645 (N_7645,N_7367,N_6867);
xor U7646 (N_7646,N_6888,N_7447);
and U7647 (N_7647,N_7129,N_7067);
nand U7648 (N_7648,N_6849,N_7010);
and U7649 (N_7649,N_6824,N_6997);
nor U7650 (N_7650,N_7034,N_6763);
xnor U7651 (N_7651,N_7014,N_6766);
nand U7652 (N_7652,N_6816,N_7269);
and U7653 (N_7653,N_7133,N_7267);
or U7654 (N_7654,N_7385,N_7404);
and U7655 (N_7655,N_7234,N_7387);
nor U7656 (N_7656,N_7243,N_7258);
nor U7657 (N_7657,N_7217,N_7245);
and U7658 (N_7658,N_7408,N_6786);
nor U7659 (N_7659,N_7275,N_7402);
xor U7660 (N_7660,N_7095,N_7464);
nor U7661 (N_7661,N_6803,N_6984);
nand U7662 (N_7662,N_6907,N_6812);
and U7663 (N_7663,N_7225,N_6876);
xnor U7664 (N_7664,N_7066,N_7090);
nor U7665 (N_7665,N_7436,N_6846);
and U7666 (N_7666,N_6830,N_7493);
xor U7667 (N_7667,N_7028,N_7130);
and U7668 (N_7668,N_6827,N_6943);
nor U7669 (N_7669,N_7381,N_6914);
or U7670 (N_7670,N_7420,N_6808);
or U7671 (N_7671,N_6850,N_7416);
nand U7672 (N_7672,N_6938,N_7154);
nand U7673 (N_7673,N_7083,N_7071);
and U7674 (N_7674,N_6797,N_7047);
and U7675 (N_7675,N_7491,N_7465);
and U7676 (N_7676,N_7305,N_6779);
nor U7677 (N_7677,N_6800,N_6757);
nor U7678 (N_7678,N_6832,N_7142);
and U7679 (N_7679,N_7253,N_6853);
and U7680 (N_7680,N_7003,N_7053);
and U7681 (N_7681,N_6962,N_6751);
nor U7682 (N_7682,N_7069,N_6767);
and U7683 (N_7683,N_7369,N_6991);
and U7684 (N_7684,N_6825,N_6959);
and U7685 (N_7685,N_6884,N_7159);
nor U7686 (N_7686,N_6917,N_7429);
nand U7687 (N_7687,N_7448,N_7140);
or U7688 (N_7688,N_6921,N_7137);
or U7689 (N_7689,N_6772,N_7373);
and U7690 (N_7690,N_7030,N_7313);
and U7691 (N_7691,N_7304,N_7359);
xor U7692 (N_7692,N_7055,N_7254);
and U7693 (N_7693,N_7363,N_7490);
nand U7694 (N_7694,N_7241,N_7403);
xnor U7695 (N_7695,N_6967,N_6807);
xor U7696 (N_7696,N_6784,N_7108);
or U7697 (N_7697,N_7100,N_7233);
and U7698 (N_7698,N_7421,N_6838);
or U7699 (N_7699,N_6912,N_7153);
nor U7700 (N_7700,N_7312,N_6873);
or U7701 (N_7701,N_7321,N_6859);
and U7702 (N_7702,N_7042,N_6920);
xor U7703 (N_7703,N_6911,N_7289);
or U7704 (N_7704,N_6793,N_7223);
nor U7705 (N_7705,N_7306,N_7214);
or U7706 (N_7706,N_7432,N_6947);
and U7707 (N_7707,N_6810,N_7000);
and U7708 (N_7708,N_7147,N_7190);
or U7709 (N_7709,N_7007,N_7460);
nand U7710 (N_7710,N_7101,N_6883);
xnor U7711 (N_7711,N_7232,N_6820);
nor U7712 (N_7712,N_7409,N_7266);
xnor U7713 (N_7713,N_6865,N_6869);
or U7714 (N_7714,N_7188,N_7462);
or U7715 (N_7715,N_7169,N_6840);
xor U7716 (N_7716,N_6999,N_6780);
xnor U7717 (N_7717,N_7191,N_6944);
and U7718 (N_7718,N_7411,N_7202);
nand U7719 (N_7719,N_7105,N_7057);
nand U7720 (N_7720,N_7110,N_7138);
xor U7721 (N_7721,N_7206,N_7256);
or U7722 (N_7722,N_7430,N_7372);
xnor U7723 (N_7723,N_7031,N_7417);
and U7724 (N_7724,N_7080,N_6776);
nand U7725 (N_7725,N_7213,N_7335);
and U7726 (N_7726,N_7355,N_7021);
xor U7727 (N_7727,N_7497,N_6910);
and U7728 (N_7728,N_7060,N_7300);
and U7729 (N_7729,N_7445,N_6992);
nand U7730 (N_7730,N_7343,N_6822);
or U7731 (N_7731,N_7422,N_7450);
nor U7732 (N_7732,N_7350,N_6941);
xor U7733 (N_7733,N_7131,N_7161);
or U7734 (N_7734,N_7437,N_6994);
nor U7735 (N_7735,N_7494,N_6926);
or U7736 (N_7736,N_6833,N_6781);
or U7737 (N_7737,N_7446,N_6874);
nand U7738 (N_7738,N_7341,N_7194);
nand U7739 (N_7739,N_7172,N_6836);
or U7740 (N_7740,N_7017,N_6936);
and U7741 (N_7741,N_7231,N_7283);
and U7742 (N_7742,N_6886,N_7315);
or U7743 (N_7743,N_6796,N_6852);
or U7744 (N_7744,N_7349,N_7237);
and U7745 (N_7745,N_7328,N_7151);
nand U7746 (N_7746,N_7235,N_7309);
and U7747 (N_7747,N_7486,N_7050);
nand U7748 (N_7748,N_6954,N_7498);
and U7749 (N_7749,N_7157,N_6783);
nand U7750 (N_7750,N_7041,N_7122);
and U7751 (N_7751,N_7444,N_7352);
nor U7752 (N_7752,N_7492,N_7473);
or U7753 (N_7753,N_6801,N_7148);
nor U7754 (N_7754,N_6870,N_7145);
nand U7755 (N_7755,N_7284,N_6847);
nor U7756 (N_7756,N_7469,N_7262);
nor U7757 (N_7757,N_7399,N_7048);
nor U7758 (N_7758,N_7039,N_7059);
or U7759 (N_7759,N_7370,N_7391);
nor U7760 (N_7760,N_7279,N_7368);
nand U7761 (N_7761,N_7193,N_7009);
nand U7762 (N_7762,N_7166,N_7092);
nor U7763 (N_7763,N_6753,N_7397);
nor U7764 (N_7764,N_7259,N_7348);
and U7765 (N_7765,N_7164,N_7358);
nand U7766 (N_7766,N_7249,N_7251);
nor U7767 (N_7767,N_6989,N_7297);
or U7768 (N_7768,N_7483,N_6758);
or U7769 (N_7769,N_6872,N_7215);
and U7770 (N_7770,N_6913,N_7163);
or U7771 (N_7771,N_7184,N_7295);
or U7772 (N_7772,N_7176,N_6875);
nor U7773 (N_7773,N_7096,N_6982);
nand U7774 (N_7774,N_7286,N_7362);
or U7775 (N_7775,N_7155,N_7054);
or U7776 (N_7776,N_7189,N_6815);
and U7777 (N_7777,N_7144,N_7024);
or U7778 (N_7778,N_7418,N_6864);
nor U7779 (N_7779,N_7405,N_7248);
nand U7780 (N_7780,N_7277,N_7324);
and U7781 (N_7781,N_6863,N_6896);
or U7782 (N_7782,N_7102,N_7392);
xnor U7783 (N_7783,N_7123,N_7126);
nor U7784 (N_7784,N_7201,N_7175);
nor U7785 (N_7785,N_7120,N_7091);
nand U7786 (N_7786,N_6956,N_6951);
nor U7787 (N_7787,N_6899,N_7423);
and U7788 (N_7788,N_7187,N_7479);
or U7789 (N_7789,N_7263,N_7287);
and U7790 (N_7790,N_7317,N_6940);
xor U7791 (N_7791,N_7260,N_6762);
nand U7792 (N_7792,N_7171,N_6862);
xnor U7793 (N_7793,N_7093,N_7182);
and U7794 (N_7794,N_6843,N_6844);
and U7795 (N_7795,N_7011,N_7179);
nand U7796 (N_7796,N_7484,N_7004);
and U7797 (N_7797,N_6949,N_7401);
xor U7798 (N_7798,N_7064,N_7294);
and U7799 (N_7799,N_6790,N_7208);
nor U7800 (N_7800,N_6972,N_7051);
nand U7801 (N_7801,N_7078,N_7495);
nor U7802 (N_7802,N_7496,N_7211);
or U7803 (N_7803,N_7236,N_7077);
nand U7804 (N_7804,N_7472,N_7121);
nand U7805 (N_7805,N_7081,N_6935);
or U7806 (N_7806,N_6881,N_7196);
nor U7807 (N_7807,N_7480,N_7386);
or U7808 (N_7808,N_7244,N_7485);
or U7809 (N_7809,N_7380,N_6765);
nor U7810 (N_7810,N_7183,N_7002);
nor U7811 (N_7811,N_7347,N_7438);
nor U7812 (N_7812,N_6752,N_7340);
nand U7813 (N_7813,N_6754,N_6861);
nand U7814 (N_7814,N_7318,N_6930);
and U7815 (N_7815,N_7394,N_7216);
nor U7816 (N_7816,N_7146,N_7371);
and U7817 (N_7817,N_6828,N_7471);
or U7818 (N_7818,N_7125,N_6976);
or U7819 (N_7819,N_7227,N_7150);
or U7820 (N_7820,N_6969,N_6775);
nand U7821 (N_7821,N_7378,N_7167);
and U7822 (N_7822,N_6802,N_7426);
xor U7823 (N_7823,N_7354,N_6966);
and U7824 (N_7824,N_6837,N_7383);
or U7825 (N_7825,N_6795,N_7046);
nor U7826 (N_7826,N_6892,N_6868);
nand U7827 (N_7827,N_7112,N_7278);
or U7828 (N_7828,N_6945,N_7006);
and U7829 (N_7829,N_7442,N_7449);
nand U7830 (N_7830,N_7210,N_7104);
nor U7831 (N_7831,N_7094,N_7322);
and U7832 (N_7832,N_7376,N_7428);
nor U7833 (N_7833,N_7319,N_7356);
or U7834 (N_7834,N_7476,N_6900);
nand U7835 (N_7835,N_7134,N_6963);
nor U7836 (N_7836,N_7168,N_7115);
nand U7837 (N_7837,N_7365,N_7458);
or U7838 (N_7838,N_6770,N_7099);
nand U7839 (N_7839,N_7062,N_7303);
or U7840 (N_7840,N_7482,N_6905);
or U7841 (N_7841,N_7012,N_7185);
nand U7842 (N_7842,N_6952,N_7265);
nand U7843 (N_7843,N_7474,N_7043);
nor U7844 (N_7844,N_7199,N_7082);
or U7845 (N_7845,N_7027,N_7020);
nor U7846 (N_7846,N_7478,N_6834);
nand U7847 (N_7847,N_7407,N_6937);
nand U7848 (N_7848,N_7195,N_6898);
or U7849 (N_7849,N_7443,N_6895);
or U7850 (N_7850,N_7181,N_7239);
nand U7851 (N_7851,N_7351,N_7456);
and U7852 (N_7852,N_7044,N_7439);
nand U7853 (N_7853,N_6787,N_7136);
or U7854 (N_7854,N_6860,N_7457);
nand U7855 (N_7855,N_7035,N_7461);
nor U7856 (N_7856,N_7218,N_6922);
and U7857 (N_7857,N_7228,N_6978);
nor U7858 (N_7858,N_6791,N_6845);
or U7859 (N_7859,N_6915,N_7424);
or U7860 (N_7860,N_7261,N_6889);
xor U7861 (N_7861,N_7200,N_7180);
or U7862 (N_7862,N_7390,N_6764);
or U7863 (N_7863,N_6823,N_7470);
and U7864 (N_7864,N_6821,N_6782);
nor U7865 (N_7865,N_6798,N_6955);
or U7866 (N_7866,N_7302,N_6980);
and U7867 (N_7867,N_6835,N_6794);
nor U7868 (N_7868,N_7038,N_7292);
nor U7869 (N_7869,N_7431,N_6957);
or U7870 (N_7870,N_7280,N_7198);
nor U7871 (N_7871,N_7382,N_6877);
nor U7872 (N_7872,N_7149,N_7273);
nand U7873 (N_7873,N_7013,N_6974);
and U7874 (N_7874,N_7452,N_6771);
xor U7875 (N_7875,N_7344,N_7357);
nand U7876 (N_7876,N_6888,N_6896);
xor U7877 (N_7877,N_7142,N_7222);
and U7878 (N_7878,N_7301,N_7208);
nor U7879 (N_7879,N_6865,N_7080);
nand U7880 (N_7880,N_6874,N_7351);
nand U7881 (N_7881,N_7459,N_7471);
nand U7882 (N_7882,N_7089,N_7365);
nor U7883 (N_7883,N_7161,N_7491);
xnor U7884 (N_7884,N_6981,N_6870);
nand U7885 (N_7885,N_6951,N_6798);
and U7886 (N_7886,N_6988,N_7213);
nor U7887 (N_7887,N_6867,N_6988);
nand U7888 (N_7888,N_7441,N_7031);
xor U7889 (N_7889,N_7477,N_6835);
and U7890 (N_7890,N_7285,N_6858);
nor U7891 (N_7891,N_7126,N_7252);
nor U7892 (N_7892,N_6769,N_7470);
nand U7893 (N_7893,N_7410,N_7400);
or U7894 (N_7894,N_7319,N_6989);
nor U7895 (N_7895,N_7072,N_6832);
nand U7896 (N_7896,N_7263,N_7368);
nand U7897 (N_7897,N_7110,N_7393);
and U7898 (N_7898,N_7068,N_6839);
nand U7899 (N_7899,N_7049,N_7250);
or U7900 (N_7900,N_7267,N_7074);
nor U7901 (N_7901,N_7407,N_7200);
nand U7902 (N_7902,N_7098,N_6919);
nand U7903 (N_7903,N_7078,N_7499);
nand U7904 (N_7904,N_6807,N_7478);
xnor U7905 (N_7905,N_7136,N_7195);
or U7906 (N_7906,N_6974,N_7392);
nand U7907 (N_7907,N_6769,N_7348);
nand U7908 (N_7908,N_7050,N_7418);
nand U7909 (N_7909,N_6915,N_7079);
nor U7910 (N_7910,N_7016,N_7419);
nand U7911 (N_7911,N_6887,N_6944);
or U7912 (N_7912,N_6867,N_7396);
or U7913 (N_7913,N_7201,N_6942);
nand U7914 (N_7914,N_6879,N_7125);
nor U7915 (N_7915,N_7016,N_7112);
nand U7916 (N_7916,N_7473,N_7088);
nor U7917 (N_7917,N_6935,N_6781);
nor U7918 (N_7918,N_7123,N_7016);
or U7919 (N_7919,N_6999,N_6887);
nand U7920 (N_7920,N_7151,N_7079);
nand U7921 (N_7921,N_7102,N_7261);
and U7922 (N_7922,N_6755,N_7487);
and U7923 (N_7923,N_7434,N_6906);
nand U7924 (N_7924,N_6874,N_7028);
and U7925 (N_7925,N_7055,N_6790);
and U7926 (N_7926,N_7134,N_7264);
nor U7927 (N_7927,N_7043,N_7427);
xor U7928 (N_7928,N_7324,N_7097);
or U7929 (N_7929,N_6999,N_7000);
and U7930 (N_7930,N_6899,N_7274);
and U7931 (N_7931,N_7125,N_6854);
nand U7932 (N_7932,N_7190,N_7313);
nand U7933 (N_7933,N_6780,N_6993);
nand U7934 (N_7934,N_7076,N_6985);
nor U7935 (N_7935,N_7041,N_7396);
nor U7936 (N_7936,N_6912,N_7405);
nor U7937 (N_7937,N_7244,N_7282);
and U7938 (N_7938,N_7461,N_6830);
nand U7939 (N_7939,N_7261,N_7429);
and U7940 (N_7940,N_7292,N_7265);
and U7941 (N_7941,N_6953,N_7111);
nand U7942 (N_7942,N_7232,N_7380);
or U7943 (N_7943,N_7306,N_7011);
or U7944 (N_7944,N_7121,N_6955);
xor U7945 (N_7945,N_6778,N_6984);
or U7946 (N_7946,N_7005,N_6880);
and U7947 (N_7947,N_7495,N_7393);
or U7948 (N_7948,N_7223,N_7099);
nand U7949 (N_7949,N_7177,N_7036);
nor U7950 (N_7950,N_7406,N_6960);
or U7951 (N_7951,N_7363,N_7081);
or U7952 (N_7952,N_7128,N_6887);
and U7953 (N_7953,N_6782,N_6928);
nor U7954 (N_7954,N_7499,N_7468);
or U7955 (N_7955,N_6866,N_7169);
or U7956 (N_7956,N_6876,N_6857);
nor U7957 (N_7957,N_6805,N_6990);
nand U7958 (N_7958,N_6962,N_6814);
nand U7959 (N_7959,N_7080,N_7264);
nand U7960 (N_7960,N_6808,N_6885);
nor U7961 (N_7961,N_7238,N_7269);
xnor U7962 (N_7962,N_7024,N_6885);
nand U7963 (N_7963,N_7094,N_7246);
and U7964 (N_7964,N_6966,N_7133);
nand U7965 (N_7965,N_6854,N_7026);
and U7966 (N_7966,N_7177,N_7059);
xnor U7967 (N_7967,N_6899,N_6929);
nor U7968 (N_7968,N_7182,N_6962);
and U7969 (N_7969,N_7069,N_6830);
and U7970 (N_7970,N_7151,N_6873);
nand U7971 (N_7971,N_6825,N_6762);
nor U7972 (N_7972,N_7038,N_6910);
nand U7973 (N_7973,N_7020,N_7187);
nor U7974 (N_7974,N_7242,N_7011);
nand U7975 (N_7975,N_7002,N_7227);
nor U7976 (N_7976,N_7021,N_6998);
or U7977 (N_7977,N_7226,N_7360);
or U7978 (N_7978,N_6876,N_7213);
and U7979 (N_7979,N_7169,N_7405);
and U7980 (N_7980,N_7112,N_7248);
nand U7981 (N_7981,N_7069,N_7276);
nor U7982 (N_7982,N_6788,N_6787);
nor U7983 (N_7983,N_7083,N_7393);
nand U7984 (N_7984,N_7122,N_7332);
or U7985 (N_7985,N_6838,N_6796);
nand U7986 (N_7986,N_7054,N_7073);
xor U7987 (N_7987,N_7127,N_7118);
nor U7988 (N_7988,N_7193,N_7293);
nor U7989 (N_7989,N_6878,N_6773);
and U7990 (N_7990,N_6760,N_7048);
nand U7991 (N_7991,N_6866,N_7232);
xor U7992 (N_7992,N_6807,N_6843);
and U7993 (N_7993,N_7075,N_7389);
xnor U7994 (N_7994,N_6811,N_7136);
nand U7995 (N_7995,N_6986,N_6924);
nand U7996 (N_7996,N_7089,N_6764);
nor U7997 (N_7997,N_7053,N_7320);
or U7998 (N_7998,N_6950,N_6909);
or U7999 (N_7999,N_7352,N_6927);
or U8000 (N_8000,N_6889,N_7393);
or U8001 (N_8001,N_7048,N_7369);
and U8002 (N_8002,N_7261,N_7106);
and U8003 (N_8003,N_6766,N_6840);
or U8004 (N_8004,N_6864,N_6916);
nand U8005 (N_8005,N_6846,N_7028);
and U8006 (N_8006,N_7264,N_7394);
nand U8007 (N_8007,N_7246,N_7329);
and U8008 (N_8008,N_6873,N_7177);
xor U8009 (N_8009,N_7259,N_7332);
xnor U8010 (N_8010,N_6821,N_6767);
or U8011 (N_8011,N_7425,N_7344);
xor U8012 (N_8012,N_7124,N_7435);
nand U8013 (N_8013,N_6855,N_6931);
or U8014 (N_8014,N_7452,N_7074);
and U8015 (N_8015,N_7304,N_7377);
or U8016 (N_8016,N_7080,N_6760);
and U8017 (N_8017,N_7459,N_7303);
xor U8018 (N_8018,N_7385,N_6908);
nand U8019 (N_8019,N_6908,N_7125);
nor U8020 (N_8020,N_6964,N_6919);
or U8021 (N_8021,N_6864,N_7123);
and U8022 (N_8022,N_7367,N_7337);
or U8023 (N_8023,N_6872,N_7363);
and U8024 (N_8024,N_6972,N_7221);
nand U8025 (N_8025,N_7292,N_7208);
nand U8026 (N_8026,N_6805,N_7085);
nand U8027 (N_8027,N_7023,N_7464);
nor U8028 (N_8028,N_6957,N_6816);
or U8029 (N_8029,N_7370,N_6963);
xnor U8030 (N_8030,N_7003,N_7006);
and U8031 (N_8031,N_6953,N_7202);
nor U8032 (N_8032,N_7172,N_7088);
and U8033 (N_8033,N_7331,N_6816);
nand U8034 (N_8034,N_7133,N_7187);
or U8035 (N_8035,N_7028,N_7428);
and U8036 (N_8036,N_6958,N_7336);
nor U8037 (N_8037,N_6892,N_7087);
or U8038 (N_8038,N_7060,N_6948);
and U8039 (N_8039,N_6828,N_6826);
nand U8040 (N_8040,N_7004,N_7385);
nor U8041 (N_8041,N_7065,N_6886);
and U8042 (N_8042,N_6805,N_7338);
nand U8043 (N_8043,N_6958,N_7174);
xnor U8044 (N_8044,N_7272,N_7164);
xor U8045 (N_8045,N_7294,N_6853);
and U8046 (N_8046,N_7472,N_6756);
or U8047 (N_8047,N_7249,N_7050);
xnor U8048 (N_8048,N_6848,N_7215);
or U8049 (N_8049,N_7425,N_6881);
nor U8050 (N_8050,N_7323,N_7298);
nand U8051 (N_8051,N_7104,N_6936);
nand U8052 (N_8052,N_7338,N_6961);
nor U8053 (N_8053,N_6842,N_6849);
nor U8054 (N_8054,N_7258,N_7181);
or U8055 (N_8055,N_7226,N_6996);
nor U8056 (N_8056,N_7196,N_6913);
and U8057 (N_8057,N_7339,N_7171);
nor U8058 (N_8058,N_7013,N_7079);
nor U8059 (N_8059,N_7229,N_6850);
or U8060 (N_8060,N_6762,N_7414);
or U8061 (N_8061,N_7276,N_7029);
or U8062 (N_8062,N_7184,N_7447);
nand U8063 (N_8063,N_7052,N_6926);
nand U8064 (N_8064,N_7344,N_6936);
nor U8065 (N_8065,N_6892,N_7467);
and U8066 (N_8066,N_6948,N_7494);
nand U8067 (N_8067,N_7225,N_6759);
and U8068 (N_8068,N_7381,N_7308);
or U8069 (N_8069,N_6865,N_7428);
nand U8070 (N_8070,N_7123,N_7222);
nor U8071 (N_8071,N_6963,N_7442);
xnor U8072 (N_8072,N_7058,N_6920);
and U8073 (N_8073,N_6989,N_6770);
and U8074 (N_8074,N_7222,N_7389);
and U8075 (N_8075,N_6875,N_7322);
or U8076 (N_8076,N_6906,N_7036);
or U8077 (N_8077,N_7398,N_7000);
nand U8078 (N_8078,N_6777,N_6984);
nor U8079 (N_8079,N_7192,N_7183);
or U8080 (N_8080,N_7071,N_6801);
nor U8081 (N_8081,N_6767,N_7334);
and U8082 (N_8082,N_7276,N_7161);
or U8083 (N_8083,N_6777,N_7397);
nor U8084 (N_8084,N_6914,N_7150);
nand U8085 (N_8085,N_7043,N_7196);
nor U8086 (N_8086,N_7408,N_7073);
nor U8087 (N_8087,N_7151,N_6782);
nor U8088 (N_8088,N_7135,N_7329);
nor U8089 (N_8089,N_7227,N_6755);
nor U8090 (N_8090,N_6783,N_6750);
nor U8091 (N_8091,N_6966,N_6939);
or U8092 (N_8092,N_6900,N_7223);
nor U8093 (N_8093,N_7036,N_7173);
nor U8094 (N_8094,N_7475,N_7067);
xnor U8095 (N_8095,N_6855,N_6866);
xnor U8096 (N_8096,N_7385,N_7438);
and U8097 (N_8097,N_7245,N_7342);
xor U8098 (N_8098,N_7237,N_7153);
nand U8099 (N_8099,N_7178,N_7487);
or U8100 (N_8100,N_7282,N_7034);
xnor U8101 (N_8101,N_7320,N_7419);
and U8102 (N_8102,N_6900,N_7243);
or U8103 (N_8103,N_6920,N_6963);
or U8104 (N_8104,N_7119,N_7067);
nand U8105 (N_8105,N_6813,N_7047);
nand U8106 (N_8106,N_7411,N_7375);
nand U8107 (N_8107,N_7230,N_6807);
nor U8108 (N_8108,N_6880,N_7387);
nor U8109 (N_8109,N_7404,N_6873);
nor U8110 (N_8110,N_7388,N_7010);
nand U8111 (N_8111,N_6985,N_7092);
or U8112 (N_8112,N_7196,N_7328);
and U8113 (N_8113,N_7448,N_7265);
or U8114 (N_8114,N_7377,N_6824);
or U8115 (N_8115,N_7081,N_7406);
or U8116 (N_8116,N_7487,N_6867);
xnor U8117 (N_8117,N_7402,N_7228);
nor U8118 (N_8118,N_7428,N_7153);
nor U8119 (N_8119,N_7313,N_7297);
and U8120 (N_8120,N_7397,N_7027);
and U8121 (N_8121,N_7319,N_7084);
nand U8122 (N_8122,N_7231,N_6896);
nor U8123 (N_8123,N_7340,N_6955);
or U8124 (N_8124,N_7387,N_7271);
or U8125 (N_8125,N_6811,N_7145);
xor U8126 (N_8126,N_6874,N_7369);
nor U8127 (N_8127,N_7233,N_7376);
xnor U8128 (N_8128,N_7175,N_7124);
xor U8129 (N_8129,N_6798,N_7046);
nor U8130 (N_8130,N_6999,N_7070);
or U8131 (N_8131,N_7090,N_7488);
or U8132 (N_8132,N_6980,N_7092);
nor U8133 (N_8133,N_7237,N_7054);
or U8134 (N_8134,N_7183,N_7455);
or U8135 (N_8135,N_7376,N_6879);
and U8136 (N_8136,N_7430,N_7101);
xor U8137 (N_8137,N_7222,N_6792);
nor U8138 (N_8138,N_7407,N_7001);
xor U8139 (N_8139,N_7176,N_7110);
xnor U8140 (N_8140,N_7085,N_7432);
or U8141 (N_8141,N_7288,N_7105);
and U8142 (N_8142,N_6781,N_7194);
nand U8143 (N_8143,N_7336,N_7384);
nor U8144 (N_8144,N_7033,N_7306);
nand U8145 (N_8145,N_7207,N_7241);
nor U8146 (N_8146,N_7247,N_7374);
or U8147 (N_8147,N_6824,N_7177);
xor U8148 (N_8148,N_7179,N_7477);
and U8149 (N_8149,N_7283,N_7048);
nor U8150 (N_8150,N_7495,N_7217);
or U8151 (N_8151,N_6882,N_6821);
or U8152 (N_8152,N_7411,N_6970);
and U8153 (N_8153,N_7077,N_7253);
nor U8154 (N_8154,N_7131,N_7084);
and U8155 (N_8155,N_7191,N_7357);
xor U8156 (N_8156,N_7103,N_6833);
and U8157 (N_8157,N_6769,N_6995);
nand U8158 (N_8158,N_7202,N_6905);
nor U8159 (N_8159,N_7151,N_7320);
nand U8160 (N_8160,N_7438,N_7019);
and U8161 (N_8161,N_7138,N_6934);
or U8162 (N_8162,N_6999,N_6859);
or U8163 (N_8163,N_7183,N_7118);
or U8164 (N_8164,N_6797,N_7056);
xor U8165 (N_8165,N_7345,N_6829);
or U8166 (N_8166,N_7123,N_6961);
nand U8167 (N_8167,N_6821,N_7380);
nand U8168 (N_8168,N_7019,N_6778);
nand U8169 (N_8169,N_7452,N_7101);
nor U8170 (N_8170,N_7072,N_7294);
or U8171 (N_8171,N_7370,N_6864);
nand U8172 (N_8172,N_7422,N_7047);
and U8173 (N_8173,N_7340,N_6968);
nand U8174 (N_8174,N_7451,N_7061);
and U8175 (N_8175,N_7267,N_7281);
xor U8176 (N_8176,N_7376,N_7336);
or U8177 (N_8177,N_6846,N_6949);
and U8178 (N_8178,N_7447,N_7130);
nand U8179 (N_8179,N_7191,N_7286);
or U8180 (N_8180,N_7068,N_7469);
or U8181 (N_8181,N_6892,N_6965);
xor U8182 (N_8182,N_7045,N_7488);
nor U8183 (N_8183,N_7177,N_7485);
and U8184 (N_8184,N_7201,N_6785);
nand U8185 (N_8185,N_7493,N_7009);
and U8186 (N_8186,N_7176,N_7295);
nand U8187 (N_8187,N_6851,N_7105);
or U8188 (N_8188,N_7244,N_6969);
nor U8189 (N_8189,N_7171,N_7344);
or U8190 (N_8190,N_7197,N_7349);
and U8191 (N_8191,N_7262,N_6961);
or U8192 (N_8192,N_7376,N_7100);
and U8193 (N_8193,N_7320,N_7077);
nor U8194 (N_8194,N_6924,N_6906);
and U8195 (N_8195,N_6929,N_6955);
and U8196 (N_8196,N_7465,N_7190);
nor U8197 (N_8197,N_6783,N_7466);
nand U8198 (N_8198,N_6792,N_6842);
nor U8199 (N_8199,N_6917,N_6976);
or U8200 (N_8200,N_6955,N_6886);
nand U8201 (N_8201,N_7429,N_7126);
nor U8202 (N_8202,N_7405,N_7453);
and U8203 (N_8203,N_6922,N_7010);
nand U8204 (N_8204,N_6941,N_6961);
nor U8205 (N_8205,N_7137,N_7490);
nor U8206 (N_8206,N_7222,N_6880);
nor U8207 (N_8207,N_6969,N_7325);
nand U8208 (N_8208,N_7172,N_7442);
nor U8209 (N_8209,N_7240,N_7085);
nand U8210 (N_8210,N_6867,N_6926);
nand U8211 (N_8211,N_6791,N_7492);
nand U8212 (N_8212,N_7298,N_7401);
and U8213 (N_8213,N_7308,N_6802);
nor U8214 (N_8214,N_7435,N_7352);
and U8215 (N_8215,N_7022,N_6852);
xor U8216 (N_8216,N_7217,N_7146);
or U8217 (N_8217,N_7402,N_7411);
nand U8218 (N_8218,N_7170,N_7079);
or U8219 (N_8219,N_6807,N_7257);
or U8220 (N_8220,N_6985,N_6931);
nand U8221 (N_8221,N_7366,N_6886);
nand U8222 (N_8222,N_6937,N_7472);
and U8223 (N_8223,N_7059,N_7254);
xor U8224 (N_8224,N_7451,N_7333);
and U8225 (N_8225,N_7421,N_6821);
nand U8226 (N_8226,N_7004,N_6856);
or U8227 (N_8227,N_7348,N_7483);
or U8228 (N_8228,N_6981,N_6993);
nand U8229 (N_8229,N_7035,N_7150);
and U8230 (N_8230,N_7222,N_7301);
xor U8231 (N_8231,N_6969,N_6790);
or U8232 (N_8232,N_7231,N_6901);
and U8233 (N_8233,N_6879,N_6805);
nor U8234 (N_8234,N_7365,N_7407);
nand U8235 (N_8235,N_7399,N_7400);
and U8236 (N_8236,N_6906,N_7185);
or U8237 (N_8237,N_7018,N_7070);
nor U8238 (N_8238,N_7372,N_7446);
and U8239 (N_8239,N_7347,N_7409);
nand U8240 (N_8240,N_6755,N_6751);
or U8241 (N_8241,N_7489,N_7225);
xnor U8242 (N_8242,N_7252,N_6818);
nor U8243 (N_8243,N_7376,N_7364);
or U8244 (N_8244,N_7398,N_6954);
nand U8245 (N_8245,N_7165,N_7022);
or U8246 (N_8246,N_6857,N_7081);
nor U8247 (N_8247,N_7016,N_7001);
nand U8248 (N_8248,N_7119,N_7428);
nor U8249 (N_8249,N_6885,N_6836);
or U8250 (N_8250,N_7577,N_8176);
or U8251 (N_8251,N_8110,N_7813);
or U8252 (N_8252,N_7527,N_7573);
nor U8253 (N_8253,N_8213,N_7558);
nand U8254 (N_8254,N_8190,N_8015);
nor U8255 (N_8255,N_7729,N_7509);
and U8256 (N_8256,N_7682,N_8023);
or U8257 (N_8257,N_7924,N_7738);
or U8258 (N_8258,N_7585,N_8118);
and U8259 (N_8259,N_8131,N_7828);
or U8260 (N_8260,N_7647,N_7545);
or U8261 (N_8261,N_7854,N_8019);
nor U8262 (N_8262,N_7563,N_7718);
and U8263 (N_8263,N_7930,N_7763);
nand U8264 (N_8264,N_7945,N_7588);
nor U8265 (N_8265,N_7601,N_7700);
or U8266 (N_8266,N_8055,N_7937);
nand U8267 (N_8267,N_7923,N_8100);
and U8268 (N_8268,N_7826,N_8101);
and U8269 (N_8269,N_7799,N_8107);
and U8270 (N_8270,N_7995,N_8200);
or U8271 (N_8271,N_8060,N_8067);
or U8272 (N_8272,N_8208,N_7954);
nor U8273 (N_8273,N_7801,N_8069);
and U8274 (N_8274,N_7731,N_7872);
or U8275 (N_8275,N_7766,N_7897);
nor U8276 (N_8276,N_8004,N_7946);
and U8277 (N_8277,N_8172,N_7633);
or U8278 (N_8278,N_8127,N_7637);
nor U8279 (N_8279,N_7720,N_7947);
xor U8280 (N_8280,N_7579,N_7753);
nor U8281 (N_8281,N_7908,N_7519);
nor U8282 (N_8282,N_7940,N_7506);
nor U8283 (N_8283,N_8044,N_7961);
and U8284 (N_8284,N_8036,N_8026);
nor U8285 (N_8285,N_7734,N_7727);
nand U8286 (N_8286,N_7655,N_7638);
and U8287 (N_8287,N_8216,N_8064);
and U8288 (N_8288,N_8141,N_7709);
or U8289 (N_8289,N_7663,N_7909);
xnor U8290 (N_8290,N_8116,N_7855);
or U8291 (N_8291,N_8046,N_8109);
nor U8292 (N_8292,N_7825,N_7675);
nand U8293 (N_8293,N_7848,N_7530);
and U8294 (N_8294,N_7815,N_7783);
or U8295 (N_8295,N_8159,N_8029);
and U8296 (N_8296,N_7651,N_8105);
nor U8297 (N_8297,N_7972,N_7504);
nand U8298 (N_8298,N_8091,N_8011);
nor U8299 (N_8299,N_7806,N_7704);
or U8300 (N_8300,N_8113,N_7887);
or U8301 (N_8301,N_7640,N_8152);
and U8302 (N_8302,N_7877,N_8228);
and U8303 (N_8303,N_8084,N_8231);
and U8304 (N_8304,N_8239,N_8167);
or U8305 (N_8305,N_7911,N_8128);
or U8306 (N_8306,N_8016,N_7621);
xor U8307 (N_8307,N_7793,N_8063);
or U8308 (N_8308,N_7672,N_8214);
nand U8309 (N_8309,N_7539,N_7643);
or U8310 (N_8310,N_7988,N_7730);
nor U8311 (N_8311,N_7619,N_7798);
and U8312 (N_8312,N_7782,N_8248);
xnor U8313 (N_8313,N_8013,N_8197);
nand U8314 (N_8314,N_8042,N_7523);
and U8315 (N_8315,N_7977,N_7863);
nand U8316 (N_8316,N_7615,N_8249);
or U8317 (N_8317,N_8145,N_7892);
and U8318 (N_8318,N_7822,N_7610);
nand U8319 (N_8319,N_8170,N_7938);
or U8320 (N_8320,N_7850,N_7844);
nor U8321 (N_8321,N_7642,N_7973);
xnor U8322 (N_8322,N_7790,N_7811);
and U8323 (N_8323,N_7944,N_7900);
nand U8324 (N_8324,N_7551,N_7928);
and U8325 (N_8325,N_7553,N_7906);
xnor U8326 (N_8326,N_7745,N_8202);
or U8327 (N_8327,N_7544,N_7914);
or U8328 (N_8328,N_8028,N_7569);
or U8329 (N_8329,N_8241,N_8086);
nor U8330 (N_8330,N_8182,N_7732);
nand U8331 (N_8331,N_8125,N_7706);
and U8332 (N_8332,N_7598,N_7980);
or U8333 (N_8333,N_7968,N_7578);
nor U8334 (N_8334,N_8057,N_7823);
nand U8335 (N_8335,N_7883,N_8187);
or U8336 (N_8336,N_8094,N_7963);
and U8337 (N_8337,N_7628,N_7991);
nor U8338 (N_8338,N_8051,N_7532);
nand U8339 (N_8339,N_7915,N_7624);
nand U8340 (N_8340,N_7547,N_8092);
nand U8341 (N_8341,N_7531,N_8149);
and U8342 (N_8342,N_7969,N_7711);
nor U8343 (N_8343,N_7645,N_7723);
nor U8344 (N_8344,N_8158,N_7713);
xor U8345 (N_8345,N_7676,N_7851);
nor U8346 (N_8346,N_7744,N_7629);
xor U8347 (N_8347,N_7809,N_8181);
and U8348 (N_8348,N_8203,N_8043);
and U8349 (N_8349,N_7784,N_7989);
or U8350 (N_8350,N_7599,N_7898);
or U8351 (N_8351,N_7652,N_7757);
nand U8352 (N_8352,N_8192,N_8186);
and U8353 (N_8353,N_7550,N_8102);
nor U8354 (N_8354,N_7534,N_7587);
or U8355 (N_8355,N_7749,N_7511);
nor U8356 (N_8356,N_7702,N_7746);
nand U8357 (N_8357,N_7717,N_8243);
nor U8358 (N_8358,N_7699,N_8196);
nand U8359 (N_8359,N_7879,N_7810);
and U8360 (N_8360,N_8169,N_7696);
nand U8361 (N_8361,N_7878,N_7916);
or U8362 (N_8362,N_8089,N_7679);
nor U8363 (N_8363,N_7522,N_7688);
or U8364 (N_8364,N_7756,N_7864);
nand U8365 (N_8365,N_7773,N_7904);
xnor U8366 (N_8366,N_7510,N_8142);
or U8367 (N_8367,N_7890,N_8073);
nand U8368 (N_8368,N_7901,N_7902);
nand U8369 (N_8369,N_8061,N_7839);
or U8370 (N_8370,N_7994,N_7866);
nand U8371 (N_8371,N_8088,N_7568);
or U8372 (N_8372,N_7592,N_8065);
and U8373 (N_8373,N_7987,N_8081);
nor U8374 (N_8374,N_7816,N_7646);
nand U8375 (N_8375,N_7570,N_7760);
nor U8376 (N_8376,N_7884,N_7767);
and U8377 (N_8377,N_7525,N_7979);
nand U8378 (N_8378,N_7836,N_7574);
or U8379 (N_8379,N_7657,N_7934);
and U8380 (N_8380,N_7808,N_7779);
nor U8381 (N_8381,N_7742,N_8133);
or U8382 (N_8382,N_7800,N_7674);
xor U8383 (N_8383,N_7540,N_7858);
nor U8384 (N_8384,N_7956,N_8221);
nand U8385 (N_8385,N_8047,N_7560);
and U8386 (N_8386,N_7649,N_7626);
xnor U8387 (N_8387,N_7668,N_7935);
nor U8388 (N_8388,N_8104,N_7978);
or U8389 (N_8389,N_7516,N_7778);
nand U8390 (N_8390,N_7833,N_8175);
and U8391 (N_8391,N_7796,N_7533);
nand U8392 (N_8392,N_8123,N_7758);
or U8393 (N_8393,N_7959,N_8112);
and U8394 (N_8394,N_7976,N_8097);
and U8395 (N_8395,N_7571,N_7993);
nand U8396 (N_8396,N_8166,N_8022);
nor U8397 (N_8397,N_7941,N_7561);
nor U8398 (N_8398,N_7794,N_7875);
nor U8399 (N_8399,N_7590,N_8179);
nand U8400 (N_8400,N_7919,N_7846);
or U8401 (N_8401,N_7543,N_7518);
nor U8402 (N_8402,N_8134,N_7564);
nand U8403 (N_8403,N_8234,N_8014);
xor U8404 (N_8404,N_8005,N_7802);
xnor U8405 (N_8405,N_7733,N_7538);
nor U8406 (N_8406,N_7960,N_7695);
nand U8407 (N_8407,N_8080,N_8189);
nor U8408 (N_8408,N_7614,N_7775);
nand U8409 (N_8409,N_7716,N_7606);
and U8410 (N_8410,N_7739,N_8072);
or U8411 (N_8411,N_8074,N_7831);
and U8412 (N_8412,N_7684,N_7780);
nand U8413 (N_8413,N_7774,N_8225);
or U8414 (N_8414,N_7754,N_7891);
nor U8415 (N_8415,N_7795,N_7894);
nand U8416 (N_8416,N_7992,N_7971);
or U8417 (N_8417,N_8178,N_7697);
and U8418 (N_8418,N_8068,N_7520);
or U8419 (N_8419,N_7881,N_8098);
or U8420 (N_8420,N_7671,N_7936);
nor U8421 (N_8421,N_7514,N_7627);
nor U8422 (N_8422,N_8229,N_7701);
or U8423 (N_8423,N_7762,N_7860);
xor U8424 (N_8424,N_7604,N_7631);
nand U8425 (N_8425,N_7933,N_7899);
or U8426 (N_8426,N_7726,N_7841);
nor U8427 (N_8427,N_7951,N_7820);
or U8428 (N_8428,N_7856,N_7721);
or U8429 (N_8429,N_8010,N_7677);
nand U8430 (N_8430,N_8050,N_7670);
and U8431 (N_8431,N_7786,N_7982);
nor U8432 (N_8432,N_7903,N_8174);
and U8433 (N_8433,N_7787,N_8244);
or U8434 (N_8434,N_8139,N_8168);
nand U8435 (N_8435,N_8210,N_7886);
nand U8436 (N_8436,N_8031,N_7715);
xor U8437 (N_8437,N_7608,N_7920);
nand U8438 (N_8438,N_7931,N_7876);
xor U8439 (N_8439,N_7835,N_7748);
nor U8440 (N_8440,N_8218,N_8012);
or U8441 (N_8441,N_8034,N_7750);
nor U8442 (N_8442,N_7683,N_8121);
nor U8443 (N_8443,N_8151,N_7803);
nand U8444 (N_8444,N_8135,N_7636);
or U8445 (N_8445,N_7949,N_8245);
and U8446 (N_8446,N_8160,N_7535);
and U8447 (N_8447,N_7542,N_8230);
nand U8448 (N_8448,N_7764,N_8070);
nor U8449 (N_8449,N_8240,N_7623);
or U8450 (N_8450,N_8129,N_7586);
xnor U8451 (N_8451,N_7869,N_8079);
or U8452 (N_8452,N_7515,N_8163);
nor U8453 (N_8453,N_7567,N_8157);
nor U8454 (N_8454,N_8093,N_8017);
or U8455 (N_8455,N_8191,N_7616);
or U8456 (N_8456,N_7965,N_7710);
and U8457 (N_8457,N_7747,N_7639);
and U8458 (N_8458,N_8085,N_8209);
and U8459 (N_8459,N_7691,N_8008);
nand U8460 (N_8460,N_8066,N_8148);
or U8461 (N_8461,N_7630,N_8075);
nand U8462 (N_8462,N_7537,N_7611);
xnor U8463 (N_8463,N_8171,N_7557);
xor U8464 (N_8464,N_7929,N_7501);
and U8465 (N_8465,N_7853,N_7932);
or U8466 (N_8466,N_8111,N_8122);
nand U8467 (N_8467,N_8155,N_7913);
or U8468 (N_8468,N_8201,N_7505);
nor U8469 (N_8469,N_7594,N_7583);
and U8470 (N_8470,N_7528,N_7885);
or U8471 (N_8471,N_8217,N_7521);
or U8472 (N_8472,N_7759,N_7591);
nor U8473 (N_8473,N_7999,N_7769);
and U8474 (N_8474,N_7680,N_7857);
nand U8475 (N_8475,N_7985,N_7781);
and U8476 (N_8476,N_7832,N_7953);
or U8477 (N_8477,N_8049,N_8082);
and U8478 (N_8478,N_7653,N_8052);
and U8479 (N_8479,N_8180,N_8238);
and U8480 (N_8480,N_7882,N_7895);
or U8481 (N_8481,N_8144,N_7830);
or U8482 (N_8482,N_7740,N_8237);
and U8483 (N_8483,N_8056,N_8184);
or U8484 (N_8484,N_8242,N_8039);
or U8485 (N_8485,N_8233,N_7658);
and U8486 (N_8486,N_8126,N_7925);
nor U8487 (N_8487,N_8103,N_7659);
nor U8488 (N_8488,N_7641,N_7580);
nand U8489 (N_8489,N_7548,N_8037);
xnor U8490 (N_8490,N_7772,N_7785);
nand U8491 (N_8491,N_7613,N_8194);
xor U8492 (N_8492,N_8173,N_7595);
or U8493 (N_8493,N_7536,N_7554);
and U8494 (N_8494,N_7765,N_7955);
xor U8495 (N_8495,N_7681,N_7603);
or U8496 (N_8496,N_7893,N_8223);
or U8497 (N_8497,N_7958,N_7998);
and U8498 (N_8498,N_7669,N_7689);
or U8499 (N_8499,N_7654,N_7950);
and U8500 (N_8500,N_7888,N_7735);
or U8501 (N_8501,N_8143,N_7634);
nand U8502 (N_8502,N_8120,N_7792);
nor U8503 (N_8503,N_7562,N_7648);
nand U8504 (N_8504,N_7566,N_7970);
or U8505 (N_8505,N_7698,N_8235);
nor U8506 (N_8506,N_7865,N_7752);
and U8507 (N_8507,N_7797,N_7849);
nand U8508 (N_8508,N_7771,N_7687);
or U8509 (N_8509,N_7556,N_7843);
xor U8510 (N_8510,N_8077,N_8040);
and U8511 (N_8511,N_7593,N_7804);
and U8512 (N_8512,N_7814,N_8027);
or U8513 (N_8513,N_8018,N_8021);
and U8514 (N_8514,N_8211,N_8124);
and U8515 (N_8515,N_7575,N_8002);
nor U8516 (N_8516,N_7708,N_8071);
or U8517 (N_8517,N_8222,N_8154);
or U8518 (N_8518,N_8032,N_8224);
nor U8519 (N_8519,N_8035,N_7777);
nand U8520 (N_8520,N_7724,N_7600);
nor U8521 (N_8521,N_8038,N_7705);
xnor U8522 (N_8522,N_8099,N_8076);
or U8523 (N_8523,N_8054,N_8045);
and U8524 (N_8524,N_7817,N_7905);
xor U8525 (N_8525,N_7555,N_8087);
nand U8526 (N_8526,N_7622,N_7807);
or U8527 (N_8527,N_7874,N_7620);
nor U8528 (N_8528,N_8236,N_7660);
or U8529 (N_8529,N_7662,N_8146);
nor U8530 (N_8530,N_7625,N_8185);
nor U8531 (N_8531,N_7819,N_7990);
nor U8532 (N_8532,N_8007,N_8137);
or U8533 (N_8533,N_8183,N_8205);
and U8534 (N_8534,N_8246,N_7728);
or U8535 (N_8535,N_8115,N_7829);
nor U8536 (N_8536,N_7840,N_8083);
nor U8537 (N_8537,N_7852,N_7939);
xor U8538 (N_8538,N_8193,N_7644);
or U8539 (N_8539,N_7859,N_7975);
nand U8540 (N_8540,N_7867,N_8132);
and U8541 (N_8541,N_8001,N_7719);
xor U8542 (N_8542,N_8095,N_8062);
xor U8543 (N_8543,N_8164,N_8108);
nand U8544 (N_8544,N_7943,N_7910);
nand U8545 (N_8545,N_7589,N_7983);
and U8546 (N_8546,N_8206,N_7690);
nor U8547 (N_8547,N_7948,N_7743);
xor U8548 (N_8548,N_7692,N_7552);
nor U8549 (N_8549,N_8215,N_7576);
and U8550 (N_8550,N_7707,N_7736);
and U8551 (N_8551,N_8058,N_8106);
and U8552 (N_8552,N_7596,N_7703);
nor U8553 (N_8553,N_7678,N_7693);
nand U8554 (N_8554,N_8247,N_7838);
xnor U8555 (N_8555,N_7612,N_7751);
and U8556 (N_8556,N_8207,N_7981);
xnor U8557 (N_8557,N_8226,N_7605);
xor U8558 (N_8558,N_7686,N_7529);
nor U8559 (N_8559,N_8220,N_8161);
nor U8560 (N_8560,N_8177,N_8212);
or U8561 (N_8561,N_7776,N_7962);
xor U8562 (N_8562,N_7837,N_7755);
or U8563 (N_8563,N_7650,N_7685);
or U8564 (N_8564,N_7673,N_7896);
and U8565 (N_8565,N_7952,N_7761);
nor U8566 (N_8566,N_7957,N_8096);
nor U8567 (N_8567,N_7805,N_7834);
nand U8568 (N_8568,N_7845,N_7712);
and U8569 (N_8569,N_7513,N_7526);
nor U8570 (N_8570,N_7821,N_7609);
nor U8571 (N_8571,N_7912,N_7559);
and U8572 (N_8572,N_8219,N_7665);
nand U8573 (N_8573,N_7635,N_7788);
nand U8574 (N_8574,N_7602,N_7926);
xor U8575 (N_8575,N_7927,N_7964);
xor U8576 (N_8576,N_7607,N_7597);
nor U8577 (N_8577,N_8059,N_7984);
or U8578 (N_8578,N_7541,N_8138);
xnor U8579 (N_8579,N_7812,N_7870);
nor U8580 (N_8580,N_7921,N_8020);
nand U8581 (N_8581,N_7789,N_7986);
or U8582 (N_8582,N_7827,N_7996);
and U8583 (N_8583,N_7880,N_8114);
nand U8584 (N_8584,N_7791,N_7967);
nor U8585 (N_8585,N_7664,N_8188);
and U8586 (N_8586,N_7502,N_8140);
and U8587 (N_8587,N_7889,N_7618);
or U8588 (N_8588,N_8009,N_7572);
nand U8589 (N_8589,N_7661,N_7966);
or U8590 (N_8590,N_7818,N_7517);
nor U8591 (N_8591,N_8195,N_7632);
xor U8592 (N_8592,N_7667,N_7584);
or U8593 (N_8593,N_7871,N_7768);
nand U8594 (N_8594,N_7524,N_7549);
nand U8595 (N_8595,N_8165,N_7997);
or U8596 (N_8596,N_7770,N_7873);
and U8597 (N_8597,N_8130,N_7714);
or U8598 (N_8598,N_7741,N_7508);
xor U8599 (N_8599,N_7861,N_7666);
xnor U8600 (N_8600,N_7847,N_7656);
xor U8601 (N_8601,N_7507,N_8153);
or U8602 (N_8602,N_8053,N_8162);
or U8603 (N_8603,N_7503,N_8006);
or U8604 (N_8604,N_8119,N_8227);
nand U8605 (N_8605,N_8204,N_8000);
and U8606 (N_8606,N_8078,N_8048);
xor U8607 (N_8607,N_7922,N_7500);
nor U8608 (N_8608,N_7942,N_7725);
nor U8609 (N_8609,N_7546,N_7582);
and U8610 (N_8610,N_7918,N_8117);
or U8611 (N_8611,N_7722,N_8147);
and U8612 (N_8612,N_8136,N_8025);
and U8613 (N_8613,N_7974,N_7737);
xor U8614 (N_8614,N_8090,N_7917);
and U8615 (N_8615,N_8024,N_7824);
and U8616 (N_8616,N_7617,N_8199);
nor U8617 (N_8617,N_8041,N_8150);
nand U8618 (N_8618,N_7842,N_7581);
nand U8619 (N_8619,N_7868,N_7907);
nor U8620 (N_8620,N_8030,N_7565);
nand U8621 (N_8621,N_7862,N_8198);
and U8622 (N_8622,N_8003,N_8156);
and U8623 (N_8623,N_7512,N_7694);
nor U8624 (N_8624,N_8232,N_8033);
or U8625 (N_8625,N_7535,N_7651);
and U8626 (N_8626,N_7715,N_8249);
and U8627 (N_8627,N_7956,N_8003);
or U8628 (N_8628,N_8103,N_7984);
and U8629 (N_8629,N_7998,N_7503);
nor U8630 (N_8630,N_7539,N_7725);
nand U8631 (N_8631,N_8205,N_8012);
nor U8632 (N_8632,N_7906,N_7904);
and U8633 (N_8633,N_8198,N_8116);
and U8634 (N_8634,N_7588,N_7522);
or U8635 (N_8635,N_7602,N_7604);
nor U8636 (N_8636,N_7957,N_7872);
or U8637 (N_8637,N_7919,N_8178);
and U8638 (N_8638,N_8157,N_8060);
or U8639 (N_8639,N_8217,N_7727);
and U8640 (N_8640,N_7770,N_8074);
xor U8641 (N_8641,N_8106,N_7685);
and U8642 (N_8642,N_7879,N_7593);
nand U8643 (N_8643,N_7595,N_7795);
nand U8644 (N_8644,N_7547,N_7535);
nand U8645 (N_8645,N_8023,N_8079);
or U8646 (N_8646,N_8100,N_8249);
or U8647 (N_8647,N_7919,N_7562);
nor U8648 (N_8648,N_7761,N_7630);
or U8649 (N_8649,N_7590,N_8153);
and U8650 (N_8650,N_7664,N_7769);
and U8651 (N_8651,N_7984,N_7956);
or U8652 (N_8652,N_7774,N_8053);
nor U8653 (N_8653,N_8079,N_7664);
nand U8654 (N_8654,N_8155,N_7574);
nand U8655 (N_8655,N_7626,N_7541);
nand U8656 (N_8656,N_8065,N_7645);
nand U8657 (N_8657,N_7747,N_7680);
xor U8658 (N_8658,N_8133,N_8029);
or U8659 (N_8659,N_8057,N_7564);
nand U8660 (N_8660,N_8098,N_7515);
nand U8661 (N_8661,N_7856,N_7998);
nand U8662 (N_8662,N_8204,N_8165);
nand U8663 (N_8663,N_7727,N_7543);
nor U8664 (N_8664,N_7743,N_7850);
nor U8665 (N_8665,N_7586,N_7935);
nand U8666 (N_8666,N_7571,N_7654);
or U8667 (N_8667,N_7777,N_7943);
nand U8668 (N_8668,N_7918,N_7787);
nand U8669 (N_8669,N_7601,N_7785);
and U8670 (N_8670,N_8073,N_7650);
or U8671 (N_8671,N_7723,N_7954);
and U8672 (N_8672,N_8075,N_8099);
or U8673 (N_8673,N_8068,N_8103);
nand U8674 (N_8674,N_8097,N_7541);
nand U8675 (N_8675,N_8106,N_7691);
xnor U8676 (N_8676,N_7660,N_7644);
and U8677 (N_8677,N_7697,N_8239);
and U8678 (N_8678,N_7824,N_7989);
nand U8679 (N_8679,N_8205,N_8030);
nor U8680 (N_8680,N_7775,N_7885);
xnor U8681 (N_8681,N_7817,N_7926);
nor U8682 (N_8682,N_7592,N_7873);
nand U8683 (N_8683,N_7700,N_8220);
nor U8684 (N_8684,N_7628,N_7578);
or U8685 (N_8685,N_7897,N_7536);
or U8686 (N_8686,N_8103,N_8110);
nor U8687 (N_8687,N_8194,N_7592);
nand U8688 (N_8688,N_8042,N_8120);
and U8689 (N_8689,N_8087,N_7686);
nand U8690 (N_8690,N_7916,N_7656);
or U8691 (N_8691,N_7899,N_7887);
nand U8692 (N_8692,N_7655,N_7772);
or U8693 (N_8693,N_8185,N_7863);
nor U8694 (N_8694,N_7811,N_8211);
and U8695 (N_8695,N_8187,N_7500);
nor U8696 (N_8696,N_7976,N_7707);
nand U8697 (N_8697,N_8175,N_7893);
and U8698 (N_8698,N_7548,N_7965);
or U8699 (N_8699,N_7700,N_8026);
nand U8700 (N_8700,N_7983,N_7765);
nand U8701 (N_8701,N_7987,N_8057);
nor U8702 (N_8702,N_8154,N_7937);
or U8703 (N_8703,N_8112,N_7911);
nand U8704 (N_8704,N_7517,N_8153);
and U8705 (N_8705,N_7804,N_7585);
or U8706 (N_8706,N_7611,N_7796);
nor U8707 (N_8707,N_8057,N_7567);
or U8708 (N_8708,N_8163,N_7985);
and U8709 (N_8709,N_7851,N_7655);
or U8710 (N_8710,N_8035,N_8022);
nand U8711 (N_8711,N_7954,N_7776);
nand U8712 (N_8712,N_8224,N_7804);
nor U8713 (N_8713,N_8153,N_7873);
nand U8714 (N_8714,N_7867,N_7721);
nor U8715 (N_8715,N_7583,N_7989);
xor U8716 (N_8716,N_8149,N_7691);
nand U8717 (N_8717,N_8099,N_8086);
xor U8718 (N_8718,N_7958,N_7733);
xor U8719 (N_8719,N_8049,N_7617);
and U8720 (N_8720,N_8096,N_7765);
or U8721 (N_8721,N_7859,N_8213);
or U8722 (N_8722,N_8137,N_7607);
nor U8723 (N_8723,N_8090,N_7923);
and U8724 (N_8724,N_7853,N_8017);
nor U8725 (N_8725,N_7786,N_7856);
and U8726 (N_8726,N_7673,N_7696);
or U8727 (N_8727,N_7687,N_7764);
or U8728 (N_8728,N_8038,N_7785);
nand U8729 (N_8729,N_7848,N_8064);
nand U8730 (N_8730,N_7760,N_7518);
and U8731 (N_8731,N_8120,N_7833);
nor U8732 (N_8732,N_8203,N_7525);
and U8733 (N_8733,N_7582,N_7504);
nand U8734 (N_8734,N_8078,N_7704);
nand U8735 (N_8735,N_7956,N_7810);
nand U8736 (N_8736,N_8062,N_7709);
and U8737 (N_8737,N_8218,N_7954);
and U8738 (N_8738,N_8188,N_8104);
nand U8739 (N_8739,N_7986,N_7990);
nand U8740 (N_8740,N_8242,N_7643);
nor U8741 (N_8741,N_7948,N_8181);
nand U8742 (N_8742,N_7654,N_7785);
or U8743 (N_8743,N_7793,N_7936);
nand U8744 (N_8744,N_8113,N_7657);
nand U8745 (N_8745,N_8112,N_7607);
nand U8746 (N_8746,N_7933,N_7602);
and U8747 (N_8747,N_7553,N_8160);
and U8748 (N_8748,N_7704,N_7826);
and U8749 (N_8749,N_8108,N_7581);
and U8750 (N_8750,N_7791,N_7890);
or U8751 (N_8751,N_7847,N_7962);
or U8752 (N_8752,N_7510,N_7818);
or U8753 (N_8753,N_7585,N_7798);
and U8754 (N_8754,N_7747,N_7595);
nor U8755 (N_8755,N_7628,N_7879);
nor U8756 (N_8756,N_7824,N_7932);
xnor U8757 (N_8757,N_7696,N_7695);
and U8758 (N_8758,N_7825,N_7535);
or U8759 (N_8759,N_8235,N_7652);
or U8760 (N_8760,N_7661,N_7596);
and U8761 (N_8761,N_7628,N_8030);
and U8762 (N_8762,N_7525,N_7976);
or U8763 (N_8763,N_7899,N_8093);
nand U8764 (N_8764,N_7689,N_7623);
or U8765 (N_8765,N_8065,N_7583);
or U8766 (N_8766,N_7956,N_8211);
xor U8767 (N_8767,N_7607,N_7551);
nor U8768 (N_8768,N_7760,N_7877);
or U8769 (N_8769,N_8074,N_8246);
and U8770 (N_8770,N_8192,N_7569);
xor U8771 (N_8771,N_8058,N_7952);
or U8772 (N_8772,N_8105,N_7567);
xor U8773 (N_8773,N_7660,N_7745);
and U8774 (N_8774,N_7954,N_7936);
nor U8775 (N_8775,N_8142,N_7852);
or U8776 (N_8776,N_8109,N_8157);
and U8777 (N_8777,N_8235,N_7961);
or U8778 (N_8778,N_7976,N_7855);
xor U8779 (N_8779,N_7684,N_7650);
or U8780 (N_8780,N_7897,N_7916);
or U8781 (N_8781,N_8210,N_7893);
nor U8782 (N_8782,N_8197,N_7547);
and U8783 (N_8783,N_8190,N_8217);
and U8784 (N_8784,N_7694,N_8240);
or U8785 (N_8785,N_8117,N_7900);
nor U8786 (N_8786,N_8111,N_7907);
nor U8787 (N_8787,N_7983,N_7699);
or U8788 (N_8788,N_7806,N_7803);
and U8789 (N_8789,N_7904,N_7661);
or U8790 (N_8790,N_7654,N_8233);
nand U8791 (N_8791,N_8038,N_8125);
and U8792 (N_8792,N_7635,N_8150);
nor U8793 (N_8793,N_8028,N_8081);
nand U8794 (N_8794,N_7515,N_7639);
nor U8795 (N_8795,N_7529,N_7717);
nand U8796 (N_8796,N_7767,N_7959);
nand U8797 (N_8797,N_7923,N_8018);
nand U8798 (N_8798,N_7696,N_7921);
and U8799 (N_8799,N_7781,N_8233);
nand U8800 (N_8800,N_7866,N_8200);
nand U8801 (N_8801,N_8080,N_7667);
and U8802 (N_8802,N_7583,N_8242);
or U8803 (N_8803,N_7882,N_8160);
and U8804 (N_8804,N_7574,N_7711);
xnor U8805 (N_8805,N_8143,N_7819);
and U8806 (N_8806,N_7915,N_7816);
and U8807 (N_8807,N_7968,N_8054);
and U8808 (N_8808,N_8114,N_7851);
nor U8809 (N_8809,N_7927,N_8243);
or U8810 (N_8810,N_7584,N_8139);
and U8811 (N_8811,N_8153,N_8249);
or U8812 (N_8812,N_7591,N_8033);
nor U8813 (N_8813,N_8218,N_7786);
and U8814 (N_8814,N_8080,N_8182);
and U8815 (N_8815,N_7905,N_7630);
and U8816 (N_8816,N_7658,N_7872);
xnor U8817 (N_8817,N_7690,N_7697);
nand U8818 (N_8818,N_7823,N_8134);
or U8819 (N_8819,N_7628,N_7998);
nor U8820 (N_8820,N_7626,N_7548);
nor U8821 (N_8821,N_7978,N_7756);
nor U8822 (N_8822,N_7632,N_7963);
and U8823 (N_8823,N_7708,N_7885);
and U8824 (N_8824,N_7647,N_7728);
and U8825 (N_8825,N_8230,N_8191);
nand U8826 (N_8826,N_8117,N_7747);
and U8827 (N_8827,N_8052,N_8058);
nor U8828 (N_8828,N_8184,N_8119);
and U8829 (N_8829,N_7903,N_8158);
or U8830 (N_8830,N_7819,N_8152);
nand U8831 (N_8831,N_7891,N_7989);
nand U8832 (N_8832,N_7894,N_8110);
nor U8833 (N_8833,N_8245,N_7600);
or U8834 (N_8834,N_8015,N_7522);
or U8835 (N_8835,N_7917,N_7879);
or U8836 (N_8836,N_7867,N_7946);
and U8837 (N_8837,N_8156,N_8113);
or U8838 (N_8838,N_8004,N_7559);
or U8839 (N_8839,N_7606,N_7686);
and U8840 (N_8840,N_7631,N_7507);
and U8841 (N_8841,N_8123,N_7716);
nor U8842 (N_8842,N_7518,N_8159);
nand U8843 (N_8843,N_7917,N_7849);
xnor U8844 (N_8844,N_7672,N_8217);
nor U8845 (N_8845,N_8215,N_7638);
or U8846 (N_8846,N_7958,N_7863);
nand U8847 (N_8847,N_8158,N_7926);
nor U8848 (N_8848,N_7952,N_8099);
xnor U8849 (N_8849,N_8074,N_7875);
and U8850 (N_8850,N_8199,N_7760);
and U8851 (N_8851,N_7720,N_8118);
or U8852 (N_8852,N_7878,N_8010);
and U8853 (N_8853,N_8025,N_7706);
xor U8854 (N_8854,N_8216,N_7607);
nand U8855 (N_8855,N_7534,N_7894);
nand U8856 (N_8856,N_7580,N_7920);
and U8857 (N_8857,N_7818,N_7644);
nor U8858 (N_8858,N_7980,N_7676);
nor U8859 (N_8859,N_7942,N_7698);
nand U8860 (N_8860,N_7517,N_8237);
or U8861 (N_8861,N_7778,N_8129);
xnor U8862 (N_8862,N_7518,N_7566);
nand U8863 (N_8863,N_8237,N_7743);
or U8864 (N_8864,N_7506,N_7954);
or U8865 (N_8865,N_7941,N_8117);
nand U8866 (N_8866,N_8247,N_8147);
xor U8867 (N_8867,N_8123,N_7928);
nand U8868 (N_8868,N_7741,N_7845);
nor U8869 (N_8869,N_7628,N_7632);
nor U8870 (N_8870,N_8227,N_7606);
xor U8871 (N_8871,N_7629,N_7586);
xor U8872 (N_8872,N_7982,N_7519);
nand U8873 (N_8873,N_8110,N_7754);
and U8874 (N_8874,N_8034,N_7923);
xor U8875 (N_8875,N_7866,N_7586);
nand U8876 (N_8876,N_8113,N_7782);
nor U8877 (N_8877,N_8215,N_7766);
nand U8878 (N_8878,N_7964,N_8057);
nor U8879 (N_8879,N_7797,N_7907);
nand U8880 (N_8880,N_7582,N_7622);
xor U8881 (N_8881,N_7663,N_8136);
nand U8882 (N_8882,N_7781,N_8164);
nor U8883 (N_8883,N_7733,N_7753);
or U8884 (N_8884,N_8158,N_7770);
nand U8885 (N_8885,N_7581,N_8243);
xnor U8886 (N_8886,N_7886,N_7977);
or U8887 (N_8887,N_7915,N_8123);
and U8888 (N_8888,N_8160,N_7974);
and U8889 (N_8889,N_8142,N_7888);
nor U8890 (N_8890,N_7798,N_7811);
or U8891 (N_8891,N_7984,N_7735);
or U8892 (N_8892,N_7747,N_7839);
or U8893 (N_8893,N_7803,N_8196);
nand U8894 (N_8894,N_7625,N_7735);
nand U8895 (N_8895,N_7828,N_8056);
and U8896 (N_8896,N_8097,N_7829);
nor U8897 (N_8897,N_8022,N_8038);
and U8898 (N_8898,N_7614,N_8150);
nor U8899 (N_8899,N_7513,N_8085);
and U8900 (N_8900,N_7541,N_7636);
nand U8901 (N_8901,N_7537,N_8165);
or U8902 (N_8902,N_7995,N_7779);
and U8903 (N_8903,N_8166,N_8062);
or U8904 (N_8904,N_8094,N_8015);
nand U8905 (N_8905,N_7739,N_8066);
and U8906 (N_8906,N_7878,N_8062);
nor U8907 (N_8907,N_7723,N_7815);
xor U8908 (N_8908,N_7613,N_7676);
nand U8909 (N_8909,N_8021,N_8189);
xor U8910 (N_8910,N_7998,N_8002);
nor U8911 (N_8911,N_7647,N_7823);
and U8912 (N_8912,N_8020,N_7679);
nand U8913 (N_8913,N_7991,N_7575);
or U8914 (N_8914,N_7901,N_7571);
or U8915 (N_8915,N_7973,N_8193);
and U8916 (N_8916,N_8227,N_8218);
and U8917 (N_8917,N_8019,N_7817);
or U8918 (N_8918,N_7667,N_7894);
or U8919 (N_8919,N_8170,N_7801);
or U8920 (N_8920,N_7815,N_8037);
nor U8921 (N_8921,N_7565,N_7543);
nand U8922 (N_8922,N_8067,N_8184);
nand U8923 (N_8923,N_7963,N_7822);
xnor U8924 (N_8924,N_7852,N_7672);
nor U8925 (N_8925,N_7932,N_8198);
and U8926 (N_8926,N_7799,N_7748);
and U8927 (N_8927,N_7515,N_8085);
nor U8928 (N_8928,N_7965,N_7903);
or U8929 (N_8929,N_8167,N_8172);
nor U8930 (N_8930,N_7987,N_7981);
xnor U8931 (N_8931,N_8044,N_7600);
and U8932 (N_8932,N_8186,N_7530);
nor U8933 (N_8933,N_7658,N_8146);
nand U8934 (N_8934,N_7688,N_7668);
and U8935 (N_8935,N_7822,N_8027);
and U8936 (N_8936,N_8092,N_7863);
xor U8937 (N_8937,N_8035,N_7706);
nand U8938 (N_8938,N_8010,N_7901);
nand U8939 (N_8939,N_8031,N_7866);
xnor U8940 (N_8940,N_8071,N_8009);
and U8941 (N_8941,N_7620,N_7860);
or U8942 (N_8942,N_7598,N_7638);
xor U8943 (N_8943,N_7687,N_7788);
xnor U8944 (N_8944,N_8064,N_8161);
nand U8945 (N_8945,N_7973,N_7936);
or U8946 (N_8946,N_7677,N_7581);
xnor U8947 (N_8947,N_7880,N_7783);
nand U8948 (N_8948,N_8001,N_7745);
nand U8949 (N_8949,N_7708,N_8044);
nand U8950 (N_8950,N_8139,N_8096);
nand U8951 (N_8951,N_7989,N_7531);
xnor U8952 (N_8952,N_7842,N_8009);
or U8953 (N_8953,N_8083,N_7829);
nand U8954 (N_8954,N_8132,N_7789);
xor U8955 (N_8955,N_7825,N_7517);
nand U8956 (N_8956,N_7971,N_7633);
nand U8957 (N_8957,N_7872,N_7613);
or U8958 (N_8958,N_8248,N_7772);
nor U8959 (N_8959,N_7778,N_7527);
xor U8960 (N_8960,N_8201,N_7635);
nor U8961 (N_8961,N_8109,N_7724);
and U8962 (N_8962,N_7722,N_7730);
nor U8963 (N_8963,N_8201,N_7875);
nand U8964 (N_8964,N_8085,N_8037);
xnor U8965 (N_8965,N_7884,N_7962);
nor U8966 (N_8966,N_7687,N_7520);
nor U8967 (N_8967,N_7592,N_7857);
nor U8968 (N_8968,N_7866,N_8247);
nand U8969 (N_8969,N_8163,N_7896);
nand U8970 (N_8970,N_7798,N_8034);
and U8971 (N_8971,N_8225,N_8203);
xnor U8972 (N_8972,N_7607,N_7985);
nor U8973 (N_8973,N_7788,N_7539);
nand U8974 (N_8974,N_7995,N_8171);
nand U8975 (N_8975,N_7772,N_7525);
nand U8976 (N_8976,N_7649,N_7637);
or U8977 (N_8977,N_8150,N_7655);
and U8978 (N_8978,N_7768,N_8238);
nor U8979 (N_8979,N_7926,N_7913);
nand U8980 (N_8980,N_7964,N_7549);
or U8981 (N_8981,N_8071,N_7856);
and U8982 (N_8982,N_7736,N_7986);
nor U8983 (N_8983,N_7729,N_8009);
nor U8984 (N_8984,N_7890,N_7516);
nor U8985 (N_8985,N_8032,N_7606);
nor U8986 (N_8986,N_8171,N_7730);
nor U8987 (N_8987,N_7717,N_8175);
and U8988 (N_8988,N_8090,N_7869);
xnor U8989 (N_8989,N_7514,N_7995);
or U8990 (N_8990,N_7565,N_7700);
and U8991 (N_8991,N_7914,N_7747);
nand U8992 (N_8992,N_8006,N_7794);
xor U8993 (N_8993,N_8227,N_7662);
and U8994 (N_8994,N_7539,N_7707);
or U8995 (N_8995,N_7508,N_7824);
or U8996 (N_8996,N_7698,N_7592);
and U8997 (N_8997,N_7986,N_8105);
nand U8998 (N_8998,N_7596,N_7704);
nand U8999 (N_8999,N_7975,N_7682);
and U9000 (N_9000,N_8366,N_8684);
nand U9001 (N_9001,N_8291,N_8799);
nand U9002 (N_9002,N_8692,N_8616);
or U9003 (N_9003,N_8800,N_8896);
xnor U9004 (N_9004,N_8642,N_8961);
xnor U9005 (N_9005,N_8995,N_8258);
xnor U9006 (N_9006,N_8831,N_8839);
and U9007 (N_9007,N_8857,N_8486);
and U9008 (N_9008,N_8308,N_8749);
or U9009 (N_9009,N_8666,N_8524);
nand U9010 (N_9010,N_8992,N_8891);
or U9011 (N_9011,N_8456,N_8461);
and U9012 (N_9012,N_8370,N_8444);
or U9013 (N_9013,N_8359,N_8372);
nor U9014 (N_9014,N_8780,N_8647);
or U9015 (N_9015,N_8882,N_8421);
or U9016 (N_9016,N_8336,N_8863);
and U9017 (N_9017,N_8674,N_8369);
and U9018 (N_9018,N_8253,N_8260);
nand U9019 (N_9019,N_8655,N_8742);
and U9020 (N_9020,N_8887,N_8406);
xor U9021 (N_9021,N_8789,N_8886);
and U9022 (N_9022,N_8772,N_8871);
or U9023 (N_9023,N_8631,N_8535);
xnor U9024 (N_9024,N_8250,N_8310);
xnor U9025 (N_9025,N_8404,N_8453);
and U9026 (N_9026,N_8256,N_8516);
or U9027 (N_9027,N_8259,N_8694);
xnor U9028 (N_9028,N_8855,N_8747);
and U9029 (N_9029,N_8832,N_8737);
or U9030 (N_9030,N_8661,N_8895);
or U9031 (N_9031,N_8822,N_8299);
nand U9032 (N_9032,N_8670,N_8521);
nor U9033 (N_9033,N_8880,N_8411);
nor U9034 (N_9034,N_8893,N_8779);
nand U9035 (N_9035,N_8858,N_8339);
and U9036 (N_9036,N_8526,N_8835);
and U9037 (N_9037,N_8695,N_8628);
nor U9038 (N_9038,N_8989,N_8614);
or U9039 (N_9039,N_8617,N_8301);
or U9040 (N_9040,N_8335,N_8463);
or U9041 (N_9041,N_8905,N_8571);
nand U9042 (N_9042,N_8271,N_8615);
and U9043 (N_9043,N_8788,N_8763);
and U9044 (N_9044,N_8562,N_8506);
nand U9045 (N_9045,N_8469,N_8813);
nor U9046 (N_9046,N_8445,N_8828);
nor U9047 (N_9047,N_8881,N_8251);
nor U9048 (N_9048,N_8906,N_8594);
and U9049 (N_9049,N_8622,N_8733);
nand U9050 (N_9050,N_8848,N_8932);
and U9051 (N_9051,N_8558,N_8326);
xor U9052 (N_9052,N_8588,N_8940);
and U9053 (N_9053,N_8634,N_8610);
or U9054 (N_9054,N_8542,N_8413);
nor U9055 (N_9055,N_8541,N_8644);
nor U9056 (N_9056,N_8830,N_8707);
or U9057 (N_9057,N_8685,N_8890);
nor U9058 (N_9058,N_8374,N_8424);
nand U9059 (N_9059,N_8270,N_8876);
nor U9060 (N_9060,N_8719,N_8912);
nor U9061 (N_9061,N_8522,N_8909);
nor U9062 (N_9062,N_8701,N_8547);
nand U9063 (N_9063,N_8637,N_8651);
nor U9064 (N_9064,N_8990,N_8405);
nor U9065 (N_9065,N_8317,N_8282);
nand U9066 (N_9066,N_8630,N_8430);
nor U9067 (N_9067,N_8868,N_8650);
or U9068 (N_9068,N_8298,N_8660);
and U9069 (N_9069,N_8416,N_8609);
or U9070 (N_9070,N_8947,N_8755);
or U9071 (N_9071,N_8693,N_8738);
nor U9072 (N_9072,N_8477,N_8636);
nor U9073 (N_9073,N_8309,N_8540);
nor U9074 (N_9074,N_8466,N_8946);
or U9075 (N_9075,N_8389,N_8409);
nor U9076 (N_9076,N_8587,N_8375);
and U9077 (N_9077,N_8425,N_8812);
xor U9078 (N_9078,N_8752,N_8872);
nand U9079 (N_9079,N_8302,N_8343);
and U9080 (N_9080,N_8801,N_8586);
nand U9081 (N_9081,N_8266,N_8728);
nand U9082 (N_9082,N_8826,N_8934);
xnor U9083 (N_9083,N_8635,N_8294);
nand U9084 (N_9084,N_8619,N_8705);
or U9085 (N_9085,N_8460,N_8681);
nor U9086 (N_9086,N_8816,N_8724);
nand U9087 (N_9087,N_8915,N_8980);
nand U9088 (N_9088,N_8950,N_8750);
nor U9089 (N_9089,N_8548,N_8532);
nor U9090 (N_9090,N_8504,N_8804);
nor U9091 (N_9091,N_8697,N_8396);
or U9092 (N_9092,N_8398,N_8721);
and U9093 (N_9093,N_8722,N_8613);
or U9094 (N_9094,N_8386,N_8585);
and U9095 (N_9095,N_8467,N_8696);
nor U9096 (N_9096,N_8774,N_8295);
or U9097 (N_9097,N_8479,N_8446);
or U9098 (N_9098,N_8926,N_8796);
or U9099 (N_9099,N_8972,N_8423);
or U9100 (N_9100,N_8599,N_8354);
xor U9101 (N_9101,N_8760,N_8536);
nor U9102 (N_9102,N_8623,N_8531);
nand U9103 (N_9103,N_8380,N_8889);
nand U9104 (N_9104,N_8598,N_8385);
nand U9105 (N_9105,N_8808,N_8546);
nor U9106 (N_9106,N_8952,N_8714);
nand U9107 (N_9107,N_8777,N_8982);
xnor U9108 (N_9108,N_8443,N_8589);
nor U9109 (N_9109,N_8713,N_8928);
or U9110 (N_9110,N_8363,N_8471);
nand U9111 (N_9111,N_8361,N_8328);
nor U9112 (N_9112,N_8323,N_8795);
nor U9113 (N_9113,N_8440,N_8407);
nand U9114 (N_9114,N_8279,N_8296);
or U9115 (N_9115,N_8347,N_8307);
nor U9116 (N_9116,N_8480,N_8942);
and U9117 (N_9117,N_8759,N_8641);
nor U9118 (N_9118,N_8392,N_8959);
nand U9119 (N_9119,N_8447,N_8803);
nand U9120 (N_9120,N_8508,N_8340);
or U9121 (N_9121,N_8578,N_8938);
nor U9122 (N_9122,N_8770,N_8873);
nand U9123 (N_9123,N_8809,N_8576);
nor U9124 (N_9124,N_8781,N_8758);
or U9125 (N_9125,N_8529,N_8498);
nand U9126 (N_9126,N_8303,N_8640);
or U9127 (N_9127,N_8496,N_8330);
or U9128 (N_9128,N_8785,N_8315);
or U9129 (N_9129,N_8358,N_8678);
and U9130 (N_9130,N_8274,N_8457);
nor U9131 (N_9131,N_8931,N_8606);
and U9132 (N_9132,N_8512,N_8807);
nand U9133 (N_9133,N_8957,N_8331);
or U9134 (N_9134,N_8834,N_8859);
xor U9135 (N_9135,N_8633,N_8936);
nand U9136 (N_9136,N_8690,N_8948);
and U9137 (N_9137,N_8493,N_8820);
nor U9138 (N_9138,N_8350,N_8953);
or U9139 (N_9139,N_8740,N_8273);
nand U9140 (N_9140,N_8514,N_8861);
or U9141 (N_9141,N_8907,N_8378);
xor U9142 (N_9142,N_8561,N_8709);
or U9143 (N_9143,N_8865,N_8679);
and U9144 (N_9144,N_8550,N_8762);
nor U9145 (N_9145,N_8341,N_8643);
nor U9146 (N_9146,N_8884,N_8929);
and U9147 (N_9147,N_8963,N_8794);
nand U9148 (N_9148,N_8439,N_8904);
or U9149 (N_9149,N_8680,N_8402);
nor U9150 (N_9150,N_8517,N_8817);
and U9151 (N_9151,N_8838,N_8559);
or U9152 (N_9152,N_8793,N_8723);
xor U9153 (N_9153,N_8659,N_8657);
or U9154 (N_9154,N_8941,N_8272);
and U9155 (N_9155,N_8582,N_8580);
nor U9156 (N_9156,N_8786,N_8870);
xor U9157 (N_9157,N_8492,N_8744);
xnor U9158 (N_9158,N_8533,N_8564);
and U9159 (N_9159,N_8263,N_8283);
or U9160 (N_9160,N_8527,N_8388);
and U9161 (N_9161,N_8844,N_8883);
and U9162 (N_9162,N_8491,N_8284);
and U9163 (N_9163,N_8811,N_8365);
or U9164 (N_9164,N_8729,N_8746);
nand U9165 (N_9165,N_8280,N_8700);
nor U9166 (N_9166,N_8824,N_8662);
nor U9167 (N_9167,N_8499,N_8939);
nand U9168 (N_9168,N_8327,N_8268);
nor U9169 (N_9169,N_8487,N_8316);
and U9170 (N_9170,N_8716,N_8821);
nor U9171 (N_9171,N_8376,N_8797);
and U9172 (N_9172,N_8583,N_8682);
nor U9173 (N_9173,N_8654,N_8265);
nor U9174 (N_9174,N_8910,N_8437);
nor U9175 (N_9175,N_8408,N_8579);
nor U9176 (N_9176,N_8379,N_8290);
nor U9177 (N_9177,N_8903,N_8563);
xnor U9178 (N_9178,N_8414,N_8255);
and U9179 (N_9179,N_8879,N_8393);
nor U9180 (N_9180,N_8567,N_8304);
nand U9181 (N_9181,N_8625,N_8656);
nor U9182 (N_9182,N_8885,N_8373);
xor U9183 (N_9183,N_8462,N_8289);
or U9184 (N_9184,N_8352,N_8761);
nand U9185 (N_9185,N_8554,N_8590);
and U9186 (N_9186,N_8305,N_8448);
or U9187 (N_9187,N_8787,N_8267);
nor U9188 (N_9188,N_8851,N_8632);
nor U9189 (N_9189,N_8484,N_8683);
and U9190 (N_9190,N_8954,N_8987);
nand U9191 (N_9191,N_8687,N_8551);
or U9192 (N_9192,N_8911,N_8669);
and U9193 (N_9193,N_8720,N_8287);
nand U9194 (N_9194,N_8704,N_8967);
nor U9195 (N_9195,N_8566,N_8814);
nor U9196 (N_9196,N_8433,N_8964);
nor U9197 (N_9197,N_8325,N_8538);
nand U9198 (N_9198,N_8739,N_8648);
and U9199 (N_9199,N_8897,N_8332);
nand U9200 (N_9200,N_8269,N_8577);
nor U9201 (N_9201,N_8845,N_8297);
nor U9202 (N_9202,N_8962,N_8856);
xnor U9203 (N_9203,N_8766,N_8502);
xnor U9204 (N_9204,N_8600,N_8288);
xor U9205 (N_9205,N_8483,N_8275);
and U9206 (N_9206,N_8968,N_8390);
and U9207 (N_9207,N_8412,N_8689);
and U9208 (N_9208,N_8410,N_8584);
or U9209 (N_9209,N_8311,N_8511);
or U9210 (N_9210,N_8557,N_8306);
nor U9211 (N_9211,N_8639,N_8473);
nor U9212 (N_9212,N_8769,N_8918);
and U9213 (N_9213,N_8397,N_8658);
nand U9214 (N_9214,N_8741,N_8878);
and U9215 (N_9215,N_8649,N_8920);
and U9216 (N_9216,N_8877,N_8348);
or U9217 (N_9217,N_8543,N_8994);
and U9218 (N_9218,N_8970,N_8368);
or U9219 (N_9219,N_8875,N_8565);
nand U9220 (N_9220,N_8537,N_8699);
or U9221 (N_9221,N_8925,N_8252);
nor U9222 (N_9222,N_8745,N_8459);
xnor U9223 (N_9223,N_8837,N_8450);
and U9224 (N_9224,N_8509,N_8474);
or U9225 (N_9225,N_8349,N_8977);
xor U9226 (N_9226,N_8342,N_8849);
xnor U9227 (N_9227,N_8597,N_8956);
nand U9228 (N_9228,N_8802,N_8555);
or U9229 (N_9229,N_8735,N_8528);
xnor U9230 (N_9230,N_8382,N_8570);
and U9231 (N_9231,N_8334,N_8346);
nand U9232 (N_9232,N_8850,N_8978);
and U9233 (N_9233,N_8998,N_8629);
and U9234 (N_9234,N_8815,N_8481);
or U9235 (N_9235,N_8573,N_8281);
or U9236 (N_9236,N_8322,N_8677);
nand U9237 (N_9237,N_8711,N_8549);
and U9238 (N_9238,N_8264,N_8703);
xor U9239 (N_9239,N_8892,N_8277);
and U9240 (N_9240,N_8778,N_8403);
nor U9241 (N_9241,N_8751,N_8494);
and U9242 (N_9242,N_8899,N_8362);
and U9243 (N_9243,N_8428,N_8596);
and U9244 (N_9244,N_8869,N_8966);
and U9245 (N_9245,N_8991,N_8426);
nor U9246 (N_9246,N_8353,N_8698);
nand U9247 (N_9247,N_8853,N_8441);
nand U9248 (N_9248,N_8922,N_8923);
or U9249 (N_9249,N_8672,N_8624);
nand U9250 (N_9250,N_8996,N_8530);
nand U9251 (N_9251,N_8860,N_8431);
nor U9252 (N_9252,N_8611,N_8556);
nand U9253 (N_9253,N_8731,N_8454);
and U9254 (N_9254,N_8429,N_8924);
and U9255 (N_9255,N_8974,N_8686);
or U9256 (N_9256,N_8945,N_8836);
xor U9257 (N_9257,N_8455,N_8621);
and U9258 (N_9258,N_8344,N_8901);
nand U9259 (N_9259,N_8917,N_8312);
nand U9260 (N_9260,N_8329,N_8846);
xor U9261 (N_9261,N_8475,N_8394);
nor U9262 (N_9262,N_8665,N_8377);
and U9263 (N_9263,N_8574,N_8999);
nor U9264 (N_9264,N_8653,N_8773);
nor U9265 (N_9265,N_8452,N_8691);
xnor U9266 (N_9266,N_8612,N_8706);
nand U9267 (N_9267,N_8935,N_8688);
xnor U9268 (N_9268,N_8485,N_8607);
xor U9269 (N_9269,N_8333,N_8864);
nor U9270 (N_9270,N_8360,N_8489);
and U9271 (N_9271,N_8320,N_8783);
nor U9272 (N_9272,N_8427,N_8627);
nand U9273 (N_9273,N_8618,N_8293);
and U9274 (N_9274,N_8958,N_8419);
nand U9275 (N_9275,N_8507,N_8927);
nor U9276 (N_9276,N_8510,N_8449);
and U9277 (N_9277,N_8842,N_8422);
and U9278 (N_9278,N_8472,N_8908);
and U9279 (N_9279,N_8673,N_8732);
nor U9280 (N_9280,N_8357,N_8768);
nor U9281 (N_9281,N_8717,N_8754);
nand U9282 (N_9282,N_8519,N_8988);
nor U9283 (N_9283,N_8791,N_8983);
or U9284 (N_9284,N_8604,N_8979);
and U9285 (N_9285,N_8726,N_8545);
nor U9286 (N_9286,N_8725,N_8417);
nand U9287 (N_9287,N_8888,N_8663);
nand U9288 (N_9288,N_8592,N_8539);
nor U9289 (N_9289,N_8748,N_8285);
or U9290 (N_9290,N_8438,N_8652);
and U9291 (N_9291,N_8810,N_8949);
xnor U9292 (N_9292,N_8675,N_8337);
and U9293 (N_9293,N_8708,N_8399);
and U9294 (N_9294,N_8490,N_8261);
nor U9295 (N_9295,N_8765,N_8391);
and U9296 (N_9296,N_8960,N_8933);
and U9297 (N_9297,N_8667,N_8913);
nand U9298 (N_9298,N_8965,N_8854);
xor U9299 (N_9299,N_8985,N_8847);
and U9300 (N_9300,N_8513,N_8955);
and U9301 (N_9301,N_8418,N_8458);
xnor U9302 (N_9302,N_8664,N_8442);
and U9303 (N_9303,N_8381,N_8645);
or U9304 (N_9304,N_8944,N_8560);
and U9305 (N_9305,N_8552,N_8862);
nor U9306 (N_9306,N_8603,N_8488);
or U9307 (N_9307,N_8367,N_8501);
or U9308 (N_9308,N_8262,N_8771);
and U9309 (N_9309,N_8401,N_8806);
xor U9310 (N_9310,N_8400,N_8436);
and U9311 (N_9311,N_8736,N_8668);
nand U9312 (N_9312,N_8916,N_8525);
nand U9313 (N_9313,N_8278,N_8395);
and U9314 (N_9314,N_8646,N_8568);
xnor U9315 (N_9315,N_8257,N_8843);
nand U9316 (N_9316,N_8495,N_8470);
nand U9317 (N_9317,N_8523,N_8753);
nand U9318 (N_9318,N_8825,N_8969);
and U9319 (N_9319,N_8318,N_8819);
nor U9320 (N_9320,N_8757,N_8581);
or U9321 (N_9321,N_8914,N_8727);
or U9322 (N_9322,N_8798,N_8671);
xnor U9323 (N_9323,N_8314,N_8482);
or U9324 (N_9324,N_8345,N_8432);
or U9325 (N_9325,N_8715,N_8503);
or U9326 (N_9326,N_8718,N_8608);
xor U9327 (N_9327,N_8971,N_8937);
nand U9328 (N_9328,N_8784,N_8321);
or U9329 (N_9329,N_8544,N_8993);
nor U9330 (N_9330,N_8833,N_8605);
or U9331 (N_9331,N_8902,N_8364);
or U9332 (N_9332,N_8792,N_8730);
nor U9333 (N_9333,N_8823,N_8973);
or U9334 (N_9334,N_8313,N_8601);
or U9335 (N_9335,N_8894,N_8767);
nor U9336 (N_9336,N_8841,N_8286);
nor U9337 (N_9337,N_8435,N_8775);
nand U9338 (N_9338,N_8593,N_8984);
nor U9339 (N_9339,N_8919,N_8702);
nand U9340 (N_9340,N_8930,N_8986);
and U9341 (N_9341,N_8776,N_8371);
nand U9342 (N_9342,N_8921,N_8569);
nor U9343 (N_9343,N_8976,N_8712);
and U9344 (N_9344,N_8324,N_8602);
nand U9345 (N_9345,N_8338,N_8829);
and U9346 (N_9346,N_8415,N_8451);
nand U9347 (N_9347,N_8874,N_8975);
nand U9348 (N_9348,N_8943,N_8319);
nor U9349 (N_9349,N_8534,N_8790);
nand U9350 (N_9350,N_8852,N_8827);
or U9351 (N_9351,N_8734,N_8898);
xnor U9352 (N_9352,N_8292,N_8505);
or U9353 (N_9353,N_8638,N_8387);
or U9354 (N_9354,N_8900,N_8997);
nor U9355 (N_9355,N_8300,N_8867);
and U9356 (N_9356,N_8626,N_8840);
nand U9357 (N_9357,N_8743,N_8981);
nor U9358 (N_9358,N_8866,N_8951);
nor U9359 (N_9359,N_8468,N_8355);
nor U9360 (N_9360,N_8676,N_8276);
and U9361 (N_9361,N_8515,N_8254);
nor U9362 (N_9362,N_8620,N_8434);
nor U9363 (N_9363,N_8575,N_8518);
nor U9364 (N_9364,N_8805,N_8591);
nand U9365 (N_9365,N_8476,N_8710);
nor U9366 (N_9366,N_8497,N_8764);
nor U9367 (N_9367,N_8478,N_8384);
and U9368 (N_9368,N_8383,N_8520);
or U9369 (N_9369,N_8351,N_8465);
nand U9370 (N_9370,N_8595,N_8553);
nor U9371 (N_9371,N_8420,N_8782);
and U9372 (N_9372,N_8572,N_8500);
nor U9373 (N_9373,N_8464,N_8356);
nor U9374 (N_9374,N_8756,N_8818);
or U9375 (N_9375,N_8667,N_8817);
or U9376 (N_9376,N_8387,N_8448);
nor U9377 (N_9377,N_8889,N_8892);
nor U9378 (N_9378,N_8840,N_8821);
and U9379 (N_9379,N_8526,N_8701);
nor U9380 (N_9380,N_8925,N_8397);
and U9381 (N_9381,N_8657,N_8618);
nand U9382 (N_9382,N_8875,N_8475);
nor U9383 (N_9383,N_8437,N_8342);
nor U9384 (N_9384,N_8756,N_8972);
or U9385 (N_9385,N_8433,N_8825);
xnor U9386 (N_9386,N_8604,N_8660);
nand U9387 (N_9387,N_8560,N_8764);
and U9388 (N_9388,N_8463,N_8964);
or U9389 (N_9389,N_8847,N_8895);
and U9390 (N_9390,N_8872,N_8823);
xor U9391 (N_9391,N_8857,N_8900);
xnor U9392 (N_9392,N_8378,N_8422);
nor U9393 (N_9393,N_8974,N_8699);
nor U9394 (N_9394,N_8290,N_8299);
xnor U9395 (N_9395,N_8656,N_8900);
or U9396 (N_9396,N_8329,N_8957);
and U9397 (N_9397,N_8385,N_8283);
and U9398 (N_9398,N_8589,N_8250);
nand U9399 (N_9399,N_8547,N_8605);
nand U9400 (N_9400,N_8693,N_8622);
nand U9401 (N_9401,N_8848,N_8516);
xor U9402 (N_9402,N_8966,N_8902);
and U9403 (N_9403,N_8843,N_8988);
and U9404 (N_9404,N_8591,N_8931);
or U9405 (N_9405,N_8331,N_8401);
or U9406 (N_9406,N_8724,N_8922);
or U9407 (N_9407,N_8654,N_8410);
and U9408 (N_9408,N_8691,N_8474);
nor U9409 (N_9409,N_8551,N_8673);
nand U9410 (N_9410,N_8612,N_8373);
nor U9411 (N_9411,N_8803,N_8954);
nand U9412 (N_9412,N_8507,N_8628);
or U9413 (N_9413,N_8822,N_8894);
nand U9414 (N_9414,N_8259,N_8384);
nor U9415 (N_9415,N_8627,N_8695);
nor U9416 (N_9416,N_8434,N_8390);
nand U9417 (N_9417,N_8940,N_8423);
and U9418 (N_9418,N_8998,N_8894);
or U9419 (N_9419,N_8437,N_8630);
and U9420 (N_9420,N_8366,N_8582);
nor U9421 (N_9421,N_8544,N_8468);
xor U9422 (N_9422,N_8644,N_8683);
or U9423 (N_9423,N_8267,N_8303);
nand U9424 (N_9424,N_8830,N_8336);
and U9425 (N_9425,N_8890,N_8615);
and U9426 (N_9426,N_8936,N_8729);
xor U9427 (N_9427,N_8516,N_8549);
nor U9428 (N_9428,N_8417,N_8679);
xor U9429 (N_9429,N_8701,N_8523);
and U9430 (N_9430,N_8644,N_8266);
or U9431 (N_9431,N_8519,N_8564);
nand U9432 (N_9432,N_8991,N_8380);
and U9433 (N_9433,N_8333,N_8806);
xnor U9434 (N_9434,N_8645,N_8829);
or U9435 (N_9435,N_8681,N_8908);
xor U9436 (N_9436,N_8809,N_8504);
and U9437 (N_9437,N_8961,N_8697);
xor U9438 (N_9438,N_8603,N_8499);
nand U9439 (N_9439,N_8802,N_8753);
nor U9440 (N_9440,N_8961,N_8381);
nand U9441 (N_9441,N_8576,N_8964);
xor U9442 (N_9442,N_8377,N_8983);
xor U9443 (N_9443,N_8964,N_8812);
or U9444 (N_9444,N_8973,N_8319);
xor U9445 (N_9445,N_8390,N_8640);
or U9446 (N_9446,N_8367,N_8259);
or U9447 (N_9447,N_8690,N_8668);
or U9448 (N_9448,N_8747,N_8757);
and U9449 (N_9449,N_8499,N_8396);
or U9450 (N_9450,N_8605,N_8462);
xnor U9451 (N_9451,N_8597,N_8865);
and U9452 (N_9452,N_8691,N_8587);
nand U9453 (N_9453,N_8760,N_8876);
nor U9454 (N_9454,N_8523,N_8666);
nor U9455 (N_9455,N_8925,N_8930);
xnor U9456 (N_9456,N_8282,N_8445);
or U9457 (N_9457,N_8835,N_8583);
or U9458 (N_9458,N_8614,N_8470);
nand U9459 (N_9459,N_8936,N_8342);
nor U9460 (N_9460,N_8534,N_8285);
nor U9461 (N_9461,N_8663,N_8531);
and U9462 (N_9462,N_8882,N_8334);
nor U9463 (N_9463,N_8838,N_8795);
or U9464 (N_9464,N_8637,N_8995);
or U9465 (N_9465,N_8601,N_8563);
nand U9466 (N_9466,N_8890,N_8755);
nand U9467 (N_9467,N_8441,N_8985);
nor U9468 (N_9468,N_8853,N_8504);
nand U9469 (N_9469,N_8706,N_8523);
nor U9470 (N_9470,N_8783,N_8474);
nor U9471 (N_9471,N_8965,N_8563);
and U9472 (N_9472,N_8833,N_8980);
nand U9473 (N_9473,N_8290,N_8367);
nor U9474 (N_9474,N_8780,N_8964);
or U9475 (N_9475,N_8634,N_8874);
nor U9476 (N_9476,N_8253,N_8362);
nand U9477 (N_9477,N_8310,N_8930);
nand U9478 (N_9478,N_8568,N_8394);
and U9479 (N_9479,N_8317,N_8943);
nor U9480 (N_9480,N_8800,N_8437);
xnor U9481 (N_9481,N_8768,N_8399);
nor U9482 (N_9482,N_8559,N_8622);
and U9483 (N_9483,N_8755,N_8879);
nor U9484 (N_9484,N_8499,N_8783);
nand U9485 (N_9485,N_8395,N_8575);
and U9486 (N_9486,N_8823,N_8828);
nor U9487 (N_9487,N_8550,N_8765);
nor U9488 (N_9488,N_8863,N_8831);
nor U9489 (N_9489,N_8484,N_8357);
nand U9490 (N_9490,N_8299,N_8890);
and U9491 (N_9491,N_8534,N_8799);
xnor U9492 (N_9492,N_8609,N_8769);
and U9493 (N_9493,N_8771,N_8873);
nand U9494 (N_9494,N_8548,N_8381);
xnor U9495 (N_9495,N_8963,N_8422);
or U9496 (N_9496,N_8981,N_8725);
nand U9497 (N_9497,N_8843,N_8439);
xnor U9498 (N_9498,N_8788,N_8648);
xor U9499 (N_9499,N_8811,N_8946);
and U9500 (N_9500,N_8881,N_8693);
and U9501 (N_9501,N_8530,N_8613);
and U9502 (N_9502,N_8296,N_8908);
or U9503 (N_9503,N_8349,N_8478);
and U9504 (N_9504,N_8530,N_8429);
nand U9505 (N_9505,N_8261,N_8369);
xor U9506 (N_9506,N_8435,N_8770);
nand U9507 (N_9507,N_8611,N_8839);
or U9508 (N_9508,N_8818,N_8628);
xnor U9509 (N_9509,N_8661,N_8901);
and U9510 (N_9510,N_8630,N_8800);
or U9511 (N_9511,N_8544,N_8504);
and U9512 (N_9512,N_8960,N_8905);
nor U9513 (N_9513,N_8623,N_8587);
nor U9514 (N_9514,N_8400,N_8800);
nand U9515 (N_9515,N_8727,N_8376);
or U9516 (N_9516,N_8883,N_8787);
or U9517 (N_9517,N_8507,N_8808);
nand U9518 (N_9518,N_8693,N_8787);
and U9519 (N_9519,N_8763,N_8948);
and U9520 (N_9520,N_8417,N_8497);
nand U9521 (N_9521,N_8555,N_8953);
or U9522 (N_9522,N_8599,N_8973);
nand U9523 (N_9523,N_8832,N_8963);
and U9524 (N_9524,N_8520,N_8951);
or U9525 (N_9525,N_8711,N_8699);
nand U9526 (N_9526,N_8536,N_8935);
nand U9527 (N_9527,N_8866,N_8355);
and U9528 (N_9528,N_8813,N_8913);
and U9529 (N_9529,N_8278,N_8512);
nand U9530 (N_9530,N_8368,N_8917);
and U9531 (N_9531,N_8915,N_8875);
nor U9532 (N_9532,N_8699,N_8987);
or U9533 (N_9533,N_8305,N_8996);
and U9534 (N_9534,N_8445,N_8780);
nand U9535 (N_9535,N_8778,N_8583);
nand U9536 (N_9536,N_8335,N_8393);
and U9537 (N_9537,N_8803,N_8547);
xor U9538 (N_9538,N_8699,N_8328);
or U9539 (N_9539,N_8607,N_8414);
or U9540 (N_9540,N_8911,N_8901);
nor U9541 (N_9541,N_8259,N_8595);
nor U9542 (N_9542,N_8723,N_8508);
nor U9543 (N_9543,N_8391,N_8734);
or U9544 (N_9544,N_8651,N_8613);
nand U9545 (N_9545,N_8280,N_8406);
nor U9546 (N_9546,N_8737,N_8960);
nand U9547 (N_9547,N_8456,N_8780);
nand U9548 (N_9548,N_8529,N_8609);
or U9549 (N_9549,N_8888,N_8864);
nand U9550 (N_9550,N_8468,N_8374);
and U9551 (N_9551,N_8402,N_8314);
or U9552 (N_9552,N_8395,N_8329);
and U9553 (N_9553,N_8445,N_8881);
nor U9554 (N_9554,N_8485,N_8984);
nor U9555 (N_9555,N_8767,N_8828);
nor U9556 (N_9556,N_8631,N_8450);
nor U9557 (N_9557,N_8563,N_8845);
nor U9558 (N_9558,N_8370,N_8320);
nor U9559 (N_9559,N_8518,N_8872);
and U9560 (N_9560,N_8976,N_8446);
nand U9561 (N_9561,N_8505,N_8772);
xor U9562 (N_9562,N_8989,N_8271);
and U9563 (N_9563,N_8981,N_8436);
nor U9564 (N_9564,N_8783,N_8870);
xnor U9565 (N_9565,N_8538,N_8584);
or U9566 (N_9566,N_8816,N_8674);
nor U9567 (N_9567,N_8318,N_8893);
or U9568 (N_9568,N_8784,N_8634);
or U9569 (N_9569,N_8297,N_8901);
nand U9570 (N_9570,N_8799,N_8833);
and U9571 (N_9571,N_8419,N_8931);
and U9572 (N_9572,N_8366,N_8981);
xor U9573 (N_9573,N_8337,N_8681);
nor U9574 (N_9574,N_8343,N_8520);
and U9575 (N_9575,N_8889,N_8418);
and U9576 (N_9576,N_8741,N_8666);
nand U9577 (N_9577,N_8387,N_8590);
nor U9578 (N_9578,N_8549,N_8545);
nor U9579 (N_9579,N_8331,N_8538);
and U9580 (N_9580,N_8904,N_8518);
and U9581 (N_9581,N_8556,N_8512);
and U9582 (N_9582,N_8556,N_8544);
nand U9583 (N_9583,N_8871,N_8886);
or U9584 (N_9584,N_8685,N_8930);
or U9585 (N_9585,N_8325,N_8876);
and U9586 (N_9586,N_8510,N_8430);
nor U9587 (N_9587,N_8396,N_8784);
and U9588 (N_9588,N_8433,N_8655);
and U9589 (N_9589,N_8768,N_8532);
nor U9590 (N_9590,N_8937,N_8791);
and U9591 (N_9591,N_8913,N_8768);
and U9592 (N_9592,N_8778,N_8312);
nand U9593 (N_9593,N_8340,N_8333);
xor U9594 (N_9594,N_8584,N_8840);
xnor U9595 (N_9595,N_8643,N_8344);
xnor U9596 (N_9596,N_8843,N_8735);
xor U9597 (N_9597,N_8597,N_8774);
and U9598 (N_9598,N_8684,N_8763);
nand U9599 (N_9599,N_8556,N_8587);
or U9600 (N_9600,N_8325,N_8912);
xnor U9601 (N_9601,N_8380,N_8852);
xor U9602 (N_9602,N_8700,N_8660);
or U9603 (N_9603,N_8887,N_8563);
or U9604 (N_9604,N_8660,N_8911);
nand U9605 (N_9605,N_8439,N_8542);
nand U9606 (N_9606,N_8540,N_8891);
nor U9607 (N_9607,N_8446,N_8636);
nor U9608 (N_9608,N_8592,N_8566);
or U9609 (N_9609,N_8401,N_8410);
or U9610 (N_9610,N_8507,N_8790);
or U9611 (N_9611,N_8298,N_8260);
nor U9612 (N_9612,N_8803,N_8262);
and U9613 (N_9613,N_8596,N_8584);
nand U9614 (N_9614,N_8683,N_8366);
and U9615 (N_9615,N_8850,N_8991);
nor U9616 (N_9616,N_8976,N_8874);
or U9617 (N_9617,N_8797,N_8844);
nor U9618 (N_9618,N_8250,N_8448);
and U9619 (N_9619,N_8277,N_8928);
and U9620 (N_9620,N_8505,N_8551);
or U9621 (N_9621,N_8331,N_8746);
or U9622 (N_9622,N_8393,N_8928);
or U9623 (N_9623,N_8401,N_8663);
or U9624 (N_9624,N_8691,N_8441);
nand U9625 (N_9625,N_8963,N_8922);
nand U9626 (N_9626,N_8420,N_8568);
or U9627 (N_9627,N_8991,N_8776);
nand U9628 (N_9628,N_8743,N_8628);
nand U9629 (N_9629,N_8294,N_8318);
and U9630 (N_9630,N_8880,N_8567);
nor U9631 (N_9631,N_8467,N_8288);
nand U9632 (N_9632,N_8524,N_8956);
nor U9633 (N_9633,N_8639,N_8534);
nand U9634 (N_9634,N_8807,N_8566);
nand U9635 (N_9635,N_8704,N_8341);
nor U9636 (N_9636,N_8565,N_8939);
xor U9637 (N_9637,N_8748,N_8517);
or U9638 (N_9638,N_8535,N_8559);
and U9639 (N_9639,N_8813,N_8302);
nor U9640 (N_9640,N_8499,N_8313);
nand U9641 (N_9641,N_8911,N_8924);
nand U9642 (N_9642,N_8619,N_8261);
and U9643 (N_9643,N_8486,N_8719);
or U9644 (N_9644,N_8283,N_8551);
and U9645 (N_9645,N_8944,N_8898);
and U9646 (N_9646,N_8256,N_8548);
nand U9647 (N_9647,N_8735,N_8637);
nand U9648 (N_9648,N_8343,N_8345);
and U9649 (N_9649,N_8584,N_8975);
xnor U9650 (N_9650,N_8477,N_8706);
or U9651 (N_9651,N_8945,N_8497);
nand U9652 (N_9652,N_8496,N_8730);
and U9653 (N_9653,N_8610,N_8770);
nand U9654 (N_9654,N_8846,N_8976);
xor U9655 (N_9655,N_8900,N_8326);
or U9656 (N_9656,N_8724,N_8793);
nand U9657 (N_9657,N_8727,N_8817);
and U9658 (N_9658,N_8527,N_8387);
and U9659 (N_9659,N_8508,N_8436);
nor U9660 (N_9660,N_8421,N_8566);
and U9661 (N_9661,N_8917,N_8883);
and U9662 (N_9662,N_8867,N_8516);
nor U9663 (N_9663,N_8873,N_8864);
nand U9664 (N_9664,N_8984,N_8678);
nand U9665 (N_9665,N_8974,N_8774);
and U9666 (N_9666,N_8948,N_8710);
nand U9667 (N_9667,N_8383,N_8847);
nor U9668 (N_9668,N_8555,N_8275);
xor U9669 (N_9669,N_8588,N_8837);
nor U9670 (N_9670,N_8823,N_8731);
nand U9671 (N_9671,N_8933,N_8538);
or U9672 (N_9672,N_8337,N_8997);
nand U9673 (N_9673,N_8418,N_8897);
nand U9674 (N_9674,N_8866,N_8676);
and U9675 (N_9675,N_8543,N_8649);
or U9676 (N_9676,N_8262,N_8558);
nor U9677 (N_9677,N_8865,N_8589);
xor U9678 (N_9678,N_8697,N_8557);
nand U9679 (N_9679,N_8623,N_8584);
nand U9680 (N_9680,N_8862,N_8404);
or U9681 (N_9681,N_8486,N_8325);
nand U9682 (N_9682,N_8625,N_8520);
nand U9683 (N_9683,N_8524,N_8487);
and U9684 (N_9684,N_8521,N_8726);
or U9685 (N_9685,N_8604,N_8727);
nor U9686 (N_9686,N_8329,N_8381);
nand U9687 (N_9687,N_8739,N_8594);
and U9688 (N_9688,N_8816,N_8938);
nand U9689 (N_9689,N_8400,N_8446);
nor U9690 (N_9690,N_8482,N_8772);
nand U9691 (N_9691,N_8610,N_8632);
and U9692 (N_9692,N_8861,N_8737);
or U9693 (N_9693,N_8343,N_8630);
or U9694 (N_9694,N_8541,N_8717);
or U9695 (N_9695,N_8333,N_8459);
and U9696 (N_9696,N_8262,N_8706);
nor U9697 (N_9697,N_8901,N_8432);
xor U9698 (N_9698,N_8717,N_8423);
and U9699 (N_9699,N_8980,N_8394);
and U9700 (N_9700,N_8466,N_8652);
nand U9701 (N_9701,N_8967,N_8715);
or U9702 (N_9702,N_8411,N_8390);
or U9703 (N_9703,N_8801,N_8695);
nor U9704 (N_9704,N_8520,N_8305);
xnor U9705 (N_9705,N_8338,N_8748);
nor U9706 (N_9706,N_8838,N_8464);
and U9707 (N_9707,N_8719,N_8588);
and U9708 (N_9708,N_8492,N_8367);
xnor U9709 (N_9709,N_8741,N_8783);
and U9710 (N_9710,N_8732,N_8599);
nor U9711 (N_9711,N_8570,N_8639);
and U9712 (N_9712,N_8773,N_8752);
or U9713 (N_9713,N_8524,N_8294);
nor U9714 (N_9714,N_8487,N_8327);
xor U9715 (N_9715,N_8403,N_8387);
nand U9716 (N_9716,N_8743,N_8585);
or U9717 (N_9717,N_8612,N_8657);
or U9718 (N_9718,N_8825,N_8917);
nor U9719 (N_9719,N_8580,N_8331);
nor U9720 (N_9720,N_8632,N_8385);
nor U9721 (N_9721,N_8771,N_8344);
nand U9722 (N_9722,N_8274,N_8745);
and U9723 (N_9723,N_8627,N_8776);
nor U9724 (N_9724,N_8684,N_8486);
xor U9725 (N_9725,N_8874,N_8641);
or U9726 (N_9726,N_8593,N_8460);
nor U9727 (N_9727,N_8620,N_8869);
nor U9728 (N_9728,N_8871,N_8289);
or U9729 (N_9729,N_8916,N_8506);
or U9730 (N_9730,N_8770,N_8959);
and U9731 (N_9731,N_8448,N_8283);
nor U9732 (N_9732,N_8620,N_8866);
and U9733 (N_9733,N_8992,N_8689);
and U9734 (N_9734,N_8680,N_8384);
nand U9735 (N_9735,N_8450,N_8541);
and U9736 (N_9736,N_8340,N_8646);
nand U9737 (N_9737,N_8393,N_8740);
nand U9738 (N_9738,N_8320,N_8997);
nand U9739 (N_9739,N_8464,N_8806);
and U9740 (N_9740,N_8594,N_8550);
nor U9741 (N_9741,N_8956,N_8489);
nor U9742 (N_9742,N_8426,N_8453);
nor U9743 (N_9743,N_8949,N_8801);
xor U9744 (N_9744,N_8771,N_8371);
and U9745 (N_9745,N_8794,N_8912);
and U9746 (N_9746,N_8398,N_8927);
or U9747 (N_9747,N_8452,N_8839);
or U9748 (N_9748,N_8835,N_8928);
nand U9749 (N_9749,N_8536,N_8609);
nand U9750 (N_9750,N_9122,N_9177);
and U9751 (N_9751,N_9555,N_9529);
nand U9752 (N_9752,N_9330,N_9183);
nor U9753 (N_9753,N_9028,N_9577);
xnor U9754 (N_9754,N_9109,N_9352);
nor U9755 (N_9755,N_9245,N_9171);
and U9756 (N_9756,N_9656,N_9651);
xor U9757 (N_9757,N_9269,N_9460);
and U9758 (N_9758,N_9632,N_9483);
and U9759 (N_9759,N_9433,N_9251);
and U9760 (N_9760,N_9542,N_9070);
nor U9761 (N_9761,N_9075,N_9221);
and U9762 (N_9762,N_9061,N_9337);
nand U9763 (N_9763,N_9504,N_9107);
and U9764 (N_9764,N_9021,N_9272);
nor U9765 (N_9765,N_9519,N_9489);
or U9766 (N_9766,N_9151,N_9682);
or U9767 (N_9767,N_9304,N_9267);
nor U9768 (N_9768,N_9455,N_9486);
nand U9769 (N_9769,N_9132,N_9194);
nand U9770 (N_9770,N_9643,N_9633);
or U9771 (N_9771,N_9142,N_9627);
nor U9772 (N_9772,N_9473,N_9017);
nand U9773 (N_9773,N_9408,N_9226);
or U9774 (N_9774,N_9650,N_9378);
nor U9775 (N_9775,N_9724,N_9383);
xnor U9776 (N_9776,N_9457,N_9260);
nor U9777 (N_9777,N_9343,N_9686);
and U9778 (N_9778,N_9363,N_9299);
or U9779 (N_9779,N_9339,N_9557);
and U9780 (N_9780,N_9034,N_9647);
and U9781 (N_9781,N_9141,N_9564);
nor U9782 (N_9782,N_9406,N_9289);
and U9783 (N_9783,N_9749,N_9691);
nor U9784 (N_9784,N_9083,N_9032);
nand U9785 (N_9785,N_9574,N_9683);
nor U9786 (N_9786,N_9192,N_9409);
nand U9787 (N_9787,N_9106,N_9035);
nand U9788 (N_9788,N_9273,N_9618);
nand U9789 (N_9789,N_9646,N_9582);
or U9790 (N_9790,N_9156,N_9560);
or U9791 (N_9791,N_9162,N_9741);
nand U9792 (N_9792,N_9305,N_9105);
nor U9793 (N_9793,N_9585,N_9625);
nand U9794 (N_9794,N_9392,N_9456);
and U9795 (N_9795,N_9622,N_9572);
xor U9796 (N_9796,N_9197,N_9354);
nand U9797 (N_9797,N_9620,N_9131);
nor U9798 (N_9798,N_9054,N_9401);
nor U9799 (N_9799,N_9018,N_9187);
nand U9800 (N_9800,N_9371,N_9550);
and U9801 (N_9801,N_9563,N_9702);
and U9802 (N_9802,N_9502,N_9246);
or U9803 (N_9803,N_9279,N_9041);
nand U9804 (N_9804,N_9224,N_9199);
nor U9805 (N_9805,N_9638,N_9206);
nand U9806 (N_9806,N_9748,N_9518);
xor U9807 (N_9807,N_9358,N_9700);
nor U9808 (N_9808,N_9520,N_9480);
or U9809 (N_9809,N_9710,N_9499);
and U9810 (N_9810,N_9076,N_9185);
nor U9811 (N_9811,N_9393,N_9575);
or U9812 (N_9812,N_9303,N_9368);
or U9813 (N_9813,N_9482,N_9168);
and U9814 (N_9814,N_9008,N_9324);
nand U9815 (N_9815,N_9096,N_9616);
nor U9816 (N_9816,N_9362,N_9009);
or U9817 (N_9817,N_9191,N_9039);
nor U9818 (N_9818,N_9531,N_9711);
nor U9819 (N_9819,N_9495,N_9416);
nand U9820 (N_9820,N_9101,N_9088);
or U9821 (N_9821,N_9341,N_9373);
and U9822 (N_9822,N_9715,N_9268);
nor U9823 (N_9823,N_9115,N_9503);
nand U9824 (N_9824,N_9287,N_9612);
nor U9825 (N_9825,N_9025,N_9441);
and U9826 (N_9826,N_9325,N_9739);
nand U9827 (N_9827,N_9628,N_9584);
and U9828 (N_9828,N_9117,N_9227);
xor U9829 (N_9829,N_9551,N_9006);
nand U9830 (N_9830,N_9188,N_9547);
nor U9831 (N_9831,N_9410,N_9218);
and U9832 (N_9832,N_9467,N_9478);
nand U9833 (N_9833,N_9400,N_9522);
nor U9834 (N_9834,N_9728,N_9334);
or U9835 (N_9835,N_9417,N_9309);
nor U9836 (N_9836,N_9357,N_9022);
nand U9837 (N_9837,N_9615,N_9641);
or U9838 (N_9838,N_9234,N_9443);
and U9839 (N_9839,N_9621,N_9252);
xor U9840 (N_9840,N_9385,N_9386);
nand U9841 (N_9841,N_9461,N_9387);
nand U9842 (N_9842,N_9228,N_9326);
xnor U9843 (N_9843,N_9388,N_9698);
xnor U9844 (N_9844,N_9462,N_9669);
and U9845 (N_9845,N_9327,N_9716);
or U9846 (N_9846,N_9244,N_9573);
or U9847 (N_9847,N_9554,N_9605);
nor U9848 (N_9848,N_9202,N_9587);
nand U9849 (N_9849,N_9237,N_9431);
nand U9850 (N_9850,N_9578,N_9422);
nand U9851 (N_9851,N_9407,N_9336);
and U9852 (N_9852,N_9614,N_9681);
nor U9853 (N_9853,N_9254,N_9005);
and U9854 (N_9854,N_9674,N_9415);
nand U9855 (N_9855,N_9182,N_9404);
nor U9856 (N_9856,N_9207,N_9571);
and U9857 (N_9857,N_9723,N_9003);
xnor U9858 (N_9858,N_9536,N_9212);
or U9859 (N_9859,N_9527,N_9057);
xor U9860 (N_9860,N_9316,N_9544);
nor U9861 (N_9861,N_9217,N_9219);
or U9862 (N_9862,N_9720,N_9013);
nand U9863 (N_9863,N_9498,N_9423);
nor U9864 (N_9864,N_9263,N_9127);
or U9865 (N_9865,N_9428,N_9320);
and U9866 (N_9866,N_9421,N_9617);
nand U9867 (N_9867,N_9747,N_9049);
or U9868 (N_9868,N_9092,N_9258);
nand U9869 (N_9869,N_9538,N_9328);
nor U9870 (N_9870,N_9414,N_9223);
or U9871 (N_9871,N_9033,N_9012);
nand U9872 (N_9872,N_9155,N_9465);
or U9873 (N_9873,N_9568,N_9562);
xnor U9874 (N_9874,N_9277,N_9434);
or U9875 (N_9875,N_9082,N_9174);
and U9876 (N_9876,N_9446,N_9472);
or U9877 (N_9877,N_9089,N_9660);
nand U9878 (N_9878,N_9190,N_9173);
and U9879 (N_9879,N_9093,N_9319);
xor U9880 (N_9880,N_9559,N_9042);
nor U9881 (N_9881,N_9055,N_9610);
and U9882 (N_9882,N_9491,N_9001);
nor U9883 (N_9883,N_9528,N_9290);
or U9884 (N_9884,N_9595,N_9425);
and U9885 (N_9885,N_9717,N_9043);
nand U9886 (N_9886,N_9470,N_9379);
or U9887 (N_9887,N_9126,N_9091);
or U9888 (N_9888,N_9654,N_9133);
nor U9889 (N_9889,N_9360,N_9344);
or U9890 (N_9890,N_9271,N_9424);
nor U9891 (N_9891,N_9721,N_9558);
xnor U9892 (N_9892,N_9213,N_9347);
nand U9893 (N_9893,N_9149,N_9052);
nand U9894 (N_9894,N_9231,N_9589);
or U9895 (N_9895,N_9230,N_9448);
nand U9896 (N_9896,N_9282,N_9350);
and U9897 (N_9897,N_9604,N_9514);
and U9898 (N_9898,N_9007,N_9077);
nor U9899 (N_9899,N_9023,N_9210);
nor U9900 (N_9900,N_9157,N_9186);
and U9901 (N_9901,N_9275,N_9016);
nand U9902 (N_9902,N_9725,N_9069);
or U9903 (N_9903,N_9123,N_9592);
nand U9904 (N_9904,N_9450,N_9530);
nand U9905 (N_9905,N_9624,N_9214);
nor U9906 (N_9906,N_9100,N_9429);
or U9907 (N_9907,N_9736,N_9015);
nand U9908 (N_9908,N_9160,N_9338);
xnor U9909 (N_9909,N_9479,N_9137);
nand U9910 (N_9910,N_9420,N_9738);
or U9911 (N_9911,N_9667,N_9389);
or U9912 (N_9912,N_9639,N_9209);
or U9913 (N_9913,N_9685,N_9180);
and U9914 (N_9914,N_9349,N_9477);
xor U9915 (N_9915,N_9636,N_9073);
nand U9916 (N_9916,N_9678,N_9361);
and U9917 (N_9917,N_9516,N_9570);
nor U9918 (N_9918,N_9014,N_9204);
nor U9919 (N_9919,N_9024,N_9356);
nand U9920 (N_9920,N_9283,N_9597);
nor U9921 (N_9921,N_9644,N_9537);
or U9922 (N_9922,N_9545,N_9637);
nor U9923 (N_9923,N_9493,N_9611);
nand U9924 (N_9924,N_9232,N_9040);
nand U9925 (N_9925,N_9068,N_9376);
and U9926 (N_9926,N_9193,N_9098);
and U9927 (N_9927,N_9200,N_9458);
nor U9928 (N_9928,N_9038,N_9048);
and U9929 (N_9929,N_9340,N_9552);
nor U9930 (N_9930,N_9265,N_9364);
and U9931 (N_9931,N_9099,N_9619);
and U9932 (N_9932,N_9395,N_9118);
or U9933 (N_9933,N_9261,N_9418);
and U9934 (N_9934,N_9136,N_9445);
and U9935 (N_9935,N_9694,N_9047);
and U9936 (N_9936,N_9238,N_9381);
or U9937 (N_9937,N_9313,N_9242);
nand U9938 (N_9938,N_9396,N_9648);
xor U9939 (N_9939,N_9399,N_9342);
nor U9940 (N_9940,N_9085,N_9487);
nor U9941 (N_9941,N_9439,N_9044);
nand U9942 (N_9942,N_9285,N_9300);
nand U9943 (N_9943,N_9590,N_9365);
xnor U9944 (N_9944,N_9152,N_9072);
nor U9945 (N_9945,N_9317,N_9284);
or U9946 (N_9946,N_9370,N_9440);
and U9947 (N_9947,N_9066,N_9010);
and U9948 (N_9948,N_9121,N_9372);
xor U9949 (N_9949,N_9634,N_9293);
and U9950 (N_9950,N_9134,N_9201);
xnor U9951 (N_9951,N_9384,N_9288);
nor U9952 (N_9952,N_9655,N_9394);
or U9953 (N_9953,N_9027,N_9144);
nor U9954 (N_9954,N_9463,N_9466);
nor U9955 (N_9955,N_9081,N_9524);
and U9956 (N_9956,N_9129,N_9161);
and U9957 (N_9957,N_9707,N_9490);
nand U9958 (N_9958,N_9247,N_9566);
or U9959 (N_9959,N_9124,N_9167);
nand U9960 (N_9960,N_9703,N_9579);
xnor U9961 (N_9961,N_9642,N_9561);
or U9962 (N_9962,N_9256,N_9084);
or U9963 (N_9963,N_9539,N_9355);
or U9964 (N_9964,N_9153,N_9526);
and U9965 (N_9965,N_9169,N_9146);
or U9966 (N_9966,N_9494,N_9172);
or U9967 (N_9967,N_9278,N_9074);
nand U9968 (N_9968,N_9517,N_9509);
xor U9969 (N_9969,N_9398,N_9672);
or U9970 (N_9970,N_9195,N_9053);
and U9971 (N_9971,N_9645,N_9591);
or U9972 (N_9972,N_9189,N_9351);
or U9973 (N_9973,N_9692,N_9664);
and U9974 (N_9974,N_9332,N_9405);
nand U9975 (N_9975,N_9501,N_9427);
or U9976 (N_9976,N_9020,N_9159);
or U9977 (N_9977,N_9451,N_9744);
nor U9978 (N_9978,N_9165,N_9110);
nor U9979 (N_9979,N_9497,N_9150);
nand U9980 (N_9980,N_9178,N_9203);
nor U9981 (N_9981,N_9447,N_9649);
nor U9982 (N_9982,N_9500,N_9696);
nand U9983 (N_9983,N_9732,N_9248);
and U9984 (N_9984,N_9143,N_9062);
nor U9985 (N_9985,N_9059,N_9629);
nor U9986 (N_9986,N_9170,N_9176);
nor U9987 (N_9987,N_9481,N_9496);
and U9988 (N_9988,N_9080,N_9255);
nor U9989 (N_9989,N_9525,N_9154);
and U9990 (N_9990,N_9051,N_9546);
and U9991 (N_9991,N_9593,N_9659);
and U9992 (N_9992,N_9452,N_9677);
nor U9993 (N_9993,N_9603,N_9046);
xnor U9994 (N_9994,N_9704,N_9216);
nand U9995 (N_9995,N_9735,N_9484);
or U9996 (N_9996,N_9722,N_9366);
and U9997 (N_9997,N_9719,N_9543);
nor U9998 (N_9998,N_9274,N_9331);
and U9999 (N_9999,N_9145,N_9222);
nor U10000 (N_10000,N_9270,N_9097);
nand U10001 (N_10001,N_9599,N_9454);
and U10002 (N_10002,N_9468,N_9179);
nor U10003 (N_10003,N_9130,N_9158);
nand U10004 (N_10004,N_9588,N_9050);
nand U10005 (N_10005,N_9631,N_9243);
xor U10006 (N_10006,N_9679,N_9662);
or U10007 (N_10007,N_9533,N_9166);
nor U10008 (N_10008,N_9689,N_9291);
and U10009 (N_10009,N_9281,N_9652);
xnor U10010 (N_10010,N_9675,N_9019);
or U10011 (N_10011,N_9184,N_9580);
or U10012 (N_10012,N_9321,N_9567);
nor U10013 (N_10013,N_9714,N_9112);
nand U10014 (N_10014,N_9147,N_9469);
xor U10015 (N_10015,N_9163,N_9506);
xnor U10016 (N_10016,N_9532,N_9708);
xor U10017 (N_10017,N_9727,N_9430);
nand U10018 (N_10018,N_9078,N_9437);
or U10019 (N_10019,N_9128,N_9556);
nand U10020 (N_10020,N_9307,N_9485);
and U10021 (N_10021,N_9064,N_9310);
and U10022 (N_10022,N_9175,N_9718);
nand U10023 (N_10023,N_9668,N_9280);
nor U10024 (N_10024,N_9004,N_9297);
nand U10025 (N_10025,N_9693,N_9402);
nand U10026 (N_10026,N_9276,N_9390);
nand U10027 (N_10027,N_9298,N_9581);
or U10028 (N_10028,N_9635,N_9507);
or U10029 (N_10029,N_9374,N_9661);
nand U10030 (N_10030,N_9476,N_9333);
or U10031 (N_10031,N_9239,N_9671);
nor U10032 (N_10032,N_9412,N_9094);
nand U10033 (N_10033,N_9695,N_9598);
and U10034 (N_10034,N_9111,N_9295);
nor U10035 (N_10035,N_9548,N_9697);
nand U10036 (N_10036,N_9733,N_9135);
and U10037 (N_10037,N_9680,N_9623);
and U10038 (N_10038,N_9726,N_9712);
xnor U10039 (N_10039,N_9391,N_9535);
or U10040 (N_10040,N_9444,N_9000);
or U10041 (N_10041,N_9515,N_9250);
or U10042 (N_10042,N_9541,N_9403);
and U10043 (N_10043,N_9116,N_9030);
nor U10044 (N_10044,N_9138,N_9508);
and U10045 (N_10045,N_9011,N_9653);
nand U10046 (N_10046,N_9240,N_9318);
nand U10047 (N_10047,N_9449,N_9411);
nor U10048 (N_10048,N_9488,N_9353);
nand U10049 (N_10049,N_9513,N_9253);
and U10050 (N_10050,N_9065,N_9583);
and U10051 (N_10051,N_9308,N_9380);
or U10052 (N_10052,N_9346,N_9302);
or U10053 (N_10053,N_9464,N_9705);
nor U10054 (N_10054,N_9676,N_9067);
and U10055 (N_10055,N_9139,N_9596);
and U10056 (N_10056,N_9459,N_9103);
or U10057 (N_10057,N_9348,N_9225);
nand U10058 (N_10058,N_9731,N_9315);
nor U10059 (N_10059,N_9257,N_9684);
nor U10060 (N_10060,N_9262,N_9523);
and U10061 (N_10061,N_9699,N_9148);
xnor U10062 (N_10062,N_9296,N_9534);
nor U10063 (N_10063,N_9688,N_9301);
xnor U10064 (N_10064,N_9345,N_9211);
nand U10065 (N_10065,N_9569,N_9602);
nor U10066 (N_10066,N_9323,N_9215);
xnor U10067 (N_10067,N_9576,N_9229);
nor U10068 (N_10068,N_9663,N_9397);
nor U10069 (N_10069,N_9438,N_9521);
and U10070 (N_10070,N_9031,N_9036);
nor U10071 (N_10071,N_9613,N_9037);
nand U10072 (N_10072,N_9367,N_9670);
or U10073 (N_10073,N_9474,N_9745);
and U10074 (N_10074,N_9071,N_9312);
nor U10075 (N_10075,N_9586,N_9549);
xnor U10076 (N_10076,N_9090,N_9140);
xnor U10077 (N_10077,N_9594,N_9359);
and U10078 (N_10078,N_9746,N_9426);
nor U10079 (N_10079,N_9119,N_9259);
and U10080 (N_10080,N_9264,N_9233);
xnor U10081 (N_10081,N_9294,N_9609);
nor U10082 (N_10082,N_9730,N_9164);
nor U10083 (N_10083,N_9235,N_9492);
or U10084 (N_10084,N_9181,N_9079);
or U10085 (N_10085,N_9205,N_9029);
nand U10086 (N_10086,N_9740,N_9512);
and U10087 (N_10087,N_9286,N_9666);
nor U10088 (N_10088,N_9442,N_9436);
nand U10089 (N_10089,N_9087,N_9737);
xnor U10090 (N_10090,N_9208,N_9060);
xnor U10091 (N_10091,N_9220,N_9435);
nand U10092 (N_10092,N_9553,N_9673);
or U10093 (N_10093,N_9665,N_9102);
xor U10094 (N_10094,N_9026,N_9640);
nand U10095 (N_10095,N_9058,N_9236);
xnor U10096 (N_10096,N_9505,N_9565);
nand U10097 (N_10097,N_9729,N_9113);
nand U10098 (N_10098,N_9056,N_9314);
nand U10099 (N_10099,N_9453,N_9742);
nand U10100 (N_10100,N_9600,N_9329);
or U10101 (N_10101,N_9095,N_9292);
and U10102 (N_10102,N_9630,N_9657);
and U10103 (N_10103,N_9601,N_9306);
and U10104 (N_10104,N_9713,N_9377);
or U10105 (N_10105,N_9086,N_9241);
nor U10106 (N_10106,N_9249,N_9413);
nor U10107 (N_10107,N_9607,N_9701);
nor U10108 (N_10108,N_9322,N_9432);
nor U10109 (N_10109,N_9734,N_9690);
nand U10110 (N_10110,N_9311,N_9125);
nor U10111 (N_10111,N_9196,N_9335);
and U10112 (N_10112,N_9510,N_9114);
nor U10113 (N_10113,N_9687,N_9419);
and U10114 (N_10114,N_9104,N_9471);
xor U10115 (N_10115,N_9540,N_9375);
nor U10116 (N_10116,N_9120,N_9608);
and U10117 (N_10117,N_9475,N_9382);
xnor U10118 (N_10118,N_9063,N_9369);
xor U10119 (N_10119,N_9709,N_9658);
or U10120 (N_10120,N_9626,N_9743);
and U10121 (N_10121,N_9108,N_9511);
nand U10122 (N_10122,N_9198,N_9002);
or U10123 (N_10123,N_9706,N_9606);
nand U10124 (N_10124,N_9045,N_9266);
nand U10125 (N_10125,N_9322,N_9134);
nand U10126 (N_10126,N_9725,N_9249);
nand U10127 (N_10127,N_9270,N_9014);
nand U10128 (N_10128,N_9749,N_9567);
and U10129 (N_10129,N_9410,N_9393);
xnor U10130 (N_10130,N_9279,N_9031);
or U10131 (N_10131,N_9367,N_9120);
and U10132 (N_10132,N_9222,N_9200);
nand U10133 (N_10133,N_9496,N_9256);
nor U10134 (N_10134,N_9160,N_9302);
nor U10135 (N_10135,N_9393,N_9274);
or U10136 (N_10136,N_9556,N_9104);
nand U10137 (N_10137,N_9415,N_9704);
xor U10138 (N_10138,N_9126,N_9182);
or U10139 (N_10139,N_9351,N_9049);
or U10140 (N_10140,N_9463,N_9365);
nand U10141 (N_10141,N_9174,N_9595);
nor U10142 (N_10142,N_9000,N_9016);
nor U10143 (N_10143,N_9618,N_9506);
nand U10144 (N_10144,N_9338,N_9337);
xor U10145 (N_10145,N_9266,N_9293);
or U10146 (N_10146,N_9450,N_9490);
nand U10147 (N_10147,N_9529,N_9649);
or U10148 (N_10148,N_9491,N_9561);
and U10149 (N_10149,N_9454,N_9073);
or U10150 (N_10150,N_9196,N_9688);
nor U10151 (N_10151,N_9050,N_9287);
nor U10152 (N_10152,N_9170,N_9738);
nor U10153 (N_10153,N_9624,N_9309);
and U10154 (N_10154,N_9360,N_9350);
nand U10155 (N_10155,N_9566,N_9629);
and U10156 (N_10156,N_9041,N_9242);
and U10157 (N_10157,N_9489,N_9398);
and U10158 (N_10158,N_9179,N_9091);
xnor U10159 (N_10159,N_9033,N_9421);
and U10160 (N_10160,N_9569,N_9433);
or U10161 (N_10161,N_9153,N_9113);
and U10162 (N_10162,N_9405,N_9748);
or U10163 (N_10163,N_9196,N_9451);
and U10164 (N_10164,N_9392,N_9278);
nand U10165 (N_10165,N_9011,N_9557);
or U10166 (N_10166,N_9081,N_9718);
and U10167 (N_10167,N_9155,N_9519);
nand U10168 (N_10168,N_9268,N_9104);
nand U10169 (N_10169,N_9498,N_9367);
and U10170 (N_10170,N_9179,N_9139);
xor U10171 (N_10171,N_9159,N_9638);
nor U10172 (N_10172,N_9305,N_9193);
and U10173 (N_10173,N_9304,N_9286);
or U10174 (N_10174,N_9678,N_9017);
or U10175 (N_10175,N_9198,N_9011);
nor U10176 (N_10176,N_9145,N_9440);
and U10177 (N_10177,N_9270,N_9110);
nor U10178 (N_10178,N_9556,N_9654);
or U10179 (N_10179,N_9086,N_9437);
nor U10180 (N_10180,N_9387,N_9732);
nand U10181 (N_10181,N_9318,N_9146);
xor U10182 (N_10182,N_9270,N_9133);
nor U10183 (N_10183,N_9037,N_9464);
xnor U10184 (N_10184,N_9024,N_9394);
nand U10185 (N_10185,N_9592,N_9210);
nand U10186 (N_10186,N_9605,N_9242);
and U10187 (N_10187,N_9718,N_9203);
and U10188 (N_10188,N_9366,N_9698);
and U10189 (N_10189,N_9134,N_9060);
nand U10190 (N_10190,N_9625,N_9682);
and U10191 (N_10191,N_9097,N_9469);
nor U10192 (N_10192,N_9736,N_9349);
nor U10193 (N_10193,N_9690,N_9422);
or U10194 (N_10194,N_9207,N_9458);
or U10195 (N_10195,N_9533,N_9056);
or U10196 (N_10196,N_9275,N_9380);
nand U10197 (N_10197,N_9054,N_9720);
and U10198 (N_10198,N_9610,N_9057);
nor U10199 (N_10199,N_9647,N_9104);
or U10200 (N_10200,N_9093,N_9298);
xor U10201 (N_10201,N_9285,N_9301);
nor U10202 (N_10202,N_9253,N_9331);
and U10203 (N_10203,N_9197,N_9618);
or U10204 (N_10204,N_9171,N_9697);
nor U10205 (N_10205,N_9434,N_9227);
and U10206 (N_10206,N_9659,N_9742);
nand U10207 (N_10207,N_9173,N_9378);
or U10208 (N_10208,N_9562,N_9478);
or U10209 (N_10209,N_9399,N_9201);
and U10210 (N_10210,N_9262,N_9403);
and U10211 (N_10211,N_9423,N_9142);
and U10212 (N_10212,N_9350,N_9320);
nand U10213 (N_10213,N_9308,N_9741);
and U10214 (N_10214,N_9616,N_9543);
nand U10215 (N_10215,N_9338,N_9172);
nand U10216 (N_10216,N_9461,N_9403);
nand U10217 (N_10217,N_9235,N_9179);
nor U10218 (N_10218,N_9334,N_9571);
nand U10219 (N_10219,N_9405,N_9153);
or U10220 (N_10220,N_9678,N_9302);
and U10221 (N_10221,N_9334,N_9499);
nor U10222 (N_10222,N_9136,N_9363);
and U10223 (N_10223,N_9050,N_9522);
and U10224 (N_10224,N_9022,N_9283);
nor U10225 (N_10225,N_9720,N_9503);
and U10226 (N_10226,N_9280,N_9640);
nor U10227 (N_10227,N_9726,N_9286);
nor U10228 (N_10228,N_9661,N_9045);
xnor U10229 (N_10229,N_9404,N_9660);
nand U10230 (N_10230,N_9129,N_9589);
or U10231 (N_10231,N_9699,N_9690);
nor U10232 (N_10232,N_9169,N_9623);
nand U10233 (N_10233,N_9185,N_9094);
and U10234 (N_10234,N_9536,N_9165);
nor U10235 (N_10235,N_9323,N_9445);
nor U10236 (N_10236,N_9310,N_9206);
and U10237 (N_10237,N_9551,N_9072);
nor U10238 (N_10238,N_9313,N_9325);
or U10239 (N_10239,N_9498,N_9586);
nor U10240 (N_10240,N_9274,N_9558);
and U10241 (N_10241,N_9700,N_9256);
nand U10242 (N_10242,N_9703,N_9298);
or U10243 (N_10243,N_9730,N_9395);
nor U10244 (N_10244,N_9145,N_9742);
or U10245 (N_10245,N_9061,N_9446);
nand U10246 (N_10246,N_9250,N_9368);
nand U10247 (N_10247,N_9054,N_9623);
and U10248 (N_10248,N_9499,N_9347);
nor U10249 (N_10249,N_9394,N_9260);
or U10250 (N_10250,N_9347,N_9076);
nor U10251 (N_10251,N_9489,N_9652);
or U10252 (N_10252,N_9448,N_9099);
nand U10253 (N_10253,N_9450,N_9043);
or U10254 (N_10254,N_9592,N_9261);
nor U10255 (N_10255,N_9045,N_9314);
nor U10256 (N_10256,N_9116,N_9548);
and U10257 (N_10257,N_9259,N_9489);
nor U10258 (N_10258,N_9445,N_9313);
xor U10259 (N_10259,N_9146,N_9113);
or U10260 (N_10260,N_9341,N_9019);
xnor U10261 (N_10261,N_9023,N_9201);
and U10262 (N_10262,N_9176,N_9734);
xnor U10263 (N_10263,N_9742,N_9470);
or U10264 (N_10264,N_9161,N_9085);
or U10265 (N_10265,N_9169,N_9637);
xor U10266 (N_10266,N_9425,N_9125);
nor U10267 (N_10267,N_9201,N_9054);
and U10268 (N_10268,N_9495,N_9376);
nor U10269 (N_10269,N_9596,N_9723);
nor U10270 (N_10270,N_9190,N_9308);
nand U10271 (N_10271,N_9733,N_9598);
nand U10272 (N_10272,N_9362,N_9051);
and U10273 (N_10273,N_9715,N_9475);
and U10274 (N_10274,N_9409,N_9527);
nor U10275 (N_10275,N_9743,N_9631);
and U10276 (N_10276,N_9480,N_9404);
and U10277 (N_10277,N_9278,N_9605);
nand U10278 (N_10278,N_9187,N_9243);
and U10279 (N_10279,N_9147,N_9029);
xnor U10280 (N_10280,N_9692,N_9738);
nor U10281 (N_10281,N_9036,N_9278);
or U10282 (N_10282,N_9218,N_9330);
nor U10283 (N_10283,N_9300,N_9188);
nor U10284 (N_10284,N_9376,N_9074);
or U10285 (N_10285,N_9462,N_9154);
nor U10286 (N_10286,N_9024,N_9028);
nand U10287 (N_10287,N_9522,N_9452);
nand U10288 (N_10288,N_9364,N_9661);
or U10289 (N_10289,N_9180,N_9202);
nand U10290 (N_10290,N_9349,N_9503);
xnor U10291 (N_10291,N_9542,N_9224);
or U10292 (N_10292,N_9718,N_9477);
nand U10293 (N_10293,N_9746,N_9421);
nor U10294 (N_10294,N_9071,N_9491);
and U10295 (N_10295,N_9653,N_9128);
nand U10296 (N_10296,N_9193,N_9036);
nor U10297 (N_10297,N_9360,N_9603);
nor U10298 (N_10298,N_9529,N_9489);
and U10299 (N_10299,N_9083,N_9317);
xnor U10300 (N_10300,N_9060,N_9643);
and U10301 (N_10301,N_9387,N_9027);
or U10302 (N_10302,N_9711,N_9423);
and U10303 (N_10303,N_9741,N_9291);
or U10304 (N_10304,N_9527,N_9464);
nor U10305 (N_10305,N_9368,N_9616);
nand U10306 (N_10306,N_9524,N_9555);
and U10307 (N_10307,N_9614,N_9705);
and U10308 (N_10308,N_9123,N_9604);
nor U10309 (N_10309,N_9408,N_9158);
or U10310 (N_10310,N_9304,N_9025);
nor U10311 (N_10311,N_9059,N_9403);
and U10312 (N_10312,N_9624,N_9745);
and U10313 (N_10313,N_9017,N_9348);
xor U10314 (N_10314,N_9233,N_9596);
or U10315 (N_10315,N_9058,N_9483);
nor U10316 (N_10316,N_9140,N_9431);
or U10317 (N_10317,N_9248,N_9501);
and U10318 (N_10318,N_9650,N_9314);
nor U10319 (N_10319,N_9202,N_9177);
xor U10320 (N_10320,N_9723,N_9117);
nor U10321 (N_10321,N_9255,N_9627);
nand U10322 (N_10322,N_9254,N_9298);
and U10323 (N_10323,N_9464,N_9558);
nand U10324 (N_10324,N_9177,N_9685);
or U10325 (N_10325,N_9003,N_9058);
nor U10326 (N_10326,N_9173,N_9697);
and U10327 (N_10327,N_9639,N_9175);
xor U10328 (N_10328,N_9387,N_9283);
nor U10329 (N_10329,N_9704,N_9505);
and U10330 (N_10330,N_9369,N_9064);
or U10331 (N_10331,N_9164,N_9470);
xor U10332 (N_10332,N_9270,N_9481);
nor U10333 (N_10333,N_9177,N_9307);
xor U10334 (N_10334,N_9369,N_9343);
and U10335 (N_10335,N_9214,N_9642);
nand U10336 (N_10336,N_9537,N_9748);
nand U10337 (N_10337,N_9017,N_9469);
and U10338 (N_10338,N_9204,N_9481);
nor U10339 (N_10339,N_9523,N_9455);
nand U10340 (N_10340,N_9616,N_9594);
nor U10341 (N_10341,N_9623,N_9161);
or U10342 (N_10342,N_9116,N_9731);
and U10343 (N_10343,N_9224,N_9348);
nand U10344 (N_10344,N_9363,N_9009);
nor U10345 (N_10345,N_9112,N_9095);
or U10346 (N_10346,N_9039,N_9113);
or U10347 (N_10347,N_9446,N_9673);
and U10348 (N_10348,N_9524,N_9170);
nand U10349 (N_10349,N_9511,N_9313);
or U10350 (N_10350,N_9461,N_9368);
and U10351 (N_10351,N_9133,N_9010);
or U10352 (N_10352,N_9274,N_9397);
nand U10353 (N_10353,N_9463,N_9539);
nor U10354 (N_10354,N_9508,N_9460);
nor U10355 (N_10355,N_9478,N_9017);
nand U10356 (N_10356,N_9061,N_9049);
xor U10357 (N_10357,N_9654,N_9419);
and U10358 (N_10358,N_9250,N_9274);
or U10359 (N_10359,N_9191,N_9031);
and U10360 (N_10360,N_9354,N_9366);
xnor U10361 (N_10361,N_9515,N_9733);
nor U10362 (N_10362,N_9047,N_9730);
and U10363 (N_10363,N_9667,N_9611);
nand U10364 (N_10364,N_9710,N_9573);
or U10365 (N_10365,N_9628,N_9626);
or U10366 (N_10366,N_9105,N_9500);
nand U10367 (N_10367,N_9274,N_9247);
or U10368 (N_10368,N_9114,N_9639);
nor U10369 (N_10369,N_9634,N_9567);
xor U10370 (N_10370,N_9465,N_9231);
nor U10371 (N_10371,N_9498,N_9016);
nor U10372 (N_10372,N_9497,N_9534);
nor U10373 (N_10373,N_9032,N_9391);
nand U10374 (N_10374,N_9710,N_9315);
nand U10375 (N_10375,N_9220,N_9599);
nand U10376 (N_10376,N_9065,N_9144);
xnor U10377 (N_10377,N_9321,N_9370);
and U10378 (N_10378,N_9264,N_9102);
and U10379 (N_10379,N_9676,N_9605);
and U10380 (N_10380,N_9468,N_9004);
and U10381 (N_10381,N_9518,N_9438);
or U10382 (N_10382,N_9655,N_9164);
or U10383 (N_10383,N_9478,N_9689);
nor U10384 (N_10384,N_9417,N_9640);
nand U10385 (N_10385,N_9644,N_9138);
and U10386 (N_10386,N_9704,N_9089);
nor U10387 (N_10387,N_9658,N_9626);
nor U10388 (N_10388,N_9351,N_9435);
nor U10389 (N_10389,N_9733,N_9327);
and U10390 (N_10390,N_9560,N_9616);
and U10391 (N_10391,N_9463,N_9235);
or U10392 (N_10392,N_9110,N_9185);
or U10393 (N_10393,N_9331,N_9469);
or U10394 (N_10394,N_9618,N_9699);
nand U10395 (N_10395,N_9268,N_9628);
and U10396 (N_10396,N_9395,N_9686);
nand U10397 (N_10397,N_9699,N_9510);
nand U10398 (N_10398,N_9480,N_9566);
and U10399 (N_10399,N_9332,N_9171);
nor U10400 (N_10400,N_9335,N_9248);
nor U10401 (N_10401,N_9027,N_9061);
or U10402 (N_10402,N_9436,N_9596);
and U10403 (N_10403,N_9329,N_9375);
nor U10404 (N_10404,N_9259,N_9437);
nand U10405 (N_10405,N_9541,N_9747);
xnor U10406 (N_10406,N_9116,N_9285);
or U10407 (N_10407,N_9746,N_9080);
or U10408 (N_10408,N_9402,N_9441);
and U10409 (N_10409,N_9184,N_9501);
nor U10410 (N_10410,N_9712,N_9149);
and U10411 (N_10411,N_9062,N_9499);
and U10412 (N_10412,N_9325,N_9667);
or U10413 (N_10413,N_9342,N_9281);
xor U10414 (N_10414,N_9092,N_9204);
nor U10415 (N_10415,N_9028,N_9725);
or U10416 (N_10416,N_9249,N_9290);
nor U10417 (N_10417,N_9748,N_9221);
nand U10418 (N_10418,N_9463,N_9284);
and U10419 (N_10419,N_9304,N_9144);
xnor U10420 (N_10420,N_9511,N_9330);
or U10421 (N_10421,N_9637,N_9692);
and U10422 (N_10422,N_9575,N_9492);
nor U10423 (N_10423,N_9015,N_9311);
or U10424 (N_10424,N_9479,N_9391);
or U10425 (N_10425,N_9311,N_9726);
nor U10426 (N_10426,N_9244,N_9382);
nor U10427 (N_10427,N_9112,N_9657);
nor U10428 (N_10428,N_9733,N_9457);
and U10429 (N_10429,N_9504,N_9490);
xor U10430 (N_10430,N_9688,N_9427);
nor U10431 (N_10431,N_9159,N_9602);
and U10432 (N_10432,N_9186,N_9277);
or U10433 (N_10433,N_9117,N_9745);
xor U10434 (N_10434,N_9735,N_9665);
or U10435 (N_10435,N_9135,N_9301);
or U10436 (N_10436,N_9641,N_9411);
nor U10437 (N_10437,N_9071,N_9118);
nand U10438 (N_10438,N_9193,N_9032);
nor U10439 (N_10439,N_9478,N_9571);
or U10440 (N_10440,N_9582,N_9287);
nand U10441 (N_10441,N_9529,N_9048);
nand U10442 (N_10442,N_9398,N_9270);
nand U10443 (N_10443,N_9539,N_9345);
or U10444 (N_10444,N_9736,N_9507);
or U10445 (N_10445,N_9689,N_9500);
and U10446 (N_10446,N_9456,N_9674);
xor U10447 (N_10447,N_9501,N_9233);
nor U10448 (N_10448,N_9570,N_9290);
and U10449 (N_10449,N_9434,N_9189);
or U10450 (N_10450,N_9731,N_9563);
nand U10451 (N_10451,N_9456,N_9524);
nor U10452 (N_10452,N_9282,N_9626);
nand U10453 (N_10453,N_9256,N_9070);
and U10454 (N_10454,N_9489,N_9342);
or U10455 (N_10455,N_9616,N_9383);
or U10456 (N_10456,N_9584,N_9106);
and U10457 (N_10457,N_9337,N_9726);
and U10458 (N_10458,N_9389,N_9372);
and U10459 (N_10459,N_9488,N_9665);
or U10460 (N_10460,N_9399,N_9245);
and U10461 (N_10461,N_9718,N_9253);
nor U10462 (N_10462,N_9661,N_9037);
or U10463 (N_10463,N_9617,N_9550);
and U10464 (N_10464,N_9513,N_9290);
nor U10465 (N_10465,N_9032,N_9574);
nor U10466 (N_10466,N_9534,N_9379);
nand U10467 (N_10467,N_9728,N_9250);
nand U10468 (N_10468,N_9336,N_9097);
nand U10469 (N_10469,N_9257,N_9019);
nor U10470 (N_10470,N_9318,N_9089);
nor U10471 (N_10471,N_9646,N_9290);
xor U10472 (N_10472,N_9556,N_9259);
xnor U10473 (N_10473,N_9290,N_9542);
nor U10474 (N_10474,N_9618,N_9308);
nor U10475 (N_10475,N_9694,N_9626);
or U10476 (N_10476,N_9447,N_9554);
and U10477 (N_10477,N_9634,N_9708);
nor U10478 (N_10478,N_9027,N_9165);
nor U10479 (N_10479,N_9502,N_9285);
nand U10480 (N_10480,N_9397,N_9748);
and U10481 (N_10481,N_9104,N_9635);
xor U10482 (N_10482,N_9748,N_9255);
nand U10483 (N_10483,N_9660,N_9632);
and U10484 (N_10484,N_9328,N_9497);
and U10485 (N_10485,N_9509,N_9460);
and U10486 (N_10486,N_9233,N_9205);
nand U10487 (N_10487,N_9492,N_9421);
or U10488 (N_10488,N_9586,N_9597);
nand U10489 (N_10489,N_9047,N_9688);
nor U10490 (N_10490,N_9612,N_9051);
xnor U10491 (N_10491,N_9673,N_9508);
nand U10492 (N_10492,N_9176,N_9391);
or U10493 (N_10493,N_9279,N_9603);
and U10494 (N_10494,N_9473,N_9472);
nand U10495 (N_10495,N_9159,N_9520);
or U10496 (N_10496,N_9052,N_9655);
nand U10497 (N_10497,N_9213,N_9685);
xnor U10498 (N_10498,N_9737,N_9230);
nor U10499 (N_10499,N_9610,N_9369);
nor U10500 (N_10500,N_10067,N_10479);
nor U10501 (N_10501,N_9955,N_10338);
or U10502 (N_10502,N_10088,N_10426);
or U10503 (N_10503,N_10093,N_10268);
nand U10504 (N_10504,N_9947,N_10474);
and U10505 (N_10505,N_10347,N_9840);
nand U10506 (N_10506,N_10096,N_10113);
nor U10507 (N_10507,N_10138,N_10133);
nand U10508 (N_10508,N_10069,N_10361);
nor U10509 (N_10509,N_10380,N_10490);
nand U10510 (N_10510,N_10124,N_10345);
nor U10511 (N_10511,N_10022,N_10107);
and U10512 (N_10512,N_10484,N_9877);
and U10513 (N_10513,N_10005,N_9874);
or U10514 (N_10514,N_10452,N_10074);
and U10515 (N_10515,N_9987,N_9882);
and U10516 (N_10516,N_9858,N_10368);
and U10517 (N_10517,N_9920,N_9883);
nor U10518 (N_10518,N_10171,N_9907);
nor U10519 (N_10519,N_10386,N_10416);
nand U10520 (N_10520,N_10343,N_10421);
xnor U10521 (N_10521,N_10495,N_10125);
or U10522 (N_10522,N_10436,N_10434);
nor U10523 (N_10523,N_10390,N_10132);
xor U10524 (N_10524,N_10139,N_10020);
or U10525 (N_10525,N_10265,N_10085);
nand U10526 (N_10526,N_10425,N_10051);
and U10527 (N_10527,N_9752,N_9948);
or U10528 (N_10528,N_10378,N_10038);
xor U10529 (N_10529,N_9972,N_10059);
or U10530 (N_10530,N_9782,N_10234);
xnor U10531 (N_10531,N_10236,N_10207);
xnor U10532 (N_10532,N_9884,N_10325);
or U10533 (N_10533,N_10470,N_9838);
nor U10534 (N_10534,N_9846,N_10449);
or U10535 (N_10535,N_10097,N_10217);
nand U10536 (N_10536,N_10087,N_10428);
xnor U10537 (N_10537,N_10057,N_10246);
nor U10538 (N_10538,N_10204,N_10066);
xor U10539 (N_10539,N_10457,N_10205);
and U10540 (N_10540,N_10120,N_10092);
xor U10541 (N_10541,N_10017,N_9985);
nor U10542 (N_10542,N_10257,N_10456);
or U10543 (N_10543,N_9962,N_9945);
and U10544 (N_10544,N_10279,N_10342);
and U10545 (N_10545,N_10458,N_10135);
or U10546 (N_10546,N_9906,N_10160);
xnor U10547 (N_10547,N_9901,N_10102);
nand U10548 (N_10548,N_10350,N_10369);
nor U10549 (N_10549,N_9779,N_10154);
and U10550 (N_10550,N_9844,N_9815);
and U10551 (N_10551,N_9759,N_10199);
nand U10552 (N_10552,N_10100,N_10267);
or U10553 (N_10553,N_10036,N_10188);
and U10554 (N_10554,N_9814,N_10251);
or U10555 (N_10555,N_10134,N_9809);
and U10556 (N_10556,N_10119,N_10219);
nor U10557 (N_10557,N_10404,N_10394);
nand U10558 (N_10558,N_9892,N_9876);
or U10559 (N_10559,N_10300,N_10318);
nor U10560 (N_10560,N_10354,N_10001);
or U10561 (N_10561,N_9850,N_10213);
and U10562 (N_10562,N_10221,N_9848);
and U10563 (N_10563,N_10179,N_10043);
and U10564 (N_10564,N_10168,N_10237);
and U10565 (N_10565,N_10060,N_9761);
nand U10566 (N_10566,N_9764,N_10439);
and U10567 (N_10567,N_10052,N_10231);
and U10568 (N_10568,N_10025,N_9956);
and U10569 (N_10569,N_10376,N_10109);
and U10570 (N_10570,N_9821,N_9810);
nand U10571 (N_10571,N_10482,N_9767);
or U10572 (N_10572,N_9750,N_9903);
nand U10573 (N_10573,N_10201,N_10453);
nand U10574 (N_10574,N_9833,N_10131);
xor U10575 (N_10575,N_9989,N_9834);
and U10576 (N_10576,N_10411,N_10061);
or U10577 (N_10577,N_10117,N_10090);
and U10578 (N_10578,N_9781,N_10371);
xor U10579 (N_10579,N_9860,N_10169);
xnor U10580 (N_10580,N_10245,N_10389);
nor U10581 (N_10581,N_10370,N_9842);
xor U10582 (N_10582,N_9847,N_10225);
or U10583 (N_10583,N_9852,N_9983);
and U10584 (N_10584,N_10309,N_10098);
nor U10585 (N_10585,N_9916,N_10110);
or U10586 (N_10586,N_9953,N_10095);
nor U10587 (N_10587,N_9885,N_9942);
nand U10588 (N_10588,N_10270,N_10483);
nor U10589 (N_10589,N_10152,N_9855);
nand U10590 (N_10590,N_10004,N_9902);
nor U10591 (N_10591,N_10491,N_10239);
or U10592 (N_10592,N_9872,N_10336);
xor U10593 (N_10593,N_10140,N_10281);
nor U10594 (N_10594,N_10377,N_10280);
nor U10595 (N_10595,N_10356,N_9856);
and U10596 (N_10596,N_9946,N_10312);
or U10597 (N_10597,N_10197,N_9992);
or U10598 (N_10598,N_10299,N_9836);
or U10599 (N_10599,N_10297,N_9961);
and U10600 (N_10600,N_10012,N_10030);
or U10601 (N_10601,N_10327,N_10071);
or U10602 (N_10602,N_10282,N_9807);
and U10603 (N_10603,N_10202,N_10193);
and U10604 (N_10604,N_10401,N_10405);
or U10605 (N_10605,N_9918,N_10435);
nor U10606 (N_10606,N_10487,N_10230);
nor U10607 (N_10607,N_10332,N_10440);
nor U10608 (N_10608,N_9830,N_9870);
nor U10609 (N_10609,N_10162,N_10349);
nand U10610 (N_10610,N_9887,N_10247);
and U10611 (N_10611,N_10399,N_9880);
and U10612 (N_10612,N_10116,N_10341);
nand U10613 (N_10613,N_10142,N_10015);
and U10614 (N_10614,N_9954,N_9806);
or U10615 (N_10615,N_9969,N_10497);
or U10616 (N_10616,N_10387,N_10208);
nor U10617 (N_10617,N_10407,N_9811);
nor U10618 (N_10618,N_10126,N_9762);
xnor U10619 (N_10619,N_10419,N_9952);
and U10620 (N_10620,N_9853,N_10240);
nand U10621 (N_10621,N_10473,N_10478);
or U10622 (N_10622,N_9801,N_9826);
xor U10623 (N_10623,N_10464,N_9968);
nand U10624 (N_10624,N_10210,N_10146);
and U10625 (N_10625,N_10235,N_9794);
nor U10626 (N_10626,N_10010,N_10460);
and U10627 (N_10627,N_10198,N_10226);
nor U10628 (N_10628,N_9775,N_10330);
or U10629 (N_10629,N_9827,N_10329);
nand U10630 (N_10630,N_10196,N_10224);
nand U10631 (N_10631,N_10252,N_10437);
nor U10632 (N_10632,N_9912,N_9974);
nor U10633 (N_10633,N_10200,N_9758);
nand U10634 (N_10634,N_10469,N_10155);
and U10635 (N_10635,N_9819,N_10291);
nor U10636 (N_10636,N_10047,N_9997);
nor U10637 (N_10637,N_10447,N_9949);
nand U10638 (N_10638,N_9756,N_9796);
and U10639 (N_10639,N_10393,N_10078);
nor U10640 (N_10640,N_9891,N_10159);
or U10641 (N_10641,N_9973,N_10357);
and U10642 (N_10642,N_9793,N_10276);
or U10643 (N_10643,N_9965,N_10072);
nor U10644 (N_10644,N_10333,N_10158);
nand U10645 (N_10645,N_10054,N_9982);
or U10646 (N_10646,N_9923,N_9932);
nor U10647 (N_10647,N_10311,N_10148);
nand U10648 (N_10648,N_9790,N_10170);
xnor U10649 (N_10649,N_10499,N_10422);
xnor U10650 (N_10650,N_10278,N_10304);
nand U10651 (N_10651,N_9928,N_10128);
or U10652 (N_10652,N_10182,N_10056);
nand U10653 (N_10653,N_9929,N_10438);
and U10654 (N_10654,N_9978,N_9986);
or U10655 (N_10655,N_9879,N_10101);
nor U10656 (N_10656,N_10408,N_10151);
and U10657 (N_10657,N_10454,N_9958);
or U10658 (N_10658,N_10445,N_10122);
nor U10659 (N_10659,N_9957,N_10150);
nor U10660 (N_10660,N_10335,N_10303);
nor U10661 (N_10661,N_9890,N_10053);
nand U10662 (N_10662,N_10307,N_9896);
nand U10663 (N_10663,N_10292,N_10014);
or U10664 (N_10664,N_9990,N_10396);
and U10665 (N_10665,N_9805,N_10023);
and U10666 (N_10666,N_10352,N_10403);
nand U10667 (N_10667,N_10383,N_10033);
nand U10668 (N_10668,N_10076,N_9754);
nand U10669 (N_10669,N_10018,N_10286);
or U10670 (N_10670,N_10176,N_10398);
nor U10671 (N_10671,N_9924,N_10242);
and U10672 (N_10672,N_10415,N_9869);
nor U10673 (N_10673,N_10021,N_10183);
and U10674 (N_10674,N_9976,N_9895);
and U10675 (N_10675,N_10254,N_10039);
or U10676 (N_10676,N_10147,N_10353);
nor U10677 (N_10677,N_9977,N_9996);
and U10678 (N_10678,N_9820,N_10256);
or U10679 (N_10679,N_10189,N_10358);
and U10680 (N_10680,N_10296,N_10472);
nor U10681 (N_10681,N_10273,N_10156);
nand U10682 (N_10682,N_10003,N_10264);
and U10683 (N_10683,N_10326,N_10105);
xor U10684 (N_10684,N_9888,N_10498);
nor U10685 (N_10685,N_9886,N_10123);
or U10686 (N_10686,N_9785,N_9894);
nand U10687 (N_10687,N_10164,N_10400);
or U10688 (N_10688,N_10448,N_9900);
xnor U10689 (N_10689,N_10184,N_10143);
or U10690 (N_10690,N_10418,N_10375);
nand U10691 (N_10691,N_10442,N_10459);
and U10692 (N_10692,N_9919,N_10190);
or U10693 (N_10693,N_10172,N_10037);
xor U10694 (N_10694,N_9934,N_9927);
and U10695 (N_10695,N_10175,N_10044);
and U10696 (N_10696,N_10410,N_9898);
nand U10697 (N_10697,N_10395,N_10379);
and U10698 (N_10698,N_10374,N_9849);
and U10699 (N_10699,N_9913,N_9998);
nand U10700 (N_10700,N_10082,N_10322);
xnor U10701 (N_10701,N_10366,N_10382);
nand U10702 (N_10702,N_9795,N_10244);
nand U10703 (N_10703,N_10417,N_10137);
nor U10704 (N_10704,N_10058,N_9800);
or U10705 (N_10705,N_9915,N_9950);
xor U10706 (N_10706,N_9993,N_10424);
or U10707 (N_10707,N_9798,N_10228);
nor U10708 (N_10708,N_10465,N_10446);
xnor U10709 (N_10709,N_9802,N_9763);
and U10710 (N_10710,N_10262,N_10463);
nor U10711 (N_10711,N_10181,N_10372);
and U10712 (N_10712,N_10191,N_9804);
nor U10713 (N_10713,N_10031,N_10480);
nor U10714 (N_10714,N_9788,N_10289);
and U10715 (N_10715,N_10091,N_9936);
or U10716 (N_10716,N_9831,N_10308);
nor U10717 (N_10717,N_9816,N_10255);
or U10718 (N_10718,N_9937,N_9959);
nand U10719 (N_10719,N_10315,N_10272);
and U10720 (N_10720,N_10466,N_10359);
or U10721 (N_10721,N_10346,N_9864);
and U10722 (N_10722,N_9889,N_10223);
nand U10723 (N_10723,N_10263,N_10388);
or U10724 (N_10724,N_10266,N_10063);
and U10725 (N_10725,N_10227,N_10314);
and U10726 (N_10726,N_10385,N_10130);
nor U10727 (N_10727,N_10046,N_9941);
nand U10728 (N_10728,N_10024,N_10178);
and U10729 (N_10729,N_10032,N_10215);
or U10730 (N_10730,N_9975,N_10310);
nand U10731 (N_10731,N_9921,N_10451);
nor U10732 (N_10732,N_10153,N_10000);
nor U10733 (N_10733,N_10002,N_9818);
or U10734 (N_10734,N_9862,N_9935);
and U10735 (N_10735,N_9765,N_9873);
or U10736 (N_10736,N_10313,N_9881);
nor U10737 (N_10737,N_9766,N_10209);
or U10738 (N_10738,N_9909,N_9971);
or U10739 (N_10739,N_9780,N_10115);
nand U10740 (N_10740,N_10261,N_9940);
nor U10741 (N_10741,N_10136,N_9784);
nor U10742 (N_10742,N_9776,N_10049);
nand U10743 (N_10743,N_10080,N_10275);
nor U10744 (N_10744,N_10174,N_10145);
or U10745 (N_10745,N_10064,N_9861);
nor U10746 (N_10746,N_10355,N_10402);
or U10747 (N_10747,N_10218,N_9899);
nand U10748 (N_10748,N_10269,N_9843);
nor U10749 (N_10749,N_9812,N_10441);
nand U10750 (N_10750,N_9813,N_10492);
nand U10751 (N_10751,N_10250,N_9837);
xor U10752 (N_10752,N_10035,N_10086);
nor U10753 (N_10753,N_10420,N_9803);
or U10754 (N_10754,N_10290,N_10238);
or U10755 (N_10755,N_10042,N_10485);
or U10756 (N_10756,N_10328,N_9773);
nor U10757 (N_10757,N_9772,N_10302);
and U10758 (N_10758,N_10344,N_9925);
nor U10759 (N_10759,N_10323,N_10362);
and U10760 (N_10760,N_9966,N_10229);
nand U10761 (N_10761,N_10011,N_10481);
and U10762 (N_10762,N_9867,N_10287);
or U10763 (N_10763,N_10099,N_10214);
nand U10764 (N_10764,N_10065,N_10206);
nor U10765 (N_10765,N_9823,N_10180);
nor U10766 (N_10766,N_9854,N_10277);
nand U10767 (N_10767,N_9979,N_9777);
and U10768 (N_10768,N_10443,N_10381);
nand U10769 (N_10769,N_10427,N_9917);
and U10770 (N_10770,N_9770,N_10008);
and U10771 (N_10771,N_10186,N_9994);
nor U10772 (N_10772,N_10055,N_10319);
and U10773 (N_10773,N_9751,N_10489);
and U10774 (N_10774,N_9865,N_9839);
or U10775 (N_10775,N_10108,N_9768);
and U10776 (N_10776,N_10103,N_9753);
nand U10777 (N_10777,N_10127,N_9963);
nor U10778 (N_10778,N_9951,N_9905);
nand U10779 (N_10779,N_10141,N_9980);
nand U10780 (N_10780,N_9991,N_10249);
and U10781 (N_10781,N_10121,N_10461);
nand U10782 (N_10782,N_10073,N_10391);
nand U10783 (N_10783,N_10195,N_10433);
xor U10784 (N_10784,N_10365,N_10019);
or U10785 (N_10785,N_9931,N_9789);
nand U10786 (N_10786,N_9859,N_9944);
nor U10787 (N_10787,N_10294,N_10432);
and U10788 (N_10788,N_10129,N_10455);
and U10789 (N_10789,N_10271,N_9995);
or U10790 (N_10790,N_9755,N_9845);
nand U10791 (N_10791,N_10337,N_10194);
nor U10792 (N_10792,N_10165,N_10360);
and U10793 (N_10793,N_10173,N_10177);
or U10794 (N_10794,N_10166,N_10295);
nor U10795 (N_10795,N_9797,N_10468);
or U10796 (N_10796,N_9787,N_9964);
and U10797 (N_10797,N_9970,N_9868);
xnor U10798 (N_10798,N_10029,N_10274);
and U10799 (N_10799,N_10077,N_10027);
or U10800 (N_10800,N_10351,N_9757);
nand U10801 (N_10801,N_10144,N_10111);
or U10802 (N_10802,N_10094,N_10306);
nor U10803 (N_10803,N_10081,N_9967);
and U10804 (N_10804,N_10423,N_10222);
nor U10805 (N_10805,N_10112,N_10348);
nor U10806 (N_10806,N_9825,N_9933);
or U10807 (N_10807,N_10041,N_10187);
nor U10808 (N_10808,N_10104,N_10471);
nand U10809 (N_10809,N_9893,N_9835);
nor U10810 (N_10810,N_9897,N_10476);
nand U10811 (N_10811,N_10317,N_9769);
nand U10812 (N_10812,N_9904,N_10488);
or U10813 (N_10813,N_10211,N_9943);
or U10814 (N_10814,N_10493,N_10192);
nand U10815 (N_10815,N_10414,N_10450);
nand U10816 (N_10816,N_9832,N_10431);
or U10817 (N_10817,N_10384,N_9792);
nor U10818 (N_10818,N_10006,N_10157);
nor U10819 (N_10819,N_9878,N_10233);
xnor U10820 (N_10820,N_10334,N_10494);
nand U10821 (N_10821,N_10232,N_9926);
or U10822 (N_10822,N_10301,N_10203);
or U10823 (N_10823,N_10028,N_10373);
and U10824 (N_10824,N_9817,N_9981);
xnor U10825 (N_10825,N_9938,N_10084);
nor U10826 (N_10826,N_10253,N_10367);
nor U10827 (N_10827,N_9922,N_10009);
nor U10828 (N_10828,N_10293,N_9908);
nor U10829 (N_10829,N_9774,N_10406);
nand U10830 (N_10830,N_9851,N_9871);
nor U10831 (N_10831,N_10486,N_9999);
xnor U10832 (N_10832,N_10324,N_10259);
and U10833 (N_10833,N_10161,N_9857);
or U10834 (N_10834,N_9791,N_10475);
or U10835 (N_10835,N_10339,N_10106);
nor U10836 (N_10836,N_10220,N_10185);
and U10837 (N_10837,N_10075,N_10007);
nor U10838 (N_10838,N_9984,N_10284);
nor U10839 (N_10839,N_9799,N_10243);
or U10840 (N_10840,N_10114,N_10430);
or U10841 (N_10841,N_10167,N_10045);
and U10842 (N_10842,N_10040,N_10413);
nand U10843 (N_10843,N_10258,N_10016);
or U10844 (N_10844,N_10392,N_10363);
and U10845 (N_10845,N_10477,N_10068);
nand U10846 (N_10846,N_10397,N_9822);
nand U10847 (N_10847,N_10285,N_9778);
or U10848 (N_10848,N_9786,N_10079);
or U10849 (N_10849,N_10089,N_10283);
or U10850 (N_10850,N_10163,N_10062);
nor U10851 (N_10851,N_10026,N_9914);
nor U10852 (N_10852,N_9783,N_9911);
xor U10853 (N_10853,N_9910,N_10070);
nor U10854 (N_10854,N_10340,N_10118);
nor U10855 (N_10855,N_9875,N_10305);
nor U10856 (N_10856,N_10320,N_10212);
and U10857 (N_10857,N_9863,N_9760);
nor U10858 (N_10858,N_9866,N_10467);
nor U10859 (N_10859,N_9829,N_10331);
nand U10860 (N_10860,N_10241,N_10321);
xor U10861 (N_10861,N_10462,N_10050);
nor U10862 (N_10862,N_10429,N_10409);
nor U10863 (N_10863,N_10083,N_9988);
xnor U10864 (N_10864,N_9841,N_10288);
nor U10865 (N_10865,N_10248,N_10444);
nand U10866 (N_10866,N_9808,N_10316);
nand U10867 (N_10867,N_9828,N_10496);
or U10868 (N_10868,N_9930,N_10013);
nand U10869 (N_10869,N_10412,N_10298);
and U10870 (N_10870,N_10216,N_9939);
or U10871 (N_10871,N_10149,N_10364);
and U10872 (N_10872,N_9960,N_10260);
and U10873 (N_10873,N_10048,N_9771);
and U10874 (N_10874,N_10034,N_9824);
or U10875 (N_10875,N_10416,N_10173);
and U10876 (N_10876,N_10277,N_9839);
and U10877 (N_10877,N_10336,N_10461);
nor U10878 (N_10878,N_9812,N_10045);
nor U10879 (N_10879,N_10223,N_9998);
or U10880 (N_10880,N_10319,N_10455);
nor U10881 (N_10881,N_10243,N_10065);
nand U10882 (N_10882,N_10080,N_10418);
and U10883 (N_10883,N_9752,N_10477);
nand U10884 (N_10884,N_10049,N_10184);
and U10885 (N_10885,N_9989,N_10052);
nand U10886 (N_10886,N_10263,N_9923);
nand U10887 (N_10887,N_10341,N_10130);
nor U10888 (N_10888,N_10440,N_10214);
xnor U10889 (N_10889,N_9969,N_10473);
nand U10890 (N_10890,N_10349,N_10371);
or U10891 (N_10891,N_9762,N_9960);
xor U10892 (N_10892,N_10340,N_10130);
nor U10893 (N_10893,N_10154,N_9750);
nor U10894 (N_10894,N_10339,N_10365);
and U10895 (N_10895,N_10285,N_10258);
nor U10896 (N_10896,N_10314,N_10128);
or U10897 (N_10897,N_9834,N_9870);
nor U10898 (N_10898,N_9935,N_10022);
or U10899 (N_10899,N_10003,N_9979);
or U10900 (N_10900,N_10253,N_10116);
xnor U10901 (N_10901,N_9789,N_9884);
and U10902 (N_10902,N_9783,N_10176);
nand U10903 (N_10903,N_10458,N_10325);
nand U10904 (N_10904,N_10437,N_10210);
nor U10905 (N_10905,N_9925,N_10446);
xor U10906 (N_10906,N_10119,N_10102);
nor U10907 (N_10907,N_10088,N_9950);
or U10908 (N_10908,N_10112,N_9826);
nand U10909 (N_10909,N_9780,N_10418);
and U10910 (N_10910,N_9829,N_10409);
or U10911 (N_10911,N_10386,N_10081);
nand U10912 (N_10912,N_10492,N_10043);
or U10913 (N_10913,N_9764,N_10032);
nand U10914 (N_10914,N_10066,N_10137);
nor U10915 (N_10915,N_10159,N_10051);
and U10916 (N_10916,N_10211,N_10253);
nor U10917 (N_10917,N_10220,N_10089);
nor U10918 (N_10918,N_9787,N_10481);
or U10919 (N_10919,N_9775,N_9861);
and U10920 (N_10920,N_10326,N_9971);
nor U10921 (N_10921,N_9785,N_9994);
nand U10922 (N_10922,N_10221,N_10290);
and U10923 (N_10923,N_9760,N_10176);
nor U10924 (N_10924,N_10116,N_10292);
nor U10925 (N_10925,N_10233,N_9765);
and U10926 (N_10926,N_9969,N_9853);
and U10927 (N_10927,N_10256,N_10359);
or U10928 (N_10928,N_10355,N_10357);
nor U10929 (N_10929,N_10499,N_9960);
nor U10930 (N_10930,N_9889,N_9940);
and U10931 (N_10931,N_10376,N_9787);
or U10932 (N_10932,N_9996,N_9921);
xor U10933 (N_10933,N_9973,N_10432);
or U10934 (N_10934,N_9980,N_10485);
or U10935 (N_10935,N_9941,N_10428);
or U10936 (N_10936,N_10159,N_10129);
nand U10937 (N_10937,N_10089,N_9971);
xor U10938 (N_10938,N_10443,N_9926);
and U10939 (N_10939,N_10208,N_9798);
or U10940 (N_10940,N_10400,N_10076);
or U10941 (N_10941,N_10477,N_10138);
and U10942 (N_10942,N_9853,N_10266);
nand U10943 (N_10943,N_9832,N_10007);
nand U10944 (N_10944,N_10320,N_10421);
nor U10945 (N_10945,N_10263,N_9765);
or U10946 (N_10946,N_10353,N_9762);
nor U10947 (N_10947,N_9956,N_9909);
or U10948 (N_10948,N_9803,N_9898);
nor U10949 (N_10949,N_9969,N_9813);
nand U10950 (N_10950,N_9758,N_10467);
xnor U10951 (N_10951,N_9887,N_10268);
and U10952 (N_10952,N_9880,N_10276);
nand U10953 (N_10953,N_10296,N_10179);
nand U10954 (N_10954,N_10244,N_9936);
or U10955 (N_10955,N_10066,N_10361);
and U10956 (N_10956,N_10149,N_9885);
nor U10957 (N_10957,N_10162,N_10161);
nand U10958 (N_10958,N_10084,N_10387);
nor U10959 (N_10959,N_9818,N_10410);
and U10960 (N_10960,N_9945,N_10242);
and U10961 (N_10961,N_10472,N_10073);
nand U10962 (N_10962,N_10435,N_10400);
nand U10963 (N_10963,N_9759,N_10249);
or U10964 (N_10964,N_10282,N_10478);
nand U10965 (N_10965,N_9944,N_10383);
nor U10966 (N_10966,N_9962,N_10262);
nand U10967 (N_10967,N_10479,N_9775);
or U10968 (N_10968,N_9979,N_10445);
nand U10969 (N_10969,N_10409,N_9968);
and U10970 (N_10970,N_10022,N_10439);
nor U10971 (N_10971,N_9897,N_10403);
nand U10972 (N_10972,N_10031,N_10163);
nor U10973 (N_10973,N_10148,N_10401);
and U10974 (N_10974,N_10271,N_10366);
xnor U10975 (N_10975,N_10191,N_9890);
and U10976 (N_10976,N_10223,N_10399);
xnor U10977 (N_10977,N_10288,N_9833);
and U10978 (N_10978,N_9916,N_10284);
and U10979 (N_10979,N_9752,N_10094);
and U10980 (N_10980,N_9865,N_10206);
nor U10981 (N_10981,N_10030,N_10136);
and U10982 (N_10982,N_10247,N_10140);
or U10983 (N_10983,N_10348,N_9931);
nand U10984 (N_10984,N_10250,N_10413);
and U10985 (N_10985,N_10348,N_9849);
nor U10986 (N_10986,N_10041,N_10042);
or U10987 (N_10987,N_10214,N_10054);
nor U10988 (N_10988,N_10299,N_10111);
nor U10989 (N_10989,N_9956,N_9960);
and U10990 (N_10990,N_9944,N_10250);
xnor U10991 (N_10991,N_10380,N_10454);
and U10992 (N_10992,N_10130,N_10215);
xnor U10993 (N_10993,N_9847,N_10499);
nor U10994 (N_10994,N_10443,N_9834);
nor U10995 (N_10995,N_10307,N_10097);
or U10996 (N_10996,N_9835,N_10178);
nor U10997 (N_10997,N_10421,N_9928);
nand U10998 (N_10998,N_9885,N_10272);
nand U10999 (N_10999,N_10139,N_10495);
or U11000 (N_11000,N_10347,N_9794);
and U11001 (N_11001,N_10144,N_10096);
and U11002 (N_11002,N_10172,N_9828);
or U11003 (N_11003,N_9903,N_10484);
and U11004 (N_11004,N_10318,N_10455);
and U11005 (N_11005,N_10349,N_10194);
or U11006 (N_11006,N_10092,N_10072);
and U11007 (N_11007,N_10218,N_10296);
nand U11008 (N_11008,N_10054,N_10429);
xor U11009 (N_11009,N_9837,N_10217);
nor U11010 (N_11010,N_10186,N_10431);
nor U11011 (N_11011,N_10450,N_10110);
nand U11012 (N_11012,N_10422,N_9957);
or U11013 (N_11013,N_9943,N_9867);
nor U11014 (N_11014,N_9920,N_10302);
nand U11015 (N_11015,N_9770,N_10486);
xnor U11016 (N_11016,N_10305,N_10394);
nand U11017 (N_11017,N_10092,N_10179);
and U11018 (N_11018,N_10051,N_10078);
or U11019 (N_11019,N_10022,N_10060);
or U11020 (N_11020,N_10226,N_9950);
nand U11021 (N_11021,N_10358,N_9844);
nor U11022 (N_11022,N_10025,N_9999);
and U11023 (N_11023,N_10431,N_9949);
nor U11024 (N_11024,N_9878,N_10115);
nand U11025 (N_11025,N_9998,N_10021);
nand U11026 (N_11026,N_10204,N_10449);
and U11027 (N_11027,N_10490,N_10248);
or U11028 (N_11028,N_10340,N_9953);
nand U11029 (N_11029,N_9800,N_10106);
nor U11030 (N_11030,N_10127,N_10142);
nand U11031 (N_11031,N_10052,N_9950);
nor U11032 (N_11032,N_9864,N_10167);
and U11033 (N_11033,N_9914,N_9949);
xnor U11034 (N_11034,N_10282,N_9827);
nand U11035 (N_11035,N_10462,N_10113);
nand U11036 (N_11036,N_10075,N_9837);
nor U11037 (N_11037,N_10171,N_10086);
nor U11038 (N_11038,N_10265,N_10050);
nor U11039 (N_11039,N_10132,N_10170);
xor U11040 (N_11040,N_10312,N_10389);
nand U11041 (N_11041,N_10436,N_9870);
and U11042 (N_11042,N_10394,N_10486);
nand U11043 (N_11043,N_10043,N_10088);
or U11044 (N_11044,N_10436,N_10181);
or U11045 (N_11045,N_10473,N_9843);
nor U11046 (N_11046,N_10378,N_10140);
nand U11047 (N_11047,N_10384,N_9793);
nand U11048 (N_11048,N_10264,N_10390);
xnor U11049 (N_11049,N_10158,N_9777);
or U11050 (N_11050,N_10359,N_10471);
and U11051 (N_11051,N_9870,N_9828);
or U11052 (N_11052,N_10471,N_10472);
or U11053 (N_11053,N_10321,N_10264);
nor U11054 (N_11054,N_10227,N_10162);
and U11055 (N_11055,N_10317,N_10391);
nand U11056 (N_11056,N_10471,N_10139);
nor U11057 (N_11057,N_10038,N_10491);
nand U11058 (N_11058,N_10381,N_10060);
nor U11059 (N_11059,N_10019,N_10062);
or U11060 (N_11060,N_10489,N_9843);
and U11061 (N_11061,N_10458,N_9776);
nand U11062 (N_11062,N_9827,N_10264);
nor U11063 (N_11063,N_10410,N_9765);
and U11064 (N_11064,N_9756,N_9761);
or U11065 (N_11065,N_9953,N_10079);
nor U11066 (N_11066,N_10462,N_10153);
or U11067 (N_11067,N_10153,N_9781);
nand U11068 (N_11068,N_9831,N_10476);
and U11069 (N_11069,N_10278,N_9763);
nand U11070 (N_11070,N_10261,N_10398);
or U11071 (N_11071,N_10382,N_10244);
nor U11072 (N_11072,N_10164,N_10380);
nor U11073 (N_11073,N_10306,N_9785);
nand U11074 (N_11074,N_10161,N_10310);
xor U11075 (N_11075,N_10259,N_9760);
and U11076 (N_11076,N_10051,N_9846);
nand U11077 (N_11077,N_10339,N_9752);
and U11078 (N_11078,N_9899,N_10057);
xor U11079 (N_11079,N_10257,N_10390);
or U11080 (N_11080,N_10219,N_9929);
nor U11081 (N_11081,N_10058,N_10182);
nand U11082 (N_11082,N_10066,N_10261);
nor U11083 (N_11083,N_10052,N_10389);
and U11084 (N_11084,N_10170,N_9772);
nor U11085 (N_11085,N_10216,N_10005);
or U11086 (N_11086,N_10374,N_9885);
nand U11087 (N_11087,N_10053,N_9762);
and U11088 (N_11088,N_9895,N_10363);
or U11089 (N_11089,N_10046,N_9798);
or U11090 (N_11090,N_10183,N_10359);
or U11091 (N_11091,N_9762,N_10047);
nor U11092 (N_11092,N_10307,N_10353);
xnor U11093 (N_11093,N_10080,N_10268);
and U11094 (N_11094,N_10388,N_9947);
and U11095 (N_11095,N_9846,N_9924);
nor U11096 (N_11096,N_9880,N_10370);
nor U11097 (N_11097,N_10062,N_9801);
and U11098 (N_11098,N_10085,N_10361);
nor U11099 (N_11099,N_10140,N_10239);
and U11100 (N_11100,N_9805,N_9817);
nand U11101 (N_11101,N_9947,N_10015);
or U11102 (N_11102,N_10363,N_9930);
nand U11103 (N_11103,N_9858,N_10061);
or U11104 (N_11104,N_10339,N_9822);
and U11105 (N_11105,N_10161,N_9998);
or U11106 (N_11106,N_10436,N_9774);
nor U11107 (N_11107,N_9996,N_10422);
nand U11108 (N_11108,N_10338,N_10464);
or U11109 (N_11109,N_10419,N_10274);
nor U11110 (N_11110,N_9877,N_10141);
nor U11111 (N_11111,N_10378,N_9932);
nor U11112 (N_11112,N_10061,N_10443);
and U11113 (N_11113,N_9824,N_9847);
and U11114 (N_11114,N_10218,N_10124);
xnor U11115 (N_11115,N_10009,N_10167);
and U11116 (N_11116,N_9793,N_10281);
nand U11117 (N_11117,N_10105,N_9957);
and U11118 (N_11118,N_9811,N_9872);
nand U11119 (N_11119,N_10374,N_10376);
and U11120 (N_11120,N_9880,N_10389);
nand U11121 (N_11121,N_10455,N_10499);
xnor U11122 (N_11122,N_9763,N_9798);
and U11123 (N_11123,N_9923,N_10303);
or U11124 (N_11124,N_10172,N_10247);
or U11125 (N_11125,N_10308,N_10207);
nand U11126 (N_11126,N_9972,N_10042);
and U11127 (N_11127,N_10139,N_10229);
xor U11128 (N_11128,N_9940,N_9922);
and U11129 (N_11129,N_10013,N_10257);
nand U11130 (N_11130,N_9851,N_10363);
nor U11131 (N_11131,N_9896,N_9983);
or U11132 (N_11132,N_10377,N_10479);
and U11133 (N_11133,N_10220,N_10460);
nand U11134 (N_11134,N_10250,N_10225);
and U11135 (N_11135,N_10410,N_9966);
nand U11136 (N_11136,N_10339,N_10248);
and U11137 (N_11137,N_9839,N_10388);
and U11138 (N_11138,N_10197,N_9886);
and U11139 (N_11139,N_10499,N_9838);
and U11140 (N_11140,N_9894,N_9836);
nor U11141 (N_11141,N_9988,N_10244);
and U11142 (N_11142,N_10162,N_10120);
nand U11143 (N_11143,N_9894,N_9838);
nand U11144 (N_11144,N_9890,N_9913);
nor U11145 (N_11145,N_10176,N_10305);
nor U11146 (N_11146,N_10302,N_10044);
or U11147 (N_11147,N_10061,N_9802);
nor U11148 (N_11148,N_10382,N_10282);
nor U11149 (N_11149,N_9973,N_10095);
nor U11150 (N_11150,N_9921,N_10081);
or U11151 (N_11151,N_10398,N_10155);
nor U11152 (N_11152,N_10436,N_10358);
or U11153 (N_11153,N_10345,N_10374);
and U11154 (N_11154,N_9991,N_9781);
or U11155 (N_11155,N_9972,N_10023);
nor U11156 (N_11156,N_10331,N_10108);
nand U11157 (N_11157,N_10022,N_10256);
nor U11158 (N_11158,N_10233,N_10225);
or U11159 (N_11159,N_9921,N_10389);
nand U11160 (N_11160,N_10493,N_9810);
or U11161 (N_11161,N_10006,N_9942);
nor U11162 (N_11162,N_10126,N_10035);
nand U11163 (N_11163,N_10220,N_9782);
nor U11164 (N_11164,N_9867,N_10075);
and U11165 (N_11165,N_10330,N_10381);
and U11166 (N_11166,N_9859,N_10332);
nand U11167 (N_11167,N_9918,N_10483);
or U11168 (N_11168,N_10435,N_10446);
nor U11169 (N_11169,N_10344,N_10091);
and U11170 (N_11170,N_10330,N_10282);
nor U11171 (N_11171,N_10400,N_10118);
or U11172 (N_11172,N_10124,N_9884);
and U11173 (N_11173,N_10009,N_9839);
nor U11174 (N_11174,N_10408,N_9871);
nand U11175 (N_11175,N_10357,N_9927);
nand U11176 (N_11176,N_9881,N_9852);
or U11177 (N_11177,N_9941,N_10398);
nor U11178 (N_11178,N_10257,N_10012);
nand U11179 (N_11179,N_9824,N_10021);
nand U11180 (N_11180,N_9785,N_10280);
nor U11181 (N_11181,N_10352,N_10163);
and U11182 (N_11182,N_10442,N_10136);
or U11183 (N_11183,N_10135,N_10123);
nor U11184 (N_11184,N_10389,N_10370);
and U11185 (N_11185,N_10205,N_10448);
and U11186 (N_11186,N_9884,N_10148);
nor U11187 (N_11187,N_10222,N_9762);
nand U11188 (N_11188,N_10370,N_9971);
or U11189 (N_11189,N_10304,N_10325);
nor U11190 (N_11190,N_9758,N_10163);
xnor U11191 (N_11191,N_10240,N_10211);
and U11192 (N_11192,N_10363,N_9952);
nand U11193 (N_11193,N_10425,N_10436);
nor U11194 (N_11194,N_9792,N_10258);
or U11195 (N_11195,N_10147,N_10245);
or U11196 (N_11196,N_9890,N_10294);
nor U11197 (N_11197,N_10034,N_10133);
and U11198 (N_11198,N_10275,N_9792);
or U11199 (N_11199,N_10106,N_10107);
nand U11200 (N_11200,N_10387,N_10122);
xor U11201 (N_11201,N_9850,N_10436);
nand U11202 (N_11202,N_10105,N_10086);
and U11203 (N_11203,N_9763,N_10435);
xnor U11204 (N_11204,N_10411,N_9921);
nand U11205 (N_11205,N_9849,N_10098);
nand U11206 (N_11206,N_10093,N_9958);
and U11207 (N_11207,N_9798,N_10381);
nand U11208 (N_11208,N_9951,N_10465);
nand U11209 (N_11209,N_9774,N_10126);
or U11210 (N_11210,N_10128,N_10493);
nor U11211 (N_11211,N_9923,N_10106);
or U11212 (N_11212,N_10328,N_9935);
nor U11213 (N_11213,N_9762,N_9894);
nor U11214 (N_11214,N_10275,N_9765);
nand U11215 (N_11215,N_10448,N_9804);
nand U11216 (N_11216,N_10231,N_10345);
and U11217 (N_11217,N_9947,N_9792);
nor U11218 (N_11218,N_10047,N_9910);
nor U11219 (N_11219,N_9785,N_9963);
nor U11220 (N_11220,N_10309,N_9875);
nand U11221 (N_11221,N_10257,N_10441);
xnor U11222 (N_11222,N_10318,N_9775);
nand U11223 (N_11223,N_9866,N_10151);
nand U11224 (N_11224,N_10074,N_10172);
or U11225 (N_11225,N_10410,N_10491);
nand U11226 (N_11226,N_9948,N_10264);
and U11227 (N_11227,N_9794,N_10099);
nand U11228 (N_11228,N_10081,N_10230);
nor U11229 (N_11229,N_9832,N_9787);
nand U11230 (N_11230,N_9753,N_10276);
nand U11231 (N_11231,N_9954,N_9851);
nor U11232 (N_11232,N_9762,N_9764);
and U11233 (N_11233,N_10061,N_10038);
or U11234 (N_11234,N_10428,N_10360);
or U11235 (N_11235,N_9998,N_10119);
nand U11236 (N_11236,N_9924,N_10061);
xor U11237 (N_11237,N_10494,N_10251);
nand U11238 (N_11238,N_9940,N_10125);
nor U11239 (N_11239,N_10168,N_10062);
nor U11240 (N_11240,N_10489,N_10235);
nor U11241 (N_11241,N_9875,N_10038);
nand U11242 (N_11242,N_9938,N_9978);
or U11243 (N_11243,N_10473,N_10080);
nor U11244 (N_11244,N_10276,N_10198);
or U11245 (N_11245,N_9791,N_10460);
and U11246 (N_11246,N_10250,N_10121);
nand U11247 (N_11247,N_10154,N_9805);
nor U11248 (N_11248,N_10258,N_10379);
and U11249 (N_11249,N_10083,N_9977);
and U11250 (N_11250,N_10850,N_10929);
and U11251 (N_11251,N_10551,N_11072);
nor U11252 (N_11252,N_11023,N_11150);
nor U11253 (N_11253,N_11065,N_10859);
nor U11254 (N_11254,N_10677,N_11070);
nand U11255 (N_11255,N_10982,N_10856);
or U11256 (N_11256,N_11112,N_10963);
nor U11257 (N_11257,N_10645,N_10699);
nand U11258 (N_11258,N_10997,N_10989);
nand U11259 (N_11259,N_11044,N_10832);
or U11260 (N_11260,N_10539,N_10580);
xor U11261 (N_11261,N_10570,N_10624);
nor U11262 (N_11262,N_10992,N_10755);
nor U11263 (N_11263,N_11181,N_10999);
or U11264 (N_11264,N_10939,N_10904);
nand U11265 (N_11265,N_10796,N_10512);
nand U11266 (N_11266,N_10771,N_11013);
or U11267 (N_11267,N_11046,N_11061);
and U11268 (N_11268,N_11184,N_10530);
or U11269 (N_11269,N_10778,N_10532);
and U11270 (N_11270,N_10650,N_11050);
xnor U11271 (N_11271,N_10791,N_10646);
or U11272 (N_11272,N_10502,N_11141);
or U11273 (N_11273,N_11094,N_10666);
nand U11274 (N_11274,N_11039,N_11106);
or U11275 (N_11275,N_10739,N_10990);
xnor U11276 (N_11276,N_10901,N_11178);
or U11277 (N_11277,N_11096,N_10880);
nor U11278 (N_11278,N_10720,N_10722);
nand U11279 (N_11279,N_11155,N_10566);
nand U11280 (N_11280,N_11245,N_11089);
nand U11281 (N_11281,N_10634,N_11152);
and U11282 (N_11282,N_10881,N_10806);
or U11283 (N_11283,N_10531,N_11228);
xor U11284 (N_11284,N_10770,N_11071);
or U11285 (N_11285,N_11002,N_11114);
nand U11286 (N_11286,N_10785,N_11129);
nand U11287 (N_11287,N_10697,N_11135);
xor U11288 (N_11288,N_11171,N_11032);
nand U11289 (N_11289,N_11220,N_10775);
and U11290 (N_11290,N_10964,N_10648);
xnor U11291 (N_11291,N_10729,N_10845);
xnor U11292 (N_11292,N_11001,N_10702);
nor U11293 (N_11293,N_11248,N_10550);
nand U11294 (N_11294,N_10657,N_11077);
or U11295 (N_11295,N_10979,N_11103);
nor U11296 (N_11296,N_10540,N_10672);
nor U11297 (N_11297,N_10740,N_11014);
nand U11298 (N_11298,N_10841,N_10782);
nor U11299 (N_11299,N_10886,N_10520);
or U11300 (N_11300,N_10756,N_11237);
nand U11301 (N_11301,N_11052,N_10581);
xor U11302 (N_11302,N_11203,N_10575);
xor U11303 (N_11303,N_10994,N_11038);
or U11304 (N_11304,N_11239,N_10734);
or U11305 (N_11305,N_10553,N_11127);
nand U11306 (N_11306,N_11108,N_11067);
nor U11307 (N_11307,N_10565,N_11175);
nand U11308 (N_11308,N_10829,N_10714);
xor U11309 (N_11309,N_11113,N_11147);
or U11310 (N_11310,N_10956,N_11043);
nand U11311 (N_11311,N_10940,N_11012);
or U11312 (N_11312,N_10589,N_11142);
or U11313 (N_11313,N_10944,N_10847);
nand U11314 (N_11314,N_10693,N_10788);
or U11315 (N_11315,N_11185,N_11231);
or U11316 (N_11316,N_10594,N_10690);
nor U11317 (N_11317,N_11095,N_10554);
nor U11318 (N_11318,N_10733,N_10779);
or U11319 (N_11319,N_10737,N_10597);
nor U11320 (N_11320,N_10749,N_10644);
xor U11321 (N_11321,N_10925,N_11194);
xor U11322 (N_11322,N_11172,N_11207);
nor U11323 (N_11323,N_10613,N_10932);
or U11324 (N_11324,N_10958,N_10680);
or U11325 (N_11325,N_10808,N_10614);
and U11326 (N_11326,N_11230,N_10849);
and U11327 (N_11327,N_11160,N_10916);
nand U11328 (N_11328,N_10833,N_11235);
nand U11329 (N_11329,N_10587,N_11057);
nand U11330 (N_11330,N_11020,N_10687);
nand U11331 (N_11331,N_11030,N_10935);
nor U11332 (N_11332,N_11107,N_10518);
nor U11333 (N_11333,N_11056,N_11166);
xnor U11334 (N_11334,N_11022,N_11078);
nor U11335 (N_11335,N_10821,N_10988);
nor U11336 (N_11336,N_11041,N_11085);
nand U11337 (N_11337,N_10781,N_11005);
nand U11338 (N_11338,N_10662,N_11159);
nor U11339 (N_11339,N_10574,N_11176);
and U11340 (N_11340,N_10688,N_11051);
or U11341 (N_11341,N_11027,N_11145);
or U11342 (N_11342,N_10804,N_11092);
or U11343 (N_11343,N_10941,N_10567);
and U11344 (N_11344,N_10758,N_10920);
and U11345 (N_11345,N_10903,N_10834);
and U11346 (N_11346,N_10899,N_10772);
nand U11347 (N_11347,N_10857,N_10652);
nor U11348 (N_11348,N_10838,N_11111);
nand U11349 (N_11349,N_10913,N_10765);
nand U11350 (N_11350,N_10534,N_10840);
or U11351 (N_11351,N_10759,N_10651);
and U11352 (N_11352,N_10768,N_10736);
nor U11353 (N_11353,N_10789,N_10527);
nor U11354 (N_11354,N_11209,N_10555);
nor U11355 (N_11355,N_11211,N_10603);
nor U11356 (N_11356,N_11074,N_10980);
nor U11357 (N_11357,N_10953,N_10584);
or U11358 (N_11358,N_11125,N_10908);
and U11359 (N_11359,N_11153,N_10757);
or U11360 (N_11360,N_10800,N_10748);
or U11361 (N_11361,N_11060,N_10893);
nand U11362 (N_11362,N_10607,N_10952);
nor U11363 (N_11363,N_10577,N_10503);
and U11364 (N_11364,N_11218,N_11162);
and U11365 (N_11365,N_11164,N_10541);
nand U11366 (N_11366,N_10767,N_11109);
nand U11367 (N_11367,N_10810,N_11163);
nor U11368 (N_11368,N_11242,N_10803);
and U11369 (N_11369,N_10544,N_10854);
or U11370 (N_11370,N_10728,N_10822);
nor U11371 (N_11371,N_10605,N_10762);
and U11372 (N_11372,N_10863,N_11182);
nand U11373 (N_11373,N_10716,N_10891);
or U11374 (N_11374,N_10787,N_10723);
nand U11375 (N_11375,N_11206,N_10816);
and U11376 (N_11376,N_10921,N_10561);
nand U11377 (N_11377,N_10855,N_10609);
or U11378 (N_11378,N_10673,N_10717);
nand U11379 (N_11379,N_10704,N_11091);
nand U11380 (N_11380,N_11024,N_10922);
or U11381 (N_11381,N_11167,N_11130);
nor U11382 (N_11382,N_11008,N_10823);
or U11383 (N_11383,N_10970,N_11177);
nand U11384 (N_11384,N_10814,N_11154);
or U11385 (N_11385,N_10815,N_10637);
nor U11386 (N_11386,N_10996,N_10504);
and U11387 (N_11387,N_10725,N_11034);
and U11388 (N_11388,N_10967,N_10957);
nor U11389 (N_11389,N_11186,N_10844);
nor U11390 (N_11390,N_10851,N_10521);
or U11391 (N_11391,N_10861,N_10627);
xnor U11392 (N_11392,N_10546,N_11204);
nand U11393 (N_11393,N_10514,N_11007);
nor U11394 (N_11394,N_10835,N_10689);
nand U11395 (N_11395,N_11139,N_10852);
nand U11396 (N_11396,N_11165,N_10978);
nor U11397 (N_11397,N_11076,N_10578);
nor U11398 (N_11398,N_10926,N_10965);
nand U11399 (N_11399,N_10865,N_10593);
and U11400 (N_11400,N_10612,N_11009);
or U11401 (N_11401,N_10653,N_10793);
or U11402 (N_11402,N_10710,N_10905);
nor U11403 (N_11403,N_10522,N_11118);
and U11404 (N_11404,N_10786,N_10910);
nand U11405 (N_11405,N_10862,N_11063);
or U11406 (N_11406,N_10985,N_11098);
or U11407 (N_11407,N_11033,N_10776);
or U11408 (N_11408,N_10611,N_10811);
nor U11409 (N_11409,N_10911,N_10703);
xnor U11410 (N_11410,N_10632,N_10515);
and U11411 (N_11411,N_10797,N_10831);
or U11412 (N_11412,N_10820,N_10635);
nor U11413 (N_11413,N_10509,N_11210);
xnor U11414 (N_11414,N_10727,N_10643);
nor U11415 (N_11415,N_10516,N_11244);
nor U11416 (N_11416,N_10602,N_10558);
nand U11417 (N_11417,N_10973,N_10507);
nor U11418 (N_11418,N_10508,N_10706);
or U11419 (N_11419,N_10638,N_10827);
xnor U11420 (N_11420,N_10933,N_10528);
and U11421 (N_11421,N_10923,N_11062);
nor U11422 (N_11422,N_10713,N_11080);
xnor U11423 (N_11423,N_10513,N_10930);
nand U11424 (N_11424,N_10919,N_10542);
or U11425 (N_11425,N_11031,N_10887);
or U11426 (N_11426,N_11240,N_10735);
and U11427 (N_11427,N_11227,N_11003);
nor U11428 (N_11428,N_10655,N_11134);
nor U11429 (N_11429,N_10981,N_10897);
and U11430 (N_11430,N_10525,N_10912);
and U11431 (N_11431,N_11156,N_11119);
or U11432 (N_11432,N_10694,N_11083);
nor U11433 (N_11433,N_10777,N_11081);
nor U11434 (N_11434,N_11201,N_10871);
nor U11435 (N_11435,N_11016,N_10962);
nor U11436 (N_11436,N_10890,N_10568);
and U11437 (N_11437,N_10585,N_10548);
nor U11438 (N_11438,N_11102,N_10661);
nand U11439 (N_11439,N_10902,N_10701);
nor U11440 (N_11440,N_10595,N_11213);
and U11441 (N_11441,N_10617,N_10937);
or U11442 (N_11442,N_10681,N_11126);
and U11443 (N_11443,N_10591,N_11053);
and U11444 (N_11444,N_11199,N_11088);
and U11445 (N_11445,N_11226,N_10676);
nand U11446 (N_11446,N_10642,N_10959);
and U11447 (N_11447,N_11087,N_11028);
or U11448 (N_11448,N_11232,N_11138);
or U11449 (N_11449,N_10885,N_10761);
or U11450 (N_11450,N_10828,N_11189);
nor U11451 (N_11451,N_11058,N_10955);
or U11452 (N_11452,N_11011,N_10600);
or U11453 (N_11453,N_10543,N_10741);
nor U11454 (N_11454,N_10836,N_10631);
and U11455 (N_11455,N_10560,N_10914);
nand U11456 (N_11456,N_10623,N_11086);
and U11457 (N_11457,N_10895,N_10692);
and U11458 (N_11458,N_10524,N_10569);
nor U11459 (N_11459,N_10711,N_10984);
nor U11460 (N_11460,N_10620,N_10685);
or U11461 (N_11461,N_11068,N_11191);
nand U11462 (N_11462,N_11040,N_10817);
and U11463 (N_11463,N_10691,N_10715);
and U11464 (N_11464,N_10819,N_11148);
and U11465 (N_11465,N_10742,N_11122);
nand U11466 (N_11466,N_11222,N_11132);
nor U11467 (N_11467,N_10869,N_11223);
nand U11468 (N_11468,N_10529,N_11158);
or U11469 (N_11469,N_10995,N_10824);
and U11470 (N_11470,N_10658,N_10698);
nor U11471 (N_11471,N_10738,N_11133);
nand U11472 (N_11472,N_10971,N_11174);
or U11473 (N_11473,N_10807,N_10679);
nor U11474 (N_11474,N_11249,N_11079);
nor U11475 (N_11475,N_10745,N_10928);
and U11476 (N_11476,N_10876,N_11090);
nand U11477 (N_11477,N_10942,N_10889);
and U11478 (N_11478,N_10538,N_11198);
or U11479 (N_11479,N_10654,N_10573);
and U11480 (N_11480,N_11173,N_10860);
or U11481 (N_11481,N_11208,N_10976);
xor U11482 (N_11482,N_10667,N_11042);
or U11483 (N_11483,N_10754,N_10721);
and U11484 (N_11484,N_10682,N_10906);
nor U11485 (N_11485,N_10946,N_11029);
nor U11486 (N_11486,N_10536,N_10559);
nand U11487 (N_11487,N_10760,N_10802);
nor U11488 (N_11488,N_10991,N_10986);
and U11489 (N_11489,N_11202,N_10874);
nor U11490 (N_11490,N_10656,N_11214);
xnor U11491 (N_11491,N_10830,N_11116);
xor U11492 (N_11492,N_10545,N_11017);
or U11493 (N_11493,N_10664,N_11059);
or U11494 (N_11494,N_10647,N_11151);
nor U11495 (N_11495,N_10630,N_10663);
nand U11496 (N_11496,N_10948,N_10752);
nand U11497 (N_11497,N_10795,N_10537);
nand U11498 (N_11498,N_10763,N_10974);
nor U11499 (N_11499,N_10696,N_10853);
nand U11500 (N_11500,N_10608,N_11128);
and U11501 (N_11501,N_10780,N_11161);
or U11502 (N_11502,N_10649,N_10858);
nor U11503 (N_11503,N_10882,N_11019);
or U11504 (N_11504,N_10628,N_11149);
or U11505 (N_11505,N_10724,N_11136);
nor U11506 (N_11506,N_10812,N_10619);
and U11507 (N_11507,N_11246,N_10511);
and U11508 (N_11508,N_10883,N_11015);
nor U11509 (N_11509,N_10626,N_10907);
and U11510 (N_11510,N_10671,N_10753);
or U11511 (N_11511,N_10938,N_11247);
nor U11512 (N_11512,N_11110,N_11004);
or U11513 (N_11513,N_10764,N_10813);
nor U11514 (N_11514,N_10870,N_11236);
nor U11515 (N_11515,N_10535,N_11121);
or U11516 (N_11516,N_11216,N_10888);
and U11517 (N_11517,N_11099,N_11073);
or U11518 (N_11518,N_10506,N_10934);
or U11519 (N_11519,N_10500,N_11075);
and U11520 (N_11520,N_10894,N_11105);
nand U11521 (N_11521,N_11018,N_10563);
or U11522 (N_11522,N_10629,N_11234);
or U11523 (N_11523,N_10927,N_11026);
nor U11524 (N_11524,N_11010,N_10968);
and U11525 (N_11525,N_11193,N_10571);
nor U11526 (N_11526,N_10879,N_10826);
nand U11527 (N_11527,N_11205,N_11233);
xnor U11528 (N_11528,N_10665,N_10798);
nand U11529 (N_11529,N_10625,N_10750);
nand U11530 (N_11530,N_10640,N_10809);
and U11531 (N_11531,N_10588,N_11225);
nand U11532 (N_11532,N_10872,N_10659);
or U11533 (N_11533,N_11143,N_11082);
or U11534 (N_11534,N_10825,N_10866);
or U11535 (N_11535,N_10744,N_10517);
and U11536 (N_11536,N_10726,N_11243);
or U11537 (N_11537,N_10949,N_10633);
nor U11538 (N_11538,N_10839,N_11192);
or U11539 (N_11539,N_11229,N_11047);
and U11540 (N_11540,N_10868,N_10562);
and U11541 (N_11541,N_10526,N_10719);
nand U11542 (N_11542,N_10686,N_11049);
and U11543 (N_11543,N_11157,N_11037);
nand U11544 (N_11544,N_11115,N_10945);
or U11545 (N_11545,N_11212,N_10572);
nor U11546 (N_11546,N_10792,N_11195);
or U11547 (N_11547,N_10936,N_10805);
and U11548 (N_11548,N_10900,N_10684);
or U11549 (N_11549,N_10966,N_10732);
or U11550 (N_11550,N_11170,N_11224);
and U11551 (N_11551,N_11100,N_10975);
nor U11552 (N_11552,N_10843,N_10769);
and U11553 (N_11553,N_10898,N_11146);
and U11554 (N_11554,N_10917,N_10924);
nor U11555 (N_11555,N_11196,N_10993);
and U11556 (N_11556,N_11124,N_10877);
xor U11557 (N_11557,N_10718,N_10751);
and U11558 (N_11558,N_11101,N_10896);
nand U11559 (N_11559,N_10873,N_11179);
or U11560 (N_11560,N_10675,N_10700);
nand U11561 (N_11561,N_10641,N_11217);
nand U11562 (N_11562,N_11131,N_10766);
and U11563 (N_11563,N_11221,N_10519);
and U11564 (N_11564,N_11180,N_10998);
nand U11565 (N_11565,N_11021,N_10954);
nand U11566 (N_11566,N_11006,N_10712);
and U11567 (N_11567,N_10818,N_10969);
nand U11568 (N_11568,N_10576,N_11048);
and U11569 (N_11569,N_11120,N_10616);
and U11570 (N_11570,N_11140,N_11035);
nor U11571 (N_11571,N_10943,N_10909);
and U11572 (N_11572,N_11117,N_10884);
nand U11573 (N_11573,N_11000,N_10582);
or U11574 (N_11574,N_10864,N_10784);
and U11575 (N_11575,N_11187,N_11097);
nand U11576 (N_11576,N_10557,N_10552);
xor U11577 (N_11577,N_10583,N_10556);
nand U11578 (N_11578,N_10615,N_10730);
nor U11579 (N_11579,N_10950,N_10794);
nor U11580 (N_11580,N_10639,N_11241);
and U11581 (N_11581,N_10878,N_11036);
or U11582 (N_11582,N_10621,N_11168);
nand U11583 (N_11583,N_10695,N_10579);
and U11584 (N_11584,N_10983,N_10915);
nand U11585 (N_11585,N_10601,N_10783);
nand U11586 (N_11586,N_10708,N_11183);
nor U11587 (N_11587,N_11054,N_10842);
and U11588 (N_11588,N_10972,N_10731);
nor U11589 (N_11589,N_11025,N_10747);
nor U11590 (N_11590,N_11093,N_11064);
and U11591 (N_11591,N_10669,N_10707);
nor U11592 (N_11592,N_10848,N_10564);
nand U11593 (N_11593,N_10668,N_10678);
nor U11594 (N_11594,N_10590,N_10918);
nand U11595 (N_11595,N_10505,N_10596);
nand U11596 (N_11596,N_10799,N_10867);
or U11597 (N_11597,N_10947,N_10961);
nand U11598 (N_11598,N_10846,N_10746);
nand U11599 (N_11599,N_10592,N_10604);
or U11600 (N_11600,N_10773,N_11104);
and U11601 (N_11601,N_10523,N_11169);
or U11602 (N_11602,N_10533,N_10683);
and U11603 (N_11603,N_11238,N_11084);
nor U11604 (N_11604,N_10951,N_10549);
or U11605 (N_11605,N_11137,N_10960);
nor U11606 (N_11606,N_10705,N_10774);
or U11607 (N_11607,N_10547,N_11123);
nand U11608 (N_11608,N_11066,N_11055);
and U11609 (N_11609,N_10837,N_10674);
and U11610 (N_11610,N_10606,N_11144);
nand U11611 (N_11611,N_10618,N_10743);
nand U11612 (N_11612,N_10610,N_10875);
nand U11613 (N_11613,N_11069,N_10987);
and U11614 (N_11614,N_10977,N_10660);
nor U11615 (N_11615,N_10622,N_10790);
nand U11616 (N_11616,N_11215,N_10501);
or U11617 (N_11617,N_10636,N_10670);
nor U11618 (N_11618,N_11197,N_10510);
nand U11619 (N_11619,N_10892,N_10598);
nand U11620 (N_11620,N_10586,N_10931);
nand U11621 (N_11621,N_11190,N_11188);
or U11622 (N_11622,N_10801,N_11200);
xor U11623 (N_11623,N_11045,N_10599);
and U11624 (N_11624,N_11219,N_10709);
and U11625 (N_11625,N_11023,N_10978);
and U11626 (N_11626,N_10843,N_11054);
nand U11627 (N_11627,N_10666,N_11041);
xnor U11628 (N_11628,N_10668,N_10854);
and U11629 (N_11629,N_11064,N_11033);
or U11630 (N_11630,N_10628,N_10865);
nand U11631 (N_11631,N_11120,N_11243);
nand U11632 (N_11632,N_10936,N_11048);
nand U11633 (N_11633,N_11023,N_10587);
nor U11634 (N_11634,N_10883,N_10607);
or U11635 (N_11635,N_10665,N_11137);
xor U11636 (N_11636,N_10575,N_11174);
nand U11637 (N_11637,N_10613,N_10632);
and U11638 (N_11638,N_11143,N_10545);
and U11639 (N_11639,N_10685,N_10768);
and U11640 (N_11640,N_11046,N_10701);
xnor U11641 (N_11641,N_10606,N_10743);
nand U11642 (N_11642,N_11001,N_10827);
nor U11643 (N_11643,N_11211,N_10690);
nor U11644 (N_11644,N_10783,N_11194);
nand U11645 (N_11645,N_11079,N_10709);
nor U11646 (N_11646,N_10649,N_11108);
nand U11647 (N_11647,N_10948,N_10865);
nor U11648 (N_11648,N_10958,N_10626);
or U11649 (N_11649,N_10508,N_11172);
and U11650 (N_11650,N_10801,N_10929);
nand U11651 (N_11651,N_11155,N_10949);
or U11652 (N_11652,N_10768,N_11090);
or U11653 (N_11653,N_10758,N_11099);
nand U11654 (N_11654,N_11075,N_11170);
xor U11655 (N_11655,N_10850,N_11118);
nand U11656 (N_11656,N_10928,N_10656);
and U11657 (N_11657,N_10810,N_10805);
or U11658 (N_11658,N_10936,N_10669);
or U11659 (N_11659,N_10970,N_11215);
nor U11660 (N_11660,N_10653,N_11022);
nor U11661 (N_11661,N_10513,N_10627);
and U11662 (N_11662,N_10757,N_11202);
and U11663 (N_11663,N_10781,N_10871);
xor U11664 (N_11664,N_11153,N_10856);
nor U11665 (N_11665,N_10649,N_11202);
or U11666 (N_11666,N_11236,N_11107);
nor U11667 (N_11667,N_11018,N_10628);
nor U11668 (N_11668,N_10640,N_10758);
nand U11669 (N_11669,N_10537,N_10880);
nand U11670 (N_11670,N_10740,N_11228);
nand U11671 (N_11671,N_10565,N_10563);
nor U11672 (N_11672,N_10951,N_10901);
or U11673 (N_11673,N_11151,N_10776);
nand U11674 (N_11674,N_10570,N_10917);
or U11675 (N_11675,N_11163,N_10833);
nand U11676 (N_11676,N_11133,N_10576);
nor U11677 (N_11677,N_10522,N_11179);
nand U11678 (N_11678,N_10959,N_10685);
xor U11679 (N_11679,N_11162,N_10539);
xor U11680 (N_11680,N_11045,N_11064);
and U11681 (N_11681,N_10680,N_10798);
and U11682 (N_11682,N_10569,N_10618);
nand U11683 (N_11683,N_10816,N_11079);
nand U11684 (N_11684,N_10563,N_10901);
or U11685 (N_11685,N_11208,N_11215);
and U11686 (N_11686,N_11030,N_10500);
and U11687 (N_11687,N_11126,N_10694);
or U11688 (N_11688,N_11069,N_11149);
and U11689 (N_11689,N_10552,N_11117);
or U11690 (N_11690,N_10777,N_10595);
nor U11691 (N_11691,N_10921,N_10692);
nand U11692 (N_11692,N_10508,N_10875);
nand U11693 (N_11693,N_10895,N_11171);
and U11694 (N_11694,N_10968,N_10755);
or U11695 (N_11695,N_10689,N_11068);
nand U11696 (N_11696,N_10556,N_10742);
nand U11697 (N_11697,N_10740,N_11002);
nor U11698 (N_11698,N_10734,N_10527);
nor U11699 (N_11699,N_10778,N_10534);
nand U11700 (N_11700,N_11215,N_10801);
nor U11701 (N_11701,N_10513,N_10551);
nand U11702 (N_11702,N_11148,N_10962);
or U11703 (N_11703,N_10519,N_10647);
nand U11704 (N_11704,N_10531,N_10895);
or U11705 (N_11705,N_11216,N_10783);
nor U11706 (N_11706,N_11246,N_11104);
or U11707 (N_11707,N_11246,N_11160);
xor U11708 (N_11708,N_10629,N_11031);
and U11709 (N_11709,N_11137,N_11148);
or U11710 (N_11710,N_10642,N_10863);
or U11711 (N_11711,N_10830,N_10533);
and U11712 (N_11712,N_10783,N_11025);
xnor U11713 (N_11713,N_10860,N_11045);
nand U11714 (N_11714,N_10951,N_10562);
nor U11715 (N_11715,N_10855,N_10949);
or U11716 (N_11716,N_10668,N_11066);
nand U11717 (N_11717,N_10890,N_10616);
or U11718 (N_11718,N_10823,N_10907);
and U11719 (N_11719,N_11212,N_10873);
nand U11720 (N_11720,N_10689,N_10658);
nand U11721 (N_11721,N_10931,N_11168);
and U11722 (N_11722,N_11110,N_11031);
nor U11723 (N_11723,N_11195,N_10865);
or U11724 (N_11724,N_11138,N_11024);
or U11725 (N_11725,N_10515,N_10612);
nor U11726 (N_11726,N_10874,N_11233);
or U11727 (N_11727,N_10845,N_11108);
nand U11728 (N_11728,N_10670,N_10573);
and U11729 (N_11729,N_10783,N_10979);
nand U11730 (N_11730,N_10888,N_11165);
and U11731 (N_11731,N_10602,N_10757);
nand U11732 (N_11732,N_11165,N_10965);
and U11733 (N_11733,N_10647,N_10627);
or U11734 (N_11734,N_10607,N_11232);
or U11735 (N_11735,N_11119,N_11018);
nand U11736 (N_11736,N_10881,N_10601);
nand U11737 (N_11737,N_11112,N_10579);
or U11738 (N_11738,N_10634,N_11080);
or U11739 (N_11739,N_10919,N_10897);
or U11740 (N_11740,N_11069,N_10752);
nor U11741 (N_11741,N_11005,N_10978);
or U11742 (N_11742,N_10916,N_11168);
nand U11743 (N_11743,N_10672,N_10972);
or U11744 (N_11744,N_10735,N_10519);
xnor U11745 (N_11745,N_11055,N_10982);
and U11746 (N_11746,N_10555,N_10565);
or U11747 (N_11747,N_10847,N_11163);
or U11748 (N_11748,N_10677,N_10917);
nor U11749 (N_11749,N_11194,N_10793);
nor U11750 (N_11750,N_10527,N_10967);
nor U11751 (N_11751,N_11100,N_10635);
nand U11752 (N_11752,N_10912,N_11081);
nand U11753 (N_11753,N_10700,N_11168);
and U11754 (N_11754,N_11205,N_11074);
nor U11755 (N_11755,N_10773,N_10761);
and U11756 (N_11756,N_10837,N_11087);
nand U11757 (N_11757,N_10746,N_11181);
or U11758 (N_11758,N_10840,N_10714);
or U11759 (N_11759,N_10745,N_10527);
xor U11760 (N_11760,N_10760,N_11066);
nor U11761 (N_11761,N_10865,N_10740);
nor U11762 (N_11762,N_10936,N_11152);
nor U11763 (N_11763,N_11105,N_11239);
and U11764 (N_11764,N_11086,N_10899);
nand U11765 (N_11765,N_11223,N_10928);
xnor U11766 (N_11766,N_10623,N_10518);
or U11767 (N_11767,N_10601,N_11225);
nor U11768 (N_11768,N_10633,N_10990);
or U11769 (N_11769,N_10805,N_11133);
or U11770 (N_11770,N_10733,N_10657);
nand U11771 (N_11771,N_10879,N_10520);
or U11772 (N_11772,N_10817,N_10725);
xnor U11773 (N_11773,N_10687,N_10892);
nor U11774 (N_11774,N_11037,N_10973);
nand U11775 (N_11775,N_10613,N_10839);
and U11776 (N_11776,N_10675,N_10915);
nand U11777 (N_11777,N_10664,N_11089);
or U11778 (N_11778,N_10894,N_11019);
nand U11779 (N_11779,N_11117,N_10890);
nor U11780 (N_11780,N_10977,N_10644);
nor U11781 (N_11781,N_11158,N_10575);
nor U11782 (N_11782,N_10850,N_10611);
nor U11783 (N_11783,N_10837,N_10589);
and U11784 (N_11784,N_10983,N_10819);
and U11785 (N_11785,N_10599,N_10808);
or U11786 (N_11786,N_10981,N_10871);
nor U11787 (N_11787,N_10796,N_11176);
or U11788 (N_11788,N_10831,N_10734);
nand U11789 (N_11789,N_11037,N_10504);
nand U11790 (N_11790,N_11088,N_10562);
and U11791 (N_11791,N_10967,N_10949);
nor U11792 (N_11792,N_11120,N_10514);
nor U11793 (N_11793,N_11043,N_10654);
nand U11794 (N_11794,N_10724,N_11175);
nor U11795 (N_11795,N_10626,N_10936);
or U11796 (N_11796,N_11092,N_10889);
xor U11797 (N_11797,N_10668,N_11248);
and U11798 (N_11798,N_10887,N_11095);
nand U11799 (N_11799,N_10833,N_11004);
and U11800 (N_11800,N_11152,N_11064);
nand U11801 (N_11801,N_10824,N_10999);
and U11802 (N_11802,N_10605,N_10805);
nand U11803 (N_11803,N_10563,N_11172);
nand U11804 (N_11804,N_11071,N_11167);
nand U11805 (N_11805,N_10699,N_10857);
and U11806 (N_11806,N_10574,N_10696);
or U11807 (N_11807,N_10869,N_11080);
or U11808 (N_11808,N_10742,N_10515);
nand U11809 (N_11809,N_10667,N_10924);
nand U11810 (N_11810,N_11003,N_10843);
nand U11811 (N_11811,N_11086,N_11194);
or U11812 (N_11812,N_11139,N_10758);
nand U11813 (N_11813,N_10917,N_10688);
nand U11814 (N_11814,N_11085,N_10563);
or U11815 (N_11815,N_11071,N_11129);
or U11816 (N_11816,N_10709,N_10906);
nor U11817 (N_11817,N_10790,N_10629);
nor U11818 (N_11818,N_10910,N_10973);
nand U11819 (N_11819,N_11178,N_10503);
or U11820 (N_11820,N_10674,N_10646);
nor U11821 (N_11821,N_11235,N_11188);
or U11822 (N_11822,N_10513,N_10705);
and U11823 (N_11823,N_11161,N_11107);
nor U11824 (N_11824,N_11215,N_11194);
and U11825 (N_11825,N_10723,N_11169);
and U11826 (N_11826,N_10824,N_10605);
nor U11827 (N_11827,N_10638,N_10839);
xor U11828 (N_11828,N_10529,N_11011);
or U11829 (N_11829,N_11220,N_11199);
nand U11830 (N_11830,N_11089,N_10602);
nor U11831 (N_11831,N_10874,N_10500);
or U11832 (N_11832,N_11122,N_10524);
or U11833 (N_11833,N_10914,N_11140);
or U11834 (N_11834,N_10648,N_11137);
nand U11835 (N_11835,N_11048,N_11106);
xor U11836 (N_11836,N_11206,N_10915);
nor U11837 (N_11837,N_10680,N_10509);
or U11838 (N_11838,N_10877,N_11230);
nand U11839 (N_11839,N_10668,N_10631);
nor U11840 (N_11840,N_10883,N_10569);
or U11841 (N_11841,N_10763,N_10891);
and U11842 (N_11842,N_10699,N_10548);
or U11843 (N_11843,N_11238,N_10808);
and U11844 (N_11844,N_10937,N_11193);
and U11845 (N_11845,N_11036,N_11116);
or U11846 (N_11846,N_10830,N_11154);
or U11847 (N_11847,N_10873,N_10827);
or U11848 (N_11848,N_10972,N_11062);
nor U11849 (N_11849,N_10595,N_10794);
and U11850 (N_11850,N_10872,N_10744);
and U11851 (N_11851,N_11111,N_11218);
and U11852 (N_11852,N_10795,N_10661);
and U11853 (N_11853,N_11036,N_10704);
nand U11854 (N_11854,N_10901,N_10726);
or U11855 (N_11855,N_10995,N_10900);
nand U11856 (N_11856,N_11193,N_10685);
or U11857 (N_11857,N_11046,N_10553);
nand U11858 (N_11858,N_10857,N_11248);
or U11859 (N_11859,N_11033,N_10974);
nor U11860 (N_11860,N_11164,N_11138);
or U11861 (N_11861,N_11032,N_11209);
or U11862 (N_11862,N_11159,N_10974);
and U11863 (N_11863,N_11007,N_10928);
and U11864 (N_11864,N_11125,N_10951);
or U11865 (N_11865,N_10981,N_10582);
or U11866 (N_11866,N_10769,N_11156);
and U11867 (N_11867,N_10724,N_10805);
or U11868 (N_11868,N_11141,N_10972);
nor U11869 (N_11869,N_11166,N_10593);
or U11870 (N_11870,N_10822,N_10985);
or U11871 (N_11871,N_10537,N_11196);
nor U11872 (N_11872,N_10512,N_10761);
and U11873 (N_11873,N_10592,N_10944);
or U11874 (N_11874,N_10543,N_10686);
nand U11875 (N_11875,N_10508,N_11214);
nor U11876 (N_11876,N_10756,N_10621);
or U11877 (N_11877,N_10831,N_11199);
nor U11878 (N_11878,N_10850,N_11223);
and U11879 (N_11879,N_10710,N_10895);
and U11880 (N_11880,N_10974,N_10889);
nor U11881 (N_11881,N_11195,N_10828);
nand U11882 (N_11882,N_11094,N_11030);
and U11883 (N_11883,N_10961,N_11058);
and U11884 (N_11884,N_10937,N_11093);
nand U11885 (N_11885,N_11099,N_11040);
or U11886 (N_11886,N_10769,N_11071);
and U11887 (N_11887,N_10551,N_10636);
xnor U11888 (N_11888,N_11155,N_11214);
or U11889 (N_11889,N_10707,N_10689);
nor U11890 (N_11890,N_11123,N_10558);
nor U11891 (N_11891,N_11130,N_10947);
and U11892 (N_11892,N_10551,N_11112);
xor U11893 (N_11893,N_11031,N_10813);
nor U11894 (N_11894,N_10592,N_10904);
and U11895 (N_11895,N_11156,N_10563);
and U11896 (N_11896,N_10993,N_11065);
nand U11897 (N_11897,N_10928,N_10546);
nand U11898 (N_11898,N_11248,N_11245);
xnor U11899 (N_11899,N_11234,N_11054);
nor U11900 (N_11900,N_11058,N_10661);
or U11901 (N_11901,N_10860,N_11215);
and U11902 (N_11902,N_10665,N_10872);
nor U11903 (N_11903,N_10790,N_10550);
or U11904 (N_11904,N_11175,N_11217);
nor U11905 (N_11905,N_10754,N_11161);
nor U11906 (N_11906,N_10945,N_11088);
nor U11907 (N_11907,N_10915,N_10988);
and U11908 (N_11908,N_10741,N_10562);
or U11909 (N_11909,N_10536,N_10857);
or U11910 (N_11910,N_11166,N_10778);
or U11911 (N_11911,N_11087,N_10928);
xnor U11912 (N_11912,N_10657,N_11239);
and U11913 (N_11913,N_10995,N_10988);
nor U11914 (N_11914,N_10516,N_10659);
nand U11915 (N_11915,N_10711,N_11130);
nand U11916 (N_11916,N_11059,N_10897);
or U11917 (N_11917,N_10774,N_10585);
nor U11918 (N_11918,N_10898,N_10577);
and U11919 (N_11919,N_10767,N_10586);
nand U11920 (N_11920,N_10812,N_11042);
xor U11921 (N_11921,N_11191,N_10702);
or U11922 (N_11922,N_10786,N_11067);
and U11923 (N_11923,N_10631,N_10534);
and U11924 (N_11924,N_10762,N_10641);
and U11925 (N_11925,N_10530,N_10684);
nor U11926 (N_11926,N_10983,N_11180);
nand U11927 (N_11927,N_10935,N_10637);
or U11928 (N_11928,N_10777,N_10536);
or U11929 (N_11929,N_11046,N_10949);
nand U11930 (N_11930,N_11208,N_11049);
nor U11931 (N_11931,N_11109,N_10802);
nor U11932 (N_11932,N_11031,N_10642);
or U11933 (N_11933,N_10953,N_10562);
nor U11934 (N_11934,N_11089,N_11122);
nor U11935 (N_11935,N_10685,N_11248);
xnor U11936 (N_11936,N_10610,N_10841);
nor U11937 (N_11937,N_10689,N_10768);
nand U11938 (N_11938,N_10654,N_10512);
xor U11939 (N_11939,N_11011,N_10569);
and U11940 (N_11940,N_10959,N_10749);
nor U11941 (N_11941,N_11079,N_10631);
or U11942 (N_11942,N_10743,N_10854);
nand U11943 (N_11943,N_10622,N_11228);
nand U11944 (N_11944,N_10693,N_10552);
and U11945 (N_11945,N_11247,N_10989);
and U11946 (N_11946,N_10769,N_10963);
and U11947 (N_11947,N_10823,N_10502);
and U11948 (N_11948,N_10883,N_11033);
nor U11949 (N_11949,N_10800,N_11167);
xor U11950 (N_11950,N_10730,N_10968);
nor U11951 (N_11951,N_10514,N_11188);
nor U11952 (N_11952,N_10961,N_11078);
or U11953 (N_11953,N_10987,N_10908);
xor U11954 (N_11954,N_11155,N_10666);
or U11955 (N_11955,N_10689,N_10981);
xnor U11956 (N_11956,N_10666,N_10563);
xnor U11957 (N_11957,N_10745,N_11090);
nand U11958 (N_11958,N_11068,N_11091);
and U11959 (N_11959,N_10757,N_10904);
and U11960 (N_11960,N_10729,N_11008);
nor U11961 (N_11961,N_11035,N_10500);
nor U11962 (N_11962,N_10675,N_10800);
and U11963 (N_11963,N_10638,N_10714);
and U11964 (N_11964,N_10842,N_10821);
or U11965 (N_11965,N_10738,N_10937);
and U11966 (N_11966,N_10715,N_10806);
xor U11967 (N_11967,N_10740,N_11008);
and U11968 (N_11968,N_11228,N_10943);
nand U11969 (N_11969,N_10997,N_11082);
or U11970 (N_11970,N_11144,N_10623);
nor U11971 (N_11971,N_10811,N_10553);
nand U11972 (N_11972,N_10651,N_10818);
and U11973 (N_11973,N_11243,N_10942);
nand U11974 (N_11974,N_10966,N_10869);
nor U11975 (N_11975,N_11037,N_11060);
or U11976 (N_11976,N_10844,N_11129);
xnor U11977 (N_11977,N_10831,N_10584);
or U11978 (N_11978,N_11082,N_10783);
or U11979 (N_11979,N_10513,N_10731);
xor U11980 (N_11980,N_10678,N_11056);
and U11981 (N_11981,N_10783,N_10898);
xnor U11982 (N_11982,N_11239,N_10605);
and U11983 (N_11983,N_10701,N_10575);
xnor U11984 (N_11984,N_10753,N_10604);
or U11985 (N_11985,N_10917,N_10673);
nand U11986 (N_11986,N_10786,N_10715);
or U11987 (N_11987,N_10999,N_10737);
and U11988 (N_11988,N_11062,N_10728);
nand U11989 (N_11989,N_11206,N_11093);
nor U11990 (N_11990,N_10692,N_11220);
xnor U11991 (N_11991,N_11165,N_10518);
and U11992 (N_11992,N_11232,N_11117);
nor U11993 (N_11993,N_10652,N_10813);
xor U11994 (N_11994,N_10841,N_10803);
or U11995 (N_11995,N_10641,N_11225);
xor U11996 (N_11996,N_10879,N_10546);
nand U11997 (N_11997,N_10871,N_11093);
nor U11998 (N_11998,N_10939,N_10568);
nand U11999 (N_11999,N_11192,N_11004);
nand U12000 (N_12000,N_11734,N_11949);
nand U12001 (N_12001,N_11480,N_11772);
and U12002 (N_12002,N_11961,N_11631);
nand U12003 (N_12003,N_11604,N_11917);
nand U12004 (N_12004,N_11743,N_11569);
nor U12005 (N_12005,N_11648,N_11972);
nand U12006 (N_12006,N_11284,N_11442);
and U12007 (N_12007,N_11377,N_11849);
nand U12008 (N_12008,N_11291,N_11730);
nand U12009 (N_12009,N_11558,N_11798);
nor U12010 (N_12010,N_11292,N_11955);
nor U12011 (N_12011,N_11775,N_11898);
nand U12012 (N_12012,N_11826,N_11708);
nor U12013 (N_12013,N_11928,N_11492);
or U12014 (N_12014,N_11266,N_11953);
and U12015 (N_12015,N_11706,N_11767);
and U12016 (N_12016,N_11739,N_11540);
xnor U12017 (N_12017,N_11787,N_11516);
nor U12018 (N_12018,N_11904,N_11658);
nor U12019 (N_12019,N_11453,N_11645);
nor U12020 (N_12020,N_11446,N_11286);
nor U12021 (N_12021,N_11966,N_11725);
or U12022 (N_12022,N_11590,N_11400);
nand U12023 (N_12023,N_11287,N_11721);
or U12024 (N_12024,N_11547,N_11525);
nor U12025 (N_12025,N_11383,N_11894);
and U12026 (N_12026,N_11555,N_11983);
nor U12027 (N_12027,N_11689,N_11663);
or U12028 (N_12028,N_11533,N_11654);
and U12029 (N_12029,N_11923,N_11507);
and U12030 (N_12030,N_11448,N_11926);
or U12031 (N_12031,N_11384,N_11500);
xor U12032 (N_12032,N_11445,N_11799);
nand U12033 (N_12033,N_11583,N_11840);
and U12034 (N_12034,N_11574,N_11831);
xor U12035 (N_12035,N_11549,N_11333);
nor U12036 (N_12036,N_11657,N_11993);
xor U12037 (N_12037,N_11581,N_11834);
nand U12038 (N_12038,N_11825,N_11944);
and U12039 (N_12039,N_11603,N_11539);
and U12040 (N_12040,N_11815,N_11587);
nor U12041 (N_12041,N_11874,N_11495);
or U12042 (N_12042,N_11762,N_11548);
and U12043 (N_12043,N_11577,N_11885);
and U12044 (N_12044,N_11807,N_11842);
and U12045 (N_12045,N_11477,N_11372);
and U12046 (N_12046,N_11634,N_11561);
nor U12047 (N_12047,N_11393,N_11309);
and U12048 (N_12048,N_11370,N_11951);
nand U12049 (N_12049,N_11550,N_11310);
nand U12050 (N_12050,N_11502,N_11353);
or U12051 (N_12051,N_11943,N_11594);
nand U12052 (N_12052,N_11674,N_11413);
or U12053 (N_12053,N_11638,N_11864);
xor U12054 (N_12054,N_11470,N_11295);
nand U12055 (N_12055,N_11314,N_11343);
nor U12056 (N_12056,N_11978,N_11395);
nand U12057 (N_12057,N_11858,N_11436);
or U12058 (N_12058,N_11366,N_11302);
nor U12059 (N_12059,N_11910,N_11509);
nor U12060 (N_12060,N_11911,N_11935);
and U12061 (N_12061,N_11726,N_11999);
nand U12062 (N_12062,N_11850,N_11356);
nand U12063 (N_12063,N_11802,N_11852);
nor U12064 (N_12064,N_11979,N_11407);
or U12065 (N_12065,N_11890,N_11636);
xnor U12066 (N_12066,N_11256,N_11683);
nor U12067 (N_12067,N_11897,N_11680);
nor U12068 (N_12068,N_11731,N_11348);
or U12069 (N_12069,N_11293,N_11517);
nor U12070 (N_12070,N_11260,N_11913);
or U12071 (N_12071,N_11289,N_11559);
nand U12072 (N_12072,N_11253,N_11780);
or U12073 (N_12073,N_11317,N_11661);
nor U12074 (N_12074,N_11791,N_11626);
and U12075 (N_12075,N_11740,N_11675);
or U12076 (N_12076,N_11524,N_11833);
nand U12077 (N_12077,N_11820,N_11251);
nand U12078 (N_12078,N_11347,N_11932);
nand U12079 (N_12079,N_11929,N_11279);
or U12080 (N_12080,N_11272,N_11766);
xnor U12081 (N_12081,N_11434,N_11705);
or U12082 (N_12082,N_11596,N_11744);
nor U12083 (N_12083,N_11489,N_11963);
xor U12084 (N_12084,N_11992,N_11461);
nor U12085 (N_12085,N_11429,N_11591);
or U12086 (N_12086,N_11968,N_11883);
or U12087 (N_12087,N_11622,N_11670);
or U12088 (N_12088,N_11467,N_11867);
nor U12089 (N_12089,N_11621,N_11403);
nor U12090 (N_12090,N_11554,N_11985);
or U12091 (N_12091,N_11936,N_11582);
nor U12092 (N_12092,N_11350,N_11805);
nand U12093 (N_12093,N_11769,N_11456);
and U12094 (N_12094,N_11496,N_11484);
xnor U12095 (N_12095,N_11494,N_11564);
or U12096 (N_12096,N_11651,N_11427);
nor U12097 (N_12097,N_11504,N_11482);
nand U12098 (N_12098,N_11886,N_11503);
nor U12099 (N_12099,N_11270,N_11940);
nand U12100 (N_12100,N_11315,N_11649);
and U12101 (N_12101,N_11971,N_11324);
or U12102 (N_12102,N_11981,N_11598);
nand U12103 (N_12103,N_11462,N_11385);
nor U12104 (N_12104,N_11946,N_11746);
nor U12105 (N_12105,N_11602,N_11501);
or U12106 (N_12106,N_11712,N_11685);
nor U12107 (N_12107,N_11511,N_11280);
nor U12108 (N_12108,N_11514,N_11557);
nand U12109 (N_12109,N_11584,N_11902);
xor U12110 (N_12110,N_11303,N_11551);
or U12111 (N_12111,N_11488,N_11877);
or U12112 (N_12112,N_11457,N_11363);
nand U12113 (N_12113,N_11401,N_11392);
nor U12114 (N_12114,N_11778,N_11782);
nand U12115 (N_12115,N_11531,N_11522);
nand U12116 (N_12116,N_11320,N_11471);
nand U12117 (N_12117,N_11640,N_11790);
nand U12118 (N_12118,N_11696,N_11747);
xnor U12119 (N_12119,N_11515,N_11274);
and U12120 (N_12120,N_11956,N_11793);
nor U12121 (N_12121,N_11571,N_11465);
nand U12122 (N_12122,N_11854,N_11642);
and U12123 (N_12123,N_11472,N_11837);
and U12124 (N_12124,N_11757,N_11847);
and U12125 (N_12125,N_11727,N_11311);
nor U12126 (N_12126,N_11633,N_11318);
and U12127 (N_12127,N_11433,N_11895);
nor U12128 (N_12128,N_11773,N_11869);
or U12129 (N_12129,N_11610,N_11258);
xnor U12130 (N_12130,N_11358,N_11312);
or U12131 (N_12131,N_11447,N_11960);
or U12132 (N_12132,N_11728,N_11655);
nand U12133 (N_12133,N_11475,N_11637);
nand U12134 (N_12134,N_11485,N_11327);
and U12135 (N_12135,N_11693,N_11466);
or U12136 (N_12136,N_11975,N_11454);
and U12137 (N_12137,N_11277,N_11824);
nand U12138 (N_12138,N_11268,N_11296);
xor U12139 (N_12139,N_11276,N_11952);
and U12140 (N_12140,N_11964,N_11271);
nand U12141 (N_12141,N_11828,N_11694);
nand U12142 (N_12142,N_11255,N_11907);
or U12143 (N_12143,N_11529,N_11418);
or U12144 (N_12144,N_11829,N_11662);
and U12145 (N_12145,N_11821,N_11337);
or U12146 (N_12146,N_11543,N_11659);
and U12147 (N_12147,N_11660,N_11424);
nor U12148 (N_12148,N_11570,N_11681);
and U12149 (N_12149,N_11534,N_11360);
nand U12150 (N_12150,N_11437,N_11893);
nand U12151 (N_12151,N_11779,N_11459);
xnor U12152 (N_12152,N_11801,N_11553);
or U12153 (N_12153,N_11924,N_11394);
nor U12154 (N_12154,N_11860,N_11933);
nand U12155 (N_12155,N_11408,N_11344);
nor U12156 (N_12156,N_11367,N_11761);
or U12157 (N_12157,N_11439,N_11668);
nor U12158 (N_12158,N_11856,N_11733);
or U12159 (N_12159,N_11735,N_11717);
xnor U12160 (N_12160,N_11378,N_11892);
nor U12161 (N_12161,N_11716,N_11566);
or U12162 (N_12162,N_11901,N_11490);
and U12163 (N_12163,N_11617,N_11464);
nor U12164 (N_12164,N_11977,N_11411);
and U12165 (N_12165,N_11425,N_11947);
or U12166 (N_12166,N_11781,N_11868);
and U12167 (N_12167,N_11756,N_11764);
or U12168 (N_12168,N_11493,N_11299);
and U12169 (N_12169,N_11386,N_11530);
or U12170 (N_12170,N_11812,N_11723);
or U12171 (N_12171,N_11593,N_11941);
or U12172 (N_12172,N_11599,N_11380);
nand U12173 (N_12173,N_11455,N_11714);
and U12174 (N_12174,N_11752,N_11934);
nand U12175 (N_12175,N_11352,N_11770);
or U12176 (N_12176,N_11745,N_11510);
or U12177 (N_12177,N_11600,N_11758);
xnor U12178 (N_12178,N_11405,N_11342);
and U12179 (N_12179,N_11967,N_11345);
xnor U12180 (N_12180,N_11871,N_11519);
nand U12181 (N_12181,N_11688,N_11612);
nand U12182 (N_12182,N_11406,N_11989);
or U12183 (N_12183,N_11635,N_11435);
or U12184 (N_12184,N_11639,N_11281);
or U12185 (N_12185,N_11261,N_11959);
nor U12186 (N_12186,N_11387,N_11891);
and U12187 (N_12187,N_11597,N_11527);
nand U12188 (N_12188,N_11646,N_11699);
nor U12189 (N_12189,N_11653,N_11449);
and U12190 (N_12190,N_11544,N_11374);
nand U12191 (N_12191,N_11879,N_11682);
or U12192 (N_12192,N_11800,N_11285);
nand U12193 (N_12193,N_11803,N_11322);
nand U12194 (N_12194,N_11351,N_11873);
or U12195 (N_12195,N_11664,N_11468);
nand U12196 (N_12196,N_11925,N_11718);
and U12197 (N_12197,N_11278,N_11986);
and U12198 (N_12198,N_11753,N_11880);
xnor U12199 (N_12199,N_11722,N_11938);
xnor U12200 (N_12200,N_11580,N_11866);
xnor U12201 (N_12201,N_11578,N_11263);
and U12202 (N_12202,N_11630,N_11573);
and U12203 (N_12203,N_11912,N_11476);
xor U12204 (N_12204,N_11373,N_11592);
or U12205 (N_12205,N_11538,N_11520);
nand U12206 (N_12206,N_11795,N_11273);
nor U12207 (N_12207,N_11836,N_11995);
nand U12208 (N_12208,N_11861,N_11336);
and U12209 (N_12209,N_11368,N_11789);
or U12210 (N_12210,N_11361,N_11818);
xnor U12211 (N_12211,N_11676,N_11264);
nand U12212 (N_12212,N_11528,N_11665);
nor U12213 (N_12213,N_11294,N_11497);
and U12214 (N_12214,N_11498,N_11632);
nor U12215 (N_12215,N_11624,N_11369);
nand U12216 (N_12216,N_11809,N_11410);
xor U12217 (N_12217,N_11896,N_11915);
or U12218 (N_12218,N_11765,N_11341);
nand U12219 (N_12219,N_11875,N_11774);
and U12220 (N_12220,N_11629,N_11754);
nor U12221 (N_12221,N_11398,N_11474);
nor U12222 (N_12222,N_11419,N_11338);
and U12223 (N_12223,N_11729,N_11922);
and U12224 (N_12224,N_11323,N_11613);
nand U12225 (N_12225,N_11397,N_11703);
nor U12226 (N_12226,N_11463,N_11997);
or U12227 (N_12227,N_11257,N_11505);
or U12228 (N_12228,N_11313,N_11865);
nand U12229 (N_12229,N_11620,N_11939);
xor U12230 (N_12230,N_11556,N_11267);
or U12231 (N_12231,N_11623,N_11863);
and U12232 (N_12232,N_11487,N_11331);
nor U12233 (N_12233,N_11346,N_11432);
xnor U12234 (N_12234,N_11908,N_11919);
and U12235 (N_12235,N_11671,N_11980);
and U12236 (N_12236,N_11563,N_11823);
nor U12237 (N_12237,N_11948,N_11857);
nand U12238 (N_12238,N_11878,N_11950);
xor U12239 (N_12239,N_11822,N_11269);
nand U12240 (N_12240,N_11567,N_11720);
and U12241 (N_12241,N_11585,N_11452);
xnor U12242 (N_12242,N_11469,N_11399);
and U12243 (N_12243,N_11641,N_11698);
nand U12244 (N_12244,N_11513,N_11381);
nand U12245 (N_12245,N_11644,N_11316);
nand U12246 (N_12246,N_11576,N_11535);
nor U12247 (N_12247,N_11304,N_11987);
xnor U12248 (N_12248,N_11816,N_11458);
or U12249 (N_12249,N_11899,N_11389);
nor U12250 (N_12250,N_11307,N_11954);
nand U12251 (N_12251,N_11562,N_11297);
and U12252 (N_12252,N_11859,N_11990);
nor U12253 (N_12253,N_11627,N_11450);
and U12254 (N_12254,N_11426,N_11738);
nor U12255 (N_12255,N_11423,N_11906);
or U12256 (N_12256,N_11306,N_11262);
or U12257 (N_12257,N_11308,N_11619);
nand U12258 (N_12258,N_11927,N_11460);
nand U12259 (N_12259,N_11958,N_11918);
and U12260 (N_12260,N_11330,N_11788);
and U12261 (N_12261,N_11499,N_11444);
nor U12262 (N_12262,N_11512,N_11546);
or U12263 (N_12263,N_11695,N_11250);
or U12264 (N_12264,N_11914,N_11305);
or U12265 (N_12265,N_11532,N_11937);
nand U12266 (N_12266,N_11719,N_11813);
or U12267 (N_12267,N_11855,N_11900);
nand U12268 (N_12268,N_11541,N_11428);
and U12269 (N_12269,N_11830,N_11608);
and U12270 (N_12270,N_11707,N_11486);
nand U12271 (N_12271,N_11969,N_11376);
and U12272 (N_12272,N_11652,N_11526);
or U12273 (N_12273,N_11355,N_11785);
nand U12274 (N_12274,N_11827,N_11996);
or U12275 (N_12275,N_11382,N_11814);
xor U12276 (N_12276,N_11364,N_11690);
and U12277 (N_12277,N_11905,N_11290);
and U12278 (N_12278,N_11396,N_11390);
and U12279 (N_12279,N_11677,N_11838);
nor U12280 (N_12280,N_11970,N_11848);
nor U12281 (N_12281,N_11794,N_11841);
and U12282 (N_12282,N_11884,N_11328);
and U12283 (N_12283,N_11870,N_11702);
and U12284 (N_12284,N_11988,N_11379);
nand U12285 (N_12285,N_11441,N_11768);
and U12286 (N_12286,N_11365,N_11810);
nor U12287 (N_12287,N_11615,N_11736);
or U12288 (N_12288,N_11991,N_11611);
xnor U12289 (N_12289,N_11252,N_11711);
xnor U12290 (N_12290,N_11962,N_11672);
or U12291 (N_12291,N_11973,N_11760);
nand U12292 (N_12292,N_11930,N_11876);
xor U12293 (N_12293,N_11568,N_11942);
or U12294 (N_12294,N_11982,N_11412);
or U12295 (N_12295,N_11404,N_11518);
and U12296 (N_12296,N_11804,N_11371);
or U12297 (N_12297,N_11420,N_11416);
nor U12298 (N_12298,N_11832,N_11375);
nor U12299 (N_12299,N_11438,N_11771);
nand U12300 (N_12300,N_11391,N_11616);
xnor U12301 (N_12301,N_11715,N_11422);
or U12302 (N_12302,N_11325,N_11796);
and U12303 (N_12303,N_11440,N_11692);
nor U12304 (N_12304,N_11319,N_11483);
and U12305 (N_12305,N_11750,N_11254);
nor U12306 (N_12306,N_11606,N_11650);
nand U12307 (N_12307,N_11552,N_11326);
or U12308 (N_12308,N_11508,N_11839);
nand U12309 (N_12309,N_11409,N_11421);
nand U12310 (N_12310,N_11321,N_11339);
and U12311 (N_12311,N_11759,N_11607);
or U12312 (N_12312,N_11872,N_11340);
xnor U12313 (N_12313,N_11710,N_11984);
xnor U12314 (N_12314,N_11301,N_11862);
xnor U12315 (N_12315,N_11362,N_11579);
and U12316 (N_12316,N_11354,N_11853);
nor U12317 (N_12317,N_11565,N_11601);
or U12318 (N_12318,N_11595,N_11335);
nand U12319 (N_12319,N_11537,N_11784);
nand U12320 (N_12320,N_11491,N_11835);
or U12321 (N_12321,N_11275,N_11618);
nor U12322 (N_12322,N_11845,N_11687);
and U12323 (N_12323,N_11588,N_11334);
nor U12324 (N_12324,N_11763,N_11732);
or U12325 (N_12325,N_11819,N_11776);
and U12326 (N_12326,N_11300,N_11713);
nor U12327 (N_12327,N_11415,N_11283);
nand U12328 (N_12328,N_11625,N_11402);
nor U12329 (N_12329,N_11589,N_11332);
nand U12330 (N_12330,N_11755,N_11282);
or U12331 (N_12331,N_11605,N_11786);
nor U12332 (N_12332,N_11749,N_11451);
nand U12333 (N_12333,N_11536,N_11572);
or U12334 (N_12334,N_11976,N_11542);
nand U12335 (N_12335,N_11560,N_11851);
nand U12336 (N_12336,N_11417,N_11521);
or U12337 (N_12337,N_11298,N_11479);
nand U12338 (N_12338,N_11817,N_11945);
or U12339 (N_12339,N_11478,N_11349);
nand U12340 (N_12340,N_11704,N_11888);
or U12341 (N_12341,N_11742,N_11414);
or U12342 (N_12342,N_11473,N_11903);
and U12343 (N_12343,N_11709,N_11669);
or U12344 (N_12344,N_11443,N_11887);
or U12345 (N_12345,N_11679,N_11697);
or U12346 (N_12346,N_11724,N_11647);
xnor U12347 (N_12347,N_11931,N_11751);
nand U12348 (N_12348,N_11609,N_11921);
xnor U12349 (N_12349,N_11737,N_11889);
nor U12350 (N_12350,N_11974,N_11701);
nand U12351 (N_12351,N_11666,N_11792);
and U12352 (N_12352,N_11686,N_11748);
xnor U12353 (N_12353,N_11843,N_11643);
nor U12354 (N_12354,N_11359,N_11684);
nor U12355 (N_12355,N_11265,N_11673);
nand U12356 (N_12356,N_11741,N_11909);
nor U12357 (N_12357,N_11523,N_11882);
nor U12358 (N_12358,N_11783,N_11808);
nand U12359 (N_12359,N_11431,N_11678);
or U12360 (N_12360,N_11811,N_11656);
or U12361 (N_12361,N_11700,N_11994);
and U12362 (N_12362,N_11998,N_11575);
nor U12363 (N_12363,N_11481,N_11965);
nor U12364 (N_12364,N_11545,N_11586);
nor U12365 (N_12365,N_11329,N_11777);
nand U12366 (N_12366,N_11506,N_11357);
nand U12367 (N_12367,N_11881,N_11806);
nand U12368 (N_12368,N_11259,N_11846);
nor U12369 (N_12369,N_11957,N_11916);
or U12370 (N_12370,N_11614,N_11388);
and U12371 (N_12371,N_11844,N_11628);
and U12372 (N_12372,N_11430,N_11691);
or U12373 (N_12373,N_11797,N_11288);
nor U12374 (N_12374,N_11920,N_11667);
or U12375 (N_12375,N_11906,N_11603);
xor U12376 (N_12376,N_11793,N_11405);
xor U12377 (N_12377,N_11575,N_11519);
nand U12378 (N_12378,N_11252,N_11584);
and U12379 (N_12379,N_11612,N_11757);
nand U12380 (N_12380,N_11995,N_11687);
nand U12381 (N_12381,N_11294,N_11832);
xor U12382 (N_12382,N_11444,N_11582);
and U12383 (N_12383,N_11559,N_11640);
xor U12384 (N_12384,N_11947,N_11872);
xor U12385 (N_12385,N_11946,N_11366);
nor U12386 (N_12386,N_11271,N_11807);
or U12387 (N_12387,N_11794,N_11720);
xor U12388 (N_12388,N_11380,N_11593);
and U12389 (N_12389,N_11951,N_11746);
nor U12390 (N_12390,N_11637,N_11293);
or U12391 (N_12391,N_11419,N_11992);
or U12392 (N_12392,N_11984,N_11573);
nand U12393 (N_12393,N_11658,N_11292);
nand U12394 (N_12394,N_11265,N_11824);
and U12395 (N_12395,N_11943,N_11551);
nand U12396 (N_12396,N_11497,N_11507);
and U12397 (N_12397,N_11833,N_11356);
nor U12398 (N_12398,N_11413,N_11570);
nand U12399 (N_12399,N_11992,N_11287);
nand U12400 (N_12400,N_11576,N_11253);
nor U12401 (N_12401,N_11486,N_11662);
or U12402 (N_12402,N_11259,N_11857);
nor U12403 (N_12403,N_11692,N_11607);
and U12404 (N_12404,N_11429,N_11687);
nand U12405 (N_12405,N_11416,N_11948);
xnor U12406 (N_12406,N_11617,N_11824);
nand U12407 (N_12407,N_11993,N_11359);
and U12408 (N_12408,N_11826,N_11452);
and U12409 (N_12409,N_11983,N_11891);
and U12410 (N_12410,N_11446,N_11961);
nor U12411 (N_12411,N_11909,N_11410);
or U12412 (N_12412,N_11995,N_11372);
and U12413 (N_12413,N_11304,N_11314);
nand U12414 (N_12414,N_11844,N_11796);
nor U12415 (N_12415,N_11984,N_11516);
nand U12416 (N_12416,N_11895,N_11404);
xor U12417 (N_12417,N_11780,N_11713);
and U12418 (N_12418,N_11495,N_11298);
or U12419 (N_12419,N_11268,N_11948);
nand U12420 (N_12420,N_11627,N_11299);
or U12421 (N_12421,N_11276,N_11270);
xor U12422 (N_12422,N_11381,N_11911);
or U12423 (N_12423,N_11550,N_11895);
or U12424 (N_12424,N_11676,N_11270);
and U12425 (N_12425,N_11785,N_11913);
nor U12426 (N_12426,N_11250,N_11743);
or U12427 (N_12427,N_11886,N_11749);
nand U12428 (N_12428,N_11633,N_11295);
or U12429 (N_12429,N_11962,N_11654);
nand U12430 (N_12430,N_11388,N_11440);
nor U12431 (N_12431,N_11956,N_11390);
nor U12432 (N_12432,N_11361,N_11301);
or U12433 (N_12433,N_11932,N_11634);
or U12434 (N_12434,N_11856,N_11329);
nand U12435 (N_12435,N_11310,N_11560);
xor U12436 (N_12436,N_11901,N_11924);
or U12437 (N_12437,N_11477,N_11277);
nand U12438 (N_12438,N_11620,N_11671);
xnor U12439 (N_12439,N_11896,N_11592);
or U12440 (N_12440,N_11876,N_11443);
or U12441 (N_12441,N_11651,N_11667);
xnor U12442 (N_12442,N_11854,N_11931);
or U12443 (N_12443,N_11651,N_11409);
nand U12444 (N_12444,N_11436,N_11653);
and U12445 (N_12445,N_11622,N_11790);
or U12446 (N_12446,N_11904,N_11621);
or U12447 (N_12447,N_11346,N_11749);
or U12448 (N_12448,N_11322,N_11648);
nor U12449 (N_12449,N_11944,N_11945);
nor U12450 (N_12450,N_11747,N_11892);
and U12451 (N_12451,N_11787,N_11938);
or U12452 (N_12452,N_11916,N_11816);
nand U12453 (N_12453,N_11805,N_11813);
and U12454 (N_12454,N_11291,N_11520);
or U12455 (N_12455,N_11439,N_11637);
or U12456 (N_12456,N_11252,N_11464);
nor U12457 (N_12457,N_11725,N_11638);
nand U12458 (N_12458,N_11694,N_11944);
nor U12459 (N_12459,N_11761,N_11513);
nor U12460 (N_12460,N_11333,N_11625);
nor U12461 (N_12461,N_11704,N_11804);
or U12462 (N_12462,N_11425,N_11821);
nand U12463 (N_12463,N_11599,N_11730);
and U12464 (N_12464,N_11986,N_11635);
and U12465 (N_12465,N_11305,N_11813);
xnor U12466 (N_12466,N_11909,N_11330);
or U12467 (N_12467,N_11344,N_11306);
xnor U12468 (N_12468,N_11286,N_11934);
or U12469 (N_12469,N_11272,N_11512);
nor U12470 (N_12470,N_11421,N_11877);
or U12471 (N_12471,N_11610,N_11593);
or U12472 (N_12472,N_11930,N_11481);
nand U12473 (N_12473,N_11274,N_11595);
xor U12474 (N_12474,N_11488,N_11432);
nand U12475 (N_12475,N_11868,N_11943);
or U12476 (N_12476,N_11826,N_11398);
nor U12477 (N_12477,N_11826,N_11298);
xor U12478 (N_12478,N_11615,N_11966);
nor U12479 (N_12479,N_11400,N_11465);
or U12480 (N_12480,N_11547,N_11763);
and U12481 (N_12481,N_11948,N_11347);
nand U12482 (N_12482,N_11758,N_11894);
nor U12483 (N_12483,N_11503,N_11333);
or U12484 (N_12484,N_11930,N_11437);
nand U12485 (N_12485,N_11926,N_11646);
nor U12486 (N_12486,N_11330,N_11997);
or U12487 (N_12487,N_11864,N_11355);
xor U12488 (N_12488,N_11883,N_11258);
and U12489 (N_12489,N_11747,N_11488);
nor U12490 (N_12490,N_11603,N_11979);
nand U12491 (N_12491,N_11453,N_11839);
xor U12492 (N_12492,N_11772,N_11389);
nand U12493 (N_12493,N_11317,N_11272);
nor U12494 (N_12494,N_11437,N_11441);
nor U12495 (N_12495,N_11960,N_11615);
or U12496 (N_12496,N_11597,N_11567);
or U12497 (N_12497,N_11962,N_11756);
nand U12498 (N_12498,N_11807,N_11475);
and U12499 (N_12499,N_11410,N_11670);
and U12500 (N_12500,N_11637,N_11849);
nor U12501 (N_12501,N_11695,N_11816);
or U12502 (N_12502,N_11649,N_11516);
nand U12503 (N_12503,N_11926,N_11485);
and U12504 (N_12504,N_11977,N_11764);
and U12505 (N_12505,N_11535,N_11684);
nand U12506 (N_12506,N_11311,N_11885);
and U12507 (N_12507,N_11341,N_11972);
or U12508 (N_12508,N_11317,N_11415);
and U12509 (N_12509,N_11911,N_11262);
nand U12510 (N_12510,N_11679,N_11916);
nor U12511 (N_12511,N_11793,N_11751);
xor U12512 (N_12512,N_11630,N_11295);
or U12513 (N_12513,N_11534,N_11845);
and U12514 (N_12514,N_11561,N_11609);
nor U12515 (N_12515,N_11320,N_11457);
nand U12516 (N_12516,N_11856,N_11370);
or U12517 (N_12517,N_11629,N_11916);
nand U12518 (N_12518,N_11687,N_11636);
or U12519 (N_12519,N_11274,N_11484);
or U12520 (N_12520,N_11694,N_11257);
and U12521 (N_12521,N_11587,N_11375);
xnor U12522 (N_12522,N_11398,N_11442);
or U12523 (N_12523,N_11865,N_11270);
or U12524 (N_12524,N_11797,N_11712);
or U12525 (N_12525,N_11462,N_11303);
nor U12526 (N_12526,N_11691,N_11776);
or U12527 (N_12527,N_11551,N_11965);
nor U12528 (N_12528,N_11403,N_11321);
xnor U12529 (N_12529,N_11961,N_11558);
nor U12530 (N_12530,N_11431,N_11260);
nor U12531 (N_12531,N_11432,N_11476);
or U12532 (N_12532,N_11918,N_11884);
nor U12533 (N_12533,N_11376,N_11888);
nor U12534 (N_12534,N_11584,N_11250);
nor U12535 (N_12535,N_11675,N_11844);
nor U12536 (N_12536,N_11671,N_11875);
nand U12537 (N_12537,N_11542,N_11682);
nand U12538 (N_12538,N_11999,N_11404);
or U12539 (N_12539,N_11514,N_11279);
or U12540 (N_12540,N_11486,N_11255);
nand U12541 (N_12541,N_11528,N_11794);
nand U12542 (N_12542,N_11643,N_11652);
nor U12543 (N_12543,N_11710,N_11813);
nor U12544 (N_12544,N_11350,N_11383);
xnor U12545 (N_12545,N_11263,N_11710);
nor U12546 (N_12546,N_11294,N_11582);
or U12547 (N_12547,N_11503,N_11475);
nand U12548 (N_12548,N_11643,N_11911);
and U12549 (N_12549,N_11865,N_11876);
and U12550 (N_12550,N_11361,N_11753);
nor U12551 (N_12551,N_11328,N_11867);
or U12552 (N_12552,N_11369,N_11692);
nand U12553 (N_12553,N_11402,N_11755);
and U12554 (N_12554,N_11459,N_11765);
nand U12555 (N_12555,N_11717,N_11826);
nand U12556 (N_12556,N_11548,N_11552);
or U12557 (N_12557,N_11378,N_11261);
nor U12558 (N_12558,N_11573,N_11597);
or U12559 (N_12559,N_11525,N_11587);
nand U12560 (N_12560,N_11776,N_11354);
or U12561 (N_12561,N_11290,N_11260);
nor U12562 (N_12562,N_11483,N_11750);
nor U12563 (N_12563,N_11838,N_11990);
and U12564 (N_12564,N_11459,N_11922);
and U12565 (N_12565,N_11930,N_11848);
or U12566 (N_12566,N_11313,N_11430);
or U12567 (N_12567,N_11789,N_11703);
or U12568 (N_12568,N_11950,N_11470);
nand U12569 (N_12569,N_11253,N_11799);
nand U12570 (N_12570,N_11488,N_11558);
nor U12571 (N_12571,N_11618,N_11496);
nor U12572 (N_12572,N_11516,N_11264);
nor U12573 (N_12573,N_11578,N_11347);
or U12574 (N_12574,N_11417,N_11704);
nand U12575 (N_12575,N_11969,N_11617);
nand U12576 (N_12576,N_11775,N_11375);
nand U12577 (N_12577,N_11723,N_11424);
nand U12578 (N_12578,N_11263,N_11290);
nor U12579 (N_12579,N_11956,N_11965);
nand U12580 (N_12580,N_11438,N_11927);
nor U12581 (N_12581,N_11587,N_11683);
or U12582 (N_12582,N_11910,N_11600);
nor U12583 (N_12583,N_11633,N_11876);
and U12584 (N_12584,N_11726,N_11286);
nor U12585 (N_12585,N_11614,N_11906);
or U12586 (N_12586,N_11286,N_11527);
nand U12587 (N_12587,N_11436,N_11688);
nand U12588 (N_12588,N_11274,N_11492);
or U12589 (N_12589,N_11285,N_11936);
nor U12590 (N_12590,N_11295,N_11744);
nor U12591 (N_12591,N_11817,N_11843);
xnor U12592 (N_12592,N_11370,N_11350);
nand U12593 (N_12593,N_11854,N_11699);
nor U12594 (N_12594,N_11273,N_11367);
or U12595 (N_12595,N_11321,N_11602);
or U12596 (N_12596,N_11713,N_11474);
or U12597 (N_12597,N_11343,N_11414);
nor U12598 (N_12598,N_11896,N_11744);
and U12599 (N_12599,N_11730,N_11366);
or U12600 (N_12600,N_11584,N_11393);
and U12601 (N_12601,N_11953,N_11328);
nand U12602 (N_12602,N_11961,N_11656);
or U12603 (N_12603,N_11826,N_11943);
nand U12604 (N_12604,N_11806,N_11840);
nand U12605 (N_12605,N_11261,N_11811);
nor U12606 (N_12606,N_11489,N_11881);
or U12607 (N_12607,N_11908,N_11825);
xnor U12608 (N_12608,N_11596,N_11407);
and U12609 (N_12609,N_11281,N_11285);
and U12610 (N_12610,N_11339,N_11425);
and U12611 (N_12611,N_11764,N_11532);
nor U12612 (N_12612,N_11756,N_11352);
nand U12613 (N_12613,N_11386,N_11614);
nor U12614 (N_12614,N_11771,N_11891);
or U12615 (N_12615,N_11670,N_11782);
or U12616 (N_12616,N_11580,N_11740);
nor U12617 (N_12617,N_11366,N_11900);
or U12618 (N_12618,N_11545,N_11984);
or U12619 (N_12619,N_11466,N_11938);
and U12620 (N_12620,N_11402,N_11379);
or U12621 (N_12621,N_11292,N_11497);
or U12622 (N_12622,N_11884,N_11329);
xor U12623 (N_12623,N_11715,N_11900);
and U12624 (N_12624,N_11963,N_11555);
nor U12625 (N_12625,N_11680,N_11392);
and U12626 (N_12626,N_11588,N_11846);
and U12627 (N_12627,N_11515,N_11851);
xor U12628 (N_12628,N_11700,N_11488);
or U12629 (N_12629,N_11893,N_11257);
nor U12630 (N_12630,N_11529,N_11887);
nor U12631 (N_12631,N_11550,N_11524);
nor U12632 (N_12632,N_11623,N_11661);
nand U12633 (N_12633,N_11543,N_11586);
nand U12634 (N_12634,N_11753,N_11888);
or U12635 (N_12635,N_11601,N_11980);
and U12636 (N_12636,N_11347,N_11905);
nor U12637 (N_12637,N_11895,N_11757);
or U12638 (N_12638,N_11414,N_11545);
xor U12639 (N_12639,N_11795,N_11508);
nor U12640 (N_12640,N_11376,N_11618);
xor U12641 (N_12641,N_11603,N_11568);
nand U12642 (N_12642,N_11499,N_11611);
nand U12643 (N_12643,N_11817,N_11450);
nor U12644 (N_12644,N_11485,N_11393);
and U12645 (N_12645,N_11743,N_11692);
and U12646 (N_12646,N_11361,N_11337);
nor U12647 (N_12647,N_11308,N_11793);
and U12648 (N_12648,N_11547,N_11986);
nand U12649 (N_12649,N_11406,N_11448);
and U12650 (N_12650,N_11315,N_11812);
nand U12651 (N_12651,N_11871,N_11473);
or U12652 (N_12652,N_11562,N_11940);
nand U12653 (N_12653,N_11307,N_11432);
nor U12654 (N_12654,N_11839,N_11447);
or U12655 (N_12655,N_11587,N_11580);
nor U12656 (N_12656,N_11531,N_11577);
or U12657 (N_12657,N_11665,N_11793);
and U12658 (N_12658,N_11837,N_11275);
or U12659 (N_12659,N_11545,N_11580);
nand U12660 (N_12660,N_11966,N_11986);
and U12661 (N_12661,N_11539,N_11540);
nand U12662 (N_12662,N_11663,N_11961);
xnor U12663 (N_12663,N_11958,N_11643);
or U12664 (N_12664,N_11888,N_11423);
and U12665 (N_12665,N_11738,N_11675);
and U12666 (N_12666,N_11960,N_11553);
nand U12667 (N_12667,N_11952,N_11416);
or U12668 (N_12668,N_11733,N_11284);
or U12669 (N_12669,N_11998,N_11798);
or U12670 (N_12670,N_11907,N_11454);
and U12671 (N_12671,N_11992,N_11687);
nor U12672 (N_12672,N_11705,N_11677);
nand U12673 (N_12673,N_11280,N_11723);
nand U12674 (N_12674,N_11252,N_11601);
and U12675 (N_12675,N_11580,N_11921);
or U12676 (N_12676,N_11682,N_11806);
nor U12677 (N_12677,N_11976,N_11714);
xnor U12678 (N_12678,N_11390,N_11370);
xor U12679 (N_12679,N_11480,N_11315);
and U12680 (N_12680,N_11272,N_11793);
or U12681 (N_12681,N_11515,N_11427);
nor U12682 (N_12682,N_11419,N_11538);
nor U12683 (N_12683,N_11412,N_11379);
nand U12684 (N_12684,N_11270,N_11700);
nor U12685 (N_12685,N_11898,N_11322);
or U12686 (N_12686,N_11760,N_11534);
or U12687 (N_12687,N_11958,N_11465);
nor U12688 (N_12688,N_11959,N_11436);
or U12689 (N_12689,N_11389,N_11347);
nor U12690 (N_12690,N_11665,N_11829);
nand U12691 (N_12691,N_11889,N_11658);
or U12692 (N_12692,N_11780,N_11558);
nor U12693 (N_12693,N_11491,N_11352);
nand U12694 (N_12694,N_11267,N_11905);
and U12695 (N_12695,N_11731,N_11781);
nor U12696 (N_12696,N_11960,N_11589);
nand U12697 (N_12697,N_11432,N_11617);
nor U12698 (N_12698,N_11344,N_11933);
and U12699 (N_12699,N_11745,N_11525);
or U12700 (N_12700,N_11790,N_11457);
or U12701 (N_12701,N_11597,N_11962);
nor U12702 (N_12702,N_11996,N_11593);
and U12703 (N_12703,N_11906,N_11526);
nor U12704 (N_12704,N_11708,N_11937);
and U12705 (N_12705,N_11526,N_11943);
nor U12706 (N_12706,N_11844,N_11422);
nor U12707 (N_12707,N_11751,N_11366);
nand U12708 (N_12708,N_11914,N_11309);
and U12709 (N_12709,N_11642,N_11571);
nor U12710 (N_12710,N_11788,N_11709);
xor U12711 (N_12711,N_11780,N_11952);
nor U12712 (N_12712,N_11481,N_11798);
or U12713 (N_12713,N_11658,N_11997);
xnor U12714 (N_12714,N_11520,N_11476);
and U12715 (N_12715,N_11644,N_11825);
nand U12716 (N_12716,N_11886,N_11356);
and U12717 (N_12717,N_11336,N_11847);
or U12718 (N_12718,N_11722,N_11895);
nor U12719 (N_12719,N_11365,N_11611);
nand U12720 (N_12720,N_11757,N_11824);
nand U12721 (N_12721,N_11925,N_11296);
xor U12722 (N_12722,N_11415,N_11828);
and U12723 (N_12723,N_11590,N_11626);
and U12724 (N_12724,N_11876,N_11526);
nor U12725 (N_12725,N_11508,N_11706);
and U12726 (N_12726,N_11316,N_11685);
or U12727 (N_12727,N_11594,N_11705);
nor U12728 (N_12728,N_11777,N_11799);
or U12729 (N_12729,N_11888,N_11999);
or U12730 (N_12730,N_11575,N_11490);
or U12731 (N_12731,N_11675,N_11548);
nand U12732 (N_12732,N_11437,N_11460);
nand U12733 (N_12733,N_11624,N_11572);
and U12734 (N_12734,N_11936,N_11461);
nand U12735 (N_12735,N_11863,N_11583);
nor U12736 (N_12736,N_11519,N_11593);
nand U12737 (N_12737,N_11789,N_11604);
and U12738 (N_12738,N_11674,N_11724);
nor U12739 (N_12739,N_11895,N_11351);
nor U12740 (N_12740,N_11304,N_11563);
and U12741 (N_12741,N_11930,N_11881);
nor U12742 (N_12742,N_11452,N_11387);
nor U12743 (N_12743,N_11443,N_11719);
or U12744 (N_12744,N_11370,N_11801);
or U12745 (N_12745,N_11440,N_11795);
nand U12746 (N_12746,N_11862,N_11962);
and U12747 (N_12747,N_11661,N_11527);
nor U12748 (N_12748,N_11558,N_11319);
and U12749 (N_12749,N_11964,N_11934);
xnor U12750 (N_12750,N_12012,N_12718);
nor U12751 (N_12751,N_12740,N_12246);
nor U12752 (N_12752,N_12702,N_12721);
or U12753 (N_12753,N_12212,N_12434);
and U12754 (N_12754,N_12198,N_12079);
xnor U12755 (N_12755,N_12714,N_12114);
nand U12756 (N_12756,N_12509,N_12228);
nor U12757 (N_12757,N_12322,N_12288);
or U12758 (N_12758,N_12572,N_12338);
and U12759 (N_12759,N_12620,N_12112);
or U12760 (N_12760,N_12124,N_12449);
or U12761 (N_12761,N_12276,N_12379);
nand U12762 (N_12762,N_12329,N_12066);
or U12763 (N_12763,N_12463,N_12367);
nand U12764 (N_12764,N_12452,N_12497);
nand U12765 (N_12765,N_12700,N_12389);
nor U12766 (N_12766,N_12024,N_12745);
or U12767 (N_12767,N_12377,N_12106);
and U12768 (N_12768,N_12720,N_12581);
nor U12769 (N_12769,N_12340,N_12564);
and U12770 (N_12770,N_12319,N_12400);
xor U12771 (N_12771,N_12614,N_12643);
or U12772 (N_12772,N_12371,N_12505);
nor U12773 (N_12773,N_12619,N_12575);
or U12774 (N_12774,N_12381,N_12680);
nand U12775 (N_12775,N_12477,N_12454);
nor U12776 (N_12776,N_12421,N_12468);
nor U12777 (N_12777,N_12683,N_12391);
nor U12778 (N_12778,N_12084,N_12686);
or U12779 (N_12779,N_12384,N_12334);
nor U12780 (N_12780,N_12439,N_12610);
xor U12781 (N_12781,N_12677,N_12524);
or U12782 (N_12782,N_12744,N_12169);
nor U12783 (N_12783,N_12215,N_12146);
or U12784 (N_12784,N_12107,N_12177);
or U12785 (N_12785,N_12690,N_12027);
xor U12786 (N_12786,N_12646,N_12402);
nor U12787 (N_12787,N_12166,N_12602);
or U12788 (N_12788,N_12360,N_12093);
nor U12789 (N_12789,N_12672,N_12474);
and U12790 (N_12790,N_12020,N_12021);
xor U12791 (N_12791,N_12386,N_12019);
nand U12792 (N_12792,N_12733,N_12565);
nor U12793 (N_12793,N_12137,N_12260);
xor U12794 (N_12794,N_12179,N_12640);
nand U12795 (N_12795,N_12015,N_12275);
and U12796 (N_12796,N_12070,N_12354);
nor U12797 (N_12797,N_12430,N_12533);
or U12798 (N_12798,N_12550,N_12213);
nor U12799 (N_12799,N_12647,N_12387);
or U12800 (N_12800,N_12577,N_12139);
and U12801 (N_12801,N_12111,N_12290);
nor U12802 (N_12802,N_12685,N_12715);
and U12803 (N_12803,N_12285,N_12464);
nand U12804 (N_12804,N_12521,N_12448);
nand U12805 (N_12805,N_12237,N_12703);
nor U12806 (N_12806,N_12664,N_12332);
nand U12807 (N_12807,N_12385,N_12480);
nor U12808 (N_12808,N_12182,N_12618);
nor U12809 (N_12809,N_12372,N_12238);
nor U12810 (N_12810,N_12206,N_12221);
nand U12811 (N_12811,N_12236,N_12369);
and U12812 (N_12812,N_12201,N_12743);
nand U12813 (N_12813,N_12002,N_12350);
nor U12814 (N_12814,N_12214,N_12692);
or U12815 (N_12815,N_12675,N_12525);
nor U12816 (N_12816,N_12028,N_12586);
nand U12817 (N_12817,N_12345,N_12527);
or U12818 (N_12818,N_12045,N_12574);
nor U12819 (N_12819,N_12348,N_12623);
nor U12820 (N_12820,N_12425,N_12063);
or U12821 (N_12821,N_12080,N_12263);
or U12822 (N_12822,N_12141,N_12416);
nor U12823 (N_12823,N_12712,N_12014);
xnor U12824 (N_12824,N_12138,N_12209);
nor U12825 (N_12825,N_12708,N_12711);
xnor U12826 (N_12826,N_12248,N_12026);
nor U12827 (N_12827,N_12540,N_12731);
and U12828 (N_12828,N_12053,N_12247);
nand U12829 (N_12829,N_12417,N_12515);
nor U12830 (N_12830,N_12038,N_12304);
and U12831 (N_12831,N_12429,N_12408);
nand U12832 (N_12832,N_12437,N_12520);
and U12833 (N_12833,N_12362,N_12481);
and U12834 (N_12834,N_12227,N_12202);
xnor U12835 (N_12835,N_12473,N_12424);
nor U12836 (N_12836,N_12398,N_12394);
nor U12837 (N_12837,N_12626,N_12642);
and U12838 (N_12838,N_12678,N_12067);
or U12839 (N_12839,N_12397,N_12605);
nor U12840 (N_12840,N_12644,N_12529);
and U12841 (N_12841,N_12055,N_12253);
nand U12842 (N_12842,N_12071,N_12608);
nand U12843 (N_12843,N_12327,N_12484);
and U12844 (N_12844,N_12315,N_12719);
or U12845 (N_12845,N_12735,N_12666);
nand U12846 (N_12846,N_12585,N_12631);
nor U12847 (N_12847,N_12530,N_12560);
and U12848 (N_12848,N_12208,N_12062);
nor U12849 (N_12849,N_12018,N_12162);
and U12850 (N_12850,N_12159,N_12029);
nand U12851 (N_12851,N_12134,N_12291);
and U12852 (N_12852,N_12493,N_12170);
nand U12853 (N_12853,N_12301,N_12030);
nor U12854 (N_12854,N_12051,N_12099);
nand U12855 (N_12855,N_12210,N_12292);
and U12856 (N_12856,N_12355,N_12578);
nand U12857 (N_12857,N_12659,N_12189);
nand U12858 (N_12858,N_12637,N_12031);
nand U12859 (N_12859,N_12219,N_12662);
or U12860 (N_12860,N_12569,N_12413);
nand U12861 (N_12861,N_12671,N_12616);
nand U12862 (N_12862,N_12097,N_12121);
xor U12863 (N_12863,N_12044,N_12503);
and U12864 (N_12864,N_12399,N_12588);
nor U12865 (N_12865,N_12042,N_12230);
and U12866 (N_12866,N_12054,N_12274);
or U12867 (N_12867,N_12440,N_12092);
or U12868 (N_12868,N_12245,N_12544);
nor U12869 (N_12869,N_12073,N_12115);
or U12870 (N_12870,N_12641,N_12376);
and U12871 (N_12871,N_12695,N_12669);
xnor U12872 (N_12872,N_12172,N_12725);
xnor U12873 (N_12873,N_12551,N_12010);
nand U12874 (N_12874,N_12232,N_12336);
nor U12875 (N_12875,N_12450,N_12507);
nand U12876 (N_12876,N_12432,N_12592);
nor U12877 (N_12877,N_12280,N_12059);
nand U12878 (N_12878,N_12052,N_12705);
and U12879 (N_12879,N_12456,N_12270);
nor U12880 (N_12880,N_12239,N_12240);
nor U12881 (N_12881,N_12127,N_12392);
nand U12882 (N_12882,N_12546,N_12074);
nand U12883 (N_12883,N_12674,N_12220);
xor U12884 (N_12884,N_12654,N_12483);
or U12885 (N_12885,N_12635,N_12361);
and U12886 (N_12886,N_12613,N_12748);
xnor U12887 (N_12887,N_12266,N_12258);
nand U12888 (N_12888,N_12118,N_12352);
or U12889 (N_12889,N_12409,N_12171);
or U12890 (N_12890,N_12086,N_12231);
and U12891 (N_12891,N_12412,N_12383);
or U12892 (N_12892,N_12682,N_12064);
or U12893 (N_12893,N_12713,N_12414);
nand U12894 (N_12894,N_12061,N_12607);
nand U12895 (N_12895,N_12341,N_12188);
or U12896 (N_12896,N_12007,N_12528);
nand U12897 (N_12897,N_12200,N_12223);
or U12898 (N_12898,N_12517,N_12005);
nor U12899 (N_12899,N_12296,N_12186);
and U12900 (N_12900,N_12445,N_12330);
nand U12901 (N_12901,N_12157,N_12308);
and U12902 (N_12902,N_12472,N_12536);
nor U12903 (N_12903,N_12573,N_12282);
or U12904 (N_12904,N_12289,N_12254);
xnor U12905 (N_12905,N_12558,N_12512);
nand U12906 (N_12906,N_12256,N_12150);
nor U12907 (N_12907,N_12582,N_12465);
nor U12908 (N_12908,N_12076,N_12023);
nand U12909 (N_12909,N_12225,N_12563);
nand U12910 (N_12910,N_12370,N_12504);
or U12911 (N_12911,N_12382,N_12511);
and U12912 (N_12912,N_12321,N_12749);
nor U12913 (N_12913,N_12436,N_12167);
or U12914 (N_12914,N_12668,N_12297);
or U12915 (N_12915,N_12462,N_12145);
or U12916 (N_12916,N_12155,N_12140);
and U12917 (N_12917,N_12226,N_12175);
nor U12918 (N_12918,N_12604,N_12197);
nand U12919 (N_12919,N_12309,N_12008);
nand U12920 (N_12920,N_12482,N_12455);
or U12921 (N_12921,N_12651,N_12557);
xor U12922 (N_12922,N_12670,N_12158);
or U12923 (N_12923,N_12707,N_12418);
and U12924 (N_12924,N_12621,N_12535);
nand U12925 (N_12925,N_12541,N_12013);
nand U12926 (N_12926,N_12698,N_12470);
and U12927 (N_12927,N_12571,N_12365);
or U12928 (N_12928,N_12595,N_12691);
or U12929 (N_12929,N_12356,N_12298);
or U12930 (N_12930,N_12261,N_12726);
or U12931 (N_12931,N_12277,N_12609);
or U12932 (N_12932,N_12148,N_12634);
nand U12933 (N_12933,N_12144,N_12438);
xnor U12934 (N_12934,N_12089,N_12344);
nor U12935 (N_12935,N_12057,N_12142);
and U12936 (N_12936,N_12469,N_12006);
and U12937 (N_12937,N_12410,N_12081);
or U12938 (N_12938,N_12694,N_12545);
or U12939 (N_12939,N_12561,N_12318);
or U12940 (N_12940,N_12194,N_12657);
nor U12941 (N_12941,N_12234,N_12443);
nand U12942 (N_12942,N_12229,N_12428);
and U12943 (N_12943,N_12181,N_12599);
nor U12944 (N_12944,N_12596,N_12326);
and U12945 (N_12945,N_12043,N_12101);
nand U12946 (N_12946,N_12501,N_12331);
xor U12947 (N_12947,N_12004,N_12629);
nand U12948 (N_12948,N_12730,N_12684);
and U12949 (N_12949,N_12312,N_12519);
or U12950 (N_12950,N_12126,N_12583);
and U12951 (N_12951,N_12192,N_12523);
and U12952 (N_12952,N_12632,N_12125);
or U12953 (N_12953,N_12660,N_12306);
or U12954 (N_12954,N_12034,N_12724);
nand U12955 (N_12955,N_12611,N_12337);
nor U12956 (N_12956,N_12153,N_12704);
and U12957 (N_12957,N_12508,N_12163);
nor U12958 (N_12958,N_12060,N_12050);
or U12959 (N_12959,N_12548,N_12461);
and U12960 (N_12960,N_12487,N_12349);
xnor U12961 (N_12961,N_12490,N_12269);
nand U12962 (N_12962,N_12734,N_12273);
nand U12963 (N_12963,N_12601,N_12451);
nand U12964 (N_12964,N_12267,N_12624);
and U12965 (N_12965,N_12491,N_12459);
or U12966 (N_12966,N_12554,N_12658);
nand U12967 (N_12967,N_12697,N_12593);
nor U12968 (N_12968,N_12078,N_12143);
or U12969 (N_12969,N_12566,N_12268);
nand U12970 (N_12970,N_12278,N_12420);
and U12971 (N_12971,N_12396,N_12555);
xnor U12972 (N_12972,N_12222,N_12403);
or U12973 (N_12973,N_12077,N_12722);
and U12974 (N_12974,N_12109,N_12591);
and U12975 (N_12975,N_12262,N_12532);
and U12976 (N_12976,N_12346,N_12649);
nor U12977 (N_12977,N_12590,N_12307);
or U12978 (N_12978,N_12617,N_12553);
nor U12979 (N_12979,N_12102,N_12040);
nor U12980 (N_12980,N_12567,N_12211);
xnor U12981 (N_12981,N_12305,N_12218);
nand U12982 (N_12982,N_12333,N_12217);
nand U12983 (N_12983,N_12184,N_12320);
and U12984 (N_12984,N_12423,N_12036);
and U12985 (N_12985,N_12688,N_12589);
nor U12986 (N_12986,N_12294,N_12736);
and U12987 (N_12987,N_12244,N_12747);
or U12988 (N_12988,N_12287,N_12363);
nor U12989 (N_12989,N_12433,N_12467);
nor U12990 (N_12990,N_12016,N_12046);
or U12991 (N_12991,N_12576,N_12131);
nor U12992 (N_12992,N_12441,N_12195);
xnor U12993 (N_12993,N_12281,N_12368);
or U12994 (N_12994,N_12233,N_12117);
or U12995 (N_12995,N_12009,N_12119);
nand U12996 (N_12996,N_12494,N_12580);
xor U12997 (N_12997,N_12431,N_12096);
or U12998 (N_12998,N_12375,N_12130);
and U12999 (N_12999,N_12422,N_12325);
nand U13000 (N_13000,N_12732,N_12500);
or U13001 (N_13001,N_12539,N_12559);
nand U13002 (N_13002,N_12098,N_12444);
and U13003 (N_13003,N_12435,N_12205);
or U13004 (N_13004,N_12633,N_12390);
nor U13005 (N_13005,N_12252,N_12068);
nand U13006 (N_13006,N_12419,N_12359);
nor U13007 (N_13007,N_12739,N_12627);
nand U13008 (N_13008,N_12286,N_12404);
xor U13009 (N_13009,N_12001,N_12011);
and U13010 (N_13010,N_12492,N_12049);
nand U13011 (N_13011,N_12639,N_12537);
nor U13012 (N_13012,N_12173,N_12105);
nor U13013 (N_13013,N_12295,N_12128);
nand U13014 (N_13014,N_12568,N_12056);
or U13015 (N_13015,N_12395,N_12082);
and U13016 (N_13016,N_12405,N_12193);
nand U13017 (N_13017,N_12625,N_12584);
and U13018 (N_13018,N_12693,N_12094);
or U13019 (N_13019,N_12090,N_12190);
xor U13020 (N_13020,N_12570,N_12699);
and U13021 (N_13021,N_12339,N_12709);
nand U13022 (N_13022,N_12746,N_12284);
and U13023 (N_13023,N_12710,N_12661);
nor U13024 (N_13024,N_12516,N_12676);
or U13025 (N_13025,N_12415,N_12513);
xnor U13026 (N_13026,N_12187,N_12207);
or U13027 (N_13027,N_12406,N_12728);
or U13028 (N_13028,N_12606,N_12191);
nand U13029 (N_13029,N_12265,N_12122);
nor U13030 (N_13030,N_12149,N_12241);
or U13031 (N_13031,N_12742,N_12185);
nand U13032 (N_13032,N_12302,N_12518);
nand U13033 (N_13033,N_12380,N_12579);
nor U13034 (N_13034,N_12072,N_12648);
nand U13035 (N_13035,N_12154,N_12120);
or U13036 (N_13036,N_12047,N_12499);
or U13037 (N_13037,N_12168,N_12108);
and U13038 (N_13038,N_12035,N_12373);
nor U13039 (N_13039,N_12393,N_12113);
xnor U13040 (N_13040,N_12314,N_12374);
nor U13041 (N_13041,N_12324,N_12317);
xor U13042 (N_13042,N_12542,N_12630);
or U13043 (N_13043,N_12135,N_12264);
nor U13044 (N_13044,N_12538,N_12032);
nand U13045 (N_13045,N_12116,N_12401);
or U13046 (N_13046,N_12594,N_12663);
and U13047 (N_13047,N_12597,N_12316);
nand U13048 (N_13048,N_12178,N_12033);
nand U13049 (N_13049,N_12272,N_12065);
nor U13050 (N_13050,N_12727,N_12151);
nor U13051 (N_13051,N_12347,N_12681);
xor U13052 (N_13052,N_12132,N_12510);
nand U13053 (N_13053,N_12088,N_12299);
or U13054 (N_13054,N_12216,N_12645);
xnor U13055 (N_13055,N_12471,N_12652);
or U13056 (N_13056,N_12453,N_12123);
nand U13057 (N_13057,N_12407,N_12242);
and U13058 (N_13058,N_12737,N_12095);
nand U13059 (N_13059,N_12104,N_12311);
and U13060 (N_13060,N_12701,N_12696);
or U13061 (N_13061,N_12328,N_12650);
xor U13062 (N_13062,N_12458,N_12196);
nand U13063 (N_13063,N_12653,N_12638);
or U13064 (N_13064,N_12343,N_12679);
nor U13065 (N_13065,N_12498,N_12156);
and U13066 (N_13066,N_12335,N_12665);
or U13067 (N_13067,N_12486,N_12488);
nor U13068 (N_13068,N_12556,N_12447);
and U13069 (N_13069,N_12534,N_12103);
nor U13070 (N_13070,N_12183,N_12017);
nand U13071 (N_13071,N_12723,N_12489);
nor U13072 (N_13072,N_12531,N_12366);
and U13073 (N_13073,N_12717,N_12543);
nand U13074 (N_13074,N_12475,N_12204);
nand U13075 (N_13075,N_12514,N_12176);
and U13076 (N_13076,N_12476,N_12075);
nor U13077 (N_13077,N_12741,N_12257);
nor U13078 (N_13078,N_12160,N_12342);
nor U13079 (N_13079,N_12037,N_12041);
xnor U13080 (N_13080,N_12495,N_12224);
and U13081 (N_13081,N_12351,N_12426);
or U13082 (N_13082,N_12069,N_12025);
and U13083 (N_13083,N_12249,N_12485);
and U13084 (N_13084,N_12587,N_12478);
nand U13085 (N_13085,N_12293,N_12667);
and U13086 (N_13086,N_12358,N_12378);
or U13087 (N_13087,N_12255,N_12243);
or U13088 (N_13088,N_12235,N_12622);
nand U13089 (N_13089,N_12313,N_12303);
nand U13090 (N_13090,N_12615,N_12388);
xnor U13091 (N_13091,N_12673,N_12110);
xor U13092 (N_13092,N_12522,N_12549);
and U13093 (N_13093,N_12048,N_12039);
nand U13094 (N_13094,N_12427,N_12457);
nor U13095 (N_13095,N_12600,N_12506);
and U13096 (N_13096,N_12687,N_12100);
or U13097 (N_13097,N_12466,N_12091);
and U13098 (N_13098,N_12655,N_12706);
nand U13099 (N_13099,N_12323,N_12562);
or U13100 (N_13100,N_12000,N_12628);
or U13101 (N_13101,N_12442,N_12598);
or U13102 (N_13102,N_12729,N_12129);
nor U13103 (N_13103,N_12259,N_12738);
nor U13104 (N_13104,N_12547,N_12526);
nand U13105 (N_13105,N_12460,N_12411);
nand U13106 (N_13106,N_12203,N_12003);
and U13107 (N_13107,N_12133,N_12174);
nor U13108 (N_13108,N_12085,N_12689);
nand U13109 (N_13109,N_12603,N_12310);
or U13110 (N_13110,N_12283,N_12612);
nor U13111 (N_13111,N_12300,N_12353);
or U13112 (N_13112,N_12656,N_12147);
nand U13113 (N_13113,N_12161,N_12446);
nand U13114 (N_13114,N_12087,N_12716);
xor U13115 (N_13115,N_12199,N_12022);
or U13116 (N_13116,N_12636,N_12152);
xor U13117 (N_13117,N_12279,N_12058);
or U13118 (N_13118,N_12479,N_12136);
and U13119 (N_13119,N_12502,N_12180);
or U13120 (N_13120,N_12552,N_12271);
and U13121 (N_13121,N_12250,N_12083);
and U13122 (N_13122,N_12496,N_12357);
nor U13123 (N_13123,N_12251,N_12165);
nand U13124 (N_13124,N_12364,N_12164);
or U13125 (N_13125,N_12394,N_12438);
xor U13126 (N_13126,N_12610,N_12621);
or U13127 (N_13127,N_12127,N_12540);
nand U13128 (N_13128,N_12446,N_12415);
and U13129 (N_13129,N_12544,N_12657);
nor U13130 (N_13130,N_12663,N_12238);
or U13131 (N_13131,N_12736,N_12361);
nor U13132 (N_13132,N_12160,N_12062);
and U13133 (N_13133,N_12450,N_12561);
or U13134 (N_13134,N_12434,N_12151);
nor U13135 (N_13135,N_12538,N_12552);
xor U13136 (N_13136,N_12722,N_12075);
nand U13137 (N_13137,N_12607,N_12240);
and U13138 (N_13138,N_12652,N_12607);
nand U13139 (N_13139,N_12651,N_12454);
nor U13140 (N_13140,N_12104,N_12724);
nor U13141 (N_13141,N_12735,N_12161);
nor U13142 (N_13142,N_12411,N_12678);
nor U13143 (N_13143,N_12093,N_12235);
nor U13144 (N_13144,N_12562,N_12329);
xor U13145 (N_13145,N_12174,N_12377);
and U13146 (N_13146,N_12572,N_12479);
or U13147 (N_13147,N_12610,N_12322);
and U13148 (N_13148,N_12084,N_12567);
and U13149 (N_13149,N_12489,N_12611);
or U13150 (N_13150,N_12282,N_12643);
or U13151 (N_13151,N_12700,N_12223);
nor U13152 (N_13152,N_12547,N_12478);
or U13153 (N_13153,N_12050,N_12635);
nor U13154 (N_13154,N_12346,N_12005);
or U13155 (N_13155,N_12577,N_12150);
nand U13156 (N_13156,N_12028,N_12029);
nand U13157 (N_13157,N_12037,N_12607);
and U13158 (N_13158,N_12478,N_12618);
and U13159 (N_13159,N_12122,N_12628);
nand U13160 (N_13160,N_12636,N_12568);
nand U13161 (N_13161,N_12600,N_12477);
or U13162 (N_13162,N_12257,N_12332);
and U13163 (N_13163,N_12233,N_12461);
and U13164 (N_13164,N_12524,N_12139);
and U13165 (N_13165,N_12414,N_12580);
and U13166 (N_13166,N_12023,N_12707);
or U13167 (N_13167,N_12566,N_12717);
nand U13168 (N_13168,N_12379,N_12155);
and U13169 (N_13169,N_12245,N_12227);
nand U13170 (N_13170,N_12681,N_12256);
and U13171 (N_13171,N_12358,N_12444);
and U13172 (N_13172,N_12564,N_12339);
and U13173 (N_13173,N_12286,N_12204);
nor U13174 (N_13174,N_12720,N_12223);
nand U13175 (N_13175,N_12077,N_12383);
xnor U13176 (N_13176,N_12315,N_12586);
xnor U13177 (N_13177,N_12712,N_12241);
and U13178 (N_13178,N_12415,N_12545);
nor U13179 (N_13179,N_12443,N_12589);
nand U13180 (N_13180,N_12513,N_12706);
or U13181 (N_13181,N_12214,N_12507);
or U13182 (N_13182,N_12590,N_12310);
or U13183 (N_13183,N_12448,N_12090);
nand U13184 (N_13184,N_12038,N_12715);
or U13185 (N_13185,N_12204,N_12426);
or U13186 (N_13186,N_12222,N_12711);
nand U13187 (N_13187,N_12559,N_12594);
nor U13188 (N_13188,N_12131,N_12065);
nand U13189 (N_13189,N_12253,N_12228);
and U13190 (N_13190,N_12049,N_12024);
nand U13191 (N_13191,N_12152,N_12507);
and U13192 (N_13192,N_12160,N_12441);
or U13193 (N_13193,N_12578,N_12058);
nor U13194 (N_13194,N_12363,N_12528);
nand U13195 (N_13195,N_12072,N_12246);
nand U13196 (N_13196,N_12156,N_12158);
nand U13197 (N_13197,N_12289,N_12708);
or U13198 (N_13198,N_12632,N_12552);
xor U13199 (N_13199,N_12416,N_12331);
nand U13200 (N_13200,N_12032,N_12424);
nand U13201 (N_13201,N_12212,N_12088);
or U13202 (N_13202,N_12591,N_12487);
or U13203 (N_13203,N_12572,N_12370);
xor U13204 (N_13204,N_12343,N_12084);
nand U13205 (N_13205,N_12555,N_12463);
xnor U13206 (N_13206,N_12500,N_12328);
nand U13207 (N_13207,N_12678,N_12508);
and U13208 (N_13208,N_12280,N_12370);
xor U13209 (N_13209,N_12063,N_12013);
and U13210 (N_13210,N_12241,N_12075);
or U13211 (N_13211,N_12577,N_12360);
or U13212 (N_13212,N_12329,N_12455);
and U13213 (N_13213,N_12610,N_12465);
or U13214 (N_13214,N_12243,N_12265);
and U13215 (N_13215,N_12062,N_12221);
and U13216 (N_13216,N_12071,N_12382);
and U13217 (N_13217,N_12089,N_12003);
and U13218 (N_13218,N_12141,N_12467);
nand U13219 (N_13219,N_12474,N_12212);
xor U13220 (N_13220,N_12386,N_12233);
or U13221 (N_13221,N_12681,N_12465);
and U13222 (N_13222,N_12264,N_12121);
or U13223 (N_13223,N_12061,N_12150);
or U13224 (N_13224,N_12103,N_12585);
or U13225 (N_13225,N_12420,N_12182);
and U13226 (N_13226,N_12569,N_12368);
or U13227 (N_13227,N_12679,N_12726);
or U13228 (N_13228,N_12691,N_12610);
and U13229 (N_13229,N_12722,N_12213);
nor U13230 (N_13230,N_12596,N_12511);
and U13231 (N_13231,N_12144,N_12025);
nand U13232 (N_13232,N_12480,N_12076);
xnor U13233 (N_13233,N_12526,N_12567);
nor U13234 (N_13234,N_12722,N_12418);
nand U13235 (N_13235,N_12213,N_12052);
nand U13236 (N_13236,N_12497,N_12407);
nor U13237 (N_13237,N_12195,N_12671);
or U13238 (N_13238,N_12630,N_12638);
nor U13239 (N_13239,N_12643,N_12537);
nand U13240 (N_13240,N_12148,N_12437);
and U13241 (N_13241,N_12533,N_12023);
or U13242 (N_13242,N_12266,N_12534);
and U13243 (N_13243,N_12701,N_12357);
or U13244 (N_13244,N_12172,N_12676);
nand U13245 (N_13245,N_12353,N_12528);
nand U13246 (N_13246,N_12700,N_12735);
nand U13247 (N_13247,N_12320,N_12615);
and U13248 (N_13248,N_12738,N_12024);
nor U13249 (N_13249,N_12733,N_12031);
nor U13250 (N_13250,N_12620,N_12277);
and U13251 (N_13251,N_12414,N_12572);
and U13252 (N_13252,N_12504,N_12394);
and U13253 (N_13253,N_12112,N_12616);
and U13254 (N_13254,N_12336,N_12425);
nor U13255 (N_13255,N_12729,N_12743);
xnor U13256 (N_13256,N_12580,N_12512);
and U13257 (N_13257,N_12710,N_12719);
and U13258 (N_13258,N_12276,N_12007);
or U13259 (N_13259,N_12693,N_12226);
nor U13260 (N_13260,N_12506,N_12318);
and U13261 (N_13261,N_12308,N_12259);
and U13262 (N_13262,N_12267,N_12070);
or U13263 (N_13263,N_12514,N_12741);
or U13264 (N_13264,N_12746,N_12523);
or U13265 (N_13265,N_12040,N_12298);
nor U13266 (N_13266,N_12077,N_12643);
nor U13267 (N_13267,N_12094,N_12470);
nor U13268 (N_13268,N_12409,N_12519);
and U13269 (N_13269,N_12045,N_12143);
or U13270 (N_13270,N_12244,N_12243);
nor U13271 (N_13271,N_12171,N_12367);
nor U13272 (N_13272,N_12718,N_12495);
and U13273 (N_13273,N_12035,N_12305);
nor U13274 (N_13274,N_12340,N_12585);
or U13275 (N_13275,N_12639,N_12672);
and U13276 (N_13276,N_12160,N_12593);
nand U13277 (N_13277,N_12069,N_12245);
nand U13278 (N_13278,N_12515,N_12378);
or U13279 (N_13279,N_12588,N_12221);
and U13280 (N_13280,N_12611,N_12295);
and U13281 (N_13281,N_12522,N_12582);
and U13282 (N_13282,N_12061,N_12133);
or U13283 (N_13283,N_12054,N_12244);
nor U13284 (N_13284,N_12534,N_12685);
nand U13285 (N_13285,N_12020,N_12099);
or U13286 (N_13286,N_12546,N_12215);
xor U13287 (N_13287,N_12424,N_12018);
nand U13288 (N_13288,N_12719,N_12065);
or U13289 (N_13289,N_12586,N_12057);
nand U13290 (N_13290,N_12685,N_12070);
or U13291 (N_13291,N_12622,N_12471);
nor U13292 (N_13292,N_12344,N_12106);
nand U13293 (N_13293,N_12154,N_12111);
nor U13294 (N_13294,N_12396,N_12623);
and U13295 (N_13295,N_12447,N_12136);
nor U13296 (N_13296,N_12177,N_12113);
nand U13297 (N_13297,N_12291,N_12144);
xnor U13298 (N_13298,N_12057,N_12090);
or U13299 (N_13299,N_12745,N_12462);
nor U13300 (N_13300,N_12397,N_12570);
or U13301 (N_13301,N_12379,N_12629);
nor U13302 (N_13302,N_12698,N_12493);
or U13303 (N_13303,N_12149,N_12604);
or U13304 (N_13304,N_12496,N_12390);
and U13305 (N_13305,N_12294,N_12517);
or U13306 (N_13306,N_12332,N_12223);
nor U13307 (N_13307,N_12573,N_12036);
or U13308 (N_13308,N_12105,N_12389);
nand U13309 (N_13309,N_12325,N_12482);
and U13310 (N_13310,N_12119,N_12128);
and U13311 (N_13311,N_12473,N_12232);
nor U13312 (N_13312,N_12193,N_12575);
nand U13313 (N_13313,N_12131,N_12320);
and U13314 (N_13314,N_12291,N_12682);
nor U13315 (N_13315,N_12505,N_12735);
and U13316 (N_13316,N_12326,N_12263);
xnor U13317 (N_13317,N_12749,N_12208);
or U13318 (N_13318,N_12539,N_12260);
and U13319 (N_13319,N_12006,N_12112);
or U13320 (N_13320,N_12552,N_12487);
and U13321 (N_13321,N_12480,N_12403);
xnor U13322 (N_13322,N_12207,N_12006);
nand U13323 (N_13323,N_12362,N_12596);
nand U13324 (N_13324,N_12349,N_12465);
and U13325 (N_13325,N_12232,N_12536);
nor U13326 (N_13326,N_12620,N_12427);
nor U13327 (N_13327,N_12249,N_12365);
nor U13328 (N_13328,N_12144,N_12433);
nor U13329 (N_13329,N_12739,N_12001);
xnor U13330 (N_13330,N_12693,N_12276);
nand U13331 (N_13331,N_12003,N_12251);
nor U13332 (N_13332,N_12132,N_12002);
nor U13333 (N_13333,N_12208,N_12379);
and U13334 (N_13334,N_12577,N_12053);
or U13335 (N_13335,N_12217,N_12626);
and U13336 (N_13336,N_12148,N_12542);
nand U13337 (N_13337,N_12659,N_12589);
and U13338 (N_13338,N_12554,N_12164);
or U13339 (N_13339,N_12011,N_12322);
nor U13340 (N_13340,N_12705,N_12114);
and U13341 (N_13341,N_12746,N_12706);
nand U13342 (N_13342,N_12177,N_12447);
xnor U13343 (N_13343,N_12253,N_12459);
nand U13344 (N_13344,N_12216,N_12629);
xor U13345 (N_13345,N_12304,N_12590);
and U13346 (N_13346,N_12544,N_12578);
nor U13347 (N_13347,N_12211,N_12694);
or U13348 (N_13348,N_12405,N_12053);
or U13349 (N_13349,N_12675,N_12716);
nand U13350 (N_13350,N_12353,N_12256);
or U13351 (N_13351,N_12351,N_12693);
nand U13352 (N_13352,N_12366,N_12019);
or U13353 (N_13353,N_12423,N_12123);
nand U13354 (N_13354,N_12427,N_12487);
or U13355 (N_13355,N_12748,N_12029);
nor U13356 (N_13356,N_12317,N_12205);
nand U13357 (N_13357,N_12499,N_12217);
nor U13358 (N_13358,N_12740,N_12461);
nand U13359 (N_13359,N_12574,N_12230);
nor U13360 (N_13360,N_12642,N_12308);
or U13361 (N_13361,N_12654,N_12407);
and U13362 (N_13362,N_12384,N_12178);
or U13363 (N_13363,N_12056,N_12495);
nand U13364 (N_13364,N_12395,N_12747);
nand U13365 (N_13365,N_12585,N_12502);
nor U13366 (N_13366,N_12269,N_12577);
or U13367 (N_13367,N_12714,N_12585);
nand U13368 (N_13368,N_12434,N_12351);
xor U13369 (N_13369,N_12231,N_12233);
nand U13370 (N_13370,N_12646,N_12059);
and U13371 (N_13371,N_12175,N_12285);
and U13372 (N_13372,N_12611,N_12173);
nand U13373 (N_13373,N_12464,N_12461);
nand U13374 (N_13374,N_12195,N_12498);
nor U13375 (N_13375,N_12173,N_12394);
or U13376 (N_13376,N_12088,N_12744);
and U13377 (N_13377,N_12567,N_12155);
and U13378 (N_13378,N_12433,N_12667);
nor U13379 (N_13379,N_12702,N_12221);
and U13380 (N_13380,N_12066,N_12459);
nor U13381 (N_13381,N_12425,N_12713);
or U13382 (N_13382,N_12210,N_12080);
nor U13383 (N_13383,N_12095,N_12583);
nand U13384 (N_13384,N_12042,N_12633);
xnor U13385 (N_13385,N_12303,N_12550);
and U13386 (N_13386,N_12094,N_12118);
nor U13387 (N_13387,N_12055,N_12452);
and U13388 (N_13388,N_12369,N_12091);
nor U13389 (N_13389,N_12712,N_12574);
or U13390 (N_13390,N_12252,N_12143);
nor U13391 (N_13391,N_12406,N_12211);
nand U13392 (N_13392,N_12540,N_12646);
nand U13393 (N_13393,N_12522,N_12547);
nand U13394 (N_13394,N_12241,N_12147);
or U13395 (N_13395,N_12615,N_12510);
xnor U13396 (N_13396,N_12345,N_12398);
and U13397 (N_13397,N_12634,N_12098);
nor U13398 (N_13398,N_12237,N_12620);
xnor U13399 (N_13399,N_12301,N_12586);
nor U13400 (N_13400,N_12462,N_12714);
or U13401 (N_13401,N_12129,N_12485);
and U13402 (N_13402,N_12725,N_12736);
nand U13403 (N_13403,N_12605,N_12744);
nand U13404 (N_13404,N_12034,N_12619);
and U13405 (N_13405,N_12209,N_12396);
or U13406 (N_13406,N_12391,N_12740);
or U13407 (N_13407,N_12068,N_12051);
or U13408 (N_13408,N_12073,N_12672);
nor U13409 (N_13409,N_12347,N_12521);
nor U13410 (N_13410,N_12526,N_12497);
nor U13411 (N_13411,N_12091,N_12265);
and U13412 (N_13412,N_12598,N_12049);
nor U13413 (N_13413,N_12131,N_12366);
and U13414 (N_13414,N_12191,N_12656);
nand U13415 (N_13415,N_12671,N_12450);
and U13416 (N_13416,N_12231,N_12602);
and U13417 (N_13417,N_12527,N_12517);
nor U13418 (N_13418,N_12372,N_12220);
nor U13419 (N_13419,N_12474,N_12477);
and U13420 (N_13420,N_12680,N_12168);
or U13421 (N_13421,N_12476,N_12504);
nor U13422 (N_13422,N_12452,N_12105);
nor U13423 (N_13423,N_12001,N_12154);
nand U13424 (N_13424,N_12611,N_12291);
or U13425 (N_13425,N_12049,N_12604);
xor U13426 (N_13426,N_12618,N_12641);
nor U13427 (N_13427,N_12609,N_12338);
nor U13428 (N_13428,N_12624,N_12205);
and U13429 (N_13429,N_12537,N_12588);
or U13430 (N_13430,N_12353,N_12257);
or U13431 (N_13431,N_12225,N_12174);
nand U13432 (N_13432,N_12570,N_12087);
and U13433 (N_13433,N_12470,N_12652);
and U13434 (N_13434,N_12262,N_12585);
and U13435 (N_13435,N_12724,N_12022);
nand U13436 (N_13436,N_12678,N_12721);
or U13437 (N_13437,N_12370,N_12083);
xnor U13438 (N_13438,N_12639,N_12581);
and U13439 (N_13439,N_12709,N_12155);
and U13440 (N_13440,N_12427,N_12630);
and U13441 (N_13441,N_12435,N_12698);
nor U13442 (N_13442,N_12492,N_12430);
or U13443 (N_13443,N_12602,N_12647);
or U13444 (N_13444,N_12446,N_12220);
nand U13445 (N_13445,N_12289,N_12260);
nor U13446 (N_13446,N_12086,N_12344);
xor U13447 (N_13447,N_12542,N_12726);
nor U13448 (N_13448,N_12258,N_12324);
and U13449 (N_13449,N_12465,N_12549);
or U13450 (N_13450,N_12471,N_12502);
nor U13451 (N_13451,N_12645,N_12507);
nand U13452 (N_13452,N_12481,N_12124);
nor U13453 (N_13453,N_12305,N_12716);
nor U13454 (N_13454,N_12528,N_12428);
and U13455 (N_13455,N_12648,N_12101);
and U13456 (N_13456,N_12037,N_12696);
and U13457 (N_13457,N_12225,N_12598);
and U13458 (N_13458,N_12550,N_12513);
nand U13459 (N_13459,N_12199,N_12245);
or U13460 (N_13460,N_12700,N_12055);
and U13461 (N_13461,N_12424,N_12214);
nand U13462 (N_13462,N_12034,N_12376);
nand U13463 (N_13463,N_12686,N_12447);
nor U13464 (N_13464,N_12235,N_12458);
nand U13465 (N_13465,N_12457,N_12306);
nand U13466 (N_13466,N_12334,N_12675);
and U13467 (N_13467,N_12222,N_12473);
nand U13468 (N_13468,N_12683,N_12394);
and U13469 (N_13469,N_12247,N_12010);
xor U13470 (N_13470,N_12444,N_12701);
and U13471 (N_13471,N_12099,N_12475);
nand U13472 (N_13472,N_12570,N_12712);
nor U13473 (N_13473,N_12039,N_12717);
and U13474 (N_13474,N_12574,N_12498);
or U13475 (N_13475,N_12686,N_12660);
or U13476 (N_13476,N_12306,N_12699);
nor U13477 (N_13477,N_12154,N_12749);
nor U13478 (N_13478,N_12233,N_12405);
nor U13479 (N_13479,N_12416,N_12702);
or U13480 (N_13480,N_12612,N_12093);
nand U13481 (N_13481,N_12109,N_12110);
nand U13482 (N_13482,N_12471,N_12705);
nor U13483 (N_13483,N_12650,N_12003);
or U13484 (N_13484,N_12656,N_12709);
nor U13485 (N_13485,N_12440,N_12590);
and U13486 (N_13486,N_12534,N_12519);
nand U13487 (N_13487,N_12543,N_12015);
and U13488 (N_13488,N_12717,N_12255);
nor U13489 (N_13489,N_12350,N_12200);
nand U13490 (N_13490,N_12062,N_12461);
nor U13491 (N_13491,N_12382,N_12133);
or U13492 (N_13492,N_12311,N_12085);
nor U13493 (N_13493,N_12259,N_12527);
nand U13494 (N_13494,N_12124,N_12739);
or U13495 (N_13495,N_12114,N_12124);
xnor U13496 (N_13496,N_12145,N_12483);
nand U13497 (N_13497,N_12607,N_12690);
nor U13498 (N_13498,N_12706,N_12478);
nand U13499 (N_13499,N_12206,N_12661);
nor U13500 (N_13500,N_13143,N_12823);
and U13501 (N_13501,N_13057,N_13369);
nor U13502 (N_13502,N_13333,N_12880);
nor U13503 (N_13503,N_13210,N_12911);
nor U13504 (N_13504,N_13317,N_13176);
and U13505 (N_13505,N_13257,N_13116);
or U13506 (N_13506,N_13404,N_12955);
nand U13507 (N_13507,N_13073,N_12957);
nand U13508 (N_13508,N_13277,N_13487);
nand U13509 (N_13509,N_13020,N_13008);
xnor U13510 (N_13510,N_13196,N_12865);
nand U13511 (N_13511,N_12815,N_13035);
nand U13512 (N_13512,N_13198,N_13163);
xor U13513 (N_13513,N_13131,N_12978);
and U13514 (N_13514,N_12894,N_13078);
nand U13515 (N_13515,N_13280,N_12867);
xnor U13516 (N_13516,N_13040,N_13119);
nor U13517 (N_13517,N_13009,N_13170);
nor U13518 (N_13518,N_13217,N_12993);
nand U13519 (N_13519,N_13301,N_13357);
nand U13520 (N_13520,N_12877,N_12977);
and U13521 (N_13521,N_13000,N_13449);
nor U13522 (N_13522,N_12839,N_13265);
or U13523 (N_13523,N_13007,N_13208);
nor U13524 (N_13524,N_12754,N_13160);
nor U13525 (N_13525,N_12797,N_13367);
xnor U13526 (N_13526,N_12898,N_12924);
and U13527 (N_13527,N_13370,N_12936);
and U13528 (N_13528,N_13183,N_13074);
nor U13529 (N_13529,N_12963,N_13106);
nor U13530 (N_13530,N_12767,N_12775);
xor U13531 (N_13531,N_12975,N_12835);
nand U13532 (N_13532,N_13383,N_13118);
xor U13533 (N_13533,N_13019,N_13068);
or U13534 (N_13534,N_13394,N_13438);
or U13535 (N_13535,N_12989,N_13366);
and U13536 (N_13536,N_12812,N_12793);
or U13537 (N_13537,N_13085,N_12813);
or U13538 (N_13538,N_13220,N_12832);
nor U13539 (N_13539,N_13485,N_13330);
nor U13540 (N_13540,N_13016,N_13222);
nor U13541 (N_13541,N_12984,N_13046);
nand U13542 (N_13542,N_13410,N_12808);
or U13543 (N_13543,N_12805,N_12946);
nor U13544 (N_13544,N_12872,N_12964);
and U13545 (N_13545,N_13181,N_12971);
nor U13546 (N_13546,N_13060,N_13308);
and U13547 (N_13547,N_12822,N_13499);
nand U13548 (N_13548,N_12795,N_13380);
and U13549 (N_13549,N_13470,N_12926);
xor U13550 (N_13550,N_13031,N_13364);
or U13551 (N_13551,N_13336,N_13407);
xnor U13552 (N_13552,N_12837,N_13032);
xnor U13553 (N_13553,N_13324,N_13295);
nor U13554 (N_13554,N_13150,N_13134);
nand U13555 (N_13555,N_13197,N_13465);
xor U13556 (N_13556,N_13092,N_13152);
nand U13557 (N_13557,N_12856,N_13224);
nor U13558 (N_13558,N_13123,N_13193);
nor U13559 (N_13559,N_13023,N_13212);
or U13560 (N_13560,N_12786,N_13345);
nand U13561 (N_13561,N_13065,N_12902);
nand U13562 (N_13562,N_13325,N_12806);
and U13563 (N_13563,N_13294,N_13088);
nand U13564 (N_13564,N_13115,N_13351);
or U13565 (N_13565,N_12962,N_12779);
and U13566 (N_13566,N_12966,N_12769);
nor U13567 (N_13567,N_12937,N_13232);
nand U13568 (N_13568,N_13080,N_13406);
nor U13569 (N_13569,N_12969,N_13390);
or U13570 (N_13570,N_13296,N_13306);
or U13571 (N_13571,N_12914,N_13273);
nand U13572 (N_13572,N_13056,N_13275);
or U13573 (N_13573,N_12776,N_13488);
nor U13574 (N_13574,N_13248,N_13025);
or U13575 (N_13575,N_13493,N_13077);
or U13576 (N_13576,N_12942,N_12884);
nand U13577 (N_13577,N_13028,N_13148);
or U13578 (N_13578,N_12757,N_13090);
nand U13579 (N_13579,N_13043,N_13290);
or U13580 (N_13580,N_13192,N_13200);
xnor U13581 (N_13581,N_12860,N_13374);
and U13582 (N_13582,N_13014,N_12778);
nor U13583 (N_13583,N_13352,N_13135);
nor U13584 (N_13584,N_12829,N_13133);
and U13585 (N_13585,N_13162,N_13399);
nand U13586 (N_13586,N_13318,N_13288);
nor U13587 (N_13587,N_13376,N_13218);
and U13588 (N_13588,N_12974,N_12930);
and U13589 (N_13589,N_13356,N_12932);
and U13590 (N_13590,N_13066,N_12929);
or U13591 (N_13591,N_12782,N_13262);
or U13592 (N_13592,N_13342,N_12814);
nor U13593 (N_13593,N_13417,N_13063);
nand U13594 (N_13594,N_13484,N_12997);
nor U13595 (N_13595,N_13483,N_13423);
or U13596 (N_13596,N_13132,N_13076);
nor U13597 (N_13597,N_13253,N_13221);
and U13598 (N_13598,N_12792,N_13419);
xor U13599 (N_13599,N_13079,N_13363);
or U13600 (N_13600,N_13326,N_13069);
nand U13601 (N_13601,N_13051,N_13332);
and U13602 (N_13602,N_12934,N_12896);
or U13603 (N_13603,N_12887,N_12931);
nor U13604 (N_13604,N_12922,N_13486);
nor U13605 (N_13605,N_13034,N_13341);
or U13606 (N_13606,N_13395,N_12921);
and U13607 (N_13607,N_12999,N_12770);
and U13608 (N_13608,N_13256,N_13497);
and U13609 (N_13609,N_13124,N_13282);
nor U13610 (N_13610,N_13235,N_12824);
or U13611 (N_13611,N_13434,N_13234);
and U13612 (N_13612,N_12866,N_13393);
and U13613 (N_13613,N_13489,N_12892);
and U13614 (N_13614,N_12886,N_13409);
or U13615 (N_13615,N_13446,N_13140);
xnor U13616 (N_13616,N_13316,N_13284);
xnor U13617 (N_13617,N_13379,N_13418);
nand U13618 (N_13618,N_13261,N_12842);
or U13619 (N_13619,N_13474,N_13071);
nor U13620 (N_13620,N_13335,N_12980);
nand U13621 (N_13621,N_12817,N_13315);
or U13622 (N_13622,N_13189,N_13471);
nor U13623 (N_13623,N_13044,N_13378);
nor U13624 (N_13624,N_13322,N_13203);
and U13625 (N_13625,N_12952,N_13178);
xnor U13626 (N_13626,N_13155,N_12855);
nor U13627 (N_13627,N_12753,N_13024);
or U13628 (N_13628,N_12756,N_13478);
xor U13629 (N_13629,N_13440,N_13302);
nand U13630 (N_13630,N_13182,N_13303);
nand U13631 (N_13631,N_13084,N_13388);
nor U13632 (N_13632,N_12983,N_13297);
and U13633 (N_13633,N_13445,N_12916);
nor U13634 (N_13634,N_13236,N_12882);
nand U13635 (N_13635,N_13039,N_12816);
and U13636 (N_13636,N_13138,N_13319);
nor U13637 (N_13637,N_13067,N_13139);
xnor U13638 (N_13638,N_13185,N_13444);
nand U13639 (N_13639,N_13095,N_12825);
nor U13640 (N_13640,N_12947,N_13158);
or U13641 (N_13641,N_12888,N_12958);
nor U13642 (N_13642,N_12994,N_13225);
nor U13643 (N_13643,N_12927,N_13207);
nor U13644 (N_13644,N_12986,N_13100);
nand U13645 (N_13645,N_13242,N_12948);
nand U13646 (N_13646,N_12868,N_13396);
or U13647 (N_13647,N_13012,N_13428);
nand U13648 (N_13648,N_12871,N_13432);
and U13649 (N_13649,N_13430,N_13146);
or U13650 (N_13650,N_12920,N_13001);
or U13651 (N_13651,N_13172,N_13006);
or U13652 (N_13652,N_13168,N_12838);
nand U13653 (N_13653,N_12833,N_12849);
xnor U13654 (N_13654,N_13350,N_12847);
nand U13655 (N_13655,N_13461,N_13015);
and U13656 (N_13656,N_12878,N_12939);
and U13657 (N_13657,N_12979,N_13424);
and U13658 (N_13658,N_13468,N_12845);
or U13659 (N_13659,N_13433,N_12961);
and U13660 (N_13660,N_13187,N_13425);
or U13661 (N_13661,N_12791,N_13223);
or U13662 (N_13662,N_13002,N_12897);
xnor U13663 (N_13663,N_13266,N_12843);
and U13664 (N_13664,N_13321,N_13018);
xor U13665 (N_13665,N_13269,N_12900);
nand U13666 (N_13666,N_13102,N_13191);
nand U13667 (N_13667,N_13400,N_13240);
nand U13668 (N_13668,N_12945,N_13239);
nand U13669 (N_13669,N_12834,N_13128);
nor U13670 (N_13670,N_13287,N_13070);
nor U13671 (N_13671,N_12876,N_13348);
nor U13672 (N_13672,N_13258,N_13320);
or U13673 (N_13673,N_12774,N_12850);
nand U13674 (N_13674,N_13202,N_13246);
or U13675 (N_13675,N_13346,N_13021);
and U13676 (N_13676,N_12851,N_13011);
nand U13677 (N_13677,N_12803,N_12827);
or U13678 (N_13678,N_13405,N_13227);
xnor U13679 (N_13679,N_13381,N_13270);
nand U13680 (N_13680,N_13099,N_12991);
nor U13681 (N_13681,N_13205,N_13122);
and U13682 (N_13682,N_13129,N_13037);
nand U13683 (N_13683,N_13004,N_13165);
or U13684 (N_13684,N_13450,N_12759);
nor U13685 (N_13685,N_13110,N_12996);
or U13686 (N_13686,N_13447,N_12809);
xnor U13687 (N_13687,N_13451,N_13293);
or U13688 (N_13688,N_13403,N_12857);
nand U13689 (N_13689,N_12826,N_12790);
nand U13690 (N_13690,N_13490,N_13093);
nor U13691 (N_13691,N_12773,N_12766);
or U13692 (N_13692,N_12982,N_13109);
nand U13693 (N_13693,N_13286,N_13309);
and U13694 (N_13694,N_13173,N_12933);
and U13695 (N_13695,N_13368,N_13384);
xor U13696 (N_13696,N_13463,N_12819);
and U13697 (N_13697,N_13121,N_13083);
nand U13698 (N_13698,N_12859,N_12828);
or U13699 (N_13699,N_12789,N_13130);
or U13700 (N_13700,N_13199,N_13114);
nand U13701 (N_13701,N_12893,N_12970);
or U13702 (N_13702,N_12908,N_12863);
and U13703 (N_13703,N_13254,N_13229);
and U13704 (N_13704,N_13372,N_13473);
or U13705 (N_13705,N_13245,N_13142);
nor U13706 (N_13706,N_13094,N_13312);
xnor U13707 (N_13707,N_13013,N_13408);
or U13708 (N_13708,N_13375,N_13492);
nor U13709 (N_13709,N_13010,N_13329);
nor U13710 (N_13710,N_13355,N_12919);
and U13711 (N_13711,N_12990,N_13300);
and U13712 (N_13712,N_13476,N_13215);
nor U13713 (N_13713,N_13491,N_13052);
and U13714 (N_13714,N_13081,N_12917);
nand U13715 (N_13715,N_13310,N_13238);
xnor U13716 (N_13716,N_12804,N_13264);
xor U13717 (N_13717,N_12821,N_13059);
nor U13718 (N_13718,N_12788,N_13371);
nand U13719 (N_13719,N_13125,N_13331);
and U13720 (N_13720,N_12903,N_13214);
and U13721 (N_13721,N_12846,N_13481);
and U13722 (N_13722,N_12852,N_12771);
nand U13723 (N_13723,N_13472,N_13112);
nor U13724 (N_13724,N_12895,N_13382);
nor U13725 (N_13725,N_13047,N_13340);
and U13726 (N_13726,N_13460,N_12758);
nand U13727 (N_13727,N_13454,N_13466);
and U13728 (N_13728,N_13111,N_12784);
xnor U13729 (N_13729,N_13360,N_13285);
or U13730 (N_13730,N_13219,N_13443);
and U13731 (N_13731,N_13086,N_13391);
nor U13732 (N_13732,N_12940,N_13108);
nor U13733 (N_13733,N_13030,N_13247);
nand U13734 (N_13734,N_13343,N_13036);
and U13735 (N_13735,N_13482,N_13347);
xnor U13736 (N_13736,N_13353,N_13233);
or U13737 (N_13737,N_13213,N_13190);
nor U13738 (N_13738,N_13464,N_12915);
xnor U13739 (N_13739,N_13278,N_13362);
nand U13740 (N_13740,N_12901,N_13361);
xor U13741 (N_13741,N_13276,N_13429);
and U13742 (N_13742,N_12765,N_12751);
nand U13743 (N_13743,N_12889,N_13026);
and U13744 (N_13744,N_13274,N_13082);
and U13745 (N_13745,N_13305,N_13180);
or U13746 (N_13746,N_13103,N_12874);
nand U13747 (N_13747,N_13201,N_12883);
nor U13748 (N_13748,N_13439,N_13050);
or U13749 (N_13749,N_12862,N_13149);
nor U13750 (N_13750,N_13249,N_12972);
nor U13751 (N_13751,N_13161,N_12885);
nand U13752 (N_13752,N_12909,N_13053);
nand U13753 (N_13753,N_12953,N_12956);
and U13754 (N_13754,N_12800,N_12905);
and U13755 (N_13755,N_12959,N_12841);
or U13756 (N_13756,N_13027,N_13412);
nor U13757 (N_13757,N_12910,N_12873);
nand U13758 (N_13758,N_12864,N_12950);
or U13759 (N_13759,N_12985,N_13307);
nor U13760 (N_13760,N_13153,N_12807);
nand U13761 (N_13761,N_13188,N_13064);
nor U13762 (N_13762,N_13328,N_13054);
xor U13763 (N_13763,N_12987,N_13281);
xnor U13764 (N_13764,N_13147,N_12879);
nand U13765 (N_13765,N_13091,N_13255);
nor U13766 (N_13766,N_12943,N_12907);
and U13767 (N_13767,N_13211,N_12935);
or U13768 (N_13768,N_12928,N_13299);
nor U13769 (N_13769,N_12861,N_13479);
and U13770 (N_13770,N_13292,N_13159);
or U13771 (N_13771,N_13387,N_12798);
nor U13772 (N_13772,N_12763,N_12944);
nor U13773 (N_13773,N_13107,N_13174);
nand U13774 (N_13774,N_12941,N_12760);
or U13775 (N_13775,N_13414,N_13420);
nor U13776 (N_13776,N_12768,N_13327);
xnor U13777 (N_13777,N_12906,N_13459);
or U13778 (N_13778,N_12870,N_13415);
nand U13779 (N_13779,N_13096,N_13113);
nor U13780 (N_13780,N_13137,N_12831);
xor U13781 (N_13781,N_13061,N_13151);
nand U13782 (N_13782,N_12891,N_13386);
xor U13783 (N_13783,N_13228,N_12811);
nand U13784 (N_13784,N_13045,N_13495);
and U13785 (N_13785,N_13055,N_13344);
nand U13786 (N_13786,N_13298,N_13283);
xnor U13787 (N_13787,N_13049,N_12787);
xnor U13788 (N_13788,N_13421,N_13475);
or U13789 (N_13789,N_13209,N_13365);
xnor U13790 (N_13790,N_12995,N_13494);
xor U13791 (N_13791,N_12976,N_13289);
nand U13792 (N_13792,N_13029,N_13177);
nor U13793 (N_13793,N_13260,N_13358);
xor U13794 (N_13794,N_13338,N_12992);
xor U13795 (N_13795,N_13157,N_13042);
nor U13796 (N_13796,N_12918,N_12899);
or U13797 (N_13797,N_12780,N_12848);
nor U13798 (N_13798,N_13455,N_13431);
nor U13799 (N_13799,N_13437,N_13272);
nand U13800 (N_13800,N_13164,N_12853);
or U13801 (N_13801,N_12912,N_13398);
or U13802 (N_13802,N_13003,N_13062);
nand U13803 (N_13803,N_13075,N_12783);
nand U13804 (N_13804,N_13349,N_12761);
nor U13805 (N_13805,N_12799,N_13268);
or U13806 (N_13806,N_13204,N_13373);
nor U13807 (N_13807,N_13462,N_12794);
and U13808 (N_13808,N_13104,N_13179);
nand U13809 (N_13809,N_12954,N_13435);
or U13810 (N_13810,N_13105,N_13477);
and U13811 (N_13811,N_13101,N_12810);
nand U13812 (N_13812,N_13279,N_13389);
nand U13813 (N_13813,N_12781,N_13154);
nand U13814 (N_13814,N_13456,N_13231);
nand U13815 (N_13815,N_13314,N_12973);
nor U13816 (N_13816,N_12836,N_12796);
or U13817 (N_13817,N_13156,N_13241);
or U13818 (N_13818,N_13167,N_13136);
nor U13819 (N_13819,N_13498,N_12802);
nand U13820 (N_13820,N_13041,N_12777);
nor U13821 (N_13821,N_13145,N_13448);
nand U13822 (N_13822,N_13359,N_13323);
or U13823 (N_13823,N_13243,N_12960);
and U13824 (N_13824,N_12904,N_13097);
nand U13825 (N_13825,N_12830,N_13339);
nor U13826 (N_13826,N_13033,N_13271);
xor U13827 (N_13827,N_13291,N_13457);
and U13828 (N_13828,N_13166,N_13171);
nor U13829 (N_13829,N_12925,N_12875);
or U13830 (N_13830,N_13117,N_13252);
and U13831 (N_13831,N_13126,N_12801);
nand U13832 (N_13832,N_12755,N_12968);
nor U13833 (N_13833,N_13397,N_13334);
nand U13834 (N_13834,N_13251,N_12890);
and U13835 (N_13835,N_13442,N_12750);
nor U13836 (N_13836,N_13127,N_13458);
nand U13837 (N_13837,N_12844,N_12840);
and U13838 (N_13838,N_13402,N_13226);
and U13839 (N_13839,N_13436,N_13422);
or U13840 (N_13840,N_13392,N_13230);
and U13841 (N_13841,N_13195,N_13496);
xnor U13842 (N_13842,N_13005,N_12998);
nor U13843 (N_13843,N_13048,N_13141);
nand U13844 (N_13844,N_12938,N_13263);
or U13845 (N_13845,N_13022,N_12772);
xnor U13846 (N_13846,N_13377,N_13206);
or U13847 (N_13847,N_13089,N_13441);
and U13848 (N_13848,N_13267,N_13144);
or U13849 (N_13849,N_13186,N_12988);
nor U13850 (N_13850,N_13237,N_13453);
nand U13851 (N_13851,N_13216,N_13244);
nor U13852 (N_13852,N_13427,N_13480);
and U13853 (N_13853,N_12854,N_12820);
and U13854 (N_13854,N_13426,N_12762);
nor U13855 (N_13855,N_13017,N_13194);
and U13856 (N_13856,N_13467,N_12981);
nor U13857 (N_13857,N_13385,N_12965);
nor U13858 (N_13858,N_13304,N_12869);
or U13859 (N_13859,N_13354,N_12967);
xnor U13860 (N_13860,N_13072,N_13098);
nand U13861 (N_13861,N_12949,N_13169);
xor U13862 (N_13862,N_12785,N_12752);
nor U13863 (N_13863,N_13469,N_12923);
nor U13864 (N_13864,N_12858,N_13250);
nor U13865 (N_13865,N_13038,N_12818);
and U13866 (N_13866,N_12913,N_12881);
nor U13867 (N_13867,N_13452,N_13120);
or U13868 (N_13868,N_13175,N_12951);
nor U13869 (N_13869,N_13411,N_12764);
xnor U13870 (N_13870,N_13413,N_13311);
and U13871 (N_13871,N_13313,N_13058);
nand U13872 (N_13872,N_13416,N_13087);
nor U13873 (N_13873,N_13401,N_13259);
xor U13874 (N_13874,N_13184,N_13337);
nand U13875 (N_13875,N_12854,N_13341);
and U13876 (N_13876,N_12964,N_13272);
xor U13877 (N_13877,N_12857,N_13061);
nand U13878 (N_13878,N_13042,N_12755);
nand U13879 (N_13879,N_13418,N_12872);
nor U13880 (N_13880,N_13181,N_13205);
xnor U13881 (N_13881,N_13335,N_13338);
nand U13882 (N_13882,N_13155,N_12787);
and U13883 (N_13883,N_13240,N_13245);
nand U13884 (N_13884,N_12934,N_13297);
nor U13885 (N_13885,N_12924,N_13390);
nand U13886 (N_13886,N_13014,N_13212);
nand U13887 (N_13887,N_12894,N_13138);
xnor U13888 (N_13888,N_12844,N_13262);
nor U13889 (N_13889,N_13026,N_13350);
nand U13890 (N_13890,N_13332,N_12910);
nor U13891 (N_13891,N_13005,N_13358);
or U13892 (N_13892,N_13463,N_12762);
nand U13893 (N_13893,N_13229,N_12812);
nor U13894 (N_13894,N_13147,N_12834);
xor U13895 (N_13895,N_13369,N_13473);
nand U13896 (N_13896,N_13137,N_13329);
nand U13897 (N_13897,N_12990,N_13321);
and U13898 (N_13898,N_13359,N_12887);
xnor U13899 (N_13899,N_12889,N_12876);
and U13900 (N_13900,N_12861,N_13054);
nor U13901 (N_13901,N_13350,N_13496);
nor U13902 (N_13902,N_12852,N_12839);
nor U13903 (N_13903,N_12792,N_12933);
nor U13904 (N_13904,N_12918,N_13100);
nand U13905 (N_13905,N_12910,N_13330);
or U13906 (N_13906,N_13373,N_13226);
and U13907 (N_13907,N_13024,N_13137);
or U13908 (N_13908,N_13401,N_12937);
or U13909 (N_13909,N_12917,N_12935);
xor U13910 (N_13910,N_13071,N_13115);
and U13911 (N_13911,N_13439,N_13494);
nand U13912 (N_13912,N_13121,N_13040);
nor U13913 (N_13913,N_13013,N_13427);
nand U13914 (N_13914,N_13297,N_13426);
nor U13915 (N_13915,N_12811,N_13409);
nand U13916 (N_13916,N_12974,N_12852);
and U13917 (N_13917,N_13458,N_13185);
xnor U13918 (N_13918,N_13440,N_13107);
and U13919 (N_13919,N_13391,N_13022);
nand U13920 (N_13920,N_12920,N_12767);
and U13921 (N_13921,N_12865,N_12902);
and U13922 (N_13922,N_12856,N_12804);
nor U13923 (N_13923,N_12991,N_13461);
nand U13924 (N_13924,N_13104,N_12983);
or U13925 (N_13925,N_13215,N_13207);
nor U13926 (N_13926,N_12964,N_12781);
nor U13927 (N_13927,N_12951,N_13406);
xnor U13928 (N_13928,N_13082,N_12894);
xor U13929 (N_13929,N_12983,N_13125);
nor U13930 (N_13930,N_13283,N_13070);
nand U13931 (N_13931,N_13147,N_12919);
nand U13932 (N_13932,N_13012,N_13165);
or U13933 (N_13933,N_13407,N_13161);
and U13934 (N_13934,N_13127,N_12933);
or U13935 (N_13935,N_13177,N_13489);
and U13936 (N_13936,N_12753,N_13170);
nor U13937 (N_13937,N_13436,N_12849);
nor U13938 (N_13938,N_13395,N_13270);
or U13939 (N_13939,N_13262,N_13238);
or U13940 (N_13940,N_13121,N_13044);
nand U13941 (N_13941,N_13216,N_13338);
and U13942 (N_13942,N_12913,N_13104);
xor U13943 (N_13943,N_12856,N_13244);
xor U13944 (N_13944,N_13094,N_13105);
or U13945 (N_13945,N_13364,N_13304);
or U13946 (N_13946,N_12780,N_12766);
nand U13947 (N_13947,N_13444,N_13323);
nor U13948 (N_13948,N_13037,N_12927);
or U13949 (N_13949,N_12922,N_12864);
nor U13950 (N_13950,N_13485,N_12761);
nand U13951 (N_13951,N_12899,N_13433);
xnor U13952 (N_13952,N_12946,N_13257);
nand U13953 (N_13953,N_13326,N_12791);
nor U13954 (N_13954,N_13177,N_13122);
xor U13955 (N_13955,N_12854,N_12802);
and U13956 (N_13956,N_12982,N_13080);
nand U13957 (N_13957,N_12982,N_13102);
and U13958 (N_13958,N_13457,N_12953);
or U13959 (N_13959,N_13489,N_13448);
and U13960 (N_13960,N_13133,N_13458);
or U13961 (N_13961,N_13424,N_13095);
and U13962 (N_13962,N_13215,N_12884);
nand U13963 (N_13963,N_13142,N_13256);
nand U13964 (N_13964,N_13287,N_12847);
nor U13965 (N_13965,N_12992,N_13016);
or U13966 (N_13966,N_13148,N_13261);
nand U13967 (N_13967,N_13341,N_13489);
or U13968 (N_13968,N_12793,N_13214);
nand U13969 (N_13969,N_12974,N_13372);
xor U13970 (N_13970,N_13474,N_13316);
and U13971 (N_13971,N_12818,N_13100);
or U13972 (N_13972,N_12849,N_13172);
nand U13973 (N_13973,N_13433,N_13022);
nand U13974 (N_13974,N_13191,N_12895);
nor U13975 (N_13975,N_13137,N_13228);
and U13976 (N_13976,N_13328,N_13329);
nor U13977 (N_13977,N_13133,N_12862);
nor U13978 (N_13978,N_13272,N_13405);
nor U13979 (N_13979,N_12848,N_13036);
xor U13980 (N_13980,N_12840,N_12913);
and U13981 (N_13981,N_13375,N_12889);
or U13982 (N_13982,N_13477,N_12762);
and U13983 (N_13983,N_12838,N_13150);
nand U13984 (N_13984,N_13290,N_13215);
xnor U13985 (N_13985,N_12931,N_13122);
xor U13986 (N_13986,N_12945,N_13383);
nand U13987 (N_13987,N_12835,N_13257);
or U13988 (N_13988,N_13142,N_13487);
and U13989 (N_13989,N_13257,N_13021);
nor U13990 (N_13990,N_13000,N_13365);
nor U13991 (N_13991,N_12799,N_13186);
or U13992 (N_13992,N_12815,N_13117);
and U13993 (N_13993,N_13142,N_12804);
xnor U13994 (N_13994,N_12911,N_12783);
nor U13995 (N_13995,N_12774,N_13011);
nand U13996 (N_13996,N_13410,N_13335);
nand U13997 (N_13997,N_13239,N_12868);
or U13998 (N_13998,N_13076,N_13121);
and U13999 (N_13999,N_13347,N_13256);
or U14000 (N_14000,N_12806,N_12903);
nand U14001 (N_14001,N_13182,N_13133);
or U14002 (N_14002,N_13025,N_12951);
and U14003 (N_14003,N_13336,N_12975);
and U14004 (N_14004,N_12768,N_12946);
nand U14005 (N_14005,N_12833,N_12982);
nor U14006 (N_14006,N_12839,N_13147);
nand U14007 (N_14007,N_13476,N_12805);
xnor U14008 (N_14008,N_13318,N_13033);
or U14009 (N_14009,N_13137,N_13084);
nand U14010 (N_14010,N_13003,N_12950);
and U14011 (N_14011,N_13225,N_12766);
xnor U14012 (N_14012,N_13284,N_12839);
nand U14013 (N_14013,N_13314,N_13097);
nand U14014 (N_14014,N_13089,N_13057);
or U14015 (N_14015,N_13208,N_13165);
and U14016 (N_14016,N_12835,N_12921);
and U14017 (N_14017,N_12808,N_12872);
and U14018 (N_14018,N_13366,N_12993);
nor U14019 (N_14019,N_13467,N_12771);
nand U14020 (N_14020,N_13235,N_12755);
or U14021 (N_14021,N_13086,N_13156);
and U14022 (N_14022,N_13222,N_12853);
nand U14023 (N_14023,N_12961,N_13058);
or U14024 (N_14024,N_12960,N_13048);
nor U14025 (N_14025,N_13442,N_12983);
or U14026 (N_14026,N_13181,N_13266);
and U14027 (N_14027,N_13252,N_13032);
nor U14028 (N_14028,N_12862,N_13219);
nand U14029 (N_14029,N_13041,N_13088);
nor U14030 (N_14030,N_13112,N_13174);
or U14031 (N_14031,N_13333,N_12851);
nor U14032 (N_14032,N_12779,N_12785);
nand U14033 (N_14033,N_13126,N_12951);
nor U14034 (N_14034,N_13253,N_12958);
nand U14035 (N_14035,N_12798,N_13140);
and U14036 (N_14036,N_12763,N_13218);
or U14037 (N_14037,N_12896,N_13214);
or U14038 (N_14038,N_12883,N_12971);
or U14039 (N_14039,N_13039,N_13033);
nor U14040 (N_14040,N_13007,N_12959);
nor U14041 (N_14041,N_13151,N_13174);
nand U14042 (N_14042,N_13044,N_12811);
and U14043 (N_14043,N_13184,N_13393);
and U14044 (N_14044,N_13014,N_12922);
xor U14045 (N_14045,N_13074,N_13188);
nand U14046 (N_14046,N_13343,N_12833);
nor U14047 (N_14047,N_13155,N_13009);
and U14048 (N_14048,N_13339,N_13200);
or U14049 (N_14049,N_13383,N_12919);
or U14050 (N_14050,N_13428,N_13135);
nand U14051 (N_14051,N_13378,N_13497);
or U14052 (N_14052,N_13430,N_13041);
nor U14053 (N_14053,N_12963,N_13244);
and U14054 (N_14054,N_13258,N_13303);
nand U14055 (N_14055,N_12901,N_13226);
xnor U14056 (N_14056,N_12751,N_12862);
and U14057 (N_14057,N_13456,N_12754);
nand U14058 (N_14058,N_13188,N_13108);
or U14059 (N_14059,N_13496,N_13327);
xnor U14060 (N_14060,N_12913,N_12756);
and U14061 (N_14061,N_12916,N_12896);
nand U14062 (N_14062,N_12870,N_13341);
or U14063 (N_14063,N_12961,N_13417);
or U14064 (N_14064,N_13033,N_13143);
nand U14065 (N_14065,N_13397,N_13405);
nand U14066 (N_14066,N_13395,N_13252);
and U14067 (N_14067,N_12788,N_13315);
nand U14068 (N_14068,N_13421,N_13191);
nor U14069 (N_14069,N_12945,N_12770);
and U14070 (N_14070,N_13069,N_13098);
nor U14071 (N_14071,N_13447,N_12842);
and U14072 (N_14072,N_12881,N_13404);
nor U14073 (N_14073,N_13439,N_13045);
and U14074 (N_14074,N_13340,N_13292);
xor U14075 (N_14075,N_13460,N_13181);
nor U14076 (N_14076,N_13418,N_12873);
xnor U14077 (N_14077,N_13273,N_13272);
nor U14078 (N_14078,N_13275,N_13168);
nand U14079 (N_14079,N_13186,N_13477);
nor U14080 (N_14080,N_12870,N_12781);
or U14081 (N_14081,N_13204,N_13000);
and U14082 (N_14082,N_13191,N_13261);
nor U14083 (N_14083,N_12926,N_13072);
or U14084 (N_14084,N_13355,N_13131);
and U14085 (N_14085,N_13043,N_13376);
or U14086 (N_14086,N_12884,N_12754);
or U14087 (N_14087,N_13360,N_13433);
nand U14088 (N_14088,N_13432,N_13226);
nand U14089 (N_14089,N_13210,N_12994);
or U14090 (N_14090,N_13261,N_13154);
nor U14091 (N_14091,N_13277,N_13483);
nor U14092 (N_14092,N_12966,N_13413);
or U14093 (N_14093,N_13129,N_13243);
or U14094 (N_14094,N_13113,N_12750);
or U14095 (N_14095,N_13327,N_13253);
nor U14096 (N_14096,N_13141,N_12952);
or U14097 (N_14097,N_12853,N_13187);
and U14098 (N_14098,N_13209,N_13070);
and U14099 (N_14099,N_13394,N_12908);
nor U14100 (N_14100,N_12896,N_12974);
nor U14101 (N_14101,N_13260,N_13199);
or U14102 (N_14102,N_13192,N_13303);
and U14103 (N_14103,N_13315,N_13168);
and U14104 (N_14104,N_13285,N_13314);
nand U14105 (N_14105,N_12851,N_13009);
and U14106 (N_14106,N_13292,N_13143);
or U14107 (N_14107,N_13286,N_12964);
or U14108 (N_14108,N_13120,N_13084);
and U14109 (N_14109,N_13327,N_13435);
or U14110 (N_14110,N_12817,N_13063);
and U14111 (N_14111,N_13241,N_12829);
nand U14112 (N_14112,N_13248,N_13313);
nand U14113 (N_14113,N_13451,N_13274);
xnor U14114 (N_14114,N_12843,N_13449);
nand U14115 (N_14115,N_13499,N_13165);
nor U14116 (N_14116,N_13189,N_13074);
xor U14117 (N_14117,N_13347,N_13064);
or U14118 (N_14118,N_12873,N_13331);
nor U14119 (N_14119,N_13015,N_13190);
and U14120 (N_14120,N_13043,N_13257);
nand U14121 (N_14121,N_13462,N_13183);
or U14122 (N_14122,N_13310,N_13272);
or U14123 (N_14123,N_13435,N_13149);
and U14124 (N_14124,N_13372,N_13392);
xnor U14125 (N_14125,N_13392,N_13068);
nor U14126 (N_14126,N_12988,N_13331);
nor U14127 (N_14127,N_13074,N_13083);
or U14128 (N_14128,N_13200,N_13142);
nor U14129 (N_14129,N_13260,N_13134);
nor U14130 (N_14130,N_12951,N_13354);
and U14131 (N_14131,N_12848,N_13264);
nor U14132 (N_14132,N_12966,N_13388);
nand U14133 (N_14133,N_13272,N_13149);
or U14134 (N_14134,N_12879,N_12921);
nor U14135 (N_14135,N_12827,N_13332);
xnor U14136 (N_14136,N_13027,N_12897);
and U14137 (N_14137,N_12945,N_13240);
nand U14138 (N_14138,N_12924,N_13215);
nand U14139 (N_14139,N_13307,N_12962);
nor U14140 (N_14140,N_13000,N_12966);
nand U14141 (N_14141,N_12887,N_13321);
nor U14142 (N_14142,N_13483,N_12842);
xnor U14143 (N_14143,N_13363,N_13254);
nor U14144 (N_14144,N_13336,N_13377);
nor U14145 (N_14145,N_13489,N_13068);
xnor U14146 (N_14146,N_13331,N_13152);
and U14147 (N_14147,N_13272,N_12797);
xnor U14148 (N_14148,N_13318,N_13363);
nor U14149 (N_14149,N_12905,N_13162);
and U14150 (N_14150,N_13431,N_13159);
and U14151 (N_14151,N_12966,N_13481);
nor U14152 (N_14152,N_13228,N_13441);
nor U14153 (N_14153,N_12776,N_13282);
nand U14154 (N_14154,N_13377,N_13026);
nand U14155 (N_14155,N_13257,N_13256);
nand U14156 (N_14156,N_13122,N_13077);
nor U14157 (N_14157,N_12810,N_12905);
or U14158 (N_14158,N_13236,N_12947);
or U14159 (N_14159,N_13392,N_12975);
and U14160 (N_14160,N_13197,N_13447);
nand U14161 (N_14161,N_12993,N_13307);
nor U14162 (N_14162,N_12965,N_13071);
xnor U14163 (N_14163,N_12997,N_12821);
or U14164 (N_14164,N_13083,N_13263);
nand U14165 (N_14165,N_13401,N_12995);
and U14166 (N_14166,N_13407,N_13060);
and U14167 (N_14167,N_12759,N_13419);
nor U14168 (N_14168,N_12871,N_12795);
nand U14169 (N_14169,N_13334,N_12875);
nor U14170 (N_14170,N_12901,N_13214);
or U14171 (N_14171,N_13375,N_13017);
or U14172 (N_14172,N_13118,N_12868);
xnor U14173 (N_14173,N_12839,N_12751);
and U14174 (N_14174,N_12873,N_12854);
xor U14175 (N_14175,N_13015,N_13434);
or U14176 (N_14176,N_13268,N_13408);
nand U14177 (N_14177,N_13041,N_13302);
or U14178 (N_14178,N_13285,N_13028);
nor U14179 (N_14179,N_12776,N_13457);
and U14180 (N_14180,N_13015,N_13228);
nand U14181 (N_14181,N_12793,N_12871);
and U14182 (N_14182,N_13135,N_13318);
or U14183 (N_14183,N_13339,N_12944);
and U14184 (N_14184,N_13169,N_12950);
and U14185 (N_14185,N_13264,N_13084);
or U14186 (N_14186,N_12812,N_13135);
xor U14187 (N_14187,N_12826,N_13055);
nand U14188 (N_14188,N_13212,N_13026);
and U14189 (N_14189,N_13258,N_13087);
nor U14190 (N_14190,N_12768,N_12797);
or U14191 (N_14191,N_13093,N_12799);
nor U14192 (N_14192,N_13436,N_13276);
nor U14193 (N_14193,N_13327,N_12937);
nor U14194 (N_14194,N_13227,N_12878);
or U14195 (N_14195,N_13244,N_13055);
nand U14196 (N_14196,N_13154,N_12775);
nand U14197 (N_14197,N_12825,N_13044);
nand U14198 (N_14198,N_13271,N_13120);
nor U14199 (N_14199,N_13298,N_13231);
or U14200 (N_14200,N_12953,N_13295);
or U14201 (N_14201,N_13448,N_13485);
nor U14202 (N_14202,N_13177,N_13167);
or U14203 (N_14203,N_12779,N_13041);
or U14204 (N_14204,N_13266,N_12854);
xnor U14205 (N_14205,N_12942,N_13254);
and U14206 (N_14206,N_12763,N_13345);
nor U14207 (N_14207,N_13391,N_12981);
xnor U14208 (N_14208,N_12801,N_13349);
nand U14209 (N_14209,N_13477,N_13026);
nor U14210 (N_14210,N_13054,N_13418);
nand U14211 (N_14211,N_13049,N_12763);
and U14212 (N_14212,N_13212,N_13131);
nor U14213 (N_14213,N_13306,N_12763);
or U14214 (N_14214,N_13010,N_13291);
nand U14215 (N_14215,N_13282,N_12916);
or U14216 (N_14216,N_12979,N_13339);
xor U14217 (N_14217,N_12795,N_12964);
nand U14218 (N_14218,N_12933,N_13249);
xnor U14219 (N_14219,N_13115,N_12892);
and U14220 (N_14220,N_12957,N_12978);
or U14221 (N_14221,N_13274,N_13428);
nor U14222 (N_14222,N_12856,N_13213);
or U14223 (N_14223,N_13162,N_13028);
and U14224 (N_14224,N_13090,N_12904);
or U14225 (N_14225,N_12960,N_12837);
or U14226 (N_14226,N_13417,N_13432);
nor U14227 (N_14227,N_13130,N_13315);
nor U14228 (N_14228,N_13055,N_12905);
nor U14229 (N_14229,N_12828,N_13234);
nor U14230 (N_14230,N_13024,N_13327);
xor U14231 (N_14231,N_12985,N_13442);
xnor U14232 (N_14232,N_13392,N_13444);
or U14233 (N_14233,N_13111,N_13105);
xnor U14234 (N_14234,N_12989,N_12761);
and U14235 (N_14235,N_12996,N_12903);
nand U14236 (N_14236,N_13009,N_12956);
nand U14237 (N_14237,N_12960,N_13459);
or U14238 (N_14238,N_13143,N_13490);
and U14239 (N_14239,N_13483,N_13175);
xnor U14240 (N_14240,N_13344,N_13323);
nand U14241 (N_14241,N_12779,N_12834);
nand U14242 (N_14242,N_12996,N_12974);
nor U14243 (N_14243,N_12844,N_13164);
nand U14244 (N_14244,N_13349,N_13330);
nand U14245 (N_14245,N_13271,N_13414);
and U14246 (N_14246,N_13366,N_13147);
and U14247 (N_14247,N_12851,N_12752);
or U14248 (N_14248,N_13462,N_13352);
nand U14249 (N_14249,N_12969,N_12784);
or U14250 (N_14250,N_13592,N_13832);
nor U14251 (N_14251,N_13600,N_13655);
and U14252 (N_14252,N_13939,N_13801);
nor U14253 (N_14253,N_13649,N_13741);
nor U14254 (N_14254,N_13734,N_13959);
and U14255 (N_14255,N_14062,N_13578);
nand U14256 (N_14256,N_13763,N_13597);
or U14257 (N_14257,N_13598,N_13602);
and U14258 (N_14258,N_13569,N_13586);
or U14259 (N_14259,N_13718,N_13761);
nand U14260 (N_14260,N_13888,N_14202);
nand U14261 (N_14261,N_13962,N_13944);
nor U14262 (N_14262,N_13582,N_13704);
or U14263 (N_14263,N_13806,N_13587);
nor U14264 (N_14264,N_13816,N_13936);
and U14265 (N_14265,N_13781,N_14088);
nor U14266 (N_14266,N_13844,N_13515);
and U14267 (N_14267,N_13839,N_13966);
nand U14268 (N_14268,N_13957,N_13529);
or U14269 (N_14269,N_14086,N_13846);
nor U14270 (N_14270,N_13681,N_13548);
nor U14271 (N_14271,N_13782,N_13774);
and U14272 (N_14272,N_14130,N_14229);
and U14273 (N_14273,N_13794,N_13532);
nand U14274 (N_14274,N_14230,N_13986);
or U14275 (N_14275,N_13983,N_14096);
xor U14276 (N_14276,N_13510,N_13715);
nand U14277 (N_14277,N_13685,N_14220);
nand U14278 (N_14278,N_13500,N_13536);
nor U14279 (N_14279,N_13948,N_13893);
xor U14280 (N_14280,N_13615,N_14067);
or U14281 (N_14281,N_14239,N_13753);
nor U14282 (N_14282,N_13621,N_13706);
or U14283 (N_14283,N_14007,N_14002);
and U14284 (N_14284,N_13736,N_14189);
nor U14285 (N_14285,N_14206,N_13691);
or U14286 (N_14286,N_14053,N_14183);
or U14287 (N_14287,N_13538,N_13512);
and U14288 (N_14288,N_13778,N_13757);
nand U14289 (N_14289,N_14033,N_13735);
and U14290 (N_14290,N_13814,N_14232);
nor U14291 (N_14291,N_13988,N_13863);
or U14292 (N_14292,N_13932,N_14186);
nand U14293 (N_14293,N_13913,N_13656);
or U14294 (N_14294,N_13915,N_14208);
and U14295 (N_14295,N_13613,N_14029);
nand U14296 (N_14296,N_13584,N_14132);
and U14297 (N_14297,N_13564,N_13835);
nor U14298 (N_14298,N_14171,N_14081);
and U14299 (N_14299,N_13730,N_13777);
and U14300 (N_14300,N_13865,N_14050);
nor U14301 (N_14301,N_13698,N_13935);
or U14302 (N_14302,N_13511,N_14179);
nor U14303 (N_14303,N_13754,N_14082);
or U14304 (N_14304,N_13747,N_13544);
nor U14305 (N_14305,N_13560,N_13922);
nand U14306 (N_14306,N_13599,N_13501);
or U14307 (N_14307,N_13860,N_13993);
and U14308 (N_14308,N_13628,N_13851);
nand U14309 (N_14309,N_13738,N_13834);
xnor U14310 (N_14310,N_13841,N_14187);
and U14311 (N_14311,N_14219,N_14165);
xor U14312 (N_14312,N_13929,N_14175);
nand U14313 (N_14313,N_14017,N_13967);
or U14314 (N_14314,N_14172,N_14233);
nand U14315 (N_14315,N_14091,N_13750);
and U14316 (N_14316,N_13588,N_13854);
nand U14317 (N_14317,N_14238,N_14185);
and U14318 (N_14318,N_13696,N_13953);
nand U14319 (N_14319,N_13614,N_13881);
or U14320 (N_14320,N_14072,N_13815);
xnor U14321 (N_14321,N_13675,N_13665);
nor U14322 (N_14322,N_13961,N_13596);
or U14323 (N_14323,N_14222,N_14032);
nor U14324 (N_14324,N_14008,N_13925);
or U14325 (N_14325,N_13687,N_13508);
nand U14326 (N_14326,N_13629,N_13589);
nor U14327 (N_14327,N_13673,N_13910);
xnor U14328 (N_14328,N_13810,N_14076);
xnor U14329 (N_14329,N_14136,N_14163);
or U14330 (N_14330,N_14031,N_13987);
nand U14331 (N_14331,N_14043,N_14231);
nand U14332 (N_14332,N_14077,N_13612);
xnor U14333 (N_14333,N_13547,N_14237);
nand U14334 (N_14334,N_14235,N_13573);
nor U14335 (N_14335,N_13697,N_13765);
nor U14336 (N_14336,N_13688,N_13693);
or U14337 (N_14337,N_14041,N_13570);
nand U14338 (N_14338,N_13581,N_14228);
nor U14339 (N_14339,N_13566,N_13633);
xnor U14340 (N_14340,N_14169,N_14211);
or U14341 (N_14341,N_13772,N_13546);
nand U14342 (N_14342,N_13620,N_13768);
nand U14343 (N_14343,N_13965,N_13664);
nor U14344 (N_14344,N_13514,N_13800);
nand U14345 (N_14345,N_13686,N_14184);
nand U14346 (N_14346,N_14097,N_13767);
and U14347 (N_14347,N_14178,N_13574);
nand U14348 (N_14348,N_14010,N_13725);
nand U14349 (N_14349,N_14161,N_13904);
and U14350 (N_14350,N_13876,N_13674);
nor U14351 (N_14351,N_14193,N_13836);
or U14352 (N_14352,N_13700,N_13997);
nor U14353 (N_14353,N_13733,N_14103);
nor U14354 (N_14354,N_13912,N_13737);
nand U14355 (N_14355,N_13504,N_13606);
nand U14356 (N_14356,N_13891,N_14106);
xnor U14357 (N_14357,N_14071,N_13872);
and U14358 (N_14358,N_14117,N_14047);
nor U14359 (N_14359,N_13918,N_13792);
xor U14360 (N_14360,N_13521,N_14131);
and U14361 (N_14361,N_13684,N_13826);
nand U14362 (N_14362,N_14196,N_14110);
nand U14363 (N_14363,N_13603,N_13857);
and U14364 (N_14364,N_13746,N_14099);
or U14365 (N_14365,N_13722,N_13954);
or U14366 (N_14366,N_14013,N_13601);
nand U14367 (N_14367,N_14227,N_14123);
nor U14368 (N_14368,N_13678,N_13712);
or U14369 (N_14369,N_13805,N_14248);
xnor U14370 (N_14370,N_13727,N_13917);
or U14371 (N_14371,N_13642,N_13764);
nor U14372 (N_14372,N_13632,N_13883);
nand U14373 (N_14373,N_13644,N_13790);
nor U14374 (N_14374,N_14079,N_13553);
nand U14375 (N_14375,N_14061,N_14089);
nand U14376 (N_14376,N_13695,N_14138);
xor U14377 (N_14377,N_14129,N_14141);
or U14378 (N_14378,N_14027,N_13776);
nor U14379 (N_14379,N_13568,N_14157);
nand U14380 (N_14380,N_13523,N_14014);
nand U14381 (N_14381,N_14118,N_13923);
or U14382 (N_14382,N_13880,N_14198);
nand U14383 (N_14383,N_14162,N_14003);
nor U14384 (N_14384,N_13572,N_14217);
nand U14385 (N_14385,N_13847,N_13711);
or U14386 (N_14386,N_13975,N_13540);
and U14387 (N_14387,N_13769,N_13518);
nor U14388 (N_14388,N_14149,N_14052);
nor U14389 (N_14389,N_13797,N_14034);
and U14390 (N_14390,N_14153,N_13885);
or U14391 (N_14391,N_13676,N_13626);
xnor U14392 (N_14392,N_13899,N_14049);
or U14393 (N_14393,N_13634,N_13969);
nand U14394 (N_14394,N_14207,N_13978);
nor U14395 (N_14395,N_14212,N_13798);
or U14396 (N_14396,N_13989,N_13580);
and U14397 (N_14397,N_13622,N_13624);
nor U14398 (N_14398,N_13985,N_13946);
nor U14399 (N_14399,N_14016,N_14065);
nor U14400 (N_14400,N_13708,N_13701);
and U14401 (N_14401,N_14126,N_13562);
and U14402 (N_14402,N_13783,N_13709);
xor U14403 (N_14403,N_13808,N_13981);
xor U14404 (N_14404,N_13551,N_13831);
and U14405 (N_14405,N_14009,N_13739);
nor U14406 (N_14406,N_13611,N_13968);
and U14407 (N_14407,N_13575,N_13652);
nor U14408 (N_14408,N_13856,N_13919);
or U14409 (N_14409,N_13577,N_13550);
nor U14410 (N_14410,N_13503,N_13623);
or U14411 (N_14411,N_13920,N_14194);
nor U14412 (N_14412,N_13994,N_13963);
nand U14413 (N_14413,N_14001,N_13571);
nor U14414 (N_14414,N_13554,N_13583);
or U14415 (N_14415,N_13506,N_14226);
and U14416 (N_14416,N_13639,N_13533);
nor U14417 (N_14417,N_13534,N_13850);
or U14418 (N_14418,N_13972,N_13648);
nor U14419 (N_14419,N_13595,N_14063);
xor U14420 (N_14420,N_14215,N_14247);
nor U14421 (N_14421,N_14104,N_13990);
nand U14422 (N_14422,N_14214,N_13974);
or U14423 (N_14423,N_13998,N_13682);
nor U14424 (N_14424,N_14221,N_14024);
nor U14425 (N_14425,N_13822,N_14197);
nor U14426 (N_14426,N_13567,N_13666);
or U14427 (N_14427,N_14241,N_14135);
and U14428 (N_14428,N_13813,N_13819);
nor U14429 (N_14429,N_13887,N_13651);
nand U14430 (N_14430,N_13619,N_14018);
nor U14431 (N_14431,N_13520,N_14218);
or U14432 (N_14432,N_13896,N_13947);
and U14433 (N_14433,N_13517,N_14203);
and U14434 (N_14434,N_13977,N_14160);
or U14435 (N_14435,N_14245,N_13799);
xor U14436 (N_14436,N_13849,N_14200);
xor U14437 (N_14437,N_13837,N_13852);
xnor U14438 (N_14438,N_13809,N_13579);
nand U14439 (N_14439,N_13627,N_14026);
nor U14440 (N_14440,N_13661,N_14045);
nand U14441 (N_14441,N_14069,N_13759);
or U14442 (N_14442,N_13535,N_13662);
or U14443 (N_14443,N_13758,N_13549);
and U14444 (N_14444,N_13869,N_13667);
xnor U14445 (N_14445,N_13779,N_14058);
nand U14446 (N_14446,N_14246,N_13565);
nor U14447 (N_14447,N_13949,N_13672);
and U14448 (N_14448,N_13898,N_13690);
nand U14449 (N_14449,N_13890,N_14124);
nor U14450 (N_14450,N_13911,N_14073);
and U14451 (N_14451,N_13897,N_14068);
and U14452 (N_14452,N_13559,N_13663);
nand U14453 (N_14453,N_13650,N_13745);
xor U14454 (N_14454,N_13970,N_14121);
and U14455 (N_14455,N_13821,N_14119);
nand U14456 (N_14456,N_14087,N_14066);
or U14457 (N_14457,N_14075,N_13740);
xor U14458 (N_14458,N_13960,N_13908);
or U14459 (N_14459,N_13845,N_13921);
or U14460 (N_14460,N_14039,N_13882);
nand U14461 (N_14461,N_14225,N_14004);
nand U14462 (N_14462,N_14036,N_13552);
and U14463 (N_14463,N_14152,N_14107);
nor U14464 (N_14464,N_14191,N_13817);
or U14465 (N_14465,N_14046,N_13771);
or U14466 (N_14466,N_14105,N_13905);
nand U14467 (N_14467,N_13964,N_13631);
xnor U14468 (N_14468,N_13607,N_13909);
or U14469 (N_14469,N_13900,N_13755);
or U14470 (N_14470,N_14000,N_13996);
and U14471 (N_14471,N_14108,N_14064);
and U14472 (N_14472,N_13829,N_13720);
or U14473 (N_14473,N_13749,N_14127);
and U14474 (N_14474,N_14120,N_13884);
or U14475 (N_14475,N_13812,N_13762);
nor U14476 (N_14476,N_13940,N_13509);
and U14477 (N_14477,N_13732,N_13717);
and U14478 (N_14478,N_14173,N_13956);
or U14479 (N_14479,N_13542,N_13907);
nor U14480 (N_14480,N_14112,N_13878);
nand U14481 (N_14481,N_14057,N_13843);
nor U14482 (N_14482,N_14240,N_14177);
and U14483 (N_14483,N_13557,N_13543);
or U14484 (N_14484,N_14020,N_14051);
or U14485 (N_14485,N_13903,N_14180);
and U14486 (N_14486,N_14122,N_14040);
and U14487 (N_14487,N_13502,N_14114);
nand U14488 (N_14488,N_13645,N_13770);
nand U14489 (N_14489,N_14216,N_14090);
xor U14490 (N_14490,N_14054,N_14195);
or U14491 (N_14491,N_14182,N_13505);
nor U14492 (N_14492,N_13958,N_13855);
nor U14493 (N_14493,N_13945,N_14011);
or U14494 (N_14494,N_14098,N_14085);
and U14495 (N_14495,N_14174,N_13724);
or U14496 (N_14496,N_13630,N_13933);
or U14497 (N_14497,N_13680,N_13669);
or U14498 (N_14498,N_13729,N_14224);
nor U14499 (N_14499,N_13721,N_13530);
or U14500 (N_14500,N_13636,N_14125);
or U14501 (N_14501,N_13823,N_13892);
and U14502 (N_14502,N_14151,N_13980);
or U14503 (N_14503,N_13604,N_14201);
or U14504 (N_14504,N_14059,N_14145);
or U14505 (N_14505,N_13618,N_13751);
and U14506 (N_14506,N_13833,N_14060);
nor U14507 (N_14507,N_13874,N_14167);
nor U14508 (N_14508,N_14137,N_14015);
or U14509 (N_14509,N_13943,N_13756);
or U14510 (N_14510,N_14249,N_14115);
nand U14511 (N_14511,N_13802,N_13976);
and U14512 (N_14512,N_14094,N_13830);
nor U14513 (N_14513,N_13694,N_13657);
and U14514 (N_14514,N_13563,N_13522);
or U14515 (N_14515,N_13924,N_13643);
or U14516 (N_14516,N_14134,N_14170);
nor U14517 (N_14517,N_13877,N_14150);
nand U14518 (N_14518,N_13894,N_14144);
nor U14519 (N_14519,N_13610,N_13616);
nand U14520 (N_14520,N_13828,N_14012);
nand U14521 (N_14521,N_13979,N_14213);
nor U14522 (N_14522,N_14159,N_13660);
or U14523 (N_14523,N_14181,N_13689);
nor U14524 (N_14524,N_13524,N_13605);
nor U14525 (N_14525,N_13941,N_13807);
xor U14526 (N_14526,N_13901,N_13784);
and U14527 (N_14527,N_13906,N_14210);
and U14528 (N_14528,N_13519,N_13545);
or U14529 (N_14529,N_13513,N_13640);
or U14530 (N_14530,N_13973,N_13995);
and U14531 (N_14531,N_14158,N_13786);
xnor U14532 (N_14532,N_14190,N_13991);
nor U14533 (N_14533,N_14102,N_14209);
nand U14534 (N_14534,N_14168,N_14155);
and U14535 (N_14535,N_13971,N_13710);
and U14536 (N_14536,N_14044,N_13902);
or U14537 (N_14537,N_13683,N_13795);
or U14538 (N_14538,N_14022,N_13593);
xor U14539 (N_14539,N_13594,N_13713);
and U14540 (N_14540,N_13789,N_13537);
or U14541 (N_14541,N_13950,N_14139);
xnor U14542 (N_14542,N_14023,N_14028);
or U14543 (N_14543,N_13525,N_13528);
and U14544 (N_14544,N_13641,N_13742);
and U14545 (N_14545,N_13654,N_13951);
nor U14546 (N_14546,N_13791,N_13707);
or U14547 (N_14547,N_13864,N_13842);
and U14548 (N_14548,N_14147,N_14204);
xor U14549 (N_14549,N_13827,N_13527);
and U14550 (N_14550,N_14142,N_13820);
or U14551 (N_14551,N_14038,N_14113);
nor U14552 (N_14552,N_13558,N_13866);
and U14553 (N_14553,N_13803,N_14116);
nand U14554 (N_14554,N_13931,N_13539);
xnor U14555 (N_14555,N_14084,N_13785);
and U14556 (N_14556,N_13590,N_13576);
and U14557 (N_14557,N_14111,N_13895);
and U14558 (N_14558,N_13942,N_13916);
and U14559 (N_14559,N_13952,N_14164);
or U14560 (N_14560,N_14199,N_13659);
xnor U14561 (N_14561,N_14048,N_13818);
nor U14562 (N_14562,N_13699,N_14166);
or U14563 (N_14563,N_13875,N_13671);
or U14564 (N_14564,N_13926,N_13561);
nor U14565 (N_14565,N_13824,N_13862);
or U14566 (N_14566,N_14244,N_13927);
or U14567 (N_14567,N_14140,N_13677);
or U14568 (N_14568,N_13608,N_13859);
nand U14569 (N_14569,N_13752,N_14143);
nand U14570 (N_14570,N_14025,N_13638);
and U14571 (N_14571,N_14006,N_13728);
or U14572 (N_14572,N_13930,N_13646);
or U14573 (N_14573,N_13714,N_13609);
nand U14574 (N_14574,N_14095,N_13934);
and U14575 (N_14575,N_13637,N_13748);
nor U14576 (N_14576,N_13796,N_14093);
nor U14577 (N_14577,N_13955,N_13938);
or U14578 (N_14578,N_14234,N_13744);
or U14579 (N_14579,N_13670,N_14070);
nand U14580 (N_14580,N_14109,N_13999);
xor U14581 (N_14581,N_14192,N_14019);
and U14582 (N_14582,N_14236,N_14055);
and U14583 (N_14583,N_13658,N_14148);
nand U14584 (N_14584,N_13838,N_13914);
or U14585 (N_14585,N_13591,N_13788);
nand U14586 (N_14586,N_13775,N_14083);
or U14587 (N_14587,N_14205,N_13743);
or U14588 (N_14588,N_13937,N_13531);
nor U14589 (N_14589,N_13858,N_13635);
or U14590 (N_14590,N_13647,N_13679);
nor U14591 (N_14591,N_14074,N_13867);
xnor U14592 (N_14592,N_13780,N_13825);
nand U14593 (N_14593,N_13541,N_13731);
nor U14594 (N_14594,N_14188,N_13992);
and U14595 (N_14595,N_13811,N_13507);
and U14596 (N_14596,N_13625,N_13653);
nor U14597 (N_14597,N_13873,N_13889);
nor U14598 (N_14598,N_13692,N_13787);
nor U14599 (N_14599,N_13870,N_14078);
nor U14600 (N_14600,N_13702,N_13526);
xnor U14601 (N_14601,N_14243,N_14092);
nor U14602 (N_14602,N_14154,N_13793);
and U14603 (N_14603,N_14042,N_14037);
or U14604 (N_14604,N_14156,N_14146);
nand U14605 (N_14605,N_13984,N_13760);
nor U14606 (N_14606,N_14035,N_13804);
and U14607 (N_14607,N_14223,N_13716);
and U14608 (N_14608,N_13868,N_14101);
nor U14609 (N_14609,N_13555,N_14056);
nand U14610 (N_14610,N_13928,N_14128);
nand U14611 (N_14611,N_13703,N_13982);
nor U14612 (N_14612,N_13886,N_14005);
and U14613 (N_14613,N_13723,N_13726);
nor U14614 (N_14614,N_13840,N_14133);
or U14615 (N_14615,N_13853,N_14176);
nand U14616 (N_14616,N_13773,N_13668);
nand U14617 (N_14617,N_13705,N_14030);
nand U14618 (N_14618,N_13719,N_13516);
nand U14619 (N_14619,N_14021,N_13871);
nand U14620 (N_14620,N_14100,N_13879);
xor U14621 (N_14621,N_13556,N_13861);
or U14622 (N_14622,N_14242,N_13585);
nor U14623 (N_14623,N_13617,N_13766);
or U14624 (N_14624,N_13848,N_14080);
and U14625 (N_14625,N_14016,N_14104);
or U14626 (N_14626,N_14190,N_13571);
nor U14627 (N_14627,N_13580,N_13538);
nor U14628 (N_14628,N_13687,N_13745);
or U14629 (N_14629,N_14045,N_13831);
nor U14630 (N_14630,N_13716,N_14225);
or U14631 (N_14631,N_13846,N_13948);
or U14632 (N_14632,N_14146,N_14126);
nand U14633 (N_14633,N_14235,N_14204);
or U14634 (N_14634,N_14121,N_13852);
or U14635 (N_14635,N_13908,N_13779);
and U14636 (N_14636,N_14109,N_13943);
nand U14637 (N_14637,N_13683,N_13776);
and U14638 (N_14638,N_13693,N_14053);
nand U14639 (N_14639,N_13742,N_14107);
or U14640 (N_14640,N_13755,N_13517);
nand U14641 (N_14641,N_13654,N_14151);
and U14642 (N_14642,N_13643,N_14180);
nand U14643 (N_14643,N_14030,N_13628);
nand U14644 (N_14644,N_13995,N_14152);
nand U14645 (N_14645,N_13745,N_13970);
or U14646 (N_14646,N_13579,N_13766);
xor U14647 (N_14647,N_14169,N_14066);
and U14648 (N_14648,N_13500,N_14020);
nand U14649 (N_14649,N_14195,N_14023);
nor U14650 (N_14650,N_13906,N_13543);
or U14651 (N_14651,N_14081,N_14239);
nand U14652 (N_14652,N_13792,N_13993);
nand U14653 (N_14653,N_14073,N_13574);
nor U14654 (N_14654,N_13838,N_14043);
or U14655 (N_14655,N_13788,N_14208);
and U14656 (N_14656,N_13662,N_14211);
nand U14657 (N_14657,N_13985,N_13738);
and U14658 (N_14658,N_13692,N_13728);
nand U14659 (N_14659,N_13672,N_14041);
and U14660 (N_14660,N_13857,N_14067);
nand U14661 (N_14661,N_13542,N_14026);
nor U14662 (N_14662,N_13551,N_13837);
or U14663 (N_14663,N_13813,N_13858);
nor U14664 (N_14664,N_13963,N_14029);
xor U14665 (N_14665,N_13787,N_14179);
nand U14666 (N_14666,N_13705,N_13528);
nand U14667 (N_14667,N_13800,N_13991);
nand U14668 (N_14668,N_13624,N_14080);
nand U14669 (N_14669,N_13944,N_13922);
or U14670 (N_14670,N_13540,N_13717);
or U14671 (N_14671,N_14086,N_14172);
nor U14672 (N_14672,N_13743,N_14091);
nor U14673 (N_14673,N_13689,N_13837);
nor U14674 (N_14674,N_13566,N_14056);
xnor U14675 (N_14675,N_13519,N_14234);
or U14676 (N_14676,N_13825,N_14023);
nand U14677 (N_14677,N_14054,N_13799);
nand U14678 (N_14678,N_14020,N_13990);
nand U14679 (N_14679,N_13664,N_14226);
nor U14680 (N_14680,N_14124,N_13561);
and U14681 (N_14681,N_14215,N_13537);
xnor U14682 (N_14682,N_13816,N_13687);
nor U14683 (N_14683,N_14011,N_13958);
and U14684 (N_14684,N_13868,N_14227);
nor U14685 (N_14685,N_13874,N_13976);
and U14686 (N_14686,N_13846,N_14024);
and U14687 (N_14687,N_13672,N_13859);
nand U14688 (N_14688,N_13878,N_13678);
nand U14689 (N_14689,N_13832,N_13937);
and U14690 (N_14690,N_13910,N_13778);
or U14691 (N_14691,N_13821,N_14067);
nand U14692 (N_14692,N_14093,N_13537);
nand U14693 (N_14693,N_14032,N_14223);
or U14694 (N_14694,N_13784,N_14069);
xnor U14695 (N_14695,N_13506,N_14168);
nand U14696 (N_14696,N_14184,N_14116);
nor U14697 (N_14697,N_13660,N_14083);
xor U14698 (N_14698,N_13901,N_13961);
nand U14699 (N_14699,N_13895,N_14050);
nand U14700 (N_14700,N_14198,N_13740);
or U14701 (N_14701,N_13799,N_13810);
xor U14702 (N_14702,N_13939,N_14068);
and U14703 (N_14703,N_13700,N_14001);
nand U14704 (N_14704,N_13728,N_13511);
nand U14705 (N_14705,N_13752,N_13509);
xnor U14706 (N_14706,N_13991,N_13849);
nor U14707 (N_14707,N_13976,N_13769);
nand U14708 (N_14708,N_13937,N_13548);
xnor U14709 (N_14709,N_14097,N_13809);
nand U14710 (N_14710,N_13865,N_13823);
nor U14711 (N_14711,N_13662,N_13587);
and U14712 (N_14712,N_13902,N_13725);
and U14713 (N_14713,N_14027,N_13801);
and U14714 (N_14714,N_13852,N_14011);
or U14715 (N_14715,N_13628,N_13662);
nand U14716 (N_14716,N_14090,N_14183);
xor U14717 (N_14717,N_13751,N_13962);
nor U14718 (N_14718,N_14210,N_13699);
and U14719 (N_14719,N_13824,N_14013);
and U14720 (N_14720,N_14066,N_13704);
xnor U14721 (N_14721,N_13835,N_13972);
and U14722 (N_14722,N_13964,N_14054);
nand U14723 (N_14723,N_14200,N_13755);
or U14724 (N_14724,N_13958,N_13552);
and U14725 (N_14725,N_14034,N_13634);
nor U14726 (N_14726,N_14246,N_14015);
xor U14727 (N_14727,N_13942,N_14133);
and U14728 (N_14728,N_13992,N_14245);
and U14729 (N_14729,N_14165,N_13777);
nor U14730 (N_14730,N_13851,N_13787);
and U14731 (N_14731,N_13978,N_13670);
or U14732 (N_14732,N_13934,N_13515);
or U14733 (N_14733,N_13803,N_13845);
nand U14734 (N_14734,N_13990,N_14093);
nand U14735 (N_14735,N_13772,N_13582);
and U14736 (N_14736,N_13561,N_13659);
and U14737 (N_14737,N_13762,N_13581);
and U14738 (N_14738,N_14122,N_13526);
xnor U14739 (N_14739,N_13717,N_14212);
nor U14740 (N_14740,N_13631,N_13526);
and U14741 (N_14741,N_13544,N_14051);
xor U14742 (N_14742,N_13515,N_13645);
or U14743 (N_14743,N_14033,N_13989);
nand U14744 (N_14744,N_13886,N_13847);
nand U14745 (N_14745,N_14228,N_13723);
xnor U14746 (N_14746,N_13622,N_13808);
and U14747 (N_14747,N_13926,N_14224);
nand U14748 (N_14748,N_14236,N_14104);
and U14749 (N_14749,N_13620,N_13553);
or U14750 (N_14750,N_13749,N_13618);
xor U14751 (N_14751,N_13710,N_14247);
or U14752 (N_14752,N_14141,N_14006);
or U14753 (N_14753,N_13855,N_14213);
xnor U14754 (N_14754,N_13810,N_14123);
nand U14755 (N_14755,N_14012,N_13663);
nand U14756 (N_14756,N_14234,N_14113);
or U14757 (N_14757,N_14106,N_13902);
or U14758 (N_14758,N_13720,N_13825);
or U14759 (N_14759,N_14023,N_14225);
nor U14760 (N_14760,N_14156,N_13985);
and U14761 (N_14761,N_14002,N_14109);
nand U14762 (N_14762,N_13777,N_13686);
nor U14763 (N_14763,N_13577,N_13889);
nor U14764 (N_14764,N_13748,N_13714);
or U14765 (N_14765,N_13633,N_14176);
nor U14766 (N_14766,N_14216,N_13793);
nand U14767 (N_14767,N_13620,N_13967);
or U14768 (N_14768,N_13574,N_14017);
or U14769 (N_14769,N_13669,N_14187);
and U14770 (N_14770,N_14123,N_13963);
nor U14771 (N_14771,N_14147,N_14084);
nor U14772 (N_14772,N_13842,N_13894);
and U14773 (N_14773,N_14004,N_14066);
nand U14774 (N_14774,N_14138,N_14016);
or U14775 (N_14775,N_14099,N_14180);
nor U14776 (N_14776,N_14194,N_13753);
nor U14777 (N_14777,N_14094,N_14081);
nand U14778 (N_14778,N_13515,N_14085);
and U14779 (N_14779,N_13925,N_13664);
and U14780 (N_14780,N_13769,N_13992);
nand U14781 (N_14781,N_13725,N_14210);
nand U14782 (N_14782,N_14065,N_13767);
nor U14783 (N_14783,N_13924,N_13610);
nand U14784 (N_14784,N_13556,N_14092);
nor U14785 (N_14785,N_13870,N_13700);
xor U14786 (N_14786,N_13653,N_13935);
or U14787 (N_14787,N_14176,N_13963);
nand U14788 (N_14788,N_14180,N_13876);
or U14789 (N_14789,N_13695,N_13816);
and U14790 (N_14790,N_13922,N_14180);
nand U14791 (N_14791,N_13518,N_13513);
nor U14792 (N_14792,N_13768,N_14119);
and U14793 (N_14793,N_13899,N_13796);
and U14794 (N_14794,N_14034,N_13557);
nand U14795 (N_14795,N_14022,N_13879);
and U14796 (N_14796,N_14182,N_13569);
nand U14797 (N_14797,N_14152,N_13700);
nand U14798 (N_14798,N_13564,N_13747);
nand U14799 (N_14799,N_14211,N_13740);
or U14800 (N_14800,N_13831,N_14013);
xnor U14801 (N_14801,N_13794,N_14055);
or U14802 (N_14802,N_13897,N_13752);
xor U14803 (N_14803,N_14232,N_13631);
or U14804 (N_14804,N_13840,N_13793);
and U14805 (N_14805,N_13850,N_13688);
nor U14806 (N_14806,N_13881,N_13631);
or U14807 (N_14807,N_13955,N_13816);
and U14808 (N_14808,N_13541,N_13755);
nor U14809 (N_14809,N_13865,N_13803);
and U14810 (N_14810,N_13906,N_14042);
or U14811 (N_14811,N_14016,N_14046);
xor U14812 (N_14812,N_13525,N_13833);
or U14813 (N_14813,N_13596,N_14159);
and U14814 (N_14814,N_14039,N_14228);
nand U14815 (N_14815,N_14223,N_14079);
or U14816 (N_14816,N_13869,N_13531);
or U14817 (N_14817,N_13970,N_13536);
nand U14818 (N_14818,N_14128,N_13697);
and U14819 (N_14819,N_14094,N_13683);
and U14820 (N_14820,N_14235,N_14148);
nor U14821 (N_14821,N_14238,N_14178);
nor U14822 (N_14822,N_13577,N_13959);
or U14823 (N_14823,N_13711,N_13680);
xnor U14824 (N_14824,N_13813,N_13908);
nor U14825 (N_14825,N_14114,N_13878);
nand U14826 (N_14826,N_13509,N_14159);
nor U14827 (N_14827,N_13615,N_13791);
nand U14828 (N_14828,N_14195,N_13736);
or U14829 (N_14829,N_13553,N_14109);
nor U14830 (N_14830,N_14213,N_14229);
and U14831 (N_14831,N_13801,N_13685);
nor U14832 (N_14832,N_13598,N_13962);
nand U14833 (N_14833,N_13731,N_13682);
nor U14834 (N_14834,N_13859,N_13804);
or U14835 (N_14835,N_13904,N_13586);
xor U14836 (N_14836,N_13695,N_14164);
and U14837 (N_14837,N_13692,N_14082);
or U14838 (N_14838,N_14187,N_13681);
nor U14839 (N_14839,N_13921,N_13976);
xor U14840 (N_14840,N_13914,N_13548);
or U14841 (N_14841,N_13592,N_13572);
or U14842 (N_14842,N_14022,N_14074);
and U14843 (N_14843,N_14083,N_14097);
nand U14844 (N_14844,N_13644,N_13806);
nand U14845 (N_14845,N_13875,N_13777);
nor U14846 (N_14846,N_13715,N_13615);
xor U14847 (N_14847,N_14048,N_14098);
xnor U14848 (N_14848,N_13955,N_13616);
nor U14849 (N_14849,N_13528,N_13891);
nor U14850 (N_14850,N_13857,N_13611);
nor U14851 (N_14851,N_13745,N_13903);
xor U14852 (N_14852,N_14058,N_13539);
xor U14853 (N_14853,N_13544,N_14215);
xor U14854 (N_14854,N_14054,N_14227);
nor U14855 (N_14855,N_14133,N_14149);
or U14856 (N_14856,N_13887,N_14044);
and U14857 (N_14857,N_13592,N_13602);
nor U14858 (N_14858,N_14166,N_14095);
nor U14859 (N_14859,N_13807,N_13594);
and U14860 (N_14860,N_13988,N_13763);
nor U14861 (N_14861,N_13620,N_14222);
nand U14862 (N_14862,N_13999,N_13803);
xnor U14863 (N_14863,N_13856,N_13967);
nand U14864 (N_14864,N_13910,N_13636);
or U14865 (N_14865,N_14116,N_13732);
nor U14866 (N_14866,N_13902,N_14218);
nand U14867 (N_14867,N_13647,N_14219);
nor U14868 (N_14868,N_13679,N_13681);
xor U14869 (N_14869,N_13864,N_13936);
nor U14870 (N_14870,N_14173,N_13510);
and U14871 (N_14871,N_13799,N_13664);
nand U14872 (N_14872,N_13815,N_14111);
or U14873 (N_14873,N_13761,N_13628);
or U14874 (N_14874,N_13944,N_13961);
nor U14875 (N_14875,N_13698,N_13561);
nor U14876 (N_14876,N_14113,N_13937);
and U14877 (N_14877,N_14165,N_14059);
nand U14878 (N_14878,N_13589,N_14176);
nor U14879 (N_14879,N_14143,N_14154);
or U14880 (N_14880,N_14002,N_14162);
xnor U14881 (N_14881,N_13661,N_13856);
nand U14882 (N_14882,N_14213,N_13623);
nor U14883 (N_14883,N_13787,N_13601);
nand U14884 (N_14884,N_14142,N_13765);
and U14885 (N_14885,N_14105,N_13651);
xnor U14886 (N_14886,N_14011,N_13821);
xor U14887 (N_14887,N_13890,N_13981);
or U14888 (N_14888,N_13569,N_13716);
xnor U14889 (N_14889,N_13866,N_14235);
and U14890 (N_14890,N_14074,N_13894);
nand U14891 (N_14891,N_13613,N_13668);
nor U14892 (N_14892,N_13872,N_13669);
or U14893 (N_14893,N_13909,N_13531);
or U14894 (N_14894,N_14163,N_13952);
or U14895 (N_14895,N_14158,N_14052);
xnor U14896 (N_14896,N_13899,N_14072);
xor U14897 (N_14897,N_13832,N_13813);
nor U14898 (N_14898,N_14183,N_13671);
and U14899 (N_14899,N_13974,N_14037);
nand U14900 (N_14900,N_14082,N_14078);
nor U14901 (N_14901,N_14016,N_14080);
or U14902 (N_14902,N_13988,N_14144);
nand U14903 (N_14903,N_14186,N_13717);
or U14904 (N_14904,N_13817,N_13827);
and U14905 (N_14905,N_14026,N_13614);
or U14906 (N_14906,N_13887,N_14022);
or U14907 (N_14907,N_13584,N_13630);
nand U14908 (N_14908,N_14049,N_14084);
or U14909 (N_14909,N_13736,N_14157);
or U14910 (N_14910,N_13643,N_13806);
nor U14911 (N_14911,N_13830,N_13597);
or U14912 (N_14912,N_14145,N_13611);
or U14913 (N_14913,N_13535,N_13762);
and U14914 (N_14914,N_13664,N_13849);
nand U14915 (N_14915,N_14124,N_13732);
nor U14916 (N_14916,N_13970,N_13792);
xnor U14917 (N_14917,N_14115,N_13793);
and U14918 (N_14918,N_13987,N_13888);
nand U14919 (N_14919,N_13794,N_14070);
and U14920 (N_14920,N_13851,N_13714);
and U14921 (N_14921,N_13777,N_13641);
nor U14922 (N_14922,N_14223,N_14121);
and U14923 (N_14923,N_13823,N_13759);
or U14924 (N_14924,N_13871,N_13763);
nand U14925 (N_14925,N_14222,N_14054);
nand U14926 (N_14926,N_13970,N_13722);
or U14927 (N_14927,N_13824,N_13715);
nand U14928 (N_14928,N_13779,N_13599);
or U14929 (N_14929,N_13541,N_13551);
and U14930 (N_14930,N_13614,N_13915);
nor U14931 (N_14931,N_14196,N_13941);
or U14932 (N_14932,N_13698,N_13526);
nand U14933 (N_14933,N_13796,N_14194);
nand U14934 (N_14934,N_13512,N_13949);
and U14935 (N_14935,N_13790,N_13995);
and U14936 (N_14936,N_14030,N_13756);
or U14937 (N_14937,N_13744,N_14091);
nor U14938 (N_14938,N_14138,N_14050);
nand U14939 (N_14939,N_14184,N_13565);
and U14940 (N_14940,N_13566,N_13977);
xor U14941 (N_14941,N_13561,N_14017);
nor U14942 (N_14942,N_14164,N_13604);
or U14943 (N_14943,N_13893,N_13748);
nor U14944 (N_14944,N_14239,N_13607);
nor U14945 (N_14945,N_13901,N_13791);
and U14946 (N_14946,N_13808,N_14074);
nand U14947 (N_14947,N_13526,N_13996);
xor U14948 (N_14948,N_13572,N_14202);
nand U14949 (N_14949,N_13740,N_13659);
nor U14950 (N_14950,N_14228,N_13613);
nand U14951 (N_14951,N_13892,N_14076);
nor U14952 (N_14952,N_13615,N_14214);
or U14953 (N_14953,N_13631,N_13993);
or U14954 (N_14954,N_14122,N_14233);
and U14955 (N_14955,N_13517,N_13962);
xnor U14956 (N_14956,N_14086,N_14239);
nor U14957 (N_14957,N_14190,N_13508);
and U14958 (N_14958,N_14101,N_13984);
nor U14959 (N_14959,N_14029,N_13698);
or U14960 (N_14960,N_14070,N_13555);
and U14961 (N_14961,N_14219,N_13906);
or U14962 (N_14962,N_13516,N_14124);
xnor U14963 (N_14963,N_13769,N_14230);
nand U14964 (N_14964,N_13556,N_14044);
and U14965 (N_14965,N_13899,N_14189);
nor U14966 (N_14966,N_14185,N_14101);
nor U14967 (N_14967,N_13703,N_13679);
or U14968 (N_14968,N_13737,N_13995);
nand U14969 (N_14969,N_13866,N_14167);
nor U14970 (N_14970,N_13976,N_13502);
and U14971 (N_14971,N_13613,N_13510);
or U14972 (N_14972,N_14119,N_13935);
or U14973 (N_14973,N_14227,N_13711);
nor U14974 (N_14974,N_14173,N_13919);
and U14975 (N_14975,N_13973,N_14232);
nand U14976 (N_14976,N_13996,N_13990);
xor U14977 (N_14977,N_13664,N_13700);
nor U14978 (N_14978,N_14245,N_13522);
xnor U14979 (N_14979,N_13854,N_13998);
and U14980 (N_14980,N_14164,N_13949);
or U14981 (N_14981,N_13578,N_14169);
nand U14982 (N_14982,N_14113,N_13951);
or U14983 (N_14983,N_14052,N_14200);
nand U14984 (N_14984,N_13757,N_13774);
or U14985 (N_14985,N_13870,N_13986);
nand U14986 (N_14986,N_14055,N_13769);
xor U14987 (N_14987,N_13932,N_13579);
nand U14988 (N_14988,N_14086,N_14249);
nand U14989 (N_14989,N_14240,N_13625);
nor U14990 (N_14990,N_13542,N_13853);
and U14991 (N_14991,N_13857,N_13902);
xor U14992 (N_14992,N_13753,N_14099);
nand U14993 (N_14993,N_13696,N_14057);
nand U14994 (N_14994,N_13739,N_14147);
nand U14995 (N_14995,N_14122,N_13946);
nand U14996 (N_14996,N_13648,N_13960);
nor U14997 (N_14997,N_14067,N_13523);
and U14998 (N_14998,N_13616,N_14234);
or U14999 (N_14999,N_14168,N_14088);
nor UO_0 (O_0,N_14545,N_14819);
nor UO_1 (O_1,N_14530,N_14678);
or UO_2 (O_2,N_14750,N_14301);
nand UO_3 (O_3,N_14659,N_14486);
nand UO_4 (O_4,N_14492,N_14499);
and UO_5 (O_5,N_14980,N_14946);
xor UO_6 (O_6,N_14693,N_14336);
nand UO_7 (O_7,N_14978,N_14908);
nand UO_8 (O_8,N_14307,N_14781);
or UO_9 (O_9,N_14446,N_14661);
nand UO_10 (O_10,N_14809,N_14812);
nand UO_11 (O_11,N_14982,N_14601);
and UO_12 (O_12,N_14565,N_14599);
or UO_13 (O_13,N_14363,N_14835);
and UO_14 (O_14,N_14947,N_14421);
or UO_15 (O_15,N_14483,N_14293);
or UO_16 (O_16,N_14430,N_14490);
or UO_17 (O_17,N_14801,N_14451);
or UO_18 (O_18,N_14616,N_14692);
and UO_19 (O_19,N_14620,N_14452);
or UO_20 (O_20,N_14785,N_14264);
or UO_21 (O_21,N_14808,N_14869);
nand UO_22 (O_22,N_14383,N_14425);
nand UO_23 (O_23,N_14881,N_14780);
nor UO_24 (O_24,N_14584,N_14871);
nand UO_25 (O_25,N_14256,N_14755);
xor UO_26 (O_26,N_14969,N_14501);
nor UO_27 (O_27,N_14830,N_14314);
nand UO_28 (O_28,N_14368,N_14393);
xor UO_29 (O_29,N_14807,N_14289);
nand UO_30 (O_30,N_14358,N_14909);
nor UO_31 (O_31,N_14444,N_14502);
nor UO_32 (O_32,N_14382,N_14720);
or UO_33 (O_33,N_14511,N_14274);
or UO_34 (O_34,N_14943,N_14321);
xor UO_35 (O_35,N_14811,N_14743);
nand UO_36 (O_36,N_14291,N_14742);
nor UO_37 (O_37,N_14284,N_14267);
or UO_38 (O_38,N_14974,N_14656);
and UO_39 (O_39,N_14298,N_14261);
nor UO_40 (O_40,N_14642,N_14255);
nor UO_41 (O_41,N_14457,N_14603);
nand UO_42 (O_42,N_14259,N_14863);
and UO_43 (O_43,N_14715,N_14318);
xor UO_44 (O_44,N_14919,N_14448);
or UO_45 (O_45,N_14398,N_14397);
nand UO_46 (O_46,N_14939,N_14664);
nor UO_47 (O_47,N_14543,N_14898);
and UO_48 (O_48,N_14837,N_14832);
nor UO_49 (O_49,N_14381,N_14370);
nand UO_50 (O_50,N_14766,N_14254);
nand UO_51 (O_51,N_14561,N_14300);
nor UO_52 (O_52,N_14675,N_14280);
or UO_53 (O_53,N_14331,N_14450);
nand UO_54 (O_54,N_14705,N_14774);
nand UO_55 (O_55,N_14414,N_14756);
nand UO_56 (O_56,N_14663,N_14641);
nand UO_57 (O_57,N_14416,N_14672);
and UO_58 (O_58,N_14602,N_14341);
nor UO_59 (O_59,N_14698,N_14953);
nor UO_60 (O_60,N_14771,N_14462);
nor UO_61 (O_61,N_14480,N_14296);
nor UO_62 (O_62,N_14660,N_14708);
or UO_63 (O_63,N_14328,N_14729);
and UO_64 (O_64,N_14555,N_14359);
nand UO_65 (O_65,N_14690,N_14573);
xnor UO_66 (O_66,N_14657,N_14569);
or UO_67 (O_67,N_14349,N_14442);
xor UO_68 (O_68,N_14332,N_14695);
nand UO_69 (O_69,N_14864,N_14907);
and UO_70 (O_70,N_14391,N_14784);
nor UO_71 (O_71,N_14670,N_14831);
and UO_72 (O_72,N_14822,N_14882);
nand UO_73 (O_73,N_14913,N_14803);
xnor UO_74 (O_74,N_14282,N_14445);
nor UO_75 (O_75,N_14709,N_14515);
or UO_76 (O_76,N_14921,N_14631);
nand UO_77 (O_77,N_14392,N_14551);
nand UO_78 (O_78,N_14966,N_14400);
and UO_79 (O_79,N_14302,N_14773);
nand UO_80 (O_80,N_14987,N_14879);
and UO_81 (O_81,N_14748,N_14873);
xnor UO_82 (O_82,N_14554,N_14717);
nor UO_83 (O_83,N_14345,N_14304);
nand UO_84 (O_84,N_14783,N_14677);
and UO_85 (O_85,N_14776,N_14329);
nor UO_86 (O_86,N_14266,N_14374);
nand UO_87 (O_87,N_14814,N_14993);
and UO_88 (O_88,N_14932,N_14582);
nand UO_89 (O_89,N_14853,N_14440);
and UO_90 (O_90,N_14997,N_14722);
or UO_91 (O_91,N_14481,N_14648);
or UO_92 (O_92,N_14322,N_14817);
nand UO_93 (O_93,N_14523,N_14458);
nand UO_94 (O_94,N_14860,N_14733);
nand UO_95 (O_95,N_14734,N_14253);
nor UO_96 (O_96,N_14567,N_14961);
nand UO_97 (O_97,N_14892,N_14310);
and UO_98 (O_98,N_14439,N_14948);
nor UO_99 (O_99,N_14357,N_14745);
nand UO_100 (O_100,N_14962,N_14806);
nand UO_101 (O_101,N_14360,N_14920);
xor UO_102 (O_102,N_14754,N_14372);
and UO_103 (O_103,N_14638,N_14721);
nand UO_104 (O_104,N_14403,N_14759);
nand UO_105 (O_105,N_14257,N_14852);
nor UO_106 (O_106,N_14612,N_14277);
nor UO_107 (O_107,N_14687,N_14682);
xnor UO_108 (O_108,N_14688,N_14799);
nand UO_109 (O_109,N_14662,N_14900);
xor UO_110 (O_110,N_14885,N_14354);
or UO_111 (O_111,N_14593,N_14968);
nand UO_112 (O_112,N_14598,N_14384);
nor UO_113 (O_113,N_14741,N_14681);
nor UO_114 (O_114,N_14294,N_14668);
nand UO_115 (O_115,N_14834,N_14376);
or UO_116 (O_116,N_14471,N_14855);
nand UO_117 (O_117,N_14726,N_14958);
nand UO_118 (O_118,N_14699,N_14487);
or UO_119 (O_119,N_14265,N_14517);
nand UO_120 (O_120,N_14614,N_14923);
or UO_121 (O_121,N_14607,N_14676);
xnor UO_122 (O_122,N_14258,N_14408);
nand UO_123 (O_123,N_14506,N_14926);
nand UO_124 (O_124,N_14903,N_14433);
xnor UO_125 (O_125,N_14821,N_14883);
nor UO_126 (O_126,N_14604,N_14977);
nor UO_127 (O_127,N_14348,N_14438);
or UO_128 (O_128,N_14609,N_14320);
nor UO_129 (O_129,N_14521,N_14972);
nor UO_130 (O_130,N_14531,N_14586);
and UO_131 (O_131,N_14417,N_14665);
nand UO_132 (O_132,N_14933,N_14880);
xnor UO_133 (O_133,N_14537,N_14610);
xnor UO_134 (O_134,N_14299,N_14477);
and UO_135 (O_135,N_14611,N_14538);
or UO_136 (O_136,N_14469,N_14658);
or UO_137 (O_137,N_14976,N_14454);
nand UO_138 (O_138,N_14824,N_14333);
xnor UO_139 (O_139,N_14666,N_14279);
nand UO_140 (O_140,N_14934,N_14394);
or UO_141 (O_141,N_14632,N_14262);
xor UO_142 (O_142,N_14833,N_14644);
xnor UO_143 (O_143,N_14495,N_14423);
xor UO_144 (O_144,N_14574,N_14366);
and UO_145 (O_145,N_14390,N_14325);
and UO_146 (O_146,N_14347,N_14870);
nor UO_147 (O_147,N_14878,N_14588);
nor UO_148 (O_148,N_14906,N_14550);
and UO_149 (O_149,N_14330,N_14557);
or UO_150 (O_150,N_14412,N_14522);
nand UO_151 (O_151,N_14981,N_14410);
xor UO_152 (O_152,N_14500,N_14411);
nor UO_153 (O_153,N_14305,N_14983);
xor UO_154 (O_154,N_14753,N_14991);
and UO_155 (O_155,N_14749,N_14367);
or UO_156 (O_156,N_14624,N_14804);
nand UO_157 (O_157,N_14769,N_14988);
and UO_158 (O_158,N_14912,N_14914);
or UO_159 (O_159,N_14449,N_14590);
xor UO_160 (O_160,N_14649,N_14790);
or UO_161 (O_161,N_14514,N_14570);
nand UO_162 (O_162,N_14866,N_14889);
nor UO_163 (O_163,N_14459,N_14704);
or UO_164 (O_164,N_14475,N_14396);
nand UO_165 (O_165,N_14546,N_14399);
nor UO_166 (O_166,N_14989,N_14536);
or UO_167 (O_167,N_14793,N_14655);
and UO_168 (O_168,N_14512,N_14850);
and UO_169 (O_169,N_14539,N_14472);
nand UO_170 (O_170,N_14434,N_14952);
nand UO_171 (O_171,N_14549,N_14591);
nor UO_172 (O_172,N_14973,N_14994);
or UO_173 (O_173,N_14736,N_14760);
and UO_174 (O_174,N_14957,N_14849);
or UO_175 (O_175,N_14904,N_14971);
nor UO_176 (O_176,N_14409,N_14292);
nand UO_177 (O_177,N_14303,N_14875);
and UO_178 (O_178,N_14455,N_14918);
nor UO_179 (O_179,N_14419,N_14563);
nor UO_180 (O_180,N_14541,N_14437);
and UO_181 (O_181,N_14826,N_14847);
nor UO_182 (O_182,N_14975,N_14746);
or UO_183 (O_183,N_14465,N_14606);
nor UO_184 (O_184,N_14772,N_14429);
nor UO_185 (O_185,N_14626,N_14813);
nand UO_186 (O_186,N_14380,N_14556);
nand UO_187 (O_187,N_14577,N_14851);
nor UO_188 (O_188,N_14694,N_14525);
and UO_189 (O_189,N_14542,N_14615);
xnor UO_190 (O_190,N_14273,N_14323);
or UO_191 (O_191,N_14911,N_14636);
or UO_192 (O_192,N_14316,N_14581);
nor UO_193 (O_193,N_14470,N_14510);
xnor UO_194 (O_194,N_14944,N_14639);
and UO_195 (O_195,N_14825,N_14757);
and UO_196 (O_196,N_14810,N_14424);
nor UO_197 (O_197,N_14418,N_14422);
and UO_198 (O_198,N_14867,N_14956);
and UO_199 (O_199,N_14990,N_14967);
and UO_200 (O_200,N_14874,N_14401);
nor UO_201 (O_201,N_14897,N_14605);
nor UO_202 (O_202,N_14628,N_14778);
or UO_203 (O_203,N_14361,N_14818);
and UO_204 (O_204,N_14317,N_14377);
xnor UO_205 (O_205,N_14667,N_14697);
nand UO_206 (O_206,N_14585,N_14985);
and UO_207 (O_207,N_14456,N_14959);
or UO_208 (O_208,N_14365,N_14637);
or UO_209 (O_209,N_14895,N_14707);
nand UO_210 (O_210,N_14580,N_14640);
nand UO_211 (O_211,N_14558,N_14735);
nand UO_212 (O_212,N_14738,N_14650);
and UO_213 (O_213,N_14752,N_14560);
nand UO_214 (O_214,N_14443,N_14405);
or UO_215 (O_215,N_14575,N_14992);
and UO_216 (O_216,N_14276,N_14485);
nand UO_217 (O_217,N_14728,N_14886);
nor UO_218 (O_218,N_14751,N_14356);
or UO_219 (O_219,N_14768,N_14829);
nand UO_220 (O_220,N_14868,N_14592);
and UO_221 (O_221,N_14902,N_14950);
nor UO_222 (O_222,N_14689,N_14540);
nor UO_223 (O_223,N_14406,N_14899);
and UO_224 (O_224,N_14508,N_14589);
or UO_225 (O_225,N_14686,N_14696);
or UO_226 (O_226,N_14576,N_14789);
nor UO_227 (O_227,N_14435,N_14362);
or UO_228 (O_228,N_14386,N_14338);
nand UO_229 (O_229,N_14463,N_14857);
or UO_230 (O_230,N_14836,N_14364);
or UO_231 (O_231,N_14489,N_14353);
and UO_232 (O_232,N_14260,N_14679);
or UO_233 (O_233,N_14770,N_14998);
and UO_234 (O_234,N_14427,N_14767);
and UO_235 (O_235,N_14378,N_14845);
and UO_236 (O_236,N_14520,N_14805);
or UO_237 (O_237,N_14597,N_14281);
and UO_238 (O_238,N_14319,N_14740);
nand UO_239 (O_239,N_14395,N_14643);
nor UO_240 (O_240,N_14290,N_14937);
nor UO_241 (O_241,N_14653,N_14464);
or UO_242 (O_242,N_14838,N_14796);
and UO_243 (O_243,N_14352,N_14691);
nand UO_244 (O_244,N_14827,N_14685);
xnor UO_245 (O_245,N_14795,N_14724);
nor UO_246 (O_246,N_14263,N_14782);
nor UO_247 (O_247,N_14671,N_14504);
nand UO_248 (O_248,N_14617,N_14578);
or UO_249 (O_249,N_14351,N_14714);
nor UO_250 (O_250,N_14816,N_14940);
and UO_251 (O_251,N_14840,N_14859);
and UO_252 (O_252,N_14621,N_14371);
and UO_253 (O_253,N_14548,N_14493);
or UO_254 (O_254,N_14622,N_14646);
or UO_255 (O_255,N_14441,N_14865);
nor UO_256 (O_256,N_14928,N_14797);
nor UO_257 (O_257,N_14669,N_14788);
and UO_258 (O_258,N_14716,N_14503);
nor UO_259 (O_259,N_14564,N_14547);
or UO_260 (O_260,N_14713,N_14802);
nor UO_261 (O_261,N_14596,N_14858);
and UO_262 (O_262,N_14888,N_14613);
nor UO_263 (O_263,N_14623,N_14529);
or UO_264 (O_264,N_14775,N_14327);
and UO_265 (O_265,N_14700,N_14758);
and UO_266 (O_266,N_14474,N_14527);
and UO_267 (O_267,N_14630,N_14798);
nor UO_268 (O_268,N_14730,N_14711);
nor UO_269 (O_269,N_14343,N_14910);
and UO_270 (O_270,N_14732,N_14278);
nor UO_271 (O_271,N_14286,N_14929);
or UO_272 (O_272,N_14497,N_14634);
xor UO_273 (O_273,N_14927,N_14562);
and UO_274 (O_274,N_14413,N_14633);
and UO_275 (O_275,N_14308,N_14792);
or UO_276 (O_276,N_14269,N_14507);
xnor UO_277 (O_277,N_14635,N_14762);
or UO_278 (O_278,N_14369,N_14984);
or UO_279 (O_279,N_14848,N_14701);
nand UO_280 (O_280,N_14568,N_14553);
and UO_281 (O_281,N_14960,N_14526);
nor UO_282 (O_282,N_14498,N_14887);
or UO_283 (O_283,N_14731,N_14823);
and UO_284 (O_284,N_14468,N_14744);
nand UO_285 (O_285,N_14915,N_14916);
or UO_286 (O_286,N_14673,N_14986);
xnor UO_287 (O_287,N_14930,N_14389);
or UO_288 (O_288,N_14476,N_14295);
and UO_289 (O_289,N_14571,N_14706);
nand UO_290 (O_290,N_14373,N_14828);
nand UO_291 (O_291,N_14519,N_14272);
nand UO_292 (O_292,N_14941,N_14629);
nand UO_293 (O_293,N_14884,N_14467);
nand UO_294 (O_294,N_14275,N_14432);
nor UO_295 (O_295,N_14251,N_14938);
nor UO_296 (O_296,N_14288,N_14618);
nor UO_297 (O_297,N_14339,N_14608);
nor UO_298 (O_298,N_14651,N_14936);
and UO_299 (O_299,N_14344,N_14727);
or UO_300 (O_300,N_14544,N_14509);
or UO_301 (O_301,N_14342,N_14862);
xnor UO_302 (O_302,N_14896,N_14533);
nor UO_303 (O_303,N_14787,N_14552);
nor UO_304 (O_304,N_14625,N_14763);
nor UO_305 (O_305,N_14528,N_14340);
nand UO_306 (O_306,N_14963,N_14482);
xor UO_307 (O_307,N_14777,N_14285);
nand UO_308 (O_308,N_14312,N_14794);
nor UO_309 (O_309,N_14703,N_14645);
and UO_310 (O_310,N_14428,N_14496);
and UO_311 (O_311,N_14979,N_14964);
nand UO_312 (O_312,N_14516,N_14846);
and UO_313 (O_313,N_14872,N_14306);
and UO_314 (O_314,N_14765,N_14385);
nand UO_315 (O_315,N_14922,N_14315);
or UO_316 (O_316,N_14791,N_14524);
xnor UO_317 (O_317,N_14619,N_14877);
and UO_318 (O_318,N_14856,N_14839);
xor UO_319 (O_319,N_14283,N_14627);
or UO_320 (O_320,N_14488,N_14324);
nand UO_321 (O_321,N_14252,N_14479);
and UO_322 (O_322,N_14595,N_14718);
nor UO_323 (O_323,N_14945,N_14402);
nor UO_324 (O_324,N_14297,N_14996);
or UO_325 (O_325,N_14844,N_14583);
nor UO_326 (O_326,N_14407,N_14737);
xnor UO_327 (O_327,N_14250,N_14420);
and UO_328 (O_328,N_14861,N_14894);
nand UO_329 (O_329,N_14587,N_14335);
or UO_330 (O_330,N_14905,N_14854);
nor UO_331 (O_331,N_14725,N_14447);
nor UO_332 (O_332,N_14478,N_14559);
nand UO_333 (O_333,N_14346,N_14494);
or UO_334 (O_334,N_14702,N_14935);
xor UO_335 (O_335,N_14566,N_14466);
or UO_336 (O_336,N_14313,N_14999);
nand UO_337 (O_337,N_14761,N_14491);
nor UO_338 (O_338,N_14779,N_14925);
nor UO_339 (O_339,N_14901,N_14815);
and UO_340 (O_340,N_14484,N_14951);
nand UO_341 (O_341,N_14579,N_14931);
nand UO_342 (O_342,N_14891,N_14415);
and UO_343 (O_343,N_14955,N_14594);
and UO_344 (O_344,N_14518,N_14431);
nor UO_345 (O_345,N_14820,N_14942);
and UO_346 (O_346,N_14924,N_14843);
or UO_347 (O_347,N_14712,N_14311);
or UO_348 (O_348,N_14513,N_14387);
nand UO_349 (O_349,N_14684,N_14337);
nand UO_350 (O_350,N_14534,N_14647);
nor UO_351 (O_351,N_14505,N_14764);
and UO_352 (O_352,N_14841,N_14842);
xnor UO_353 (O_353,N_14287,N_14461);
nor UO_354 (O_354,N_14473,N_14786);
and UO_355 (O_355,N_14453,N_14426);
or UO_356 (O_356,N_14739,N_14654);
nor UO_357 (O_357,N_14350,N_14710);
xnor UO_358 (O_358,N_14893,N_14404);
nor UO_359 (O_359,N_14890,N_14723);
nand UO_360 (O_360,N_14876,N_14268);
and UO_361 (O_361,N_14460,N_14355);
nor UO_362 (O_362,N_14965,N_14326);
nand UO_363 (O_363,N_14532,N_14334);
and UO_364 (O_364,N_14375,N_14747);
and UO_365 (O_365,N_14379,N_14270);
nor UO_366 (O_366,N_14954,N_14917);
or UO_367 (O_367,N_14719,N_14680);
nor UO_368 (O_368,N_14970,N_14388);
or UO_369 (O_369,N_14572,N_14309);
or UO_370 (O_370,N_14535,N_14652);
or UO_371 (O_371,N_14949,N_14800);
nor UO_372 (O_372,N_14436,N_14995);
or UO_373 (O_373,N_14271,N_14674);
or UO_374 (O_374,N_14600,N_14683);
xor UO_375 (O_375,N_14418,N_14789);
nor UO_376 (O_376,N_14423,N_14289);
or UO_377 (O_377,N_14319,N_14721);
nand UO_378 (O_378,N_14479,N_14757);
or UO_379 (O_379,N_14872,N_14488);
xor UO_380 (O_380,N_14314,N_14833);
and UO_381 (O_381,N_14573,N_14582);
nand UO_382 (O_382,N_14838,N_14478);
and UO_383 (O_383,N_14461,N_14812);
xor UO_384 (O_384,N_14406,N_14988);
or UO_385 (O_385,N_14804,N_14404);
and UO_386 (O_386,N_14288,N_14854);
or UO_387 (O_387,N_14768,N_14557);
and UO_388 (O_388,N_14569,N_14424);
nand UO_389 (O_389,N_14516,N_14693);
and UO_390 (O_390,N_14355,N_14915);
nor UO_391 (O_391,N_14679,N_14474);
or UO_392 (O_392,N_14639,N_14921);
and UO_393 (O_393,N_14300,N_14316);
nor UO_394 (O_394,N_14581,N_14606);
nand UO_395 (O_395,N_14885,N_14418);
nand UO_396 (O_396,N_14690,N_14251);
or UO_397 (O_397,N_14567,N_14692);
and UO_398 (O_398,N_14661,N_14876);
or UO_399 (O_399,N_14604,N_14793);
nand UO_400 (O_400,N_14251,N_14379);
nand UO_401 (O_401,N_14739,N_14768);
nand UO_402 (O_402,N_14918,N_14771);
xor UO_403 (O_403,N_14364,N_14612);
nor UO_404 (O_404,N_14428,N_14383);
nand UO_405 (O_405,N_14524,N_14612);
nand UO_406 (O_406,N_14682,N_14276);
or UO_407 (O_407,N_14501,N_14514);
or UO_408 (O_408,N_14865,N_14711);
or UO_409 (O_409,N_14334,N_14504);
and UO_410 (O_410,N_14779,N_14327);
or UO_411 (O_411,N_14749,N_14474);
and UO_412 (O_412,N_14911,N_14829);
and UO_413 (O_413,N_14284,N_14850);
and UO_414 (O_414,N_14674,N_14534);
or UO_415 (O_415,N_14619,N_14439);
xor UO_416 (O_416,N_14507,N_14327);
and UO_417 (O_417,N_14347,N_14634);
nor UO_418 (O_418,N_14668,N_14360);
xor UO_419 (O_419,N_14440,N_14496);
or UO_420 (O_420,N_14412,N_14942);
and UO_421 (O_421,N_14574,N_14544);
and UO_422 (O_422,N_14493,N_14714);
nor UO_423 (O_423,N_14397,N_14427);
nor UO_424 (O_424,N_14574,N_14556);
nand UO_425 (O_425,N_14940,N_14773);
xor UO_426 (O_426,N_14622,N_14446);
nor UO_427 (O_427,N_14816,N_14785);
and UO_428 (O_428,N_14663,N_14760);
and UO_429 (O_429,N_14683,N_14467);
or UO_430 (O_430,N_14435,N_14364);
nand UO_431 (O_431,N_14484,N_14362);
xor UO_432 (O_432,N_14562,N_14345);
nor UO_433 (O_433,N_14312,N_14603);
nand UO_434 (O_434,N_14810,N_14562);
and UO_435 (O_435,N_14999,N_14847);
or UO_436 (O_436,N_14906,N_14960);
or UO_437 (O_437,N_14547,N_14779);
xor UO_438 (O_438,N_14879,N_14647);
xor UO_439 (O_439,N_14509,N_14626);
nand UO_440 (O_440,N_14284,N_14376);
nand UO_441 (O_441,N_14955,N_14644);
nand UO_442 (O_442,N_14349,N_14308);
nor UO_443 (O_443,N_14762,N_14652);
or UO_444 (O_444,N_14452,N_14370);
xor UO_445 (O_445,N_14441,N_14952);
nor UO_446 (O_446,N_14997,N_14281);
and UO_447 (O_447,N_14610,N_14869);
and UO_448 (O_448,N_14877,N_14263);
and UO_449 (O_449,N_14349,N_14753);
nor UO_450 (O_450,N_14435,N_14613);
or UO_451 (O_451,N_14978,N_14341);
nand UO_452 (O_452,N_14793,N_14562);
and UO_453 (O_453,N_14514,N_14585);
and UO_454 (O_454,N_14423,N_14959);
xnor UO_455 (O_455,N_14719,N_14504);
xor UO_456 (O_456,N_14339,N_14709);
or UO_457 (O_457,N_14687,N_14837);
and UO_458 (O_458,N_14831,N_14981);
or UO_459 (O_459,N_14735,N_14332);
nor UO_460 (O_460,N_14809,N_14484);
nor UO_461 (O_461,N_14418,N_14271);
or UO_462 (O_462,N_14736,N_14959);
nand UO_463 (O_463,N_14668,N_14484);
and UO_464 (O_464,N_14480,N_14421);
nor UO_465 (O_465,N_14508,N_14915);
nand UO_466 (O_466,N_14865,N_14848);
and UO_467 (O_467,N_14656,N_14899);
nor UO_468 (O_468,N_14354,N_14953);
nand UO_469 (O_469,N_14666,N_14712);
nor UO_470 (O_470,N_14930,N_14408);
or UO_471 (O_471,N_14653,N_14446);
xor UO_472 (O_472,N_14674,N_14282);
and UO_473 (O_473,N_14412,N_14802);
nand UO_474 (O_474,N_14626,N_14974);
and UO_475 (O_475,N_14724,N_14515);
nor UO_476 (O_476,N_14675,N_14921);
nand UO_477 (O_477,N_14801,N_14271);
and UO_478 (O_478,N_14510,N_14835);
nand UO_479 (O_479,N_14627,N_14380);
or UO_480 (O_480,N_14632,N_14289);
nor UO_481 (O_481,N_14409,N_14911);
and UO_482 (O_482,N_14264,N_14936);
nand UO_483 (O_483,N_14326,N_14862);
nand UO_484 (O_484,N_14350,N_14358);
and UO_485 (O_485,N_14355,N_14506);
xor UO_486 (O_486,N_14591,N_14505);
nand UO_487 (O_487,N_14907,N_14883);
nand UO_488 (O_488,N_14768,N_14370);
and UO_489 (O_489,N_14836,N_14283);
or UO_490 (O_490,N_14955,N_14912);
and UO_491 (O_491,N_14547,N_14847);
and UO_492 (O_492,N_14350,N_14562);
or UO_493 (O_493,N_14285,N_14677);
or UO_494 (O_494,N_14588,N_14339);
nor UO_495 (O_495,N_14995,N_14577);
and UO_496 (O_496,N_14830,N_14374);
or UO_497 (O_497,N_14617,N_14406);
or UO_498 (O_498,N_14452,N_14260);
xnor UO_499 (O_499,N_14610,N_14520);
and UO_500 (O_500,N_14748,N_14444);
xnor UO_501 (O_501,N_14937,N_14557);
nand UO_502 (O_502,N_14830,N_14841);
and UO_503 (O_503,N_14880,N_14355);
and UO_504 (O_504,N_14923,N_14714);
or UO_505 (O_505,N_14491,N_14616);
and UO_506 (O_506,N_14725,N_14267);
or UO_507 (O_507,N_14601,N_14650);
xor UO_508 (O_508,N_14601,N_14683);
nor UO_509 (O_509,N_14723,N_14307);
and UO_510 (O_510,N_14730,N_14386);
and UO_511 (O_511,N_14982,N_14318);
nor UO_512 (O_512,N_14977,N_14830);
nor UO_513 (O_513,N_14871,N_14495);
and UO_514 (O_514,N_14268,N_14739);
or UO_515 (O_515,N_14733,N_14759);
nand UO_516 (O_516,N_14814,N_14954);
or UO_517 (O_517,N_14785,N_14562);
and UO_518 (O_518,N_14755,N_14891);
xnor UO_519 (O_519,N_14952,N_14624);
or UO_520 (O_520,N_14460,N_14553);
or UO_521 (O_521,N_14431,N_14779);
or UO_522 (O_522,N_14771,N_14391);
or UO_523 (O_523,N_14457,N_14942);
xnor UO_524 (O_524,N_14981,N_14873);
nand UO_525 (O_525,N_14643,N_14897);
and UO_526 (O_526,N_14917,N_14521);
or UO_527 (O_527,N_14747,N_14782);
or UO_528 (O_528,N_14365,N_14859);
and UO_529 (O_529,N_14405,N_14848);
and UO_530 (O_530,N_14601,N_14594);
xor UO_531 (O_531,N_14498,N_14565);
nor UO_532 (O_532,N_14852,N_14641);
xor UO_533 (O_533,N_14388,N_14498);
xnor UO_534 (O_534,N_14957,N_14707);
nor UO_535 (O_535,N_14543,N_14371);
nand UO_536 (O_536,N_14484,N_14369);
nand UO_537 (O_537,N_14469,N_14709);
and UO_538 (O_538,N_14461,N_14999);
nor UO_539 (O_539,N_14761,N_14367);
nor UO_540 (O_540,N_14369,N_14619);
xnor UO_541 (O_541,N_14740,N_14981);
or UO_542 (O_542,N_14997,N_14381);
nor UO_543 (O_543,N_14729,N_14964);
nor UO_544 (O_544,N_14683,N_14452);
nand UO_545 (O_545,N_14917,N_14748);
nor UO_546 (O_546,N_14407,N_14659);
nand UO_547 (O_547,N_14803,N_14508);
xnor UO_548 (O_548,N_14756,N_14430);
and UO_549 (O_549,N_14774,N_14587);
nor UO_550 (O_550,N_14997,N_14824);
nand UO_551 (O_551,N_14998,N_14411);
xnor UO_552 (O_552,N_14314,N_14405);
or UO_553 (O_553,N_14818,N_14556);
nor UO_554 (O_554,N_14547,N_14927);
nor UO_555 (O_555,N_14470,N_14529);
or UO_556 (O_556,N_14292,N_14702);
nand UO_557 (O_557,N_14976,N_14813);
nand UO_558 (O_558,N_14711,N_14758);
xnor UO_559 (O_559,N_14428,N_14280);
nand UO_560 (O_560,N_14618,N_14549);
or UO_561 (O_561,N_14408,N_14700);
nand UO_562 (O_562,N_14472,N_14938);
or UO_563 (O_563,N_14897,N_14523);
xnor UO_564 (O_564,N_14286,N_14783);
nand UO_565 (O_565,N_14708,N_14579);
xor UO_566 (O_566,N_14438,N_14735);
nand UO_567 (O_567,N_14835,N_14447);
and UO_568 (O_568,N_14775,N_14270);
nand UO_569 (O_569,N_14972,N_14310);
and UO_570 (O_570,N_14496,N_14433);
or UO_571 (O_571,N_14418,N_14953);
and UO_572 (O_572,N_14870,N_14710);
nand UO_573 (O_573,N_14302,N_14955);
nor UO_574 (O_574,N_14444,N_14621);
nor UO_575 (O_575,N_14991,N_14343);
nand UO_576 (O_576,N_14326,N_14278);
nor UO_577 (O_577,N_14548,N_14401);
nor UO_578 (O_578,N_14958,N_14756);
nor UO_579 (O_579,N_14468,N_14797);
xnor UO_580 (O_580,N_14717,N_14988);
nand UO_581 (O_581,N_14649,N_14607);
nand UO_582 (O_582,N_14503,N_14727);
nor UO_583 (O_583,N_14659,N_14772);
or UO_584 (O_584,N_14337,N_14532);
or UO_585 (O_585,N_14677,N_14329);
and UO_586 (O_586,N_14715,N_14946);
nor UO_587 (O_587,N_14634,N_14863);
or UO_588 (O_588,N_14473,N_14579);
or UO_589 (O_589,N_14833,N_14477);
xor UO_590 (O_590,N_14903,N_14991);
xnor UO_591 (O_591,N_14573,N_14757);
and UO_592 (O_592,N_14298,N_14834);
or UO_593 (O_593,N_14448,N_14693);
nor UO_594 (O_594,N_14488,N_14391);
nand UO_595 (O_595,N_14551,N_14708);
or UO_596 (O_596,N_14997,N_14285);
nand UO_597 (O_597,N_14448,N_14804);
or UO_598 (O_598,N_14473,N_14573);
or UO_599 (O_599,N_14719,N_14834);
or UO_600 (O_600,N_14788,N_14652);
nand UO_601 (O_601,N_14573,N_14369);
nor UO_602 (O_602,N_14985,N_14768);
nand UO_603 (O_603,N_14570,N_14381);
or UO_604 (O_604,N_14764,N_14598);
or UO_605 (O_605,N_14581,N_14553);
or UO_606 (O_606,N_14698,N_14625);
xnor UO_607 (O_607,N_14949,N_14983);
or UO_608 (O_608,N_14919,N_14643);
or UO_609 (O_609,N_14795,N_14951);
or UO_610 (O_610,N_14624,N_14336);
nor UO_611 (O_611,N_14533,N_14961);
xor UO_612 (O_612,N_14472,N_14796);
or UO_613 (O_613,N_14477,N_14898);
or UO_614 (O_614,N_14581,N_14863);
nor UO_615 (O_615,N_14270,N_14547);
xor UO_616 (O_616,N_14498,N_14338);
and UO_617 (O_617,N_14503,N_14651);
nor UO_618 (O_618,N_14970,N_14852);
nand UO_619 (O_619,N_14277,N_14994);
xnor UO_620 (O_620,N_14895,N_14983);
or UO_621 (O_621,N_14848,N_14612);
or UO_622 (O_622,N_14693,N_14659);
nor UO_623 (O_623,N_14314,N_14289);
and UO_624 (O_624,N_14480,N_14918);
nand UO_625 (O_625,N_14330,N_14583);
nor UO_626 (O_626,N_14314,N_14728);
and UO_627 (O_627,N_14547,N_14398);
nand UO_628 (O_628,N_14465,N_14700);
and UO_629 (O_629,N_14729,N_14852);
nand UO_630 (O_630,N_14291,N_14654);
nor UO_631 (O_631,N_14374,N_14674);
or UO_632 (O_632,N_14837,N_14487);
and UO_633 (O_633,N_14369,N_14403);
xor UO_634 (O_634,N_14657,N_14650);
or UO_635 (O_635,N_14549,N_14396);
nand UO_636 (O_636,N_14421,N_14869);
or UO_637 (O_637,N_14656,N_14299);
nor UO_638 (O_638,N_14735,N_14391);
nand UO_639 (O_639,N_14622,N_14366);
or UO_640 (O_640,N_14614,N_14557);
nor UO_641 (O_641,N_14711,N_14801);
and UO_642 (O_642,N_14501,N_14709);
nand UO_643 (O_643,N_14274,N_14565);
or UO_644 (O_644,N_14831,N_14862);
and UO_645 (O_645,N_14525,N_14676);
nand UO_646 (O_646,N_14982,N_14316);
xor UO_647 (O_647,N_14546,N_14858);
nand UO_648 (O_648,N_14948,N_14767);
or UO_649 (O_649,N_14683,N_14635);
nor UO_650 (O_650,N_14549,N_14493);
nor UO_651 (O_651,N_14579,N_14813);
nor UO_652 (O_652,N_14788,N_14894);
nand UO_653 (O_653,N_14258,N_14984);
or UO_654 (O_654,N_14726,N_14956);
and UO_655 (O_655,N_14828,N_14332);
and UO_656 (O_656,N_14887,N_14358);
and UO_657 (O_657,N_14501,N_14813);
nor UO_658 (O_658,N_14277,N_14815);
and UO_659 (O_659,N_14630,N_14822);
nor UO_660 (O_660,N_14516,N_14953);
and UO_661 (O_661,N_14722,N_14961);
nand UO_662 (O_662,N_14673,N_14588);
and UO_663 (O_663,N_14887,N_14858);
nor UO_664 (O_664,N_14797,N_14505);
and UO_665 (O_665,N_14275,N_14660);
and UO_666 (O_666,N_14445,N_14417);
nand UO_667 (O_667,N_14551,N_14939);
or UO_668 (O_668,N_14646,N_14540);
nand UO_669 (O_669,N_14699,N_14360);
nor UO_670 (O_670,N_14933,N_14281);
xnor UO_671 (O_671,N_14632,N_14567);
nand UO_672 (O_672,N_14806,N_14951);
or UO_673 (O_673,N_14526,N_14605);
nand UO_674 (O_674,N_14699,N_14490);
nor UO_675 (O_675,N_14620,N_14638);
and UO_676 (O_676,N_14464,N_14823);
or UO_677 (O_677,N_14299,N_14835);
nor UO_678 (O_678,N_14602,N_14906);
or UO_679 (O_679,N_14940,N_14423);
xnor UO_680 (O_680,N_14373,N_14630);
nand UO_681 (O_681,N_14592,N_14430);
nor UO_682 (O_682,N_14478,N_14299);
nor UO_683 (O_683,N_14323,N_14397);
and UO_684 (O_684,N_14651,N_14794);
nand UO_685 (O_685,N_14568,N_14907);
xnor UO_686 (O_686,N_14887,N_14821);
nand UO_687 (O_687,N_14535,N_14266);
xnor UO_688 (O_688,N_14865,N_14505);
xor UO_689 (O_689,N_14448,N_14554);
or UO_690 (O_690,N_14565,N_14696);
and UO_691 (O_691,N_14438,N_14521);
nor UO_692 (O_692,N_14990,N_14802);
nand UO_693 (O_693,N_14931,N_14601);
nor UO_694 (O_694,N_14552,N_14535);
or UO_695 (O_695,N_14330,N_14991);
or UO_696 (O_696,N_14277,N_14963);
nand UO_697 (O_697,N_14674,N_14359);
or UO_698 (O_698,N_14988,N_14736);
nor UO_699 (O_699,N_14691,N_14782);
or UO_700 (O_700,N_14841,N_14366);
nor UO_701 (O_701,N_14744,N_14891);
or UO_702 (O_702,N_14438,N_14470);
and UO_703 (O_703,N_14550,N_14649);
and UO_704 (O_704,N_14967,N_14478);
xor UO_705 (O_705,N_14732,N_14314);
nand UO_706 (O_706,N_14862,N_14769);
and UO_707 (O_707,N_14322,N_14706);
and UO_708 (O_708,N_14304,N_14855);
nor UO_709 (O_709,N_14957,N_14691);
or UO_710 (O_710,N_14951,N_14941);
xor UO_711 (O_711,N_14698,N_14991);
xor UO_712 (O_712,N_14379,N_14974);
nand UO_713 (O_713,N_14800,N_14522);
nor UO_714 (O_714,N_14723,N_14732);
xnor UO_715 (O_715,N_14986,N_14614);
nor UO_716 (O_716,N_14910,N_14983);
xor UO_717 (O_717,N_14388,N_14314);
nand UO_718 (O_718,N_14754,N_14280);
nand UO_719 (O_719,N_14660,N_14514);
or UO_720 (O_720,N_14302,N_14253);
or UO_721 (O_721,N_14480,N_14778);
or UO_722 (O_722,N_14503,N_14256);
and UO_723 (O_723,N_14639,N_14589);
xor UO_724 (O_724,N_14462,N_14736);
or UO_725 (O_725,N_14307,N_14692);
and UO_726 (O_726,N_14396,N_14465);
or UO_727 (O_727,N_14845,N_14351);
nor UO_728 (O_728,N_14413,N_14787);
or UO_729 (O_729,N_14582,N_14687);
nand UO_730 (O_730,N_14547,N_14504);
nand UO_731 (O_731,N_14675,N_14403);
and UO_732 (O_732,N_14408,N_14632);
nand UO_733 (O_733,N_14966,N_14627);
or UO_734 (O_734,N_14282,N_14682);
nor UO_735 (O_735,N_14548,N_14690);
and UO_736 (O_736,N_14915,N_14480);
nand UO_737 (O_737,N_14640,N_14550);
or UO_738 (O_738,N_14704,N_14789);
or UO_739 (O_739,N_14425,N_14980);
nor UO_740 (O_740,N_14796,N_14544);
xor UO_741 (O_741,N_14597,N_14360);
and UO_742 (O_742,N_14885,N_14624);
or UO_743 (O_743,N_14302,N_14298);
and UO_744 (O_744,N_14330,N_14937);
xor UO_745 (O_745,N_14466,N_14672);
or UO_746 (O_746,N_14551,N_14461);
nor UO_747 (O_747,N_14837,N_14683);
and UO_748 (O_748,N_14373,N_14942);
and UO_749 (O_749,N_14583,N_14261);
and UO_750 (O_750,N_14255,N_14843);
nor UO_751 (O_751,N_14264,N_14331);
or UO_752 (O_752,N_14913,N_14534);
nor UO_753 (O_753,N_14339,N_14682);
and UO_754 (O_754,N_14628,N_14943);
or UO_755 (O_755,N_14272,N_14800);
and UO_756 (O_756,N_14360,N_14843);
or UO_757 (O_757,N_14866,N_14325);
xor UO_758 (O_758,N_14690,N_14683);
nor UO_759 (O_759,N_14309,N_14419);
nor UO_760 (O_760,N_14930,N_14330);
nor UO_761 (O_761,N_14689,N_14456);
nand UO_762 (O_762,N_14313,N_14564);
or UO_763 (O_763,N_14901,N_14677);
xor UO_764 (O_764,N_14293,N_14749);
and UO_765 (O_765,N_14428,N_14467);
nand UO_766 (O_766,N_14454,N_14996);
and UO_767 (O_767,N_14784,N_14998);
xor UO_768 (O_768,N_14473,N_14316);
nor UO_769 (O_769,N_14663,N_14814);
or UO_770 (O_770,N_14532,N_14491);
nor UO_771 (O_771,N_14820,N_14680);
or UO_772 (O_772,N_14359,N_14676);
nor UO_773 (O_773,N_14330,N_14269);
nor UO_774 (O_774,N_14811,N_14504);
or UO_775 (O_775,N_14486,N_14279);
xor UO_776 (O_776,N_14713,N_14445);
xnor UO_777 (O_777,N_14930,N_14762);
or UO_778 (O_778,N_14512,N_14920);
xor UO_779 (O_779,N_14877,N_14798);
or UO_780 (O_780,N_14429,N_14740);
nand UO_781 (O_781,N_14620,N_14542);
or UO_782 (O_782,N_14383,N_14452);
xor UO_783 (O_783,N_14438,N_14851);
or UO_784 (O_784,N_14297,N_14459);
nor UO_785 (O_785,N_14866,N_14560);
and UO_786 (O_786,N_14821,N_14373);
or UO_787 (O_787,N_14527,N_14975);
or UO_788 (O_788,N_14763,N_14918);
xnor UO_789 (O_789,N_14843,N_14654);
nand UO_790 (O_790,N_14717,N_14421);
nand UO_791 (O_791,N_14810,N_14790);
or UO_792 (O_792,N_14329,N_14903);
and UO_793 (O_793,N_14813,N_14686);
nand UO_794 (O_794,N_14309,N_14285);
nand UO_795 (O_795,N_14738,N_14320);
and UO_796 (O_796,N_14549,N_14338);
and UO_797 (O_797,N_14766,N_14464);
and UO_798 (O_798,N_14769,N_14956);
and UO_799 (O_799,N_14868,N_14436);
nor UO_800 (O_800,N_14647,N_14593);
or UO_801 (O_801,N_14572,N_14957);
or UO_802 (O_802,N_14993,N_14623);
or UO_803 (O_803,N_14769,N_14504);
and UO_804 (O_804,N_14432,N_14507);
nor UO_805 (O_805,N_14554,N_14801);
or UO_806 (O_806,N_14284,N_14457);
nor UO_807 (O_807,N_14641,N_14478);
xor UO_808 (O_808,N_14443,N_14789);
nor UO_809 (O_809,N_14769,N_14962);
nor UO_810 (O_810,N_14270,N_14604);
nand UO_811 (O_811,N_14750,N_14361);
and UO_812 (O_812,N_14772,N_14740);
nor UO_813 (O_813,N_14803,N_14652);
and UO_814 (O_814,N_14993,N_14867);
nor UO_815 (O_815,N_14505,N_14499);
nor UO_816 (O_816,N_14850,N_14326);
and UO_817 (O_817,N_14436,N_14522);
nand UO_818 (O_818,N_14595,N_14521);
or UO_819 (O_819,N_14710,N_14980);
nand UO_820 (O_820,N_14864,N_14386);
or UO_821 (O_821,N_14534,N_14564);
nor UO_822 (O_822,N_14503,N_14298);
and UO_823 (O_823,N_14388,N_14729);
xnor UO_824 (O_824,N_14783,N_14676);
or UO_825 (O_825,N_14966,N_14620);
nand UO_826 (O_826,N_14557,N_14793);
and UO_827 (O_827,N_14820,N_14943);
nor UO_828 (O_828,N_14398,N_14353);
xor UO_829 (O_829,N_14748,N_14789);
nor UO_830 (O_830,N_14304,N_14518);
nand UO_831 (O_831,N_14451,N_14677);
nand UO_832 (O_832,N_14491,N_14763);
nand UO_833 (O_833,N_14726,N_14854);
or UO_834 (O_834,N_14421,N_14988);
and UO_835 (O_835,N_14765,N_14608);
nand UO_836 (O_836,N_14537,N_14307);
and UO_837 (O_837,N_14397,N_14639);
or UO_838 (O_838,N_14647,N_14457);
nor UO_839 (O_839,N_14870,N_14790);
nand UO_840 (O_840,N_14361,N_14345);
nand UO_841 (O_841,N_14576,N_14301);
nor UO_842 (O_842,N_14739,N_14771);
or UO_843 (O_843,N_14909,N_14536);
nor UO_844 (O_844,N_14879,N_14968);
nand UO_845 (O_845,N_14978,N_14311);
or UO_846 (O_846,N_14837,N_14531);
nand UO_847 (O_847,N_14525,N_14881);
nor UO_848 (O_848,N_14714,N_14752);
and UO_849 (O_849,N_14786,N_14891);
and UO_850 (O_850,N_14755,N_14898);
nand UO_851 (O_851,N_14511,N_14674);
nor UO_852 (O_852,N_14483,N_14313);
xor UO_853 (O_853,N_14288,N_14740);
and UO_854 (O_854,N_14428,N_14478);
and UO_855 (O_855,N_14700,N_14570);
nor UO_856 (O_856,N_14251,N_14540);
or UO_857 (O_857,N_14476,N_14965);
nand UO_858 (O_858,N_14936,N_14941);
xor UO_859 (O_859,N_14384,N_14622);
nand UO_860 (O_860,N_14911,N_14305);
nor UO_861 (O_861,N_14503,N_14323);
nand UO_862 (O_862,N_14614,N_14590);
and UO_863 (O_863,N_14294,N_14464);
nand UO_864 (O_864,N_14780,N_14593);
nor UO_865 (O_865,N_14621,N_14887);
or UO_866 (O_866,N_14282,N_14587);
or UO_867 (O_867,N_14984,N_14699);
xor UO_868 (O_868,N_14349,N_14250);
nor UO_869 (O_869,N_14426,N_14449);
or UO_870 (O_870,N_14407,N_14872);
or UO_871 (O_871,N_14265,N_14676);
and UO_872 (O_872,N_14373,N_14980);
nand UO_873 (O_873,N_14360,N_14869);
and UO_874 (O_874,N_14582,N_14698);
and UO_875 (O_875,N_14811,N_14398);
and UO_876 (O_876,N_14580,N_14592);
xnor UO_877 (O_877,N_14735,N_14952);
and UO_878 (O_878,N_14296,N_14753);
nand UO_879 (O_879,N_14772,N_14724);
or UO_880 (O_880,N_14417,N_14438);
nand UO_881 (O_881,N_14443,N_14711);
or UO_882 (O_882,N_14469,N_14729);
and UO_883 (O_883,N_14846,N_14798);
and UO_884 (O_884,N_14375,N_14973);
nand UO_885 (O_885,N_14775,N_14937);
and UO_886 (O_886,N_14892,N_14379);
xor UO_887 (O_887,N_14962,N_14971);
and UO_888 (O_888,N_14447,N_14763);
nor UO_889 (O_889,N_14817,N_14581);
xor UO_890 (O_890,N_14982,N_14335);
and UO_891 (O_891,N_14569,N_14802);
and UO_892 (O_892,N_14462,N_14466);
or UO_893 (O_893,N_14436,N_14649);
or UO_894 (O_894,N_14559,N_14278);
nor UO_895 (O_895,N_14646,N_14725);
or UO_896 (O_896,N_14584,N_14379);
nand UO_897 (O_897,N_14956,N_14639);
nor UO_898 (O_898,N_14525,N_14273);
or UO_899 (O_899,N_14490,N_14990);
and UO_900 (O_900,N_14705,N_14607);
nor UO_901 (O_901,N_14956,N_14757);
nor UO_902 (O_902,N_14885,N_14571);
nand UO_903 (O_903,N_14265,N_14908);
and UO_904 (O_904,N_14397,N_14476);
or UO_905 (O_905,N_14302,N_14654);
nand UO_906 (O_906,N_14280,N_14480);
and UO_907 (O_907,N_14286,N_14548);
nor UO_908 (O_908,N_14690,N_14442);
nand UO_909 (O_909,N_14257,N_14948);
or UO_910 (O_910,N_14871,N_14854);
nor UO_911 (O_911,N_14767,N_14403);
nor UO_912 (O_912,N_14813,N_14912);
nor UO_913 (O_913,N_14766,N_14413);
and UO_914 (O_914,N_14813,N_14506);
nand UO_915 (O_915,N_14445,N_14250);
xnor UO_916 (O_916,N_14716,N_14304);
nor UO_917 (O_917,N_14457,N_14428);
nor UO_918 (O_918,N_14738,N_14350);
or UO_919 (O_919,N_14710,N_14401);
and UO_920 (O_920,N_14800,N_14892);
or UO_921 (O_921,N_14267,N_14454);
nor UO_922 (O_922,N_14775,N_14296);
nand UO_923 (O_923,N_14884,N_14894);
nand UO_924 (O_924,N_14799,N_14684);
nand UO_925 (O_925,N_14573,N_14360);
and UO_926 (O_926,N_14406,N_14574);
nand UO_927 (O_927,N_14807,N_14724);
or UO_928 (O_928,N_14870,N_14599);
and UO_929 (O_929,N_14581,N_14383);
and UO_930 (O_930,N_14346,N_14924);
and UO_931 (O_931,N_14554,N_14553);
nor UO_932 (O_932,N_14439,N_14682);
and UO_933 (O_933,N_14377,N_14891);
nand UO_934 (O_934,N_14621,N_14423);
or UO_935 (O_935,N_14558,N_14580);
nand UO_936 (O_936,N_14568,N_14562);
xor UO_937 (O_937,N_14368,N_14770);
nand UO_938 (O_938,N_14884,N_14269);
nand UO_939 (O_939,N_14256,N_14603);
and UO_940 (O_940,N_14967,N_14302);
and UO_941 (O_941,N_14769,N_14756);
or UO_942 (O_942,N_14748,N_14922);
and UO_943 (O_943,N_14487,N_14538);
nand UO_944 (O_944,N_14987,N_14404);
and UO_945 (O_945,N_14685,N_14638);
xor UO_946 (O_946,N_14776,N_14900);
nand UO_947 (O_947,N_14833,N_14572);
nor UO_948 (O_948,N_14265,N_14554);
nor UO_949 (O_949,N_14453,N_14365);
nand UO_950 (O_950,N_14904,N_14671);
nand UO_951 (O_951,N_14965,N_14624);
xor UO_952 (O_952,N_14323,N_14313);
nor UO_953 (O_953,N_14392,N_14375);
or UO_954 (O_954,N_14880,N_14491);
and UO_955 (O_955,N_14999,N_14784);
xnor UO_956 (O_956,N_14401,N_14266);
xnor UO_957 (O_957,N_14881,N_14545);
or UO_958 (O_958,N_14618,N_14329);
and UO_959 (O_959,N_14754,N_14275);
and UO_960 (O_960,N_14851,N_14678);
or UO_961 (O_961,N_14477,N_14621);
and UO_962 (O_962,N_14307,N_14893);
xnor UO_963 (O_963,N_14381,N_14412);
nor UO_964 (O_964,N_14468,N_14450);
and UO_965 (O_965,N_14945,N_14273);
or UO_966 (O_966,N_14929,N_14566);
nor UO_967 (O_967,N_14322,N_14551);
or UO_968 (O_968,N_14767,N_14283);
and UO_969 (O_969,N_14682,N_14886);
xnor UO_970 (O_970,N_14505,N_14271);
nand UO_971 (O_971,N_14309,N_14326);
nand UO_972 (O_972,N_14335,N_14357);
or UO_973 (O_973,N_14804,N_14337);
and UO_974 (O_974,N_14933,N_14353);
nand UO_975 (O_975,N_14400,N_14705);
and UO_976 (O_976,N_14649,N_14812);
and UO_977 (O_977,N_14893,N_14748);
nor UO_978 (O_978,N_14981,N_14904);
or UO_979 (O_979,N_14891,N_14989);
nor UO_980 (O_980,N_14810,N_14309);
and UO_981 (O_981,N_14533,N_14381);
nand UO_982 (O_982,N_14735,N_14286);
and UO_983 (O_983,N_14942,N_14626);
or UO_984 (O_984,N_14520,N_14757);
and UO_985 (O_985,N_14628,N_14261);
and UO_986 (O_986,N_14460,N_14608);
nor UO_987 (O_987,N_14759,N_14637);
nor UO_988 (O_988,N_14917,N_14438);
and UO_989 (O_989,N_14664,N_14686);
nor UO_990 (O_990,N_14345,N_14277);
and UO_991 (O_991,N_14317,N_14822);
nand UO_992 (O_992,N_14668,N_14959);
and UO_993 (O_993,N_14780,N_14874);
nor UO_994 (O_994,N_14330,N_14431);
and UO_995 (O_995,N_14512,N_14683);
nand UO_996 (O_996,N_14312,N_14705);
nor UO_997 (O_997,N_14995,N_14940);
xnor UO_998 (O_998,N_14528,N_14296);
nand UO_999 (O_999,N_14993,N_14337);
or UO_1000 (O_1000,N_14389,N_14985);
nand UO_1001 (O_1001,N_14433,N_14751);
or UO_1002 (O_1002,N_14828,N_14736);
nor UO_1003 (O_1003,N_14752,N_14691);
and UO_1004 (O_1004,N_14562,N_14631);
nor UO_1005 (O_1005,N_14976,N_14354);
xnor UO_1006 (O_1006,N_14747,N_14333);
xor UO_1007 (O_1007,N_14775,N_14747);
and UO_1008 (O_1008,N_14509,N_14723);
or UO_1009 (O_1009,N_14961,N_14752);
nor UO_1010 (O_1010,N_14563,N_14446);
and UO_1011 (O_1011,N_14701,N_14270);
nor UO_1012 (O_1012,N_14408,N_14473);
or UO_1013 (O_1013,N_14947,N_14589);
nand UO_1014 (O_1014,N_14565,N_14736);
nor UO_1015 (O_1015,N_14827,N_14800);
nand UO_1016 (O_1016,N_14299,N_14996);
nand UO_1017 (O_1017,N_14709,N_14720);
nand UO_1018 (O_1018,N_14457,N_14350);
nor UO_1019 (O_1019,N_14973,N_14938);
xor UO_1020 (O_1020,N_14737,N_14467);
or UO_1021 (O_1021,N_14761,N_14991);
and UO_1022 (O_1022,N_14381,N_14741);
nor UO_1023 (O_1023,N_14880,N_14764);
nor UO_1024 (O_1024,N_14730,N_14968);
nor UO_1025 (O_1025,N_14703,N_14723);
nor UO_1026 (O_1026,N_14669,N_14617);
and UO_1027 (O_1027,N_14970,N_14418);
nand UO_1028 (O_1028,N_14419,N_14791);
nand UO_1029 (O_1029,N_14660,N_14309);
xor UO_1030 (O_1030,N_14685,N_14253);
or UO_1031 (O_1031,N_14871,N_14915);
nand UO_1032 (O_1032,N_14942,N_14650);
and UO_1033 (O_1033,N_14910,N_14417);
and UO_1034 (O_1034,N_14814,N_14526);
xnor UO_1035 (O_1035,N_14876,N_14479);
nor UO_1036 (O_1036,N_14446,N_14539);
or UO_1037 (O_1037,N_14804,N_14578);
or UO_1038 (O_1038,N_14430,N_14274);
nor UO_1039 (O_1039,N_14749,N_14974);
nand UO_1040 (O_1040,N_14926,N_14740);
and UO_1041 (O_1041,N_14445,N_14561);
or UO_1042 (O_1042,N_14837,N_14892);
or UO_1043 (O_1043,N_14583,N_14518);
and UO_1044 (O_1044,N_14599,N_14637);
nand UO_1045 (O_1045,N_14541,N_14747);
or UO_1046 (O_1046,N_14592,N_14493);
xor UO_1047 (O_1047,N_14270,N_14317);
or UO_1048 (O_1048,N_14397,N_14492);
nand UO_1049 (O_1049,N_14252,N_14695);
or UO_1050 (O_1050,N_14636,N_14882);
xor UO_1051 (O_1051,N_14293,N_14728);
or UO_1052 (O_1052,N_14908,N_14665);
nand UO_1053 (O_1053,N_14288,N_14269);
nand UO_1054 (O_1054,N_14834,N_14997);
nand UO_1055 (O_1055,N_14803,N_14268);
nand UO_1056 (O_1056,N_14769,N_14815);
or UO_1057 (O_1057,N_14531,N_14922);
nor UO_1058 (O_1058,N_14534,N_14530);
nand UO_1059 (O_1059,N_14635,N_14978);
and UO_1060 (O_1060,N_14329,N_14828);
nand UO_1061 (O_1061,N_14342,N_14700);
or UO_1062 (O_1062,N_14313,N_14926);
xor UO_1063 (O_1063,N_14597,N_14979);
nor UO_1064 (O_1064,N_14961,N_14939);
and UO_1065 (O_1065,N_14484,N_14906);
nor UO_1066 (O_1066,N_14493,N_14826);
and UO_1067 (O_1067,N_14955,N_14481);
or UO_1068 (O_1068,N_14869,N_14380);
or UO_1069 (O_1069,N_14989,N_14986);
nand UO_1070 (O_1070,N_14293,N_14939);
or UO_1071 (O_1071,N_14394,N_14774);
nor UO_1072 (O_1072,N_14691,N_14779);
nand UO_1073 (O_1073,N_14404,N_14473);
or UO_1074 (O_1074,N_14419,N_14706);
or UO_1075 (O_1075,N_14365,N_14577);
and UO_1076 (O_1076,N_14303,N_14559);
nand UO_1077 (O_1077,N_14779,N_14821);
nand UO_1078 (O_1078,N_14676,N_14720);
nand UO_1079 (O_1079,N_14713,N_14433);
or UO_1080 (O_1080,N_14878,N_14538);
and UO_1081 (O_1081,N_14380,N_14386);
nor UO_1082 (O_1082,N_14977,N_14851);
nand UO_1083 (O_1083,N_14855,N_14498);
or UO_1084 (O_1084,N_14878,N_14800);
and UO_1085 (O_1085,N_14319,N_14307);
and UO_1086 (O_1086,N_14847,N_14803);
and UO_1087 (O_1087,N_14350,N_14762);
nor UO_1088 (O_1088,N_14318,N_14826);
nand UO_1089 (O_1089,N_14365,N_14689);
xnor UO_1090 (O_1090,N_14257,N_14391);
and UO_1091 (O_1091,N_14634,N_14928);
and UO_1092 (O_1092,N_14326,N_14300);
nand UO_1093 (O_1093,N_14348,N_14807);
and UO_1094 (O_1094,N_14447,N_14703);
or UO_1095 (O_1095,N_14909,N_14779);
and UO_1096 (O_1096,N_14360,N_14974);
and UO_1097 (O_1097,N_14698,N_14767);
or UO_1098 (O_1098,N_14861,N_14592);
xnor UO_1099 (O_1099,N_14749,N_14485);
and UO_1100 (O_1100,N_14475,N_14401);
nand UO_1101 (O_1101,N_14478,N_14601);
and UO_1102 (O_1102,N_14255,N_14401);
and UO_1103 (O_1103,N_14263,N_14674);
or UO_1104 (O_1104,N_14829,N_14807);
or UO_1105 (O_1105,N_14570,N_14463);
nor UO_1106 (O_1106,N_14559,N_14356);
nand UO_1107 (O_1107,N_14722,N_14662);
and UO_1108 (O_1108,N_14894,N_14737);
and UO_1109 (O_1109,N_14297,N_14573);
or UO_1110 (O_1110,N_14941,N_14750);
nor UO_1111 (O_1111,N_14660,N_14270);
and UO_1112 (O_1112,N_14419,N_14699);
nor UO_1113 (O_1113,N_14932,N_14376);
nor UO_1114 (O_1114,N_14867,N_14437);
and UO_1115 (O_1115,N_14947,N_14652);
or UO_1116 (O_1116,N_14540,N_14431);
and UO_1117 (O_1117,N_14541,N_14753);
xor UO_1118 (O_1118,N_14451,N_14623);
nor UO_1119 (O_1119,N_14421,N_14540);
nor UO_1120 (O_1120,N_14305,N_14370);
nand UO_1121 (O_1121,N_14966,N_14911);
nand UO_1122 (O_1122,N_14850,N_14375);
nor UO_1123 (O_1123,N_14718,N_14801);
or UO_1124 (O_1124,N_14671,N_14365);
nor UO_1125 (O_1125,N_14564,N_14726);
nand UO_1126 (O_1126,N_14531,N_14780);
nor UO_1127 (O_1127,N_14939,N_14849);
nor UO_1128 (O_1128,N_14337,N_14564);
or UO_1129 (O_1129,N_14380,N_14693);
nor UO_1130 (O_1130,N_14776,N_14349);
xnor UO_1131 (O_1131,N_14406,N_14486);
nand UO_1132 (O_1132,N_14468,N_14824);
nand UO_1133 (O_1133,N_14680,N_14268);
xor UO_1134 (O_1134,N_14575,N_14374);
xnor UO_1135 (O_1135,N_14614,N_14561);
nor UO_1136 (O_1136,N_14975,N_14650);
nor UO_1137 (O_1137,N_14673,N_14791);
and UO_1138 (O_1138,N_14788,N_14707);
or UO_1139 (O_1139,N_14527,N_14664);
nand UO_1140 (O_1140,N_14870,N_14420);
and UO_1141 (O_1141,N_14825,N_14285);
or UO_1142 (O_1142,N_14711,N_14671);
nor UO_1143 (O_1143,N_14830,N_14819);
nor UO_1144 (O_1144,N_14401,N_14514);
or UO_1145 (O_1145,N_14903,N_14391);
xor UO_1146 (O_1146,N_14935,N_14439);
nor UO_1147 (O_1147,N_14890,N_14970);
or UO_1148 (O_1148,N_14649,N_14840);
nand UO_1149 (O_1149,N_14565,N_14321);
nand UO_1150 (O_1150,N_14258,N_14850);
nand UO_1151 (O_1151,N_14788,N_14739);
or UO_1152 (O_1152,N_14890,N_14813);
or UO_1153 (O_1153,N_14407,N_14438);
nor UO_1154 (O_1154,N_14838,N_14929);
nor UO_1155 (O_1155,N_14721,N_14823);
and UO_1156 (O_1156,N_14981,N_14540);
or UO_1157 (O_1157,N_14264,N_14541);
or UO_1158 (O_1158,N_14252,N_14397);
nand UO_1159 (O_1159,N_14426,N_14897);
and UO_1160 (O_1160,N_14355,N_14370);
and UO_1161 (O_1161,N_14255,N_14533);
and UO_1162 (O_1162,N_14477,N_14423);
nor UO_1163 (O_1163,N_14562,N_14952);
and UO_1164 (O_1164,N_14705,N_14421);
and UO_1165 (O_1165,N_14472,N_14580);
nor UO_1166 (O_1166,N_14764,N_14408);
and UO_1167 (O_1167,N_14314,N_14653);
xor UO_1168 (O_1168,N_14918,N_14538);
or UO_1169 (O_1169,N_14803,N_14865);
and UO_1170 (O_1170,N_14279,N_14451);
nand UO_1171 (O_1171,N_14480,N_14340);
and UO_1172 (O_1172,N_14572,N_14779);
nor UO_1173 (O_1173,N_14510,N_14294);
or UO_1174 (O_1174,N_14742,N_14974);
or UO_1175 (O_1175,N_14260,N_14638);
nor UO_1176 (O_1176,N_14327,N_14734);
and UO_1177 (O_1177,N_14928,N_14807);
nand UO_1178 (O_1178,N_14924,N_14978);
xor UO_1179 (O_1179,N_14366,N_14963);
nor UO_1180 (O_1180,N_14257,N_14323);
nand UO_1181 (O_1181,N_14524,N_14296);
and UO_1182 (O_1182,N_14973,N_14836);
nor UO_1183 (O_1183,N_14926,N_14424);
xor UO_1184 (O_1184,N_14954,N_14336);
and UO_1185 (O_1185,N_14287,N_14780);
or UO_1186 (O_1186,N_14980,N_14669);
nor UO_1187 (O_1187,N_14362,N_14258);
nor UO_1188 (O_1188,N_14875,N_14997);
xnor UO_1189 (O_1189,N_14589,N_14252);
nand UO_1190 (O_1190,N_14762,N_14333);
xor UO_1191 (O_1191,N_14457,N_14966);
nand UO_1192 (O_1192,N_14841,N_14598);
nand UO_1193 (O_1193,N_14778,N_14796);
nor UO_1194 (O_1194,N_14690,N_14637);
nand UO_1195 (O_1195,N_14760,N_14933);
or UO_1196 (O_1196,N_14409,N_14810);
nand UO_1197 (O_1197,N_14506,N_14858);
nand UO_1198 (O_1198,N_14624,N_14890);
nand UO_1199 (O_1199,N_14929,N_14705);
nand UO_1200 (O_1200,N_14707,N_14399);
nand UO_1201 (O_1201,N_14436,N_14700);
nor UO_1202 (O_1202,N_14630,N_14640);
nor UO_1203 (O_1203,N_14414,N_14684);
nor UO_1204 (O_1204,N_14300,N_14309);
nor UO_1205 (O_1205,N_14884,N_14285);
or UO_1206 (O_1206,N_14720,N_14652);
xnor UO_1207 (O_1207,N_14656,N_14854);
nand UO_1208 (O_1208,N_14961,N_14739);
xor UO_1209 (O_1209,N_14648,N_14500);
and UO_1210 (O_1210,N_14816,N_14477);
nand UO_1211 (O_1211,N_14680,N_14510);
nand UO_1212 (O_1212,N_14928,N_14547);
nor UO_1213 (O_1213,N_14663,N_14827);
or UO_1214 (O_1214,N_14442,N_14979);
and UO_1215 (O_1215,N_14440,N_14867);
nand UO_1216 (O_1216,N_14996,N_14689);
or UO_1217 (O_1217,N_14836,N_14785);
nand UO_1218 (O_1218,N_14568,N_14361);
and UO_1219 (O_1219,N_14645,N_14803);
or UO_1220 (O_1220,N_14772,N_14957);
and UO_1221 (O_1221,N_14766,N_14478);
nand UO_1222 (O_1222,N_14576,N_14821);
nor UO_1223 (O_1223,N_14670,N_14265);
nand UO_1224 (O_1224,N_14607,N_14869);
xnor UO_1225 (O_1225,N_14700,N_14614);
nor UO_1226 (O_1226,N_14515,N_14304);
nand UO_1227 (O_1227,N_14894,N_14985);
xor UO_1228 (O_1228,N_14528,N_14890);
nand UO_1229 (O_1229,N_14505,N_14949);
or UO_1230 (O_1230,N_14494,N_14850);
xnor UO_1231 (O_1231,N_14586,N_14593);
or UO_1232 (O_1232,N_14433,N_14499);
xor UO_1233 (O_1233,N_14576,N_14420);
nand UO_1234 (O_1234,N_14701,N_14692);
or UO_1235 (O_1235,N_14586,N_14568);
nor UO_1236 (O_1236,N_14957,N_14535);
nor UO_1237 (O_1237,N_14717,N_14297);
and UO_1238 (O_1238,N_14431,N_14755);
nor UO_1239 (O_1239,N_14489,N_14865);
and UO_1240 (O_1240,N_14533,N_14969);
nor UO_1241 (O_1241,N_14469,N_14938);
or UO_1242 (O_1242,N_14907,N_14718);
nor UO_1243 (O_1243,N_14831,N_14285);
and UO_1244 (O_1244,N_14423,N_14726);
and UO_1245 (O_1245,N_14690,N_14649);
and UO_1246 (O_1246,N_14438,N_14658);
nor UO_1247 (O_1247,N_14312,N_14775);
and UO_1248 (O_1248,N_14398,N_14467);
and UO_1249 (O_1249,N_14631,N_14898);
and UO_1250 (O_1250,N_14950,N_14865);
nor UO_1251 (O_1251,N_14618,N_14317);
or UO_1252 (O_1252,N_14845,N_14623);
nor UO_1253 (O_1253,N_14361,N_14550);
nor UO_1254 (O_1254,N_14260,N_14677);
nand UO_1255 (O_1255,N_14688,N_14496);
nor UO_1256 (O_1256,N_14843,N_14887);
and UO_1257 (O_1257,N_14683,N_14563);
xnor UO_1258 (O_1258,N_14896,N_14828);
nand UO_1259 (O_1259,N_14338,N_14508);
nor UO_1260 (O_1260,N_14684,N_14279);
nor UO_1261 (O_1261,N_14400,N_14973);
and UO_1262 (O_1262,N_14619,N_14631);
or UO_1263 (O_1263,N_14607,N_14320);
nor UO_1264 (O_1264,N_14891,N_14426);
nor UO_1265 (O_1265,N_14570,N_14312);
nor UO_1266 (O_1266,N_14381,N_14718);
or UO_1267 (O_1267,N_14826,N_14422);
nand UO_1268 (O_1268,N_14345,N_14997);
nand UO_1269 (O_1269,N_14732,N_14569);
nand UO_1270 (O_1270,N_14469,N_14604);
and UO_1271 (O_1271,N_14467,N_14918);
nor UO_1272 (O_1272,N_14394,N_14601);
nor UO_1273 (O_1273,N_14421,N_14747);
nor UO_1274 (O_1274,N_14552,N_14998);
and UO_1275 (O_1275,N_14508,N_14301);
nor UO_1276 (O_1276,N_14347,N_14275);
and UO_1277 (O_1277,N_14282,N_14581);
or UO_1278 (O_1278,N_14732,N_14429);
or UO_1279 (O_1279,N_14466,N_14433);
nand UO_1280 (O_1280,N_14871,N_14933);
and UO_1281 (O_1281,N_14549,N_14448);
or UO_1282 (O_1282,N_14340,N_14532);
nand UO_1283 (O_1283,N_14700,N_14561);
and UO_1284 (O_1284,N_14902,N_14952);
nand UO_1285 (O_1285,N_14821,N_14862);
nand UO_1286 (O_1286,N_14304,N_14615);
nor UO_1287 (O_1287,N_14481,N_14631);
nand UO_1288 (O_1288,N_14365,N_14570);
nor UO_1289 (O_1289,N_14461,N_14505);
nor UO_1290 (O_1290,N_14622,N_14504);
or UO_1291 (O_1291,N_14522,N_14387);
nor UO_1292 (O_1292,N_14392,N_14461);
and UO_1293 (O_1293,N_14953,N_14961);
nor UO_1294 (O_1294,N_14435,N_14343);
and UO_1295 (O_1295,N_14585,N_14563);
and UO_1296 (O_1296,N_14440,N_14953);
nor UO_1297 (O_1297,N_14790,N_14890);
or UO_1298 (O_1298,N_14501,N_14973);
and UO_1299 (O_1299,N_14574,N_14733);
xnor UO_1300 (O_1300,N_14308,N_14476);
or UO_1301 (O_1301,N_14934,N_14876);
and UO_1302 (O_1302,N_14898,N_14888);
nand UO_1303 (O_1303,N_14957,N_14687);
and UO_1304 (O_1304,N_14403,N_14318);
or UO_1305 (O_1305,N_14523,N_14354);
or UO_1306 (O_1306,N_14848,N_14598);
and UO_1307 (O_1307,N_14552,N_14261);
and UO_1308 (O_1308,N_14309,N_14743);
and UO_1309 (O_1309,N_14930,N_14388);
nand UO_1310 (O_1310,N_14615,N_14262);
and UO_1311 (O_1311,N_14262,N_14932);
nand UO_1312 (O_1312,N_14326,N_14961);
nor UO_1313 (O_1313,N_14641,N_14596);
or UO_1314 (O_1314,N_14321,N_14603);
nand UO_1315 (O_1315,N_14634,N_14823);
nand UO_1316 (O_1316,N_14484,N_14548);
or UO_1317 (O_1317,N_14546,N_14822);
nand UO_1318 (O_1318,N_14757,N_14631);
nand UO_1319 (O_1319,N_14964,N_14297);
nand UO_1320 (O_1320,N_14930,N_14972);
and UO_1321 (O_1321,N_14825,N_14363);
nor UO_1322 (O_1322,N_14306,N_14428);
nand UO_1323 (O_1323,N_14736,N_14396);
and UO_1324 (O_1324,N_14737,N_14506);
and UO_1325 (O_1325,N_14765,N_14271);
xnor UO_1326 (O_1326,N_14545,N_14935);
and UO_1327 (O_1327,N_14503,N_14550);
or UO_1328 (O_1328,N_14442,N_14667);
or UO_1329 (O_1329,N_14943,N_14301);
or UO_1330 (O_1330,N_14977,N_14460);
and UO_1331 (O_1331,N_14872,N_14593);
and UO_1332 (O_1332,N_14648,N_14554);
or UO_1333 (O_1333,N_14694,N_14717);
or UO_1334 (O_1334,N_14846,N_14320);
or UO_1335 (O_1335,N_14294,N_14264);
xnor UO_1336 (O_1336,N_14749,N_14302);
nand UO_1337 (O_1337,N_14345,N_14941);
and UO_1338 (O_1338,N_14346,N_14702);
xor UO_1339 (O_1339,N_14450,N_14570);
xnor UO_1340 (O_1340,N_14291,N_14964);
nand UO_1341 (O_1341,N_14995,N_14288);
xnor UO_1342 (O_1342,N_14408,N_14817);
and UO_1343 (O_1343,N_14786,N_14425);
or UO_1344 (O_1344,N_14834,N_14461);
nand UO_1345 (O_1345,N_14594,N_14960);
nand UO_1346 (O_1346,N_14908,N_14654);
or UO_1347 (O_1347,N_14754,N_14705);
and UO_1348 (O_1348,N_14274,N_14623);
or UO_1349 (O_1349,N_14350,N_14915);
nand UO_1350 (O_1350,N_14387,N_14890);
xor UO_1351 (O_1351,N_14552,N_14533);
nand UO_1352 (O_1352,N_14696,N_14713);
and UO_1353 (O_1353,N_14298,N_14289);
nor UO_1354 (O_1354,N_14754,N_14790);
nor UO_1355 (O_1355,N_14965,N_14906);
xnor UO_1356 (O_1356,N_14856,N_14766);
and UO_1357 (O_1357,N_14648,N_14355);
nor UO_1358 (O_1358,N_14765,N_14753);
and UO_1359 (O_1359,N_14435,N_14873);
and UO_1360 (O_1360,N_14883,N_14532);
or UO_1361 (O_1361,N_14465,N_14269);
nand UO_1362 (O_1362,N_14826,N_14590);
and UO_1363 (O_1363,N_14503,N_14261);
nor UO_1364 (O_1364,N_14441,N_14730);
or UO_1365 (O_1365,N_14678,N_14789);
and UO_1366 (O_1366,N_14862,N_14762);
nor UO_1367 (O_1367,N_14513,N_14356);
or UO_1368 (O_1368,N_14721,N_14255);
xor UO_1369 (O_1369,N_14663,N_14940);
nor UO_1370 (O_1370,N_14563,N_14428);
nand UO_1371 (O_1371,N_14661,N_14599);
or UO_1372 (O_1372,N_14503,N_14585);
nand UO_1373 (O_1373,N_14562,N_14351);
nor UO_1374 (O_1374,N_14824,N_14623);
nand UO_1375 (O_1375,N_14409,N_14663);
or UO_1376 (O_1376,N_14259,N_14253);
nor UO_1377 (O_1377,N_14731,N_14900);
nor UO_1378 (O_1378,N_14910,N_14508);
nand UO_1379 (O_1379,N_14735,N_14375);
or UO_1380 (O_1380,N_14884,N_14702);
nand UO_1381 (O_1381,N_14682,N_14955);
nor UO_1382 (O_1382,N_14311,N_14538);
or UO_1383 (O_1383,N_14428,N_14416);
nand UO_1384 (O_1384,N_14848,N_14485);
and UO_1385 (O_1385,N_14360,N_14256);
nor UO_1386 (O_1386,N_14525,N_14549);
nand UO_1387 (O_1387,N_14426,N_14527);
nand UO_1388 (O_1388,N_14764,N_14978);
and UO_1389 (O_1389,N_14400,N_14753);
nand UO_1390 (O_1390,N_14721,N_14378);
and UO_1391 (O_1391,N_14360,N_14847);
xor UO_1392 (O_1392,N_14289,N_14740);
nor UO_1393 (O_1393,N_14961,N_14641);
nand UO_1394 (O_1394,N_14363,N_14728);
nor UO_1395 (O_1395,N_14881,N_14467);
nor UO_1396 (O_1396,N_14875,N_14931);
nor UO_1397 (O_1397,N_14976,N_14630);
or UO_1398 (O_1398,N_14603,N_14551);
nor UO_1399 (O_1399,N_14572,N_14461);
nand UO_1400 (O_1400,N_14818,N_14965);
nand UO_1401 (O_1401,N_14665,N_14685);
or UO_1402 (O_1402,N_14760,N_14268);
nand UO_1403 (O_1403,N_14401,N_14841);
nand UO_1404 (O_1404,N_14790,N_14577);
and UO_1405 (O_1405,N_14253,N_14681);
and UO_1406 (O_1406,N_14776,N_14446);
and UO_1407 (O_1407,N_14979,N_14864);
nor UO_1408 (O_1408,N_14391,N_14356);
nand UO_1409 (O_1409,N_14451,N_14597);
nand UO_1410 (O_1410,N_14329,N_14325);
nor UO_1411 (O_1411,N_14477,N_14957);
nor UO_1412 (O_1412,N_14748,N_14250);
nand UO_1413 (O_1413,N_14714,N_14312);
or UO_1414 (O_1414,N_14406,N_14772);
or UO_1415 (O_1415,N_14747,N_14299);
nand UO_1416 (O_1416,N_14541,N_14643);
or UO_1417 (O_1417,N_14721,N_14770);
nor UO_1418 (O_1418,N_14819,N_14508);
xnor UO_1419 (O_1419,N_14368,N_14727);
xor UO_1420 (O_1420,N_14755,N_14737);
nand UO_1421 (O_1421,N_14487,N_14584);
xnor UO_1422 (O_1422,N_14825,N_14514);
and UO_1423 (O_1423,N_14697,N_14768);
nor UO_1424 (O_1424,N_14495,N_14500);
nor UO_1425 (O_1425,N_14675,N_14894);
or UO_1426 (O_1426,N_14752,N_14768);
xor UO_1427 (O_1427,N_14617,N_14423);
or UO_1428 (O_1428,N_14710,N_14990);
nand UO_1429 (O_1429,N_14738,N_14568);
and UO_1430 (O_1430,N_14523,N_14710);
nor UO_1431 (O_1431,N_14991,N_14365);
nand UO_1432 (O_1432,N_14271,N_14452);
or UO_1433 (O_1433,N_14898,N_14468);
nand UO_1434 (O_1434,N_14263,N_14750);
xnor UO_1435 (O_1435,N_14423,N_14489);
nand UO_1436 (O_1436,N_14728,N_14838);
and UO_1437 (O_1437,N_14738,N_14389);
xor UO_1438 (O_1438,N_14883,N_14351);
nor UO_1439 (O_1439,N_14374,N_14648);
nor UO_1440 (O_1440,N_14713,N_14794);
and UO_1441 (O_1441,N_14250,N_14310);
and UO_1442 (O_1442,N_14412,N_14397);
or UO_1443 (O_1443,N_14357,N_14455);
and UO_1444 (O_1444,N_14499,N_14413);
or UO_1445 (O_1445,N_14553,N_14879);
nor UO_1446 (O_1446,N_14624,N_14653);
and UO_1447 (O_1447,N_14294,N_14574);
or UO_1448 (O_1448,N_14719,N_14847);
nand UO_1449 (O_1449,N_14574,N_14848);
nor UO_1450 (O_1450,N_14582,N_14781);
nor UO_1451 (O_1451,N_14292,N_14888);
nand UO_1452 (O_1452,N_14282,N_14276);
nor UO_1453 (O_1453,N_14312,N_14972);
nor UO_1454 (O_1454,N_14331,N_14925);
and UO_1455 (O_1455,N_14389,N_14707);
xor UO_1456 (O_1456,N_14994,N_14764);
nand UO_1457 (O_1457,N_14388,N_14743);
xor UO_1458 (O_1458,N_14576,N_14620);
or UO_1459 (O_1459,N_14609,N_14490);
xnor UO_1460 (O_1460,N_14568,N_14403);
nor UO_1461 (O_1461,N_14891,N_14290);
and UO_1462 (O_1462,N_14431,N_14821);
and UO_1463 (O_1463,N_14525,N_14990);
nand UO_1464 (O_1464,N_14335,N_14607);
and UO_1465 (O_1465,N_14286,N_14676);
or UO_1466 (O_1466,N_14518,N_14396);
nor UO_1467 (O_1467,N_14946,N_14484);
nor UO_1468 (O_1468,N_14479,N_14409);
nor UO_1469 (O_1469,N_14709,N_14410);
xnor UO_1470 (O_1470,N_14252,N_14870);
and UO_1471 (O_1471,N_14939,N_14991);
or UO_1472 (O_1472,N_14363,N_14635);
xor UO_1473 (O_1473,N_14600,N_14539);
nand UO_1474 (O_1474,N_14336,N_14762);
or UO_1475 (O_1475,N_14386,N_14808);
and UO_1476 (O_1476,N_14571,N_14854);
nor UO_1477 (O_1477,N_14792,N_14307);
or UO_1478 (O_1478,N_14684,N_14322);
nand UO_1479 (O_1479,N_14715,N_14513);
or UO_1480 (O_1480,N_14904,N_14989);
nand UO_1481 (O_1481,N_14332,N_14668);
xor UO_1482 (O_1482,N_14593,N_14475);
or UO_1483 (O_1483,N_14889,N_14578);
nor UO_1484 (O_1484,N_14415,N_14276);
and UO_1485 (O_1485,N_14687,N_14357);
and UO_1486 (O_1486,N_14951,N_14966);
xor UO_1487 (O_1487,N_14922,N_14903);
and UO_1488 (O_1488,N_14614,N_14754);
and UO_1489 (O_1489,N_14467,N_14689);
and UO_1490 (O_1490,N_14411,N_14840);
nor UO_1491 (O_1491,N_14796,N_14395);
or UO_1492 (O_1492,N_14296,N_14667);
or UO_1493 (O_1493,N_14453,N_14658);
or UO_1494 (O_1494,N_14467,N_14924);
xnor UO_1495 (O_1495,N_14754,N_14761);
or UO_1496 (O_1496,N_14300,N_14576);
nor UO_1497 (O_1497,N_14981,N_14779);
nor UO_1498 (O_1498,N_14621,N_14767);
and UO_1499 (O_1499,N_14512,N_14650);
nor UO_1500 (O_1500,N_14957,N_14953);
and UO_1501 (O_1501,N_14667,N_14604);
nand UO_1502 (O_1502,N_14409,N_14492);
and UO_1503 (O_1503,N_14447,N_14995);
or UO_1504 (O_1504,N_14502,N_14922);
nand UO_1505 (O_1505,N_14324,N_14251);
nor UO_1506 (O_1506,N_14425,N_14830);
nand UO_1507 (O_1507,N_14434,N_14762);
nor UO_1508 (O_1508,N_14418,N_14850);
and UO_1509 (O_1509,N_14526,N_14531);
and UO_1510 (O_1510,N_14725,N_14969);
or UO_1511 (O_1511,N_14692,N_14721);
and UO_1512 (O_1512,N_14882,N_14515);
xnor UO_1513 (O_1513,N_14260,N_14496);
or UO_1514 (O_1514,N_14481,N_14793);
nor UO_1515 (O_1515,N_14911,N_14795);
nand UO_1516 (O_1516,N_14950,N_14516);
nand UO_1517 (O_1517,N_14321,N_14755);
nor UO_1518 (O_1518,N_14278,N_14677);
or UO_1519 (O_1519,N_14532,N_14372);
xnor UO_1520 (O_1520,N_14281,N_14256);
nand UO_1521 (O_1521,N_14633,N_14820);
nand UO_1522 (O_1522,N_14662,N_14497);
nor UO_1523 (O_1523,N_14597,N_14866);
nor UO_1524 (O_1524,N_14744,N_14385);
or UO_1525 (O_1525,N_14580,N_14853);
nand UO_1526 (O_1526,N_14393,N_14275);
nand UO_1527 (O_1527,N_14893,N_14911);
and UO_1528 (O_1528,N_14543,N_14802);
or UO_1529 (O_1529,N_14498,N_14906);
or UO_1530 (O_1530,N_14362,N_14307);
xnor UO_1531 (O_1531,N_14783,N_14542);
and UO_1532 (O_1532,N_14533,N_14671);
nand UO_1533 (O_1533,N_14812,N_14381);
and UO_1534 (O_1534,N_14577,N_14305);
and UO_1535 (O_1535,N_14687,N_14429);
xnor UO_1536 (O_1536,N_14577,N_14908);
or UO_1537 (O_1537,N_14604,N_14778);
nor UO_1538 (O_1538,N_14507,N_14981);
nor UO_1539 (O_1539,N_14574,N_14285);
or UO_1540 (O_1540,N_14565,N_14548);
nand UO_1541 (O_1541,N_14522,N_14625);
nor UO_1542 (O_1542,N_14786,N_14347);
or UO_1543 (O_1543,N_14887,N_14656);
nor UO_1544 (O_1544,N_14527,N_14666);
and UO_1545 (O_1545,N_14301,N_14463);
nand UO_1546 (O_1546,N_14287,N_14539);
and UO_1547 (O_1547,N_14499,N_14738);
and UO_1548 (O_1548,N_14730,N_14321);
nand UO_1549 (O_1549,N_14927,N_14721);
nor UO_1550 (O_1550,N_14713,N_14505);
and UO_1551 (O_1551,N_14353,N_14257);
or UO_1552 (O_1552,N_14796,N_14750);
nor UO_1553 (O_1553,N_14745,N_14941);
nand UO_1554 (O_1554,N_14292,N_14759);
or UO_1555 (O_1555,N_14969,N_14846);
nor UO_1556 (O_1556,N_14682,N_14853);
nand UO_1557 (O_1557,N_14895,N_14655);
or UO_1558 (O_1558,N_14489,N_14582);
nand UO_1559 (O_1559,N_14346,N_14777);
nand UO_1560 (O_1560,N_14875,N_14832);
nand UO_1561 (O_1561,N_14639,N_14700);
nand UO_1562 (O_1562,N_14452,N_14706);
or UO_1563 (O_1563,N_14407,N_14963);
nand UO_1564 (O_1564,N_14672,N_14797);
and UO_1565 (O_1565,N_14279,N_14437);
xor UO_1566 (O_1566,N_14507,N_14494);
nor UO_1567 (O_1567,N_14732,N_14366);
nor UO_1568 (O_1568,N_14318,N_14465);
or UO_1569 (O_1569,N_14405,N_14299);
xnor UO_1570 (O_1570,N_14625,N_14938);
nor UO_1571 (O_1571,N_14685,N_14333);
and UO_1572 (O_1572,N_14262,N_14457);
nor UO_1573 (O_1573,N_14661,N_14905);
and UO_1574 (O_1574,N_14536,N_14919);
or UO_1575 (O_1575,N_14458,N_14588);
nand UO_1576 (O_1576,N_14990,N_14883);
and UO_1577 (O_1577,N_14662,N_14418);
and UO_1578 (O_1578,N_14621,N_14304);
or UO_1579 (O_1579,N_14699,N_14315);
nor UO_1580 (O_1580,N_14496,N_14954);
nand UO_1581 (O_1581,N_14668,N_14917);
and UO_1582 (O_1582,N_14844,N_14466);
xor UO_1583 (O_1583,N_14279,N_14867);
nand UO_1584 (O_1584,N_14779,N_14931);
nor UO_1585 (O_1585,N_14872,N_14985);
xor UO_1586 (O_1586,N_14763,N_14402);
nand UO_1587 (O_1587,N_14777,N_14605);
nand UO_1588 (O_1588,N_14563,N_14572);
or UO_1589 (O_1589,N_14944,N_14757);
and UO_1590 (O_1590,N_14836,N_14665);
or UO_1591 (O_1591,N_14752,N_14679);
nor UO_1592 (O_1592,N_14477,N_14310);
nor UO_1593 (O_1593,N_14567,N_14938);
nand UO_1594 (O_1594,N_14959,N_14551);
or UO_1595 (O_1595,N_14975,N_14707);
and UO_1596 (O_1596,N_14412,N_14426);
nand UO_1597 (O_1597,N_14313,N_14550);
nand UO_1598 (O_1598,N_14788,N_14699);
nand UO_1599 (O_1599,N_14485,N_14809);
xor UO_1600 (O_1600,N_14292,N_14981);
xnor UO_1601 (O_1601,N_14456,N_14481);
or UO_1602 (O_1602,N_14900,N_14864);
nand UO_1603 (O_1603,N_14321,N_14262);
nor UO_1604 (O_1604,N_14960,N_14687);
xnor UO_1605 (O_1605,N_14903,N_14890);
or UO_1606 (O_1606,N_14269,N_14893);
nand UO_1607 (O_1607,N_14619,N_14603);
xor UO_1608 (O_1608,N_14695,N_14573);
nor UO_1609 (O_1609,N_14881,N_14264);
or UO_1610 (O_1610,N_14724,N_14919);
and UO_1611 (O_1611,N_14507,N_14552);
nand UO_1612 (O_1612,N_14361,N_14922);
and UO_1613 (O_1613,N_14821,N_14626);
nand UO_1614 (O_1614,N_14593,N_14472);
and UO_1615 (O_1615,N_14466,N_14471);
and UO_1616 (O_1616,N_14644,N_14501);
and UO_1617 (O_1617,N_14867,N_14991);
or UO_1618 (O_1618,N_14384,N_14602);
or UO_1619 (O_1619,N_14898,N_14731);
nor UO_1620 (O_1620,N_14907,N_14367);
and UO_1621 (O_1621,N_14711,N_14368);
xor UO_1622 (O_1622,N_14898,N_14552);
nor UO_1623 (O_1623,N_14675,N_14807);
or UO_1624 (O_1624,N_14579,N_14254);
xnor UO_1625 (O_1625,N_14405,N_14404);
nor UO_1626 (O_1626,N_14325,N_14886);
or UO_1627 (O_1627,N_14704,N_14494);
nor UO_1628 (O_1628,N_14448,N_14603);
nand UO_1629 (O_1629,N_14546,N_14603);
and UO_1630 (O_1630,N_14952,N_14662);
and UO_1631 (O_1631,N_14399,N_14999);
and UO_1632 (O_1632,N_14962,N_14554);
or UO_1633 (O_1633,N_14737,N_14580);
and UO_1634 (O_1634,N_14617,N_14627);
nand UO_1635 (O_1635,N_14771,N_14899);
and UO_1636 (O_1636,N_14929,N_14406);
nand UO_1637 (O_1637,N_14250,N_14641);
nor UO_1638 (O_1638,N_14358,N_14890);
or UO_1639 (O_1639,N_14514,N_14477);
or UO_1640 (O_1640,N_14792,N_14485);
or UO_1641 (O_1641,N_14624,N_14926);
and UO_1642 (O_1642,N_14555,N_14532);
xnor UO_1643 (O_1643,N_14958,N_14895);
nand UO_1644 (O_1644,N_14974,N_14459);
nand UO_1645 (O_1645,N_14836,N_14282);
nand UO_1646 (O_1646,N_14937,N_14374);
or UO_1647 (O_1647,N_14750,N_14982);
nand UO_1648 (O_1648,N_14908,N_14286);
nand UO_1649 (O_1649,N_14953,N_14348);
nand UO_1650 (O_1650,N_14858,N_14480);
and UO_1651 (O_1651,N_14388,N_14656);
nor UO_1652 (O_1652,N_14682,N_14974);
xor UO_1653 (O_1653,N_14469,N_14384);
nand UO_1654 (O_1654,N_14835,N_14737);
or UO_1655 (O_1655,N_14371,N_14482);
nand UO_1656 (O_1656,N_14926,N_14816);
or UO_1657 (O_1657,N_14762,N_14515);
or UO_1658 (O_1658,N_14637,N_14953);
nand UO_1659 (O_1659,N_14940,N_14253);
and UO_1660 (O_1660,N_14911,N_14806);
or UO_1661 (O_1661,N_14787,N_14395);
xnor UO_1662 (O_1662,N_14937,N_14946);
and UO_1663 (O_1663,N_14827,N_14865);
nand UO_1664 (O_1664,N_14655,N_14782);
xnor UO_1665 (O_1665,N_14571,N_14461);
nor UO_1666 (O_1666,N_14834,N_14616);
xor UO_1667 (O_1667,N_14838,N_14868);
nor UO_1668 (O_1668,N_14513,N_14308);
nand UO_1669 (O_1669,N_14356,N_14279);
or UO_1670 (O_1670,N_14980,N_14343);
nor UO_1671 (O_1671,N_14435,N_14575);
and UO_1672 (O_1672,N_14274,N_14596);
and UO_1673 (O_1673,N_14645,N_14801);
nand UO_1674 (O_1674,N_14811,N_14327);
and UO_1675 (O_1675,N_14995,N_14338);
or UO_1676 (O_1676,N_14381,N_14584);
xor UO_1677 (O_1677,N_14770,N_14561);
nor UO_1678 (O_1678,N_14505,N_14645);
or UO_1679 (O_1679,N_14533,N_14935);
xnor UO_1680 (O_1680,N_14994,N_14908);
nand UO_1681 (O_1681,N_14916,N_14675);
and UO_1682 (O_1682,N_14336,N_14960);
nand UO_1683 (O_1683,N_14271,N_14835);
nand UO_1684 (O_1684,N_14855,N_14299);
nand UO_1685 (O_1685,N_14523,N_14415);
and UO_1686 (O_1686,N_14307,N_14780);
nor UO_1687 (O_1687,N_14928,N_14282);
xor UO_1688 (O_1688,N_14597,N_14298);
or UO_1689 (O_1689,N_14555,N_14401);
nand UO_1690 (O_1690,N_14450,N_14293);
or UO_1691 (O_1691,N_14673,N_14547);
and UO_1692 (O_1692,N_14947,N_14448);
and UO_1693 (O_1693,N_14753,N_14251);
nor UO_1694 (O_1694,N_14766,N_14489);
or UO_1695 (O_1695,N_14430,N_14432);
nand UO_1696 (O_1696,N_14421,N_14616);
or UO_1697 (O_1697,N_14620,N_14912);
nand UO_1698 (O_1698,N_14501,N_14453);
or UO_1699 (O_1699,N_14828,N_14893);
or UO_1700 (O_1700,N_14803,N_14333);
and UO_1701 (O_1701,N_14264,N_14791);
nand UO_1702 (O_1702,N_14555,N_14665);
or UO_1703 (O_1703,N_14391,N_14679);
nor UO_1704 (O_1704,N_14935,N_14694);
xor UO_1705 (O_1705,N_14400,N_14309);
nor UO_1706 (O_1706,N_14783,N_14432);
nand UO_1707 (O_1707,N_14966,N_14465);
or UO_1708 (O_1708,N_14695,N_14998);
and UO_1709 (O_1709,N_14511,N_14902);
nand UO_1710 (O_1710,N_14889,N_14780);
nand UO_1711 (O_1711,N_14321,N_14546);
and UO_1712 (O_1712,N_14873,N_14294);
or UO_1713 (O_1713,N_14366,N_14419);
nand UO_1714 (O_1714,N_14288,N_14725);
nand UO_1715 (O_1715,N_14914,N_14832);
and UO_1716 (O_1716,N_14433,N_14612);
and UO_1717 (O_1717,N_14449,N_14480);
nand UO_1718 (O_1718,N_14484,N_14507);
and UO_1719 (O_1719,N_14739,N_14919);
and UO_1720 (O_1720,N_14566,N_14293);
and UO_1721 (O_1721,N_14994,N_14883);
nand UO_1722 (O_1722,N_14693,N_14290);
or UO_1723 (O_1723,N_14337,N_14827);
nand UO_1724 (O_1724,N_14950,N_14885);
nand UO_1725 (O_1725,N_14545,N_14917);
or UO_1726 (O_1726,N_14397,N_14513);
nand UO_1727 (O_1727,N_14291,N_14950);
nor UO_1728 (O_1728,N_14977,N_14969);
and UO_1729 (O_1729,N_14677,N_14899);
nand UO_1730 (O_1730,N_14599,N_14993);
nand UO_1731 (O_1731,N_14335,N_14668);
or UO_1732 (O_1732,N_14406,N_14927);
and UO_1733 (O_1733,N_14790,N_14571);
and UO_1734 (O_1734,N_14578,N_14803);
nand UO_1735 (O_1735,N_14580,N_14411);
nand UO_1736 (O_1736,N_14513,N_14316);
nor UO_1737 (O_1737,N_14631,N_14262);
nor UO_1738 (O_1738,N_14317,N_14927);
and UO_1739 (O_1739,N_14587,N_14467);
nand UO_1740 (O_1740,N_14986,N_14275);
or UO_1741 (O_1741,N_14623,N_14891);
xor UO_1742 (O_1742,N_14480,N_14361);
nor UO_1743 (O_1743,N_14979,N_14817);
nand UO_1744 (O_1744,N_14418,N_14521);
and UO_1745 (O_1745,N_14693,N_14715);
nand UO_1746 (O_1746,N_14975,N_14876);
nor UO_1747 (O_1747,N_14455,N_14777);
and UO_1748 (O_1748,N_14868,N_14671);
nor UO_1749 (O_1749,N_14640,N_14519);
nor UO_1750 (O_1750,N_14884,N_14540);
nand UO_1751 (O_1751,N_14838,N_14823);
or UO_1752 (O_1752,N_14319,N_14742);
and UO_1753 (O_1753,N_14881,N_14928);
nor UO_1754 (O_1754,N_14970,N_14462);
nand UO_1755 (O_1755,N_14302,N_14848);
nor UO_1756 (O_1756,N_14712,N_14817);
nor UO_1757 (O_1757,N_14616,N_14685);
and UO_1758 (O_1758,N_14779,N_14595);
nor UO_1759 (O_1759,N_14728,N_14869);
or UO_1760 (O_1760,N_14381,N_14665);
nand UO_1761 (O_1761,N_14975,N_14896);
and UO_1762 (O_1762,N_14763,N_14822);
or UO_1763 (O_1763,N_14293,N_14364);
nor UO_1764 (O_1764,N_14681,N_14552);
nand UO_1765 (O_1765,N_14932,N_14596);
nand UO_1766 (O_1766,N_14993,N_14615);
or UO_1767 (O_1767,N_14356,N_14341);
nand UO_1768 (O_1768,N_14444,N_14512);
or UO_1769 (O_1769,N_14794,N_14805);
and UO_1770 (O_1770,N_14567,N_14589);
and UO_1771 (O_1771,N_14704,N_14432);
and UO_1772 (O_1772,N_14292,N_14939);
xor UO_1773 (O_1773,N_14530,N_14392);
and UO_1774 (O_1774,N_14973,N_14365);
xor UO_1775 (O_1775,N_14934,N_14250);
or UO_1776 (O_1776,N_14387,N_14786);
nand UO_1777 (O_1777,N_14483,N_14928);
nand UO_1778 (O_1778,N_14915,N_14456);
nor UO_1779 (O_1779,N_14913,N_14820);
nand UO_1780 (O_1780,N_14574,N_14489);
nor UO_1781 (O_1781,N_14907,N_14383);
nor UO_1782 (O_1782,N_14929,N_14691);
and UO_1783 (O_1783,N_14681,N_14510);
nor UO_1784 (O_1784,N_14853,N_14961);
or UO_1785 (O_1785,N_14834,N_14456);
nor UO_1786 (O_1786,N_14466,N_14893);
nand UO_1787 (O_1787,N_14799,N_14304);
nor UO_1788 (O_1788,N_14484,N_14297);
xor UO_1789 (O_1789,N_14747,N_14481);
and UO_1790 (O_1790,N_14870,N_14407);
nor UO_1791 (O_1791,N_14703,N_14632);
and UO_1792 (O_1792,N_14816,N_14447);
nor UO_1793 (O_1793,N_14956,N_14502);
or UO_1794 (O_1794,N_14562,N_14285);
nor UO_1795 (O_1795,N_14969,N_14382);
and UO_1796 (O_1796,N_14672,N_14518);
nor UO_1797 (O_1797,N_14964,N_14283);
or UO_1798 (O_1798,N_14780,N_14940);
or UO_1799 (O_1799,N_14995,N_14252);
or UO_1800 (O_1800,N_14281,N_14658);
and UO_1801 (O_1801,N_14566,N_14324);
nor UO_1802 (O_1802,N_14811,N_14265);
xnor UO_1803 (O_1803,N_14399,N_14937);
nor UO_1804 (O_1804,N_14443,N_14628);
or UO_1805 (O_1805,N_14358,N_14812);
and UO_1806 (O_1806,N_14459,N_14340);
or UO_1807 (O_1807,N_14325,N_14251);
or UO_1808 (O_1808,N_14489,N_14427);
or UO_1809 (O_1809,N_14500,N_14840);
nand UO_1810 (O_1810,N_14732,N_14838);
nand UO_1811 (O_1811,N_14759,N_14833);
nor UO_1812 (O_1812,N_14856,N_14888);
and UO_1813 (O_1813,N_14452,N_14495);
and UO_1814 (O_1814,N_14893,N_14329);
and UO_1815 (O_1815,N_14759,N_14252);
nand UO_1816 (O_1816,N_14315,N_14817);
nand UO_1817 (O_1817,N_14513,N_14692);
or UO_1818 (O_1818,N_14561,N_14722);
nor UO_1819 (O_1819,N_14419,N_14271);
and UO_1820 (O_1820,N_14647,N_14737);
nand UO_1821 (O_1821,N_14653,N_14642);
and UO_1822 (O_1822,N_14717,N_14437);
xor UO_1823 (O_1823,N_14886,N_14865);
or UO_1824 (O_1824,N_14987,N_14516);
nor UO_1825 (O_1825,N_14626,N_14475);
or UO_1826 (O_1826,N_14428,N_14881);
nand UO_1827 (O_1827,N_14705,N_14420);
nor UO_1828 (O_1828,N_14997,N_14517);
or UO_1829 (O_1829,N_14301,N_14427);
or UO_1830 (O_1830,N_14508,N_14963);
nor UO_1831 (O_1831,N_14266,N_14933);
nand UO_1832 (O_1832,N_14347,N_14832);
nand UO_1833 (O_1833,N_14976,N_14549);
and UO_1834 (O_1834,N_14882,N_14926);
and UO_1835 (O_1835,N_14464,N_14404);
nand UO_1836 (O_1836,N_14908,N_14832);
nand UO_1837 (O_1837,N_14434,N_14370);
and UO_1838 (O_1838,N_14871,N_14739);
nand UO_1839 (O_1839,N_14926,N_14515);
xnor UO_1840 (O_1840,N_14752,N_14541);
and UO_1841 (O_1841,N_14362,N_14686);
and UO_1842 (O_1842,N_14763,N_14530);
nand UO_1843 (O_1843,N_14830,N_14493);
nor UO_1844 (O_1844,N_14673,N_14699);
nor UO_1845 (O_1845,N_14463,N_14908);
nor UO_1846 (O_1846,N_14385,N_14786);
nand UO_1847 (O_1847,N_14342,N_14958);
nand UO_1848 (O_1848,N_14565,N_14646);
and UO_1849 (O_1849,N_14964,N_14586);
nor UO_1850 (O_1850,N_14689,N_14328);
nor UO_1851 (O_1851,N_14534,N_14593);
nand UO_1852 (O_1852,N_14354,N_14512);
and UO_1853 (O_1853,N_14690,N_14964);
xor UO_1854 (O_1854,N_14861,N_14996);
nand UO_1855 (O_1855,N_14621,N_14777);
or UO_1856 (O_1856,N_14882,N_14682);
and UO_1857 (O_1857,N_14805,N_14738);
nand UO_1858 (O_1858,N_14529,N_14554);
and UO_1859 (O_1859,N_14572,N_14301);
nand UO_1860 (O_1860,N_14600,N_14597);
nor UO_1861 (O_1861,N_14876,N_14977);
or UO_1862 (O_1862,N_14444,N_14875);
and UO_1863 (O_1863,N_14815,N_14418);
nor UO_1864 (O_1864,N_14931,N_14614);
nand UO_1865 (O_1865,N_14319,N_14680);
and UO_1866 (O_1866,N_14857,N_14842);
nor UO_1867 (O_1867,N_14909,N_14565);
nor UO_1868 (O_1868,N_14766,N_14788);
and UO_1869 (O_1869,N_14395,N_14411);
nor UO_1870 (O_1870,N_14848,N_14681);
nor UO_1871 (O_1871,N_14896,N_14451);
nand UO_1872 (O_1872,N_14783,N_14485);
or UO_1873 (O_1873,N_14647,N_14753);
and UO_1874 (O_1874,N_14937,N_14505);
xnor UO_1875 (O_1875,N_14646,N_14576);
nand UO_1876 (O_1876,N_14864,N_14426);
nor UO_1877 (O_1877,N_14524,N_14277);
and UO_1878 (O_1878,N_14426,N_14647);
xor UO_1879 (O_1879,N_14644,N_14522);
or UO_1880 (O_1880,N_14685,N_14873);
or UO_1881 (O_1881,N_14312,N_14750);
nand UO_1882 (O_1882,N_14411,N_14812);
and UO_1883 (O_1883,N_14460,N_14414);
and UO_1884 (O_1884,N_14442,N_14793);
and UO_1885 (O_1885,N_14724,N_14468);
or UO_1886 (O_1886,N_14842,N_14401);
and UO_1887 (O_1887,N_14725,N_14813);
and UO_1888 (O_1888,N_14419,N_14718);
and UO_1889 (O_1889,N_14990,N_14721);
xnor UO_1890 (O_1890,N_14333,N_14633);
nor UO_1891 (O_1891,N_14821,N_14793);
and UO_1892 (O_1892,N_14276,N_14260);
or UO_1893 (O_1893,N_14539,N_14308);
and UO_1894 (O_1894,N_14642,N_14693);
nand UO_1895 (O_1895,N_14718,N_14818);
and UO_1896 (O_1896,N_14637,N_14344);
and UO_1897 (O_1897,N_14671,N_14675);
nor UO_1898 (O_1898,N_14478,N_14522);
or UO_1899 (O_1899,N_14380,N_14488);
nand UO_1900 (O_1900,N_14570,N_14318);
nor UO_1901 (O_1901,N_14977,N_14502);
nand UO_1902 (O_1902,N_14505,N_14327);
or UO_1903 (O_1903,N_14623,N_14425);
nand UO_1904 (O_1904,N_14695,N_14721);
or UO_1905 (O_1905,N_14803,N_14907);
and UO_1906 (O_1906,N_14854,N_14735);
nor UO_1907 (O_1907,N_14741,N_14430);
and UO_1908 (O_1908,N_14605,N_14837);
nand UO_1909 (O_1909,N_14282,N_14802);
xor UO_1910 (O_1910,N_14363,N_14873);
nor UO_1911 (O_1911,N_14294,N_14412);
nor UO_1912 (O_1912,N_14512,N_14835);
and UO_1913 (O_1913,N_14809,N_14706);
or UO_1914 (O_1914,N_14716,N_14637);
nand UO_1915 (O_1915,N_14502,N_14809);
nand UO_1916 (O_1916,N_14638,N_14268);
or UO_1917 (O_1917,N_14660,N_14889);
nand UO_1918 (O_1918,N_14877,N_14312);
or UO_1919 (O_1919,N_14692,N_14544);
and UO_1920 (O_1920,N_14774,N_14302);
nand UO_1921 (O_1921,N_14328,N_14596);
nor UO_1922 (O_1922,N_14839,N_14564);
nand UO_1923 (O_1923,N_14592,N_14609);
nand UO_1924 (O_1924,N_14406,N_14958);
and UO_1925 (O_1925,N_14627,N_14976);
nand UO_1926 (O_1926,N_14603,N_14707);
nand UO_1927 (O_1927,N_14264,N_14775);
or UO_1928 (O_1928,N_14650,N_14678);
nand UO_1929 (O_1929,N_14475,N_14951);
or UO_1930 (O_1930,N_14530,N_14997);
nor UO_1931 (O_1931,N_14745,N_14630);
nand UO_1932 (O_1932,N_14864,N_14747);
nor UO_1933 (O_1933,N_14613,N_14518);
or UO_1934 (O_1934,N_14999,N_14719);
nand UO_1935 (O_1935,N_14984,N_14461);
nand UO_1936 (O_1936,N_14875,N_14993);
xnor UO_1937 (O_1937,N_14770,N_14589);
nand UO_1938 (O_1938,N_14367,N_14538);
nand UO_1939 (O_1939,N_14992,N_14541);
nor UO_1940 (O_1940,N_14986,N_14335);
nor UO_1941 (O_1941,N_14535,N_14507);
or UO_1942 (O_1942,N_14869,N_14787);
nor UO_1943 (O_1943,N_14993,N_14317);
and UO_1944 (O_1944,N_14957,N_14705);
or UO_1945 (O_1945,N_14612,N_14414);
nand UO_1946 (O_1946,N_14800,N_14527);
or UO_1947 (O_1947,N_14876,N_14530);
nand UO_1948 (O_1948,N_14321,N_14706);
nand UO_1949 (O_1949,N_14631,N_14737);
and UO_1950 (O_1950,N_14513,N_14757);
xnor UO_1951 (O_1951,N_14595,N_14482);
nand UO_1952 (O_1952,N_14723,N_14719);
nand UO_1953 (O_1953,N_14555,N_14723);
and UO_1954 (O_1954,N_14984,N_14470);
or UO_1955 (O_1955,N_14316,N_14846);
nand UO_1956 (O_1956,N_14328,N_14394);
and UO_1957 (O_1957,N_14483,N_14440);
nor UO_1958 (O_1958,N_14857,N_14689);
nand UO_1959 (O_1959,N_14994,N_14494);
nand UO_1960 (O_1960,N_14425,N_14593);
or UO_1961 (O_1961,N_14474,N_14295);
nand UO_1962 (O_1962,N_14269,N_14353);
or UO_1963 (O_1963,N_14480,N_14380);
or UO_1964 (O_1964,N_14432,N_14323);
or UO_1965 (O_1965,N_14628,N_14716);
and UO_1966 (O_1966,N_14676,N_14989);
and UO_1967 (O_1967,N_14318,N_14363);
or UO_1968 (O_1968,N_14520,N_14871);
xor UO_1969 (O_1969,N_14674,N_14965);
and UO_1970 (O_1970,N_14385,N_14403);
and UO_1971 (O_1971,N_14341,N_14858);
or UO_1972 (O_1972,N_14688,N_14332);
nor UO_1973 (O_1973,N_14478,N_14467);
xor UO_1974 (O_1974,N_14483,N_14934);
nand UO_1975 (O_1975,N_14635,N_14455);
and UO_1976 (O_1976,N_14406,N_14720);
nor UO_1977 (O_1977,N_14375,N_14575);
xnor UO_1978 (O_1978,N_14706,N_14530);
nor UO_1979 (O_1979,N_14822,N_14656);
nand UO_1980 (O_1980,N_14812,N_14347);
nand UO_1981 (O_1981,N_14854,N_14479);
or UO_1982 (O_1982,N_14389,N_14945);
or UO_1983 (O_1983,N_14312,N_14440);
nor UO_1984 (O_1984,N_14278,N_14843);
or UO_1985 (O_1985,N_14666,N_14473);
and UO_1986 (O_1986,N_14812,N_14657);
nand UO_1987 (O_1987,N_14725,N_14636);
nand UO_1988 (O_1988,N_14613,N_14356);
nor UO_1989 (O_1989,N_14485,N_14710);
nor UO_1990 (O_1990,N_14817,N_14683);
nand UO_1991 (O_1991,N_14376,N_14297);
and UO_1992 (O_1992,N_14835,N_14387);
and UO_1993 (O_1993,N_14800,N_14746);
nor UO_1994 (O_1994,N_14877,N_14491);
nand UO_1995 (O_1995,N_14311,N_14658);
nor UO_1996 (O_1996,N_14775,N_14360);
xnor UO_1997 (O_1997,N_14977,N_14677);
and UO_1998 (O_1998,N_14573,N_14699);
nand UO_1999 (O_1999,N_14410,N_14951);
endmodule