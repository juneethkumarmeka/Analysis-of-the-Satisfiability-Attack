module basic_1500_15000_2000_20_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nand U0 (N_0,In_504,In_1026);
or U1 (N_1,In_523,In_512);
nand U2 (N_2,In_196,In_859);
nor U3 (N_3,In_437,In_1057);
and U4 (N_4,In_372,In_48);
nand U5 (N_5,In_339,In_945);
and U6 (N_6,In_726,In_1473);
xnor U7 (N_7,In_389,In_375);
xor U8 (N_8,In_684,In_1127);
xor U9 (N_9,In_842,In_1114);
and U10 (N_10,In_1226,In_1218);
xor U11 (N_11,In_1009,In_1496);
and U12 (N_12,In_45,In_325);
or U13 (N_13,In_176,In_97);
nor U14 (N_14,In_377,In_970);
or U15 (N_15,In_787,In_431);
nor U16 (N_16,In_204,In_661);
or U17 (N_17,In_317,In_526);
nand U18 (N_18,In_588,In_876);
or U19 (N_19,In_995,In_1340);
and U20 (N_20,In_1411,In_1086);
nand U21 (N_21,In_770,In_591);
nor U22 (N_22,In_1069,In_595);
and U23 (N_23,In_1171,In_484);
and U24 (N_24,In_1314,In_1157);
and U25 (N_25,In_471,In_709);
or U26 (N_26,In_1083,In_1214);
nor U27 (N_27,In_837,In_302);
nand U28 (N_28,In_1084,In_1391);
or U29 (N_29,In_1184,In_756);
xnor U30 (N_30,In_7,In_1401);
or U31 (N_31,In_1284,In_1134);
or U32 (N_32,In_956,In_486);
nor U33 (N_33,In_229,In_1358);
nor U34 (N_34,In_269,In_566);
and U35 (N_35,In_1167,In_1356);
nor U36 (N_36,In_965,In_906);
or U37 (N_37,In_332,In_259);
nor U38 (N_38,In_1308,In_346);
and U39 (N_39,In_524,In_16);
and U40 (N_40,In_489,In_134);
or U41 (N_41,In_1387,In_1395);
nor U42 (N_42,In_92,In_345);
and U43 (N_43,In_42,In_1166);
nand U44 (N_44,In_503,In_1095);
and U45 (N_45,In_112,In_470);
or U46 (N_46,In_386,In_133);
nor U47 (N_47,In_1475,In_1079);
nand U48 (N_48,In_1379,In_1264);
nor U49 (N_49,In_147,In_931);
and U50 (N_50,In_115,In_746);
nor U51 (N_51,In_2,In_232);
and U52 (N_52,In_505,In_208);
or U53 (N_53,In_950,In_579);
nand U54 (N_54,In_899,In_412);
xnor U55 (N_55,In_43,In_1372);
and U56 (N_56,In_8,In_458);
nand U57 (N_57,In_828,In_193);
or U58 (N_58,In_5,In_1062);
nor U59 (N_59,In_773,In_795);
nor U60 (N_60,In_334,In_1036);
nand U61 (N_61,In_1266,In_1326);
nor U62 (N_62,In_407,In_761);
nand U63 (N_63,In_29,In_933);
nand U64 (N_64,In_264,In_285);
and U65 (N_65,In_953,In_319);
and U66 (N_66,In_844,In_780);
nand U67 (N_67,In_515,In_442);
or U68 (N_68,In_1133,In_910);
xor U69 (N_69,In_20,In_144);
nand U70 (N_70,In_974,In_573);
nand U71 (N_71,In_741,In_1193);
or U72 (N_72,In_1149,In_1113);
and U73 (N_73,In_693,In_559);
nand U74 (N_74,In_744,In_501);
nor U75 (N_75,In_668,In_1003);
nor U76 (N_76,In_767,In_1495);
or U77 (N_77,In_294,In_1025);
nor U78 (N_78,In_478,In_1354);
nor U79 (N_79,In_244,In_1389);
or U80 (N_80,In_823,In_301);
and U81 (N_81,In_13,In_877);
xor U82 (N_82,In_628,In_18);
nor U83 (N_83,In_1229,In_1492);
nand U84 (N_84,In_9,In_1038);
nand U85 (N_85,In_649,In_641);
or U86 (N_86,In_961,In_104);
nor U87 (N_87,In_316,In_1111);
nor U88 (N_88,In_242,In_251);
xnor U89 (N_89,In_1055,In_1408);
or U90 (N_90,In_398,In_256);
nand U91 (N_91,In_131,In_711);
or U92 (N_92,In_1257,In_519);
nand U93 (N_93,In_885,In_587);
nand U94 (N_94,In_141,In_195);
or U95 (N_95,In_280,In_1047);
and U96 (N_96,In_1219,In_1393);
or U97 (N_97,In_1405,In_882);
or U98 (N_98,In_827,In_1309);
nor U99 (N_99,In_420,In_89);
or U100 (N_100,In_1297,In_593);
nand U101 (N_101,In_297,In_660);
or U102 (N_102,In_718,In_646);
nand U103 (N_103,In_93,In_26);
nor U104 (N_104,In_771,In_76);
nand U105 (N_105,In_1263,In_1353);
or U106 (N_106,In_1454,In_1285);
nand U107 (N_107,In_1165,In_794);
and U108 (N_108,In_373,In_769);
and U109 (N_109,In_1472,In_288);
or U110 (N_110,In_1436,In_328);
nor U111 (N_111,In_967,In_686);
and U112 (N_112,In_1082,In_198);
and U113 (N_113,In_142,In_1203);
and U114 (N_114,In_1190,In_27);
or U115 (N_115,In_311,In_333);
nand U116 (N_116,In_1331,In_562);
or U117 (N_117,In_962,In_1129);
nor U118 (N_118,In_154,In_781);
and U119 (N_119,In_463,In_1078);
nand U120 (N_120,In_922,In_243);
and U121 (N_121,In_1279,In_347);
nand U122 (N_122,In_1359,In_450);
nand U123 (N_123,In_62,In_1092);
nor U124 (N_124,In_582,In_749);
nand U125 (N_125,In_949,In_1384);
and U126 (N_126,In_534,In_1247);
nor U127 (N_127,In_103,In_1020);
xor U128 (N_128,In_19,In_617);
nand U129 (N_129,In_283,In_991);
nor U130 (N_130,In_1256,In_202);
or U131 (N_131,In_905,In_127);
nor U132 (N_132,In_447,In_890);
xnor U133 (N_133,In_1346,In_396);
or U134 (N_134,In_1231,In_577);
or U135 (N_135,In_875,In_541);
nand U136 (N_136,In_988,In_1216);
nor U137 (N_137,In_1132,In_1243);
and U138 (N_138,In_1146,In_723);
xor U139 (N_139,In_427,In_1463);
or U140 (N_140,In_779,In_122);
nand U141 (N_141,In_737,In_706);
xor U142 (N_142,In_547,In_710);
nor U143 (N_143,In_629,In_639);
xnor U144 (N_144,In_344,In_1435);
nor U145 (N_145,In_804,In_246);
nor U146 (N_146,In_535,In_155);
xor U147 (N_147,In_410,In_1105);
nand U148 (N_148,In_1179,In_1089);
or U149 (N_149,In_370,In_776);
or U150 (N_150,In_192,In_1310);
nor U151 (N_151,In_214,In_327);
nand U152 (N_152,In_607,In_531);
nand U153 (N_153,In_934,In_125);
and U154 (N_154,In_847,In_1438);
nand U155 (N_155,In_772,In_262);
or U156 (N_156,In_855,In_15);
and U157 (N_157,In_453,In_209);
nand U158 (N_158,In_455,In_1017);
and U159 (N_159,In_382,In_762);
nor U160 (N_160,In_1224,In_464);
and U161 (N_161,In_1059,In_1427);
xor U162 (N_162,In_1160,In_932);
nor U163 (N_163,In_221,In_1044);
nor U164 (N_164,In_331,In_1298);
nand U165 (N_165,In_1470,In_376);
and U166 (N_166,In_704,In_355);
nor U167 (N_167,In_1367,In_1209);
and U168 (N_168,In_391,In_581);
nand U169 (N_169,In_1324,In_1177);
xnor U170 (N_170,In_436,In_378);
and U171 (N_171,In_850,In_1434);
or U172 (N_172,In_1148,In_830);
nand U173 (N_173,In_1156,In_1428);
nand U174 (N_174,In_615,In_439);
and U175 (N_175,In_1011,In_201);
or U176 (N_176,In_1103,In_782);
nor U177 (N_177,In_49,In_969);
xor U178 (N_178,In_492,In_477);
nand U179 (N_179,In_656,In_529);
nand U180 (N_180,In_895,In_1251);
nand U181 (N_181,In_819,In_96);
or U182 (N_182,In_879,In_241);
and U183 (N_183,In_408,In_400);
or U184 (N_184,In_1422,In_696);
or U185 (N_185,In_1242,In_338);
nor U186 (N_186,In_824,In_921);
or U187 (N_187,In_1466,In_924);
and U188 (N_188,In_1468,In_100);
and U189 (N_189,In_691,In_1016);
and U190 (N_190,In_496,In_465);
and U191 (N_191,In_444,In_483);
and U192 (N_192,In_1029,In_1345);
nand U193 (N_193,In_665,In_371);
and U194 (N_194,In_799,In_894);
or U195 (N_195,In_688,In_1106);
or U196 (N_196,In_912,In_226);
nand U197 (N_197,In_203,In_145);
nor U198 (N_198,In_1291,In_360);
nand U199 (N_199,In_1486,In_669);
and U200 (N_200,In_831,In_871);
nand U201 (N_201,In_1325,In_25);
nand U202 (N_202,In_816,In_815);
nand U203 (N_203,In_1212,In_1151);
or U204 (N_204,In_1043,In_1090);
xnor U205 (N_205,In_733,In_1338);
and U206 (N_206,In_1437,In_1108);
and U207 (N_207,In_1474,In_809);
or U208 (N_208,In_705,In_1123);
nand U209 (N_209,In_755,In_1244);
or U210 (N_210,In_715,In_643);
or U211 (N_211,In_296,In_516);
xor U212 (N_212,In_1066,In_1006);
or U213 (N_213,In_468,In_521);
and U214 (N_214,In_250,In_887);
nand U215 (N_215,In_1211,In_681);
nand U216 (N_216,In_735,In_888);
nand U217 (N_217,In_168,In_110);
xor U218 (N_218,In_884,In_1339);
xnor U219 (N_219,In_1176,In_774);
or U220 (N_220,In_611,In_724);
or U221 (N_221,In_1140,In_286);
nand U222 (N_222,In_12,In_846);
and U223 (N_223,In_1420,In_307);
nor U224 (N_224,In_305,In_68);
nor U225 (N_225,In_1,In_653);
nand U226 (N_226,In_1164,In_758);
or U227 (N_227,In_275,In_182);
or U228 (N_228,In_475,In_367);
nand U229 (N_229,In_1377,In_443);
and U230 (N_230,In_699,In_1077);
and U231 (N_231,In_445,In_1144);
and U232 (N_232,In_676,In_982);
nor U233 (N_233,In_151,In_480);
xnor U234 (N_234,In_36,In_536);
or U235 (N_235,In_1450,In_1227);
nor U236 (N_236,In_146,In_1259);
nand U237 (N_237,In_864,In_1099);
nand U238 (N_238,In_109,In_449);
nor U239 (N_239,In_261,In_1185);
and U240 (N_240,In_1199,In_1444);
or U241 (N_241,In_171,In_813);
nand U242 (N_242,In_1058,In_1478);
nand U243 (N_243,In_1008,In_948);
and U244 (N_244,In_231,In_418);
nor U245 (N_245,In_754,In_1252);
nor U246 (N_246,In_245,In_268);
or U247 (N_247,In_1366,In_1415);
nor U248 (N_248,In_395,In_1225);
nor U249 (N_249,In_1182,In_805);
and U250 (N_250,In_272,In_654);
nor U251 (N_251,In_690,In_188);
nor U252 (N_252,In_1052,In_517);
nand U253 (N_253,In_732,In_760);
nand U254 (N_254,In_1121,In_191);
nor U255 (N_255,In_1471,In_568);
or U256 (N_256,In_609,In_1183);
xor U257 (N_257,In_152,In_971);
nor U258 (N_258,In_1406,In_648);
xor U259 (N_259,In_357,In_1054);
and U260 (N_260,In_1485,In_658);
nand U261 (N_261,In_700,In_543);
nor U262 (N_262,In_6,In_598);
and U263 (N_263,In_935,In_81);
or U264 (N_264,In_409,In_989);
nand U265 (N_265,In_817,In_768);
and U266 (N_266,In_1142,In_1030);
xor U267 (N_267,In_289,In_322);
xnor U268 (N_268,In_807,In_987);
nor U269 (N_269,In_1490,In_585);
or U270 (N_270,In_549,In_603);
nor U271 (N_271,In_140,In_834);
and U272 (N_272,In_321,In_349);
and U273 (N_273,In_403,In_1497);
and U274 (N_274,In_1131,In_116);
xor U275 (N_275,In_55,In_1031);
nor U276 (N_276,In_401,In_342);
and U277 (N_277,In_175,In_960);
or U278 (N_278,In_814,In_1155);
and U279 (N_279,In_793,In_941);
nor U280 (N_280,In_1425,In_329);
and U281 (N_281,In_337,In_954);
or U282 (N_282,In_228,In_385);
nand U283 (N_283,In_466,In_1289);
and U284 (N_284,In_542,In_1323);
and U285 (N_285,In_796,In_139);
and U286 (N_286,In_1409,In_254);
nor U287 (N_287,In_467,In_605);
nand U288 (N_288,In_1320,In_249);
or U289 (N_289,In_720,In_1137);
and U290 (N_290,In_1396,In_1018);
nand U291 (N_291,In_1400,In_1382);
nor U292 (N_292,In_1154,In_1388);
nand U293 (N_293,In_120,In_1322);
or U294 (N_294,In_765,In_900);
or U295 (N_295,In_299,In_1014);
or U296 (N_296,In_273,In_734);
or U297 (N_297,In_1001,In_1376);
or U298 (N_298,In_1007,In_348);
nor U299 (N_299,In_1085,In_490);
nand U300 (N_300,In_1276,In_502);
nand U301 (N_301,In_22,In_964);
and U302 (N_302,In_40,In_1128);
nor U303 (N_303,In_1306,In_60);
and U304 (N_304,In_930,In_390);
nor U305 (N_305,In_1056,In_1081);
or U306 (N_306,In_858,In_1365);
and U307 (N_307,In_1236,In_24);
nor U308 (N_308,In_728,In_163);
nor U309 (N_309,In_619,In_53);
nand U310 (N_310,In_87,In_1168);
and U311 (N_311,In_752,In_1414);
and U312 (N_312,In_742,In_892);
or U313 (N_313,In_1241,In_1398);
nor U314 (N_314,In_1073,In_618);
and U315 (N_315,In_622,In_560);
and U316 (N_316,In_826,In_118);
nor U317 (N_317,In_865,In_1201);
and U318 (N_318,In_1392,In_1210);
nand U319 (N_319,In_841,In_430);
and U320 (N_320,In_359,In_1307);
nor U321 (N_321,In_800,In_1273);
nor U322 (N_322,In_197,In_896);
or U323 (N_323,In_1368,In_128);
and U324 (N_324,In_35,In_1337);
nand U325 (N_325,In_1431,In_156);
nor U326 (N_326,In_940,In_363);
xor U327 (N_327,In_835,In_1163);
nor U328 (N_328,In_323,In_454);
and U329 (N_329,In_532,In_1024);
and U330 (N_330,In_34,In_205);
nor U331 (N_331,In_432,In_223);
nand U332 (N_332,In_966,In_1068);
nor U333 (N_333,In_998,In_633);
or U334 (N_334,In_4,In_50);
xor U335 (N_335,In_1443,In_680);
nand U336 (N_336,In_341,In_1220);
and U337 (N_337,In_1002,In_747);
nand U338 (N_338,In_608,In_1493);
and U339 (N_339,In_1035,In_1363);
or U340 (N_340,In_73,In_1397);
nor U341 (N_341,In_644,In_1378);
nand U342 (N_342,In_525,In_672);
nand U343 (N_343,In_1100,In_220);
xor U344 (N_344,In_157,In_227);
and U345 (N_345,In_1413,In_891);
nand U346 (N_346,In_240,In_507);
and U347 (N_347,In_999,In_576);
or U348 (N_348,In_851,In_1453);
and U349 (N_349,In_31,In_200);
nand U350 (N_350,In_778,In_544);
and U351 (N_351,In_1407,In_1332);
or U352 (N_352,In_414,In_763);
and U353 (N_353,In_821,In_1188);
nor U354 (N_354,In_736,In_584);
or U355 (N_355,In_263,In_1268);
nand U356 (N_356,In_1311,In_627);
and U357 (N_357,In_843,In_1223);
nor U358 (N_358,In_149,In_153);
nor U359 (N_359,In_624,In_101);
nor U360 (N_360,In_32,In_513);
xnor U361 (N_361,In_1249,In_172);
and U362 (N_362,In_1094,In_567);
xor U363 (N_363,In_279,In_897);
nor U364 (N_364,In_1027,In_257);
nor U365 (N_365,In_753,In_1304);
xnor U366 (N_366,In_494,In_1233);
nor U367 (N_367,In_889,In_1370);
or U368 (N_368,In_369,In_224);
and U369 (N_369,In_539,In_271);
or U370 (N_370,In_440,In_248);
nand U371 (N_371,In_1299,In_992);
nor U372 (N_372,In_1101,In_822);
nand U373 (N_373,In_39,In_862);
and U374 (N_374,In_417,In_267);
nor U375 (N_375,In_255,In_571);
nand U376 (N_376,In_137,In_1491);
nor U377 (N_377,In_985,In_506);
nand U378 (N_378,In_1041,In_599);
and U379 (N_379,In_57,In_708);
and U380 (N_380,In_1296,In_947);
and U381 (N_381,In_1159,In_474);
and U382 (N_382,In_1278,In_867);
nand U383 (N_383,In_1245,In_1102);
nand U384 (N_384,In_148,In_58);
nor U385 (N_385,In_739,In_413);
and U386 (N_386,In_350,In_1204);
or U387 (N_387,In_687,In_918);
nand U388 (N_388,In_1088,In_743);
and U389 (N_389,In_167,In_434);
or U390 (N_390,In_1375,In_199);
and U391 (N_391,In_1173,In_685);
nor U392 (N_392,In_872,In_482);
or U393 (N_393,In_902,In_51);
nor U394 (N_394,In_136,In_554);
nor U395 (N_395,In_703,In_469);
or U396 (N_396,In_487,In_287);
or U397 (N_397,In_1022,In_186);
or U398 (N_398,In_1360,In_1302);
nand U399 (N_399,In_551,In_613);
and U400 (N_400,In_586,In_738);
and U401 (N_401,In_1487,In_1093);
and U402 (N_402,In_1333,In_1476);
nand U403 (N_403,In_225,In_1248);
nor U404 (N_404,In_215,In_1499);
and U405 (N_405,In_485,In_247);
or U406 (N_406,In_1118,In_1112);
nand U407 (N_407,In_411,In_1412);
nand U408 (N_408,In_1239,In_790);
xor U409 (N_409,In_85,In_1373);
nand U410 (N_410,In_1120,In_997);
or U411 (N_411,In_1246,In_491);
nand U412 (N_412,In_1399,In_281);
nor U413 (N_413,In_1446,In_1228);
and U414 (N_414,In_561,In_590);
nand U415 (N_415,In_510,In_354);
nor U416 (N_416,In_917,In_1186);
or U417 (N_417,In_206,In_493);
nand U418 (N_418,In_1048,In_1442);
or U419 (N_419,In_671,In_786);
nand U420 (N_420,In_592,In_266);
and U421 (N_421,In_419,In_1357);
or U422 (N_422,In_79,In_1232);
nand U423 (N_423,In_1040,In_1091);
xnor U424 (N_424,In_580,In_694);
nand U425 (N_425,In_803,In_707);
or U426 (N_426,In_252,In_785);
nand U427 (N_427,In_30,In_1341);
and U428 (N_428,In_1458,In_300);
nand U429 (N_429,In_1023,In_1390);
nand U430 (N_430,In_1217,In_901);
nor U431 (N_431,In_392,In_1277);
nor U432 (N_432,In_1104,In_1275);
nand U433 (N_433,In_330,In_569);
nor U434 (N_434,In_219,In_614);
nand U435 (N_435,In_1192,In_878);
xnor U436 (N_436,In_1064,In_424);
and U437 (N_437,In_28,In_1464);
nor U438 (N_438,In_833,In_438);
nor U439 (N_439,In_939,In_518);
or U440 (N_440,In_1313,In_1350);
and U441 (N_441,In_682,In_1362);
xor U442 (N_442,In_473,In_159);
xor U443 (N_443,In_1385,In_958);
nor U444 (N_444,In_488,In_1290);
or U445 (N_445,In_218,In_113);
nand U446 (N_446,In_234,In_604);
and U447 (N_447,In_425,In_546);
nor U448 (N_448,In_1139,In_1033);
xor U449 (N_449,In_238,In_938);
and U450 (N_450,In_959,In_1281);
and U451 (N_451,In_797,In_67);
and U452 (N_452,In_365,In_725);
and U453 (N_453,In_784,In_919);
and U454 (N_454,In_213,In_84);
nand U455 (N_455,In_1303,In_1288);
xnor U456 (N_456,In_1433,In_177);
and U457 (N_457,In_1369,In_689);
nor U458 (N_458,In_472,In_435);
and U459 (N_459,In_393,In_1178);
nor U460 (N_460,In_1348,In_634);
nor U461 (N_461,In_1404,In_83);
xnor U462 (N_462,In_190,In_82);
and U463 (N_463,In_973,In_1152);
or U464 (N_464,In_1330,In_714);
nor U465 (N_465,In_597,In_655);
nor U466 (N_466,In_1342,In_636);
nor U467 (N_467,In_235,In_1004);
or U468 (N_468,In_913,In_426);
or U469 (N_469,In_1355,In_1187);
nor U470 (N_470,In_132,In_384);
or U471 (N_471,In_1045,In_1448);
nand U472 (N_472,In_91,In_1280);
nor U473 (N_473,In_358,In_1200);
or U474 (N_474,In_886,In_1050);
nor U475 (N_475,In_1381,In_150);
nor U476 (N_476,In_812,In_849);
or U477 (N_477,In_351,In_38);
and U478 (N_478,In_740,In_916);
nand U479 (N_479,In_1270,In_1230);
and U480 (N_480,In_457,In_119);
or U481 (N_481,In_1189,In_537);
nor U482 (N_482,In_1250,In_41);
and U483 (N_483,In_664,In_1195);
nor U484 (N_484,In_678,In_1202);
or U485 (N_485,In_399,In_169);
or U486 (N_486,In_852,In_102);
nand U487 (N_487,In_1046,In_866);
or U488 (N_488,In_381,In_236);
nand U489 (N_489,In_174,In_1271);
nor U490 (N_490,In_1107,In_589);
nand U491 (N_491,In_1457,In_368);
or U492 (N_492,In_335,In_1028);
or U493 (N_493,In_679,In_565);
nand U494 (N_494,In_1125,In_1080);
and U495 (N_495,In_364,In_1070);
nor U496 (N_496,In_652,In_563);
nand U497 (N_497,In_1126,In_343);
and U498 (N_498,In_379,In_1198);
nor U499 (N_499,In_986,In_1117);
and U500 (N_500,In_77,In_558);
nand U501 (N_501,In_129,In_929);
xnor U502 (N_502,In_667,In_853);
nand U503 (N_503,In_840,In_1145);
or U504 (N_504,In_1207,In_983);
and U505 (N_505,In_1005,In_1419);
nor U506 (N_506,In_904,In_1426);
and U507 (N_507,In_572,In_1261);
or U508 (N_508,In_123,In_1096);
nor U509 (N_509,In_759,In_861);
nand U510 (N_510,In_915,In_1253);
nor U511 (N_511,In_404,In_1380);
nor U512 (N_512,In_911,In_388);
or U513 (N_513,In_320,In_920);
nor U514 (N_514,In_1410,In_459);
or U515 (N_515,In_162,In_161);
nor U516 (N_516,In_479,In_1447);
and U517 (N_517,In_1467,In_1429);
nand U518 (N_518,In_1465,In_907);
nor U519 (N_519,In_270,In_1424);
xnor U520 (N_520,In_0,In_675);
or U521 (N_521,In_1205,In_751);
or U522 (N_522,In_1394,In_1000);
or U523 (N_523,In_702,In_54);
or U524 (N_524,In_868,In_1215);
nand U525 (N_525,In_1484,In_721);
nor U526 (N_526,In_59,In_550);
or U527 (N_527,In_274,In_1075);
or U528 (N_528,In_1042,In_90);
nor U529 (N_529,In_836,In_557);
and U530 (N_530,In_909,In_303);
nand U531 (N_531,In_863,In_845);
or U532 (N_532,In_697,In_143);
and U533 (N_533,In_651,In_306);
or U534 (N_534,In_312,In_1254);
nor U535 (N_535,In_421,In_698);
or U536 (N_536,In_1265,In_522);
and U537 (N_537,In_583,In_423);
or U538 (N_538,In_352,In_1116);
and U539 (N_539,In_23,In_1130);
nand U540 (N_540,In_207,In_1300);
nand U541 (N_541,In_80,In_448);
or U542 (N_542,In_857,In_64);
and U543 (N_543,In_121,In_944);
and U544 (N_544,In_955,In_1460);
xnor U545 (N_545,In_514,In_1122);
nor U546 (N_546,In_284,In_446);
or U547 (N_547,In_75,In_239);
nor U548 (N_548,In_429,In_570);
nor U549 (N_549,In_1032,In_336);
nand U550 (N_550,In_511,In_1282);
or U551 (N_551,In_71,In_1074);
nor U552 (N_552,In_1021,In_1498);
and U553 (N_553,In_1161,In_1461);
and U554 (N_554,In_1272,In_1439);
nand U555 (N_555,In_86,In_1352);
nor U556 (N_556,In_1483,In_1286);
nor U557 (N_557,In_462,In_1034);
and U558 (N_558,In_722,In_258);
and U559 (N_559,In_1110,In_716);
nor U560 (N_560,In_625,In_111);
nand U561 (N_561,In_1262,In_61);
nand U562 (N_562,In_497,In_662);
nor U563 (N_563,In_292,In_854);
nor U564 (N_564,In_730,In_291);
nor U565 (N_565,In_1076,In_642);
or U566 (N_566,In_820,In_78);
or U567 (N_567,In_165,In_838);
or U568 (N_568,In_719,In_353);
or U569 (N_569,In_647,In_356);
or U570 (N_570,In_277,In_495);
nor U571 (N_571,In_783,In_1482);
nand U572 (N_572,In_187,In_873);
or U573 (N_573,In_626,In_308);
nor U574 (N_574,In_1162,In_105);
and U575 (N_575,In_540,In_810);
or U576 (N_576,In_1430,In_374);
nor U577 (N_577,In_1010,In_976);
nor U578 (N_578,In_977,In_1235);
xor U579 (N_579,In_880,In_1175);
nor U580 (N_580,In_11,In_757);
nand U581 (N_581,In_748,In_282);
nand U582 (N_582,In_1459,In_1301);
or U583 (N_583,In_623,In_415);
or U584 (N_584,In_160,In_926);
nand U585 (N_585,In_717,In_315);
or U586 (N_586,In_387,In_1455);
nor U587 (N_587,In_775,In_575);
and U588 (N_588,In_278,In_1221);
and U589 (N_589,In_1344,In_1053);
and U590 (N_590,In_1124,In_1206);
and U591 (N_591,In_383,In_166);
nand U592 (N_592,In_1488,In_46);
and U593 (N_593,In_63,In_789);
nor U594 (N_594,In_692,In_304);
or U595 (N_595,In_185,In_290);
nand U596 (N_596,In_638,In_1452);
and U597 (N_597,In_107,In_1019);
xnor U598 (N_598,In_1319,In_1295);
and U599 (N_599,In_1260,In_340);
nor U600 (N_600,In_1462,In_402);
nand U601 (N_601,In_1364,In_394);
nand U602 (N_602,In_1072,In_1418);
nand U603 (N_603,In_481,In_731);
and U604 (N_604,In_1138,In_1237);
nor U605 (N_605,In_44,In_1143);
nand U606 (N_606,In_1267,In_397);
or U607 (N_607,In_666,In_1119);
or U608 (N_608,In_712,In_928);
or U609 (N_609,In_1312,In_276);
nand U610 (N_610,In_1449,In_222);
nor U611 (N_611,In_806,In_135);
nand U612 (N_612,In_181,In_460);
nand U613 (N_613,In_1321,In_914);
or U614 (N_614,In_972,In_683);
or U615 (N_615,In_637,In_791);
and U616 (N_616,In_553,In_980);
and U617 (N_617,In_1269,In_674);
nand U618 (N_618,In_1061,In_600);
or U619 (N_619,In_237,In_313);
nand U620 (N_620,In_766,In_1481);
xor U621 (N_621,In_456,In_217);
nand U622 (N_622,In_179,In_975);
and U623 (N_623,In_260,In_361);
xor U624 (N_624,In_1158,In_114);
and U625 (N_625,In_1222,In_451);
xor U626 (N_626,In_94,In_829);
xor U627 (N_627,In_310,In_996);
xor U628 (N_628,In_1274,In_194);
or U629 (N_629,In_777,In_1292);
and U630 (N_630,In_211,In_1283);
or U631 (N_631,In_180,In_1317);
nand U632 (N_632,In_1255,In_527);
nand U633 (N_633,In_881,In_1315);
nor U634 (N_634,In_3,In_898);
and U635 (N_635,In_1421,In_677);
nor U636 (N_636,In_602,In_818);
and U637 (N_637,In_318,In_33);
or U638 (N_638,In_37,In_126);
nand U639 (N_639,In_839,In_1169);
nand U640 (N_640,In_640,In_552);
nand U641 (N_641,In_1097,In_574);
or U642 (N_642,In_14,In_309);
xor U643 (N_643,In_792,In_903);
nand U644 (N_644,In_663,In_1456);
xor U645 (N_645,In_1335,In_957);
and U646 (N_646,In_212,In_713);
xnor U647 (N_647,In_1489,In_893);
and U648 (N_648,In_788,In_298);
xnor U649 (N_649,In_461,In_874);
nor U650 (N_650,In_1196,In_798);
nor U651 (N_651,In_164,In_1213);
nor U652 (N_652,In_88,In_99);
xnor U653 (N_653,In_832,In_990);
and U654 (N_654,In_994,In_936);
xor U655 (N_655,In_1012,In_993);
and U656 (N_656,In_825,In_1063);
and U657 (N_657,In_1240,In_1037);
nor U658 (N_658,In_870,In_937);
and U659 (N_659,In_17,In_499);
nor U660 (N_660,In_856,In_695);
nand U661 (N_661,In_1294,In_253);
nand U662 (N_662,In_52,In_1477);
or U663 (N_663,In_943,In_476);
nor U664 (N_664,In_95,In_631);
nor U665 (N_665,In_1371,In_1349);
or U666 (N_666,In_645,In_366);
nand U667 (N_667,In_1445,In_811);
and U668 (N_668,In_621,In_1327);
xor U669 (N_669,In_158,In_764);
and U670 (N_670,In_416,In_1440);
or U671 (N_671,In_1174,In_1067);
nor U672 (N_672,In_1318,In_1238);
nor U673 (N_673,In_596,In_968);
or U674 (N_674,In_981,In_1109);
nand U675 (N_675,In_612,In_1098);
and U676 (N_676,In_441,In_428);
or U677 (N_677,In_265,In_1258);
and U678 (N_678,In_1469,In_545);
nand U679 (N_679,In_1402,In_509);
nor U680 (N_680,In_1374,In_946);
xor U681 (N_681,In_173,In_942);
or U682 (N_682,In_1403,In_908);
or U683 (N_683,In_555,In_500);
nand U684 (N_684,In_530,In_508);
nor U685 (N_685,In_56,In_1141);
xnor U686 (N_686,In_98,In_659);
and U687 (N_687,In_701,In_452);
nand U688 (N_688,In_610,In_47);
and U689 (N_689,In_433,In_745);
or U690 (N_690,In_520,In_601);
and U691 (N_691,In_230,In_293);
and U692 (N_692,In_801,In_1361);
nor U693 (N_693,In_620,In_1441);
and U694 (N_694,In_1060,In_1172);
or U695 (N_695,In_1417,In_594);
or U696 (N_696,In_170,In_632);
nand U697 (N_697,In_750,In_1181);
nor U698 (N_698,In_498,In_1383);
nor U699 (N_699,In_606,In_1336);
nor U700 (N_700,In_1115,In_189);
nor U701 (N_701,In_1191,In_295);
or U702 (N_702,In_178,In_670);
nand U703 (N_703,In_1293,In_673);
nor U704 (N_704,In_927,In_1386);
xor U705 (N_705,In_978,In_1347);
nor U706 (N_706,In_1334,In_405);
nor U707 (N_707,In_1015,In_183);
or U708 (N_708,In_1479,In_616);
nand U709 (N_709,In_70,In_184);
and U710 (N_710,In_1087,In_1194);
xnor U711 (N_711,In_1208,In_578);
nor U712 (N_712,In_650,In_1065);
and U713 (N_713,In_117,In_538);
xnor U714 (N_714,In_106,In_1351);
nor U715 (N_715,In_1328,In_1416);
or U716 (N_716,In_124,In_1480);
and U717 (N_717,In_406,In_951);
nand U718 (N_718,In_74,In_630);
nor U719 (N_719,In_1494,In_808);
nor U720 (N_720,In_923,In_326);
nor U721 (N_721,In_802,In_1197);
nor U722 (N_722,In_422,In_1051);
nand U723 (N_723,In_1316,In_883);
nand U724 (N_724,In_66,In_10);
and U725 (N_725,In_1136,In_528);
nand U726 (N_726,In_72,In_548);
nand U727 (N_727,In_1432,In_1147);
xor U728 (N_728,In_1135,In_952);
nand U729 (N_729,In_727,In_1180);
and U730 (N_730,In_635,In_65);
nor U731 (N_731,In_21,In_1287);
or U732 (N_732,In_233,In_1423);
nand U733 (N_733,In_108,In_556);
nor U734 (N_734,In_210,In_1451);
and U735 (N_735,In_314,In_860);
nand U736 (N_736,In_979,In_1049);
nand U737 (N_737,In_362,In_380);
or U738 (N_738,In_963,In_1343);
nand U739 (N_739,In_1305,In_1013);
nand U740 (N_740,In_1170,In_1153);
nor U741 (N_741,In_848,In_657);
and U742 (N_742,In_1071,In_1150);
and U743 (N_743,In_869,In_729);
or U744 (N_744,In_564,In_533);
and U745 (N_745,In_1329,In_130);
nor U746 (N_746,In_984,In_216);
or U747 (N_747,In_1039,In_925);
nand U748 (N_748,In_138,In_324);
or U749 (N_749,In_1234,In_69);
nor U750 (N_750,N_358,N_69);
or U751 (N_751,N_373,N_510);
nor U752 (N_752,N_53,N_726);
nor U753 (N_753,N_57,N_423);
or U754 (N_754,N_678,N_507);
xnor U755 (N_755,N_17,N_707);
nor U756 (N_756,N_715,N_741);
nand U757 (N_757,N_431,N_309);
or U758 (N_758,N_696,N_52);
nor U759 (N_759,N_213,N_483);
nor U760 (N_760,N_607,N_180);
or U761 (N_761,N_603,N_2);
nand U762 (N_762,N_391,N_545);
nor U763 (N_763,N_725,N_746);
nor U764 (N_764,N_37,N_645);
nand U765 (N_765,N_666,N_230);
or U766 (N_766,N_305,N_64);
nand U767 (N_767,N_129,N_196);
or U768 (N_768,N_118,N_271);
xnor U769 (N_769,N_125,N_106);
nand U770 (N_770,N_269,N_415);
nor U771 (N_771,N_341,N_235);
or U772 (N_772,N_455,N_380);
nor U773 (N_773,N_504,N_31);
nand U774 (N_774,N_495,N_291);
or U775 (N_775,N_332,N_710);
nand U776 (N_776,N_225,N_281);
nand U777 (N_777,N_200,N_685);
nor U778 (N_778,N_40,N_62);
nor U779 (N_779,N_246,N_314);
nand U780 (N_780,N_708,N_290);
or U781 (N_781,N_232,N_537);
nand U782 (N_782,N_739,N_534);
nor U783 (N_783,N_1,N_387);
nor U784 (N_784,N_335,N_458);
nand U785 (N_785,N_193,N_647);
xnor U786 (N_786,N_326,N_721);
nor U787 (N_787,N_593,N_469);
xnor U788 (N_788,N_153,N_498);
nand U789 (N_789,N_299,N_158);
nand U790 (N_790,N_195,N_462);
and U791 (N_791,N_749,N_82);
and U792 (N_792,N_83,N_352);
or U793 (N_793,N_508,N_436);
and U794 (N_794,N_591,N_437);
and U795 (N_795,N_240,N_533);
nor U796 (N_796,N_347,N_527);
and U797 (N_797,N_698,N_744);
or U798 (N_798,N_171,N_25);
xor U799 (N_799,N_105,N_124);
nand U800 (N_800,N_137,N_688);
and U801 (N_801,N_419,N_306);
nor U802 (N_802,N_218,N_632);
nor U803 (N_803,N_544,N_134);
and U804 (N_804,N_207,N_642);
nand U805 (N_805,N_18,N_11);
nor U806 (N_806,N_536,N_747);
or U807 (N_807,N_107,N_98);
or U808 (N_808,N_110,N_610);
and U809 (N_809,N_452,N_425);
nor U810 (N_810,N_327,N_297);
and U811 (N_811,N_717,N_737);
nor U812 (N_812,N_531,N_432);
xor U813 (N_813,N_628,N_587);
nand U814 (N_814,N_517,N_165);
nand U815 (N_815,N_637,N_712);
nor U816 (N_816,N_101,N_569);
nor U817 (N_817,N_461,N_427);
xnor U818 (N_818,N_679,N_173);
and U819 (N_819,N_417,N_585);
and U820 (N_820,N_266,N_443);
and U821 (N_821,N_278,N_264);
nand U822 (N_822,N_621,N_261);
nand U823 (N_823,N_476,N_449);
and U824 (N_824,N_192,N_377);
nor U825 (N_825,N_93,N_234);
nand U826 (N_826,N_694,N_275);
and U827 (N_827,N_71,N_668);
nand U828 (N_828,N_651,N_304);
nand U829 (N_829,N_548,N_280);
and U830 (N_830,N_86,N_238);
nor U831 (N_831,N_518,N_4);
and U832 (N_832,N_185,N_252);
and U833 (N_833,N_372,N_606);
nor U834 (N_834,N_114,N_614);
or U835 (N_835,N_677,N_657);
nand U836 (N_836,N_35,N_95);
nor U837 (N_837,N_487,N_7);
nor U838 (N_838,N_374,N_549);
or U839 (N_839,N_72,N_10);
nor U840 (N_840,N_295,N_638);
or U841 (N_841,N_426,N_402);
nand U842 (N_842,N_223,N_538);
nand U843 (N_843,N_430,N_486);
xor U844 (N_844,N_499,N_579);
nand U845 (N_845,N_478,N_220);
nor U846 (N_846,N_468,N_568);
nor U847 (N_847,N_90,N_67);
or U848 (N_848,N_515,N_578);
xor U849 (N_849,N_338,N_100);
and U850 (N_850,N_308,N_683);
and U851 (N_851,N_144,N_420);
xor U852 (N_852,N_321,N_277);
nor U853 (N_853,N_539,N_214);
nor U854 (N_854,N_520,N_355);
nor U855 (N_855,N_599,N_547);
and U856 (N_856,N_215,N_732);
xor U857 (N_857,N_346,N_369);
nor U858 (N_858,N_244,N_169);
nand U859 (N_859,N_328,N_640);
nand U860 (N_860,N_617,N_655);
and U861 (N_861,N_160,N_514);
nor U862 (N_862,N_401,N_345);
or U863 (N_863,N_550,N_320);
or U864 (N_864,N_582,N_0);
or U865 (N_865,N_600,N_413);
nand U866 (N_866,N_245,N_51);
and U867 (N_867,N_279,N_263);
or U868 (N_868,N_382,N_87);
nor U869 (N_869,N_644,N_650);
nor U870 (N_870,N_674,N_664);
and U871 (N_871,N_485,N_268);
or U872 (N_872,N_285,N_604);
nand U873 (N_873,N_396,N_294);
nand U874 (N_874,N_697,N_581);
xnor U875 (N_875,N_699,N_8);
nor U876 (N_876,N_130,N_172);
or U877 (N_877,N_13,N_360);
and U878 (N_878,N_170,N_388);
nand U879 (N_879,N_745,N_466);
nand U880 (N_880,N_557,N_331);
or U881 (N_881,N_284,N_108);
xnor U882 (N_882,N_247,N_140);
or U883 (N_883,N_625,N_639);
or U884 (N_884,N_505,N_113);
and U885 (N_885,N_684,N_14);
or U886 (N_886,N_257,N_590);
nor U887 (N_887,N_602,N_734);
nand U888 (N_888,N_342,N_555);
nor U889 (N_889,N_561,N_733);
and U890 (N_890,N_571,N_411);
or U891 (N_891,N_633,N_143);
nand U892 (N_892,N_509,N_330);
and U893 (N_893,N_334,N_404);
nand U894 (N_894,N_724,N_667);
nor U895 (N_895,N_283,N_670);
and U896 (N_896,N_339,N_700);
and U897 (N_897,N_258,N_528);
and U898 (N_898,N_233,N_151);
and U899 (N_899,N_65,N_94);
xnor U900 (N_900,N_723,N_139);
and U901 (N_901,N_325,N_318);
nor U902 (N_902,N_611,N_484);
and U903 (N_903,N_46,N_208);
nor U904 (N_904,N_618,N_109);
nor U905 (N_905,N_652,N_322);
nand U906 (N_906,N_671,N_177);
nand U907 (N_907,N_378,N_159);
and U908 (N_908,N_658,N_711);
or U909 (N_909,N_410,N_634);
and U910 (N_910,N_78,N_577);
and U911 (N_911,N_622,N_643);
or U912 (N_912,N_502,N_75);
nor U913 (N_913,N_259,N_526);
nor U914 (N_914,N_722,N_97);
nand U915 (N_915,N_164,N_435);
nor U916 (N_916,N_654,N_190);
and U917 (N_917,N_237,N_201);
nand U918 (N_918,N_250,N_738);
nand U919 (N_919,N_481,N_359);
nor U920 (N_920,N_79,N_641);
nor U921 (N_921,N_61,N_501);
nor U922 (N_922,N_28,N_84);
nand U923 (N_923,N_400,N_273);
xor U924 (N_924,N_563,N_523);
nor U925 (N_925,N_748,N_687);
and U926 (N_926,N_442,N_301);
nor U927 (N_927,N_150,N_68);
nand U928 (N_928,N_660,N_624);
nand U929 (N_929,N_690,N_669);
and U930 (N_930,N_102,N_530);
or U931 (N_931,N_421,N_231);
or U932 (N_932,N_274,N_370);
nor U933 (N_933,N_228,N_197);
and U934 (N_934,N_50,N_613);
nand U935 (N_935,N_511,N_15);
xor U936 (N_936,N_80,N_399);
and U937 (N_937,N_210,N_112);
nor U938 (N_938,N_189,N_99);
or U939 (N_939,N_663,N_479);
xor U940 (N_940,N_146,N_96);
nand U941 (N_941,N_390,N_619);
nor U942 (N_942,N_543,N_574);
or U943 (N_943,N_298,N_540);
nor U944 (N_944,N_16,N_88);
or U945 (N_945,N_608,N_253);
xor U946 (N_946,N_519,N_312);
nand U947 (N_947,N_313,N_251);
or U948 (N_948,N_116,N_541);
nor U949 (N_949,N_292,N_248);
and U950 (N_950,N_262,N_605);
nand U951 (N_951,N_542,N_76);
and U952 (N_952,N_293,N_546);
nand U953 (N_953,N_242,N_727);
nor U954 (N_954,N_202,N_365);
and U955 (N_955,N_21,N_414);
nand U956 (N_956,N_123,N_428);
or U957 (N_957,N_142,N_296);
nor U958 (N_958,N_438,N_77);
or U959 (N_959,N_389,N_282);
and U960 (N_960,N_203,N_492);
nor U961 (N_961,N_205,N_467);
nor U962 (N_962,N_128,N_363);
or U963 (N_963,N_592,N_300);
nor U964 (N_964,N_597,N_615);
or U965 (N_965,N_513,N_454);
or U966 (N_966,N_357,N_323);
xor U967 (N_967,N_392,N_703);
or U968 (N_968,N_553,N_556);
nand U969 (N_969,N_728,N_635);
or U970 (N_970,N_89,N_315);
nand U971 (N_971,N_23,N_673);
nor U972 (N_972,N_333,N_403);
nand U973 (N_973,N_488,N_424);
or U974 (N_974,N_731,N_41);
nand U975 (N_975,N_176,N_475);
and U976 (N_976,N_489,N_702);
or U977 (N_977,N_630,N_494);
nand U978 (N_978,N_395,N_39);
nor U979 (N_979,N_450,N_689);
and U980 (N_980,N_629,N_111);
nor U981 (N_981,N_126,N_434);
nor U982 (N_982,N_535,N_224);
nor U983 (N_983,N_719,N_446);
nor U984 (N_984,N_609,N_740);
or U985 (N_985,N_705,N_70);
and U986 (N_986,N_47,N_310);
nand U987 (N_987,N_38,N_376);
nor U988 (N_988,N_287,N_525);
or U989 (N_989,N_364,N_122);
nor U990 (N_990,N_152,N_30);
nand U991 (N_991,N_289,N_366);
or U992 (N_992,N_672,N_565);
or U993 (N_993,N_361,N_337);
and U994 (N_994,N_302,N_646);
xnor U995 (N_995,N_706,N_583);
nor U996 (N_996,N_42,N_612);
nor U997 (N_997,N_491,N_272);
nor U998 (N_998,N_255,N_162);
or U999 (N_999,N_596,N_49);
or U1000 (N_1000,N_463,N_206);
nand U1001 (N_1001,N_60,N_456);
nand U1002 (N_1002,N_408,N_429);
or U1003 (N_1003,N_36,N_586);
nor U1004 (N_1004,N_324,N_209);
and U1005 (N_1005,N_691,N_58);
or U1006 (N_1006,N_656,N_490);
or U1007 (N_1007,N_659,N_199);
or U1008 (N_1008,N_26,N_63);
and U1009 (N_1009,N_136,N_343);
nor U1010 (N_1010,N_66,N_249);
nor U1011 (N_1011,N_626,N_623);
and U1012 (N_1012,N_393,N_127);
nand U1013 (N_1013,N_496,N_551);
or U1014 (N_1014,N_665,N_117);
or U1015 (N_1015,N_163,N_5);
nand U1016 (N_1016,N_336,N_219);
nand U1017 (N_1017,N_270,N_120);
nor U1018 (N_1018,N_473,N_155);
nor U1019 (N_1019,N_9,N_529);
and U1020 (N_1020,N_179,N_472);
or U1021 (N_1021,N_211,N_131);
xnor U1022 (N_1022,N_188,N_340);
or U1023 (N_1023,N_85,N_516);
xnor U1024 (N_1024,N_662,N_121);
xor U1025 (N_1025,N_24,N_439);
xor U1026 (N_1026,N_464,N_319);
nor U1027 (N_1027,N_221,N_477);
and U1028 (N_1028,N_572,N_701);
or U1029 (N_1029,N_497,N_156);
nor U1030 (N_1030,N_718,N_383);
and U1031 (N_1031,N_138,N_92);
xnor U1032 (N_1032,N_133,N_704);
or U1033 (N_1033,N_132,N_676);
nor U1034 (N_1034,N_405,N_56);
nand U1035 (N_1035,N_103,N_43);
and U1036 (N_1036,N_181,N_521);
and U1037 (N_1037,N_742,N_186);
nor U1038 (N_1038,N_34,N_441);
xnor U1039 (N_1039,N_115,N_191);
or U1040 (N_1040,N_198,N_329);
and U1041 (N_1041,N_141,N_695);
nand U1042 (N_1042,N_522,N_661);
and U1043 (N_1043,N_350,N_54);
nor U1044 (N_1044,N_567,N_500);
and U1045 (N_1045,N_532,N_166);
or U1046 (N_1046,N_381,N_12);
xor U1047 (N_1047,N_344,N_386);
xnor U1048 (N_1048,N_560,N_709);
or U1049 (N_1049,N_184,N_174);
or U1050 (N_1050,N_594,N_375);
nor U1051 (N_1051,N_575,N_471);
nor U1052 (N_1052,N_559,N_736);
and U1053 (N_1053,N_147,N_554);
nor U1054 (N_1054,N_265,N_19);
or U1055 (N_1055,N_433,N_368);
and U1056 (N_1056,N_354,N_407);
and U1057 (N_1057,N_459,N_187);
nor U1058 (N_1058,N_227,N_562);
nand U1059 (N_1059,N_254,N_448);
or U1060 (N_1060,N_743,N_267);
nor U1061 (N_1061,N_573,N_73);
and U1062 (N_1062,N_44,N_620);
nor U1063 (N_1063,N_470,N_493);
or U1064 (N_1064,N_589,N_91);
or U1065 (N_1065,N_648,N_474);
nand U1066 (N_1066,N_385,N_311);
nand U1067 (N_1067,N_482,N_348);
nand U1068 (N_1068,N_167,N_81);
xnor U1069 (N_1069,N_27,N_730);
and U1070 (N_1070,N_182,N_353);
xor U1071 (N_1071,N_276,N_409);
xor U1072 (N_1072,N_217,N_226);
nand U1073 (N_1073,N_681,N_45);
nand U1074 (N_1074,N_22,N_584);
nand U1075 (N_1075,N_349,N_627);
nand U1076 (N_1076,N_154,N_692);
and U1077 (N_1077,N_3,N_351);
nand U1078 (N_1078,N_6,N_713);
nor U1079 (N_1079,N_570,N_33);
nand U1080 (N_1080,N_564,N_241);
and U1081 (N_1081,N_576,N_236);
nand U1082 (N_1082,N_149,N_601);
nor U1083 (N_1083,N_29,N_457);
nor U1084 (N_1084,N_356,N_451);
and U1085 (N_1085,N_379,N_616);
xor U1086 (N_1086,N_183,N_720);
and U1087 (N_1087,N_631,N_714);
nand U1088 (N_1088,N_222,N_675);
and U1089 (N_1089,N_288,N_686);
xor U1090 (N_1090,N_636,N_367);
or U1091 (N_1091,N_371,N_422);
or U1092 (N_1092,N_444,N_453);
and U1093 (N_1093,N_48,N_416);
or U1094 (N_1094,N_212,N_119);
and U1095 (N_1095,N_394,N_588);
or U1096 (N_1096,N_161,N_460);
nor U1097 (N_1097,N_384,N_145);
and U1098 (N_1098,N_558,N_104);
xor U1099 (N_1099,N_307,N_682);
nand U1100 (N_1100,N_303,N_316);
or U1101 (N_1101,N_397,N_447);
or U1102 (N_1102,N_735,N_229);
xnor U1103 (N_1103,N_503,N_566);
xnor U1104 (N_1104,N_680,N_512);
nor U1105 (N_1105,N_418,N_243);
and U1106 (N_1106,N_729,N_178);
nor U1107 (N_1107,N_524,N_406);
nand U1108 (N_1108,N_239,N_362);
or U1109 (N_1109,N_204,N_412);
xnor U1110 (N_1110,N_175,N_693);
and U1111 (N_1111,N_168,N_440);
nand U1112 (N_1112,N_260,N_598);
nor U1113 (N_1113,N_398,N_506);
or U1114 (N_1114,N_552,N_317);
and U1115 (N_1115,N_256,N_74);
nand U1116 (N_1116,N_216,N_649);
nor U1117 (N_1117,N_653,N_716);
nor U1118 (N_1118,N_32,N_55);
xnor U1119 (N_1119,N_580,N_480);
nor U1120 (N_1120,N_135,N_286);
nor U1121 (N_1121,N_148,N_194);
nand U1122 (N_1122,N_59,N_465);
nor U1123 (N_1123,N_445,N_157);
xor U1124 (N_1124,N_595,N_20);
nor U1125 (N_1125,N_574,N_674);
or U1126 (N_1126,N_311,N_283);
or U1127 (N_1127,N_645,N_474);
xnor U1128 (N_1128,N_711,N_675);
or U1129 (N_1129,N_255,N_28);
nor U1130 (N_1130,N_147,N_342);
xnor U1131 (N_1131,N_370,N_586);
nor U1132 (N_1132,N_408,N_197);
or U1133 (N_1133,N_733,N_627);
and U1134 (N_1134,N_558,N_214);
nand U1135 (N_1135,N_34,N_629);
nor U1136 (N_1136,N_557,N_178);
nand U1137 (N_1137,N_325,N_287);
nand U1138 (N_1138,N_235,N_32);
and U1139 (N_1139,N_674,N_157);
xor U1140 (N_1140,N_620,N_196);
and U1141 (N_1141,N_35,N_5);
nor U1142 (N_1142,N_577,N_635);
or U1143 (N_1143,N_342,N_302);
and U1144 (N_1144,N_201,N_346);
or U1145 (N_1145,N_75,N_309);
nor U1146 (N_1146,N_163,N_318);
and U1147 (N_1147,N_656,N_209);
xnor U1148 (N_1148,N_447,N_17);
and U1149 (N_1149,N_586,N_439);
nand U1150 (N_1150,N_211,N_338);
and U1151 (N_1151,N_660,N_171);
and U1152 (N_1152,N_411,N_517);
nor U1153 (N_1153,N_373,N_155);
nand U1154 (N_1154,N_608,N_331);
nor U1155 (N_1155,N_255,N_490);
nand U1156 (N_1156,N_358,N_599);
and U1157 (N_1157,N_5,N_734);
xnor U1158 (N_1158,N_199,N_684);
or U1159 (N_1159,N_148,N_189);
nand U1160 (N_1160,N_102,N_605);
and U1161 (N_1161,N_104,N_369);
nand U1162 (N_1162,N_160,N_597);
and U1163 (N_1163,N_41,N_210);
and U1164 (N_1164,N_485,N_124);
and U1165 (N_1165,N_512,N_497);
nor U1166 (N_1166,N_59,N_591);
or U1167 (N_1167,N_307,N_630);
nand U1168 (N_1168,N_284,N_151);
nand U1169 (N_1169,N_3,N_532);
and U1170 (N_1170,N_125,N_511);
and U1171 (N_1171,N_588,N_264);
nor U1172 (N_1172,N_357,N_40);
or U1173 (N_1173,N_453,N_537);
nand U1174 (N_1174,N_394,N_329);
and U1175 (N_1175,N_245,N_635);
and U1176 (N_1176,N_484,N_137);
or U1177 (N_1177,N_246,N_639);
nor U1178 (N_1178,N_659,N_324);
nor U1179 (N_1179,N_514,N_582);
nand U1180 (N_1180,N_361,N_339);
or U1181 (N_1181,N_402,N_328);
or U1182 (N_1182,N_596,N_355);
and U1183 (N_1183,N_489,N_530);
xor U1184 (N_1184,N_200,N_228);
nand U1185 (N_1185,N_79,N_104);
or U1186 (N_1186,N_520,N_336);
and U1187 (N_1187,N_372,N_184);
and U1188 (N_1188,N_707,N_384);
or U1189 (N_1189,N_731,N_76);
nand U1190 (N_1190,N_104,N_292);
xor U1191 (N_1191,N_365,N_412);
xnor U1192 (N_1192,N_686,N_263);
or U1193 (N_1193,N_377,N_177);
or U1194 (N_1194,N_54,N_192);
xnor U1195 (N_1195,N_593,N_648);
or U1196 (N_1196,N_575,N_352);
nor U1197 (N_1197,N_543,N_218);
xnor U1198 (N_1198,N_117,N_132);
or U1199 (N_1199,N_259,N_380);
and U1200 (N_1200,N_237,N_711);
nand U1201 (N_1201,N_185,N_102);
nor U1202 (N_1202,N_467,N_674);
or U1203 (N_1203,N_471,N_243);
nor U1204 (N_1204,N_549,N_345);
xor U1205 (N_1205,N_425,N_247);
nor U1206 (N_1206,N_471,N_218);
nand U1207 (N_1207,N_131,N_627);
and U1208 (N_1208,N_106,N_649);
nor U1209 (N_1209,N_41,N_488);
and U1210 (N_1210,N_556,N_746);
nor U1211 (N_1211,N_25,N_197);
nor U1212 (N_1212,N_264,N_162);
nor U1213 (N_1213,N_342,N_0);
or U1214 (N_1214,N_533,N_747);
nand U1215 (N_1215,N_368,N_576);
nor U1216 (N_1216,N_426,N_25);
nand U1217 (N_1217,N_65,N_658);
or U1218 (N_1218,N_58,N_38);
or U1219 (N_1219,N_177,N_475);
nor U1220 (N_1220,N_297,N_658);
and U1221 (N_1221,N_130,N_150);
or U1222 (N_1222,N_150,N_345);
nor U1223 (N_1223,N_126,N_114);
nand U1224 (N_1224,N_364,N_22);
nor U1225 (N_1225,N_318,N_587);
or U1226 (N_1226,N_390,N_194);
or U1227 (N_1227,N_124,N_112);
or U1228 (N_1228,N_198,N_6);
and U1229 (N_1229,N_363,N_125);
xor U1230 (N_1230,N_317,N_70);
and U1231 (N_1231,N_307,N_532);
nand U1232 (N_1232,N_319,N_337);
nand U1233 (N_1233,N_74,N_539);
nor U1234 (N_1234,N_172,N_473);
nor U1235 (N_1235,N_60,N_573);
or U1236 (N_1236,N_695,N_147);
and U1237 (N_1237,N_25,N_442);
xor U1238 (N_1238,N_417,N_479);
nand U1239 (N_1239,N_679,N_523);
and U1240 (N_1240,N_698,N_706);
nand U1241 (N_1241,N_381,N_79);
or U1242 (N_1242,N_213,N_34);
and U1243 (N_1243,N_690,N_358);
nor U1244 (N_1244,N_671,N_679);
and U1245 (N_1245,N_39,N_59);
xor U1246 (N_1246,N_513,N_501);
xnor U1247 (N_1247,N_105,N_246);
and U1248 (N_1248,N_691,N_617);
nor U1249 (N_1249,N_621,N_536);
nor U1250 (N_1250,N_519,N_464);
nand U1251 (N_1251,N_53,N_20);
nand U1252 (N_1252,N_287,N_591);
nand U1253 (N_1253,N_249,N_748);
nand U1254 (N_1254,N_41,N_355);
or U1255 (N_1255,N_388,N_198);
nor U1256 (N_1256,N_170,N_272);
or U1257 (N_1257,N_702,N_607);
nand U1258 (N_1258,N_497,N_712);
or U1259 (N_1259,N_207,N_414);
nand U1260 (N_1260,N_60,N_280);
or U1261 (N_1261,N_376,N_81);
and U1262 (N_1262,N_441,N_529);
xnor U1263 (N_1263,N_362,N_485);
xnor U1264 (N_1264,N_293,N_679);
nor U1265 (N_1265,N_102,N_54);
and U1266 (N_1266,N_542,N_163);
xnor U1267 (N_1267,N_519,N_654);
nor U1268 (N_1268,N_158,N_70);
nand U1269 (N_1269,N_721,N_463);
xnor U1270 (N_1270,N_367,N_70);
or U1271 (N_1271,N_466,N_427);
and U1272 (N_1272,N_371,N_500);
nor U1273 (N_1273,N_646,N_341);
and U1274 (N_1274,N_372,N_365);
or U1275 (N_1275,N_87,N_155);
nor U1276 (N_1276,N_74,N_317);
nand U1277 (N_1277,N_663,N_229);
xor U1278 (N_1278,N_576,N_57);
and U1279 (N_1279,N_101,N_345);
and U1280 (N_1280,N_338,N_124);
nand U1281 (N_1281,N_601,N_221);
or U1282 (N_1282,N_548,N_138);
nor U1283 (N_1283,N_25,N_318);
or U1284 (N_1284,N_143,N_565);
nor U1285 (N_1285,N_196,N_71);
nand U1286 (N_1286,N_540,N_361);
nor U1287 (N_1287,N_66,N_311);
and U1288 (N_1288,N_411,N_499);
nor U1289 (N_1289,N_477,N_331);
nor U1290 (N_1290,N_341,N_673);
nand U1291 (N_1291,N_174,N_226);
xnor U1292 (N_1292,N_460,N_301);
nor U1293 (N_1293,N_38,N_89);
and U1294 (N_1294,N_653,N_15);
nand U1295 (N_1295,N_251,N_301);
and U1296 (N_1296,N_553,N_475);
nand U1297 (N_1297,N_719,N_112);
nor U1298 (N_1298,N_3,N_25);
and U1299 (N_1299,N_495,N_625);
nand U1300 (N_1300,N_223,N_18);
xor U1301 (N_1301,N_734,N_33);
and U1302 (N_1302,N_306,N_388);
or U1303 (N_1303,N_700,N_547);
and U1304 (N_1304,N_353,N_227);
or U1305 (N_1305,N_30,N_28);
xor U1306 (N_1306,N_26,N_519);
and U1307 (N_1307,N_488,N_515);
or U1308 (N_1308,N_612,N_702);
and U1309 (N_1309,N_427,N_167);
or U1310 (N_1310,N_369,N_459);
nor U1311 (N_1311,N_681,N_536);
or U1312 (N_1312,N_26,N_559);
nand U1313 (N_1313,N_26,N_435);
nand U1314 (N_1314,N_480,N_510);
and U1315 (N_1315,N_617,N_160);
or U1316 (N_1316,N_41,N_614);
or U1317 (N_1317,N_625,N_478);
nor U1318 (N_1318,N_130,N_330);
xnor U1319 (N_1319,N_586,N_92);
nand U1320 (N_1320,N_45,N_197);
and U1321 (N_1321,N_738,N_498);
xnor U1322 (N_1322,N_69,N_0);
nand U1323 (N_1323,N_739,N_721);
nor U1324 (N_1324,N_362,N_222);
nor U1325 (N_1325,N_251,N_131);
nand U1326 (N_1326,N_12,N_302);
or U1327 (N_1327,N_684,N_413);
nand U1328 (N_1328,N_2,N_55);
and U1329 (N_1329,N_283,N_220);
nor U1330 (N_1330,N_36,N_706);
nor U1331 (N_1331,N_640,N_461);
nand U1332 (N_1332,N_94,N_117);
xor U1333 (N_1333,N_625,N_637);
and U1334 (N_1334,N_243,N_477);
nand U1335 (N_1335,N_635,N_637);
or U1336 (N_1336,N_375,N_122);
or U1337 (N_1337,N_98,N_413);
and U1338 (N_1338,N_739,N_418);
nand U1339 (N_1339,N_204,N_721);
nand U1340 (N_1340,N_475,N_29);
or U1341 (N_1341,N_371,N_88);
nor U1342 (N_1342,N_105,N_421);
nor U1343 (N_1343,N_217,N_70);
and U1344 (N_1344,N_25,N_373);
and U1345 (N_1345,N_399,N_239);
xnor U1346 (N_1346,N_700,N_182);
and U1347 (N_1347,N_625,N_605);
nor U1348 (N_1348,N_57,N_609);
nand U1349 (N_1349,N_462,N_111);
and U1350 (N_1350,N_502,N_303);
nor U1351 (N_1351,N_480,N_562);
and U1352 (N_1352,N_497,N_440);
nand U1353 (N_1353,N_563,N_63);
and U1354 (N_1354,N_66,N_297);
and U1355 (N_1355,N_337,N_363);
and U1356 (N_1356,N_212,N_67);
nor U1357 (N_1357,N_632,N_26);
xnor U1358 (N_1358,N_531,N_220);
and U1359 (N_1359,N_536,N_88);
and U1360 (N_1360,N_122,N_272);
nand U1361 (N_1361,N_120,N_138);
and U1362 (N_1362,N_20,N_178);
nor U1363 (N_1363,N_748,N_98);
nor U1364 (N_1364,N_375,N_608);
xor U1365 (N_1365,N_444,N_142);
xnor U1366 (N_1366,N_106,N_553);
nand U1367 (N_1367,N_533,N_103);
nand U1368 (N_1368,N_78,N_85);
nand U1369 (N_1369,N_563,N_555);
or U1370 (N_1370,N_57,N_643);
and U1371 (N_1371,N_177,N_324);
xor U1372 (N_1372,N_215,N_609);
nor U1373 (N_1373,N_679,N_394);
nand U1374 (N_1374,N_701,N_746);
xnor U1375 (N_1375,N_52,N_210);
nand U1376 (N_1376,N_635,N_467);
and U1377 (N_1377,N_45,N_362);
nor U1378 (N_1378,N_143,N_168);
nand U1379 (N_1379,N_604,N_26);
nand U1380 (N_1380,N_432,N_93);
or U1381 (N_1381,N_523,N_657);
nor U1382 (N_1382,N_147,N_129);
or U1383 (N_1383,N_402,N_271);
nor U1384 (N_1384,N_730,N_43);
or U1385 (N_1385,N_694,N_436);
and U1386 (N_1386,N_203,N_220);
nor U1387 (N_1387,N_456,N_516);
or U1388 (N_1388,N_692,N_265);
nor U1389 (N_1389,N_294,N_28);
or U1390 (N_1390,N_156,N_222);
nor U1391 (N_1391,N_393,N_551);
nor U1392 (N_1392,N_722,N_147);
or U1393 (N_1393,N_176,N_665);
nor U1394 (N_1394,N_517,N_340);
nor U1395 (N_1395,N_715,N_652);
and U1396 (N_1396,N_656,N_147);
xor U1397 (N_1397,N_304,N_503);
or U1398 (N_1398,N_510,N_372);
nor U1399 (N_1399,N_688,N_124);
or U1400 (N_1400,N_377,N_369);
nand U1401 (N_1401,N_309,N_587);
nand U1402 (N_1402,N_490,N_632);
nor U1403 (N_1403,N_613,N_434);
or U1404 (N_1404,N_173,N_74);
nand U1405 (N_1405,N_597,N_197);
and U1406 (N_1406,N_462,N_62);
nor U1407 (N_1407,N_675,N_741);
or U1408 (N_1408,N_63,N_496);
or U1409 (N_1409,N_349,N_241);
nor U1410 (N_1410,N_368,N_371);
nand U1411 (N_1411,N_90,N_272);
nand U1412 (N_1412,N_86,N_671);
or U1413 (N_1413,N_365,N_197);
and U1414 (N_1414,N_166,N_316);
and U1415 (N_1415,N_320,N_55);
or U1416 (N_1416,N_233,N_95);
or U1417 (N_1417,N_147,N_387);
nand U1418 (N_1418,N_124,N_360);
and U1419 (N_1419,N_186,N_279);
and U1420 (N_1420,N_268,N_244);
nand U1421 (N_1421,N_144,N_83);
or U1422 (N_1422,N_135,N_67);
nor U1423 (N_1423,N_533,N_145);
xnor U1424 (N_1424,N_337,N_712);
and U1425 (N_1425,N_705,N_593);
xnor U1426 (N_1426,N_609,N_70);
nand U1427 (N_1427,N_433,N_0);
and U1428 (N_1428,N_518,N_576);
and U1429 (N_1429,N_28,N_206);
or U1430 (N_1430,N_301,N_231);
xor U1431 (N_1431,N_641,N_85);
nand U1432 (N_1432,N_103,N_316);
nand U1433 (N_1433,N_175,N_440);
or U1434 (N_1434,N_696,N_498);
xor U1435 (N_1435,N_70,N_18);
or U1436 (N_1436,N_671,N_478);
nor U1437 (N_1437,N_669,N_611);
nand U1438 (N_1438,N_111,N_245);
nand U1439 (N_1439,N_462,N_607);
xnor U1440 (N_1440,N_57,N_38);
or U1441 (N_1441,N_387,N_363);
or U1442 (N_1442,N_403,N_258);
xor U1443 (N_1443,N_669,N_412);
and U1444 (N_1444,N_347,N_686);
and U1445 (N_1445,N_729,N_702);
nand U1446 (N_1446,N_115,N_229);
nor U1447 (N_1447,N_65,N_121);
nor U1448 (N_1448,N_504,N_524);
or U1449 (N_1449,N_540,N_68);
and U1450 (N_1450,N_733,N_665);
and U1451 (N_1451,N_646,N_21);
or U1452 (N_1452,N_36,N_499);
nor U1453 (N_1453,N_275,N_558);
xor U1454 (N_1454,N_344,N_84);
nand U1455 (N_1455,N_182,N_397);
nor U1456 (N_1456,N_543,N_410);
or U1457 (N_1457,N_692,N_10);
nand U1458 (N_1458,N_74,N_357);
nand U1459 (N_1459,N_586,N_220);
xor U1460 (N_1460,N_587,N_70);
nor U1461 (N_1461,N_585,N_37);
and U1462 (N_1462,N_409,N_82);
and U1463 (N_1463,N_700,N_383);
nor U1464 (N_1464,N_151,N_395);
nor U1465 (N_1465,N_719,N_15);
or U1466 (N_1466,N_109,N_384);
or U1467 (N_1467,N_498,N_185);
and U1468 (N_1468,N_497,N_230);
and U1469 (N_1469,N_447,N_576);
or U1470 (N_1470,N_201,N_647);
xnor U1471 (N_1471,N_70,N_618);
nand U1472 (N_1472,N_121,N_96);
nand U1473 (N_1473,N_324,N_267);
xnor U1474 (N_1474,N_52,N_409);
nand U1475 (N_1475,N_42,N_228);
or U1476 (N_1476,N_438,N_111);
nor U1477 (N_1477,N_469,N_638);
or U1478 (N_1478,N_266,N_542);
and U1479 (N_1479,N_298,N_362);
or U1480 (N_1480,N_13,N_14);
nor U1481 (N_1481,N_715,N_77);
nand U1482 (N_1482,N_687,N_741);
and U1483 (N_1483,N_602,N_267);
nand U1484 (N_1484,N_586,N_734);
xnor U1485 (N_1485,N_480,N_165);
nor U1486 (N_1486,N_194,N_622);
and U1487 (N_1487,N_169,N_66);
nand U1488 (N_1488,N_571,N_612);
or U1489 (N_1489,N_686,N_683);
or U1490 (N_1490,N_2,N_168);
and U1491 (N_1491,N_372,N_261);
nor U1492 (N_1492,N_739,N_414);
nand U1493 (N_1493,N_434,N_661);
nor U1494 (N_1494,N_105,N_736);
nor U1495 (N_1495,N_93,N_128);
nand U1496 (N_1496,N_684,N_342);
or U1497 (N_1497,N_615,N_694);
nand U1498 (N_1498,N_129,N_394);
and U1499 (N_1499,N_8,N_673);
or U1500 (N_1500,N_1439,N_830);
nor U1501 (N_1501,N_868,N_926);
and U1502 (N_1502,N_873,N_1031);
nor U1503 (N_1503,N_1260,N_1460);
nand U1504 (N_1504,N_1087,N_1166);
or U1505 (N_1505,N_1187,N_1106);
nand U1506 (N_1506,N_810,N_1458);
nor U1507 (N_1507,N_787,N_1186);
nor U1508 (N_1508,N_1143,N_1228);
or U1509 (N_1509,N_1403,N_1318);
nor U1510 (N_1510,N_1153,N_1459);
xor U1511 (N_1511,N_1138,N_1116);
or U1512 (N_1512,N_1225,N_932);
or U1513 (N_1513,N_760,N_1472);
nand U1514 (N_1514,N_1486,N_1267);
nand U1515 (N_1515,N_1250,N_900);
nand U1516 (N_1516,N_755,N_1303);
nor U1517 (N_1517,N_1088,N_961);
and U1518 (N_1518,N_1397,N_1466);
and U1519 (N_1519,N_1162,N_1082);
and U1520 (N_1520,N_1379,N_965);
nand U1521 (N_1521,N_1323,N_1229);
nor U1522 (N_1522,N_1305,N_1287);
nor U1523 (N_1523,N_903,N_892);
nand U1524 (N_1524,N_1060,N_1333);
nor U1525 (N_1525,N_1265,N_1469);
and U1526 (N_1526,N_1112,N_1360);
nand U1527 (N_1527,N_1230,N_1408);
nand U1528 (N_1528,N_1154,N_1314);
nand U1529 (N_1529,N_1051,N_941);
xor U1530 (N_1530,N_1426,N_1131);
or U1531 (N_1531,N_1382,N_1477);
and U1532 (N_1532,N_778,N_1139);
or U1533 (N_1533,N_969,N_769);
nor U1534 (N_1534,N_834,N_988);
nand U1535 (N_1535,N_981,N_1484);
and U1536 (N_1536,N_762,N_1342);
nand U1537 (N_1537,N_1272,N_1163);
nand U1538 (N_1538,N_1384,N_1084);
nand U1539 (N_1539,N_1404,N_1134);
nand U1540 (N_1540,N_1320,N_783);
nor U1541 (N_1541,N_823,N_962);
nand U1542 (N_1542,N_831,N_915);
nor U1543 (N_1543,N_1057,N_1115);
and U1544 (N_1544,N_1209,N_1053);
and U1545 (N_1545,N_1217,N_816);
and U1546 (N_1546,N_1223,N_750);
nor U1547 (N_1547,N_1428,N_880);
and U1548 (N_1548,N_1247,N_1105);
nand U1549 (N_1549,N_1158,N_780);
or U1550 (N_1550,N_1074,N_770);
xor U1551 (N_1551,N_1117,N_1252);
and U1552 (N_1552,N_1062,N_1038);
xor U1553 (N_1553,N_1133,N_1189);
and U1554 (N_1554,N_849,N_824);
nor U1555 (N_1555,N_773,N_1248);
or U1556 (N_1556,N_1385,N_772);
nand U1557 (N_1557,N_906,N_832);
xnor U1558 (N_1558,N_1351,N_1000);
or U1559 (N_1559,N_1177,N_1258);
xor U1560 (N_1560,N_1419,N_1004);
nor U1561 (N_1561,N_1465,N_1441);
xnor U1562 (N_1562,N_1483,N_1013);
nand U1563 (N_1563,N_1271,N_1437);
nand U1564 (N_1564,N_1043,N_874);
nor U1565 (N_1565,N_1201,N_842);
or U1566 (N_1566,N_1224,N_1291);
nor U1567 (N_1567,N_1262,N_1492);
nor U1568 (N_1568,N_1415,N_1330);
or U1569 (N_1569,N_1001,N_1079);
xor U1570 (N_1570,N_1251,N_1067);
nand U1571 (N_1571,N_1028,N_1244);
nor U1572 (N_1572,N_1147,N_947);
nor U1573 (N_1573,N_923,N_1290);
nand U1574 (N_1574,N_756,N_1180);
nand U1575 (N_1575,N_1340,N_837);
nor U1576 (N_1576,N_982,N_1041);
or U1577 (N_1577,N_1192,N_929);
xor U1578 (N_1578,N_1299,N_795);
xnor U1579 (N_1579,N_1207,N_1322);
nor U1580 (N_1580,N_945,N_1071);
xnor U1581 (N_1581,N_1246,N_1034);
nand U1582 (N_1582,N_1433,N_939);
nand U1583 (N_1583,N_1480,N_885);
nand U1584 (N_1584,N_958,N_784);
or U1585 (N_1585,N_1242,N_1197);
or U1586 (N_1586,N_1454,N_1396);
or U1587 (N_1587,N_803,N_1016);
nand U1588 (N_1588,N_1080,N_1003);
and U1589 (N_1589,N_1279,N_1239);
nand U1590 (N_1590,N_897,N_835);
and U1591 (N_1591,N_1418,N_1304);
nor U1592 (N_1592,N_1378,N_853);
nand U1593 (N_1593,N_1359,N_952);
nor U1594 (N_1594,N_917,N_1414);
xnor U1595 (N_1595,N_1058,N_1107);
or U1596 (N_1596,N_771,N_1474);
nor U1597 (N_1597,N_1137,N_951);
nor U1598 (N_1598,N_893,N_1381);
xnor U1599 (N_1599,N_1461,N_1072);
nor U1600 (N_1600,N_1365,N_1331);
nor U1601 (N_1601,N_1344,N_1311);
and U1602 (N_1602,N_1356,N_1215);
nand U1603 (N_1603,N_1475,N_1049);
nor U1604 (N_1604,N_1407,N_1297);
nor U1605 (N_1605,N_1171,N_858);
nor U1606 (N_1606,N_1317,N_905);
and U1607 (N_1607,N_912,N_1152);
nor U1608 (N_1608,N_1453,N_1211);
and U1609 (N_1609,N_1094,N_799);
nand U1610 (N_1610,N_794,N_761);
nor U1611 (N_1611,N_825,N_840);
or U1612 (N_1612,N_1463,N_753);
nor U1613 (N_1613,N_1448,N_983);
or U1614 (N_1614,N_909,N_847);
or U1615 (N_1615,N_1349,N_992);
and U1616 (N_1616,N_828,N_973);
nor U1617 (N_1617,N_1431,N_1256);
nor U1618 (N_1618,N_970,N_817);
xnor U1619 (N_1619,N_1298,N_883);
or U1620 (N_1620,N_1017,N_1345);
nand U1621 (N_1621,N_1245,N_1417);
nor U1622 (N_1622,N_766,N_844);
xor U1623 (N_1623,N_768,N_1392);
nor U1624 (N_1624,N_1122,N_953);
and U1625 (N_1625,N_888,N_1168);
and U1626 (N_1626,N_1410,N_919);
or U1627 (N_1627,N_1416,N_1097);
nor U1628 (N_1628,N_1178,N_1312);
and U1629 (N_1629,N_1190,N_1332);
nand U1630 (N_1630,N_1024,N_852);
xnor U1631 (N_1631,N_980,N_896);
or U1632 (N_1632,N_1198,N_754);
xor U1633 (N_1633,N_1146,N_751);
nand U1634 (N_1634,N_845,N_894);
nor U1635 (N_1635,N_1046,N_1165);
xor U1636 (N_1636,N_1435,N_757);
nand U1637 (N_1637,N_1169,N_963);
nand U1638 (N_1638,N_1464,N_959);
nand U1639 (N_1639,N_1481,N_934);
nand U1640 (N_1640,N_1170,N_829);
nor U1641 (N_1641,N_1490,N_1130);
or U1642 (N_1642,N_856,N_937);
nand U1643 (N_1643,N_938,N_918);
nand U1644 (N_1644,N_910,N_1042);
nand U1645 (N_1645,N_1307,N_1184);
or U1646 (N_1646,N_1204,N_1280);
or U1647 (N_1647,N_857,N_1011);
nand U1648 (N_1648,N_879,N_1363);
nor U1649 (N_1649,N_819,N_1026);
nor U1650 (N_1650,N_1226,N_1039);
nand U1651 (N_1651,N_1175,N_989);
nand U1652 (N_1652,N_1052,N_1061);
nor U1653 (N_1653,N_1123,N_1015);
and U1654 (N_1654,N_1372,N_1019);
xor U1655 (N_1655,N_1254,N_1425);
or U1656 (N_1656,N_1487,N_1455);
and U1657 (N_1657,N_911,N_821);
or U1658 (N_1658,N_1236,N_1427);
nor U1659 (N_1659,N_1276,N_1327);
nor U1660 (N_1660,N_1086,N_978);
nand U1661 (N_1661,N_1350,N_1257);
nand U1662 (N_1662,N_793,N_996);
or U1663 (N_1663,N_1232,N_1253);
xor U1664 (N_1664,N_1411,N_1293);
nand U1665 (N_1665,N_935,N_836);
nor U1666 (N_1666,N_1341,N_1387);
xor U1667 (N_1667,N_1235,N_1354);
nand U1668 (N_1668,N_1282,N_1367);
and U1669 (N_1669,N_1366,N_833);
and U1670 (N_1670,N_1181,N_848);
and U1671 (N_1671,N_1399,N_1119);
xor U1672 (N_1672,N_1489,N_1240);
or U1673 (N_1673,N_1266,N_1195);
or U1674 (N_1674,N_1092,N_1135);
nand U1675 (N_1675,N_1284,N_998);
xor U1676 (N_1676,N_1149,N_1361);
and U1677 (N_1677,N_878,N_1335);
nor U1678 (N_1678,N_1479,N_1182);
nand U1679 (N_1679,N_813,N_1205);
or U1680 (N_1680,N_1144,N_1259);
or U1681 (N_1681,N_1012,N_1148);
and U1682 (N_1682,N_927,N_1173);
and U1683 (N_1683,N_1120,N_820);
nand U1684 (N_1684,N_1096,N_1334);
nand U1685 (N_1685,N_1233,N_1386);
or U1686 (N_1686,N_1045,N_1025);
nand U1687 (N_1687,N_1352,N_1377);
nand U1688 (N_1688,N_1347,N_1406);
xor U1689 (N_1689,N_1400,N_1243);
nor U1690 (N_1690,N_920,N_1485);
xnor U1691 (N_1691,N_826,N_1179);
or U1692 (N_1692,N_1413,N_801);
and U1693 (N_1693,N_1110,N_954);
or U1694 (N_1694,N_854,N_1468);
and U1695 (N_1695,N_1109,N_1277);
or U1696 (N_1696,N_944,N_765);
and U1697 (N_1697,N_811,N_1237);
nand U1698 (N_1698,N_987,N_1095);
xor U1699 (N_1699,N_1145,N_936);
and U1700 (N_1700,N_1032,N_1099);
nor U1701 (N_1701,N_1008,N_1346);
nand U1702 (N_1702,N_997,N_843);
and U1703 (N_1703,N_869,N_901);
nor U1704 (N_1704,N_1325,N_1036);
and U1705 (N_1705,N_881,N_1364);
and U1706 (N_1706,N_1362,N_884);
and U1707 (N_1707,N_955,N_1412);
nand U1708 (N_1708,N_1064,N_1129);
xnor U1709 (N_1709,N_1445,N_1430);
and U1710 (N_1710,N_890,N_964);
or U1711 (N_1711,N_863,N_798);
and U1712 (N_1712,N_1069,N_800);
or U1713 (N_1713,N_1338,N_1007);
or U1714 (N_1714,N_1376,N_1498);
or U1715 (N_1715,N_812,N_1313);
nor U1716 (N_1716,N_1124,N_1389);
nor U1717 (N_1717,N_994,N_1438);
nand U1718 (N_1718,N_1263,N_791);
and U1719 (N_1719,N_1421,N_1429);
and U1720 (N_1720,N_967,N_1050);
xor U1721 (N_1721,N_1222,N_792);
xnor U1722 (N_1722,N_1476,N_1188);
xnor U1723 (N_1723,N_1374,N_990);
and U1724 (N_1724,N_1261,N_1022);
and U1725 (N_1725,N_872,N_1447);
xor U1726 (N_1726,N_1108,N_1289);
nand U1727 (N_1727,N_976,N_1457);
nor U1728 (N_1728,N_1127,N_1373);
nor U1729 (N_1729,N_1035,N_786);
and U1730 (N_1730,N_1309,N_1434);
and U1731 (N_1731,N_1065,N_1176);
nand U1732 (N_1732,N_1398,N_1155);
or U1733 (N_1733,N_1370,N_1014);
nor U1734 (N_1734,N_1114,N_999);
nor U1735 (N_1735,N_1456,N_1212);
nand U1736 (N_1736,N_1185,N_1006);
nand U1737 (N_1737,N_889,N_1292);
or U1738 (N_1738,N_1059,N_1275);
nand U1739 (N_1739,N_986,N_928);
nor U1740 (N_1740,N_774,N_1315);
nor U1741 (N_1741,N_1473,N_1424);
or U1742 (N_1742,N_1055,N_943);
xor U1743 (N_1743,N_1339,N_1040);
and U1744 (N_1744,N_1090,N_1020);
and U1745 (N_1745,N_1118,N_1491);
nand U1746 (N_1746,N_822,N_1355);
nand U1747 (N_1747,N_763,N_1054);
nand U1748 (N_1748,N_887,N_1388);
and U1749 (N_1749,N_1156,N_809);
and U1750 (N_1750,N_942,N_946);
nor U1751 (N_1751,N_991,N_891);
xnor U1752 (N_1752,N_1393,N_1306);
and U1753 (N_1753,N_913,N_1196);
nand U1754 (N_1754,N_876,N_1241);
nor U1755 (N_1755,N_1467,N_1324);
nand U1756 (N_1756,N_1368,N_797);
xnor U1757 (N_1757,N_924,N_1023);
nor U1758 (N_1758,N_899,N_1283);
and U1759 (N_1759,N_1288,N_1113);
xor U1760 (N_1760,N_1078,N_1394);
xor U1761 (N_1761,N_972,N_1018);
xnor U1762 (N_1762,N_1450,N_1268);
or U1763 (N_1763,N_1076,N_850);
nand U1764 (N_1764,N_1140,N_1219);
nand U1765 (N_1765,N_968,N_1044);
or U1766 (N_1766,N_993,N_1183);
nand U1767 (N_1767,N_789,N_1160);
nand U1768 (N_1768,N_1255,N_1301);
xnor U1769 (N_1769,N_882,N_1056);
nor U1770 (N_1770,N_1103,N_1161);
nand U1771 (N_1771,N_1405,N_1295);
or U1772 (N_1772,N_1371,N_788);
nor U1773 (N_1773,N_1220,N_1005);
nand U1774 (N_1774,N_1157,N_1316);
or U1775 (N_1775,N_1081,N_1104);
nor U1776 (N_1776,N_1089,N_1077);
nor U1777 (N_1777,N_975,N_1422);
nor U1778 (N_1778,N_1375,N_1142);
nor U1779 (N_1779,N_1443,N_1030);
and U1780 (N_1780,N_1286,N_940);
and U1781 (N_1781,N_815,N_974);
nor U1782 (N_1782,N_950,N_1488);
or U1783 (N_1783,N_877,N_1213);
nor U1784 (N_1784,N_1451,N_971);
or U1785 (N_1785,N_1420,N_1029);
and U1786 (N_1786,N_1442,N_1302);
nand U1787 (N_1787,N_790,N_1497);
nor U1788 (N_1788,N_1264,N_1401);
nor U1789 (N_1789,N_1121,N_1021);
nor U1790 (N_1790,N_977,N_960);
or U1791 (N_1791,N_1048,N_1172);
nand U1792 (N_1792,N_1296,N_1310);
or U1793 (N_1793,N_1470,N_916);
nand U1794 (N_1794,N_805,N_1002);
and U1795 (N_1795,N_782,N_1478);
nand U1796 (N_1796,N_1353,N_851);
nand U1797 (N_1797,N_1343,N_838);
nand U1798 (N_1798,N_1100,N_1423);
nand U1799 (N_1799,N_1010,N_752);
or U1800 (N_1800,N_775,N_1126);
nor U1801 (N_1801,N_827,N_1174);
or U1802 (N_1802,N_1066,N_1319);
nor U1803 (N_1803,N_1449,N_1409);
and U1804 (N_1804,N_1070,N_907);
nor U1805 (N_1805,N_1369,N_839);
and U1806 (N_1806,N_1218,N_777);
and U1807 (N_1807,N_802,N_1326);
and U1808 (N_1808,N_1274,N_808);
nor U1809 (N_1809,N_1273,N_1164);
nor U1810 (N_1810,N_1037,N_1128);
nand U1811 (N_1811,N_1494,N_966);
nand U1812 (N_1812,N_1358,N_985);
nor U1813 (N_1813,N_1083,N_925);
or U1814 (N_1814,N_818,N_1321);
and U1815 (N_1815,N_1281,N_922);
nand U1816 (N_1816,N_1193,N_1111);
or U1817 (N_1817,N_957,N_949);
nand U1818 (N_1818,N_1191,N_865);
or U1819 (N_1819,N_1337,N_1101);
nand U1820 (N_1820,N_904,N_1194);
nand U1821 (N_1821,N_841,N_1125);
nor U1822 (N_1822,N_846,N_807);
nor U1823 (N_1823,N_1452,N_1440);
and U1824 (N_1824,N_1308,N_1210);
nand U1825 (N_1825,N_1380,N_1495);
nor U1826 (N_1826,N_933,N_1141);
xor U1827 (N_1827,N_804,N_1136);
or U1828 (N_1828,N_1269,N_796);
and U1829 (N_1829,N_1482,N_1159);
or U1830 (N_1830,N_1132,N_1329);
or U1831 (N_1831,N_1151,N_759);
and U1832 (N_1832,N_1063,N_931);
nand U1833 (N_1833,N_758,N_1278);
nor U1834 (N_1834,N_871,N_1216);
nor U1835 (N_1835,N_908,N_1249);
nand U1836 (N_1836,N_1471,N_1027);
and U1837 (N_1837,N_1395,N_1206);
and U1838 (N_1838,N_1383,N_1294);
nand U1839 (N_1839,N_948,N_886);
nand U1840 (N_1840,N_1200,N_1203);
xnor U1841 (N_1841,N_859,N_814);
nand U1842 (N_1842,N_776,N_995);
nor U1843 (N_1843,N_1234,N_902);
nand U1844 (N_1844,N_921,N_1091);
or U1845 (N_1845,N_1238,N_764);
nor U1846 (N_1846,N_1068,N_1432);
or U1847 (N_1847,N_867,N_1436);
or U1848 (N_1848,N_979,N_1009);
nand U1849 (N_1849,N_1231,N_1085);
nor U1850 (N_1850,N_861,N_875);
or U1851 (N_1851,N_1391,N_870);
and U1852 (N_1852,N_1227,N_1098);
and U1853 (N_1853,N_862,N_1499);
xnor U1854 (N_1854,N_1402,N_1270);
nor U1855 (N_1855,N_1150,N_956);
xnor U1856 (N_1856,N_1285,N_1462);
nor U1857 (N_1857,N_1493,N_1208);
nor U1858 (N_1858,N_1348,N_1496);
nor U1859 (N_1859,N_930,N_785);
nand U1860 (N_1860,N_1300,N_1328);
nor U1861 (N_1861,N_1075,N_866);
nand U1862 (N_1862,N_1357,N_1033);
xnor U1863 (N_1863,N_1221,N_1336);
nand U1864 (N_1864,N_1390,N_855);
xnor U1865 (N_1865,N_767,N_806);
nand U1866 (N_1866,N_1102,N_1073);
xnor U1867 (N_1867,N_1047,N_1167);
nor U1868 (N_1868,N_1199,N_895);
or U1869 (N_1869,N_1214,N_860);
or U1870 (N_1870,N_898,N_1446);
and U1871 (N_1871,N_779,N_914);
and U1872 (N_1872,N_1444,N_1202);
nor U1873 (N_1873,N_984,N_1093);
or U1874 (N_1874,N_864,N_781);
nor U1875 (N_1875,N_1192,N_836);
or U1876 (N_1876,N_1131,N_1412);
or U1877 (N_1877,N_814,N_1378);
nand U1878 (N_1878,N_1103,N_1305);
xnor U1879 (N_1879,N_1189,N_838);
nor U1880 (N_1880,N_1086,N_999);
nor U1881 (N_1881,N_1417,N_850);
nand U1882 (N_1882,N_1173,N_1040);
nand U1883 (N_1883,N_794,N_757);
nor U1884 (N_1884,N_1194,N_1454);
nor U1885 (N_1885,N_785,N_1281);
and U1886 (N_1886,N_921,N_887);
nor U1887 (N_1887,N_848,N_1465);
nor U1888 (N_1888,N_755,N_829);
nor U1889 (N_1889,N_1064,N_1427);
or U1890 (N_1890,N_1190,N_988);
and U1891 (N_1891,N_1245,N_1036);
or U1892 (N_1892,N_1194,N_1144);
or U1893 (N_1893,N_1138,N_978);
xor U1894 (N_1894,N_1215,N_1179);
nor U1895 (N_1895,N_982,N_977);
nand U1896 (N_1896,N_1085,N_830);
and U1897 (N_1897,N_1055,N_849);
nand U1898 (N_1898,N_1438,N_1454);
or U1899 (N_1899,N_780,N_1251);
nor U1900 (N_1900,N_1251,N_1315);
and U1901 (N_1901,N_792,N_1154);
nand U1902 (N_1902,N_833,N_1110);
and U1903 (N_1903,N_1067,N_932);
nand U1904 (N_1904,N_1149,N_838);
and U1905 (N_1905,N_1488,N_1023);
xor U1906 (N_1906,N_1069,N_1293);
xor U1907 (N_1907,N_1051,N_1318);
and U1908 (N_1908,N_959,N_1344);
nor U1909 (N_1909,N_1108,N_1009);
nand U1910 (N_1910,N_936,N_993);
and U1911 (N_1911,N_1278,N_1455);
nor U1912 (N_1912,N_821,N_816);
nand U1913 (N_1913,N_1239,N_1335);
or U1914 (N_1914,N_1220,N_990);
nand U1915 (N_1915,N_764,N_1263);
nor U1916 (N_1916,N_1245,N_1336);
and U1917 (N_1917,N_809,N_1282);
nand U1918 (N_1918,N_1465,N_1376);
or U1919 (N_1919,N_1481,N_1028);
nand U1920 (N_1920,N_1454,N_971);
or U1921 (N_1921,N_847,N_1282);
nor U1922 (N_1922,N_875,N_1291);
and U1923 (N_1923,N_1403,N_1094);
xnor U1924 (N_1924,N_1407,N_1306);
nand U1925 (N_1925,N_880,N_1390);
nand U1926 (N_1926,N_1083,N_1080);
or U1927 (N_1927,N_1061,N_1267);
nor U1928 (N_1928,N_1186,N_1313);
nor U1929 (N_1929,N_1458,N_1155);
or U1930 (N_1930,N_1371,N_883);
xor U1931 (N_1931,N_1004,N_1236);
and U1932 (N_1932,N_1054,N_758);
and U1933 (N_1933,N_977,N_890);
and U1934 (N_1934,N_854,N_1450);
and U1935 (N_1935,N_832,N_800);
xnor U1936 (N_1936,N_1210,N_1092);
or U1937 (N_1937,N_1311,N_1225);
nor U1938 (N_1938,N_1354,N_947);
nand U1939 (N_1939,N_838,N_940);
nor U1940 (N_1940,N_1460,N_1118);
or U1941 (N_1941,N_1016,N_786);
xnor U1942 (N_1942,N_971,N_1264);
or U1943 (N_1943,N_1334,N_780);
or U1944 (N_1944,N_1416,N_770);
nor U1945 (N_1945,N_793,N_1105);
nor U1946 (N_1946,N_970,N_877);
or U1947 (N_1947,N_1329,N_1181);
and U1948 (N_1948,N_1348,N_970);
nand U1949 (N_1949,N_918,N_907);
and U1950 (N_1950,N_761,N_914);
nor U1951 (N_1951,N_1355,N_1261);
or U1952 (N_1952,N_883,N_1160);
nand U1953 (N_1953,N_1266,N_1373);
nor U1954 (N_1954,N_1338,N_1174);
nand U1955 (N_1955,N_1453,N_1378);
nand U1956 (N_1956,N_1468,N_1096);
nor U1957 (N_1957,N_1218,N_1430);
and U1958 (N_1958,N_1010,N_1074);
nand U1959 (N_1959,N_914,N_795);
nor U1960 (N_1960,N_1093,N_847);
xnor U1961 (N_1961,N_947,N_1100);
and U1962 (N_1962,N_1313,N_1479);
nor U1963 (N_1963,N_1356,N_1481);
and U1964 (N_1964,N_1246,N_1270);
xor U1965 (N_1965,N_806,N_847);
xor U1966 (N_1966,N_806,N_901);
or U1967 (N_1967,N_1008,N_1005);
or U1968 (N_1968,N_959,N_801);
nand U1969 (N_1969,N_894,N_769);
or U1970 (N_1970,N_1388,N_1399);
and U1971 (N_1971,N_992,N_1173);
or U1972 (N_1972,N_1458,N_806);
nand U1973 (N_1973,N_1033,N_812);
and U1974 (N_1974,N_929,N_924);
nor U1975 (N_1975,N_1100,N_1378);
and U1976 (N_1976,N_1363,N_985);
nor U1977 (N_1977,N_985,N_925);
nor U1978 (N_1978,N_875,N_1176);
nor U1979 (N_1979,N_1149,N_1136);
nor U1980 (N_1980,N_932,N_1014);
nor U1981 (N_1981,N_1131,N_1166);
and U1982 (N_1982,N_821,N_1193);
nand U1983 (N_1983,N_1127,N_1384);
and U1984 (N_1984,N_859,N_1084);
xnor U1985 (N_1985,N_1153,N_776);
nand U1986 (N_1986,N_1416,N_924);
nor U1987 (N_1987,N_1375,N_945);
nand U1988 (N_1988,N_1073,N_951);
nor U1989 (N_1989,N_1077,N_919);
and U1990 (N_1990,N_920,N_975);
nor U1991 (N_1991,N_1463,N_1345);
and U1992 (N_1992,N_947,N_1327);
nor U1993 (N_1993,N_937,N_1032);
or U1994 (N_1994,N_1350,N_1129);
nand U1995 (N_1995,N_893,N_1033);
nand U1996 (N_1996,N_1193,N_1095);
nand U1997 (N_1997,N_1380,N_1195);
nand U1998 (N_1998,N_825,N_1392);
or U1999 (N_1999,N_918,N_1325);
and U2000 (N_2000,N_786,N_1165);
nor U2001 (N_2001,N_1304,N_1320);
or U2002 (N_2002,N_919,N_1209);
nor U2003 (N_2003,N_1281,N_1146);
nand U2004 (N_2004,N_1246,N_1349);
nor U2005 (N_2005,N_1443,N_1389);
and U2006 (N_2006,N_935,N_867);
nand U2007 (N_2007,N_1089,N_1136);
or U2008 (N_2008,N_944,N_1297);
or U2009 (N_2009,N_1326,N_1070);
nor U2010 (N_2010,N_1447,N_1414);
nor U2011 (N_2011,N_846,N_1014);
nor U2012 (N_2012,N_1191,N_1092);
nor U2013 (N_2013,N_1431,N_984);
or U2014 (N_2014,N_1289,N_1454);
xor U2015 (N_2015,N_832,N_949);
nor U2016 (N_2016,N_1026,N_1352);
and U2017 (N_2017,N_1404,N_831);
and U2018 (N_2018,N_1075,N_1330);
nor U2019 (N_2019,N_852,N_1413);
nor U2020 (N_2020,N_1194,N_962);
or U2021 (N_2021,N_1052,N_1246);
or U2022 (N_2022,N_1186,N_1317);
nor U2023 (N_2023,N_835,N_752);
and U2024 (N_2024,N_1490,N_867);
or U2025 (N_2025,N_1398,N_1272);
nand U2026 (N_2026,N_1081,N_1487);
xnor U2027 (N_2027,N_1171,N_1336);
or U2028 (N_2028,N_877,N_1301);
and U2029 (N_2029,N_1156,N_1211);
nand U2030 (N_2030,N_1214,N_964);
nor U2031 (N_2031,N_1195,N_910);
and U2032 (N_2032,N_1173,N_1168);
nor U2033 (N_2033,N_1219,N_1435);
nor U2034 (N_2034,N_1091,N_1414);
nor U2035 (N_2035,N_1430,N_1007);
nor U2036 (N_2036,N_948,N_1277);
nand U2037 (N_2037,N_834,N_1334);
or U2038 (N_2038,N_1214,N_1491);
nand U2039 (N_2039,N_1141,N_1279);
xnor U2040 (N_2040,N_1314,N_775);
or U2041 (N_2041,N_1251,N_911);
and U2042 (N_2042,N_1333,N_1264);
nand U2043 (N_2043,N_1438,N_1403);
or U2044 (N_2044,N_817,N_814);
and U2045 (N_2045,N_907,N_843);
nor U2046 (N_2046,N_763,N_837);
nor U2047 (N_2047,N_816,N_995);
or U2048 (N_2048,N_969,N_927);
and U2049 (N_2049,N_1484,N_1029);
nand U2050 (N_2050,N_1350,N_820);
nand U2051 (N_2051,N_764,N_1190);
or U2052 (N_2052,N_1012,N_996);
or U2053 (N_2053,N_1150,N_1013);
and U2054 (N_2054,N_843,N_937);
or U2055 (N_2055,N_1332,N_999);
nand U2056 (N_2056,N_1363,N_1134);
nor U2057 (N_2057,N_1409,N_1207);
nor U2058 (N_2058,N_1374,N_1070);
nor U2059 (N_2059,N_1486,N_1214);
nor U2060 (N_2060,N_762,N_838);
nand U2061 (N_2061,N_915,N_1361);
nor U2062 (N_2062,N_1454,N_1334);
nor U2063 (N_2063,N_1316,N_1353);
xnor U2064 (N_2064,N_1464,N_1324);
or U2065 (N_2065,N_1169,N_792);
nor U2066 (N_2066,N_871,N_1461);
and U2067 (N_2067,N_1317,N_823);
nand U2068 (N_2068,N_1303,N_1277);
nand U2069 (N_2069,N_1108,N_807);
nor U2070 (N_2070,N_1107,N_1399);
nand U2071 (N_2071,N_1423,N_786);
nor U2072 (N_2072,N_878,N_1397);
nand U2073 (N_2073,N_954,N_1315);
nor U2074 (N_2074,N_953,N_791);
or U2075 (N_2075,N_1118,N_1272);
and U2076 (N_2076,N_972,N_878);
nor U2077 (N_2077,N_1066,N_931);
or U2078 (N_2078,N_1425,N_998);
nand U2079 (N_2079,N_1329,N_933);
nand U2080 (N_2080,N_1009,N_1163);
nor U2081 (N_2081,N_1342,N_1267);
nand U2082 (N_2082,N_957,N_1438);
nor U2083 (N_2083,N_1362,N_1467);
xnor U2084 (N_2084,N_1296,N_1126);
or U2085 (N_2085,N_888,N_1389);
or U2086 (N_2086,N_1086,N_1106);
nand U2087 (N_2087,N_845,N_1109);
or U2088 (N_2088,N_1393,N_858);
or U2089 (N_2089,N_1029,N_1467);
and U2090 (N_2090,N_990,N_1001);
nand U2091 (N_2091,N_1159,N_1107);
or U2092 (N_2092,N_1104,N_1113);
nand U2093 (N_2093,N_1381,N_793);
or U2094 (N_2094,N_837,N_950);
nand U2095 (N_2095,N_1290,N_1413);
nand U2096 (N_2096,N_880,N_930);
and U2097 (N_2097,N_1463,N_1399);
nor U2098 (N_2098,N_837,N_989);
and U2099 (N_2099,N_1114,N_1354);
and U2100 (N_2100,N_1406,N_1480);
or U2101 (N_2101,N_1394,N_1204);
and U2102 (N_2102,N_762,N_1341);
or U2103 (N_2103,N_1274,N_1191);
or U2104 (N_2104,N_1357,N_874);
nand U2105 (N_2105,N_1017,N_1404);
nor U2106 (N_2106,N_1361,N_1023);
nor U2107 (N_2107,N_1374,N_1091);
nor U2108 (N_2108,N_843,N_818);
nor U2109 (N_2109,N_952,N_1402);
and U2110 (N_2110,N_950,N_1198);
or U2111 (N_2111,N_848,N_1097);
or U2112 (N_2112,N_915,N_914);
and U2113 (N_2113,N_1100,N_1438);
nor U2114 (N_2114,N_1403,N_1223);
and U2115 (N_2115,N_1447,N_1397);
nor U2116 (N_2116,N_998,N_1466);
nor U2117 (N_2117,N_1280,N_784);
nor U2118 (N_2118,N_1337,N_1395);
or U2119 (N_2119,N_961,N_1170);
and U2120 (N_2120,N_1285,N_875);
and U2121 (N_2121,N_893,N_1347);
and U2122 (N_2122,N_927,N_1046);
nand U2123 (N_2123,N_793,N_784);
and U2124 (N_2124,N_1420,N_1276);
or U2125 (N_2125,N_1231,N_1137);
nor U2126 (N_2126,N_1373,N_1332);
or U2127 (N_2127,N_921,N_812);
nor U2128 (N_2128,N_1486,N_909);
or U2129 (N_2129,N_1199,N_978);
nor U2130 (N_2130,N_1187,N_878);
nand U2131 (N_2131,N_1069,N_765);
nand U2132 (N_2132,N_1239,N_1146);
and U2133 (N_2133,N_751,N_1457);
or U2134 (N_2134,N_1055,N_1431);
or U2135 (N_2135,N_1443,N_1078);
nor U2136 (N_2136,N_1370,N_1241);
or U2137 (N_2137,N_822,N_1302);
nand U2138 (N_2138,N_1088,N_948);
or U2139 (N_2139,N_1446,N_1029);
nor U2140 (N_2140,N_1146,N_1477);
and U2141 (N_2141,N_1417,N_835);
xor U2142 (N_2142,N_1144,N_1012);
or U2143 (N_2143,N_1413,N_1092);
xnor U2144 (N_2144,N_857,N_1223);
or U2145 (N_2145,N_1247,N_1485);
nand U2146 (N_2146,N_1024,N_873);
and U2147 (N_2147,N_1063,N_1411);
nand U2148 (N_2148,N_1347,N_783);
or U2149 (N_2149,N_907,N_1136);
or U2150 (N_2150,N_1454,N_821);
or U2151 (N_2151,N_1142,N_944);
nor U2152 (N_2152,N_1117,N_1109);
or U2153 (N_2153,N_967,N_874);
or U2154 (N_2154,N_1144,N_855);
and U2155 (N_2155,N_806,N_1092);
and U2156 (N_2156,N_812,N_1204);
or U2157 (N_2157,N_1359,N_1281);
xor U2158 (N_2158,N_1129,N_893);
nand U2159 (N_2159,N_1459,N_990);
or U2160 (N_2160,N_1255,N_1437);
nor U2161 (N_2161,N_1495,N_978);
xnor U2162 (N_2162,N_920,N_919);
or U2163 (N_2163,N_899,N_1148);
xor U2164 (N_2164,N_834,N_1324);
nand U2165 (N_2165,N_1334,N_981);
nand U2166 (N_2166,N_1260,N_1366);
and U2167 (N_2167,N_1010,N_819);
and U2168 (N_2168,N_784,N_994);
nor U2169 (N_2169,N_840,N_1200);
nor U2170 (N_2170,N_1212,N_768);
and U2171 (N_2171,N_911,N_818);
and U2172 (N_2172,N_1242,N_1322);
nor U2173 (N_2173,N_1170,N_1048);
and U2174 (N_2174,N_971,N_1290);
and U2175 (N_2175,N_1022,N_1434);
or U2176 (N_2176,N_1101,N_1131);
and U2177 (N_2177,N_859,N_1372);
nand U2178 (N_2178,N_759,N_1190);
nand U2179 (N_2179,N_753,N_1063);
or U2180 (N_2180,N_1072,N_1287);
or U2181 (N_2181,N_1041,N_1103);
nor U2182 (N_2182,N_1191,N_1040);
xor U2183 (N_2183,N_1441,N_1155);
nor U2184 (N_2184,N_947,N_1368);
nor U2185 (N_2185,N_1071,N_1195);
or U2186 (N_2186,N_863,N_1407);
xnor U2187 (N_2187,N_1259,N_875);
nand U2188 (N_2188,N_780,N_1364);
nor U2189 (N_2189,N_938,N_815);
nand U2190 (N_2190,N_1285,N_1016);
or U2191 (N_2191,N_1062,N_1389);
nand U2192 (N_2192,N_1424,N_1369);
or U2193 (N_2193,N_1010,N_867);
nand U2194 (N_2194,N_1222,N_921);
nor U2195 (N_2195,N_1015,N_1440);
and U2196 (N_2196,N_824,N_1055);
nor U2197 (N_2197,N_1329,N_894);
nand U2198 (N_2198,N_1431,N_1015);
and U2199 (N_2199,N_1446,N_1254);
or U2200 (N_2200,N_1468,N_1296);
xor U2201 (N_2201,N_1169,N_1438);
nand U2202 (N_2202,N_1297,N_1155);
nand U2203 (N_2203,N_877,N_899);
xnor U2204 (N_2204,N_863,N_1424);
nand U2205 (N_2205,N_1240,N_1286);
nor U2206 (N_2206,N_1314,N_1169);
nor U2207 (N_2207,N_1381,N_1004);
nand U2208 (N_2208,N_1417,N_1347);
or U2209 (N_2209,N_1122,N_976);
nor U2210 (N_2210,N_1344,N_1221);
or U2211 (N_2211,N_763,N_853);
nor U2212 (N_2212,N_1017,N_991);
and U2213 (N_2213,N_1207,N_1040);
xor U2214 (N_2214,N_1095,N_1381);
nand U2215 (N_2215,N_1456,N_1060);
nor U2216 (N_2216,N_813,N_972);
nor U2217 (N_2217,N_1235,N_1420);
nor U2218 (N_2218,N_925,N_1464);
or U2219 (N_2219,N_1196,N_1267);
or U2220 (N_2220,N_976,N_1216);
or U2221 (N_2221,N_760,N_858);
and U2222 (N_2222,N_1120,N_793);
and U2223 (N_2223,N_757,N_1432);
or U2224 (N_2224,N_1084,N_1352);
or U2225 (N_2225,N_983,N_883);
or U2226 (N_2226,N_845,N_1473);
nor U2227 (N_2227,N_1002,N_812);
nor U2228 (N_2228,N_829,N_1022);
and U2229 (N_2229,N_1225,N_1170);
xnor U2230 (N_2230,N_1309,N_981);
or U2231 (N_2231,N_1258,N_959);
nor U2232 (N_2232,N_1017,N_1182);
and U2233 (N_2233,N_1062,N_952);
nor U2234 (N_2234,N_1291,N_1400);
nor U2235 (N_2235,N_1177,N_775);
nor U2236 (N_2236,N_870,N_1145);
or U2237 (N_2237,N_1262,N_1209);
nand U2238 (N_2238,N_960,N_813);
or U2239 (N_2239,N_1201,N_817);
or U2240 (N_2240,N_904,N_1109);
nand U2241 (N_2241,N_887,N_930);
nor U2242 (N_2242,N_799,N_1217);
xnor U2243 (N_2243,N_914,N_1452);
nand U2244 (N_2244,N_814,N_1305);
nand U2245 (N_2245,N_1101,N_1116);
and U2246 (N_2246,N_1325,N_846);
or U2247 (N_2247,N_986,N_1032);
or U2248 (N_2248,N_933,N_1028);
nand U2249 (N_2249,N_1005,N_923);
nand U2250 (N_2250,N_1728,N_1734);
or U2251 (N_2251,N_1855,N_1525);
xor U2252 (N_2252,N_2086,N_2131);
nand U2253 (N_2253,N_1959,N_1910);
nor U2254 (N_2254,N_2002,N_1938);
and U2255 (N_2255,N_2036,N_2158);
nor U2256 (N_2256,N_1864,N_1898);
nor U2257 (N_2257,N_1754,N_1592);
and U2258 (N_2258,N_1582,N_1552);
and U2259 (N_2259,N_2046,N_1749);
xor U2260 (N_2260,N_1936,N_2085);
or U2261 (N_2261,N_1577,N_2223);
or U2262 (N_2262,N_2205,N_1576);
and U2263 (N_2263,N_2164,N_2069);
nand U2264 (N_2264,N_2238,N_2121);
nand U2265 (N_2265,N_2109,N_1675);
xor U2266 (N_2266,N_1645,N_1685);
or U2267 (N_2267,N_1660,N_1606);
nand U2268 (N_2268,N_2072,N_2022);
nor U2269 (N_2269,N_2027,N_1639);
or U2270 (N_2270,N_1913,N_1500);
xnor U2271 (N_2271,N_1989,N_1786);
nor U2272 (N_2272,N_2242,N_2123);
nor U2273 (N_2273,N_2170,N_1671);
xnor U2274 (N_2274,N_1766,N_2004);
nor U2275 (N_2275,N_2106,N_1933);
nor U2276 (N_2276,N_1580,N_1852);
nor U2277 (N_2277,N_1862,N_2091);
nand U2278 (N_2278,N_1563,N_1968);
nand U2279 (N_2279,N_1701,N_1883);
or U2280 (N_2280,N_1543,N_1976);
nand U2281 (N_2281,N_1630,N_2044);
nor U2282 (N_2282,N_1631,N_2203);
or U2283 (N_2283,N_1511,N_1668);
nor U2284 (N_2284,N_2246,N_1775);
or U2285 (N_2285,N_1920,N_1697);
nor U2286 (N_2286,N_1653,N_2200);
nor U2287 (N_2287,N_1983,N_1847);
nor U2288 (N_2288,N_1849,N_1622);
and U2289 (N_2289,N_2077,N_1889);
or U2290 (N_2290,N_1732,N_2162);
and U2291 (N_2291,N_1941,N_1978);
nand U2292 (N_2292,N_1664,N_1969);
nor U2293 (N_2293,N_2034,N_2165);
nor U2294 (N_2294,N_2065,N_2189);
nand U2295 (N_2295,N_1584,N_1611);
xor U2296 (N_2296,N_1808,N_1863);
nand U2297 (N_2297,N_1869,N_2008);
and U2298 (N_2298,N_1906,N_1946);
nor U2299 (N_2299,N_1757,N_2110);
nor U2300 (N_2300,N_2228,N_2089);
or U2301 (N_2301,N_2060,N_1706);
nor U2302 (N_2302,N_2171,N_1939);
xor U2303 (N_2303,N_1950,N_2168);
nor U2304 (N_2304,N_2057,N_1974);
nor U2305 (N_2305,N_2145,N_1719);
xor U2306 (N_2306,N_1957,N_1598);
or U2307 (N_2307,N_1627,N_1547);
nand U2308 (N_2308,N_1878,N_2003);
xnor U2309 (N_2309,N_1851,N_2074);
xnor U2310 (N_2310,N_1517,N_2181);
nand U2311 (N_2311,N_1528,N_2218);
nor U2312 (N_2312,N_1680,N_1977);
nand U2313 (N_2313,N_1561,N_1894);
and U2314 (N_2314,N_1942,N_1635);
nand U2315 (N_2315,N_1515,N_1642);
nor U2316 (N_2316,N_1572,N_1811);
or U2317 (N_2317,N_1505,N_1794);
nor U2318 (N_2318,N_2155,N_2204);
nor U2319 (N_2319,N_2076,N_2169);
xor U2320 (N_2320,N_1996,N_2201);
nand U2321 (N_2321,N_2113,N_2220);
nor U2322 (N_2322,N_1909,N_2239);
and U2323 (N_2323,N_1566,N_1843);
or U2324 (N_2324,N_1917,N_1540);
nand U2325 (N_2325,N_2081,N_1813);
nand U2326 (N_2326,N_1601,N_2066);
xor U2327 (N_2327,N_2000,N_1982);
and U2328 (N_2328,N_1922,N_2088);
xnor U2329 (N_2329,N_1902,N_2111);
nor U2330 (N_2330,N_1778,N_1882);
nor U2331 (N_2331,N_1984,N_2177);
nand U2332 (N_2332,N_1758,N_2127);
xnor U2333 (N_2333,N_1586,N_1617);
and U2334 (N_2334,N_1814,N_1870);
or U2335 (N_2335,N_1944,N_1797);
nor U2336 (N_2336,N_1503,N_1555);
or U2337 (N_2337,N_1747,N_2064);
nor U2338 (N_2338,N_1921,N_1699);
or U2339 (N_2339,N_2068,N_2054);
and U2340 (N_2340,N_1987,N_1830);
or U2341 (N_2341,N_2222,N_1654);
and U2342 (N_2342,N_1735,N_1806);
nand U2343 (N_2343,N_1587,N_2188);
nand U2344 (N_2344,N_1823,N_1764);
nand U2345 (N_2345,N_1613,N_1911);
or U2346 (N_2346,N_1838,N_2184);
nand U2347 (N_2347,N_2151,N_1832);
and U2348 (N_2348,N_1907,N_1568);
nor U2349 (N_2349,N_2048,N_2039);
and U2350 (N_2350,N_1591,N_1824);
nor U2351 (N_2351,N_1840,N_2061);
or U2352 (N_2352,N_2167,N_1924);
nor U2353 (N_2353,N_1696,N_1967);
xnor U2354 (N_2354,N_2119,N_1925);
nor U2355 (N_2355,N_1625,N_1703);
nand U2356 (N_2356,N_1723,N_2197);
or U2357 (N_2357,N_2104,N_1844);
and U2358 (N_2358,N_1678,N_1772);
nand U2359 (N_2359,N_1704,N_1819);
nor U2360 (N_2360,N_2028,N_1776);
xor U2361 (N_2361,N_2080,N_2125);
and U2362 (N_2362,N_1537,N_2142);
nor U2363 (N_2363,N_1546,N_1663);
nor U2364 (N_2364,N_1612,N_1825);
and U2365 (N_2365,N_2118,N_1634);
nand U2366 (N_2366,N_1514,N_1585);
and U2367 (N_2367,N_1960,N_2135);
or U2368 (N_2368,N_1854,N_1655);
nor U2369 (N_2369,N_1965,N_1798);
nor U2370 (N_2370,N_1873,N_2190);
nor U2371 (N_2371,N_2139,N_1686);
nand U2372 (N_2372,N_1805,N_1698);
nor U2373 (N_2373,N_2150,N_1853);
or U2374 (N_2374,N_2143,N_1750);
nor U2375 (N_2375,N_2175,N_1979);
nand U2376 (N_2376,N_1619,N_2112);
nor U2377 (N_2377,N_1717,N_2149);
nand U2378 (N_2378,N_1770,N_1529);
and U2379 (N_2379,N_2247,N_1845);
or U2380 (N_2380,N_2172,N_2115);
xnor U2381 (N_2381,N_1994,N_1595);
nor U2382 (N_2382,N_1573,N_1539);
nor U2383 (N_2383,N_1570,N_2144);
or U2384 (N_2384,N_1709,N_1548);
nand U2385 (N_2385,N_1682,N_1952);
and U2386 (N_2386,N_2030,N_2213);
or U2387 (N_2387,N_1839,N_1677);
xor U2388 (N_2388,N_1727,N_1744);
or U2389 (N_2389,N_1650,N_1900);
nand U2390 (N_2390,N_2221,N_2100);
nand U2391 (N_2391,N_1820,N_1896);
nor U2392 (N_2392,N_2051,N_2037);
and U2393 (N_2393,N_1966,N_1940);
or U2394 (N_2394,N_2212,N_1602);
nand U2395 (N_2395,N_1518,N_2240);
nor U2396 (N_2396,N_1759,N_1662);
and U2397 (N_2397,N_2073,N_1632);
nor U2398 (N_2398,N_1509,N_2024);
nor U2399 (N_2399,N_1857,N_1885);
nand U2400 (N_2400,N_2015,N_1793);
nor U2401 (N_2401,N_1871,N_1652);
and U2402 (N_2402,N_1908,N_1624);
and U2403 (N_2403,N_2063,N_1689);
nand U2404 (N_2404,N_1707,N_1513);
and U2405 (N_2405,N_1623,N_1679);
nor U2406 (N_2406,N_2013,N_1694);
and U2407 (N_2407,N_1720,N_1599);
nor U2408 (N_2408,N_2079,N_2047);
and U2409 (N_2409,N_1519,N_1746);
or U2410 (N_2410,N_1608,N_1809);
xor U2411 (N_2411,N_1722,N_1914);
nor U2412 (N_2412,N_1904,N_2210);
nor U2413 (N_2413,N_1700,N_1716);
nor U2414 (N_2414,N_1918,N_2202);
and U2415 (N_2415,N_2192,N_1767);
or U2416 (N_2416,N_1554,N_1861);
and U2417 (N_2417,N_2237,N_1648);
or U2418 (N_2418,N_2173,N_1985);
and U2419 (N_2419,N_2154,N_2059);
and U2420 (N_2420,N_2178,N_1789);
xor U2421 (N_2421,N_1559,N_2161);
nand U2422 (N_2422,N_1783,N_2067);
nand U2423 (N_2423,N_1842,N_1616);
or U2424 (N_2424,N_1784,N_2001);
and U2425 (N_2425,N_1667,N_1866);
or U2426 (N_2426,N_1674,N_2122);
xor U2427 (N_2427,N_1708,N_2137);
and U2428 (N_2428,N_1715,N_2208);
or U2429 (N_2429,N_2095,N_2219);
and U2430 (N_2430,N_2092,N_1551);
and U2431 (N_2431,N_1726,N_1901);
or U2432 (N_2432,N_1981,N_1721);
nor U2433 (N_2433,N_1589,N_1618);
xor U2434 (N_2434,N_1567,N_2120);
nand U2435 (N_2435,N_1545,N_1964);
nand U2436 (N_2436,N_1512,N_1988);
nand U2437 (N_2437,N_1590,N_1858);
xor U2438 (N_2438,N_1741,N_2217);
and U2439 (N_2439,N_2214,N_2182);
and U2440 (N_2440,N_1995,N_1993);
xor U2441 (N_2441,N_1876,N_1737);
or U2442 (N_2442,N_1807,N_1676);
nand U2443 (N_2443,N_2019,N_2006);
nand U2444 (N_2444,N_1742,N_1868);
nor U2445 (N_2445,N_1542,N_2232);
nand U2446 (N_2446,N_1790,N_1773);
and U2447 (N_2447,N_2031,N_1693);
or U2448 (N_2448,N_2096,N_1822);
nor U2449 (N_2449,N_1571,N_1526);
nor U2450 (N_2450,N_1812,N_1533);
and U2451 (N_2451,N_2230,N_1897);
or U2452 (N_2452,N_2117,N_1986);
nand U2453 (N_2453,N_1507,N_2058);
nand U2454 (N_2454,N_1828,N_1795);
nor U2455 (N_2455,N_1597,N_1934);
nor U2456 (N_2456,N_1771,N_1818);
nor U2457 (N_2457,N_1780,N_1534);
nor U2458 (N_2458,N_2234,N_2099);
nor U2459 (N_2459,N_1927,N_2134);
nor U2460 (N_2460,N_2056,N_1739);
or U2461 (N_2461,N_1575,N_2248);
nor U2462 (N_2462,N_1769,N_1666);
or U2463 (N_2463,N_2020,N_1532);
or U2464 (N_2464,N_1998,N_1535);
nor U2465 (N_2465,N_1928,N_1801);
nor U2466 (N_2466,N_1992,N_1743);
or U2467 (N_2467,N_1804,N_1530);
and U2468 (N_2468,N_2166,N_1997);
or U2469 (N_2469,N_2009,N_2185);
nor U2470 (N_2470,N_1827,N_1796);
nor U2471 (N_2471,N_2041,N_1714);
or U2472 (N_2472,N_2207,N_2183);
or U2473 (N_2473,N_1916,N_2224);
and U2474 (N_2474,N_1765,N_1829);
and U2475 (N_2475,N_2007,N_2016);
nor U2476 (N_2476,N_1893,N_1712);
nor U2477 (N_2477,N_2045,N_2021);
nor U2478 (N_2478,N_2094,N_2071);
and U2479 (N_2479,N_1879,N_1761);
xor U2480 (N_2480,N_1629,N_2138);
or U2481 (N_2481,N_2026,N_2231);
xor U2482 (N_2482,N_1596,N_2235);
nand U2483 (N_2483,N_2244,N_1903);
xor U2484 (N_2484,N_1915,N_1673);
and U2485 (N_2485,N_1833,N_1886);
and U2486 (N_2486,N_2038,N_1640);
and U2487 (N_2487,N_1705,N_2093);
nor U2488 (N_2488,N_1508,N_1972);
nor U2489 (N_2489,N_1929,N_2102);
or U2490 (N_2490,N_1930,N_2157);
nand U2491 (N_2491,N_1651,N_2014);
and U2492 (N_2492,N_1605,N_1756);
or U2493 (N_2493,N_1877,N_1945);
nand U2494 (N_2494,N_2194,N_1541);
nor U2495 (N_2495,N_2129,N_1558);
nor U2496 (N_2496,N_2035,N_1890);
nand U2497 (N_2497,N_2160,N_1684);
or U2498 (N_2498,N_1557,N_2078);
and U2499 (N_2499,N_1755,N_1799);
nor U2500 (N_2500,N_1884,N_1949);
and U2501 (N_2501,N_1753,N_1875);
or U2502 (N_2502,N_1955,N_1791);
nand U2503 (N_2503,N_1609,N_1821);
nand U2504 (N_2504,N_1691,N_2176);
nor U2505 (N_2505,N_2032,N_1656);
and U2506 (N_2506,N_1569,N_2163);
nand U2507 (N_2507,N_2141,N_1975);
or U2508 (N_2508,N_2196,N_2108);
nor U2509 (N_2509,N_1502,N_1895);
nand U2510 (N_2510,N_1649,N_2245);
and U2511 (N_2511,N_1549,N_1725);
nand U2512 (N_2512,N_1636,N_1603);
nor U2513 (N_2513,N_2195,N_2098);
nor U2514 (N_2514,N_1961,N_1688);
or U2515 (N_2515,N_2243,N_2055);
or U2516 (N_2516,N_1657,N_1583);
and U2517 (N_2517,N_2049,N_1681);
and U2518 (N_2518,N_1637,N_2236);
nor U2519 (N_2519,N_2075,N_1520);
nand U2520 (N_2520,N_2211,N_2156);
or U2521 (N_2521,N_1850,N_1848);
and U2522 (N_2522,N_1745,N_2090);
nor U2523 (N_2523,N_2070,N_2130);
and U2524 (N_2524,N_1644,N_1579);
nand U2525 (N_2525,N_1837,N_1856);
nor U2526 (N_2526,N_2193,N_1815);
nand U2527 (N_2527,N_2082,N_1521);
or U2528 (N_2528,N_1710,N_2226);
nand U2529 (N_2529,N_1970,N_1971);
and U2530 (N_2530,N_1788,N_1553);
and U2531 (N_2531,N_1835,N_1594);
nor U2532 (N_2532,N_1779,N_2133);
or U2533 (N_2533,N_1730,N_1588);
xnor U2534 (N_2534,N_2062,N_1687);
nor U2535 (N_2535,N_1607,N_2042);
nand U2536 (N_2536,N_1792,N_1802);
or U2537 (N_2537,N_2087,N_1860);
nand U2538 (N_2538,N_1919,N_1736);
nor U2539 (N_2539,N_1956,N_2023);
or U2540 (N_2540,N_2040,N_2128);
xor U2541 (N_2541,N_2052,N_1963);
or U2542 (N_2542,N_1516,N_1556);
xor U2543 (N_2543,N_1880,N_1943);
nand U2544 (N_2544,N_2227,N_1544);
nand U2545 (N_2545,N_1810,N_1841);
or U2546 (N_2546,N_1669,N_1581);
nand U2547 (N_2547,N_1690,N_1504);
xnor U2548 (N_2548,N_1800,N_1670);
or U2549 (N_2549,N_2103,N_1641);
or U2550 (N_2550,N_1610,N_1781);
nor U2551 (N_2551,N_1932,N_1638);
and U2552 (N_2552,N_1768,N_2114);
nor U2553 (N_2553,N_1962,N_1774);
or U2554 (N_2554,N_2215,N_1643);
or U2555 (N_2555,N_1762,N_1836);
nor U2556 (N_2556,N_1931,N_1527);
xor U2557 (N_2557,N_2107,N_1522);
nor U2558 (N_2558,N_2116,N_2005);
nor U2559 (N_2559,N_1958,N_1899);
nand U2560 (N_2560,N_2018,N_1999);
nand U2561 (N_2561,N_2084,N_1887);
and U2562 (N_2562,N_1954,N_2029);
nor U2563 (N_2563,N_1752,N_1615);
and U2564 (N_2564,N_1923,N_1510);
xnor U2565 (N_2565,N_1991,N_2179);
or U2566 (N_2566,N_1817,N_1536);
and U2567 (N_2567,N_1702,N_1733);
nor U2568 (N_2568,N_1658,N_2146);
and U2569 (N_2569,N_1729,N_1738);
or U2570 (N_2570,N_1935,N_1748);
and U2571 (N_2571,N_1621,N_1633);
nand U2572 (N_2572,N_2033,N_2132);
nor U2573 (N_2573,N_1891,N_1614);
nand U2574 (N_2574,N_1523,N_1816);
and U2575 (N_2575,N_1659,N_2225);
xnor U2576 (N_2576,N_1990,N_2174);
or U2577 (N_2577,N_1626,N_1951);
or U2578 (N_2578,N_2012,N_2233);
nor U2579 (N_2579,N_2191,N_1953);
nor U2580 (N_2580,N_1565,N_1782);
nand U2581 (N_2581,N_1600,N_1531);
nor U2582 (N_2582,N_1905,N_1785);
xnor U2583 (N_2583,N_1711,N_1578);
and U2584 (N_2584,N_1646,N_1846);
nand U2585 (N_2585,N_1593,N_2198);
or U2586 (N_2586,N_2017,N_2148);
and U2587 (N_2587,N_2180,N_1724);
nand U2588 (N_2588,N_2159,N_1777);
and U2589 (N_2589,N_1665,N_1872);
and U2590 (N_2590,N_1672,N_1760);
nand U2591 (N_2591,N_2050,N_1751);
xnor U2592 (N_2592,N_1973,N_1859);
nor U2593 (N_2593,N_1506,N_1867);
or U2594 (N_2594,N_1731,N_1550);
or U2595 (N_2595,N_1948,N_1881);
or U2596 (N_2596,N_2187,N_1713);
xnor U2597 (N_2597,N_2199,N_1740);
nor U2598 (N_2598,N_1826,N_2126);
xor U2599 (N_2599,N_1874,N_2206);
or U2600 (N_2600,N_2136,N_2147);
or U2601 (N_2601,N_1501,N_2101);
nor U2602 (N_2602,N_1524,N_2053);
nor U2603 (N_2603,N_1865,N_1692);
and U2604 (N_2604,N_1628,N_1834);
nor U2605 (N_2605,N_1888,N_2152);
nor U2606 (N_2606,N_2140,N_1912);
nand U2607 (N_2607,N_1763,N_2241);
nand U2608 (N_2608,N_2229,N_2011);
nand U2609 (N_2609,N_2043,N_1831);
and U2610 (N_2610,N_1574,N_2186);
or U2611 (N_2611,N_1564,N_1695);
and U2612 (N_2612,N_1787,N_1604);
and U2613 (N_2613,N_1620,N_1803);
nand U2614 (N_2614,N_1560,N_1647);
and U2615 (N_2615,N_1947,N_2249);
nor U2616 (N_2616,N_2153,N_2025);
or U2617 (N_2617,N_1926,N_1562);
nor U2618 (N_2618,N_2083,N_1892);
or U2619 (N_2619,N_1683,N_1661);
xor U2620 (N_2620,N_1538,N_1980);
xor U2621 (N_2621,N_2105,N_2216);
and U2622 (N_2622,N_2097,N_1718);
xnor U2623 (N_2623,N_2124,N_2010);
nor U2624 (N_2624,N_2209,N_1937);
and U2625 (N_2625,N_1821,N_2167);
nand U2626 (N_2626,N_1913,N_2066);
nand U2627 (N_2627,N_1526,N_1570);
nor U2628 (N_2628,N_2242,N_1796);
and U2629 (N_2629,N_2088,N_1809);
xor U2630 (N_2630,N_1972,N_1532);
nor U2631 (N_2631,N_2176,N_2247);
and U2632 (N_2632,N_1964,N_1639);
or U2633 (N_2633,N_1970,N_1565);
or U2634 (N_2634,N_1806,N_1844);
xnor U2635 (N_2635,N_2062,N_1540);
xor U2636 (N_2636,N_1611,N_1532);
nand U2637 (N_2637,N_2224,N_1835);
or U2638 (N_2638,N_1907,N_1639);
nand U2639 (N_2639,N_2120,N_1861);
or U2640 (N_2640,N_1751,N_1516);
nand U2641 (N_2641,N_1989,N_1659);
and U2642 (N_2642,N_2217,N_1520);
nor U2643 (N_2643,N_1549,N_1578);
nand U2644 (N_2644,N_1567,N_1710);
nor U2645 (N_2645,N_1680,N_1957);
xor U2646 (N_2646,N_1864,N_1631);
or U2647 (N_2647,N_1686,N_2084);
nor U2648 (N_2648,N_1657,N_1793);
or U2649 (N_2649,N_2083,N_2050);
or U2650 (N_2650,N_2135,N_2045);
or U2651 (N_2651,N_1922,N_1638);
or U2652 (N_2652,N_1871,N_1524);
nand U2653 (N_2653,N_1862,N_1594);
nand U2654 (N_2654,N_2025,N_2124);
nor U2655 (N_2655,N_1880,N_1900);
or U2656 (N_2656,N_1765,N_2059);
nor U2657 (N_2657,N_1852,N_1610);
nor U2658 (N_2658,N_1779,N_2136);
nor U2659 (N_2659,N_1614,N_2105);
nand U2660 (N_2660,N_2203,N_2005);
or U2661 (N_2661,N_1720,N_1944);
and U2662 (N_2662,N_2061,N_2209);
nor U2663 (N_2663,N_1621,N_1936);
nor U2664 (N_2664,N_2069,N_1814);
and U2665 (N_2665,N_2244,N_2181);
xnor U2666 (N_2666,N_1827,N_1533);
nor U2667 (N_2667,N_1897,N_2212);
and U2668 (N_2668,N_1516,N_1908);
xor U2669 (N_2669,N_1928,N_1843);
nor U2670 (N_2670,N_2105,N_1860);
nand U2671 (N_2671,N_2119,N_1981);
or U2672 (N_2672,N_2230,N_1585);
and U2673 (N_2673,N_1849,N_2023);
nor U2674 (N_2674,N_2170,N_1924);
or U2675 (N_2675,N_2247,N_2194);
and U2676 (N_2676,N_2178,N_2036);
or U2677 (N_2677,N_1857,N_2048);
nand U2678 (N_2678,N_1717,N_1542);
and U2679 (N_2679,N_1745,N_1501);
xor U2680 (N_2680,N_1623,N_1605);
and U2681 (N_2681,N_2030,N_1839);
nor U2682 (N_2682,N_1800,N_1592);
or U2683 (N_2683,N_2023,N_1760);
nand U2684 (N_2684,N_1922,N_1540);
and U2685 (N_2685,N_1939,N_2246);
nor U2686 (N_2686,N_1665,N_2007);
and U2687 (N_2687,N_2065,N_2042);
nor U2688 (N_2688,N_2028,N_1709);
and U2689 (N_2689,N_2013,N_2095);
or U2690 (N_2690,N_2078,N_1927);
and U2691 (N_2691,N_2228,N_1655);
xor U2692 (N_2692,N_1786,N_1615);
or U2693 (N_2693,N_2083,N_1512);
or U2694 (N_2694,N_1670,N_2225);
nor U2695 (N_2695,N_2002,N_2119);
and U2696 (N_2696,N_1639,N_1828);
and U2697 (N_2697,N_1694,N_1530);
nand U2698 (N_2698,N_1678,N_2199);
nor U2699 (N_2699,N_2175,N_1672);
and U2700 (N_2700,N_2163,N_2000);
or U2701 (N_2701,N_1590,N_2186);
nor U2702 (N_2702,N_1737,N_2106);
nand U2703 (N_2703,N_2157,N_1781);
and U2704 (N_2704,N_1832,N_2228);
or U2705 (N_2705,N_1509,N_1920);
xor U2706 (N_2706,N_2231,N_2013);
nor U2707 (N_2707,N_1992,N_2107);
nand U2708 (N_2708,N_2174,N_2055);
nand U2709 (N_2709,N_2186,N_1648);
and U2710 (N_2710,N_2005,N_2213);
and U2711 (N_2711,N_2052,N_1857);
xor U2712 (N_2712,N_1936,N_1591);
and U2713 (N_2713,N_1720,N_1687);
or U2714 (N_2714,N_1777,N_1880);
nor U2715 (N_2715,N_2213,N_2108);
and U2716 (N_2716,N_1770,N_1642);
nand U2717 (N_2717,N_1738,N_1554);
nand U2718 (N_2718,N_1552,N_2208);
nand U2719 (N_2719,N_1933,N_1787);
xnor U2720 (N_2720,N_1809,N_1663);
or U2721 (N_2721,N_1525,N_1772);
xnor U2722 (N_2722,N_2060,N_2071);
or U2723 (N_2723,N_2044,N_1700);
and U2724 (N_2724,N_1559,N_1659);
and U2725 (N_2725,N_1866,N_1993);
nor U2726 (N_2726,N_1812,N_2098);
xor U2727 (N_2727,N_1557,N_2163);
nand U2728 (N_2728,N_2159,N_1954);
and U2729 (N_2729,N_1724,N_2015);
or U2730 (N_2730,N_2243,N_1894);
nor U2731 (N_2731,N_1587,N_2018);
and U2732 (N_2732,N_2245,N_1658);
and U2733 (N_2733,N_1839,N_1935);
nand U2734 (N_2734,N_2204,N_2187);
nor U2735 (N_2735,N_2040,N_1526);
nand U2736 (N_2736,N_1779,N_2000);
nand U2737 (N_2737,N_1661,N_2079);
nand U2738 (N_2738,N_1810,N_2042);
or U2739 (N_2739,N_1647,N_1690);
xnor U2740 (N_2740,N_2031,N_1741);
xnor U2741 (N_2741,N_1658,N_1885);
and U2742 (N_2742,N_1665,N_1698);
and U2743 (N_2743,N_2214,N_1506);
and U2744 (N_2744,N_1932,N_1604);
xnor U2745 (N_2745,N_1813,N_1843);
nand U2746 (N_2746,N_2111,N_1890);
or U2747 (N_2747,N_1848,N_2021);
nand U2748 (N_2748,N_2142,N_1945);
and U2749 (N_2749,N_1734,N_1832);
or U2750 (N_2750,N_2100,N_1608);
or U2751 (N_2751,N_1789,N_1668);
and U2752 (N_2752,N_1879,N_1783);
or U2753 (N_2753,N_1805,N_1544);
nand U2754 (N_2754,N_2021,N_2118);
nand U2755 (N_2755,N_1581,N_1638);
and U2756 (N_2756,N_1776,N_1696);
and U2757 (N_2757,N_1519,N_2075);
nand U2758 (N_2758,N_1620,N_1608);
xor U2759 (N_2759,N_2020,N_1990);
nor U2760 (N_2760,N_1584,N_2175);
or U2761 (N_2761,N_2104,N_1711);
nor U2762 (N_2762,N_1796,N_1614);
nand U2763 (N_2763,N_1542,N_2176);
xnor U2764 (N_2764,N_1657,N_1820);
nor U2765 (N_2765,N_2236,N_2090);
and U2766 (N_2766,N_1926,N_2019);
or U2767 (N_2767,N_2005,N_1514);
or U2768 (N_2768,N_2067,N_2032);
nor U2769 (N_2769,N_1591,N_1934);
nand U2770 (N_2770,N_1845,N_1811);
nand U2771 (N_2771,N_1885,N_1600);
and U2772 (N_2772,N_1763,N_1611);
nand U2773 (N_2773,N_1879,N_1758);
xnor U2774 (N_2774,N_1692,N_1524);
or U2775 (N_2775,N_1943,N_1512);
nand U2776 (N_2776,N_1824,N_1850);
or U2777 (N_2777,N_1526,N_2013);
nor U2778 (N_2778,N_2122,N_2149);
nand U2779 (N_2779,N_1749,N_2037);
nand U2780 (N_2780,N_2219,N_1788);
nand U2781 (N_2781,N_2093,N_1923);
nor U2782 (N_2782,N_1514,N_1509);
nand U2783 (N_2783,N_1549,N_1634);
and U2784 (N_2784,N_1538,N_2217);
or U2785 (N_2785,N_1959,N_1739);
and U2786 (N_2786,N_2007,N_1699);
and U2787 (N_2787,N_1560,N_1875);
xnor U2788 (N_2788,N_2008,N_1502);
nor U2789 (N_2789,N_2225,N_1621);
nor U2790 (N_2790,N_1625,N_2136);
xnor U2791 (N_2791,N_1641,N_1573);
nor U2792 (N_2792,N_1931,N_1555);
or U2793 (N_2793,N_2043,N_1558);
and U2794 (N_2794,N_2056,N_2040);
or U2795 (N_2795,N_1639,N_2062);
nand U2796 (N_2796,N_1970,N_1569);
nor U2797 (N_2797,N_2206,N_1676);
nand U2798 (N_2798,N_2153,N_1581);
nor U2799 (N_2799,N_2003,N_1964);
or U2800 (N_2800,N_1977,N_1774);
and U2801 (N_2801,N_1803,N_2241);
or U2802 (N_2802,N_1991,N_1509);
nand U2803 (N_2803,N_1863,N_1711);
nor U2804 (N_2804,N_1652,N_1974);
nand U2805 (N_2805,N_1911,N_1566);
nor U2806 (N_2806,N_1589,N_2216);
nand U2807 (N_2807,N_2100,N_1587);
nand U2808 (N_2808,N_1675,N_1876);
nand U2809 (N_2809,N_1742,N_1629);
or U2810 (N_2810,N_1943,N_1763);
nand U2811 (N_2811,N_1945,N_2063);
and U2812 (N_2812,N_1774,N_1643);
or U2813 (N_2813,N_1843,N_2087);
or U2814 (N_2814,N_1564,N_2058);
and U2815 (N_2815,N_1774,N_2247);
nand U2816 (N_2816,N_2111,N_1973);
and U2817 (N_2817,N_1669,N_1769);
and U2818 (N_2818,N_1990,N_1528);
or U2819 (N_2819,N_1983,N_1827);
and U2820 (N_2820,N_2089,N_1639);
and U2821 (N_2821,N_1972,N_1681);
or U2822 (N_2822,N_2061,N_1639);
nand U2823 (N_2823,N_1838,N_2249);
nor U2824 (N_2824,N_1837,N_2056);
nor U2825 (N_2825,N_1798,N_1915);
nand U2826 (N_2826,N_2007,N_1990);
nand U2827 (N_2827,N_2029,N_1960);
or U2828 (N_2828,N_1757,N_1947);
and U2829 (N_2829,N_1726,N_1854);
or U2830 (N_2830,N_1775,N_2231);
nand U2831 (N_2831,N_2153,N_1781);
or U2832 (N_2832,N_1717,N_1638);
and U2833 (N_2833,N_1921,N_2134);
and U2834 (N_2834,N_1924,N_1584);
nor U2835 (N_2835,N_1972,N_1840);
or U2836 (N_2836,N_1887,N_1771);
nor U2837 (N_2837,N_1767,N_1580);
nand U2838 (N_2838,N_1908,N_2168);
or U2839 (N_2839,N_1878,N_1839);
nor U2840 (N_2840,N_1946,N_2233);
or U2841 (N_2841,N_2001,N_2232);
or U2842 (N_2842,N_1636,N_1615);
xor U2843 (N_2843,N_1795,N_2151);
and U2844 (N_2844,N_2231,N_2055);
nand U2845 (N_2845,N_1820,N_1677);
nand U2846 (N_2846,N_1658,N_2215);
and U2847 (N_2847,N_2102,N_1687);
xnor U2848 (N_2848,N_1883,N_1766);
or U2849 (N_2849,N_1518,N_2218);
and U2850 (N_2850,N_1851,N_1896);
nor U2851 (N_2851,N_1564,N_2135);
nor U2852 (N_2852,N_2131,N_2152);
or U2853 (N_2853,N_1605,N_1872);
nand U2854 (N_2854,N_2198,N_2010);
xor U2855 (N_2855,N_2066,N_2220);
nor U2856 (N_2856,N_1513,N_1947);
nand U2857 (N_2857,N_1512,N_1683);
nand U2858 (N_2858,N_2191,N_1985);
nor U2859 (N_2859,N_2191,N_1680);
nor U2860 (N_2860,N_2018,N_2187);
or U2861 (N_2861,N_1766,N_2121);
or U2862 (N_2862,N_2212,N_1631);
nand U2863 (N_2863,N_1947,N_2189);
xnor U2864 (N_2864,N_2012,N_2197);
nor U2865 (N_2865,N_2106,N_1654);
or U2866 (N_2866,N_1521,N_1603);
nand U2867 (N_2867,N_2032,N_2203);
xor U2868 (N_2868,N_1776,N_1712);
nor U2869 (N_2869,N_2233,N_1518);
or U2870 (N_2870,N_1701,N_1706);
or U2871 (N_2871,N_1950,N_2218);
or U2872 (N_2872,N_1543,N_1714);
nor U2873 (N_2873,N_1738,N_1725);
or U2874 (N_2874,N_1745,N_1655);
and U2875 (N_2875,N_2204,N_1950);
nand U2876 (N_2876,N_2105,N_2239);
and U2877 (N_2877,N_2204,N_1659);
nor U2878 (N_2878,N_1704,N_1869);
nand U2879 (N_2879,N_1805,N_1758);
or U2880 (N_2880,N_1674,N_1546);
and U2881 (N_2881,N_2234,N_2057);
or U2882 (N_2882,N_2098,N_1808);
nand U2883 (N_2883,N_1863,N_2157);
and U2884 (N_2884,N_2174,N_1516);
xnor U2885 (N_2885,N_1728,N_1740);
nor U2886 (N_2886,N_1973,N_1923);
and U2887 (N_2887,N_1736,N_1590);
xnor U2888 (N_2888,N_2165,N_2051);
xor U2889 (N_2889,N_1616,N_2225);
and U2890 (N_2890,N_1682,N_2034);
and U2891 (N_2891,N_1932,N_2067);
nor U2892 (N_2892,N_1790,N_2167);
or U2893 (N_2893,N_2121,N_1903);
nor U2894 (N_2894,N_2246,N_1530);
or U2895 (N_2895,N_2001,N_2012);
xor U2896 (N_2896,N_1720,N_2222);
xor U2897 (N_2897,N_1954,N_2069);
nand U2898 (N_2898,N_1785,N_2105);
and U2899 (N_2899,N_1655,N_1818);
nand U2900 (N_2900,N_2238,N_1596);
nand U2901 (N_2901,N_1595,N_1825);
nand U2902 (N_2902,N_1981,N_1938);
nor U2903 (N_2903,N_1586,N_1777);
and U2904 (N_2904,N_1795,N_1848);
xnor U2905 (N_2905,N_1500,N_1972);
and U2906 (N_2906,N_1633,N_1629);
or U2907 (N_2907,N_2016,N_1681);
nor U2908 (N_2908,N_1779,N_1712);
and U2909 (N_2909,N_1647,N_1607);
nor U2910 (N_2910,N_2011,N_1522);
and U2911 (N_2911,N_2145,N_1526);
nand U2912 (N_2912,N_1889,N_2197);
xnor U2913 (N_2913,N_2062,N_2214);
and U2914 (N_2914,N_2021,N_2135);
nor U2915 (N_2915,N_1582,N_1996);
nor U2916 (N_2916,N_1679,N_1914);
nor U2917 (N_2917,N_1831,N_1685);
nand U2918 (N_2918,N_1871,N_1930);
or U2919 (N_2919,N_1582,N_1932);
nor U2920 (N_2920,N_2166,N_1843);
nand U2921 (N_2921,N_1692,N_1538);
xor U2922 (N_2922,N_1643,N_1689);
nand U2923 (N_2923,N_1902,N_1788);
nor U2924 (N_2924,N_1986,N_2242);
and U2925 (N_2925,N_2163,N_1889);
nand U2926 (N_2926,N_1641,N_1962);
and U2927 (N_2927,N_2095,N_2108);
or U2928 (N_2928,N_1925,N_2091);
xnor U2929 (N_2929,N_2091,N_1727);
and U2930 (N_2930,N_1572,N_2208);
or U2931 (N_2931,N_1638,N_1908);
or U2932 (N_2932,N_1940,N_2057);
and U2933 (N_2933,N_1831,N_1811);
nor U2934 (N_2934,N_1601,N_1701);
or U2935 (N_2935,N_1607,N_2073);
or U2936 (N_2936,N_2084,N_1603);
nand U2937 (N_2937,N_2101,N_1827);
nor U2938 (N_2938,N_1883,N_1969);
nand U2939 (N_2939,N_1981,N_1790);
and U2940 (N_2940,N_2138,N_1870);
or U2941 (N_2941,N_1756,N_1913);
xor U2942 (N_2942,N_2248,N_2195);
and U2943 (N_2943,N_2249,N_1582);
nand U2944 (N_2944,N_1772,N_1848);
nand U2945 (N_2945,N_1931,N_1963);
nand U2946 (N_2946,N_1549,N_1888);
nand U2947 (N_2947,N_1879,N_2141);
nand U2948 (N_2948,N_1539,N_2080);
and U2949 (N_2949,N_1881,N_1719);
or U2950 (N_2950,N_1845,N_1946);
nor U2951 (N_2951,N_2200,N_2145);
nand U2952 (N_2952,N_2127,N_2219);
and U2953 (N_2953,N_1761,N_1820);
nor U2954 (N_2954,N_2126,N_1513);
nand U2955 (N_2955,N_1742,N_1803);
nand U2956 (N_2956,N_1953,N_2076);
and U2957 (N_2957,N_1730,N_1761);
nand U2958 (N_2958,N_2157,N_1972);
nor U2959 (N_2959,N_1579,N_2152);
and U2960 (N_2960,N_2212,N_1919);
xor U2961 (N_2961,N_1952,N_2052);
nand U2962 (N_2962,N_1965,N_2177);
or U2963 (N_2963,N_2003,N_1872);
nand U2964 (N_2964,N_2237,N_1995);
or U2965 (N_2965,N_1824,N_1990);
or U2966 (N_2966,N_1907,N_1691);
xor U2967 (N_2967,N_1569,N_2236);
and U2968 (N_2968,N_2143,N_2242);
nor U2969 (N_2969,N_2104,N_1814);
nand U2970 (N_2970,N_1889,N_2066);
and U2971 (N_2971,N_2063,N_1874);
or U2972 (N_2972,N_1973,N_1895);
nor U2973 (N_2973,N_1758,N_2007);
nor U2974 (N_2974,N_1970,N_1836);
nand U2975 (N_2975,N_2100,N_1807);
nand U2976 (N_2976,N_1954,N_1977);
nor U2977 (N_2977,N_2030,N_1565);
or U2978 (N_2978,N_1747,N_1978);
nor U2979 (N_2979,N_2009,N_1867);
or U2980 (N_2980,N_1688,N_1877);
nor U2981 (N_2981,N_2118,N_2124);
nand U2982 (N_2982,N_1953,N_1994);
nand U2983 (N_2983,N_2079,N_2203);
or U2984 (N_2984,N_1646,N_1610);
and U2985 (N_2985,N_1727,N_2020);
nand U2986 (N_2986,N_1518,N_1866);
and U2987 (N_2987,N_1686,N_1734);
or U2988 (N_2988,N_1766,N_1802);
xor U2989 (N_2989,N_1735,N_1657);
or U2990 (N_2990,N_2007,N_1602);
xnor U2991 (N_2991,N_1730,N_1793);
nand U2992 (N_2992,N_1677,N_2080);
or U2993 (N_2993,N_1833,N_1724);
nor U2994 (N_2994,N_1573,N_1609);
nor U2995 (N_2995,N_1615,N_1712);
and U2996 (N_2996,N_2001,N_2020);
or U2997 (N_2997,N_2216,N_2169);
or U2998 (N_2998,N_1948,N_2014);
xor U2999 (N_2999,N_2008,N_1704);
and U3000 (N_3000,N_2720,N_2801);
nor U3001 (N_3001,N_2669,N_2849);
xor U3002 (N_3002,N_2876,N_2921);
nand U3003 (N_3003,N_2568,N_2574);
and U3004 (N_3004,N_2345,N_2803);
nor U3005 (N_3005,N_2981,N_2481);
nand U3006 (N_3006,N_2905,N_2280);
nand U3007 (N_3007,N_2368,N_2932);
or U3008 (N_3008,N_2988,N_2486);
xnor U3009 (N_3009,N_2332,N_2974);
nand U3010 (N_3010,N_2617,N_2977);
xnor U3011 (N_3011,N_2415,N_2438);
and U3012 (N_3012,N_2911,N_2753);
nand U3013 (N_3013,N_2567,N_2698);
nor U3014 (N_3014,N_2825,N_2740);
and U3015 (N_3015,N_2928,N_2756);
nor U3016 (N_3016,N_2999,N_2807);
nor U3017 (N_3017,N_2271,N_2809);
or U3018 (N_3018,N_2660,N_2786);
or U3019 (N_3019,N_2638,N_2772);
and U3020 (N_3020,N_2742,N_2830);
nor U3021 (N_3021,N_2556,N_2514);
nand U3022 (N_3022,N_2724,N_2953);
nor U3023 (N_3023,N_2730,N_2750);
or U3024 (N_3024,N_2479,N_2473);
nand U3025 (N_3025,N_2588,N_2907);
or U3026 (N_3026,N_2419,N_2987);
or U3027 (N_3027,N_2393,N_2443);
or U3028 (N_3028,N_2925,N_2603);
or U3029 (N_3029,N_2808,N_2377);
nand U3030 (N_3030,N_2894,N_2610);
xor U3031 (N_3031,N_2731,N_2872);
nand U3032 (N_3032,N_2333,N_2893);
and U3033 (N_3033,N_2755,N_2601);
nor U3034 (N_3034,N_2408,N_2549);
nand U3035 (N_3035,N_2862,N_2963);
or U3036 (N_3036,N_2676,N_2871);
nor U3037 (N_3037,N_2582,N_2653);
or U3038 (N_3038,N_2402,N_2623);
and U3039 (N_3039,N_2557,N_2275);
nand U3040 (N_3040,N_2661,N_2888);
nor U3041 (N_3041,N_2865,N_2372);
nand U3042 (N_3042,N_2650,N_2453);
and U3043 (N_3043,N_2338,N_2790);
nor U3044 (N_3044,N_2533,N_2704);
or U3045 (N_3045,N_2531,N_2655);
or U3046 (N_3046,N_2764,N_2348);
and U3047 (N_3047,N_2535,N_2499);
and U3048 (N_3048,N_2527,N_2710);
xor U3049 (N_3049,N_2708,N_2554);
xnor U3050 (N_3050,N_2477,N_2390);
nor U3051 (N_3051,N_2785,N_2880);
nand U3052 (N_3052,N_2300,N_2256);
or U3053 (N_3053,N_2885,N_2961);
nand U3054 (N_3054,N_2896,N_2856);
nor U3055 (N_3055,N_2826,N_2791);
xnor U3056 (N_3056,N_2298,N_2745);
or U3057 (N_3057,N_2648,N_2841);
nor U3058 (N_3058,N_2383,N_2428);
nor U3059 (N_3059,N_2444,N_2319);
nor U3060 (N_3060,N_2918,N_2409);
or U3061 (N_3061,N_2816,N_2917);
or U3062 (N_3062,N_2339,N_2667);
nor U3063 (N_3063,N_2451,N_2903);
or U3064 (N_3064,N_2314,N_2474);
xnor U3065 (N_3065,N_2370,N_2472);
xnor U3066 (N_3066,N_2886,N_2713);
and U3067 (N_3067,N_2551,N_2829);
nand U3068 (N_3068,N_2620,N_2813);
or U3069 (N_3069,N_2389,N_2746);
or U3070 (N_3070,N_2861,N_2290);
nand U3071 (N_3071,N_2942,N_2406);
and U3072 (N_3072,N_2435,N_2292);
nand U3073 (N_3073,N_2552,N_2553);
and U3074 (N_3074,N_2622,N_2467);
nor U3075 (N_3075,N_2421,N_2404);
or U3076 (N_3076,N_2936,N_2866);
or U3077 (N_3077,N_2874,N_2701);
nor U3078 (N_3078,N_2677,N_2986);
nor U3079 (N_3079,N_2722,N_2288);
nand U3080 (N_3080,N_2613,N_2497);
or U3081 (N_3081,N_2733,N_2575);
nand U3082 (N_3082,N_2484,N_2572);
or U3083 (N_3083,N_2837,N_2351);
and U3084 (N_3084,N_2523,N_2411);
or U3085 (N_3085,N_2328,N_2789);
and U3086 (N_3086,N_2703,N_2997);
nor U3087 (N_3087,N_2628,N_2971);
nand U3088 (N_3088,N_2504,N_2478);
nand U3089 (N_3089,N_2267,N_2686);
nand U3090 (N_3090,N_2508,N_2882);
nor U3091 (N_3091,N_2324,N_2516);
or U3092 (N_3092,N_2287,N_2394);
and U3093 (N_3093,N_2869,N_2346);
nor U3094 (N_3094,N_2639,N_2795);
or U3095 (N_3095,N_2522,N_2901);
and U3096 (N_3096,N_2923,N_2580);
and U3097 (N_3097,N_2859,N_2946);
or U3098 (N_3098,N_2458,N_2941);
nand U3099 (N_3099,N_2642,N_2855);
nor U3100 (N_3100,N_2537,N_2538);
nand U3101 (N_3101,N_2604,N_2407);
nand U3102 (N_3102,N_2565,N_2948);
nor U3103 (N_3103,N_2433,N_2299);
nor U3104 (N_3104,N_2597,N_2412);
and U3105 (N_3105,N_2329,N_2563);
and U3106 (N_3106,N_2761,N_2283);
xnor U3107 (N_3107,N_2577,N_2788);
nand U3108 (N_3108,N_2632,N_2263);
nor U3109 (N_3109,N_2985,N_2995);
and U3110 (N_3110,N_2935,N_2286);
nor U3111 (N_3111,N_2427,N_2596);
nor U3112 (N_3112,N_2425,N_2422);
xor U3113 (N_3113,N_2316,N_2943);
and U3114 (N_3114,N_2381,N_2962);
or U3115 (N_3115,N_2978,N_2831);
or U3116 (N_3116,N_2301,N_2270);
nand U3117 (N_3117,N_2920,N_2293);
and U3118 (N_3118,N_2559,N_2697);
and U3119 (N_3119,N_2681,N_2835);
and U3120 (N_3120,N_2454,N_2382);
and U3121 (N_3121,N_2700,N_2373);
nand U3122 (N_3122,N_2277,N_2496);
nand U3123 (N_3123,N_2800,N_2349);
nor U3124 (N_3124,N_2890,N_2546);
xnor U3125 (N_3125,N_2793,N_2261);
xnor U3126 (N_3126,N_2558,N_2836);
and U3127 (N_3127,N_2735,N_2250);
xor U3128 (N_3128,N_2913,N_2420);
and U3129 (N_3129,N_2327,N_2707);
nor U3130 (N_3130,N_2520,N_2476);
or U3131 (N_3131,N_2637,N_2445);
and U3132 (N_3132,N_2625,N_2939);
and U3133 (N_3133,N_2689,N_2335);
nor U3134 (N_3134,N_2358,N_2633);
and U3135 (N_3135,N_2524,N_2459);
xnor U3136 (N_3136,N_2341,N_2758);
or U3137 (N_3137,N_2611,N_2666);
xor U3138 (N_3138,N_2757,N_2464);
or U3139 (N_3139,N_2378,N_2470);
or U3140 (N_3140,N_2897,N_2282);
nor U3141 (N_3141,N_2397,N_2502);
xnor U3142 (N_3142,N_2715,N_2839);
and U3143 (N_3143,N_2822,N_2594);
or U3144 (N_3144,N_2291,N_2668);
nand U3145 (N_3145,N_2877,N_2810);
xnor U3146 (N_3146,N_2315,N_2258);
nand U3147 (N_3147,N_2851,N_2889);
nor U3148 (N_3148,N_2787,N_2881);
nor U3149 (N_3149,N_2384,N_2441);
xor U3150 (N_3150,N_2566,N_2739);
or U3151 (N_3151,N_2640,N_2507);
or U3152 (N_3152,N_2278,N_2547);
nand U3153 (N_3153,N_2706,N_2570);
or U3154 (N_3154,N_2969,N_2879);
or U3155 (N_3155,N_2654,N_2950);
nand U3156 (N_3156,N_2432,N_2992);
xor U3157 (N_3157,N_2799,N_2934);
nand U3158 (N_3158,N_2587,N_2850);
and U3159 (N_3159,N_2663,N_2457);
or U3160 (N_3160,N_2938,N_2506);
nor U3161 (N_3161,N_2904,N_2273);
nor U3162 (N_3162,N_2607,N_2498);
xnor U3163 (N_3163,N_2683,N_2262);
nand U3164 (N_3164,N_2958,N_2966);
nor U3165 (N_3165,N_2924,N_2489);
nor U3166 (N_3166,N_2721,N_2528);
nor U3167 (N_3167,N_2303,N_2356);
and U3168 (N_3168,N_2480,N_2571);
nor U3169 (N_3169,N_2386,N_2805);
nor U3170 (N_3170,N_2626,N_2624);
nand U3171 (N_3171,N_2759,N_2561);
or U3172 (N_3172,N_2437,N_2752);
or U3173 (N_3173,N_2495,N_2852);
and U3174 (N_3174,N_2276,N_2734);
nand U3175 (N_3175,N_2748,N_2847);
nand U3176 (N_3176,N_2511,N_2811);
and U3177 (N_3177,N_2854,N_2674);
nand U3178 (N_3178,N_2434,N_2766);
or U3179 (N_3179,N_2599,N_2945);
nand U3180 (N_3180,N_2929,N_2714);
and U3181 (N_3181,N_2695,N_2475);
and U3182 (N_3182,N_2781,N_2446);
nor U3183 (N_3183,N_2993,N_2670);
and U3184 (N_3184,N_2307,N_2991);
nor U3185 (N_3185,N_2331,N_2281);
and U3186 (N_3186,N_2403,N_2501);
nor U3187 (N_3187,N_2294,N_2645);
nor U3188 (N_3188,N_2774,N_2618);
and U3189 (N_3189,N_2399,N_2550);
and U3190 (N_3190,N_2780,N_2544);
nor U3191 (N_3191,N_2285,N_2926);
nand U3192 (N_3192,N_2251,N_2820);
and U3193 (N_3193,N_2452,N_2265);
and U3194 (N_3194,N_2914,N_2569);
or U3195 (N_3195,N_2728,N_2274);
or U3196 (N_3196,N_2909,N_2649);
and U3197 (N_3197,N_2843,N_2490);
nand U3198 (N_3198,N_2717,N_2823);
or U3199 (N_3199,N_2380,N_2483);
nor U3200 (N_3200,N_2777,N_2374);
or U3201 (N_3201,N_2363,N_2900);
nor U3202 (N_3202,N_2491,N_2702);
nor U3203 (N_3203,N_2529,N_2423);
and U3204 (N_3204,N_2369,N_2548);
nor U3205 (N_3205,N_2401,N_2279);
nand U3206 (N_3206,N_2469,N_2968);
or U3207 (N_3207,N_2512,N_2827);
or U3208 (N_3208,N_2796,N_2821);
nand U3209 (N_3209,N_2395,N_2982);
xnor U3210 (N_3210,N_2783,N_2584);
nand U3211 (N_3211,N_2305,N_2465);
or U3212 (N_3212,N_2614,N_2361);
xor U3213 (N_3213,N_2334,N_2818);
xor U3214 (N_3214,N_2590,N_2313);
nor U3215 (N_3215,N_2916,N_2699);
or U3216 (N_3216,N_2562,N_2268);
xor U3217 (N_3217,N_2573,N_2778);
or U3218 (N_3218,N_2848,N_2873);
and U3219 (N_3219,N_2937,N_2983);
and U3220 (N_3220,N_2804,N_2792);
and U3221 (N_3221,N_2449,N_2976);
and U3222 (N_3222,N_2712,N_2694);
and U3223 (N_3223,N_2797,N_2463);
xnor U3224 (N_3224,N_2864,N_2768);
nor U3225 (N_3225,N_2634,N_2436);
or U3226 (N_3226,N_2615,N_2947);
or U3227 (N_3227,N_2930,N_2767);
or U3228 (N_3228,N_2367,N_2542);
and U3229 (N_3229,N_2414,N_2485);
nand U3230 (N_3230,N_2364,N_2673);
or U3231 (N_3231,N_2798,N_2814);
nand U3232 (N_3232,N_2949,N_2310);
xor U3233 (N_3233,N_2892,N_2492);
and U3234 (N_3234,N_2664,N_2518);
nor U3235 (N_3235,N_2578,N_2311);
nor U3236 (N_3236,N_2692,N_2579);
nor U3237 (N_3237,N_2336,N_2429);
xnor U3238 (N_3238,N_2762,N_2672);
nor U3239 (N_3239,N_2252,N_2956);
and U3240 (N_3240,N_2545,N_2503);
and U3241 (N_3241,N_2534,N_2468);
and U3242 (N_3242,N_2906,N_2975);
and U3243 (N_3243,N_2908,N_2671);
or U3244 (N_3244,N_2899,N_2602);
nand U3245 (N_3245,N_2595,N_2760);
nand U3246 (N_3246,N_2643,N_2647);
nor U3247 (N_3247,N_2375,N_2260);
nand U3248 (N_3248,N_2255,N_2940);
or U3249 (N_3249,N_2586,N_2682);
and U3250 (N_3250,N_2853,N_2773);
nor U3251 (N_3251,N_2312,N_2998);
nand U3252 (N_3252,N_2257,N_2965);
nand U3253 (N_3253,N_2555,N_2517);
and U3254 (N_3254,N_2994,N_2355);
or U3255 (N_3255,N_2526,N_2844);
and U3256 (N_3256,N_2688,N_2641);
and U3257 (N_3257,N_2589,N_2297);
and U3258 (N_3258,N_2687,N_2605);
nor U3259 (N_3259,N_2564,N_2591);
nand U3260 (N_3260,N_2398,N_2379);
and U3261 (N_3261,N_2957,N_2424);
nand U3262 (N_3262,N_2340,N_2741);
xor U3263 (N_3263,N_2631,N_2627);
nand U3264 (N_3264,N_2505,N_2996);
and U3265 (N_3265,N_2619,N_2751);
nand U3266 (N_3266,N_2560,N_2488);
xor U3267 (N_3267,N_2858,N_2763);
or U3268 (N_3268,N_2782,N_2691);
and U3269 (N_3269,N_2754,N_2719);
nand U3270 (N_3270,N_2812,N_2418);
nor U3271 (N_3271,N_2461,N_2540);
or U3272 (N_3272,N_2284,N_2325);
nor U3273 (N_3273,N_2727,N_2466);
nand U3274 (N_3274,N_2330,N_2951);
or U3275 (N_3275,N_2984,N_2693);
and U3276 (N_3276,N_2657,N_2536);
or U3277 (N_3277,N_2343,N_2838);
nor U3278 (N_3278,N_2696,N_2430);
xnor U3279 (N_3279,N_2776,N_2659);
or U3280 (N_3280,N_2845,N_2959);
or U3281 (N_3281,N_2875,N_2658);
nand U3282 (N_3282,N_2973,N_2416);
and U3283 (N_3283,N_2616,N_2846);
nor U3284 (N_3284,N_2980,N_2306);
nand U3285 (N_3285,N_2833,N_2460);
nand U3286 (N_3286,N_2600,N_2431);
nand U3287 (N_3287,N_2738,N_2944);
and U3288 (N_3288,N_2413,N_2644);
nand U3289 (N_3289,N_2868,N_2857);
and U3290 (N_3290,N_2405,N_2442);
nand U3291 (N_3291,N_2462,N_2289);
xnor U3292 (N_3292,N_2878,N_2359);
or U3293 (N_3293,N_2576,N_2456);
and U3294 (N_3294,N_2718,N_2716);
or U3295 (N_3295,N_2598,N_2513);
nand U3296 (N_3296,N_2635,N_2606);
nand U3297 (N_3297,N_2585,N_2732);
nand U3298 (N_3298,N_2387,N_2651);
nand U3299 (N_3299,N_2592,N_2593);
nor U3300 (N_3300,N_2494,N_2519);
or U3301 (N_3301,N_2680,N_2360);
xor U3302 (N_3302,N_2802,N_2970);
or U3303 (N_3303,N_2824,N_2867);
xor U3304 (N_3304,N_2371,N_2972);
and U3305 (N_3305,N_2769,N_2309);
or U3306 (N_3306,N_2318,N_2736);
nor U3307 (N_3307,N_2832,N_2989);
and U3308 (N_3308,N_2509,N_2656);
nor U3309 (N_3309,N_2775,N_2690);
nand U3310 (N_3310,N_2352,N_2448);
nand U3311 (N_3311,N_2521,N_2828);
and U3312 (N_3312,N_2817,N_2296);
xnor U3313 (N_3313,N_2581,N_2964);
and U3314 (N_3314,N_2426,N_2493);
or U3315 (N_3315,N_2842,N_2272);
and U3316 (N_3316,N_2863,N_2539);
or U3317 (N_3317,N_2317,N_2922);
nand U3318 (N_3318,N_2410,N_2487);
xnor U3319 (N_3319,N_2322,N_2771);
nand U3320 (N_3320,N_2933,N_2834);
nand U3321 (N_3321,N_2357,N_2747);
nor U3322 (N_3322,N_2726,N_2326);
xor U3323 (N_3323,N_2902,N_2253);
and U3324 (N_3324,N_2794,N_2819);
xor U3325 (N_3325,N_2744,N_2510);
nand U3326 (N_3326,N_2678,N_2254);
xnor U3327 (N_3327,N_2530,N_2525);
or U3328 (N_3328,N_2898,N_2515);
and U3329 (N_3329,N_2685,N_2806);
xor U3330 (N_3330,N_2860,N_2447);
and U3331 (N_3331,N_2302,N_2675);
and U3332 (N_3332,N_2323,N_2636);
and U3333 (N_3333,N_2895,N_2887);
and U3334 (N_3334,N_2967,N_2500);
nand U3335 (N_3335,N_2765,N_2891);
nand U3336 (N_3336,N_2612,N_2883);
or U3337 (N_3337,N_2709,N_2684);
or U3338 (N_3338,N_2919,N_2910);
nor U3339 (N_3339,N_2955,N_2350);
nor U3340 (N_3340,N_2630,N_2912);
nand U3341 (N_3341,N_2269,N_2665);
xor U3342 (N_3342,N_2705,N_2321);
and U3343 (N_3343,N_2337,N_2629);
and U3344 (N_3344,N_2840,N_2266);
or U3345 (N_3345,N_2608,N_2679);
nor U3346 (N_3346,N_2366,N_2931);
nor U3347 (N_3347,N_2259,N_2779);
or U3348 (N_3348,N_2770,N_2609);
and U3349 (N_3349,N_2532,N_2884);
or U3350 (N_3350,N_2347,N_2737);
nor U3351 (N_3351,N_2354,N_2396);
nand U3352 (N_3352,N_2362,N_2583);
nand U3353 (N_3353,N_2979,N_2729);
and U3354 (N_3354,N_2264,N_2455);
or U3355 (N_3355,N_2927,N_2870);
nor U3356 (N_3356,N_2365,N_2417);
and U3357 (N_3357,N_2960,N_2482);
xor U3358 (N_3358,N_2400,N_2541);
or U3359 (N_3359,N_2815,N_2662);
nor U3360 (N_3360,N_2621,N_2342);
nand U3361 (N_3361,N_2646,N_2344);
xor U3362 (N_3362,N_2308,N_2749);
nand U3363 (N_3363,N_2471,N_2439);
nand U3364 (N_3364,N_2450,N_2915);
nand U3365 (N_3365,N_2725,N_2784);
and U3366 (N_3366,N_2353,N_2440);
nor U3367 (N_3367,N_2711,N_2723);
nor U3368 (N_3368,N_2385,N_2743);
or U3369 (N_3369,N_2391,N_2392);
nor U3370 (N_3370,N_2304,N_2543);
nor U3371 (N_3371,N_2295,N_2388);
xnor U3372 (N_3372,N_2320,N_2990);
and U3373 (N_3373,N_2954,N_2952);
nand U3374 (N_3374,N_2376,N_2652);
nand U3375 (N_3375,N_2525,N_2859);
xnor U3376 (N_3376,N_2952,N_2518);
nand U3377 (N_3377,N_2487,N_2964);
or U3378 (N_3378,N_2796,N_2845);
nand U3379 (N_3379,N_2399,N_2614);
or U3380 (N_3380,N_2419,N_2428);
nor U3381 (N_3381,N_2992,N_2708);
or U3382 (N_3382,N_2866,N_2784);
nor U3383 (N_3383,N_2942,N_2731);
and U3384 (N_3384,N_2917,N_2653);
or U3385 (N_3385,N_2871,N_2291);
nor U3386 (N_3386,N_2597,N_2898);
or U3387 (N_3387,N_2670,N_2465);
and U3388 (N_3388,N_2767,N_2692);
or U3389 (N_3389,N_2502,N_2986);
nand U3390 (N_3390,N_2576,N_2677);
nor U3391 (N_3391,N_2742,N_2508);
nand U3392 (N_3392,N_2668,N_2852);
or U3393 (N_3393,N_2644,N_2845);
and U3394 (N_3394,N_2985,N_2455);
nand U3395 (N_3395,N_2604,N_2697);
nor U3396 (N_3396,N_2895,N_2905);
and U3397 (N_3397,N_2670,N_2963);
nor U3398 (N_3398,N_2625,N_2311);
and U3399 (N_3399,N_2827,N_2306);
and U3400 (N_3400,N_2671,N_2718);
nor U3401 (N_3401,N_2956,N_2625);
or U3402 (N_3402,N_2455,N_2662);
and U3403 (N_3403,N_2437,N_2351);
and U3404 (N_3404,N_2716,N_2903);
nand U3405 (N_3405,N_2322,N_2856);
nand U3406 (N_3406,N_2581,N_2830);
nand U3407 (N_3407,N_2679,N_2396);
nand U3408 (N_3408,N_2447,N_2561);
and U3409 (N_3409,N_2261,N_2739);
and U3410 (N_3410,N_2753,N_2840);
nand U3411 (N_3411,N_2905,N_2662);
nor U3412 (N_3412,N_2837,N_2543);
or U3413 (N_3413,N_2496,N_2262);
and U3414 (N_3414,N_2978,N_2416);
and U3415 (N_3415,N_2880,N_2642);
nor U3416 (N_3416,N_2698,N_2875);
xnor U3417 (N_3417,N_2818,N_2411);
nor U3418 (N_3418,N_2622,N_2401);
nor U3419 (N_3419,N_2481,N_2276);
nand U3420 (N_3420,N_2955,N_2394);
nand U3421 (N_3421,N_2537,N_2753);
and U3422 (N_3422,N_2895,N_2607);
nand U3423 (N_3423,N_2868,N_2734);
or U3424 (N_3424,N_2781,N_2595);
nand U3425 (N_3425,N_2950,N_2250);
or U3426 (N_3426,N_2826,N_2304);
and U3427 (N_3427,N_2983,N_2791);
nor U3428 (N_3428,N_2341,N_2400);
or U3429 (N_3429,N_2819,N_2708);
nor U3430 (N_3430,N_2670,N_2291);
xnor U3431 (N_3431,N_2777,N_2311);
nor U3432 (N_3432,N_2330,N_2623);
nand U3433 (N_3433,N_2349,N_2575);
and U3434 (N_3434,N_2828,N_2614);
and U3435 (N_3435,N_2488,N_2809);
nand U3436 (N_3436,N_2943,N_2551);
or U3437 (N_3437,N_2357,N_2381);
nor U3438 (N_3438,N_2970,N_2529);
or U3439 (N_3439,N_2810,N_2421);
or U3440 (N_3440,N_2585,N_2367);
or U3441 (N_3441,N_2877,N_2273);
xnor U3442 (N_3442,N_2562,N_2593);
nor U3443 (N_3443,N_2452,N_2709);
nor U3444 (N_3444,N_2395,N_2505);
and U3445 (N_3445,N_2699,N_2876);
nand U3446 (N_3446,N_2268,N_2528);
or U3447 (N_3447,N_2600,N_2433);
and U3448 (N_3448,N_2540,N_2558);
nor U3449 (N_3449,N_2939,N_2450);
nor U3450 (N_3450,N_2420,N_2719);
and U3451 (N_3451,N_2680,N_2585);
and U3452 (N_3452,N_2606,N_2384);
nor U3453 (N_3453,N_2824,N_2596);
nor U3454 (N_3454,N_2289,N_2336);
and U3455 (N_3455,N_2401,N_2599);
nand U3456 (N_3456,N_2580,N_2416);
or U3457 (N_3457,N_2583,N_2833);
nand U3458 (N_3458,N_2287,N_2467);
or U3459 (N_3459,N_2750,N_2522);
or U3460 (N_3460,N_2999,N_2555);
nor U3461 (N_3461,N_2909,N_2761);
xor U3462 (N_3462,N_2787,N_2595);
nand U3463 (N_3463,N_2789,N_2623);
or U3464 (N_3464,N_2611,N_2894);
or U3465 (N_3465,N_2650,N_2912);
and U3466 (N_3466,N_2300,N_2926);
nand U3467 (N_3467,N_2276,N_2255);
xnor U3468 (N_3468,N_2346,N_2870);
and U3469 (N_3469,N_2513,N_2600);
nand U3470 (N_3470,N_2408,N_2949);
or U3471 (N_3471,N_2969,N_2920);
nor U3472 (N_3472,N_2646,N_2355);
or U3473 (N_3473,N_2887,N_2828);
xnor U3474 (N_3474,N_2549,N_2904);
nand U3475 (N_3475,N_2904,N_2552);
nand U3476 (N_3476,N_2290,N_2785);
or U3477 (N_3477,N_2644,N_2981);
or U3478 (N_3478,N_2893,N_2943);
and U3479 (N_3479,N_2280,N_2674);
and U3480 (N_3480,N_2348,N_2781);
and U3481 (N_3481,N_2374,N_2700);
or U3482 (N_3482,N_2632,N_2636);
or U3483 (N_3483,N_2873,N_2258);
nor U3484 (N_3484,N_2693,N_2413);
and U3485 (N_3485,N_2752,N_2813);
xor U3486 (N_3486,N_2820,N_2278);
and U3487 (N_3487,N_2905,N_2816);
nand U3488 (N_3488,N_2984,N_2720);
nor U3489 (N_3489,N_2940,N_2301);
nand U3490 (N_3490,N_2773,N_2987);
or U3491 (N_3491,N_2315,N_2707);
and U3492 (N_3492,N_2416,N_2661);
nand U3493 (N_3493,N_2321,N_2338);
nand U3494 (N_3494,N_2345,N_2886);
nand U3495 (N_3495,N_2724,N_2729);
and U3496 (N_3496,N_2272,N_2971);
nand U3497 (N_3497,N_2586,N_2360);
xor U3498 (N_3498,N_2429,N_2829);
nor U3499 (N_3499,N_2696,N_2613);
xnor U3500 (N_3500,N_2865,N_2321);
and U3501 (N_3501,N_2379,N_2836);
and U3502 (N_3502,N_2884,N_2644);
nor U3503 (N_3503,N_2602,N_2503);
nand U3504 (N_3504,N_2723,N_2781);
nor U3505 (N_3505,N_2764,N_2423);
and U3506 (N_3506,N_2950,N_2878);
nor U3507 (N_3507,N_2578,N_2435);
nor U3508 (N_3508,N_2520,N_2536);
and U3509 (N_3509,N_2870,N_2985);
and U3510 (N_3510,N_2492,N_2845);
or U3511 (N_3511,N_2689,N_2846);
nor U3512 (N_3512,N_2939,N_2712);
and U3513 (N_3513,N_2380,N_2553);
and U3514 (N_3514,N_2417,N_2707);
and U3515 (N_3515,N_2332,N_2435);
or U3516 (N_3516,N_2871,N_2608);
nor U3517 (N_3517,N_2628,N_2297);
nor U3518 (N_3518,N_2852,N_2475);
nand U3519 (N_3519,N_2780,N_2363);
or U3520 (N_3520,N_2798,N_2533);
and U3521 (N_3521,N_2938,N_2562);
and U3522 (N_3522,N_2297,N_2911);
nand U3523 (N_3523,N_2633,N_2695);
nand U3524 (N_3524,N_2670,N_2524);
nand U3525 (N_3525,N_2712,N_2790);
nor U3526 (N_3526,N_2797,N_2565);
and U3527 (N_3527,N_2688,N_2394);
or U3528 (N_3528,N_2434,N_2762);
nand U3529 (N_3529,N_2918,N_2445);
nand U3530 (N_3530,N_2335,N_2697);
and U3531 (N_3531,N_2359,N_2627);
nand U3532 (N_3532,N_2684,N_2986);
and U3533 (N_3533,N_2638,N_2456);
nor U3534 (N_3534,N_2716,N_2498);
or U3535 (N_3535,N_2415,N_2395);
and U3536 (N_3536,N_2641,N_2561);
xnor U3537 (N_3537,N_2951,N_2746);
and U3538 (N_3538,N_2530,N_2352);
and U3539 (N_3539,N_2871,N_2414);
nor U3540 (N_3540,N_2467,N_2823);
and U3541 (N_3541,N_2364,N_2344);
and U3542 (N_3542,N_2255,N_2648);
nand U3543 (N_3543,N_2607,N_2660);
nand U3544 (N_3544,N_2723,N_2726);
and U3545 (N_3545,N_2684,N_2544);
nor U3546 (N_3546,N_2277,N_2781);
nand U3547 (N_3547,N_2764,N_2481);
or U3548 (N_3548,N_2558,N_2276);
and U3549 (N_3549,N_2671,N_2509);
or U3550 (N_3550,N_2443,N_2585);
and U3551 (N_3551,N_2519,N_2884);
or U3552 (N_3552,N_2643,N_2925);
xor U3553 (N_3553,N_2671,N_2754);
and U3554 (N_3554,N_2795,N_2643);
and U3555 (N_3555,N_2924,N_2648);
or U3556 (N_3556,N_2755,N_2459);
nor U3557 (N_3557,N_2662,N_2512);
or U3558 (N_3558,N_2905,N_2540);
xor U3559 (N_3559,N_2873,N_2944);
nand U3560 (N_3560,N_2469,N_2335);
xnor U3561 (N_3561,N_2336,N_2656);
or U3562 (N_3562,N_2735,N_2837);
xor U3563 (N_3563,N_2921,N_2987);
nor U3564 (N_3564,N_2878,N_2768);
xnor U3565 (N_3565,N_2429,N_2756);
or U3566 (N_3566,N_2770,N_2305);
and U3567 (N_3567,N_2281,N_2887);
or U3568 (N_3568,N_2757,N_2528);
or U3569 (N_3569,N_2839,N_2302);
and U3570 (N_3570,N_2753,N_2345);
xor U3571 (N_3571,N_2615,N_2271);
and U3572 (N_3572,N_2278,N_2654);
or U3573 (N_3573,N_2477,N_2415);
nand U3574 (N_3574,N_2582,N_2508);
nand U3575 (N_3575,N_2867,N_2268);
and U3576 (N_3576,N_2863,N_2625);
and U3577 (N_3577,N_2529,N_2430);
and U3578 (N_3578,N_2937,N_2710);
nand U3579 (N_3579,N_2573,N_2843);
or U3580 (N_3580,N_2788,N_2931);
or U3581 (N_3581,N_2736,N_2519);
nand U3582 (N_3582,N_2473,N_2983);
nor U3583 (N_3583,N_2407,N_2533);
or U3584 (N_3584,N_2777,N_2630);
or U3585 (N_3585,N_2929,N_2888);
nand U3586 (N_3586,N_2801,N_2856);
nand U3587 (N_3587,N_2660,N_2681);
nand U3588 (N_3588,N_2412,N_2715);
xnor U3589 (N_3589,N_2802,N_2585);
or U3590 (N_3590,N_2920,N_2545);
and U3591 (N_3591,N_2902,N_2970);
xor U3592 (N_3592,N_2754,N_2741);
or U3593 (N_3593,N_2625,N_2698);
xor U3594 (N_3594,N_2342,N_2937);
nor U3595 (N_3595,N_2323,N_2303);
and U3596 (N_3596,N_2265,N_2529);
nand U3597 (N_3597,N_2770,N_2461);
nand U3598 (N_3598,N_2724,N_2971);
nand U3599 (N_3599,N_2751,N_2496);
nor U3600 (N_3600,N_2410,N_2799);
nor U3601 (N_3601,N_2988,N_2477);
nor U3602 (N_3602,N_2473,N_2566);
nand U3603 (N_3603,N_2431,N_2797);
xor U3604 (N_3604,N_2570,N_2640);
or U3605 (N_3605,N_2592,N_2498);
and U3606 (N_3606,N_2959,N_2923);
nand U3607 (N_3607,N_2728,N_2944);
and U3608 (N_3608,N_2267,N_2649);
nand U3609 (N_3609,N_2841,N_2998);
xnor U3610 (N_3610,N_2715,N_2922);
nand U3611 (N_3611,N_2511,N_2495);
and U3612 (N_3612,N_2540,N_2857);
and U3613 (N_3613,N_2644,N_2840);
nor U3614 (N_3614,N_2594,N_2679);
or U3615 (N_3615,N_2832,N_2279);
nand U3616 (N_3616,N_2980,N_2383);
xnor U3617 (N_3617,N_2438,N_2603);
nor U3618 (N_3618,N_2595,N_2274);
xnor U3619 (N_3619,N_2581,N_2842);
and U3620 (N_3620,N_2510,N_2375);
nor U3621 (N_3621,N_2522,N_2257);
and U3622 (N_3622,N_2533,N_2461);
nor U3623 (N_3623,N_2370,N_2553);
xor U3624 (N_3624,N_2565,N_2496);
nor U3625 (N_3625,N_2769,N_2458);
nand U3626 (N_3626,N_2428,N_2329);
nor U3627 (N_3627,N_2800,N_2771);
nand U3628 (N_3628,N_2812,N_2698);
nand U3629 (N_3629,N_2856,N_2987);
nand U3630 (N_3630,N_2877,N_2448);
and U3631 (N_3631,N_2807,N_2495);
and U3632 (N_3632,N_2786,N_2872);
xor U3633 (N_3633,N_2797,N_2635);
or U3634 (N_3634,N_2740,N_2361);
nand U3635 (N_3635,N_2515,N_2946);
and U3636 (N_3636,N_2765,N_2307);
and U3637 (N_3637,N_2843,N_2789);
nor U3638 (N_3638,N_2393,N_2564);
nor U3639 (N_3639,N_2643,N_2873);
nor U3640 (N_3640,N_2793,N_2311);
xnor U3641 (N_3641,N_2937,N_2300);
or U3642 (N_3642,N_2743,N_2311);
xor U3643 (N_3643,N_2447,N_2490);
nand U3644 (N_3644,N_2761,N_2335);
or U3645 (N_3645,N_2378,N_2589);
nor U3646 (N_3646,N_2898,N_2421);
xor U3647 (N_3647,N_2673,N_2510);
nor U3648 (N_3648,N_2780,N_2990);
nor U3649 (N_3649,N_2251,N_2625);
nor U3650 (N_3650,N_2573,N_2920);
and U3651 (N_3651,N_2595,N_2802);
nand U3652 (N_3652,N_2308,N_2547);
nand U3653 (N_3653,N_2699,N_2704);
and U3654 (N_3654,N_2558,N_2768);
xnor U3655 (N_3655,N_2571,N_2338);
nand U3656 (N_3656,N_2611,N_2299);
nor U3657 (N_3657,N_2852,N_2614);
xor U3658 (N_3658,N_2543,N_2801);
nor U3659 (N_3659,N_2976,N_2746);
nor U3660 (N_3660,N_2533,N_2715);
xor U3661 (N_3661,N_2746,N_2318);
xor U3662 (N_3662,N_2735,N_2908);
nor U3663 (N_3663,N_2733,N_2418);
or U3664 (N_3664,N_2515,N_2475);
or U3665 (N_3665,N_2815,N_2935);
and U3666 (N_3666,N_2890,N_2654);
or U3667 (N_3667,N_2956,N_2873);
xor U3668 (N_3668,N_2997,N_2497);
nor U3669 (N_3669,N_2367,N_2712);
nor U3670 (N_3670,N_2819,N_2681);
or U3671 (N_3671,N_2306,N_2722);
or U3672 (N_3672,N_2471,N_2618);
nor U3673 (N_3673,N_2780,N_2619);
and U3674 (N_3674,N_2324,N_2878);
nand U3675 (N_3675,N_2882,N_2370);
or U3676 (N_3676,N_2624,N_2858);
nor U3677 (N_3677,N_2921,N_2717);
nand U3678 (N_3678,N_2867,N_2601);
nor U3679 (N_3679,N_2394,N_2823);
nor U3680 (N_3680,N_2671,N_2929);
nand U3681 (N_3681,N_2703,N_2636);
and U3682 (N_3682,N_2597,N_2796);
nand U3683 (N_3683,N_2927,N_2553);
or U3684 (N_3684,N_2564,N_2855);
and U3685 (N_3685,N_2910,N_2789);
and U3686 (N_3686,N_2461,N_2969);
xnor U3687 (N_3687,N_2504,N_2790);
or U3688 (N_3688,N_2807,N_2259);
nand U3689 (N_3689,N_2669,N_2704);
and U3690 (N_3690,N_2821,N_2489);
nand U3691 (N_3691,N_2909,N_2568);
nand U3692 (N_3692,N_2580,N_2502);
and U3693 (N_3693,N_2825,N_2696);
or U3694 (N_3694,N_2318,N_2827);
or U3695 (N_3695,N_2993,N_2399);
nand U3696 (N_3696,N_2603,N_2588);
and U3697 (N_3697,N_2262,N_2417);
or U3698 (N_3698,N_2675,N_2591);
nor U3699 (N_3699,N_2508,N_2335);
nor U3700 (N_3700,N_2701,N_2934);
or U3701 (N_3701,N_2925,N_2806);
nand U3702 (N_3702,N_2366,N_2993);
nand U3703 (N_3703,N_2463,N_2810);
nand U3704 (N_3704,N_2761,N_2768);
nand U3705 (N_3705,N_2793,N_2636);
and U3706 (N_3706,N_2715,N_2455);
or U3707 (N_3707,N_2423,N_2728);
nor U3708 (N_3708,N_2761,N_2679);
nand U3709 (N_3709,N_2418,N_2335);
and U3710 (N_3710,N_2356,N_2275);
nor U3711 (N_3711,N_2775,N_2966);
nand U3712 (N_3712,N_2313,N_2342);
nor U3713 (N_3713,N_2446,N_2429);
nor U3714 (N_3714,N_2856,N_2686);
nor U3715 (N_3715,N_2469,N_2389);
nand U3716 (N_3716,N_2945,N_2571);
nand U3717 (N_3717,N_2940,N_2314);
and U3718 (N_3718,N_2620,N_2366);
nand U3719 (N_3719,N_2330,N_2943);
nor U3720 (N_3720,N_2611,N_2548);
or U3721 (N_3721,N_2497,N_2853);
and U3722 (N_3722,N_2989,N_2507);
nand U3723 (N_3723,N_2345,N_2698);
and U3724 (N_3724,N_2869,N_2659);
nor U3725 (N_3725,N_2865,N_2540);
xor U3726 (N_3726,N_2320,N_2515);
nor U3727 (N_3727,N_2803,N_2555);
nor U3728 (N_3728,N_2445,N_2538);
nor U3729 (N_3729,N_2436,N_2838);
nand U3730 (N_3730,N_2550,N_2764);
and U3731 (N_3731,N_2670,N_2643);
nor U3732 (N_3732,N_2943,N_2714);
nand U3733 (N_3733,N_2446,N_2951);
nor U3734 (N_3734,N_2970,N_2264);
or U3735 (N_3735,N_2844,N_2728);
nand U3736 (N_3736,N_2414,N_2947);
xor U3737 (N_3737,N_2518,N_2626);
xor U3738 (N_3738,N_2611,N_2873);
nand U3739 (N_3739,N_2856,N_2334);
nand U3740 (N_3740,N_2596,N_2684);
nand U3741 (N_3741,N_2637,N_2662);
or U3742 (N_3742,N_2888,N_2454);
or U3743 (N_3743,N_2390,N_2405);
xor U3744 (N_3744,N_2992,N_2902);
nand U3745 (N_3745,N_2934,N_2862);
xor U3746 (N_3746,N_2978,N_2680);
or U3747 (N_3747,N_2250,N_2853);
and U3748 (N_3748,N_2407,N_2852);
nand U3749 (N_3749,N_2446,N_2614);
nor U3750 (N_3750,N_3410,N_3240);
nor U3751 (N_3751,N_3309,N_3275);
and U3752 (N_3752,N_3617,N_3610);
or U3753 (N_3753,N_3312,N_3431);
or U3754 (N_3754,N_3384,N_3007);
nor U3755 (N_3755,N_3698,N_3360);
nand U3756 (N_3756,N_3140,N_3644);
nor U3757 (N_3757,N_3485,N_3719);
nor U3758 (N_3758,N_3073,N_3271);
or U3759 (N_3759,N_3123,N_3266);
or U3760 (N_3760,N_3629,N_3533);
xnor U3761 (N_3761,N_3233,N_3161);
nand U3762 (N_3762,N_3506,N_3110);
and U3763 (N_3763,N_3707,N_3370);
nand U3764 (N_3764,N_3491,N_3395);
nand U3765 (N_3765,N_3224,N_3056);
nor U3766 (N_3766,N_3427,N_3501);
and U3767 (N_3767,N_3339,N_3657);
and U3768 (N_3768,N_3613,N_3471);
nor U3769 (N_3769,N_3174,N_3682);
nor U3770 (N_3770,N_3705,N_3516);
nand U3771 (N_3771,N_3413,N_3421);
and U3772 (N_3772,N_3648,N_3594);
or U3773 (N_3773,N_3615,N_3653);
nor U3774 (N_3774,N_3397,N_3428);
nand U3775 (N_3775,N_3608,N_3106);
and U3776 (N_3776,N_3026,N_3122);
or U3777 (N_3777,N_3261,N_3481);
and U3778 (N_3778,N_3320,N_3507);
nand U3779 (N_3779,N_3453,N_3213);
nand U3780 (N_3780,N_3155,N_3674);
or U3781 (N_3781,N_3251,N_3659);
and U3782 (N_3782,N_3469,N_3628);
or U3783 (N_3783,N_3005,N_3163);
nand U3784 (N_3784,N_3525,N_3204);
or U3785 (N_3785,N_3607,N_3323);
nand U3786 (N_3786,N_3228,N_3189);
nor U3787 (N_3787,N_3436,N_3372);
xnor U3788 (N_3788,N_3134,N_3717);
or U3789 (N_3789,N_3555,N_3447);
or U3790 (N_3790,N_3253,N_3250);
and U3791 (N_3791,N_3351,N_3742);
nand U3792 (N_3792,N_3350,N_3563);
and U3793 (N_3793,N_3722,N_3346);
nand U3794 (N_3794,N_3268,N_3336);
nand U3795 (N_3795,N_3544,N_3182);
nand U3796 (N_3796,N_3435,N_3050);
nor U3797 (N_3797,N_3637,N_3284);
nand U3798 (N_3798,N_3201,N_3197);
nand U3799 (N_3799,N_3243,N_3553);
and U3800 (N_3800,N_3656,N_3241);
or U3801 (N_3801,N_3439,N_3500);
nor U3802 (N_3802,N_3156,N_3044);
nor U3803 (N_3803,N_3297,N_3735);
nor U3804 (N_3804,N_3053,N_3668);
and U3805 (N_3805,N_3542,N_3290);
nand U3806 (N_3806,N_3432,N_3305);
nand U3807 (N_3807,N_3649,N_3072);
and U3808 (N_3808,N_3064,N_3217);
and U3809 (N_3809,N_3216,N_3557);
nand U3810 (N_3810,N_3714,N_3687);
or U3811 (N_3811,N_3311,N_3573);
or U3812 (N_3812,N_3504,N_3522);
nand U3813 (N_3813,N_3405,N_3493);
nor U3814 (N_3814,N_3164,N_3376);
or U3815 (N_3815,N_3101,N_3411);
nor U3816 (N_3816,N_3468,N_3715);
and U3817 (N_3817,N_3445,N_3743);
nor U3818 (N_3818,N_3424,N_3593);
or U3819 (N_3819,N_3527,N_3093);
or U3820 (N_3820,N_3621,N_3636);
xnor U3821 (N_3821,N_3001,N_3294);
nor U3822 (N_3822,N_3448,N_3429);
nor U3823 (N_3823,N_3186,N_3623);
nand U3824 (N_3824,N_3135,N_3178);
nor U3825 (N_3825,N_3498,N_3388);
nor U3826 (N_3826,N_3539,N_3704);
and U3827 (N_3827,N_3142,N_3206);
or U3828 (N_3828,N_3152,N_3622);
and U3829 (N_3829,N_3080,N_3234);
and U3830 (N_3830,N_3661,N_3298);
nand U3831 (N_3831,N_3729,N_3558);
xnor U3832 (N_3832,N_3632,N_3132);
nand U3833 (N_3833,N_3173,N_3630);
and U3834 (N_3834,N_3166,N_3451);
and U3835 (N_3835,N_3701,N_3190);
and U3836 (N_3836,N_3015,N_3489);
nor U3837 (N_3837,N_3685,N_3292);
or U3838 (N_3838,N_3212,N_3639);
or U3839 (N_3839,N_3191,N_3452);
and U3840 (N_3840,N_3497,N_3325);
nand U3841 (N_3841,N_3300,N_3060);
nand U3842 (N_3842,N_3199,N_3078);
nor U3843 (N_3843,N_3529,N_3022);
and U3844 (N_3844,N_3021,N_3124);
xnor U3845 (N_3845,N_3009,N_3256);
nor U3846 (N_3846,N_3265,N_3499);
or U3847 (N_3847,N_3214,N_3567);
xor U3848 (N_3848,N_3699,N_3318);
nand U3849 (N_3849,N_3274,N_3449);
and U3850 (N_3850,N_3666,N_3535);
nand U3851 (N_3851,N_3128,N_3381);
or U3852 (N_3852,N_3695,N_3727);
and U3853 (N_3853,N_3720,N_3654);
nor U3854 (N_3854,N_3117,N_3277);
nor U3855 (N_3855,N_3721,N_3091);
nor U3856 (N_3856,N_3480,N_3517);
nor U3857 (N_3857,N_3012,N_3476);
nand U3858 (N_3858,N_3550,N_3502);
and U3859 (N_3859,N_3726,N_3619);
nor U3860 (N_3860,N_3092,N_3340);
xor U3861 (N_3861,N_3287,N_3108);
or U3862 (N_3862,N_3678,N_3177);
xor U3863 (N_3863,N_3129,N_3194);
nor U3864 (N_3864,N_3738,N_3231);
and U3865 (N_3865,N_3307,N_3138);
nor U3866 (N_3866,N_3441,N_3303);
nor U3867 (N_3867,N_3126,N_3302);
nand U3868 (N_3868,N_3331,N_3183);
nand U3869 (N_3869,N_3562,N_3670);
and U3870 (N_3870,N_3207,N_3523);
and U3871 (N_3871,N_3185,N_3119);
nor U3872 (N_3872,N_3412,N_3568);
nand U3873 (N_3873,N_3358,N_3546);
nand U3874 (N_3874,N_3446,N_3223);
or U3875 (N_3875,N_3642,N_3521);
or U3876 (N_3876,N_3540,N_3220);
or U3877 (N_3877,N_3671,N_3099);
and U3878 (N_3878,N_3159,N_3390);
and U3879 (N_3879,N_3130,N_3455);
and U3880 (N_3880,N_3039,N_3378);
xor U3881 (N_3881,N_3114,N_3105);
and U3882 (N_3882,N_3062,N_3651);
nor U3883 (N_3883,N_3087,N_3401);
or U3884 (N_3884,N_3181,N_3723);
nand U3885 (N_3885,N_3097,N_3147);
xnor U3886 (N_3886,N_3104,N_3718);
nand U3887 (N_3887,N_3706,N_3153);
or U3888 (N_3888,N_3203,N_3647);
and U3889 (N_3889,N_3641,N_3690);
or U3890 (N_3890,N_3430,N_3334);
nand U3891 (N_3891,N_3712,N_3450);
or U3892 (N_3892,N_3675,N_3133);
or U3893 (N_3893,N_3248,N_3590);
and U3894 (N_3894,N_3308,N_3505);
or U3895 (N_3895,N_3329,N_3354);
nor U3896 (N_3896,N_3272,N_3575);
and U3897 (N_3897,N_3548,N_3245);
nor U3898 (N_3898,N_3198,N_3025);
or U3899 (N_3899,N_3088,N_3470);
nand U3900 (N_3900,N_3328,N_3638);
or U3901 (N_3901,N_3175,N_3014);
and U3902 (N_3902,N_3255,N_3582);
or U3903 (N_3903,N_3089,N_3084);
and U3904 (N_3904,N_3725,N_3258);
and U3905 (N_3905,N_3416,N_3565);
and U3906 (N_3906,N_3232,N_3662);
nor U3907 (N_3907,N_3635,N_3665);
xnor U3908 (N_3908,N_3038,N_3676);
nor U3909 (N_3909,N_3225,N_3150);
xnor U3910 (N_3910,N_3193,N_3195);
nand U3911 (N_3911,N_3680,N_3210);
nand U3912 (N_3912,N_3343,N_3244);
or U3913 (N_3913,N_3076,N_3111);
or U3914 (N_3914,N_3222,N_3338);
xnor U3915 (N_3915,N_3154,N_3096);
or U3916 (N_3916,N_3603,N_3566);
and U3917 (N_3917,N_3696,N_3167);
or U3918 (N_3918,N_3741,N_3364);
or U3919 (N_3919,N_3465,N_3059);
nand U3920 (N_3920,N_3561,N_3393);
nor U3921 (N_3921,N_3426,N_3528);
and U3922 (N_3922,N_3524,N_3235);
nor U3923 (N_3923,N_3409,N_3747);
and U3924 (N_3924,N_3691,N_3033);
nor U3925 (N_3925,N_3732,N_3158);
nor U3926 (N_3926,N_3047,N_3374);
and U3927 (N_3927,N_3010,N_3279);
or U3928 (N_3928,N_3464,N_3180);
nor U3929 (N_3929,N_3503,N_3285);
or U3930 (N_3930,N_3237,N_3380);
nor U3931 (N_3931,N_3040,N_3744);
xnor U3932 (N_3932,N_3536,N_3655);
nor U3933 (N_3933,N_3236,N_3107);
nor U3934 (N_3934,N_3095,N_3556);
and U3935 (N_3935,N_3100,N_3362);
nor U3936 (N_3936,N_3389,N_3160);
and U3937 (N_3937,N_3466,N_3745);
nor U3938 (N_3938,N_3137,N_3440);
nand U3939 (N_3939,N_3459,N_3348);
or U3940 (N_3940,N_3202,N_3580);
or U3941 (N_3941,N_3366,N_3734);
xor U3942 (N_3942,N_3016,N_3422);
or U3943 (N_3943,N_3423,N_3564);
nand U3944 (N_3944,N_3710,N_3547);
and U3945 (N_3945,N_3262,N_3631);
and U3946 (N_3946,N_3693,N_3136);
and U3947 (N_3947,N_3205,N_3515);
nor U3948 (N_3948,N_3359,N_3403);
nand U3949 (N_3949,N_3460,N_3490);
nand U3950 (N_3950,N_3419,N_3252);
or U3951 (N_3951,N_3383,N_3749);
and U3952 (N_3952,N_3103,N_3672);
and U3953 (N_3953,N_3187,N_3008);
nand U3954 (N_3954,N_3643,N_3571);
nand U3955 (N_3955,N_3218,N_3263);
or U3956 (N_3956,N_3116,N_3322);
nor U3957 (N_3957,N_3518,N_3249);
nor U3958 (N_3958,N_3283,N_3512);
nand U3959 (N_3959,N_3043,N_3296);
or U3960 (N_3960,N_3162,N_3363);
nor U3961 (N_3961,N_3335,N_3125);
nor U3962 (N_3962,N_3463,N_3314);
nor U3963 (N_3963,N_3400,N_3355);
and U3964 (N_3964,N_3686,N_3260);
and U3965 (N_3965,N_3420,N_3324);
nand U3966 (N_3966,N_3418,N_3549);
nor U3967 (N_3967,N_3579,N_3317);
or U3968 (N_3968,N_3127,N_3634);
nor U3969 (N_3969,N_3006,N_3011);
nor U3970 (N_3970,N_3559,N_3310);
or U3971 (N_3971,N_3581,N_3077);
and U3972 (N_3972,N_3013,N_3074);
nor U3973 (N_3973,N_3692,N_3315);
nand U3974 (N_3974,N_3066,N_3192);
or U3975 (N_3975,N_3588,N_3612);
xnor U3976 (N_3976,N_3746,N_3673);
or U3977 (N_3977,N_3572,N_3689);
nor U3978 (N_3978,N_3085,N_3281);
and U3979 (N_3979,N_3375,N_3716);
nor U3980 (N_3980,N_3650,N_3034);
or U3981 (N_3981,N_3483,N_3530);
nand U3982 (N_3982,N_3369,N_3456);
or U3983 (N_3983,N_3221,N_3728);
or U3984 (N_3984,N_3569,N_3477);
and U3985 (N_3985,N_3414,N_3278);
nor U3986 (N_3986,N_3652,N_3392);
xor U3987 (N_3987,N_3574,N_3098);
nand U3988 (N_3988,N_3645,N_3664);
xnor U3989 (N_3989,N_3139,N_3737);
and U3990 (N_3990,N_3306,N_3020);
and U3991 (N_3991,N_3472,N_3002);
and U3992 (N_3992,N_3058,N_3694);
nor U3993 (N_3993,N_3264,N_3458);
nand U3994 (N_3994,N_3444,N_3023);
and U3995 (N_3995,N_3519,N_3494);
nand U3996 (N_3996,N_3538,N_3319);
nand U3997 (N_3997,N_3592,N_3049);
and U3998 (N_3998,N_3083,N_3254);
nor U3999 (N_3999,N_3229,N_3602);
xor U4000 (N_4000,N_3382,N_3377);
or U4001 (N_4001,N_3330,N_3624);
nand U4002 (N_4002,N_3230,N_3543);
nor U4003 (N_4003,N_3276,N_3144);
nand U4004 (N_4004,N_3487,N_3141);
nor U4005 (N_4005,N_3681,N_3679);
nand U4006 (N_4006,N_3585,N_3247);
nor U4007 (N_4007,N_3700,N_3611);
or U4008 (N_4008,N_3367,N_3731);
nor U4009 (N_4009,N_3570,N_3669);
nor U4010 (N_4010,N_3090,N_3663);
nor U4011 (N_4011,N_3511,N_3361);
or U4012 (N_4012,N_3626,N_3342);
and U4013 (N_4013,N_3169,N_3352);
or U4014 (N_4014,N_3478,N_3149);
or U4015 (N_4015,N_3438,N_3048);
nor U4016 (N_4016,N_3115,N_3029);
xnor U4017 (N_4017,N_3113,N_3165);
or U4018 (N_4018,N_3146,N_3660);
nor U4019 (N_4019,N_3606,N_3109);
or U4020 (N_4020,N_3604,N_3344);
and U4021 (N_4021,N_3031,N_3172);
nor U4022 (N_4022,N_3045,N_3513);
or U4023 (N_4023,N_3042,N_3291);
and U4024 (N_4024,N_3179,N_3032);
or U4025 (N_4025,N_3219,N_3176);
and U4026 (N_4026,N_3120,N_3443);
nor U4027 (N_4027,N_3055,N_3282);
nand U4028 (N_4028,N_3304,N_3475);
xor U4029 (N_4029,N_3102,N_3599);
nor U4030 (N_4030,N_3526,N_3457);
and U4031 (N_4031,N_3295,N_3442);
and U4032 (N_4032,N_3554,N_3242);
nor U4033 (N_4033,N_3531,N_3196);
and U4034 (N_4034,N_3614,N_3577);
xor U4035 (N_4035,N_3143,N_3618);
and U4036 (N_4036,N_3227,N_3560);
xor U4037 (N_4037,N_3094,N_3537);
and U4038 (N_4038,N_3299,N_3024);
and U4039 (N_4039,N_3373,N_3345);
xor U4040 (N_4040,N_3257,N_3004);
and U4041 (N_4041,N_3488,N_3684);
nand U4042 (N_4042,N_3551,N_3587);
nor U4043 (N_4043,N_3184,N_3208);
nor U4044 (N_4044,N_3037,N_3069);
nand U4045 (N_4045,N_3326,N_3417);
or U4046 (N_4046,N_3337,N_3591);
nand U4047 (N_4047,N_3702,N_3616);
and U4048 (N_4048,N_3709,N_3508);
or U4049 (N_4049,N_3396,N_3461);
or U4050 (N_4050,N_3609,N_3545);
or U4051 (N_4051,N_3000,N_3145);
nor U4052 (N_4052,N_3385,N_3589);
nand U4053 (N_4053,N_3437,N_3313);
nor U4054 (N_4054,N_3532,N_3061);
and U4055 (N_4055,N_3273,N_3269);
and U4056 (N_4056,N_3371,N_3484);
nor U4057 (N_4057,N_3586,N_3003);
nand U4058 (N_4058,N_3474,N_3688);
nor U4059 (N_4059,N_3349,N_3534);
nand U4060 (N_4060,N_3131,N_3200);
nor U4061 (N_4061,N_3598,N_3667);
or U4062 (N_4062,N_3724,N_3357);
and U4063 (N_4063,N_3711,N_3398);
and U4064 (N_4064,N_3605,N_3510);
and U4065 (N_4065,N_3065,N_3082);
nor U4066 (N_4066,N_3627,N_3368);
nor U4067 (N_4067,N_3736,N_3379);
and U4068 (N_4068,N_3052,N_3070);
or U4069 (N_4069,N_3620,N_3733);
and U4070 (N_4070,N_3270,N_3486);
xnor U4071 (N_4071,N_3118,N_3112);
xnor U4072 (N_4072,N_3402,N_3492);
or U4073 (N_4073,N_3151,N_3597);
and U4074 (N_4074,N_3697,N_3341);
nand U4075 (N_4075,N_3211,N_3467);
or U4076 (N_4076,N_3509,N_3171);
nor U4077 (N_4077,N_3541,N_3288);
and U4078 (N_4078,N_3347,N_3683);
nor U4079 (N_4079,N_3332,N_3041);
nor U4080 (N_4080,N_3425,N_3713);
nor U4081 (N_4081,N_3321,N_3293);
xor U4082 (N_4082,N_3170,N_3730);
nand U4083 (N_4083,N_3677,N_3286);
xor U4084 (N_4084,N_3267,N_3740);
nor U4085 (N_4085,N_3259,N_3054);
or U4086 (N_4086,N_3703,N_3280);
and U4087 (N_4087,N_3239,N_3079);
xor U4088 (N_4088,N_3601,N_3658);
nand U4089 (N_4089,N_3075,N_3625);
and U4090 (N_4090,N_3386,N_3454);
xnor U4091 (N_4091,N_3583,N_3394);
or U4092 (N_4092,N_3019,N_3578);
or U4093 (N_4093,N_3391,N_3552);
or U4094 (N_4094,N_3748,N_3640);
or U4095 (N_4095,N_3387,N_3353);
and U4096 (N_4096,N_3238,N_3209);
and U4097 (N_4097,N_3081,N_3051);
and U4098 (N_4098,N_3514,N_3148);
nand U4099 (N_4099,N_3646,N_3289);
or U4100 (N_4100,N_3086,N_3028);
nand U4101 (N_4101,N_3168,N_3399);
xor U4102 (N_4102,N_3067,N_3462);
nor U4103 (N_4103,N_3157,N_3121);
nor U4104 (N_4104,N_3415,N_3327);
nand U4105 (N_4105,N_3434,N_3188);
nor U4106 (N_4106,N_3036,N_3406);
or U4107 (N_4107,N_3576,N_3479);
and U4108 (N_4108,N_3404,N_3063);
or U4109 (N_4109,N_3068,N_3333);
and U4110 (N_4110,N_3046,N_3495);
nor U4111 (N_4111,N_3246,N_3017);
xor U4112 (N_4112,N_3057,N_3035);
and U4113 (N_4113,N_3316,N_3473);
and U4114 (N_4114,N_3595,N_3600);
nor U4115 (N_4115,N_3030,N_3584);
nor U4116 (N_4116,N_3071,N_3226);
nand U4117 (N_4117,N_3018,N_3408);
nor U4118 (N_4118,N_3482,N_3407);
nand U4119 (N_4119,N_3027,N_3633);
nor U4120 (N_4120,N_3596,N_3215);
and U4121 (N_4121,N_3496,N_3708);
xor U4122 (N_4122,N_3356,N_3365);
and U4123 (N_4123,N_3520,N_3301);
nand U4124 (N_4124,N_3739,N_3433);
and U4125 (N_4125,N_3552,N_3212);
and U4126 (N_4126,N_3006,N_3707);
and U4127 (N_4127,N_3245,N_3065);
and U4128 (N_4128,N_3558,N_3507);
and U4129 (N_4129,N_3434,N_3174);
xor U4130 (N_4130,N_3610,N_3111);
nand U4131 (N_4131,N_3402,N_3126);
or U4132 (N_4132,N_3114,N_3586);
nor U4133 (N_4133,N_3725,N_3026);
xor U4134 (N_4134,N_3117,N_3003);
and U4135 (N_4135,N_3245,N_3331);
and U4136 (N_4136,N_3280,N_3568);
xnor U4137 (N_4137,N_3395,N_3167);
or U4138 (N_4138,N_3382,N_3115);
or U4139 (N_4139,N_3703,N_3631);
and U4140 (N_4140,N_3514,N_3074);
nor U4141 (N_4141,N_3471,N_3242);
nand U4142 (N_4142,N_3686,N_3033);
and U4143 (N_4143,N_3355,N_3198);
and U4144 (N_4144,N_3211,N_3272);
or U4145 (N_4145,N_3143,N_3412);
nor U4146 (N_4146,N_3705,N_3230);
xnor U4147 (N_4147,N_3417,N_3227);
or U4148 (N_4148,N_3100,N_3716);
and U4149 (N_4149,N_3108,N_3288);
nand U4150 (N_4150,N_3219,N_3564);
or U4151 (N_4151,N_3433,N_3488);
xnor U4152 (N_4152,N_3740,N_3127);
nand U4153 (N_4153,N_3406,N_3701);
or U4154 (N_4154,N_3321,N_3597);
xnor U4155 (N_4155,N_3402,N_3247);
nand U4156 (N_4156,N_3249,N_3042);
xnor U4157 (N_4157,N_3225,N_3153);
xor U4158 (N_4158,N_3361,N_3142);
nand U4159 (N_4159,N_3732,N_3069);
nor U4160 (N_4160,N_3570,N_3077);
nand U4161 (N_4161,N_3444,N_3580);
and U4162 (N_4162,N_3748,N_3595);
nor U4163 (N_4163,N_3157,N_3221);
and U4164 (N_4164,N_3733,N_3470);
or U4165 (N_4165,N_3225,N_3224);
nor U4166 (N_4166,N_3468,N_3152);
and U4167 (N_4167,N_3187,N_3604);
nor U4168 (N_4168,N_3569,N_3284);
nor U4169 (N_4169,N_3309,N_3120);
or U4170 (N_4170,N_3192,N_3207);
or U4171 (N_4171,N_3152,N_3332);
nand U4172 (N_4172,N_3195,N_3109);
and U4173 (N_4173,N_3233,N_3280);
nor U4174 (N_4174,N_3458,N_3523);
or U4175 (N_4175,N_3045,N_3149);
or U4176 (N_4176,N_3493,N_3322);
nand U4177 (N_4177,N_3689,N_3682);
or U4178 (N_4178,N_3092,N_3568);
nand U4179 (N_4179,N_3500,N_3624);
nand U4180 (N_4180,N_3244,N_3281);
nand U4181 (N_4181,N_3010,N_3113);
and U4182 (N_4182,N_3387,N_3516);
or U4183 (N_4183,N_3589,N_3392);
nor U4184 (N_4184,N_3515,N_3724);
or U4185 (N_4185,N_3015,N_3415);
or U4186 (N_4186,N_3380,N_3313);
xor U4187 (N_4187,N_3634,N_3358);
or U4188 (N_4188,N_3043,N_3636);
nor U4189 (N_4189,N_3263,N_3520);
nand U4190 (N_4190,N_3087,N_3153);
nand U4191 (N_4191,N_3688,N_3749);
nor U4192 (N_4192,N_3724,N_3070);
nor U4193 (N_4193,N_3417,N_3448);
or U4194 (N_4194,N_3392,N_3721);
or U4195 (N_4195,N_3148,N_3133);
and U4196 (N_4196,N_3451,N_3076);
and U4197 (N_4197,N_3344,N_3106);
and U4198 (N_4198,N_3021,N_3642);
and U4199 (N_4199,N_3682,N_3472);
or U4200 (N_4200,N_3335,N_3662);
and U4201 (N_4201,N_3138,N_3315);
nor U4202 (N_4202,N_3124,N_3243);
or U4203 (N_4203,N_3626,N_3049);
and U4204 (N_4204,N_3135,N_3287);
and U4205 (N_4205,N_3216,N_3587);
nand U4206 (N_4206,N_3360,N_3440);
nor U4207 (N_4207,N_3101,N_3226);
nand U4208 (N_4208,N_3440,N_3013);
xnor U4209 (N_4209,N_3447,N_3478);
xor U4210 (N_4210,N_3090,N_3299);
nand U4211 (N_4211,N_3265,N_3016);
or U4212 (N_4212,N_3301,N_3387);
nor U4213 (N_4213,N_3484,N_3129);
nor U4214 (N_4214,N_3451,N_3657);
or U4215 (N_4215,N_3396,N_3344);
xnor U4216 (N_4216,N_3441,N_3053);
xnor U4217 (N_4217,N_3365,N_3227);
nor U4218 (N_4218,N_3627,N_3236);
or U4219 (N_4219,N_3500,N_3278);
or U4220 (N_4220,N_3144,N_3373);
and U4221 (N_4221,N_3109,N_3112);
or U4222 (N_4222,N_3547,N_3269);
nand U4223 (N_4223,N_3098,N_3418);
and U4224 (N_4224,N_3539,N_3567);
nand U4225 (N_4225,N_3392,N_3186);
nor U4226 (N_4226,N_3642,N_3472);
and U4227 (N_4227,N_3489,N_3109);
and U4228 (N_4228,N_3657,N_3673);
xnor U4229 (N_4229,N_3385,N_3304);
nand U4230 (N_4230,N_3670,N_3505);
nand U4231 (N_4231,N_3438,N_3228);
xnor U4232 (N_4232,N_3442,N_3252);
nand U4233 (N_4233,N_3581,N_3683);
and U4234 (N_4234,N_3326,N_3497);
or U4235 (N_4235,N_3366,N_3225);
nand U4236 (N_4236,N_3382,N_3391);
xnor U4237 (N_4237,N_3108,N_3009);
nand U4238 (N_4238,N_3392,N_3722);
or U4239 (N_4239,N_3546,N_3116);
or U4240 (N_4240,N_3410,N_3524);
nor U4241 (N_4241,N_3318,N_3549);
nor U4242 (N_4242,N_3476,N_3472);
nand U4243 (N_4243,N_3587,N_3452);
nand U4244 (N_4244,N_3456,N_3193);
nand U4245 (N_4245,N_3446,N_3529);
and U4246 (N_4246,N_3479,N_3599);
xor U4247 (N_4247,N_3467,N_3513);
nor U4248 (N_4248,N_3675,N_3450);
nand U4249 (N_4249,N_3531,N_3366);
nand U4250 (N_4250,N_3384,N_3477);
or U4251 (N_4251,N_3176,N_3675);
or U4252 (N_4252,N_3661,N_3047);
or U4253 (N_4253,N_3405,N_3382);
or U4254 (N_4254,N_3506,N_3323);
and U4255 (N_4255,N_3586,N_3060);
nor U4256 (N_4256,N_3233,N_3598);
nor U4257 (N_4257,N_3678,N_3241);
and U4258 (N_4258,N_3660,N_3639);
and U4259 (N_4259,N_3553,N_3725);
xor U4260 (N_4260,N_3586,N_3448);
or U4261 (N_4261,N_3309,N_3714);
nor U4262 (N_4262,N_3568,N_3060);
nand U4263 (N_4263,N_3648,N_3583);
nor U4264 (N_4264,N_3059,N_3691);
nor U4265 (N_4265,N_3744,N_3503);
and U4266 (N_4266,N_3624,N_3394);
xor U4267 (N_4267,N_3588,N_3494);
and U4268 (N_4268,N_3039,N_3644);
xnor U4269 (N_4269,N_3015,N_3511);
and U4270 (N_4270,N_3310,N_3618);
nor U4271 (N_4271,N_3691,N_3100);
nor U4272 (N_4272,N_3459,N_3311);
or U4273 (N_4273,N_3543,N_3489);
or U4274 (N_4274,N_3152,N_3694);
or U4275 (N_4275,N_3658,N_3161);
or U4276 (N_4276,N_3537,N_3742);
nand U4277 (N_4277,N_3114,N_3211);
nand U4278 (N_4278,N_3604,N_3133);
and U4279 (N_4279,N_3595,N_3638);
nand U4280 (N_4280,N_3373,N_3435);
and U4281 (N_4281,N_3249,N_3431);
or U4282 (N_4282,N_3623,N_3168);
nor U4283 (N_4283,N_3033,N_3478);
or U4284 (N_4284,N_3206,N_3718);
nand U4285 (N_4285,N_3237,N_3346);
or U4286 (N_4286,N_3112,N_3435);
nand U4287 (N_4287,N_3397,N_3725);
and U4288 (N_4288,N_3078,N_3226);
nor U4289 (N_4289,N_3309,N_3743);
nor U4290 (N_4290,N_3184,N_3481);
or U4291 (N_4291,N_3473,N_3143);
or U4292 (N_4292,N_3522,N_3690);
nand U4293 (N_4293,N_3621,N_3115);
nand U4294 (N_4294,N_3521,N_3655);
nor U4295 (N_4295,N_3655,N_3522);
or U4296 (N_4296,N_3261,N_3136);
xnor U4297 (N_4297,N_3486,N_3395);
nand U4298 (N_4298,N_3685,N_3483);
nor U4299 (N_4299,N_3466,N_3034);
nand U4300 (N_4300,N_3722,N_3296);
nor U4301 (N_4301,N_3130,N_3090);
nand U4302 (N_4302,N_3153,N_3589);
nor U4303 (N_4303,N_3591,N_3026);
nand U4304 (N_4304,N_3711,N_3548);
nand U4305 (N_4305,N_3298,N_3668);
nor U4306 (N_4306,N_3558,N_3470);
or U4307 (N_4307,N_3554,N_3727);
nand U4308 (N_4308,N_3596,N_3747);
and U4309 (N_4309,N_3475,N_3044);
nor U4310 (N_4310,N_3187,N_3479);
nor U4311 (N_4311,N_3308,N_3299);
nor U4312 (N_4312,N_3534,N_3434);
and U4313 (N_4313,N_3487,N_3628);
and U4314 (N_4314,N_3019,N_3478);
nor U4315 (N_4315,N_3647,N_3123);
nor U4316 (N_4316,N_3062,N_3462);
nor U4317 (N_4317,N_3135,N_3354);
nor U4318 (N_4318,N_3741,N_3501);
and U4319 (N_4319,N_3280,N_3268);
or U4320 (N_4320,N_3294,N_3078);
nand U4321 (N_4321,N_3137,N_3338);
nor U4322 (N_4322,N_3370,N_3562);
and U4323 (N_4323,N_3201,N_3576);
nand U4324 (N_4324,N_3248,N_3588);
or U4325 (N_4325,N_3461,N_3454);
or U4326 (N_4326,N_3236,N_3707);
nor U4327 (N_4327,N_3280,N_3536);
nand U4328 (N_4328,N_3190,N_3449);
nand U4329 (N_4329,N_3354,N_3129);
nor U4330 (N_4330,N_3366,N_3169);
nor U4331 (N_4331,N_3694,N_3197);
and U4332 (N_4332,N_3158,N_3607);
and U4333 (N_4333,N_3334,N_3072);
or U4334 (N_4334,N_3284,N_3508);
nor U4335 (N_4335,N_3644,N_3109);
and U4336 (N_4336,N_3430,N_3517);
nor U4337 (N_4337,N_3459,N_3491);
nand U4338 (N_4338,N_3318,N_3115);
and U4339 (N_4339,N_3338,N_3672);
and U4340 (N_4340,N_3537,N_3635);
and U4341 (N_4341,N_3110,N_3653);
nand U4342 (N_4342,N_3037,N_3401);
and U4343 (N_4343,N_3549,N_3012);
nor U4344 (N_4344,N_3344,N_3084);
and U4345 (N_4345,N_3053,N_3257);
or U4346 (N_4346,N_3348,N_3213);
and U4347 (N_4347,N_3748,N_3557);
nand U4348 (N_4348,N_3144,N_3006);
or U4349 (N_4349,N_3467,N_3287);
xnor U4350 (N_4350,N_3412,N_3254);
xor U4351 (N_4351,N_3120,N_3029);
nand U4352 (N_4352,N_3550,N_3361);
nor U4353 (N_4353,N_3299,N_3129);
xor U4354 (N_4354,N_3137,N_3309);
nand U4355 (N_4355,N_3568,N_3401);
or U4356 (N_4356,N_3164,N_3557);
nor U4357 (N_4357,N_3313,N_3452);
or U4358 (N_4358,N_3308,N_3413);
nor U4359 (N_4359,N_3552,N_3083);
nand U4360 (N_4360,N_3123,N_3711);
and U4361 (N_4361,N_3572,N_3671);
nor U4362 (N_4362,N_3131,N_3233);
nand U4363 (N_4363,N_3092,N_3313);
nand U4364 (N_4364,N_3619,N_3061);
nor U4365 (N_4365,N_3585,N_3015);
nor U4366 (N_4366,N_3470,N_3307);
and U4367 (N_4367,N_3085,N_3177);
nand U4368 (N_4368,N_3606,N_3517);
nor U4369 (N_4369,N_3198,N_3089);
nand U4370 (N_4370,N_3212,N_3242);
nor U4371 (N_4371,N_3349,N_3728);
nor U4372 (N_4372,N_3419,N_3722);
nand U4373 (N_4373,N_3747,N_3541);
and U4374 (N_4374,N_3148,N_3713);
nand U4375 (N_4375,N_3607,N_3007);
xnor U4376 (N_4376,N_3487,N_3118);
xor U4377 (N_4377,N_3620,N_3168);
nor U4378 (N_4378,N_3273,N_3195);
nand U4379 (N_4379,N_3452,N_3747);
or U4380 (N_4380,N_3680,N_3561);
nand U4381 (N_4381,N_3341,N_3238);
or U4382 (N_4382,N_3176,N_3141);
xor U4383 (N_4383,N_3165,N_3133);
and U4384 (N_4384,N_3706,N_3040);
and U4385 (N_4385,N_3505,N_3384);
nor U4386 (N_4386,N_3690,N_3449);
or U4387 (N_4387,N_3164,N_3163);
or U4388 (N_4388,N_3505,N_3261);
nor U4389 (N_4389,N_3536,N_3006);
xnor U4390 (N_4390,N_3415,N_3025);
or U4391 (N_4391,N_3407,N_3725);
nor U4392 (N_4392,N_3444,N_3161);
nand U4393 (N_4393,N_3597,N_3728);
and U4394 (N_4394,N_3176,N_3052);
nor U4395 (N_4395,N_3211,N_3609);
nand U4396 (N_4396,N_3093,N_3188);
nor U4397 (N_4397,N_3580,N_3052);
nor U4398 (N_4398,N_3308,N_3548);
and U4399 (N_4399,N_3736,N_3041);
or U4400 (N_4400,N_3456,N_3400);
or U4401 (N_4401,N_3330,N_3261);
nor U4402 (N_4402,N_3399,N_3320);
or U4403 (N_4403,N_3666,N_3496);
xnor U4404 (N_4404,N_3330,N_3235);
nor U4405 (N_4405,N_3515,N_3621);
nand U4406 (N_4406,N_3301,N_3434);
and U4407 (N_4407,N_3013,N_3241);
nor U4408 (N_4408,N_3322,N_3617);
or U4409 (N_4409,N_3070,N_3659);
and U4410 (N_4410,N_3115,N_3018);
nand U4411 (N_4411,N_3298,N_3031);
nand U4412 (N_4412,N_3343,N_3737);
xnor U4413 (N_4413,N_3264,N_3583);
or U4414 (N_4414,N_3195,N_3261);
nor U4415 (N_4415,N_3317,N_3585);
nor U4416 (N_4416,N_3382,N_3519);
nand U4417 (N_4417,N_3481,N_3536);
nor U4418 (N_4418,N_3260,N_3492);
or U4419 (N_4419,N_3251,N_3353);
or U4420 (N_4420,N_3505,N_3295);
and U4421 (N_4421,N_3206,N_3717);
and U4422 (N_4422,N_3662,N_3257);
nand U4423 (N_4423,N_3714,N_3330);
and U4424 (N_4424,N_3297,N_3321);
nand U4425 (N_4425,N_3464,N_3719);
nand U4426 (N_4426,N_3608,N_3643);
and U4427 (N_4427,N_3266,N_3246);
nand U4428 (N_4428,N_3416,N_3403);
and U4429 (N_4429,N_3664,N_3398);
nand U4430 (N_4430,N_3694,N_3021);
nor U4431 (N_4431,N_3726,N_3072);
or U4432 (N_4432,N_3527,N_3136);
or U4433 (N_4433,N_3657,N_3723);
nor U4434 (N_4434,N_3720,N_3356);
or U4435 (N_4435,N_3558,N_3612);
nand U4436 (N_4436,N_3459,N_3646);
nor U4437 (N_4437,N_3549,N_3631);
nand U4438 (N_4438,N_3235,N_3318);
nor U4439 (N_4439,N_3628,N_3598);
nand U4440 (N_4440,N_3633,N_3705);
nand U4441 (N_4441,N_3237,N_3697);
xnor U4442 (N_4442,N_3680,N_3402);
nor U4443 (N_4443,N_3261,N_3714);
and U4444 (N_4444,N_3375,N_3153);
nor U4445 (N_4445,N_3240,N_3386);
xor U4446 (N_4446,N_3540,N_3118);
nand U4447 (N_4447,N_3159,N_3650);
nor U4448 (N_4448,N_3112,N_3330);
and U4449 (N_4449,N_3354,N_3187);
and U4450 (N_4450,N_3620,N_3306);
nor U4451 (N_4451,N_3304,N_3697);
and U4452 (N_4452,N_3173,N_3470);
and U4453 (N_4453,N_3317,N_3206);
and U4454 (N_4454,N_3495,N_3563);
or U4455 (N_4455,N_3113,N_3202);
or U4456 (N_4456,N_3538,N_3638);
or U4457 (N_4457,N_3313,N_3373);
nor U4458 (N_4458,N_3454,N_3727);
nor U4459 (N_4459,N_3308,N_3234);
nand U4460 (N_4460,N_3090,N_3715);
or U4461 (N_4461,N_3660,N_3131);
xor U4462 (N_4462,N_3723,N_3640);
or U4463 (N_4463,N_3012,N_3246);
nor U4464 (N_4464,N_3018,N_3261);
or U4465 (N_4465,N_3270,N_3493);
and U4466 (N_4466,N_3080,N_3156);
nand U4467 (N_4467,N_3165,N_3331);
or U4468 (N_4468,N_3322,N_3017);
nor U4469 (N_4469,N_3518,N_3698);
nor U4470 (N_4470,N_3235,N_3224);
nor U4471 (N_4471,N_3563,N_3041);
nand U4472 (N_4472,N_3531,N_3309);
and U4473 (N_4473,N_3680,N_3182);
and U4474 (N_4474,N_3440,N_3347);
nor U4475 (N_4475,N_3562,N_3697);
or U4476 (N_4476,N_3644,N_3271);
nor U4477 (N_4477,N_3589,N_3696);
nand U4478 (N_4478,N_3143,N_3490);
or U4479 (N_4479,N_3585,N_3511);
nor U4480 (N_4480,N_3269,N_3665);
and U4481 (N_4481,N_3284,N_3243);
or U4482 (N_4482,N_3447,N_3278);
nand U4483 (N_4483,N_3102,N_3162);
nor U4484 (N_4484,N_3202,N_3719);
nand U4485 (N_4485,N_3710,N_3123);
or U4486 (N_4486,N_3112,N_3535);
nor U4487 (N_4487,N_3417,N_3128);
nand U4488 (N_4488,N_3566,N_3663);
nand U4489 (N_4489,N_3049,N_3571);
nor U4490 (N_4490,N_3048,N_3259);
and U4491 (N_4491,N_3233,N_3254);
nor U4492 (N_4492,N_3298,N_3307);
and U4493 (N_4493,N_3433,N_3490);
and U4494 (N_4494,N_3666,N_3309);
nor U4495 (N_4495,N_3146,N_3583);
and U4496 (N_4496,N_3240,N_3159);
or U4497 (N_4497,N_3542,N_3545);
nand U4498 (N_4498,N_3267,N_3669);
nand U4499 (N_4499,N_3412,N_3617);
and U4500 (N_4500,N_3804,N_4002);
and U4501 (N_4501,N_4313,N_4260);
xor U4502 (N_4502,N_4106,N_3878);
or U4503 (N_4503,N_3909,N_4471);
xor U4504 (N_4504,N_4129,N_4009);
nor U4505 (N_4505,N_4105,N_4447);
or U4506 (N_4506,N_4253,N_4239);
or U4507 (N_4507,N_4053,N_3820);
or U4508 (N_4508,N_4329,N_4376);
and U4509 (N_4509,N_4144,N_4493);
or U4510 (N_4510,N_4177,N_4265);
nor U4511 (N_4511,N_4269,N_3825);
xor U4512 (N_4512,N_4198,N_4288);
nor U4513 (N_4513,N_4403,N_4016);
and U4514 (N_4514,N_4424,N_4209);
and U4515 (N_4515,N_4461,N_4175);
xnor U4516 (N_4516,N_4130,N_4281);
and U4517 (N_4517,N_4319,N_3939);
and U4518 (N_4518,N_4217,N_4466);
or U4519 (N_4519,N_4390,N_3784);
and U4520 (N_4520,N_4399,N_4299);
or U4521 (N_4521,N_3896,N_3759);
or U4522 (N_4522,N_4490,N_4076);
nand U4523 (N_4523,N_4133,N_4131);
or U4524 (N_4524,N_4092,N_4214);
and U4525 (N_4525,N_4479,N_4311);
nor U4526 (N_4526,N_4320,N_3757);
or U4527 (N_4527,N_3867,N_3954);
and U4528 (N_4528,N_3862,N_4426);
nand U4529 (N_4529,N_4145,N_4019);
and U4530 (N_4530,N_4407,N_4441);
or U4531 (N_4531,N_4472,N_3929);
nand U4532 (N_4532,N_4344,N_4012);
nand U4533 (N_4533,N_4402,N_4374);
xor U4534 (N_4534,N_4478,N_3947);
nor U4535 (N_4535,N_4082,N_4123);
or U4536 (N_4536,N_4307,N_4210);
nor U4537 (N_4537,N_3856,N_3933);
nand U4538 (N_4538,N_4222,N_4100);
nor U4539 (N_4539,N_4388,N_4110);
nor U4540 (N_4540,N_4237,N_3777);
and U4541 (N_4541,N_4263,N_3807);
nand U4542 (N_4542,N_3767,N_4273);
and U4543 (N_4543,N_4365,N_4301);
nor U4544 (N_4544,N_4433,N_3864);
nand U4545 (N_4545,N_4404,N_3985);
and U4546 (N_4546,N_4168,N_4496);
and U4547 (N_4547,N_4090,N_3790);
nor U4548 (N_4548,N_3941,N_4430);
nor U4549 (N_4549,N_4151,N_4292);
or U4550 (N_4550,N_3756,N_3844);
nand U4551 (N_4551,N_3860,N_4346);
xor U4552 (N_4552,N_4325,N_4382);
and U4553 (N_4553,N_4314,N_4289);
nor U4554 (N_4554,N_4455,N_4272);
or U4555 (N_4555,N_4436,N_4440);
and U4556 (N_4556,N_3910,N_3801);
nand U4557 (N_4557,N_3871,N_3949);
nand U4558 (N_4558,N_3880,N_4425);
and U4559 (N_4559,N_4184,N_3932);
xor U4560 (N_4560,N_4228,N_4229);
and U4561 (N_4561,N_4484,N_4073);
xnor U4562 (N_4562,N_4003,N_4491);
or U4563 (N_4563,N_4075,N_4348);
nor U4564 (N_4564,N_3771,N_4234);
nand U4565 (N_4565,N_4206,N_4341);
nor U4566 (N_4566,N_3898,N_3779);
or U4567 (N_4567,N_4393,N_4040);
nor U4568 (N_4568,N_4457,N_4309);
nand U4569 (N_4569,N_4069,N_3964);
or U4570 (N_4570,N_4182,N_3972);
nor U4571 (N_4571,N_4026,N_4387);
nand U4572 (N_4572,N_4308,N_4164);
nand U4573 (N_4573,N_3889,N_3828);
nand U4574 (N_4574,N_4054,N_4072);
or U4575 (N_4575,N_4460,N_3931);
nor U4576 (N_4576,N_4159,N_3793);
nor U4577 (N_4577,N_4371,N_3959);
nor U4578 (N_4578,N_4302,N_3886);
and U4579 (N_4579,N_4088,N_3785);
or U4580 (N_4580,N_4071,N_3915);
and U4581 (N_4581,N_4029,N_4049);
nor U4582 (N_4582,N_4428,N_4323);
nor U4583 (N_4583,N_3965,N_4038);
or U4584 (N_4584,N_3960,N_4337);
nand U4585 (N_4585,N_4041,N_4140);
xor U4586 (N_4586,N_3796,N_4443);
or U4587 (N_4587,N_4326,N_4458);
and U4588 (N_4588,N_4095,N_4279);
and U4589 (N_4589,N_4045,N_4459);
nand U4590 (N_4590,N_4321,N_4004);
nor U4591 (N_4591,N_3925,N_4285);
or U4592 (N_4592,N_3859,N_3951);
nor U4593 (N_4593,N_4429,N_3913);
or U4594 (N_4594,N_4454,N_4275);
nor U4595 (N_4595,N_4423,N_3952);
and U4596 (N_4596,N_4333,N_4070);
and U4597 (N_4597,N_4481,N_4189);
or U4598 (N_4598,N_4103,N_3957);
xnor U4599 (N_4599,N_4287,N_4013);
xnor U4600 (N_4600,N_3837,N_4043);
and U4601 (N_4601,N_4059,N_4022);
or U4602 (N_4602,N_4120,N_4086);
nor U4603 (N_4603,N_4416,N_3927);
or U4604 (N_4604,N_3794,N_4349);
nand U4605 (N_4605,N_3845,N_4111);
and U4606 (N_4606,N_3787,N_3826);
nor U4607 (N_4607,N_4477,N_4473);
xnor U4608 (N_4608,N_4267,N_4405);
and U4609 (N_4609,N_3953,N_4453);
nand U4610 (N_4610,N_4044,N_4166);
and U4611 (N_4611,N_3866,N_4097);
nand U4612 (N_4612,N_3803,N_4354);
or U4613 (N_4613,N_4480,N_3938);
or U4614 (N_4614,N_4243,N_4383);
nand U4615 (N_4615,N_3956,N_3791);
or U4616 (N_4616,N_4055,N_3795);
or U4617 (N_4617,N_4274,N_4412);
nand U4618 (N_4618,N_4282,N_4452);
nand U4619 (N_4619,N_3919,N_3942);
nand U4620 (N_4620,N_3810,N_4137);
or U4621 (N_4621,N_4224,N_4067);
and U4622 (N_4622,N_3935,N_4396);
or U4623 (N_4623,N_4398,N_4363);
nand U4624 (N_4624,N_4257,N_4215);
nor U4625 (N_4625,N_4298,N_4352);
or U4626 (N_4626,N_4085,N_4465);
nand U4627 (N_4627,N_4271,N_4020);
nor U4628 (N_4628,N_3943,N_4468);
xor U4629 (N_4629,N_4397,N_4025);
or U4630 (N_4630,N_3870,N_4294);
nand U4631 (N_4631,N_3979,N_4023);
nand U4632 (N_4632,N_4381,N_4204);
nand U4633 (N_4633,N_3893,N_3876);
and U4634 (N_4634,N_4252,N_4027);
nand U4635 (N_4635,N_3991,N_4408);
nor U4636 (N_4636,N_3843,N_3799);
nor U4637 (N_4637,N_4445,N_4030);
and U4638 (N_4638,N_4278,N_3945);
xor U4639 (N_4639,N_4158,N_4330);
nor U4640 (N_4640,N_4091,N_4450);
nand U4641 (N_4641,N_3976,N_3924);
nand U4642 (N_4642,N_4167,N_4208);
and U4643 (N_4643,N_4211,N_4232);
nor U4644 (N_4644,N_4169,N_3821);
and U4645 (N_4645,N_4052,N_3966);
and U4646 (N_4646,N_4042,N_3881);
nor U4647 (N_4647,N_4369,N_4411);
and U4648 (N_4648,N_4197,N_3923);
nand U4649 (N_4649,N_4074,N_3763);
nor U4650 (N_4650,N_3872,N_3888);
xor U4651 (N_4651,N_3962,N_3934);
and U4652 (N_4652,N_3853,N_4225);
nand U4653 (N_4653,N_3865,N_3936);
nor U4654 (N_4654,N_3887,N_3994);
nor U4655 (N_4655,N_4149,N_4389);
nor U4656 (N_4656,N_4121,N_3921);
nor U4657 (N_4657,N_3980,N_3854);
nor U4658 (N_4658,N_3908,N_4469);
nor U4659 (N_4659,N_4375,N_3814);
and U4660 (N_4660,N_4047,N_3788);
nor U4661 (N_4661,N_4332,N_4057);
and U4662 (N_4662,N_3998,N_3797);
or U4663 (N_4663,N_3831,N_4227);
nand U4664 (N_4664,N_3869,N_4077);
or U4665 (N_4665,N_4394,N_3835);
xnor U4666 (N_4666,N_4286,N_3948);
and U4667 (N_4667,N_4226,N_4083);
nand U4668 (N_4668,N_4179,N_3805);
nor U4669 (N_4669,N_3868,N_4098);
or U4670 (N_4670,N_4081,N_4487);
and U4671 (N_4671,N_4163,N_3916);
or U4672 (N_4672,N_3895,N_4192);
or U4673 (N_4673,N_4034,N_4212);
or U4674 (N_4674,N_4128,N_3839);
xnor U4675 (N_4675,N_4270,N_4018);
nor U4676 (N_4676,N_4356,N_3775);
nand U4677 (N_4677,N_4141,N_4148);
and U4678 (N_4678,N_4361,N_4305);
nand U4679 (N_4679,N_4154,N_4122);
and U4680 (N_4680,N_3899,N_4249);
or U4681 (N_4681,N_4183,N_3848);
and U4682 (N_4682,N_4358,N_3751);
nand U4683 (N_4683,N_4261,N_4233);
or U4684 (N_4684,N_4201,N_4342);
or U4685 (N_4685,N_4199,N_3978);
nor U4686 (N_4686,N_4417,N_4293);
nand U4687 (N_4687,N_3783,N_4024);
nor U4688 (N_4688,N_4339,N_4039);
nand U4689 (N_4689,N_4380,N_4431);
nor U4690 (N_4690,N_4033,N_4345);
nor U4691 (N_4691,N_3911,N_4051);
nand U4692 (N_4692,N_4135,N_3838);
and U4693 (N_4693,N_3920,N_3928);
and U4694 (N_4694,N_3901,N_3892);
or U4695 (N_4695,N_3769,N_3829);
or U4696 (N_4696,N_4336,N_4317);
nand U4697 (N_4697,N_3782,N_4068);
xor U4698 (N_4698,N_4035,N_3841);
or U4699 (N_4699,N_4415,N_4438);
and U4700 (N_4700,N_3973,N_4011);
or U4701 (N_4701,N_4048,N_4343);
or U4702 (N_4702,N_4015,N_4079);
xor U4703 (N_4703,N_3969,N_3846);
or U4704 (N_4704,N_4221,N_3873);
nand U4705 (N_4705,N_3884,N_3778);
or U4706 (N_4706,N_4102,N_4276);
and U4707 (N_4707,N_4219,N_3832);
or U4708 (N_4708,N_4195,N_4124);
nor U4709 (N_4709,N_4060,N_3917);
xnor U4710 (N_4710,N_4118,N_4176);
nand U4711 (N_4711,N_4231,N_4291);
nand U4712 (N_4712,N_3760,N_3834);
or U4713 (N_4713,N_4372,N_4127);
or U4714 (N_4714,N_4134,N_4462);
nand U4715 (N_4715,N_4094,N_4191);
nor U4716 (N_4716,N_3905,N_4259);
and U4717 (N_4717,N_4442,N_3827);
or U4718 (N_4718,N_4364,N_4266);
or U4719 (N_4719,N_4255,N_4165);
or U4720 (N_4720,N_4017,N_4157);
xor U4721 (N_4721,N_4241,N_4084);
nand U4722 (N_4722,N_3819,N_4050);
and U4723 (N_4723,N_4482,N_4008);
nand U4724 (N_4724,N_4406,N_3768);
nor U4725 (N_4725,N_3977,N_4304);
and U4726 (N_4726,N_4032,N_4413);
nand U4727 (N_4727,N_3907,N_4193);
or U4728 (N_4728,N_3988,N_4153);
and U4729 (N_4729,N_4251,N_4155);
nand U4730 (N_4730,N_4010,N_4235);
or U4731 (N_4731,N_3753,N_4006);
nor U4732 (N_4732,N_3818,N_3971);
and U4733 (N_4733,N_3786,N_4001);
nand U4734 (N_4734,N_4400,N_4316);
xnor U4735 (N_4735,N_4242,N_4125);
and U4736 (N_4736,N_4283,N_3990);
and U4737 (N_4737,N_3912,N_3855);
and U4738 (N_4738,N_3993,N_4262);
or U4739 (N_4739,N_4119,N_4180);
and U4740 (N_4740,N_4056,N_4448);
nor U4741 (N_4741,N_3813,N_3926);
nand U4742 (N_4742,N_3766,N_4420);
xor U4743 (N_4743,N_4096,N_4114);
nand U4744 (N_4744,N_3847,N_3885);
nand U4745 (N_4745,N_3809,N_4171);
xor U4746 (N_4746,N_4456,N_4434);
nor U4747 (N_4747,N_3765,N_4203);
nor U4748 (N_4748,N_4474,N_4449);
and U4749 (N_4749,N_4421,N_4498);
or U4750 (N_4750,N_4202,N_4280);
and U4751 (N_4751,N_4046,N_3906);
nand U4752 (N_4752,N_4300,N_3902);
nand U4753 (N_4753,N_4392,N_4318);
and U4754 (N_4754,N_3824,N_3858);
and U4755 (N_4755,N_3750,N_4061);
nand U4756 (N_4756,N_4386,N_4031);
nor U4757 (N_4757,N_4037,N_3922);
nand U4758 (N_4758,N_3780,N_4277);
nor U4759 (N_4759,N_4230,N_4021);
and U4760 (N_4760,N_4470,N_3874);
xnor U4761 (N_4761,N_4451,N_4112);
or U4762 (N_4762,N_3811,N_4435);
and U4763 (N_4763,N_4492,N_3900);
xor U4764 (N_4764,N_3995,N_4126);
nor U4765 (N_4765,N_4007,N_3975);
and U4766 (N_4766,N_3989,N_4328);
nand U4767 (N_4767,N_4312,N_4246);
nand U4768 (N_4768,N_4196,N_4437);
or U4769 (N_4769,N_4258,N_4303);
or U4770 (N_4770,N_4254,N_4036);
or U4771 (N_4771,N_4338,N_3981);
and U4772 (N_4772,N_4160,N_4238);
nand U4773 (N_4773,N_4401,N_4064);
nor U4774 (N_4774,N_3772,N_4475);
nand U4775 (N_4775,N_4156,N_4066);
or U4776 (N_4776,N_4327,N_4395);
nand U4777 (N_4777,N_4324,N_4104);
nand U4778 (N_4778,N_4467,N_4216);
nor U4779 (N_4779,N_4489,N_4014);
nand U4780 (N_4780,N_4350,N_3984);
or U4781 (N_4781,N_3850,N_4264);
nor U4782 (N_4782,N_4200,N_4362);
nor U4783 (N_4783,N_4366,N_3970);
and U4784 (N_4784,N_4315,N_3776);
xnor U4785 (N_4785,N_4116,N_4297);
and U4786 (N_4786,N_4000,N_4143);
or U4787 (N_4787,N_4186,N_3918);
or U4788 (N_4788,N_3894,N_4373);
or U4789 (N_4789,N_3974,N_4244);
and U4790 (N_4790,N_4476,N_4427);
nor U4791 (N_4791,N_3955,N_4139);
or U4792 (N_4792,N_4488,N_4207);
and U4793 (N_4793,N_3997,N_4065);
and U4794 (N_4794,N_3840,N_4357);
nor U4795 (N_4795,N_4223,N_4414);
or U4796 (N_4796,N_4109,N_4432);
nor U4797 (N_4797,N_3816,N_4113);
nand U4798 (N_4798,N_4247,N_3822);
nor U4799 (N_4799,N_3792,N_3857);
nand U4800 (N_4800,N_3897,N_3982);
or U4801 (N_4801,N_4322,N_4385);
or U4802 (N_4802,N_3754,N_3781);
or U4803 (N_4803,N_4117,N_4146);
or U4804 (N_4804,N_4446,N_4409);
nor U4805 (N_4805,N_3914,N_4236);
nor U4806 (N_4806,N_4485,N_4334);
or U4807 (N_4807,N_3999,N_3861);
nand U4808 (N_4808,N_4439,N_4379);
xor U4809 (N_4809,N_3836,N_3830);
nor U4810 (N_4810,N_4367,N_4173);
nor U4811 (N_4811,N_4162,N_3996);
nand U4812 (N_4812,N_4087,N_4378);
nand U4813 (N_4813,N_4355,N_4170);
xnor U4814 (N_4814,N_4172,N_4078);
nor U4815 (N_4815,N_3817,N_4147);
xnor U4816 (N_4816,N_4132,N_3833);
nand U4817 (N_4817,N_4360,N_3968);
nand U4818 (N_4818,N_3852,N_3851);
and U4819 (N_4819,N_4384,N_3770);
nor U4820 (N_4820,N_4290,N_3903);
nand U4821 (N_4821,N_4089,N_4296);
xnor U4822 (N_4822,N_3764,N_3842);
nor U4823 (N_4823,N_3937,N_3815);
or U4824 (N_4824,N_4005,N_4250);
or U4825 (N_4825,N_3761,N_4483);
and U4826 (N_4826,N_3875,N_3946);
and U4827 (N_4827,N_3762,N_3891);
nand U4828 (N_4828,N_4181,N_4188);
and U4829 (N_4829,N_4099,N_4444);
and U4830 (N_4830,N_3877,N_3890);
nand U4831 (N_4831,N_4495,N_4138);
xnor U4832 (N_4832,N_4218,N_3808);
and U4833 (N_4833,N_3802,N_4331);
xor U4834 (N_4834,N_3983,N_3812);
and U4835 (N_4835,N_4063,N_4245);
or U4836 (N_4836,N_4284,N_4028);
nand U4837 (N_4837,N_4377,N_4093);
and U4838 (N_4838,N_4115,N_3961);
or U4839 (N_4839,N_4306,N_4391);
and U4840 (N_4840,N_4499,N_4136);
or U4841 (N_4841,N_4194,N_4152);
and U4842 (N_4842,N_3879,N_3774);
and U4843 (N_4843,N_4256,N_3806);
nand U4844 (N_4844,N_3944,N_3986);
xnor U4845 (N_4845,N_3883,N_4161);
nor U4846 (N_4846,N_4268,N_4185);
and U4847 (N_4847,N_4108,N_3849);
nor U4848 (N_4848,N_4335,N_4150);
or U4849 (N_4849,N_4295,N_3789);
and U4850 (N_4850,N_4359,N_4463);
nand U4851 (N_4851,N_3798,N_4213);
or U4852 (N_4852,N_4370,N_4101);
or U4853 (N_4853,N_3950,N_4240);
nor U4854 (N_4854,N_4107,N_3823);
nor U4855 (N_4855,N_4353,N_3967);
and U4856 (N_4856,N_4340,N_3987);
or U4857 (N_4857,N_4464,N_4205);
xor U4858 (N_4858,N_4190,N_4410);
nor U4859 (N_4859,N_4486,N_3958);
or U4860 (N_4860,N_3940,N_3882);
or U4861 (N_4861,N_4178,N_4418);
xor U4862 (N_4862,N_3963,N_4187);
xor U4863 (N_4863,N_3930,N_3773);
and U4864 (N_4864,N_4220,N_3755);
or U4865 (N_4865,N_4142,N_3992);
nor U4866 (N_4866,N_3800,N_4058);
nor U4867 (N_4867,N_4310,N_4347);
nor U4868 (N_4868,N_4497,N_4062);
or U4869 (N_4869,N_4368,N_4174);
nand U4870 (N_4870,N_4422,N_4351);
nand U4871 (N_4871,N_4248,N_4080);
or U4872 (N_4872,N_3752,N_3863);
or U4873 (N_4873,N_4419,N_4494);
xor U4874 (N_4874,N_3758,N_3904);
nand U4875 (N_4875,N_3883,N_3886);
nor U4876 (N_4876,N_3804,N_4104);
nand U4877 (N_4877,N_4311,N_4358);
nor U4878 (N_4878,N_3958,N_4160);
or U4879 (N_4879,N_4054,N_4208);
nor U4880 (N_4880,N_3838,N_3803);
nor U4881 (N_4881,N_3933,N_3864);
nor U4882 (N_4882,N_4381,N_4017);
nand U4883 (N_4883,N_4464,N_4321);
nor U4884 (N_4884,N_4208,N_3820);
and U4885 (N_4885,N_3822,N_4334);
nor U4886 (N_4886,N_4312,N_3850);
nor U4887 (N_4887,N_4464,N_4480);
and U4888 (N_4888,N_4213,N_4395);
nand U4889 (N_4889,N_3929,N_4259);
and U4890 (N_4890,N_4325,N_4102);
or U4891 (N_4891,N_3987,N_3792);
or U4892 (N_4892,N_4136,N_3904);
xnor U4893 (N_4893,N_4363,N_4302);
or U4894 (N_4894,N_3780,N_3982);
nand U4895 (N_4895,N_3868,N_3920);
nand U4896 (N_4896,N_4437,N_3894);
xnor U4897 (N_4897,N_4064,N_4105);
or U4898 (N_4898,N_4079,N_4181);
or U4899 (N_4899,N_4214,N_4405);
or U4900 (N_4900,N_3773,N_4230);
nand U4901 (N_4901,N_4202,N_4190);
nand U4902 (N_4902,N_4415,N_4167);
or U4903 (N_4903,N_4357,N_4179);
and U4904 (N_4904,N_3913,N_3895);
and U4905 (N_4905,N_4003,N_3782);
and U4906 (N_4906,N_3937,N_3949);
nand U4907 (N_4907,N_4001,N_4261);
nand U4908 (N_4908,N_4182,N_3862);
xnor U4909 (N_4909,N_4244,N_3802);
nor U4910 (N_4910,N_4134,N_3890);
or U4911 (N_4911,N_3892,N_3884);
or U4912 (N_4912,N_3844,N_4089);
nand U4913 (N_4913,N_4292,N_4018);
or U4914 (N_4914,N_3818,N_4079);
nor U4915 (N_4915,N_4239,N_4001);
xnor U4916 (N_4916,N_3833,N_4160);
nor U4917 (N_4917,N_4161,N_3798);
nand U4918 (N_4918,N_4404,N_4014);
nor U4919 (N_4919,N_4377,N_4095);
and U4920 (N_4920,N_3787,N_3838);
nor U4921 (N_4921,N_4412,N_4372);
and U4922 (N_4922,N_3880,N_4201);
nand U4923 (N_4923,N_3805,N_3835);
or U4924 (N_4924,N_4215,N_4250);
nand U4925 (N_4925,N_4352,N_4441);
and U4926 (N_4926,N_4486,N_3830);
nor U4927 (N_4927,N_4373,N_4403);
or U4928 (N_4928,N_4444,N_4350);
nand U4929 (N_4929,N_4084,N_3840);
xnor U4930 (N_4930,N_4309,N_4013);
nor U4931 (N_4931,N_4120,N_4011);
or U4932 (N_4932,N_4195,N_4353);
nor U4933 (N_4933,N_3823,N_3844);
nor U4934 (N_4934,N_4480,N_3977);
and U4935 (N_4935,N_4337,N_3854);
or U4936 (N_4936,N_4402,N_4177);
and U4937 (N_4937,N_4271,N_4077);
nand U4938 (N_4938,N_4160,N_4344);
nor U4939 (N_4939,N_4097,N_3806);
and U4940 (N_4940,N_4381,N_4479);
nor U4941 (N_4941,N_4189,N_4103);
nand U4942 (N_4942,N_4223,N_4450);
or U4943 (N_4943,N_4039,N_4145);
and U4944 (N_4944,N_4330,N_4439);
and U4945 (N_4945,N_3933,N_4090);
nand U4946 (N_4946,N_4125,N_4254);
nor U4947 (N_4947,N_3779,N_3962);
and U4948 (N_4948,N_4000,N_3956);
nand U4949 (N_4949,N_3835,N_4188);
nand U4950 (N_4950,N_4390,N_3944);
or U4951 (N_4951,N_3754,N_4041);
nor U4952 (N_4952,N_3991,N_4011);
nor U4953 (N_4953,N_4040,N_3758);
or U4954 (N_4954,N_3860,N_3940);
or U4955 (N_4955,N_4291,N_3859);
nor U4956 (N_4956,N_4468,N_4018);
or U4957 (N_4957,N_4104,N_3981);
and U4958 (N_4958,N_3883,N_3777);
and U4959 (N_4959,N_3949,N_4399);
nor U4960 (N_4960,N_4124,N_4484);
or U4961 (N_4961,N_4028,N_3785);
and U4962 (N_4962,N_4038,N_3792);
or U4963 (N_4963,N_3852,N_3977);
or U4964 (N_4964,N_4197,N_4305);
and U4965 (N_4965,N_3825,N_4254);
or U4966 (N_4966,N_4491,N_4191);
and U4967 (N_4967,N_3955,N_3961);
nor U4968 (N_4968,N_4030,N_3936);
xnor U4969 (N_4969,N_4356,N_4363);
or U4970 (N_4970,N_4014,N_4458);
and U4971 (N_4971,N_4144,N_4303);
and U4972 (N_4972,N_4063,N_4373);
xnor U4973 (N_4973,N_4445,N_4494);
nor U4974 (N_4974,N_4128,N_4444);
or U4975 (N_4975,N_4059,N_3768);
nand U4976 (N_4976,N_4094,N_3808);
and U4977 (N_4977,N_4159,N_3868);
nand U4978 (N_4978,N_4111,N_4451);
and U4979 (N_4979,N_3998,N_4374);
and U4980 (N_4980,N_4315,N_4244);
xnor U4981 (N_4981,N_4418,N_3985);
nor U4982 (N_4982,N_3853,N_4365);
and U4983 (N_4983,N_4022,N_4344);
nand U4984 (N_4984,N_4018,N_4386);
and U4985 (N_4985,N_3847,N_3951);
or U4986 (N_4986,N_3762,N_4222);
nor U4987 (N_4987,N_4125,N_3963);
nor U4988 (N_4988,N_4021,N_4054);
nor U4989 (N_4989,N_3763,N_3825);
xor U4990 (N_4990,N_4319,N_3983);
and U4991 (N_4991,N_4283,N_4484);
and U4992 (N_4992,N_4019,N_4111);
and U4993 (N_4993,N_4140,N_4294);
nor U4994 (N_4994,N_4239,N_3787);
or U4995 (N_4995,N_3840,N_4430);
and U4996 (N_4996,N_4354,N_4224);
and U4997 (N_4997,N_3774,N_4499);
nor U4998 (N_4998,N_4031,N_4268);
nor U4999 (N_4999,N_3816,N_4444);
or U5000 (N_5000,N_3754,N_4428);
and U5001 (N_5001,N_4330,N_4375);
nor U5002 (N_5002,N_4237,N_3822);
or U5003 (N_5003,N_4000,N_4338);
and U5004 (N_5004,N_3848,N_4239);
and U5005 (N_5005,N_4240,N_4191);
nand U5006 (N_5006,N_3973,N_4416);
nor U5007 (N_5007,N_3990,N_3816);
nor U5008 (N_5008,N_4271,N_3760);
nor U5009 (N_5009,N_3750,N_3831);
and U5010 (N_5010,N_3823,N_4249);
nand U5011 (N_5011,N_3836,N_4269);
nand U5012 (N_5012,N_4446,N_3895);
and U5013 (N_5013,N_3983,N_4171);
nor U5014 (N_5014,N_3927,N_4430);
and U5015 (N_5015,N_4379,N_4311);
or U5016 (N_5016,N_4412,N_4341);
nand U5017 (N_5017,N_3900,N_4308);
and U5018 (N_5018,N_3964,N_3985);
or U5019 (N_5019,N_4135,N_4003);
xor U5020 (N_5020,N_3893,N_4198);
and U5021 (N_5021,N_3899,N_4214);
nor U5022 (N_5022,N_3879,N_4016);
nand U5023 (N_5023,N_3917,N_4323);
nand U5024 (N_5024,N_4032,N_4169);
nor U5025 (N_5025,N_4410,N_3973);
and U5026 (N_5026,N_4353,N_4356);
xnor U5027 (N_5027,N_4446,N_4190);
nand U5028 (N_5028,N_4439,N_4406);
and U5029 (N_5029,N_3961,N_4011);
or U5030 (N_5030,N_4444,N_3956);
and U5031 (N_5031,N_3901,N_4199);
nand U5032 (N_5032,N_4056,N_4171);
nor U5033 (N_5033,N_4075,N_4380);
nor U5034 (N_5034,N_3996,N_4011);
nand U5035 (N_5035,N_3812,N_4146);
nor U5036 (N_5036,N_4344,N_3996);
xnor U5037 (N_5037,N_3784,N_3904);
nand U5038 (N_5038,N_4341,N_4222);
nor U5039 (N_5039,N_4007,N_3980);
nand U5040 (N_5040,N_3911,N_4300);
and U5041 (N_5041,N_4230,N_4325);
nor U5042 (N_5042,N_4080,N_4152);
and U5043 (N_5043,N_3914,N_3807);
or U5044 (N_5044,N_4103,N_4034);
or U5045 (N_5045,N_4470,N_4347);
nor U5046 (N_5046,N_3926,N_4080);
nand U5047 (N_5047,N_3914,N_4322);
nand U5048 (N_5048,N_4012,N_4313);
nand U5049 (N_5049,N_3885,N_4287);
nand U5050 (N_5050,N_4349,N_4355);
xor U5051 (N_5051,N_4387,N_4331);
and U5052 (N_5052,N_4297,N_4407);
and U5053 (N_5053,N_4040,N_4355);
and U5054 (N_5054,N_3992,N_3887);
nand U5055 (N_5055,N_4262,N_4122);
nand U5056 (N_5056,N_4240,N_4362);
or U5057 (N_5057,N_4170,N_4112);
nor U5058 (N_5058,N_3904,N_3792);
nor U5059 (N_5059,N_3874,N_4330);
nand U5060 (N_5060,N_3817,N_4294);
or U5061 (N_5061,N_4380,N_3769);
xnor U5062 (N_5062,N_4183,N_4420);
and U5063 (N_5063,N_3769,N_4135);
nor U5064 (N_5064,N_4252,N_4024);
or U5065 (N_5065,N_3868,N_4253);
or U5066 (N_5066,N_3851,N_4206);
nor U5067 (N_5067,N_4012,N_4117);
nor U5068 (N_5068,N_4019,N_4366);
nand U5069 (N_5069,N_3914,N_4073);
nor U5070 (N_5070,N_4157,N_3788);
nor U5071 (N_5071,N_4139,N_4251);
and U5072 (N_5072,N_4403,N_3760);
or U5073 (N_5073,N_4042,N_4192);
or U5074 (N_5074,N_4312,N_3946);
xor U5075 (N_5075,N_4105,N_3837);
and U5076 (N_5076,N_4057,N_4403);
or U5077 (N_5077,N_3962,N_4468);
nor U5078 (N_5078,N_4059,N_3783);
nand U5079 (N_5079,N_4223,N_4156);
and U5080 (N_5080,N_4183,N_4099);
nor U5081 (N_5081,N_4421,N_4316);
and U5082 (N_5082,N_4400,N_4009);
xor U5083 (N_5083,N_4099,N_4289);
nor U5084 (N_5084,N_3828,N_3988);
and U5085 (N_5085,N_3836,N_3901);
xnor U5086 (N_5086,N_3998,N_3780);
or U5087 (N_5087,N_4411,N_3885);
or U5088 (N_5088,N_4396,N_4414);
and U5089 (N_5089,N_4226,N_4455);
or U5090 (N_5090,N_3934,N_4260);
and U5091 (N_5091,N_4063,N_4368);
nor U5092 (N_5092,N_4353,N_4240);
nand U5093 (N_5093,N_4171,N_3853);
or U5094 (N_5094,N_4189,N_4489);
nor U5095 (N_5095,N_4071,N_3957);
and U5096 (N_5096,N_3904,N_4133);
or U5097 (N_5097,N_3892,N_4399);
or U5098 (N_5098,N_4018,N_3851);
nor U5099 (N_5099,N_3951,N_4074);
nor U5100 (N_5100,N_4344,N_4266);
nand U5101 (N_5101,N_4011,N_4119);
nor U5102 (N_5102,N_4109,N_4439);
nand U5103 (N_5103,N_3999,N_3960);
or U5104 (N_5104,N_3920,N_4110);
or U5105 (N_5105,N_3944,N_3937);
nand U5106 (N_5106,N_4126,N_4266);
and U5107 (N_5107,N_4232,N_3762);
nand U5108 (N_5108,N_4409,N_4084);
nor U5109 (N_5109,N_3783,N_3949);
nor U5110 (N_5110,N_4078,N_4315);
and U5111 (N_5111,N_4199,N_4078);
or U5112 (N_5112,N_4490,N_4361);
xor U5113 (N_5113,N_4487,N_4086);
and U5114 (N_5114,N_4487,N_4251);
nor U5115 (N_5115,N_3786,N_4262);
nand U5116 (N_5116,N_3815,N_4482);
nand U5117 (N_5117,N_3771,N_3780);
and U5118 (N_5118,N_4002,N_4162);
nor U5119 (N_5119,N_3900,N_4263);
nor U5120 (N_5120,N_4479,N_4031);
nor U5121 (N_5121,N_3962,N_4082);
nor U5122 (N_5122,N_4131,N_4389);
nand U5123 (N_5123,N_4302,N_4407);
and U5124 (N_5124,N_3834,N_4231);
and U5125 (N_5125,N_4298,N_4494);
nand U5126 (N_5126,N_4144,N_4358);
and U5127 (N_5127,N_4233,N_4065);
nor U5128 (N_5128,N_3993,N_4344);
and U5129 (N_5129,N_4191,N_3867);
nand U5130 (N_5130,N_3782,N_4495);
and U5131 (N_5131,N_3919,N_3822);
and U5132 (N_5132,N_4057,N_4486);
nor U5133 (N_5133,N_4206,N_4118);
nor U5134 (N_5134,N_4226,N_3950);
nor U5135 (N_5135,N_4049,N_4387);
nor U5136 (N_5136,N_4445,N_4417);
and U5137 (N_5137,N_4393,N_4295);
or U5138 (N_5138,N_4436,N_3883);
xor U5139 (N_5139,N_4369,N_4101);
and U5140 (N_5140,N_4197,N_3935);
nor U5141 (N_5141,N_4279,N_4197);
xor U5142 (N_5142,N_3858,N_4391);
nor U5143 (N_5143,N_4183,N_4412);
and U5144 (N_5144,N_4416,N_4015);
nor U5145 (N_5145,N_3801,N_3944);
xor U5146 (N_5146,N_3980,N_4481);
nor U5147 (N_5147,N_4215,N_4459);
or U5148 (N_5148,N_4156,N_3927);
and U5149 (N_5149,N_4204,N_4437);
nand U5150 (N_5150,N_3858,N_4423);
nand U5151 (N_5151,N_3761,N_4454);
nor U5152 (N_5152,N_4316,N_3857);
and U5153 (N_5153,N_4458,N_3839);
and U5154 (N_5154,N_3980,N_4296);
nor U5155 (N_5155,N_4472,N_3827);
nor U5156 (N_5156,N_3769,N_3934);
or U5157 (N_5157,N_4152,N_4160);
nand U5158 (N_5158,N_4442,N_3985);
nor U5159 (N_5159,N_4052,N_4110);
nand U5160 (N_5160,N_4125,N_4485);
xnor U5161 (N_5161,N_4472,N_3974);
nand U5162 (N_5162,N_4260,N_4402);
or U5163 (N_5163,N_3842,N_4199);
nand U5164 (N_5164,N_4450,N_4446);
nand U5165 (N_5165,N_3787,N_4348);
and U5166 (N_5166,N_4354,N_4120);
xnor U5167 (N_5167,N_3754,N_3791);
nand U5168 (N_5168,N_4264,N_3893);
or U5169 (N_5169,N_4167,N_4112);
nand U5170 (N_5170,N_4362,N_3942);
nand U5171 (N_5171,N_3769,N_3901);
or U5172 (N_5172,N_3868,N_3810);
xnor U5173 (N_5173,N_4296,N_4422);
or U5174 (N_5174,N_4283,N_4064);
and U5175 (N_5175,N_3786,N_4135);
or U5176 (N_5176,N_3965,N_4337);
nor U5177 (N_5177,N_4196,N_4392);
and U5178 (N_5178,N_4425,N_4497);
xnor U5179 (N_5179,N_4293,N_4414);
nand U5180 (N_5180,N_3891,N_4334);
nor U5181 (N_5181,N_4445,N_4269);
and U5182 (N_5182,N_4025,N_3944);
nand U5183 (N_5183,N_4258,N_3786);
nand U5184 (N_5184,N_4208,N_4163);
nor U5185 (N_5185,N_4324,N_4186);
xnor U5186 (N_5186,N_3839,N_3861);
nor U5187 (N_5187,N_3990,N_4070);
nor U5188 (N_5188,N_3759,N_4130);
nand U5189 (N_5189,N_4175,N_4364);
or U5190 (N_5190,N_3992,N_4303);
or U5191 (N_5191,N_3784,N_4109);
nor U5192 (N_5192,N_4207,N_3790);
or U5193 (N_5193,N_4188,N_4322);
or U5194 (N_5194,N_3947,N_4121);
xnor U5195 (N_5195,N_4022,N_4338);
nor U5196 (N_5196,N_4152,N_3963);
and U5197 (N_5197,N_4372,N_4242);
and U5198 (N_5198,N_4313,N_4069);
or U5199 (N_5199,N_4420,N_3920);
and U5200 (N_5200,N_4358,N_4226);
and U5201 (N_5201,N_4155,N_4301);
or U5202 (N_5202,N_3816,N_4393);
xor U5203 (N_5203,N_4498,N_4132);
nand U5204 (N_5204,N_3920,N_4116);
and U5205 (N_5205,N_4027,N_4357);
nor U5206 (N_5206,N_4375,N_4497);
nor U5207 (N_5207,N_4344,N_4389);
nand U5208 (N_5208,N_4291,N_4077);
nor U5209 (N_5209,N_4285,N_4088);
nor U5210 (N_5210,N_4317,N_3837);
nand U5211 (N_5211,N_4241,N_4201);
nand U5212 (N_5212,N_4463,N_4126);
xor U5213 (N_5213,N_3916,N_3786);
nor U5214 (N_5214,N_4303,N_4397);
and U5215 (N_5215,N_4488,N_4222);
nand U5216 (N_5216,N_4010,N_3855);
and U5217 (N_5217,N_4082,N_4427);
or U5218 (N_5218,N_4311,N_4435);
nand U5219 (N_5219,N_3856,N_4041);
nand U5220 (N_5220,N_3874,N_3918);
nand U5221 (N_5221,N_4425,N_3954);
nor U5222 (N_5222,N_3946,N_3866);
xor U5223 (N_5223,N_4126,N_4385);
nor U5224 (N_5224,N_3852,N_4143);
nand U5225 (N_5225,N_4015,N_4424);
or U5226 (N_5226,N_4102,N_4117);
or U5227 (N_5227,N_3800,N_4023);
nor U5228 (N_5228,N_3771,N_4187);
and U5229 (N_5229,N_4341,N_4372);
nand U5230 (N_5230,N_3851,N_4417);
and U5231 (N_5231,N_3919,N_3898);
nor U5232 (N_5232,N_3896,N_3867);
or U5233 (N_5233,N_4137,N_4096);
nand U5234 (N_5234,N_4319,N_4293);
xnor U5235 (N_5235,N_4132,N_3910);
and U5236 (N_5236,N_3954,N_3839);
nor U5237 (N_5237,N_3883,N_4001);
nor U5238 (N_5238,N_4433,N_3754);
and U5239 (N_5239,N_4442,N_4256);
xnor U5240 (N_5240,N_4380,N_3836);
or U5241 (N_5241,N_4449,N_4180);
and U5242 (N_5242,N_3933,N_3931);
nand U5243 (N_5243,N_4301,N_3936);
or U5244 (N_5244,N_4262,N_3871);
or U5245 (N_5245,N_3999,N_3755);
nor U5246 (N_5246,N_3790,N_4302);
xor U5247 (N_5247,N_4307,N_4346);
nand U5248 (N_5248,N_3884,N_4084);
nand U5249 (N_5249,N_4389,N_3805);
nand U5250 (N_5250,N_4751,N_5174);
or U5251 (N_5251,N_4780,N_4608);
nor U5252 (N_5252,N_4736,N_5004);
xnor U5253 (N_5253,N_5224,N_5147);
or U5254 (N_5254,N_4551,N_4941);
nand U5255 (N_5255,N_4837,N_5103);
and U5256 (N_5256,N_5124,N_4760);
and U5257 (N_5257,N_5222,N_5092);
or U5258 (N_5258,N_4718,N_5083);
or U5259 (N_5259,N_4516,N_4984);
nand U5260 (N_5260,N_4918,N_4985);
and U5261 (N_5261,N_5151,N_4892);
or U5262 (N_5262,N_4532,N_5178);
nor U5263 (N_5263,N_5243,N_4552);
xnor U5264 (N_5264,N_4631,N_4706);
and U5265 (N_5265,N_4740,N_4976);
and U5266 (N_5266,N_4715,N_4661);
and U5267 (N_5267,N_4783,N_5180);
nand U5268 (N_5268,N_5026,N_4929);
or U5269 (N_5269,N_4601,N_4630);
and U5270 (N_5270,N_4693,N_4928);
or U5271 (N_5271,N_5169,N_5015);
and U5272 (N_5272,N_5231,N_4714);
nor U5273 (N_5273,N_5138,N_5201);
and U5274 (N_5274,N_4776,N_4667);
nand U5275 (N_5275,N_4593,N_4959);
nand U5276 (N_5276,N_4906,N_5225);
and U5277 (N_5277,N_4807,N_4819);
nand U5278 (N_5278,N_5229,N_4996);
and U5279 (N_5279,N_4502,N_4778);
or U5280 (N_5280,N_4506,N_4610);
and U5281 (N_5281,N_5021,N_5086);
nand U5282 (N_5282,N_4820,N_5232);
or U5283 (N_5283,N_5055,N_5030);
and U5284 (N_5284,N_4901,N_4614);
and U5285 (N_5285,N_4803,N_4847);
nand U5286 (N_5286,N_5132,N_5117);
or U5287 (N_5287,N_5233,N_4798);
nand U5288 (N_5288,N_5023,N_4962);
or U5289 (N_5289,N_4720,N_4691);
or U5290 (N_5290,N_4843,N_5106);
or U5291 (N_5291,N_5212,N_5003);
and U5292 (N_5292,N_5007,N_4936);
xor U5293 (N_5293,N_4886,N_5108);
nor U5294 (N_5294,N_4653,N_5045);
nor U5295 (N_5295,N_4537,N_5089);
nor U5296 (N_5296,N_4851,N_5114);
nand U5297 (N_5297,N_4761,N_4951);
nor U5298 (N_5298,N_4569,N_4641);
nand U5299 (N_5299,N_4549,N_4701);
nor U5300 (N_5300,N_5079,N_4957);
nor U5301 (N_5301,N_4658,N_5054);
nand U5302 (N_5302,N_5125,N_5237);
or U5303 (N_5303,N_4811,N_4600);
nand U5304 (N_5304,N_4947,N_5064);
nand U5305 (N_5305,N_4595,N_4575);
nand U5306 (N_5306,N_4977,N_4559);
nand U5307 (N_5307,N_4932,N_5014);
or U5308 (N_5308,N_5056,N_4777);
nor U5309 (N_5309,N_4645,N_4558);
xor U5310 (N_5310,N_5129,N_5005);
and U5311 (N_5311,N_5139,N_4560);
or U5312 (N_5312,N_5149,N_4678);
or U5313 (N_5313,N_4562,N_4622);
nor U5314 (N_5314,N_5013,N_4915);
or U5315 (N_5315,N_4721,N_4530);
nand U5316 (N_5316,N_4746,N_5175);
nand U5317 (N_5317,N_4930,N_4881);
nor U5318 (N_5318,N_5146,N_4829);
or U5319 (N_5319,N_4876,N_4942);
and U5320 (N_5320,N_4756,N_4711);
xor U5321 (N_5321,N_4597,N_5241);
or U5322 (N_5322,N_4867,N_4578);
nor U5323 (N_5323,N_4836,N_5122);
and U5324 (N_5324,N_4913,N_4880);
or U5325 (N_5325,N_5183,N_4800);
xor U5326 (N_5326,N_5142,N_4612);
xor U5327 (N_5327,N_5027,N_4528);
nor U5328 (N_5328,N_4974,N_4512);
nor U5329 (N_5329,N_4543,N_5238);
or U5330 (N_5330,N_4589,N_4828);
or U5331 (N_5331,N_4742,N_4571);
nor U5332 (N_5332,N_4707,N_5105);
nand U5333 (N_5333,N_4853,N_5145);
nor U5334 (N_5334,N_4827,N_4663);
and U5335 (N_5335,N_5059,N_4660);
nor U5336 (N_5336,N_4577,N_4647);
nand U5337 (N_5337,N_4938,N_5182);
or U5338 (N_5338,N_4545,N_5185);
nor U5339 (N_5339,N_5155,N_4554);
and U5340 (N_5340,N_4627,N_5072);
or U5341 (N_5341,N_4970,N_4754);
and U5342 (N_5342,N_4940,N_4927);
nor U5343 (N_5343,N_5190,N_4538);
and U5344 (N_5344,N_5001,N_4665);
nor U5345 (N_5345,N_4649,N_4674);
nand U5346 (N_5346,N_4897,N_4914);
or U5347 (N_5347,N_4728,N_4770);
or U5348 (N_5348,N_5111,N_4685);
or U5349 (N_5349,N_4757,N_5050);
and U5350 (N_5350,N_4730,N_4534);
and U5351 (N_5351,N_5148,N_5066);
and U5352 (N_5352,N_4603,N_4689);
and U5353 (N_5353,N_5006,N_5172);
or U5354 (N_5354,N_4680,N_4511);
nor U5355 (N_5355,N_4990,N_4838);
and U5356 (N_5356,N_4500,N_4989);
or U5357 (N_5357,N_5100,N_4971);
nor U5358 (N_5358,N_4529,N_5235);
nor U5359 (N_5359,N_5017,N_4682);
or U5360 (N_5360,N_4594,N_5127);
xnor U5361 (N_5361,N_4619,N_4864);
or U5362 (N_5362,N_4869,N_4541);
nor U5363 (N_5363,N_5166,N_4854);
nand U5364 (N_5364,N_4925,N_5187);
nor U5365 (N_5365,N_4825,N_5074);
nor U5366 (N_5366,N_5248,N_5131);
nor U5367 (N_5367,N_4981,N_4615);
and U5368 (N_5368,N_5195,N_5084);
xnor U5369 (N_5369,N_5016,N_4686);
nor U5370 (N_5370,N_4894,N_4652);
and U5371 (N_5371,N_5215,N_4852);
nor U5372 (N_5372,N_5165,N_4911);
nor U5373 (N_5373,N_5011,N_4831);
nand U5374 (N_5374,N_5136,N_4968);
or U5375 (N_5375,N_4832,N_5249);
nand U5376 (N_5376,N_4873,N_4931);
nor U5377 (N_5377,N_4704,N_4912);
or U5378 (N_5378,N_4644,N_5159);
nand U5379 (N_5379,N_4697,N_4983);
and U5380 (N_5380,N_4584,N_4872);
nand U5381 (N_5381,N_4998,N_4802);
nand U5382 (N_5382,N_5034,N_4517);
or U5383 (N_5383,N_4585,N_4815);
nand U5384 (N_5384,N_5218,N_4963);
nand U5385 (N_5385,N_4710,N_4722);
and U5386 (N_5386,N_4969,N_4555);
or U5387 (N_5387,N_5219,N_5227);
nor U5388 (N_5388,N_4625,N_4592);
or U5389 (N_5389,N_5216,N_4564);
or U5390 (N_5390,N_4841,N_4893);
or U5391 (N_5391,N_4747,N_4596);
and U5392 (N_5392,N_4898,N_4743);
and U5393 (N_5393,N_4958,N_5120);
and U5394 (N_5394,N_5041,N_5170);
and U5395 (N_5395,N_4764,N_4514);
or U5396 (N_5396,N_5184,N_5000);
and U5397 (N_5397,N_4536,N_4733);
nor U5398 (N_5398,N_5012,N_4621);
nor U5399 (N_5399,N_4979,N_4810);
xor U5400 (N_5400,N_4548,N_4833);
or U5401 (N_5401,N_4888,N_4885);
nand U5402 (N_5402,N_4590,N_4945);
nor U5403 (N_5403,N_4671,N_4700);
nand U5404 (N_5404,N_5200,N_4848);
nand U5405 (N_5405,N_4823,N_5040);
or U5406 (N_5406,N_4961,N_5198);
nor U5407 (N_5407,N_5058,N_4973);
xnor U5408 (N_5408,N_5210,N_4527);
nand U5409 (N_5409,N_4890,N_4920);
or U5410 (N_5410,N_4698,N_5177);
and U5411 (N_5411,N_5186,N_5043);
nand U5412 (N_5412,N_4654,N_4870);
nand U5413 (N_5413,N_5053,N_5202);
xnor U5414 (N_5414,N_5093,N_4606);
xor U5415 (N_5415,N_5247,N_4907);
nor U5416 (N_5416,N_4568,N_5110);
xnor U5417 (N_5417,N_4524,N_4643);
xor U5418 (N_5418,N_4884,N_4818);
nor U5419 (N_5419,N_4813,N_4716);
xnor U5420 (N_5420,N_4503,N_4987);
and U5421 (N_5421,N_4767,N_4994);
nand U5422 (N_5422,N_4738,N_4975);
or U5423 (N_5423,N_4670,N_4581);
nand U5424 (N_5424,N_5221,N_4695);
xor U5425 (N_5425,N_4993,N_4900);
nand U5426 (N_5426,N_4570,N_4582);
nand U5427 (N_5427,N_4664,N_4874);
nand U5428 (N_5428,N_5206,N_4692);
and U5429 (N_5429,N_4574,N_4681);
nand U5430 (N_5430,N_5088,N_4895);
and U5431 (N_5431,N_4806,N_4879);
nor U5432 (N_5432,N_4588,N_5070);
nand U5433 (N_5433,N_4861,N_4626);
xnor U5434 (N_5434,N_4956,N_5140);
and U5435 (N_5435,N_4696,N_5236);
or U5436 (N_5436,N_4766,N_4840);
or U5437 (N_5437,N_5098,N_4683);
nand U5438 (N_5438,N_4955,N_4763);
nor U5439 (N_5439,N_4793,N_5246);
nand U5440 (N_5440,N_4690,N_4708);
xor U5441 (N_5441,N_4553,N_4639);
nand U5442 (N_5442,N_5168,N_4934);
nor U5443 (N_5443,N_4933,N_4850);
and U5444 (N_5444,N_4849,N_4978);
nand U5445 (N_5445,N_4583,N_4759);
xor U5446 (N_5446,N_4550,N_4732);
nor U5447 (N_5447,N_4673,N_5112);
and U5448 (N_5448,N_5102,N_4891);
xor U5449 (N_5449,N_4587,N_4679);
or U5450 (N_5450,N_5097,N_5028);
or U5451 (N_5451,N_4659,N_4839);
or U5452 (N_5452,N_5031,N_4773);
nand U5453 (N_5453,N_4817,N_5137);
and U5454 (N_5454,N_4666,N_4948);
and U5455 (N_5455,N_4628,N_5244);
and U5456 (N_5456,N_4926,N_4816);
and U5457 (N_5457,N_4518,N_4741);
nor U5458 (N_5458,N_5234,N_4781);
nor U5459 (N_5459,N_4949,N_5126);
or U5460 (N_5460,N_4633,N_4954);
and U5461 (N_5461,N_4808,N_4544);
and U5462 (N_5462,N_5068,N_4717);
or U5463 (N_5463,N_4795,N_5085);
and U5464 (N_5464,N_5203,N_5226);
or U5465 (N_5465,N_4967,N_4805);
nor U5466 (N_5466,N_4772,N_5157);
xor U5467 (N_5467,N_4771,N_4801);
or U5468 (N_5468,N_5029,N_4609);
or U5469 (N_5469,N_5022,N_4509);
xor U5470 (N_5470,N_5109,N_4713);
and U5471 (N_5471,N_5211,N_5194);
nor U5472 (N_5472,N_4507,N_4602);
and U5473 (N_5473,N_4765,N_5042);
or U5474 (N_5474,N_4782,N_4762);
nor U5475 (N_5475,N_4856,N_5193);
nor U5476 (N_5476,N_4557,N_4905);
nor U5477 (N_5477,N_5239,N_4917);
or U5478 (N_5478,N_5082,N_4877);
or U5479 (N_5479,N_5171,N_4526);
or U5480 (N_5480,N_4629,N_4919);
or U5481 (N_5481,N_5067,N_5130);
or U5482 (N_5482,N_5009,N_4943);
or U5483 (N_5483,N_5167,N_4635);
nand U5484 (N_5484,N_4573,N_4768);
nor U5485 (N_5485,N_4531,N_4889);
nor U5486 (N_5486,N_4785,N_4992);
or U5487 (N_5487,N_4676,N_4937);
and U5488 (N_5488,N_5077,N_5150);
nor U5489 (N_5489,N_5094,N_5008);
xnor U5490 (N_5490,N_5078,N_4657);
nand U5491 (N_5491,N_4788,N_4586);
nor U5492 (N_5492,N_5057,N_4519);
and U5493 (N_5493,N_4946,N_5128);
nor U5494 (N_5494,N_4579,N_5107);
nand U5495 (N_5495,N_4546,N_4774);
nor U5496 (N_5496,N_4855,N_4753);
nor U5497 (N_5497,N_4709,N_4991);
nor U5498 (N_5498,N_4752,N_4939);
or U5499 (N_5499,N_5134,N_5158);
and U5500 (N_5500,N_4640,N_5047);
nand U5501 (N_5501,N_4719,N_4637);
or U5502 (N_5502,N_5154,N_5228);
nand U5503 (N_5503,N_5035,N_4950);
xor U5504 (N_5504,N_5119,N_4623);
xnor U5505 (N_5505,N_4737,N_4896);
xnor U5506 (N_5506,N_5104,N_4505);
nand U5507 (N_5507,N_5063,N_5099);
nor U5508 (N_5508,N_4791,N_4522);
or U5509 (N_5509,N_4822,N_4547);
xnor U5510 (N_5510,N_4556,N_5173);
and U5511 (N_5511,N_5189,N_4824);
or U5512 (N_5512,N_5242,N_5071);
and U5513 (N_5513,N_4792,N_5118);
and U5514 (N_5514,N_4862,N_4540);
nand U5515 (N_5515,N_4769,N_4887);
nor U5516 (N_5516,N_4790,N_5204);
nand U5517 (N_5517,N_4668,N_5095);
nand U5518 (N_5518,N_4814,N_5135);
and U5519 (N_5519,N_5002,N_5069);
xnor U5520 (N_5520,N_4712,N_5076);
nand U5521 (N_5521,N_5153,N_4616);
nand U5522 (N_5522,N_5116,N_4703);
nand U5523 (N_5523,N_4875,N_4964);
and U5524 (N_5524,N_4857,N_4702);
nor U5525 (N_5525,N_5144,N_5101);
nand U5526 (N_5526,N_4842,N_4504);
and U5527 (N_5527,N_5192,N_5091);
or U5528 (N_5528,N_5188,N_5032);
and U5529 (N_5529,N_5113,N_4821);
or U5530 (N_5530,N_4669,N_4866);
nand U5531 (N_5531,N_4605,N_5181);
and U5532 (N_5532,N_5213,N_5196);
and U5533 (N_5533,N_4580,N_4804);
or U5534 (N_5534,N_4687,N_4699);
and U5535 (N_5535,N_5223,N_5230);
or U5536 (N_5536,N_4748,N_4909);
and U5537 (N_5537,N_4613,N_4749);
or U5538 (N_5538,N_4632,N_5061);
nand U5539 (N_5539,N_4986,N_5046);
xor U5540 (N_5540,N_5141,N_4750);
or U5541 (N_5541,N_5197,N_5176);
nor U5542 (N_5542,N_5123,N_5199);
or U5543 (N_5543,N_4539,N_4723);
or U5544 (N_5544,N_4863,N_4908);
and U5545 (N_5545,N_4944,N_4758);
nand U5546 (N_5546,N_5024,N_4520);
and U5547 (N_5547,N_4725,N_5019);
nand U5548 (N_5548,N_4830,N_5217);
or U5549 (N_5549,N_4904,N_5038);
nand U5550 (N_5550,N_4739,N_4501);
and U5551 (N_5551,N_4510,N_4789);
and U5552 (N_5552,N_4775,N_4794);
and U5553 (N_5553,N_4835,N_4724);
nor U5554 (N_5554,N_4899,N_4883);
nand U5555 (N_5555,N_5048,N_4618);
or U5556 (N_5556,N_4636,N_4634);
xor U5557 (N_5557,N_4642,N_5075);
xnor U5558 (N_5558,N_4858,N_5240);
nand U5559 (N_5559,N_5205,N_5025);
nor U5560 (N_5560,N_4980,N_4620);
and U5561 (N_5561,N_4521,N_4513);
nand U5562 (N_5562,N_5191,N_4735);
nor U5563 (N_5563,N_4672,N_4859);
and U5564 (N_5564,N_4744,N_4576);
and U5565 (N_5565,N_5062,N_4868);
or U5566 (N_5566,N_5052,N_4860);
nand U5567 (N_5567,N_4729,N_4982);
xnor U5568 (N_5568,N_4604,N_4965);
nand U5569 (N_5569,N_5208,N_4567);
xnor U5570 (N_5570,N_4655,N_4677);
and U5571 (N_5571,N_4997,N_4797);
or U5572 (N_5572,N_4542,N_4684);
nand U5573 (N_5573,N_4910,N_5065);
xor U5574 (N_5574,N_5207,N_4972);
nor U5575 (N_5575,N_5160,N_5096);
nor U5576 (N_5576,N_4865,N_4988);
and U5577 (N_5577,N_4523,N_4617);
nor U5578 (N_5578,N_5087,N_4565);
nor U5579 (N_5579,N_4882,N_5162);
or U5580 (N_5580,N_4675,N_4727);
and U5581 (N_5581,N_5220,N_5051);
nor U5582 (N_5582,N_4796,N_5163);
and U5583 (N_5583,N_4731,N_4572);
nand U5584 (N_5584,N_5143,N_4638);
and U5585 (N_5585,N_5133,N_4902);
nor U5586 (N_5586,N_4563,N_5179);
nand U5587 (N_5587,N_4662,N_4648);
nand U5588 (N_5588,N_4525,N_4960);
nand U5589 (N_5589,N_4834,N_4952);
or U5590 (N_5590,N_4812,N_5037);
or U5591 (N_5591,N_5214,N_5049);
and U5592 (N_5592,N_4688,N_4922);
nand U5593 (N_5593,N_4624,N_4694);
nor U5594 (N_5594,N_4826,N_5209);
nand U5595 (N_5595,N_4566,N_4745);
nor U5596 (N_5596,N_4726,N_4923);
and U5597 (N_5597,N_4787,N_5039);
or U5598 (N_5598,N_4846,N_5020);
and U5599 (N_5599,N_5090,N_5044);
nand U5600 (N_5600,N_4844,N_4646);
and U5601 (N_5601,N_5161,N_5010);
nand U5602 (N_5602,N_5060,N_4966);
and U5603 (N_5603,N_4871,N_5152);
nand U5604 (N_5604,N_4903,N_5018);
xnor U5605 (N_5605,N_5036,N_4779);
xnor U5606 (N_5606,N_4734,N_5033);
or U5607 (N_5607,N_4916,N_4809);
or U5608 (N_5608,N_4705,N_4995);
nand U5609 (N_5609,N_4561,N_5073);
nand U5610 (N_5610,N_4799,N_4784);
nor U5611 (N_5611,N_4786,N_4611);
nand U5612 (N_5612,N_4755,N_4515);
and U5613 (N_5613,N_4599,N_5164);
nand U5614 (N_5614,N_4535,N_5081);
xor U5615 (N_5615,N_5121,N_4533);
nor U5616 (N_5616,N_4999,N_4598);
nand U5617 (N_5617,N_5115,N_4508);
nand U5618 (N_5618,N_4924,N_4845);
nand U5619 (N_5619,N_5080,N_4921);
xor U5620 (N_5620,N_5245,N_4650);
nor U5621 (N_5621,N_4878,N_4953);
and U5622 (N_5622,N_4935,N_4656);
xor U5623 (N_5623,N_4651,N_4591);
xor U5624 (N_5624,N_4607,N_5156);
and U5625 (N_5625,N_4935,N_5139);
nand U5626 (N_5626,N_4846,N_4590);
and U5627 (N_5627,N_4586,N_4617);
and U5628 (N_5628,N_5171,N_4611);
and U5629 (N_5629,N_4726,N_5180);
or U5630 (N_5630,N_4673,N_5245);
nand U5631 (N_5631,N_4968,N_4870);
nand U5632 (N_5632,N_4837,N_5243);
or U5633 (N_5633,N_5198,N_4621);
nand U5634 (N_5634,N_5189,N_5016);
nor U5635 (N_5635,N_5175,N_5020);
and U5636 (N_5636,N_4829,N_5014);
nor U5637 (N_5637,N_4643,N_4579);
and U5638 (N_5638,N_4726,N_4869);
or U5639 (N_5639,N_5210,N_4515);
nor U5640 (N_5640,N_4773,N_5172);
nand U5641 (N_5641,N_4949,N_4862);
and U5642 (N_5642,N_4983,N_5040);
nand U5643 (N_5643,N_4650,N_4662);
nand U5644 (N_5644,N_5162,N_4608);
or U5645 (N_5645,N_5144,N_4730);
and U5646 (N_5646,N_4523,N_4546);
nand U5647 (N_5647,N_5126,N_4868);
nand U5648 (N_5648,N_4907,N_4872);
xnor U5649 (N_5649,N_5192,N_5042);
and U5650 (N_5650,N_5140,N_4645);
nand U5651 (N_5651,N_5082,N_4813);
or U5652 (N_5652,N_4652,N_4822);
nand U5653 (N_5653,N_4672,N_4988);
or U5654 (N_5654,N_5040,N_4816);
and U5655 (N_5655,N_4781,N_5210);
nor U5656 (N_5656,N_4838,N_4930);
or U5657 (N_5657,N_4837,N_4635);
or U5658 (N_5658,N_4823,N_4864);
nor U5659 (N_5659,N_4954,N_4792);
or U5660 (N_5660,N_4751,N_4680);
xor U5661 (N_5661,N_4889,N_5011);
nand U5662 (N_5662,N_4694,N_5069);
and U5663 (N_5663,N_4521,N_5173);
or U5664 (N_5664,N_4814,N_5193);
nor U5665 (N_5665,N_4928,N_5121);
and U5666 (N_5666,N_5232,N_4733);
nand U5667 (N_5667,N_4860,N_4817);
nand U5668 (N_5668,N_4916,N_4887);
or U5669 (N_5669,N_5071,N_4815);
nand U5670 (N_5670,N_5210,N_4837);
nor U5671 (N_5671,N_4732,N_4629);
and U5672 (N_5672,N_4689,N_4755);
nand U5673 (N_5673,N_4804,N_5082);
nor U5674 (N_5674,N_5006,N_4722);
and U5675 (N_5675,N_4713,N_4542);
nor U5676 (N_5676,N_4579,N_5021);
or U5677 (N_5677,N_4668,N_4591);
nand U5678 (N_5678,N_4752,N_5007);
and U5679 (N_5679,N_5212,N_4578);
nor U5680 (N_5680,N_4864,N_5206);
and U5681 (N_5681,N_4572,N_5135);
nor U5682 (N_5682,N_4641,N_4885);
nand U5683 (N_5683,N_4631,N_4810);
and U5684 (N_5684,N_5177,N_4960);
and U5685 (N_5685,N_4522,N_4781);
nor U5686 (N_5686,N_4900,N_5072);
or U5687 (N_5687,N_4672,N_4921);
xnor U5688 (N_5688,N_5103,N_5146);
nand U5689 (N_5689,N_5055,N_5159);
or U5690 (N_5690,N_4934,N_5178);
xor U5691 (N_5691,N_4977,N_4710);
and U5692 (N_5692,N_4904,N_4599);
xor U5693 (N_5693,N_4832,N_5177);
nor U5694 (N_5694,N_4772,N_5161);
or U5695 (N_5695,N_4940,N_4564);
or U5696 (N_5696,N_4681,N_5027);
and U5697 (N_5697,N_4758,N_5141);
or U5698 (N_5698,N_4606,N_4675);
and U5699 (N_5699,N_5059,N_4533);
nor U5700 (N_5700,N_4756,N_4988);
and U5701 (N_5701,N_5041,N_4657);
nor U5702 (N_5702,N_4594,N_4890);
nand U5703 (N_5703,N_4523,N_4606);
nand U5704 (N_5704,N_5090,N_4886);
nand U5705 (N_5705,N_4563,N_4664);
or U5706 (N_5706,N_5034,N_5091);
and U5707 (N_5707,N_5225,N_4869);
nand U5708 (N_5708,N_4666,N_4664);
nor U5709 (N_5709,N_5040,N_5186);
or U5710 (N_5710,N_4870,N_5067);
nor U5711 (N_5711,N_5214,N_4511);
nand U5712 (N_5712,N_4673,N_4534);
nand U5713 (N_5713,N_5105,N_4651);
nand U5714 (N_5714,N_4790,N_4555);
and U5715 (N_5715,N_4796,N_4800);
or U5716 (N_5716,N_4892,N_5012);
nor U5717 (N_5717,N_5089,N_4927);
nor U5718 (N_5718,N_5240,N_4812);
nand U5719 (N_5719,N_4720,N_5208);
nor U5720 (N_5720,N_4840,N_4538);
or U5721 (N_5721,N_4588,N_4884);
or U5722 (N_5722,N_4580,N_4567);
and U5723 (N_5723,N_4621,N_4702);
or U5724 (N_5724,N_5050,N_5195);
and U5725 (N_5725,N_4810,N_5212);
and U5726 (N_5726,N_4748,N_5018);
and U5727 (N_5727,N_4998,N_4994);
or U5728 (N_5728,N_4918,N_4821);
and U5729 (N_5729,N_4841,N_5165);
nor U5730 (N_5730,N_4870,N_4699);
nor U5731 (N_5731,N_4953,N_4581);
nand U5732 (N_5732,N_4742,N_4747);
nand U5733 (N_5733,N_4651,N_4905);
or U5734 (N_5734,N_5177,N_4688);
or U5735 (N_5735,N_4502,N_4504);
or U5736 (N_5736,N_5194,N_4681);
nor U5737 (N_5737,N_5123,N_5011);
nand U5738 (N_5738,N_5246,N_4771);
nor U5739 (N_5739,N_4942,N_4541);
nor U5740 (N_5740,N_4680,N_5209);
nor U5741 (N_5741,N_4808,N_5161);
and U5742 (N_5742,N_5200,N_4645);
nor U5743 (N_5743,N_4857,N_4917);
nor U5744 (N_5744,N_4841,N_4568);
nor U5745 (N_5745,N_4692,N_4553);
or U5746 (N_5746,N_5204,N_4701);
xor U5747 (N_5747,N_4767,N_5035);
nor U5748 (N_5748,N_5090,N_5108);
and U5749 (N_5749,N_4864,N_4672);
nor U5750 (N_5750,N_4559,N_5011);
and U5751 (N_5751,N_5244,N_5185);
nor U5752 (N_5752,N_4922,N_4959);
nor U5753 (N_5753,N_5082,N_5063);
nor U5754 (N_5754,N_5070,N_4863);
nand U5755 (N_5755,N_4800,N_5060);
nand U5756 (N_5756,N_4678,N_4605);
or U5757 (N_5757,N_4966,N_4982);
nand U5758 (N_5758,N_4890,N_4577);
xor U5759 (N_5759,N_4770,N_4805);
or U5760 (N_5760,N_4688,N_4780);
nor U5761 (N_5761,N_5223,N_5169);
or U5762 (N_5762,N_5193,N_4971);
or U5763 (N_5763,N_4516,N_4685);
nand U5764 (N_5764,N_4971,N_4865);
or U5765 (N_5765,N_4825,N_5167);
xnor U5766 (N_5766,N_4503,N_4618);
nand U5767 (N_5767,N_4971,N_4688);
or U5768 (N_5768,N_4593,N_5118);
nand U5769 (N_5769,N_4946,N_4798);
xnor U5770 (N_5770,N_4985,N_5077);
or U5771 (N_5771,N_4875,N_5066);
nand U5772 (N_5772,N_5185,N_4675);
nor U5773 (N_5773,N_4956,N_5138);
or U5774 (N_5774,N_4624,N_5070);
and U5775 (N_5775,N_5087,N_5068);
and U5776 (N_5776,N_4934,N_4963);
nor U5777 (N_5777,N_5025,N_4999);
nor U5778 (N_5778,N_5159,N_4792);
nor U5779 (N_5779,N_5210,N_5124);
nand U5780 (N_5780,N_4666,N_4801);
and U5781 (N_5781,N_4638,N_5110);
nor U5782 (N_5782,N_5025,N_4584);
or U5783 (N_5783,N_4745,N_4891);
xor U5784 (N_5784,N_5202,N_4827);
or U5785 (N_5785,N_4726,N_5093);
nor U5786 (N_5786,N_4515,N_4670);
and U5787 (N_5787,N_4884,N_5160);
nand U5788 (N_5788,N_4753,N_5091);
and U5789 (N_5789,N_5020,N_5114);
nand U5790 (N_5790,N_4558,N_4778);
nand U5791 (N_5791,N_4914,N_4510);
nor U5792 (N_5792,N_4574,N_5135);
or U5793 (N_5793,N_4711,N_5160);
or U5794 (N_5794,N_4772,N_4677);
nand U5795 (N_5795,N_4693,N_5093);
nor U5796 (N_5796,N_4517,N_4951);
and U5797 (N_5797,N_5156,N_4604);
nor U5798 (N_5798,N_5061,N_4775);
or U5799 (N_5799,N_4570,N_5242);
nor U5800 (N_5800,N_4620,N_5113);
nand U5801 (N_5801,N_4541,N_5045);
or U5802 (N_5802,N_4767,N_4939);
nor U5803 (N_5803,N_4730,N_5228);
nor U5804 (N_5804,N_5049,N_4979);
nor U5805 (N_5805,N_4954,N_5003);
and U5806 (N_5806,N_4873,N_5174);
nand U5807 (N_5807,N_5028,N_5227);
xnor U5808 (N_5808,N_4731,N_4574);
and U5809 (N_5809,N_5005,N_5141);
xnor U5810 (N_5810,N_4802,N_5040);
and U5811 (N_5811,N_4618,N_4848);
and U5812 (N_5812,N_5083,N_4882);
nand U5813 (N_5813,N_4753,N_4826);
xor U5814 (N_5814,N_4634,N_5141);
xor U5815 (N_5815,N_5210,N_5067);
and U5816 (N_5816,N_4769,N_5222);
nor U5817 (N_5817,N_4809,N_5029);
and U5818 (N_5818,N_4553,N_5099);
or U5819 (N_5819,N_5072,N_5064);
and U5820 (N_5820,N_4657,N_4698);
or U5821 (N_5821,N_5131,N_4607);
nand U5822 (N_5822,N_4510,N_4979);
and U5823 (N_5823,N_4735,N_4771);
and U5824 (N_5824,N_4846,N_4915);
or U5825 (N_5825,N_4856,N_4889);
or U5826 (N_5826,N_5231,N_4576);
and U5827 (N_5827,N_4518,N_5115);
nor U5828 (N_5828,N_4853,N_4886);
or U5829 (N_5829,N_4912,N_5200);
nor U5830 (N_5830,N_5004,N_4668);
nor U5831 (N_5831,N_4597,N_4533);
or U5832 (N_5832,N_4840,N_4731);
nor U5833 (N_5833,N_4509,N_5132);
nand U5834 (N_5834,N_5049,N_4543);
nand U5835 (N_5835,N_4670,N_4521);
xor U5836 (N_5836,N_4976,N_4993);
nor U5837 (N_5837,N_5208,N_4843);
and U5838 (N_5838,N_4718,N_4888);
xnor U5839 (N_5839,N_4687,N_4876);
xor U5840 (N_5840,N_5202,N_4512);
nand U5841 (N_5841,N_4685,N_5024);
and U5842 (N_5842,N_5107,N_4644);
or U5843 (N_5843,N_5186,N_5114);
nand U5844 (N_5844,N_4817,N_4898);
xnor U5845 (N_5845,N_4881,N_4653);
and U5846 (N_5846,N_5008,N_4807);
or U5847 (N_5847,N_5164,N_5158);
nand U5848 (N_5848,N_4819,N_5167);
or U5849 (N_5849,N_4937,N_4933);
nor U5850 (N_5850,N_4755,N_5091);
xor U5851 (N_5851,N_4876,N_5147);
xnor U5852 (N_5852,N_5016,N_4675);
nand U5853 (N_5853,N_4789,N_5043);
and U5854 (N_5854,N_5209,N_4897);
or U5855 (N_5855,N_4705,N_5003);
nand U5856 (N_5856,N_5102,N_4988);
nand U5857 (N_5857,N_4907,N_5139);
nand U5858 (N_5858,N_4952,N_4814);
or U5859 (N_5859,N_4627,N_4886);
nand U5860 (N_5860,N_4919,N_4536);
and U5861 (N_5861,N_4993,N_4799);
and U5862 (N_5862,N_4539,N_5009);
and U5863 (N_5863,N_4539,N_4778);
nor U5864 (N_5864,N_4853,N_4865);
or U5865 (N_5865,N_5172,N_5141);
nor U5866 (N_5866,N_4587,N_4762);
nor U5867 (N_5867,N_4656,N_5170);
and U5868 (N_5868,N_4956,N_4650);
nor U5869 (N_5869,N_4978,N_4971);
and U5870 (N_5870,N_4740,N_5035);
and U5871 (N_5871,N_4955,N_4962);
nor U5872 (N_5872,N_4943,N_4696);
or U5873 (N_5873,N_4594,N_4848);
and U5874 (N_5874,N_4781,N_5133);
or U5875 (N_5875,N_4824,N_4523);
nand U5876 (N_5876,N_5187,N_5179);
or U5877 (N_5877,N_4736,N_5175);
xor U5878 (N_5878,N_4748,N_4910);
nor U5879 (N_5879,N_4624,N_5239);
nand U5880 (N_5880,N_4914,N_4983);
or U5881 (N_5881,N_4785,N_4871);
xnor U5882 (N_5882,N_4603,N_5174);
or U5883 (N_5883,N_4606,N_4789);
nand U5884 (N_5884,N_4644,N_4872);
nand U5885 (N_5885,N_4624,N_4707);
nand U5886 (N_5886,N_4517,N_4961);
and U5887 (N_5887,N_5042,N_5248);
xor U5888 (N_5888,N_4953,N_4957);
nand U5889 (N_5889,N_4808,N_4888);
and U5890 (N_5890,N_4865,N_4819);
and U5891 (N_5891,N_4916,N_4832);
xnor U5892 (N_5892,N_4799,N_5056);
nand U5893 (N_5893,N_4832,N_4845);
nand U5894 (N_5894,N_5095,N_4813);
nor U5895 (N_5895,N_4607,N_4732);
and U5896 (N_5896,N_4663,N_4574);
and U5897 (N_5897,N_4771,N_4604);
or U5898 (N_5898,N_5128,N_5101);
or U5899 (N_5899,N_5194,N_5074);
nor U5900 (N_5900,N_5089,N_4888);
nor U5901 (N_5901,N_4514,N_4545);
nand U5902 (N_5902,N_4570,N_5213);
xnor U5903 (N_5903,N_4788,N_5021);
or U5904 (N_5904,N_4976,N_4512);
nor U5905 (N_5905,N_5126,N_5131);
and U5906 (N_5906,N_4884,N_4735);
and U5907 (N_5907,N_5057,N_4536);
nand U5908 (N_5908,N_4932,N_4640);
nand U5909 (N_5909,N_4808,N_5172);
nand U5910 (N_5910,N_4584,N_5220);
nor U5911 (N_5911,N_4861,N_4579);
nand U5912 (N_5912,N_4961,N_4881);
and U5913 (N_5913,N_4607,N_4705);
or U5914 (N_5914,N_4714,N_5083);
nor U5915 (N_5915,N_5052,N_5039);
and U5916 (N_5916,N_5206,N_5244);
or U5917 (N_5917,N_4953,N_4958);
or U5918 (N_5918,N_5225,N_4950);
or U5919 (N_5919,N_4753,N_5183);
nor U5920 (N_5920,N_5228,N_5033);
and U5921 (N_5921,N_4641,N_4799);
nand U5922 (N_5922,N_5097,N_4573);
nor U5923 (N_5923,N_4632,N_4528);
or U5924 (N_5924,N_4661,N_4959);
nand U5925 (N_5925,N_4671,N_4784);
or U5926 (N_5926,N_4982,N_4862);
or U5927 (N_5927,N_4666,N_5061);
nand U5928 (N_5928,N_5204,N_5085);
nor U5929 (N_5929,N_5106,N_4728);
and U5930 (N_5930,N_4570,N_4738);
xor U5931 (N_5931,N_4708,N_5049);
and U5932 (N_5932,N_4923,N_4957);
nor U5933 (N_5933,N_4678,N_4558);
or U5934 (N_5934,N_5199,N_4932);
nor U5935 (N_5935,N_4722,N_4844);
nor U5936 (N_5936,N_4881,N_5217);
nand U5937 (N_5937,N_5016,N_5122);
nand U5938 (N_5938,N_5118,N_5026);
xnor U5939 (N_5939,N_5133,N_4861);
and U5940 (N_5940,N_4943,N_4547);
nor U5941 (N_5941,N_4513,N_4647);
and U5942 (N_5942,N_4939,N_4897);
nor U5943 (N_5943,N_4980,N_5005);
xor U5944 (N_5944,N_5125,N_4502);
nand U5945 (N_5945,N_4857,N_5240);
or U5946 (N_5946,N_5024,N_5149);
xnor U5947 (N_5947,N_4540,N_4576);
nor U5948 (N_5948,N_5050,N_4516);
or U5949 (N_5949,N_4740,N_4677);
xor U5950 (N_5950,N_4696,N_5123);
nor U5951 (N_5951,N_4753,N_5066);
nor U5952 (N_5952,N_4567,N_5053);
nand U5953 (N_5953,N_4774,N_5186);
or U5954 (N_5954,N_5036,N_4657);
or U5955 (N_5955,N_5165,N_5158);
xor U5956 (N_5956,N_4988,N_4912);
nor U5957 (N_5957,N_4690,N_4944);
nor U5958 (N_5958,N_5191,N_4694);
nor U5959 (N_5959,N_4707,N_5122);
and U5960 (N_5960,N_4725,N_4685);
nor U5961 (N_5961,N_4968,N_4597);
and U5962 (N_5962,N_5211,N_5217);
or U5963 (N_5963,N_5097,N_4646);
xor U5964 (N_5964,N_4584,N_4561);
nor U5965 (N_5965,N_4578,N_5146);
or U5966 (N_5966,N_4524,N_5111);
and U5967 (N_5967,N_4507,N_4869);
nor U5968 (N_5968,N_5149,N_4987);
nor U5969 (N_5969,N_5142,N_4893);
nand U5970 (N_5970,N_4819,N_4581);
or U5971 (N_5971,N_5132,N_5068);
or U5972 (N_5972,N_5067,N_5199);
and U5973 (N_5973,N_4922,N_4631);
or U5974 (N_5974,N_4572,N_4529);
nand U5975 (N_5975,N_4985,N_4962);
and U5976 (N_5976,N_4692,N_4784);
nor U5977 (N_5977,N_5188,N_4935);
or U5978 (N_5978,N_4700,N_4524);
and U5979 (N_5979,N_4543,N_4691);
and U5980 (N_5980,N_5126,N_4871);
nand U5981 (N_5981,N_4805,N_4650);
nor U5982 (N_5982,N_4725,N_4888);
nor U5983 (N_5983,N_4721,N_5027);
nand U5984 (N_5984,N_4695,N_4987);
or U5985 (N_5985,N_5046,N_5153);
nand U5986 (N_5986,N_5101,N_4569);
and U5987 (N_5987,N_4957,N_4839);
nor U5988 (N_5988,N_5135,N_4990);
nand U5989 (N_5989,N_4720,N_5109);
nand U5990 (N_5990,N_4515,N_4656);
nor U5991 (N_5991,N_4878,N_4808);
and U5992 (N_5992,N_4872,N_5121);
and U5993 (N_5993,N_4871,N_4597);
nor U5994 (N_5994,N_5226,N_4939);
nor U5995 (N_5995,N_4503,N_4947);
xnor U5996 (N_5996,N_4619,N_4539);
nor U5997 (N_5997,N_4740,N_5138);
xor U5998 (N_5998,N_4846,N_4689);
and U5999 (N_5999,N_4921,N_4980);
nand U6000 (N_6000,N_5685,N_5303);
and U6001 (N_6001,N_5547,N_5436);
and U6002 (N_6002,N_5360,N_5649);
or U6003 (N_6003,N_5383,N_5763);
nor U6004 (N_6004,N_5972,N_5560);
nand U6005 (N_6005,N_5962,N_5361);
or U6006 (N_6006,N_5334,N_5565);
and U6007 (N_6007,N_5716,N_5664);
or U6008 (N_6008,N_5680,N_5590);
xnor U6009 (N_6009,N_5250,N_5617);
xor U6010 (N_6010,N_5351,N_5901);
nand U6011 (N_6011,N_5600,N_5465);
nor U6012 (N_6012,N_5672,N_5729);
or U6013 (N_6013,N_5792,N_5586);
nor U6014 (N_6014,N_5994,N_5985);
and U6015 (N_6015,N_5750,N_5924);
or U6016 (N_6016,N_5342,N_5853);
or U6017 (N_6017,N_5689,N_5414);
and U6018 (N_6018,N_5724,N_5842);
and U6019 (N_6019,N_5885,N_5272);
and U6020 (N_6020,N_5953,N_5951);
nor U6021 (N_6021,N_5467,N_5711);
nand U6022 (N_6022,N_5538,N_5873);
nand U6023 (N_6023,N_5852,N_5432);
or U6024 (N_6024,N_5898,N_5278);
or U6025 (N_6025,N_5738,N_5984);
or U6026 (N_6026,N_5682,N_5356);
nor U6027 (N_6027,N_5251,N_5535);
nand U6028 (N_6028,N_5376,N_5616);
nor U6029 (N_6029,N_5411,N_5948);
nor U6030 (N_6030,N_5752,N_5270);
or U6031 (N_6031,N_5891,N_5266);
and U6032 (N_6032,N_5942,N_5338);
and U6033 (N_6033,N_5983,N_5470);
nand U6034 (N_6034,N_5587,N_5969);
and U6035 (N_6035,N_5654,N_5773);
nand U6036 (N_6036,N_5859,N_5490);
and U6037 (N_6037,N_5323,N_5715);
nand U6038 (N_6038,N_5622,N_5778);
and U6039 (N_6039,N_5960,N_5977);
or U6040 (N_6040,N_5572,N_5605);
nor U6041 (N_6041,N_5700,N_5869);
xnor U6042 (N_6042,N_5775,N_5402);
and U6043 (N_6043,N_5895,N_5370);
nor U6044 (N_6044,N_5692,N_5974);
and U6045 (N_6045,N_5451,N_5846);
nand U6046 (N_6046,N_5422,N_5982);
nor U6047 (N_6047,N_5786,N_5283);
or U6048 (N_6048,N_5987,N_5428);
nor U6049 (N_6049,N_5871,N_5755);
nor U6050 (N_6050,N_5326,N_5771);
nor U6051 (N_6051,N_5311,N_5868);
nand U6052 (N_6052,N_5922,N_5263);
nor U6053 (N_6053,N_5282,N_5379);
nor U6054 (N_6054,N_5849,N_5657);
nand U6055 (N_6055,N_5667,N_5346);
or U6056 (N_6056,N_5997,N_5843);
and U6057 (N_6057,N_5992,N_5978);
nor U6058 (N_6058,N_5726,N_5864);
nand U6059 (N_6059,N_5772,N_5947);
nand U6060 (N_6060,N_5335,N_5909);
or U6061 (N_6061,N_5980,N_5395);
nand U6062 (N_6062,N_5485,N_5830);
or U6063 (N_6063,N_5517,N_5495);
and U6064 (N_6064,N_5855,N_5364);
and U6065 (N_6065,N_5387,N_5284);
xnor U6066 (N_6066,N_5513,N_5502);
or U6067 (N_6067,N_5486,N_5366);
or U6068 (N_6068,N_5975,N_5653);
or U6069 (N_6069,N_5449,N_5269);
nand U6070 (N_6070,N_5965,N_5769);
nor U6071 (N_6071,N_5807,N_5296);
and U6072 (N_6072,N_5404,N_5615);
nand U6073 (N_6073,N_5641,N_5642);
or U6074 (N_6074,N_5723,N_5998);
and U6075 (N_6075,N_5971,N_5814);
nor U6076 (N_6076,N_5584,N_5999);
or U6077 (N_6077,N_5375,N_5803);
nand U6078 (N_6078,N_5276,N_5986);
and U6079 (N_6079,N_5882,N_5546);
or U6080 (N_6080,N_5524,N_5443);
nor U6081 (N_6081,N_5452,N_5363);
and U6082 (N_6082,N_5591,N_5583);
and U6083 (N_6083,N_5904,N_5493);
or U6084 (N_6084,N_5620,N_5645);
nor U6085 (N_6085,N_5579,N_5848);
nor U6086 (N_6086,N_5862,N_5844);
and U6087 (N_6087,N_5448,N_5804);
nand U6088 (N_6088,N_5952,N_5606);
xnor U6089 (N_6089,N_5408,N_5856);
and U6090 (N_6090,N_5439,N_5393);
or U6091 (N_6091,N_5783,N_5374);
nor U6092 (N_6092,N_5480,N_5525);
or U6093 (N_6093,N_5993,N_5446);
xnor U6094 (N_6094,N_5325,N_5888);
or U6095 (N_6095,N_5371,N_5706);
and U6096 (N_6096,N_5889,N_5795);
and U6097 (N_6097,N_5258,N_5310);
xnor U6098 (N_6098,N_5466,N_5610);
nand U6099 (N_6099,N_5900,N_5267);
xnor U6100 (N_6100,N_5883,N_5793);
nand U6101 (N_6101,N_5823,N_5825);
and U6102 (N_6102,N_5633,N_5556);
and U6103 (N_6103,N_5400,N_5568);
xnor U6104 (N_6104,N_5594,N_5821);
nand U6105 (N_6105,N_5462,N_5934);
nand U6106 (N_6106,N_5920,N_5936);
nor U6107 (N_6107,N_5759,N_5413);
xor U6108 (N_6108,N_5968,N_5317);
nand U6109 (N_6109,N_5718,N_5384);
nor U6110 (N_6110,N_5892,N_5382);
xnor U6111 (N_6111,N_5939,N_5932);
or U6112 (N_6112,N_5614,N_5827);
and U6113 (N_6113,N_5813,N_5746);
nand U6114 (N_6114,N_5421,N_5324);
nor U6115 (N_6115,N_5697,N_5429);
nor U6116 (N_6116,N_5253,N_5801);
nand U6117 (N_6117,N_5959,N_5914);
nand U6118 (N_6118,N_5320,N_5693);
nand U6119 (N_6119,N_5259,N_5412);
nand U6120 (N_6120,N_5355,N_5285);
and U6121 (N_6121,N_5673,N_5534);
or U6122 (N_6122,N_5604,N_5354);
nor U6123 (N_6123,N_5703,N_5511);
nor U6124 (N_6124,N_5442,N_5650);
nor U6125 (N_6125,N_5659,N_5656);
nor U6126 (N_6126,N_5760,N_5911);
and U6127 (N_6127,N_5423,N_5540);
nand U6128 (N_6128,N_5543,N_5841);
nor U6129 (N_6129,N_5808,N_5899);
xnor U6130 (N_6130,N_5867,N_5958);
nor U6131 (N_6131,N_5598,N_5418);
or U6132 (N_6132,N_5399,N_5676);
nor U6133 (N_6133,N_5854,N_5567);
and U6134 (N_6134,N_5728,N_5555);
nor U6135 (N_6135,N_5532,N_5306);
or U6136 (N_6136,N_5632,N_5964);
or U6137 (N_6137,N_5950,N_5782);
and U6138 (N_6138,N_5407,N_5608);
or U6139 (N_6139,N_5277,N_5410);
nand U6140 (N_6140,N_5471,N_5696);
nand U6141 (N_6141,N_5928,N_5489);
nand U6142 (N_6142,N_5339,N_5787);
nand U6143 (N_6143,N_5780,N_5530);
and U6144 (N_6144,N_5357,N_5835);
or U6145 (N_6145,N_5739,N_5589);
or U6146 (N_6146,N_5397,N_5595);
or U6147 (N_6147,N_5698,N_5621);
and U6148 (N_6148,N_5943,N_5581);
or U6149 (N_6149,N_5549,N_5537);
nor U6150 (N_6150,N_5341,N_5553);
or U6151 (N_6151,N_5686,N_5764);
nor U6152 (N_6152,N_5955,N_5596);
nor U6153 (N_6153,N_5905,N_5450);
or U6154 (N_6154,N_5880,N_5369);
or U6155 (N_6155,N_5327,N_5995);
or U6156 (N_6156,N_5926,N_5874);
or U6157 (N_6157,N_5967,N_5679);
or U6158 (N_6158,N_5903,N_5603);
xor U6159 (N_6159,N_5458,N_5720);
nor U6160 (N_6160,N_5508,N_5619);
and U6161 (N_6161,N_5761,N_5732);
xor U6162 (N_6162,N_5463,N_5352);
nand U6163 (N_6163,N_5996,N_5607);
nand U6164 (N_6164,N_5504,N_5754);
nor U6165 (N_6165,N_5318,N_5365);
or U6166 (N_6166,N_5802,N_5561);
nand U6167 (N_6167,N_5748,N_5275);
or U6168 (N_6168,N_5643,N_5637);
nand U6169 (N_6169,N_5315,N_5368);
nor U6170 (N_6170,N_5665,N_5435);
xnor U6171 (N_6171,N_5714,N_5510);
nand U6172 (N_6172,N_5392,N_5858);
or U6173 (N_6173,N_5624,N_5389);
nor U6174 (N_6174,N_5481,N_5788);
nand U6175 (N_6175,N_5295,N_5668);
and U6176 (N_6176,N_5850,N_5488);
or U6177 (N_6177,N_5690,N_5694);
nor U6178 (N_6178,N_5536,N_5312);
nand U6179 (N_6179,N_5332,N_5479);
and U6180 (N_6180,N_5945,N_5290);
and U6181 (N_6181,N_5819,N_5734);
nand U6182 (N_6182,N_5875,N_5349);
and U6183 (N_6183,N_5940,N_5851);
nor U6184 (N_6184,N_5469,N_5721);
and U6185 (N_6185,N_5287,N_5430);
nor U6186 (N_6186,N_5518,N_5743);
xor U6187 (N_6187,N_5662,N_5826);
nor U6188 (N_6188,N_5316,N_5288);
nand U6189 (N_6189,N_5837,N_5491);
xnor U6190 (N_6190,N_5805,N_5331);
xor U6191 (N_6191,N_5628,N_5963);
nand U6192 (N_6192,N_5730,N_5500);
or U6193 (N_6193,N_5709,N_5542);
nor U6194 (N_6194,N_5625,N_5663);
and U6195 (N_6195,N_5539,N_5731);
or U6196 (N_6196,N_5879,N_5767);
xnor U6197 (N_6197,N_5564,N_5477);
nor U6198 (N_6198,N_5329,N_5476);
or U6199 (N_6199,N_5260,N_5487);
nand U6200 (N_6200,N_5529,N_5261);
nand U6201 (N_6201,N_5915,N_5737);
nand U6202 (N_6202,N_5523,N_5824);
nor U6203 (N_6203,N_5669,N_5431);
and U6204 (N_6204,N_5990,N_5319);
nand U6205 (N_6205,N_5507,N_5520);
nor U6206 (N_6206,N_5330,N_5478);
and U6207 (N_6207,N_5459,N_5293);
nand U6208 (N_6208,N_5946,N_5434);
and U6209 (N_6209,N_5255,N_5509);
and U6210 (N_6210,N_5699,N_5897);
or U6211 (N_6211,N_5298,N_5725);
xnor U6212 (N_6212,N_5710,N_5747);
or U6213 (N_6213,N_5403,N_5966);
and U6214 (N_6214,N_5712,N_5935);
and U6215 (N_6215,N_5372,N_5585);
and U6216 (N_6216,N_5877,N_5806);
nor U6217 (N_6217,N_5636,N_5497);
xnor U6218 (N_6218,N_5956,N_5521);
nor U6219 (N_6219,N_5790,N_5655);
or U6220 (N_6220,N_5313,N_5860);
or U6221 (N_6221,N_5822,N_5834);
nor U6222 (N_6222,N_5286,N_5575);
or U6223 (N_6223,N_5401,N_5516);
nor U6224 (N_6224,N_5713,N_5702);
nand U6225 (N_6225,N_5333,N_5563);
nand U6226 (N_6226,N_5777,N_5321);
or U6227 (N_6227,N_5727,N_5758);
and U6228 (N_6228,N_5762,N_5291);
or U6229 (N_6229,N_5776,N_5558);
nand U6230 (N_6230,N_5816,N_5570);
xor U6231 (N_6231,N_5496,N_5279);
or U6232 (N_6232,N_5840,N_5256);
xor U6233 (N_6233,N_5809,N_5612);
nand U6234 (N_6234,N_5917,N_5390);
nor U6235 (N_6235,N_5409,N_5406);
nor U6236 (N_6236,N_5944,N_5774);
or U6237 (N_6237,N_5574,N_5475);
and U6238 (N_6238,N_5639,N_5427);
nor U6239 (N_6239,N_5571,N_5501);
and U6240 (N_6240,N_5906,N_5578);
and U6241 (N_6241,N_5756,N_5894);
or U6242 (N_6242,N_5949,N_5740);
nand U6243 (N_6243,N_5681,N_5602);
nor U6244 (N_6244,N_5863,N_5677);
nor U6245 (N_6245,N_5519,N_5722);
and U6246 (N_6246,N_5265,N_5815);
nand U6247 (N_6247,N_5927,N_5811);
and U6248 (N_6248,N_5550,N_5661);
nand U6249 (N_6249,N_5799,N_5405);
or U6250 (N_6250,N_5751,N_5957);
and U6251 (N_6251,N_5593,N_5601);
nor U6252 (N_6252,N_5988,N_5770);
nand U6253 (N_6253,N_5380,N_5441);
and U6254 (N_6254,N_5872,N_5415);
xnor U6255 (N_6255,N_5857,N_5343);
nor U6256 (N_6256,N_5847,N_5300);
or U6257 (N_6257,N_5833,N_5791);
nor U6258 (N_6258,N_5396,N_5828);
and U6259 (N_6259,N_5766,N_5464);
nand U6260 (N_6260,N_5970,N_5580);
xnor U6261 (N_6261,N_5551,N_5832);
xor U6262 (N_6262,N_5425,N_5781);
nor U6263 (N_6263,N_5736,N_5741);
or U6264 (N_6264,N_5800,N_5559);
nand U6265 (N_6265,N_5634,N_5498);
or U6266 (N_6266,N_5933,N_5257);
and U6267 (N_6267,N_5254,N_5627);
xnor U6268 (N_6268,N_5707,N_5337);
or U6269 (N_6269,N_5907,N_5618);
xor U6270 (N_6270,N_5635,N_5347);
nor U6271 (N_6271,N_5494,N_5573);
nand U6272 (N_6272,N_5444,N_5908);
nor U6273 (N_6273,N_5302,N_5708);
xnor U6274 (N_6274,N_5308,N_5492);
and U6275 (N_6275,N_5447,N_5954);
nor U6276 (N_6276,N_5309,N_5268);
nor U6277 (N_6277,N_5297,N_5362);
or U6278 (N_6278,N_5328,N_5626);
nor U6279 (N_6279,N_5789,N_5902);
and U6280 (N_6280,N_5742,N_5640);
nand U6281 (N_6281,N_5701,N_5544);
nor U6282 (N_6282,N_5870,N_5599);
nor U6283 (N_6283,N_5890,N_5528);
or U6284 (N_6284,N_5886,N_5353);
xor U6285 (N_6285,N_5515,N_5541);
or U6286 (N_6286,N_5989,N_5658);
and U6287 (N_6287,N_5630,N_5836);
nand U6288 (N_6288,N_5503,N_5385);
or U6289 (N_6289,N_5735,N_5381);
xor U6290 (N_6290,N_5651,N_5744);
nand U6291 (N_6291,N_5919,N_5301);
or U6292 (N_6292,N_5484,N_5545);
and U6293 (N_6293,N_5929,N_5271);
nand U6294 (N_6294,N_5893,N_5812);
or U6295 (N_6295,N_5457,N_5533);
or U6296 (N_6296,N_5262,N_5916);
nand U6297 (N_6297,N_5930,N_5461);
and U6298 (N_6298,N_5569,N_5424);
nor U6299 (N_6299,N_5609,N_5386);
and U6300 (N_6300,N_5784,N_5440);
or U6301 (N_6301,N_5684,N_5820);
or U6302 (N_6302,N_5912,N_5839);
nor U6303 (N_6303,N_5512,N_5878);
nand U6304 (N_6304,N_5644,N_5252);
or U6305 (N_6305,N_5981,N_5582);
or U6306 (N_6306,N_5456,N_5548);
nand U6307 (N_6307,N_5896,N_5797);
and U6308 (N_6308,N_5884,N_5377);
and U6309 (N_6309,N_5671,N_5292);
and U6310 (N_6310,N_5705,N_5348);
nor U6311 (N_6311,N_5433,N_5941);
and U6312 (N_6312,N_5367,N_5876);
nand U6313 (N_6313,N_5264,N_5588);
and U6314 (N_6314,N_5861,N_5675);
nand U6315 (N_6315,N_5838,N_5526);
or U6316 (N_6316,N_5314,N_5473);
or U6317 (N_6317,N_5280,N_5391);
and U6318 (N_6318,N_5910,N_5938);
or U6319 (N_6319,N_5695,N_5416);
and U6320 (N_6320,N_5831,N_5866);
and U6321 (N_6321,N_5829,N_5281);
and U6322 (N_6322,N_5704,N_5420);
xnor U6323 (N_6323,N_5674,N_5937);
nand U6324 (N_6324,N_5768,N_5753);
xnor U6325 (N_6325,N_5505,N_5289);
xor U6326 (N_6326,N_5666,N_5394);
nor U6327 (N_6327,N_5683,N_5358);
or U6328 (N_6328,N_5438,N_5398);
nand U6329 (N_6329,N_5344,N_5388);
and U6330 (N_6330,N_5566,N_5522);
nor U6331 (N_6331,N_5373,N_5794);
and U6332 (N_6332,N_5638,N_5322);
and U6333 (N_6333,N_5976,N_5817);
nand U6334 (N_6334,N_5453,N_5881);
nand U6335 (N_6335,N_5345,N_5445);
and U6336 (N_6336,N_5991,N_5648);
nor U6337 (N_6337,N_5796,N_5597);
nor U6338 (N_6338,N_5765,N_5785);
nor U6339 (N_6339,N_5455,N_5454);
or U6340 (N_6340,N_5918,N_5307);
xor U6341 (N_6341,N_5273,N_5474);
nor U6342 (N_6342,N_5426,N_5460);
and U6343 (N_6343,N_5745,N_5554);
and U6344 (N_6344,N_5670,N_5688);
or U6345 (N_6345,N_5818,N_5629);
xor U6346 (N_6346,N_5961,N_5865);
xnor U6347 (N_6347,N_5652,N_5483);
nand U6348 (N_6348,N_5274,N_5691);
nor U6349 (N_6349,N_5719,N_5913);
or U6350 (N_6350,N_5468,N_5350);
or U6351 (N_6351,N_5687,N_5562);
and U6352 (N_6352,N_5647,N_5294);
nand U6353 (N_6353,N_5304,N_5531);
nand U6354 (N_6354,N_5845,N_5678);
nor U6355 (N_6355,N_5887,N_5299);
nand U6356 (N_6356,N_5646,N_5506);
or U6357 (N_6357,N_5577,N_5733);
or U6358 (N_6358,N_5631,N_5552);
xnor U6359 (N_6359,N_5340,N_5779);
or U6360 (N_6360,N_5810,N_5757);
and U6361 (N_6361,N_5749,N_5623);
nor U6362 (N_6362,N_5359,N_5305);
or U6363 (N_6363,N_5613,N_5611);
nand U6364 (N_6364,N_5499,N_5973);
and U6365 (N_6365,N_5576,N_5923);
or U6366 (N_6366,N_5514,N_5931);
or U6367 (N_6367,N_5437,N_5717);
or U6368 (N_6368,N_5419,N_5482);
and U6369 (N_6369,N_5557,N_5660);
xor U6370 (N_6370,N_5527,N_5336);
nor U6371 (N_6371,N_5925,N_5472);
nor U6372 (N_6372,N_5979,N_5921);
nand U6373 (N_6373,N_5378,N_5592);
and U6374 (N_6374,N_5798,N_5417);
nand U6375 (N_6375,N_5458,N_5967);
and U6376 (N_6376,N_5931,N_5957);
nand U6377 (N_6377,N_5817,N_5661);
or U6378 (N_6378,N_5268,N_5563);
and U6379 (N_6379,N_5633,N_5830);
or U6380 (N_6380,N_5854,N_5541);
nor U6381 (N_6381,N_5334,N_5405);
xor U6382 (N_6382,N_5277,N_5795);
nand U6383 (N_6383,N_5780,N_5250);
nand U6384 (N_6384,N_5348,N_5507);
or U6385 (N_6385,N_5659,N_5954);
and U6386 (N_6386,N_5545,N_5988);
or U6387 (N_6387,N_5763,N_5648);
nor U6388 (N_6388,N_5689,N_5465);
nor U6389 (N_6389,N_5591,N_5395);
and U6390 (N_6390,N_5305,N_5543);
and U6391 (N_6391,N_5325,N_5414);
nand U6392 (N_6392,N_5412,N_5385);
xnor U6393 (N_6393,N_5477,N_5690);
and U6394 (N_6394,N_5641,N_5936);
nor U6395 (N_6395,N_5531,N_5817);
nor U6396 (N_6396,N_5552,N_5712);
nand U6397 (N_6397,N_5673,N_5354);
and U6398 (N_6398,N_5889,N_5567);
or U6399 (N_6399,N_5848,N_5359);
nand U6400 (N_6400,N_5398,N_5556);
and U6401 (N_6401,N_5603,N_5260);
or U6402 (N_6402,N_5295,N_5363);
nor U6403 (N_6403,N_5689,N_5602);
or U6404 (N_6404,N_5755,N_5318);
nand U6405 (N_6405,N_5519,N_5794);
and U6406 (N_6406,N_5807,N_5504);
nand U6407 (N_6407,N_5696,N_5307);
or U6408 (N_6408,N_5394,N_5306);
nand U6409 (N_6409,N_5898,N_5803);
nor U6410 (N_6410,N_5785,N_5372);
nor U6411 (N_6411,N_5330,N_5853);
and U6412 (N_6412,N_5767,N_5667);
nor U6413 (N_6413,N_5594,N_5276);
nand U6414 (N_6414,N_5605,N_5351);
nand U6415 (N_6415,N_5417,N_5478);
nor U6416 (N_6416,N_5477,N_5280);
or U6417 (N_6417,N_5643,N_5976);
or U6418 (N_6418,N_5482,N_5714);
and U6419 (N_6419,N_5777,N_5810);
or U6420 (N_6420,N_5538,N_5568);
or U6421 (N_6421,N_5659,N_5866);
or U6422 (N_6422,N_5636,N_5460);
and U6423 (N_6423,N_5957,N_5568);
xor U6424 (N_6424,N_5642,N_5646);
nand U6425 (N_6425,N_5771,N_5814);
xnor U6426 (N_6426,N_5879,N_5302);
nand U6427 (N_6427,N_5534,N_5732);
or U6428 (N_6428,N_5585,N_5571);
nand U6429 (N_6429,N_5545,N_5466);
and U6430 (N_6430,N_5770,N_5882);
or U6431 (N_6431,N_5795,N_5709);
xor U6432 (N_6432,N_5417,N_5300);
xnor U6433 (N_6433,N_5618,N_5910);
and U6434 (N_6434,N_5559,N_5866);
or U6435 (N_6435,N_5807,N_5869);
and U6436 (N_6436,N_5722,N_5298);
or U6437 (N_6437,N_5932,N_5286);
or U6438 (N_6438,N_5326,N_5530);
nand U6439 (N_6439,N_5626,N_5840);
nor U6440 (N_6440,N_5353,N_5351);
and U6441 (N_6441,N_5358,N_5656);
and U6442 (N_6442,N_5574,N_5952);
or U6443 (N_6443,N_5645,N_5750);
xor U6444 (N_6444,N_5622,N_5870);
nor U6445 (N_6445,N_5743,N_5706);
or U6446 (N_6446,N_5839,N_5263);
nand U6447 (N_6447,N_5547,N_5290);
nor U6448 (N_6448,N_5589,N_5558);
nor U6449 (N_6449,N_5494,N_5355);
and U6450 (N_6450,N_5801,N_5502);
nand U6451 (N_6451,N_5266,N_5347);
or U6452 (N_6452,N_5825,N_5707);
or U6453 (N_6453,N_5864,N_5471);
nand U6454 (N_6454,N_5929,N_5822);
nand U6455 (N_6455,N_5350,N_5896);
and U6456 (N_6456,N_5534,N_5849);
xnor U6457 (N_6457,N_5576,N_5781);
or U6458 (N_6458,N_5923,N_5410);
nand U6459 (N_6459,N_5894,N_5416);
xnor U6460 (N_6460,N_5559,N_5869);
nor U6461 (N_6461,N_5446,N_5722);
nor U6462 (N_6462,N_5798,N_5928);
and U6463 (N_6463,N_5627,N_5918);
nand U6464 (N_6464,N_5972,N_5742);
and U6465 (N_6465,N_5977,N_5494);
and U6466 (N_6466,N_5664,N_5991);
and U6467 (N_6467,N_5846,N_5531);
nand U6468 (N_6468,N_5865,N_5785);
and U6469 (N_6469,N_5637,N_5354);
or U6470 (N_6470,N_5783,N_5522);
nor U6471 (N_6471,N_5842,N_5971);
nand U6472 (N_6472,N_5844,N_5565);
xnor U6473 (N_6473,N_5351,N_5330);
and U6474 (N_6474,N_5464,N_5469);
and U6475 (N_6475,N_5645,N_5651);
and U6476 (N_6476,N_5918,N_5559);
and U6477 (N_6477,N_5541,N_5495);
nand U6478 (N_6478,N_5809,N_5684);
nor U6479 (N_6479,N_5631,N_5466);
xnor U6480 (N_6480,N_5598,N_5564);
and U6481 (N_6481,N_5469,N_5346);
nor U6482 (N_6482,N_5600,N_5640);
xnor U6483 (N_6483,N_5665,N_5325);
nor U6484 (N_6484,N_5770,N_5273);
nand U6485 (N_6485,N_5364,N_5307);
nand U6486 (N_6486,N_5506,N_5625);
nand U6487 (N_6487,N_5944,N_5789);
xnor U6488 (N_6488,N_5589,N_5872);
or U6489 (N_6489,N_5285,N_5336);
and U6490 (N_6490,N_5949,N_5469);
nand U6491 (N_6491,N_5758,N_5303);
nor U6492 (N_6492,N_5330,N_5399);
nor U6493 (N_6493,N_5467,N_5439);
nor U6494 (N_6494,N_5351,N_5415);
xor U6495 (N_6495,N_5584,N_5712);
xnor U6496 (N_6496,N_5981,N_5713);
and U6497 (N_6497,N_5369,N_5587);
and U6498 (N_6498,N_5931,N_5741);
xor U6499 (N_6499,N_5945,N_5292);
nor U6500 (N_6500,N_5580,N_5519);
nand U6501 (N_6501,N_5264,N_5828);
xor U6502 (N_6502,N_5753,N_5520);
nor U6503 (N_6503,N_5677,N_5589);
and U6504 (N_6504,N_5336,N_5526);
xnor U6505 (N_6505,N_5869,N_5865);
or U6506 (N_6506,N_5312,N_5514);
nor U6507 (N_6507,N_5647,N_5714);
nor U6508 (N_6508,N_5506,N_5796);
or U6509 (N_6509,N_5896,N_5512);
nand U6510 (N_6510,N_5370,N_5696);
nand U6511 (N_6511,N_5623,N_5365);
nand U6512 (N_6512,N_5945,N_5866);
or U6513 (N_6513,N_5774,N_5390);
xnor U6514 (N_6514,N_5941,N_5392);
or U6515 (N_6515,N_5498,N_5265);
nand U6516 (N_6516,N_5935,N_5860);
and U6517 (N_6517,N_5574,N_5742);
and U6518 (N_6518,N_5630,N_5338);
or U6519 (N_6519,N_5827,N_5903);
nand U6520 (N_6520,N_5809,N_5552);
and U6521 (N_6521,N_5402,N_5323);
and U6522 (N_6522,N_5717,N_5967);
or U6523 (N_6523,N_5303,N_5787);
nor U6524 (N_6524,N_5556,N_5802);
or U6525 (N_6525,N_5427,N_5479);
or U6526 (N_6526,N_5720,N_5921);
nand U6527 (N_6527,N_5441,N_5512);
nand U6528 (N_6528,N_5851,N_5256);
or U6529 (N_6529,N_5773,N_5684);
xor U6530 (N_6530,N_5266,N_5615);
or U6531 (N_6531,N_5780,N_5770);
or U6532 (N_6532,N_5464,N_5721);
nor U6533 (N_6533,N_5802,N_5789);
nor U6534 (N_6534,N_5799,N_5464);
or U6535 (N_6535,N_5660,N_5936);
nand U6536 (N_6536,N_5952,N_5863);
nor U6537 (N_6537,N_5777,N_5573);
nand U6538 (N_6538,N_5680,N_5514);
or U6539 (N_6539,N_5317,N_5958);
nand U6540 (N_6540,N_5645,N_5956);
or U6541 (N_6541,N_5468,N_5914);
nor U6542 (N_6542,N_5752,N_5301);
xor U6543 (N_6543,N_5602,N_5257);
or U6544 (N_6544,N_5517,N_5687);
nor U6545 (N_6545,N_5348,N_5746);
nand U6546 (N_6546,N_5359,N_5871);
nand U6547 (N_6547,N_5972,N_5956);
nand U6548 (N_6548,N_5569,N_5355);
nor U6549 (N_6549,N_5841,N_5321);
xor U6550 (N_6550,N_5320,N_5995);
or U6551 (N_6551,N_5927,N_5708);
nor U6552 (N_6552,N_5478,N_5524);
or U6553 (N_6553,N_5358,N_5907);
and U6554 (N_6554,N_5452,N_5940);
and U6555 (N_6555,N_5992,N_5820);
nor U6556 (N_6556,N_5383,N_5513);
or U6557 (N_6557,N_5812,N_5258);
or U6558 (N_6558,N_5974,N_5711);
or U6559 (N_6559,N_5391,N_5702);
or U6560 (N_6560,N_5305,N_5879);
nor U6561 (N_6561,N_5401,N_5724);
and U6562 (N_6562,N_5255,N_5454);
and U6563 (N_6563,N_5403,N_5764);
and U6564 (N_6564,N_5401,N_5997);
and U6565 (N_6565,N_5765,N_5401);
or U6566 (N_6566,N_5374,N_5705);
or U6567 (N_6567,N_5479,N_5463);
and U6568 (N_6568,N_5895,N_5941);
and U6569 (N_6569,N_5682,N_5286);
or U6570 (N_6570,N_5665,N_5904);
nor U6571 (N_6571,N_5791,N_5423);
and U6572 (N_6572,N_5706,N_5474);
xor U6573 (N_6573,N_5673,N_5280);
nor U6574 (N_6574,N_5985,N_5808);
or U6575 (N_6575,N_5266,N_5441);
and U6576 (N_6576,N_5692,N_5964);
nand U6577 (N_6577,N_5480,N_5821);
xor U6578 (N_6578,N_5612,N_5632);
nor U6579 (N_6579,N_5503,N_5548);
and U6580 (N_6580,N_5700,N_5855);
nor U6581 (N_6581,N_5857,N_5649);
nor U6582 (N_6582,N_5665,N_5725);
nor U6583 (N_6583,N_5949,N_5889);
or U6584 (N_6584,N_5285,N_5409);
or U6585 (N_6585,N_5565,N_5649);
or U6586 (N_6586,N_5319,N_5813);
nand U6587 (N_6587,N_5557,N_5642);
nor U6588 (N_6588,N_5646,N_5573);
and U6589 (N_6589,N_5472,N_5567);
and U6590 (N_6590,N_5348,N_5614);
nand U6591 (N_6591,N_5904,N_5250);
nand U6592 (N_6592,N_5270,N_5998);
and U6593 (N_6593,N_5688,N_5315);
nand U6594 (N_6594,N_5547,N_5505);
nor U6595 (N_6595,N_5360,N_5645);
nor U6596 (N_6596,N_5415,N_5993);
and U6597 (N_6597,N_5490,N_5851);
xor U6598 (N_6598,N_5632,N_5680);
nand U6599 (N_6599,N_5764,N_5484);
and U6600 (N_6600,N_5745,N_5942);
nor U6601 (N_6601,N_5729,N_5553);
or U6602 (N_6602,N_5526,N_5351);
nor U6603 (N_6603,N_5619,N_5379);
or U6604 (N_6604,N_5378,N_5931);
or U6605 (N_6605,N_5253,N_5924);
and U6606 (N_6606,N_5515,N_5542);
or U6607 (N_6607,N_5357,N_5990);
and U6608 (N_6608,N_5921,N_5936);
xnor U6609 (N_6609,N_5635,N_5836);
nor U6610 (N_6610,N_5505,N_5788);
xor U6611 (N_6611,N_5835,N_5444);
and U6612 (N_6612,N_5374,N_5869);
and U6613 (N_6613,N_5948,N_5801);
or U6614 (N_6614,N_5525,N_5583);
nor U6615 (N_6615,N_5299,N_5839);
nor U6616 (N_6616,N_5875,N_5893);
and U6617 (N_6617,N_5797,N_5505);
and U6618 (N_6618,N_5858,N_5364);
nand U6619 (N_6619,N_5489,N_5300);
nor U6620 (N_6620,N_5591,N_5528);
nand U6621 (N_6621,N_5588,N_5490);
and U6622 (N_6622,N_5908,N_5698);
or U6623 (N_6623,N_5587,N_5334);
or U6624 (N_6624,N_5322,N_5382);
and U6625 (N_6625,N_5554,N_5405);
and U6626 (N_6626,N_5823,N_5919);
nor U6627 (N_6627,N_5391,N_5736);
nor U6628 (N_6628,N_5575,N_5412);
nand U6629 (N_6629,N_5366,N_5556);
nand U6630 (N_6630,N_5306,N_5528);
or U6631 (N_6631,N_5743,N_5718);
nor U6632 (N_6632,N_5848,N_5865);
nand U6633 (N_6633,N_5716,N_5643);
nor U6634 (N_6634,N_5513,N_5527);
nand U6635 (N_6635,N_5827,N_5379);
and U6636 (N_6636,N_5296,N_5316);
nor U6637 (N_6637,N_5324,N_5818);
or U6638 (N_6638,N_5558,N_5936);
nor U6639 (N_6639,N_5956,N_5948);
nand U6640 (N_6640,N_5842,N_5913);
nor U6641 (N_6641,N_5508,N_5708);
nor U6642 (N_6642,N_5407,N_5466);
or U6643 (N_6643,N_5915,N_5448);
nand U6644 (N_6644,N_5728,N_5650);
and U6645 (N_6645,N_5412,N_5450);
nand U6646 (N_6646,N_5667,N_5406);
nand U6647 (N_6647,N_5307,N_5368);
nand U6648 (N_6648,N_5674,N_5366);
nand U6649 (N_6649,N_5644,N_5603);
and U6650 (N_6650,N_5556,N_5492);
and U6651 (N_6651,N_5843,N_5667);
xor U6652 (N_6652,N_5576,N_5568);
or U6653 (N_6653,N_5649,N_5577);
nor U6654 (N_6654,N_5530,N_5323);
nand U6655 (N_6655,N_5407,N_5985);
nand U6656 (N_6656,N_5553,N_5450);
and U6657 (N_6657,N_5490,N_5597);
nor U6658 (N_6658,N_5973,N_5959);
and U6659 (N_6659,N_5886,N_5603);
nand U6660 (N_6660,N_5675,N_5798);
nand U6661 (N_6661,N_5616,N_5585);
nand U6662 (N_6662,N_5780,N_5898);
and U6663 (N_6663,N_5614,N_5907);
and U6664 (N_6664,N_5360,N_5577);
nand U6665 (N_6665,N_5705,N_5775);
nand U6666 (N_6666,N_5741,N_5397);
nor U6667 (N_6667,N_5578,N_5545);
nor U6668 (N_6668,N_5507,N_5995);
or U6669 (N_6669,N_5974,N_5840);
nand U6670 (N_6670,N_5871,N_5936);
nor U6671 (N_6671,N_5590,N_5989);
nand U6672 (N_6672,N_5409,N_5624);
and U6673 (N_6673,N_5516,N_5871);
nand U6674 (N_6674,N_5623,N_5431);
nand U6675 (N_6675,N_5319,N_5893);
nand U6676 (N_6676,N_5772,N_5285);
xor U6677 (N_6677,N_5930,N_5628);
and U6678 (N_6678,N_5312,N_5391);
nand U6679 (N_6679,N_5987,N_5908);
or U6680 (N_6680,N_5366,N_5494);
nor U6681 (N_6681,N_5576,N_5371);
or U6682 (N_6682,N_5522,N_5942);
and U6683 (N_6683,N_5486,N_5737);
nor U6684 (N_6684,N_5937,N_5553);
and U6685 (N_6685,N_5936,N_5886);
nor U6686 (N_6686,N_5855,N_5493);
and U6687 (N_6687,N_5626,N_5851);
nor U6688 (N_6688,N_5873,N_5521);
xnor U6689 (N_6689,N_5319,N_5773);
and U6690 (N_6690,N_5399,N_5496);
nor U6691 (N_6691,N_5504,N_5483);
nand U6692 (N_6692,N_5510,N_5322);
or U6693 (N_6693,N_5879,N_5269);
xor U6694 (N_6694,N_5450,N_5764);
and U6695 (N_6695,N_5497,N_5362);
nand U6696 (N_6696,N_5714,N_5422);
nand U6697 (N_6697,N_5383,N_5542);
or U6698 (N_6698,N_5721,N_5737);
and U6699 (N_6699,N_5594,N_5602);
nor U6700 (N_6700,N_5990,N_5793);
or U6701 (N_6701,N_5433,N_5908);
or U6702 (N_6702,N_5955,N_5631);
and U6703 (N_6703,N_5644,N_5496);
nor U6704 (N_6704,N_5372,N_5700);
xor U6705 (N_6705,N_5917,N_5685);
nor U6706 (N_6706,N_5812,N_5351);
xnor U6707 (N_6707,N_5636,N_5572);
xnor U6708 (N_6708,N_5519,N_5915);
or U6709 (N_6709,N_5758,N_5285);
and U6710 (N_6710,N_5673,N_5584);
and U6711 (N_6711,N_5480,N_5356);
xnor U6712 (N_6712,N_5434,N_5737);
nand U6713 (N_6713,N_5998,N_5283);
and U6714 (N_6714,N_5538,N_5758);
and U6715 (N_6715,N_5957,N_5614);
nor U6716 (N_6716,N_5806,N_5305);
or U6717 (N_6717,N_5610,N_5973);
nor U6718 (N_6718,N_5666,N_5268);
nand U6719 (N_6719,N_5577,N_5387);
or U6720 (N_6720,N_5437,N_5408);
nor U6721 (N_6721,N_5885,N_5311);
or U6722 (N_6722,N_5418,N_5586);
nand U6723 (N_6723,N_5504,N_5610);
and U6724 (N_6724,N_5521,N_5573);
nand U6725 (N_6725,N_5854,N_5891);
nand U6726 (N_6726,N_5709,N_5431);
nor U6727 (N_6727,N_5752,N_5272);
and U6728 (N_6728,N_5570,N_5915);
nor U6729 (N_6729,N_5582,N_5783);
and U6730 (N_6730,N_5282,N_5519);
xnor U6731 (N_6731,N_5811,N_5725);
nor U6732 (N_6732,N_5941,N_5372);
nand U6733 (N_6733,N_5268,N_5691);
nand U6734 (N_6734,N_5925,N_5596);
nor U6735 (N_6735,N_5822,N_5857);
nand U6736 (N_6736,N_5813,N_5656);
nor U6737 (N_6737,N_5817,N_5476);
nor U6738 (N_6738,N_5786,N_5611);
xor U6739 (N_6739,N_5487,N_5564);
nor U6740 (N_6740,N_5953,N_5744);
nand U6741 (N_6741,N_5572,N_5288);
xnor U6742 (N_6742,N_5618,N_5937);
and U6743 (N_6743,N_5764,N_5552);
xor U6744 (N_6744,N_5753,N_5346);
and U6745 (N_6745,N_5934,N_5913);
or U6746 (N_6746,N_5470,N_5889);
or U6747 (N_6747,N_5310,N_5761);
nor U6748 (N_6748,N_5665,N_5559);
nand U6749 (N_6749,N_5580,N_5455);
xnor U6750 (N_6750,N_6027,N_6021);
nand U6751 (N_6751,N_6487,N_6393);
or U6752 (N_6752,N_6336,N_6341);
and U6753 (N_6753,N_6479,N_6056);
nor U6754 (N_6754,N_6383,N_6627);
nand U6755 (N_6755,N_6338,N_6477);
nor U6756 (N_6756,N_6260,N_6322);
nand U6757 (N_6757,N_6580,N_6267);
nand U6758 (N_6758,N_6448,N_6149);
and U6759 (N_6759,N_6051,N_6522);
nor U6760 (N_6760,N_6211,N_6196);
xnor U6761 (N_6761,N_6095,N_6151);
or U6762 (N_6762,N_6456,N_6680);
nor U6763 (N_6763,N_6671,N_6586);
nand U6764 (N_6764,N_6483,N_6572);
nor U6765 (N_6765,N_6063,N_6692);
or U6766 (N_6766,N_6610,N_6518);
nor U6767 (N_6767,N_6141,N_6742);
or U6768 (N_6768,N_6176,N_6353);
nor U6769 (N_6769,N_6651,N_6200);
nand U6770 (N_6770,N_6375,N_6085);
nor U6771 (N_6771,N_6437,N_6689);
xnor U6772 (N_6772,N_6055,N_6065);
nand U6773 (N_6773,N_6058,N_6728);
or U6774 (N_6774,N_6428,N_6460);
and U6775 (N_6775,N_6665,N_6054);
nand U6776 (N_6776,N_6257,N_6191);
nand U6777 (N_6777,N_6486,N_6617);
xor U6778 (N_6778,N_6420,N_6184);
nor U6779 (N_6779,N_6583,N_6004);
and U6780 (N_6780,N_6395,N_6381);
nand U6781 (N_6781,N_6639,N_6521);
nor U6782 (N_6782,N_6227,N_6536);
and U6783 (N_6783,N_6668,N_6088);
xor U6784 (N_6784,N_6497,N_6575);
nand U6785 (N_6785,N_6546,N_6560);
nor U6786 (N_6786,N_6309,N_6556);
and U6787 (N_6787,N_6139,N_6441);
nand U6788 (N_6788,N_6210,N_6593);
or U6789 (N_6789,N_6140,N_6117);
nand U6790 (N_6790,N_6515,N_6024);
or U6791 (N_6791,N_6566,N_6189);
and U6792 (N_6792,N_6623,N_6120);
or U6793 (N_6793,N_6740,N_6493);
or U6794 (N_6794,N_6506,N_6710);
nand U6795 (N_6795,N_6520,N_6073);
nand U6796 (N_6796,N_6371,N_6505);
nand U6797 (N_6797,N_6242,N_6530);
xor U6798 (N_6798,N_6685,N_6635);
xnor U6799 (N_6799,N_6485,N_6165);
nand U6800 (N_6800,N_6561,N_6291);
nor U6801 (N_6801,N_6693,N_6588);
nor U6802 (N_6802,N_6606,N_6204);
nand U6803 (N_6803,N_6609,N_6256);
and U6804 (N_6804,N_6344,N_6469);
xnor U6805 (N_6805,N_6499,N_6271);
nor U6806 (N_6806,N_6724,N_6173);
nor U6807 (N_6807,N_6661,N_6299);
nand U6808 (N_6808,N_6451,N_6620);
or U6809 (N_6809,N_6453,N_6495);
nor U6810 (N_6810,N_6619,N_6007);
nor U6811 (N_6811,N_6444,N_6434);
or U6812 (N_6812,N_6013,N_6711);
and U6813 (N_6813,N_6356,N_6360);
nand U6814 (N_6814,N_6432,N_6488);
and U6815 (N_6815,N_6399,N_6239);
nand U6816 (N_6816,N_6226,N_6504);
or U6817 (N_6817,N_6333,N_6192);
and U6818 (N_6818,N_6640,N_6482);
and U6819 (N_6819,N_6747,N_6722);
nor U6820 (N_6820,N_6585,N_6134);
nand U6821 (N_6821,N_6052,N_6332);
and U6822 (N_6822,N_6070,N_6468);
nor U6823 (N_6823,N_6405,N_6167);
or U6824 (N_6824,N_6032,N_6626);
nand U6825 (N_6825,N_6442,N_6708);
and U6826 (N_6826,N_6409,N_6272);
and U6827 (N_6827,N_6224,N_6491);
nand U6828 (N_6828,N_6553,N_6337);
nor U6829 (N_6829,N_6726,N_6234);
xnor U6830 (N_6830,N_6287,N_6547);
nand U6831 (N_6831,N_6177,N_6500);
nor U6832 (N_6832,N_6737,N_6303);
xor U6833 (N_6833,N_6529,N_6046);
nor U6834 (N_6834,N_6218,N_6490);
nand U6835 (N_6835,N_6702,N_6524);
nor U6836 (N_6836,N_6069,N_6306);
nand U6837 (N_6837,N_6124,N_6372);
xor U6838 (N_6838,N_6086,N_6221);
nand U6839 (N_6839,N_6037,N_6119);
nand U6840 (N_6840,N_6125,N_6001);
nand U6841 (N_6841,N_6723,N_6185);
nor U6842 (N_6842,N_6384,N_6464);
nor U6843 (N_6843,N_6067,N_6156);
or U6844 (N_6844,N_6532,N_6305);
nor U6845 (N_6845,N_6564,N_6555);
or U6846 (N_6846,N_6285,N_6633);
and U6847 (N_6847,N_6253,N_6042);
nand U6848 (N_6848,N_6031,N_6410);
and U6849 (N_6849,N_6050,N_6208);
nand U6850 (N_6850,N_6696,N_6084);
or U6851 (N_6851,N_6354,N_6157);
and U6852 (N_6852,N_6077,N_6195);
nor U6853 (N_6853,N_6574,N_6687);
or U6854 (N_6854,N_6649,N_6352);
and U6855 (N_6855,N_6376,N_6161);
or U6856 (N_6856,N_6718,N_6461);
nor U6857 (N_6857,N_6110,N_6734);
nor U6858 (N_6858,N_6011,N_6265);
nor U6859 (N_6859,N_6153,N_6122);
or U6860 (N_6860,N_6411,N_6143);
or U6861 (N_6861,N_6092,N_6648);
nor U6862 (N_6862,N_6214,N_6193);
nor U6863 (N_6863,N_6362,N_6220);
nor U6864 (N_6864,N_6040,N_6736);
nand U6865 (N_6865,N_6596,N_6449);
nand U6866 (N_6866,N_6531,N_6599);
nor U6867 (N_6867,N_6284,N_6160);
and U6868 (N_6868,N_6652,N_6066);
or U6869 (N_6869,N_6094,N_6729);
nand U6870 (N_6870,N_6237,N_6537);
and U6871 (N_6871,N_6557,N_6594);
nor U6872 (N_6872,N_6618,N_6359);
and U6873 (N_6873,N_6080,N_6559);
or U6874 (N_6874,N_6509,N_6251);
or U6875 (N_6875,N_6012,N_6244);
and U6876 (N_6876,N_6701,N_6235);
nand U6877 (N_6877,N_6527,N_6664);
nand U6878 (N_6878,N_6517,N_6567);
nand U6879 (N_6879,N_6670,N_6343);
xnor U6880 (N_6880,N_6158,N_6201);
xor U6881 (N_6881,N_6026,N_6424);
and U6882 (N_6882,N_6462,N_6544);
or U6883 (N_6883,N_6282,N_6731);
or U6884 (N_6884,N_6390,N_6168);
and U6885 (N_6885,N_6133,N_6030);
or U6886 (N_6886,N_6459,N_6474);
or U6887 (N_6887,N_6103,N_6408);
and U6888 (N_6888,N_6415,N_6355);
nand U6889 (N_6889,N_6187,N_6015);
or U6890 (N_6890,N_6455,N_6171);
nor U6891 (N_6891,N_6089,N_6276);
nand U6892 (N_6892,N_6129,N_6053);
or U6893 (N_6893,N_6288,N_6036);
or U6894 (N_6894,N_6370,N_6502);
xor U6895 (N_6895,N_6523,N_6005);
or U6896 (N_6896,N_6528,N_6006);
xor U6897 (N_6897,N_6412,N_6166);
nand U6898 (N_6898,N_6400,N_6000);
nand U6899 (N_6899,N_6373,N_6578);
nand U6900 (N_6900,N_6535,N_6590);
and U6901 (N_6901,N_6514,N_6570);
nand U6902 (N_6902,N_6202,N_6131);
nor U6903 (N_6903,N_6057,N_6020);
and U6904 (N_6904,N_6397,N_6741);
or U6905 (N_6905,N_6159,N_6587);
and U6906 (N_6906,N_6655,N_6246);
or U6907 (N_6907,N_6183,N_6698);
nor U6908 (N_6908,N_6198,N_6392);
and U6909 (N_6909,N_6660,N_6611);
and U6910 (N_6910,N_6466,N_6388);
nand U6911 (N_6911,N_6215,N_6096);
or U6912 (N_6912,N_6114,N_6327);
nand U6913 (N_6913,N_6571,N_6098);
xor U6914 (N_6914,N_6435,N_6358);
nor U6915 (N_6915,N_6175,N_6385);
nor U6916 (N_6916,N_6207,N_6732);
nand U6917 (N_6917,N_6047,N_6289);
nand U6918 (N_6918,N_6746,N_6154);
nor U6919 (N_6919,N_6598,N_6720);
nand U6920 (N_6920,N_6714,N_6382);
xnor U6921 (N_6921,N_6060,N_6407);
or U6922 (N_6922,N_6642,N_6577);
and U6923 (N_6923,N_6262,N_6298);
nand U6924 (N_6924,N_6439,N_6179);
nor U6925 (N_6925,N_6657,N_6249);
nand U6926 (N_6926,N_6081,N_6155);
and U6927 (N_6927,N_6074,N_6645);
nor U6928 (N_6928,N_6454,N_6164);
xor U6929 (N_6929,N_6690,N_6422);
or U6930 (N_6930,N_6601,N_6169);
nand U6931 (N_6931,N_6540,N_6107);
nand U6932 (N_6932,N_6636,N_6398);
or U6933 (N_6933,N_6238,N_6433);
or U6934 (N_6934,N_6367,N_6533);
and U6935 (N_6935,N_6266,N_6130);
nor U6936 (N_6936,N_6735,N_6072);
nand U6937 (N_6937,N_6232,N_6342);
nand U6938 (N_6938,N_6075,N_6511);
or U6939 (N_6939,N_6104,N_6194);
xor U6940 (N_6940,N_6458,N_6628);
and U6941 (N_6941,N_6616,N_6034);
xnor U6942 (N_6942,N_6697,N_6132);
nor U6943 (N_6943,N_6548,N_6621);
and U6944 (N_6944,N_6709,N_6319);
nand U6945 (N_6945,N_6470,N_6414);
nand U6946 (N_6946,N_6581,N_6366);
nand U6947 (N_6947,N_6744,N_6025);
or U6948 (N_6948,N_6135,N_6002);
and U6949 (N_6949,N_6480,N_6062);
xnor U6950 (N_6950,N_6526,N_6035);
nand U6951 (N_6951,N_6427,N_6233);
nor U6952 (N_6952,N_6301,N_6592);
nand U6953 (N_6953,N_6673,N_6349);
or U6954 (N_6954,N_6730,N_6281);
nand U6955 (N_6955,N_6009,N_6662);
or U6956 (N_6956,N_6268,N_6090);
or U6957 (N_6957,N_6430,N_6315);
or U6958 (N_6958,N_6087,N_6279);
nor U6959 (N_6959,N_6261,N_6223);
nor U6960 (N_6960,N_6330,N_6018);
and U6961 (N_6961,N_6017,N_6263);
and U6962 (N_6962,N_6543,N_6181);
or U6963 (N_6963,N_6541,N_6346);
or U6964 (N_6964,N_6116,N_6209);
or U6965 (N_6965,N_6603,N_6216);
nor U6966 (N_6966,N_6615,N_6391);
nor U6967 (N_6967,N_6269,N_6387);
or U6968 (N_6968,N_6290,N_6446);
nand U6969 (N_6969,N_6247,N_6463);
and U6970 (N_6970,N_6695,N_6182);
and U6971 (N_6971,N_6705,N_6274);
or U6972 (N_6972,N_6421,N_6688);
or U6973 (N_6973,N_6038,N_6647);
and U6974 (N_6974,N_6538,N_6563);
or U6975 (N_6975,N_6363,N_6713);
or U6976 (N_6976,N_6508,N_6721);
nor U6977 (N_6977,N_6542,N_6286);
or U6978 (N_6978,N_6749,N_6314);
nor U6979 (N_6979,N_6602,N_6101);
nand U6980 (N_6980,N_6145,N_6347);
and U6981 (N_6981,N_6163,N_6059);
nand U6982 (N_6982,N_6243,N_6457);
and U6983 (N_6983,N_6076,N_6582);
and U6984 (N_6984,N_6039,N_6108);
nor U6985 (N_6985,N_6369,N_6507);
or U6986 (N_6986,N_6328,N_6492);
nand U6987 (N_6987,N_6219,N_6188);
and U6988 (N_6988,N_6643,N_6137);
nor U6989 (N_6989,N_6308,N_6252);
and U6990 (N_6990,N_6199,N_6473);
and U6991 (N_6991,N_6684,N_6484);
nand U6992 (N_6992,N_6402,N_6321);
or U6993 (N_6993,N_6307,N_6097);
nor U6994 (N_6994,N_6348,N_6245);
xor U6995 (N_6995,N_6694,N_6404);
or U6996 (N_6996,N_6739,N_6230);
or U6997 (N_6997,N_6595,N_6691);
and U6998 (N_6998,N_6498,N_6496);
nor U6999 (N_6999,N_6699,N_6440);
or U7000 (N_7000,N_6646,N_6203);
nand U7001 (N_7001,N_6357,N_6503);
and U7002 (N_7002,N_6679,N_6106);
xor U7003 (N_7003,N_6597,N_6250);
nor U7004 (N_7004,N_6677,N_6608);
nor U7005 (N_7005,N_6361,N_6656);
and U7006 (N_7006,N_6475,N_6351);
nand U7007 (N_7007,N_6653,N_6222);
nand U7008 (N_7008,N_6102,N_6300);
or U7009 (N_7009,N_6629,N_6339);
or U7010 (N_7010,N_6406,N_6278);
nor U7011 (N_7011,N_6008,N_6374);
nor U7012 (N_7012,N_6045,N_6706);
and U7013 (N_7013,N_6078,N_6667);
nor U7014 (N_7014,N_6379,N_6465);
or U7015 (N_7015,N_6568,N_6326);
and U7016 (N_7016,N_6686,N_6150);
or U7017 (N_7017,N_6419,N_6248);
and U7018 (N_7018,N_6550,N_6666);
and U7019 (N_7019,N_6186,N_6178);
xor U7020 (N_7020,N_6403,N_6501);
or U7021 (N_7021,N_6313,N_6334);
nand U7022 (N_7022,N_6048,N_6682);
nor U7023 (N_7023,N_6311,N_6478);
or U7024 (N_7024,N_6297,N_6654);
nor U7025 (N_7025,N_6283,N_6683);
nand U7026 (N_7026,N_6436,N_6712);
xor U7027 (N_7027,N_6331,N_6674);
or U7028 (N_7028,N_6118,N_6579);
or U7029 (N_7029,N_6638,N_6516);
and U7030 (N_7030,N_6109,N_6041);
xnor U7031 (N_7031,N_6650,N_6049);
and U7032 (N_7032,N_6105,N_6584);
xnor U7033 (N_7033,N_6082,N_6205);
and U7034 (N_7034,N_6071,N_6275);
xor U7035 (N_7035,N_6152,N_6064);
nand U7036 (N_7036,N_6386,N_6236);
nand U7037 (N_7037,N_6589,N_6637);
nor U7038 (N_7038,N_6554,N_6148);
nor U7039 (N_7039,N_6231,N_6228);
nand U7040 (N_7040,N_6591,N_6417);
nor U7041 (N_7041,N_6043,N_6147);
and U7042 (N_7042,N_6316,N_6573);
and U7043 (N_7043,N_6641,N_6113);
nand U7044 (N_7044,N_6121,N_6445);
nor U7045 (N_7045,N_6719,N_6631);
and U7046 (N_7046,N_6743,N_6622);
nand U7047 (N_7047,N_6425,N_6280);
nand U7048 (N_7048,N_6489,N_6068);
nor U7049 (N_7049,N_6481,N_6144);
nor U7050 (N_7050,N_6014,N_6292);
or U7051 (N_7051,N_6029,N_6431);
or U7052 (N_7052,N_6476,N_6197);
and U7053 (N_7053,N_6707,N_6254);
or U7054 (N_7054,N_6377,N_6552);
and U7055 (N_7055,N_6146,N_6551);
nor U7056 (N_7056,N_6678,N_6350);
and U7057 (N_7057,N_6378,N_6562);
or U7058 (N_7058,N_6019,N_6644);
nor U7059 (N_7059,N_6630,N_6558);
nand U7060 (N_7060,N_6325,N_6212);
nor U7061 (N_7061,N_6138,N_6128);
or U7062 (N_7062,N_6452,N_6624);
nand U7063 (N_7063,N_6123,N_6625);
nor U7064 (N_7064,N_6335,N_6126);
nand U7065 (N_7065,N_6539,N_6127);
nor U7066 (N_7066,N_6733,N_6295);
or U7067 (N_7067,N_6513,N_6494);
nor U7068 (N_7068,N_6748,N_6525);
or U7069 (N_7069,N_6091,N_6099);
nand U7070 (N_7070,N_6264,N_6061);
nor U7071 (N_7071,N_6368,N_6217);
and U7072 (N_7072,N_6044,N_6079);
or U7073 (N_7073,N_6083,N_6438);
nor U7074 (N_7074,N_6607,N_6302);
nor U7075 (N_7075,N_6028,N_6738);
and U7076 (N_7076,N_6716,N_6093);
or U7077 (N_7077,N_6293,N_6304);
and U7078 (N_7078,N_6180,N_6258);
xor U7079 (N_7079,N_6190,N_6510);
nand U7080 (N_7080,N_6663,N_6213);
nand U7081 (N_7081,N_6672,N_6416);
nor U7082 (N_7082,N_6429,N_6172);
xnor U7083 (N_7083,N_6472,N_6345);
nor U7084 (N_7084,N_6659,N_6605);
nor U7085 (N_7085,N_6115,N_6565);
nor U7086 (N_7086,N_6604,N_6447);
and U7087 (N_7087,N_6174,N_6614);
nand U7088 (N_7088,N_6329,N_6727);
and U7089 (N_7089,N_6471,N_6100);
and U7090 (N_7090,N_6022,N_6206);
nor U7091 (N_7091,N_6112,N_6576);
or U7092 (N_7092,N_6389,N_6273);
nor U7093 (N_7093,N_6162,N_6136);
nand U7094 (N_7094,N_6111,N_6401);
nand U7095 (N_7095,N_6229,N_6675);
nand U7096 (N_7096,N_6003,N_6600);
and U7097 (N_7097,N_6010,N_6569);
nand U7098 (N_7098,N_6658,N_6240);
nand U7099 (N_7099,N_6725,N_6365);
and U7100 (N_7100,N_6676,N_6340);
xnor U7101 (N_7101,N_6320,N_6413);
or U7102 (N_7102,N_6745,N_6467);
and U7103 (N_7103,N_6418,N_6443);
nand U7104 (N_7104,N_6312,N_6634);
nor U7105 (N_7105,N_6277,N_6512);
or U7106 (N_7106,N_6270,N_6318);
xnor U7107 (N_7107,N_6225,N_6704);
nand U7108 (N_7108,N_6426,N_6142);
or U7109 (N_7109,N_6612,N_6681);
nor U7110 (N_7110,N_6396,N_6310);
and U7111 (N_7111,N_6296,N_6259);
or U7112 (N_7112,N_6016,N_6394);
nor U7113 (N_7113,N_6380,N_6323);
nand U7114 (N_7114,N_6033,N_6023);
nand U7115 (N_7115,N_6423,N_6255);
nand U7116 (N_7116,N_6450,N_6170);
nand U7117 (N_7117,N_6717,N_6534);
and U7118 (N_7118,N_6324,N_6632);
or U7119 (N_7119,N_6669,N_6317);
or U7120 (N_7120,N_6703,N_6545);
nand U7121 (N_7121,N_6241,N_6519);
or U7122 (N_7122,N_6364,N_6715);
nor U7123 (N_7123,N_6549,N_6613);
or U7124 (N_7124,N_6294,N_6700);
nor U7125 (N_7125,N_6079,N_6632);
and U7126 (N_7126,N_6362,N_6042);
and U7127 (N_7127,N_6603,N_6234);
nor U7128 (N_7128,N_6377,N_6466);
or U7129 (N_7129,N_6203,N_6555);
xnor U7130 (N_7130,N_6498,N_6078);
nor U7131 (N_7131,N_6584,N_6443);
or U7132 (N_7132,N_6627,N_6683);
nor U7133 (N_7133,N_6474,N_6041);
nor U7134 (N_7134,N_6283,N_6559);
nor U7135 (N_7135,N_6382,N_6727);
and U7136 (N_7136,N_6283,N_6189);
nand U7137 (N_7137,N_6194,N_6637);
xnor U7138 (N_7138,N_6047,N_6642);
nor U7139 (N_7139,N_6071,N_6472);
nand U7140 (N_7140,N_6639,N_6539);
and U7141 (N_7141,N_6665,N_6243);
xor U7142 (N_7142,N_6536,N_6725);
nor U7143 (N_7143,N_6685,N_6052);
nand U7144 (N_7144,N_6683,N_6260);
nand U7145 (N_7145,N_6596,N_6469);
or U7146 (N_7146,N_6424,N_6745);
or U7147 (N_7147,N_6694,N_6228);
and U7148 (N_7148,N_6073,N_6494);
xnor U7149 (N_7149,N_6208,N_6488);
nand U7150 (N_7150,N_6607,N_6203);
or U7151 (N_7151,N_6537,N_6152);
xor U7152 (N_7152,N_6522,N_6491);
nand U7153 (N_7153,N_6243,N_6480);
or U7154 (N_7154,N_6499,N_6265);
nor U7155 (N_7155,N_6283,N_6514);
nor U7156 (N_7156,N_6241,N_6279);
and U7157 (N_7157,N_6462,N_6111);
or U7158 (N_7158,N_6531,N_6196);
and U7159 (N_7159,N_6720,N_6160);
and U7160 (N_7160,N_6461,N_6689);
and U7161 (N_7161,N_6624,N_6611);
or U7162 (N_7162,N_6414,N_6110);
nor U7163 (N_7163,N_6657,N_6181);
and U7164 (N_7164,N_6289,N_6190);
nor U7165 (N_7165,N_6207,N_6199);
or U7166 (N_7166,N_6024,N_6025);
and U7167 (N_7167,N_6486,N_6113);
or U7168 (N_7168,N_6006,N_6660);
and U7169 (N_7169,N_6695,N_6398);
nor U7170 (N_7170,N_6310,N_6219);
or U7171 (N_7171,N_6376,N_6196);
nor U7172 (N_7172,N_6508,N_6069);
nand U7173 (N_7173,N_6426,N_6032);
nor U7174 (N_7174,N_6209,N_6196);
xnor U7175 (N_7175,N_6517,N_6179);
or U7176 (N_7176,N_6272,N_6225);
and U7177 (N_7177,N_6322,N_6347);
or U7178 (N_7178,N_6039,N_6486);
and U7179 (N_7179,N_6339,N_6294);
nand U7180 (N_7180,N_6664,N_6490);
nand U7181 (N_7181,N_6609,N_6511);
and U7182 (N_7182,N_6597,N_6163);
and U7183 (N_7183,N_6365,N_6630);
nor U7184 (N_7184,N_6266,N_6334);
or U7185 (N_7185,N_6094,N_6714);
and U7186 (N_7186,N_6286,N_6655);
or U7187 (N_7187,N_6300,N_6532);
nand U7188 (N_7188,N_6328,N_6568);
and U7189 (N_7189,N_6687,N_6106);
nand U7190 (N_7190,N_6493,N_6037);
nand U7191 (N_7191,N_6170,N_6119);
xor U7192 (N_7192,N_6329,N_6182);
xor U7193 (N_7193,N_6269,N_6079);
and U7194 (N_7194,N_6516,N_6630);
nand U7195 (N_7195,N_6466,N_6187);
and U7196 (N_7196,N_6273,N_6523);
or U7197 (N_7197,N_6405,N_6425);
and U7198 (N_7198,N_6714,N_6725);
or U7199 (N_7199,N_6191,N_6381);
nor U7200 (N_7200,N_6073,N_6380);
or U7201 (N_7201,N_6634,N_6255);
or U7202 (N_7202,N_6031,N_6665);
nor U7203 (N_7203,N_6275,N_6509);
xor U7204 (N_7204,N_6616,N_6107);
or U7205 (N_7205,N_6582,N_6740);
nor U7206 (N_7206,N_6543,N_6703);
or U7207 (N_7207,N_6237,N_6456);
nor U7208 (N_7208,N_6640,N_6415);
or U7209 (N_7209,N_6507,N_6326);
nand U7210 (N_7210,N_6115,N_6177);
nand U7211 (N_7211,N_6440,N_6435);
or U7212 (N_7212,N_6494,N_6375);
and U7213 (N_7213,N_6294,N_6477);
and U7214 (N_7214,N_6355,N_6523);
nor U7215 (N_7215,N_6308,N_6344);
or U7216 (N_7216,N_6513,N_6239);
nor U7217 (N_7217,N_6200,N_6555);
and U7218 (N_7218,N_6127,N_6636);
xnor U7219 (N_7219,N_6158,N_6184);
nor U7220 (N_7220,N_6300,N_6667);
nor U7221 (N_7221,N_6483,N_6671);
nand U7222 (N_7222,N_6492,N_6442);
or U7223 (N_7223,N_6111,N_6441);
nand U7224 (N_7224,N_6569,N_6016);
nor U7225 (N_7225,N_6433,N_6295);
nor U7226 (N_7226,N_6253,N_6584);
nand U7227 (N_7227,N_6147,N_6693);
and U7228 (N_7228,N_6230,N_6188);
and U7229 (N_7229,N_6026,N_6709);
and U7230 (N_7230,N_6241,N_6432);
nand U7231 (N_7231,N_6154,N_6666);
nand U7232 (N_7232,N_6704,N_6248);
nand U7233 (N_7233,N_6389,N_6698);
or U7234 (N_7234,N_6491,N_6614);
and U7235 (N_7235,N_6230,N_6537);
xor U7236 (N_7236,N_6035,N_6154);
or U7237 (N_7237,N_6419,N_6618);
and U7238 (N_7238,N_6045,N_6509);
nand U7239 (N_7239,N_6484,N_6552);
nand U7240 (N_7240,N_6749,N_6411);
or U7241 (N_7241,N_6745,N_6158);
and U7242 (N_7242,N_6339,N_6348);
and U7243 (N_7243,N_6219,N_6132);
nand U7244 (N_7244,N_6483,N_6197);
or U7245 (N_7245,N_6301,N_6113);
nor U7246 (N_7246,N_6295,N_6616);
and U7247 (N_7247,N_6222,N_6685);
nor U7248 (N_7248,N_6092,N_6098);
nor U7249 (N_7249,N_6071,N_6208);
nor U7250 (N_7250,N_6138,N_6582);
and U7251 (N_7251,N_6649,N_6330);
and U7252 (N_7252,N_6404,N_6080);
nor U7253 (N_7253,N_6680,N_6278);
nor U7254 (N_7254,N_6396,N_6539);
nand U7255 (N_7255,N_6425,N_6142);
nor U7256 (N_7256,N_6189,N_6449);
or U7257 (N_7257,N_6015,N_6184);
nor U7258 (N_7258,N_6707,N_6504);
nand U7259 (N_7259,N_6139,N_6699);
nand U7260 (N_7260,N_6425,N_6034);
nor U7261 (N_7261,N_6371,N_6364);
xor U7262 (N_7262,N_6617,N_6631);
nand U7263 (N_7263,N_6594,N_6530);
or U7264 (N_7264,N_6226,N_6542);
and U7265 (N_7265,N_6556,N_6217);
nor U7266 (N_7266,N_6084,N_6259);
or U7267 (N_7267,N_6735,N_6017);
and U7268 (N_7268,N_6148,N_6014);
or U7269 (N_7269,N_6052,N_6724);
nor U7270 (N_7270,N_6100,N_6110);
xor U7271 (N_7271,N_6661,N_6115);
nor U7272 (N_7272,N_6738,N_6348);
or U7273 (N_7273,N_6321,N_6636);
nor U7274 (N_7274,N_6654,N_6623);
nand U7275 (N_7275,N_6295,N_6012);
nor U7276 (N_7276,N_6504,N_6559);
nor U7277 (N_7277,N_6071,N_6009);
or U7278 (N_7278,N_6083,N_6220);
or U7279 (N_7279,N_6455,N_6243);
nand U7280 (N_7280,N_6732,N_6287);
nor U7281 (N_7281,N_6473,N_6275);
and U7282 (N_7282,N_6029,N_6720);
and U7283 (N_7283,N_6078,N_6262);
xnor U7284 (N_7284,N_6238,N_6129);
nand U7285 (N_7285,N_6711,N_6734);
nor U7286 (N_7286,N_6670,N_6075);
nor U7287 (N_7287,N_6218,N_6144);
nor U7288 (N_7288,N_6738,N_6206);
nand U7289 (N_7289,N_6418,N_6437);
nor U7290 (N_7290,N_6311,N_6159);
xor U7291 (N_7291,N_6081,N_6709);
nand U7292 (N_7292,N_6650,N_6608);
and U7293 (N_7293,N_6049,N_6389);
nor U7294 (N_7294,N_6029,N_6544);
nand U7295 (N_7295,N_6519,N_6536);
nor U7296 (N_7296,N_6148,N_6641);
nor U7297 (N_7297,N_6208,N_6432);
nor U7298 (N_7298,N_6385,N_6331);
nand U7299 (N_7299,N_6673,N_6269);
or U7300 (N_7300,N_6618,N_6592);
xnor U7301 (N_7301,N_6510,N_6532);
nor U7302 (N_7302,N_6040,N_6199);
xnor U7303 (N_7303,N_6472,N_6052);
xnor U7304 (N_7304,N_6221,N_6254);
nand U7305 (N_7305,N_6088,N_6498);
and U7306 (N_7306,N_6454,N_6376);
or U7307 (N_7307,N_6221,N_6665);
nor U7308 (N_7308,N_6256,N_6270);
and U7309 (N_7309,N_6252,N_6659);
and U7310 (N_7310,N_6722,N_6367);
xor U7311 (N_7311,N_6126,N_6411);
or U7312 (N_7312,N_6321,N_6034);
nand U7313 (N_7313,N_6499,N_6279);
and U7314 (N_7314,N_6098,N_6167);
xor U7315 (N_7315,N_6559,N_6107);
nor U7316 (N_7316,N_6421,N_6433);
nand U7317 (N_7317,N_6419,N_6724);
nor U7318 (N_7318,N_6285,N_6181);
or U7319 (N_7319,N_6413,N_6235);
or U7320 (N_7320,N_6360,N_6611);
and U7321 (N_7321,N_6269,N_6056);
nor U7322 (N_7322,N_6713,N_6412);
nand U7323 (N_7323,N_6588,N_6450);
nor U7324 (N_7324,N_6660,N_6618);
nor U7325 (N_7325,N_6220,N_6607);
nand U7326 (N_7326,N_6408,N_6185);
nand U7327 (N_7327,N_6582,N_6455);
nand U7328 (N_7328,N_6545,N_6498);
or U7329 (N_7329,N_6231,N_6201);
nor U7330 (N_7330,N_6684,N_6735);
nand U7331 (N_7331,N_6394,N_6725);
nor U7332 (N_7332,N_6095,N_6348);
nand U7333 (N_7333,N_6210,N_6124);
nand U7334 (N_7334,N_6560,N_6451);
nor U7335 (N_7335,N_6737,N_6511);
and U7336 (N_7336,N_6185,N_6186);
or U7337 (N_7337,N_6282,N_6635);
or U7338 (N_7338,N_6578,N_6270);
and U7339 (N_7339,N_6206,N_6560);
nor U7340 (N_7340,N_6689,N_6291);
and U7341 (N_7341,N_6027,N_6265);
and U7342 (N_7342,N_6577,N_6294);
xnor U7343 (N_7343,N_6513,N_6086);
xor U7344 (N_7344,N_6243,N_6130);
and U7345 (N_7345,N_6179,N_6535);
nor U7346 (N_7346,N_6185,N_6485);
nand U7347 (N_7347,N_6235,N_6287);
xor U7348 (N_7348,N_6533,N_6652);
nand U7349 (N_7349,N_6701,N_6744);
or U7350 (N_7350,N_6444,N_6109);
nor U7351 (N_7351,N_6411,N_6215);
or U7352 (N_7352,N_6573,N_6212);
xor U7353 (N_7353,N_6320,N_6692);
nand U7354 (N_7354,N_6167,N_6699);
or U7355 (N_7355,N_6546,N_6158);
nand U7356 (N_7356,N_6203,N_6666);
nand U7357 (N_7357,N_6120,N_6055);
or U7358 (N_7358,N_6676,N_6090);
xor U7359 (N_7359,N_6184,N_6692);
nor U7360 (N_7360,N_6471,N_6621);
and U7361 (N_7361,N_6523,N_6212);
xor U7362 (N_7362,N_6082,N_6143);
and U7363 (N_7363,N_6103,N_6319);
nand U7364 (N_7364,N_6705,N_6254);
nor U7365 (N_7365,N_6281,N_6030);
xnor U7366 (N_7366,N_6338,N_6675);
xnor U7367 (N_7367,N_6000,N_6612);
xor U7368 (N_7368,N_6442,N_6383);
nand U7369 (N_7369,N_6037,N_6671);
nand U7370 (N_7370,N_6115,N_6586);
nand U7371 (N_7371,N_6113,N_6249);
xnor U7372 (N_7372,N_6287,N_6663);
xor U7373 (N_7373,N_6028,N_6468);
and U7374 (N_7374,N_6338,N_6161);
xor U7375 (N_7375,N_6505,N_6001);
and U7376 (N_7376,N_6029,N_6333);
and U7377 (N_7377,N_6036,N_6722);
nor U7378 (N_7378,N_6305,N_6457);
nand U7379 (N_7379,N_6346,N_6247);
xnor U7380 (N_7380,N_6370,N_6136);
or U7381 (N_7381,N_6162,N_6116);
or U7382 (N_7382,N_6028,N_6492);
and U7383 (N_7383,N_6075,N_6478);
nand U7384 (N_7384,N_6282,N_6218);
and U7385 (N_7385,N_6002,N_6466);
and U7386 (N_7386,N_6665,N_6453);
nand U7387 (N_7387,N_6446,N_6705);
nand U7388 (N_7388,N_6636,N_6416);
and U7389 (N_7389,N_6680,N_6604);
or U7390 (N_7390,N_6415,N_6028);
nand U7391 (N_7391,N_6130,N_6390);
nor U7392 (N_7392,N_6699,N_6094);
and U7393 (N_7393,N_6567,N_6341);
nor U7394 (N_7394,N_6307,N_6453);
and U7395 (N_7395,N_6567,N_6429);
nor U7396 (N_7396,N_6596,N_6330);
and U7397 (N_7397,N_6662,N_6622);
or U7398 (N_7398,N_6617,N_6093);
and U7399 (N_7399,N_6553,N_6459);
and U7400 (N_7400,N_6635,N_6586);
nor U7401 (N_7401,N_6134,N_6411);
xnor U7402 (N_7402,N_6541,N_6462);
nor U7403 (N_7403,N_6277,N_6041);
and U7404 (N_7404,N_6019,N_6109);
and U7405 (N_7405,N_6220,N_6140);
and U7406 (N_7406,N_6480,N_6314);
nand U7407 (N_7407,N_6635,N_6631);
and U7408 (N_7408,N_6567,N_6537);
and U7409 (N_7409,N_6518,N_6738);
nand U7410 (N_7410,N_6509,N_6601);
nor U7411 (N_7411,N_6334,N_6404);
xor U7412 (N_7412,N_6560,N_6399);
nand U7413 (N_7413,N_6020,N_6098);
and U7414 (N_7414,N_6724,N_6565);
or U7415 (N_7415,N_6510,N_6549);
nor U7416 (N_7416,N_6588,N_6075);
xor U7417 (N_7417,N_6583,N_6737);
nor U7418 (N_7418,N_6239,N_6008);
and U7419 (N_7419,N_6043,N_6602);
or U7420 (N_7420,N_6105,N_6127);
or U7421 (N_7421,N_6717,N_6581);
or U7422 (N_7422,N_6104,N_6683);
and U7423 (N_7423,N_6216,N_6215);
or U7424 (N_7424,N_6123,N_6044);
nor U7425 (N_7425,N_6289,N_6412);
nand U7426 (N_7426,N_6490,N_6514);
and U7427 (N_7427,N_6289,N_6309);
and U7428 (N_7428,N_6174,N_6234);
and U7429 (N_7429,N_6167,N_6720);
nor U7430 (N_7430,N_6493,N_6416);
and U7431 (N_7431,N_6539,N_6488);
nor U7432 (N_7432,N_6106,N_6590);
or U7433 (N_7433,N_6708,N_6448);
nand U7434 (N_7434,N_6559,N_6110);
nor U7435 (N_7435,N_6483,N_6324);
nand U7436 (N_7436,N_6333,N_6509);
xnor U7437 (N_7437,N_6262,N_6652);
nor U7438 (N_7438,N_6018,N_6499);
nand U7439 (N_7439,N_6437,N_6283);
and U7440 (N_7440,N_6661,N_6335);
xnor U7441 (N_7441,N_6738,N_6475);
nand U7442 (N_7442,N_6688,N_6693);
and U7443 (N_7443,N_6114,N_6010);
nand U7444 (N_7444,N_6386,N_6599);
nor U7445 (N_7445,N_6232,N_6011);
and U7446 (N_7446,N_6339,N_6100);
and U7447 (N_7447,N_6035,N_6322);
xor U7448 (N_7448,N_6666,N_6254);
xnor U7449 (N_7449,N_6159,N_6412);
nand U7450 (N_7450,N_6741,N_6595);
and U7451 (N_7451,N_6377,N_6744);
and U7452 (N_7452,N_6512,N_6172);
nand U7453 (N_7453,N_6347,N_6565);
nor U7454 (N_7454,N_6723,N_6128);
nand U7455 (N_7455,N_6049,N_6151);
and U7456 (N_7456,N_6149,N_6348);
nand U7457 (N_7457,N_6674,N_6601);
or U7458 (N_7458,N_6381,N_6053);
and U7459 (N_7459,N_6108,N_6114);
or U7460 (N_7460,N_6048,N_6620);
nand U7461 (N_7461,N_6531,N_6030);
and U7462 (N_7462,N_6066,N_6051);
and U7463 (N_7463,N_6036,N_6006);
nand U7464 (N_7464,N_6543,N_6151);
xnor U7465 (N_7465,N_6439,N_6694);
and U7466 (N_7466,N_6200,N_6437);
nor U7467 (N_7467,N_6668,N_6241);
and U7468 (N_7468,N_6112,N_6135);
nor U7469 (N_7469,N_6488,N_6508);
or U7470 (N_7470,N_6115,N_6459);
nor U7471 (N_7471,N_6402,N_6247);
or U7472 (N_7472,N_6028,N_6286);
or U7473 (N_7473,N_6370,N_6710);
and U7474 (N_7474,N_6437,N_6155);
nor U7475 (N_7475,N_6372,N_6573);
nand U7476 (N_7476,N_6121,N_6479);
xor U7477 (N_7477,N_6613,N_6575);
or U7478 (N_7478,N_6256,N_6086);
nand U7479 (N_7479,N_6064,N_6553);
or U7480 (N_7480,N_6529,N_6675);
and U7481 (N_7481,N_6384,N_6060);
or U7482 (N_7482,N_6471,N_6664);
xor U7483 (N_7483,N_6740,N_6038);
nand U7484 (N_7484,N_6263,N_6123);
or U7485 (N_7485,N_6267,N_6328);
and U7486 (N_7486,N_6502,N_6068);
and U7487 (N_7487,N_6712,N_6303);
and U7488 (N_7488,N_6104,N_6354);
and U7489 (N_7489,N_6129,N_6013);
nand U7490 (N_7490,N_6655,N_6596);
nand U7491 (N_7491,N_6659,N_6307);
nand U7492 (N_7492,N_6439,N_6478);
nor U7493 (N_7493,N_6057,N_6711);
nor U7494 (N_7494,N_6399,N_6309);
nor U7495 (N_7495,N_6643,N_6404);
nor U7496 (N_7496,N_6185,N_6455);
nor U7497 (N_7497,N_6278,N_6586);
xnor U7498 (N_7498,N_6710,N_6172);
nor U7499 (N_7499,N_6160,N_6144);
and U7500 (N_7500,N_7499,N_7110);
and U7501 (N_7501,N_7018,N_7376);
or U7502 (N_7502,N_7258,N_7126);
xnor U7503 (N_7503,N_7428,N_6849);
nand U7504 (N_7504,N_7341,N_7083);
or U7505 (N_7505,N_7159,N_7085);
nand U7506 (N_7506,N_7378,N_7465);
or U7507 (N_7507,N_6873,N_6824);
nor U7508 (N_7508,N_7452,N_7448);
or U7509 (N_7509,N_7449,N_7248);
nor U7510 (N_7510,N_7273,N_7160);
nand U7511 (N_7511,N_7068,N_7451);
and U7512 (N_7512,N_6818,N_7205);
and U7513 (N_7513,N_6969,N_6929);
nand U7514 (N_7514,N_7069,N_7458);
xnor U7515 (N_7515,N_7033,N_7350);
and U7516 (N_7516,N_7404,N_7087);
nand U7517 (N_7517,N_7493,N_7256);
nor U7518 (N_7518,N_7460,N_7495);
and U7519 (N_7519,N_7459,N_7268);
nand U7520 (N_7520,N_6756,N_6803);
nor U7521 (N_7521,N_7062,N_7317);
nor U7522 (N_7522,N_7360,N_7239);
and U7523 (N_7523,N_7099,N_6870);
and U7524 (N_7524,N_7130,N_7266);
and U7525 (N_7525,N_6861,N_7027);
nand U7526 (N_7526,N_7283,N_7252);
nor U7527 (N_7527,N_7461,N_7185);
or U7528 (N_7528,N_7399,N_7147);
nor U7529 (N_7529,N_6924,N_7009);
or U7530 (N_7530,N_7082,N_7468);
and U7531 (N_7531,N_7485,N_6753);
or U7532 (N_7532,N_7242,N_7154);
nor U7533 (N_7533,N_7052,N_7223);
or U7534 (N_7534,N_7107,N_7163);
nor U7535 (N_7535,N_6982,N_7080);
nand U7536 (N_7536,N_7171,N_7345);
xnor U7537 (N_7537,N_6856,N_7261);
nor U7538 (N_7538,N_7255,N_7044);
and U7539 (N_7539,N_6758,N_7078);
and U7540 (N_7540,N_7012,N_7395);
or U7541 (N_7541,N_7442,N_7333);
or U7542 (N_7542,N_7029,N_7472);
xnor U7543 (N_7543,N_6876,N_7109);
nand U7544 (N_7544,N_6999,N_6860);
nor U7545 (N_7545,N_7301,N_7422);
nor U7546 (N_7546,N_7151,N_6894);
and U7547 (N_7547,N_6775,N_6781);
nor U7548 (N_7548,N_6839,N_7455);
nand U7549 (N_7549,N_7401,N_7298);
nand U7550 (N_7550,N_7106,N_7469);
or U7551 (N_7551,N_7034,N_7431);
or U7552 (N_7552,N_7416,N_6965);
nor U7553 (N_7553,N_7381,N_6975);
and U7554 (N_7554,N_6897,N_6859);
or U7555 (N_7555,N_7432,N_7028);
or U7556 (N_7556,N_6767,N_6898);
nand U7557 (N_7557,N_7348,N_6778);
nand U7558 (N_7558,N_7128,N_6795);
nor U7559 (N_7559,N_7098,N_7066);
and U7560 (N_7560,N_7453,N_7077);
nand U7561 (N_7561,N_7419,N_6930);
nor U7562 (N_7562,N_7291,N_7129);
and U7563 (N_7563,N_7117,N_6827);
nand U7564 (N_7564,N_6954,N_6782);
and U7565 (N_7565,N_6972,N_6823);
and U7566 (N_7566,N_6939,N_7408);
or U7567 (N_7567,N_6889,N_6980);
and U7568 (N_7568,N_7338,N_7006);
xnor U7569 (N_7569,N_6857,N_6967);
xor U7570 (N_7570,N_7302,N_6991);
and U7571 (N_7571,N_6832,N_7133);
and U7572 (N_7572,N_7375,N_7280);
nor U7573 (N_7573,N_7447,N_6792);
xor U7574 (N_7574,N_7204,N_7116);
nand U7575 (N_7575,N_6874,N_7168);
or U7576 (N_7576,N_7407,N_7347);
nand U7577 (N_7577,N_7328,N_7289);
nand U7578 (N_7578,N_7364,N_6970);
and U7579 (N_7579,N_7002,N_6838);
nand U7580 (N_7580,N_7059,N_6887);
or U7581 (N_7581,N_7037,N_6928);
or U7582 (N_7582,N_7276,N_6985);
nand U7583 (N_7583,N_7307,N_7121);
nand U7584 (N_7584,N_6888,N_7072);
nor U7585 (N_7585,N_7039,N_7195);
nor U7586 (N_7586,N_7101,N_7249);
nor U7587 (N_7587,N_7220,N_6774);
or U7588 (N_7588,N_7342,N_7277);
and U7589 (N_7589,N_7245,N_7226);
xor U7590 (N_7590,N_7122,N_6987);
or U7591 (N_7591,N_6862,N_7411);
nand U7592 (N_7592,N_6846,N_7213);
nor U7593 (N_7593,N_7394,N_7303);
nor U7594 (N_7594,N_6963,N_7065);
nor U7595 (N_7595,N_7016,N_6864);
nor U7596 (N_7596,N_6937,N_6776);
and U7597 (N_7597,N_7306,N_6983);
or U7598 (N_7598,N_7471,N_7405);
nand U7599 (N_7599,N_6932,N_7490);
nand U7600 (N_7600,N_7278,N_7251);
and U7601 (N_7601,N_6953,N_6962);
or U7602 (N_7602,N_7174,N_6907);
nand U7603 (N_7603,N_7186,N_6802);
and U7604 (N_7604,N_7070,N_6808);
nor U7605 (N_7605,N_7218,N_7125);
nand U7606 (N_7606,N_7362,N_6973);
nor U7607 (N_7607,N_7021,N_6935);
or U7608 (N_7608,N_7030,N_7424);
nand U7609 (N_7609,N_6750,N_7361);
and U7610 (N_7610,N_7073,N_7315);
or U7611 (N_7611,N_7093,N_7231);
nor U7612 (N_7612,N_7373,N_7253);
nand U7613 (N_7613,N_7152,N_7353);
or U7614 (N_7614,N_6918,N_7235);
nor U7615 (N_7615,N_6994,N_7190);
nor U7616 (N_7616,N_6780,N_6919);
nor U7617 (N_7617,N_7228,N_6797);
nor U7618 (N_7618,N_6946,N_7167);
nand U7619 (N_7619,N_7118,N_7246);
nand U7620 (N_7620,N_6825,N_6988);
nor U7621 (N_7621,N_7380,N_7368);
nand U7622 (N_7622,N_7091,N_7053);
and U7623 (N_7623,N_7429,N_6942);
or U7624 (N_7624,N_6995,N_7075);
nand U7625 (N_7625,N_7300,N_6763);
or U7626 (N_7626,N_7232,N_7427);
nand U7627 (N_7627,N_7412,N_7187);
and U7628 (N_7628,N_6842,N_7288);
or U7629 (N_7629,N_7094,N_7445);
and U7630 (N_7630,N_7150,N_7135);
nand U7631 (N_7631,N_7201,N_7279);
and U7632 (N_7632,N_7247,N_7169);
and U7633 (N_7633,N_7113,N_6905);
nor U7634 (N_7634,N_7084,N_7414);
nand U7635 (N_7635,N_7036,N_7383);
xnor U7636 (N_7636,N_7095,N_7311);
and U7637 (N_7637,N_7146,N_7209);
or U7638 (N_7638,N_6976,N_7225);
and U7639 (N_7639,N_7370,N_7153);
or U7640 (N_7640,N_7259,N_7263);
and U7641 (N_7641,N_7024,N_6866);
or U7642 (N_7642,N_7346,N_7140);
or U7643 (N_7643,N_6891,N_6850);
nand U7644 (N_7644,N_7041,N_7097);
nand U7645 (N_7645,N_6852,N_7144);
nor U7646 (N_7646,N_7202,N_6977);
nand U7647 (N_7647,N_7296,N_7057);
nor U7648 (N_7648,N_6848,N_6789);
and U7649 (N_7649,N_6920,N_7477);
nand U7650 (N_7650,N_7323,N_7011);
or U7651 (N_7651,N_7271,N_7339);
nor U7652 (N_7652,N_7275,N_6810);
xor U7653 (N_7653,N_7054,N_7038);
and U7654 (N_7654,N_7064,N_7074);
or U7655 (N_7655,N_7337,N_6978);
or U7656 (N_7656,N_7352,N_6950);
nand U7657 (N_7657,N_6794,N_7270);
nand U7658 (N_7658,N_7387,N_6882);
nor U7659 (N_7659,N_6964,N_6801);
and U7660 (N_7660,N_7162,N_7181);
nor U7661 (N_7661,N_6791,N_7250);
nand U7662 (N_7662,N_7148,N_7332);
nand U7663 (N_7663,N_6817,N_7123);
xor U7664 (N_7664,N_7141,N_6771);
or U7665 (N_7665,N_7384,N_7262);
or U7666 (N_7666,N_6971,N_7003);
nand U7667 (N_7667,N_6940,N_7219);
xnor U7668 (N_7668,N_7484,N_6768);
xnor U7669 (N_7669,N_6910,N_7145);
or U7670 (N_7670,N_7287,N_7425);
nand U7671 (N_7671,N_7402,N_6865);
and U7672 (N_7672,N_7436,N_6952);
xnor U7673 (N_7673,N_7045,N_7418);
and U7674 (N_7674,N_7194,N_7216);
nor U7675 (N_7675,N_7048,N_7238);
or U7676 (N_7676,N_7388,N_7108);
or U7677 (N_7677,N_6974,N_7004);
or U7678 (N_7678,N_7481,N_7371);
nor U7679 (N_7679,N_7227,N_7055);
nor U7680 (N_7680,N_7031,N_7358);
or U7681 (N_7681,N_7413,N_6947);
or U7682 (N_7682,N_7179,N_6812);
xnor U7683 (N_7683,N_7178,N_6902);
or U7684 (N_7684,N_6908,N_6996);
and U7685 (N_7685,N_7446,N_7274);
and U7686 (N_7686,N_6958,N_6800);
nor U7687 (N_7687,N_7026,N_6949);
nor U7688 (N_7688,N_7417,N_6884);
and U7689 (N_7689,N_7096,N_6813);
and U7690 (N_7690,N_7473,N_7357);
or U7691 (N_7691,N_7184,N_7489);
or U7692 (N_7692,N_7180,N_7382);
nand U7693 (N_7693,N_6904,N_7421);
nand U7694 (N_7694,N_6868,N_7423);
xnor U7695 (N_7695,N_6843,N_7215);
and U7696 (N_7696,N_6820,N_6805);
xor U7697 (N_7697,N_7136,N_6909);
or U7698 (N_7698,N_7203,N_7139);
nand U7699 (N_7699,N_7237,N_6764);
xor U7700 (N_7700,N_7325,N_7114);
or U7701 (N_7701,N_7496,N_7229);
nand U7702 (N_7702,N_7450,N_6806);
nor U7703 (N_7703,N_7343,N_7020);
or U7704 (N_7704,N_7284,N_6811);
and U7705 (N_7705,N_7001,N_6881);
nor U7706 (N_7706,N_6793,N_6968);
or U7707 (N_7707,N_7115,N_7089);
nor U7708 (N_7708,N_7254,N_6867);
nor U7709 (N_7709,N_7119,N_7032);
or U7710 (N_7710,N_6921,N_7047);
nand U7711 (N_7711,N_7314,N_7206);
nand U7712 (N_7712,N_7243,N_7463);
or U7713 (N_7713,N_7297,N_6784);
or U7714 (N_7714,N_6804,N_7497);
nor U7715 (N_7715,N_7067,N_7088);
or U7716 (N_7716,N_7329,N_6770);
nand U7717 (N_7717,N_7340,N_6998);
nand U7718 (N_7718,N_7111,N_6913);
or U7719 (N_7719,N_6948,N_7025);
nor U7720 (N_7720,N_7158,N_7410);
and U7721 (N_7721,N_7236,N_7183);
or U7722 (N_7722,N_7486,N_6788);
and U7723 (N_7723,N_6922,N_7369);
and U7724 (N_7724,N_7155,N_6835);
nor U7725 (N_7725,N_7105,N_7050);
nor U7726 (N_7726,N_7210,N_7351);
xnor U7727 (N_7727,N_6809,N_6822);
or U7728 (N_7728,N_6834,N_7035);
or U7729 (N_7729,N_7440,N_7367);
and U7730 (N_7730,N_7157,N_6819);
xor U7731 (N_7731,N_7019,N_7389);
and U7732 (N_7732,N_6847,N_7175);
and U7733 (N_7733,N_7005,N_6993);
nand U7734 (N_7734,N_7363,N_6941);
nor U7735 (N_7735,N_7433,N_7292);
nand U7736 (N_7736,N_7426,N_7222);
nor U7737 (N_7737,N_7331,N_7170);
nand U7738 (N_7738,N_6875,N_6833);
nand U7739 (N_7739,N_6761,N_6772);
and U7740 (N_7740,N_7046,N_7334);
and U7741 (N_7741,N_6917,N_7164);
or U7742 (N_7742,N_6877,N_7304);
nand U7743 (N_7743,N_6960,N_7318);
nor U7744 (N_7744,N_7439,N_6851);
nor U7745 (N_7745,N_7349,N_7177);
nor U7746 (N_7746,N_7385,N_7198);
nand U7747 (N_7747,N_6837,N_6836);
nand U7748 (N_7748,N_6798,N_7120);
nand U7749 (N_7749,N_6777,N_6992);
or U7750 (N_7750,N_6979,N_6931);
nand U7751 (N_7751,N_7372,N_6886);
or U7752 (N_7752,N_7007,N_7308);
nor U7753 (N_7753,N_6989,N_7161);
and U7754 (N_7754,N_6906,N_7063);
or U7755 (N_7755,N_7134,N_7230);
nand U7756 (N_7756,N_7142,N_7056);
and U7757 (N_7757,N_6762,N_7386);
nor U7758 (N_7758,N_6872,N_6853);
nand U7759 (N_7759,N_6914,N_7000);
nand U7760 (N_7760,N_6844,N_7071);
nor U7761 (N_7761,N_7374,N_7359);
or U7762 (N_7762,N_6783,N_6911);
nor U7763 (N_7763,N_6769,N_7061);
and U7764 (N_7764,N_7397,N_6945);
nor U7765 (N_7765,N_7207,N_6855);
or U7766 (N_7766,N_7400,N_6934);
nand U7767 (N_7767,N_6943,N_6916);
and U7768 (N_7768,N_7430,N_7269);
and U7769 (N_7769,N_6807,N_7149);
nand U7770 (N_7770,N_7335,N_6821);
nor U7771 (N_7771,N_7293,N_6944);
nor U7772 (N_7772,N_6990,N_6830);
xor U7773 (N_7773,N_7420,N_7435);
and U7774 (N_7774,N_6893,N_7282);
nand U7775 (N_7775,N_7132,N_6936);
nor U7776 (N_7776,N_6899,N_7172);
and U7777 (N_7777,N_6869,N_7138);
nand U7778 (N_7778,N_7487,N_7467);
nor U7779 (N_7779,N_6759,N_6878);
or U7780 (N_7780,N_7354,N_7131);
or U7781 (N_7781,N_7379,N_7390);
and U7782 (N_7782,N_7299,N_7173);
nand U7783 (N_7783,N_7079,N_7010);
or U7784 (N_7784,N_7267,N_7051);
and U7785 (N_7785,N_6986,N_7244);
nand U7786 (N_7786,N_7214,N_7092);
or U7787 (N_7787,N_6752,N_6841);
or U7788 (N_7788,N_7224,N_7377);
nand U7789 (N_7789,N_7316,N_6933);
nand U7790 (N_7790,N_7112,N_6915);
and U7791 (N_7791,N_7365,N_7176);
nand U7792 (N_7792,N_6787,N_7193);
xnor U7793 (N_7793,N_7286,N_7124);
nand U7794 (N_7794,N_6923,N_6895);
nand U7795 (N_7795,N_7321,N_6892);
nand U7796 (N_7796,N_7281,N_7392);
nor U7797 (N_7797,N_7211,N_7208);
nor U7798 (N_7798,N_7441,N_6961);
or U7799 (N_7799,N_7196,N_6785);
nand U7800 (N_7800,N_7295,N_7474);
nand U7801 (N_7801,N_7454,N_7086);
xnor U7802 (N_7802,N_7366,N_7310);
and U7803 (N_7803,N_7466,N_6956);
nand U7804 (N_7804,N_7457,N_7192);
nor U7805 (N_7805,N_7217,N_6966);
or U7806 (N_7806,N_7102,N_6951);
or U7807 (N_7807,N_6845,N_6754);
nor U7808 (N_7808,N_6863,N_7438);
nor U7809 (N_7809,N_6840,N_7240);
and U7810 (N_7810,N_7494,N_7257);
nor U7811 (N_7811,N_7322,N_7188);
or U7812 (N_7812,N_7156,N_6815);
nand U7813 (N_7813,N_7103,N_7327);
or U7814 (N_7814,N_7023,N_6900);
nor U7815 (N_7815,N_6959,N_7498);
nor U7816 (N_7816,N_7393,N_7040);
nor U7817 (N_7817,N_7015,N_7464);
nor U7818 (N_7818,N_6829,N_6854);
nor U7819 (N_7819,N_6927,N_7309);
or U7820 (N_7820,N_6885,N_7391);
or U7821 (N_7821,N_6912,N_7081);
nor U7822 (N_7822,N_6799,N_6765);
nand U7823 (N_7823,N_7221,N_7189);
nor U7824 (N_7824,N_6981,N_7199);
nor U7825 (N_7825,N_6826,N_7022);
nor U7826 (N_7826,N_7415,N_7165);
and U7827 (N_7827,N_6790,N_7197);
and U7828 (N_7828,N_6955,N_6997);
nand U7829 (N_7829,N_7013,N_6883);
nor U7830 (N_7830,N_7137,N_6751);
nor U7831 (N_7831,N_6779,N_7483);
or U7832 (N_7832,N_6925,N_6828);
nand U7833 (N_7833,N_6760,N_7320);
nand U7834 (N_7834,N_7212,N_7017);
nor U7835 (N_7835,N_7492,N_7014);
or U7836 (N_7836,N_6766,N_7356);
and U7837 (N_7837,N_7488,N_7104);
or U7838 (N_7838,N_7234,N_7058);
or U7839 (N_7839,N_7478,N_6984);
and U7840 (N_7840,N_7233,N_6938);
nor U7841 (N_7841,N_7265,N_6757);
xnor U7842 (N_7842,N_7312,N_7403);
nand U7843 (N_7843,N_7042,N_7272);
and U7844 (N_7844,N_7100,N_7470);
nand U7845 (N_7845,N_7008,N_6896);
nand U7846 (N_7846,N_6903,N_6901);
nor U7847 (N_7847,N_7191,N_6773);
and U7848 (N_7848,N_7443,N_6786);
or U7849 (N_7849,N_7290,N_7182);
and U7850 (N_7850,N_7396,N_7409);
nor U7851 (N_7851,N_7294,N_7076);
nand U7852 (N_7852,N_7305,N_6755);
xnor U7853 (N_7853,N_7437,N_7406);
nand U7854 (N_7854,N_6926,N_7444);
and U7855 (N_7855,N_7049,N_7355);
and U7856 (N_7856,N_6858,N_6880);
or U7857 (N_7857,N_7398,N_7127);
nor U7858 (N_7858,N_7264,N_6814);
or U7859 (N_7859,N_7475,N_7143);
nand U7860 (N_7860,N_7479,N_6871);
or U7861 (N_7861,N_6957,N_7456);
nor U7862 (N_7862,N_7060,N_6831);
nand U7863 (N_7863,N_6796,N_6890);
nor U7864 (N_7864,N_7324,N_7319);
or U7865 (N_7865,N_7326,N_7330);
or U7866 (N_7866,N_7260,N_7344);
xor U7867 (N_7867,N_7313,N_7043);
nor U7868 (N_7868,N_7241,N_6816);
nor U7869 (N_7869,N_7166,N_7090);
xor U7870 (N_7870,N_6879,N_7491);
or U7871 (N_7871,N_7480,N_7336);
xnor U7872 (N_7872,N_7462,N_7482);
nand U7873 (N_7873,N_7285,N_7476);
and U7874 (N_7874,N_7200,N_7434);
or U7875 (N_7875,N_7327,N_7471);
or U7876 (N_7876,N_7137,N_7218);
and U7877 (N_7877,N_7442,N_7434);
nand U7878 (N_7878,N_6963,N_6803);
nand U7879 (N_7879,N_6942,N_7267);
and U7880 (N_7880,N_7267,N_6862);
and U7881 (N_7881,N_6890,N_7090);
and U7882 (N_7882,N_7258,N_7313);
and U7883 (N_7883,N_6992,N_7125);
xor U7884 (N_7884,N_7254,N_7208);
nand U7885 (N_7885,N_7155,N_7079);
or U7886 (N_7886,N_7181,N_7117);
and U7887 (N_7887,N_6843,N_6844);
and U7888 (N_7888,N_7001,N_6937);
xnor U7889 (N_7889,N_7139,N_7380);
nor U7890 (N_7890,N_7099,N_6802);
or U7891 (N_7891,N_6842,N_6755);
nor U7892 (N_7892,N_6977,N_7424);
or U7893 (N_7893,N_7324,N_7165);
and U7894 (N_7894,N_7233,N_7495);
nor U7895 (N_7895,N_7430,N_6813);
nor U7896 (N_7896,N_6916,N_6996);
nor U7897 (N_7897,N_7400,N_7407);
and U7898 (N_7898,N_7220,N_7334);
nor U7899 (N_7899,N_7128,N_7236);
and U7900 (N_7900,N_7268,N_7265);
and U7901 (N_7901,N_7451,N_7411);
and U7902 (N_7902,N_6985,N_6810);
nor U7903 (N_7903,N_7147,N_7178);
or U7904 (N_7904,N_7407,N_6956);
nor U7905 (N_7905,N_7267,N_7262);
and U7906 (N_7906,N_7013,N_7390);
nor U7907 (N_7907,N_6891,N_6883);
or U7908 (N_7908,N_6827,N_7258);
and U7909 (N_7909,N_7320,N_7251);
and U7910 (N_7910,N_7099,N_7199);
nor U7911 (N_7911,N_7370,N_7250);
or U7912 (N_7912,N_7475,N_7091);
or U7913 (N_7913,N_6772,N_7021);
or U7914 (N_7914,N_7337,N_7312);
nor U7915 (N_7915,N_7443,N_7174);
or U7916 (N_7916,N_6813,N_6904);
nor U7917 (N_7917,N_6822,N_6918);
nor U7918 (N_7918,N_7316,N_6941);
nor U7919 (N_7919,N_7189,N_6895);
xor U7920 (N_7920,N_6877,N_7203);
xor U7921 (N_7921,N_6818,N_7296);
and U7922 (N_7922,N_7421,N_7492);
xnor U7923 (N_7923,N_7241,N_7103);
and U7924 (N_7924,N_7026,N_7359);
and U7925 (N_7925,N_7351,N_6931);
nor U7926 (N_7926,N_7456,N_7102);
and U7927 (N_7927,N_6960,N_7167);
nor U7928 (N_7928,N_6884,N_6953);
nand U7929 (N_7929,N_6966,N_7481);
nor U7930 (N_7930,N_7143,N_7499);
or U7931 (N_7931,N_7289,N_7163);
xnor U7932 (N_7932,N_7233,N_7066);
and U7933 (N_7933,N_7124,N_6805);
nand U7934 (N_7934,N_6914,N_6966);
or U7935 (N_7935,N_6909,N_6993);
or U7936 (N_7936,N_7433,N_7257);
and U7937 (N_7937,N_7327,N_6777);
or U7938 (N_7938,N_7468,N_7418);
and U7939 (N_7939,N_7496,N_7440);
xnor U7940 (N_7940,N_7185,N_7117);
xnor U7941 (N_7941,N_6919,N_7375);
nand U7942 (N_7942,N_7128,N_7055);
or U7943 (N_7943,N_7130,N_7464);
xor U7944 (N_7944,N_7234,N_6917);
or U7945 (N_7945,N_6906,N_7313);
and U7946 (N_7946,N_7003,N_6859);
or U7947 (N_7947,N_6965,N_6891);
xnor U7948 (N_7948,N_7066,N_6995);
nor U7949 (N_7949,N_7322,N_7462);
nand U7950 (N_7950,N_7252,N_6871);
nand U7951 (N_7951,N_7199,N_6767);
and U7952 (N_7952,N_7360,N_7337);
nor U7953 (N_7953,N_7234,N_7413);
or U7954 (N_7954,N_7411,N_6989);
nor U7955 (N_7955,N_6979,N_6802);
nor U7956 (N_7956,N_7178,N_7045);
or U7957 (N_7957,N_7314,N_6812);
and U7958 (N_7958,N_7239,N_7199);
xnor U7959 (N_7959,N_6891,N_7458);
or U7960 (N_7960,N_7487,N_7052);
xor U7961 (N_7961,N_6839,N_6849);
and U7962 (N_7962,N_7316,N_6935);
nor U7963 (N_7963,N_7343,N_6754);
nand U7964 (N_7964,N_7429,N_7262);
nand U7965 (N_7965,N_6807,N_6764);
and U7966 (N_7966,N_6830,N_7242);
xor U7967 (N_7967,N_7265,N_7241);
xor U7968 (N_7968,N_7423,N_6873);
nand U7969 (N_7969,N_7126,N_7477);
xor U7970 (N_7970,N_6827,N_6852);
nor U7971 (N_7971,N_6802,N_7348);
xnor U7972 (N_7972,N_7106,N_7284);
or U7973 (N_7973,N_7040,N_7240);
nand U7974 (N_7974,N_6915,N_7239);
nand U7975 (N_7975,N_7472,N_7410);
xor U7976 (N_7976,N_6989,N_7332);
nor U7977 (N_7977,N_6784,N_6937);
nor U7978 (N_7978,N_7003,N_6900);
or U7979 (N_7979,N_7377,N_7223);
nor U7980 (N_7980,N_6911,N_6936);
nand U7981 (N_7981,N_6784,N_7044);
nand U7982 (N_7982,N_6975,N_7471);
or U7983 (N_7983,N_6911,N_6809);
and U7984 (N_7984,N_7444,N_7045);
or U7985 (N_7985,N_7496,N_6835);
and U7986 (N_7986,N_6856,N_7443);
or U7987 (N_7987,N_7267,N_7260);
nand U7988 (N_7988,N_7137,N_7099);
nand U7989 (N_7989,N_6999,N_7161);
and U7990 (N_7990,N_7407,N_7289);
nand U7991 (N_7991,N_6800,N_6953);
xor U7992 (N_7992,N_7250,N_6993);
nand U7993 (N_7993,N_7031,N_7308);
nor U7994 (N_7994,N_6874,N_7300);
nor U7995 (N_7995,N_7117,N_7259);
and U7996 (N_7996,N_7340,N_7133);
xor U7997 (N_7997,N_7128,N_6966);
xor U7998 (N_7998,N_6886,N_7408);
nor U7999 (N_7999,N_6770,N_6819);
or U8000 (N_8000,N_7207,N_6834);
nor U8001 (N_8001,N_7042,N_7010);
or U8002 (N_8002,N_7388,N_6973);
or U8003 (N_8003,N_7301,N_6875);
nor U8004 (N_8004,N_6846,N_7192);
nand U8005 (N_8005,N_7058,N_6783);
nand U8006 (N_8006,N_7289,N_7454);
nor U8007 (N_8007,N_7152,N_7467);
xnor U8008 (N_8008,N_6970,N_6913);
and U8009 (N_8009,N_7332,N_7159);
nor U8010 (N_8010,N_7449,N_6929);
and U8011 (N_8011,N_7014,N_7478);
and U8012 (N_8012,N_7430,N_7107);
nand U8013 (N_8013,N_7350,N_6833);
and U8014 (N_8014,N_7427,N_7146);
xnor U8015 (N_8015,N_7262,N_7207);
nand U8016 (N_8016,N_7225,N_7433);
nor U8017 (N_8017,N_7152,N_7395);
nor U8018 (N_8018,N_6804,N_7342);
or U8019 (N_8019,N_7324,N_7265);
nor U8020 (N_8020,N_7420,N_7414);
nand U8021 (N_8021,N_7190,N_6804);
nor U8022 (N_8022,N_6796,N_6912);
nor U8023 (N_8023,N_6855,N_7438);
and U8024 (N_8024,N_7109,N_7260);
and U8025 (N_8025,N_7446,N_7011);
nor U8026 (N_8026,N_6831,N_7131);
or U8027 (N_8027,N_6922,N_7446);
nand U8028 (N_8028,N_6775,N_7165);
nand U8029 (N_8029,N_7074,N_6965);
xnor U8030 (N_8030,N_6901,N_6974);
or U8031 (N_8031,N_7010,N_6922);
and U8032 (N_8032,N_6942,N_7138);
nor U8033 (N_8033,N_7055,N_7286);
nand U8034 (N_8034,N_7406,N_7110);
or U8035 (N_8035,N_7320,N_6936);
or U8036 (N_8036,N_6982,N_7348);
nor U8037 (N_8037,N_7077,N_7020);
and U8038 (N_8038,N_6914,N_6957);
nor U8039 (N_8039,N_7163,N_7421);
xnor U8040 (N_8040,N_7103,N_7294);
and U8041 (N_8041,N_7319,N_7123);
nor U8042 (N_8042,N_7103,N_7023);
nand U8043 (N_8043,N_7370,N_6851);
nand U8044 (N_8044,N_6951,N_7366);
or U8045 (N_8045,N_6856,N_7005);
or U8046 (N_8046,N_6762,N_7006);
nor U8047 (N_8047,N_6993,N_7001);
and U8048 (N_8048,N_7435,N_6778);
or U8049 (N_8049,N_7298,N_7247);
nand U8050 (N_8050,N_6841,N_7262);
and U8051 (N_8051,N_7247,N_6877);
xnor U8052 (N_8052,N_7381,N_7426);
and U8053 (N_8053,N_6778,N_7357);
or U8054 (N_8054,N_6980,N_7136);
nand U8055 (N_8055,N_7448,N_6778);
or U8056 (N_8056,N_7375,N_6988);
nand U8057 (N_8057,N_7280,N_7191);
and U8058 (N_8058,N_6948,N_6875);
nor U8059 (N_8059,N_7480,N_6835);
and U8060 (N_8060,N_7314,N_7349);
nor U8061 (N_8061,N_7189,N_7363);
nand U8062 (N_8062,N_7032,N_7410);
and U8063 (N_8063,N_7429,N_7172);
xor U8064 (N_8064,N_7157,N_6836);
nand U8065 (N_8065,N_7136,N_6998);
nor U8066 (N_8066,N_6766,N_6846);
and U8067 (N_8067,N_7252,N_7473);
or U8068 (N_8068,N_7255,N_7175);
and U8069 (N_8069,N_7420,N_7174);
nand U8070 (N_8070,N_7247,N_7401);
and U8071 (N_8071,N_6966,N_6814);
nor U8072 (N_8072,N_6884,N_7013);
and U8073 (N_8073,N_7340,N_6961);
nand U8074 (N_8074,N_7137,N_7209);
nand U8075 (N_8075,N_7166,N_6773);
xor U8076 (N_8076,N_6859,N_7150);
xor U8077 (N_8077,N_6795,N_7168);
nor U8078 (N_8078,N_7247,N_7021);
nor U8079 (N_8079,N_6904,N_7130);
nor U8080 (N_8080,N_7293,N_6861);
nor U8081 (N_8081,N_7124,N_7224);
or U8082 (N_8082,N_7368,N_6875);
nor U8083 (N_8083,N_7223,N_6875);
and U8084 (N_8084,N_7198,N_7255);
or U8085 (N_8085,N_7064,N_7435);
and U8086 (N_8086,N_7472,N_7342);
xnor U8087 (N_8087,N_6782,N_7066);
and U8088 (N_8088,N_7053,N_6750);
xnor U8089 (N_8089,N_7439,N_6767);
xnor U8090 (N_8090,N_7254,N_6814);
nand U8091 (N_8091,N_6990,N_7215);
and U8092 (N_8092,N_7153,N_7149);
nor U8093 (N_8093,N_7387,N_6753);
nor U8094 (N_8094,N_7098,N_7387);
or U8095 (N_8095,N_7178,N_6769);
xnor U8096 (N_8096,N_6931,N_6879);
nand U8097 (N_8097,N_7340,N_7042);
and U8098 (N_8098,N_7372,N_6849);
and U8099 (N_8099,N_6899,N_6844);
and U8100 (N_8100,N_7181,N_6939);
nand U8101 (N_8101,N_7270,N_7139);
or U8102 (N_8102,N_7295,N_7456);
or U8103 (N_8103,N_7294,N_6822);
nor U8104 (N_8104,N_7030,N_7197);
or U8105 (N_8105,N_6800,N_7439);
nand U8106 (N_8106,N_7297,N_7047);
or U8107 (N_8107,N_7337,N_7377);
nor U8108 (N_8108,N_7333,N_6887);
nand U8109 (N_8109,N_6988,N_6813);
or U8110 (N_8110,N_7183,N_6940);
nand U8111 (N_8111,N_7189,N_7373);
nor U8112 (N_8112,N_7181,N_7079);
xor U8113 (N_8113,N_6865,N_7245);
and U8114 (N_8114,N_6968,N_7014);
and U8115 (N_8115,N_6837,N_7237);
nand U8116 (N_8116,N_6949,N_7207);
nor U8117 (N_8117,N_7217,N_7276);
and U8118 (N_8118,N_7010,N_6813);
or U8119 (N_8119,N_7010,N_6902);
or U8120 (N_8120,N_7317,N_7280);
or U8121 (N_8121,N_7378,N_7185);
and U8122 (N_8122,N_7444,N_6958);
nor U8123 (N_8123,N_6838,N_6993);
nor U8124 (N_8124,N_6752,N_7136);
nand U8125 (N_8125,N_6765,N_7012);
nor U8126 (N_8126,N_7252,N_7420);
or U8127 (N_8127,N_7376,N_6982);
nand U8128 (N_8128,N_6973,N_7431);
nand U8129 (N_8129,N_7207,N_6849);
nand U8130 (N_8130,N_7297,N_7066);
nand U8131 (N_8131,N_7177,N_7043);
or U8132 (N_8132,N_6911,N_7315);
nor U8133 (N_8133,N_6971,N_7221);
xnor U8134 (N_8134,N_7268,N_7386);
nand U8135 (N_8135,N_7435,N_7339);
or U8136 (N_8136,N_6814,N_6957);
nand U8137 (N_8137,N_7272,N_6984);
and U8138 (N_8138,N_7027,N_6905);
nand U8139 (N_8139,N_7095,N_6928);
nand U8140 (N_8140,N_7303,N_6882);
or U8141 (N_8141,N_7245,N_6838);
nand U8142 (N_8142,N_7283,N_7221);
nor U8143 (N_8143,N_6937,N_7479);
or U8144 (N_8144,N_7154,N_7096);
or U8145 (N_8145,N_7102,N_6979);
and U8146 (N_8146,N_7287,N_7337);
and U8147 (N_8147,N_7398,N_7227);
or U8148 (N_8148,N_7467,N_7086);
nand U8149 (N_8149,N_7497,N_7041);
and U8150 (N_8150,N_7114,N_7273);
xor U8151 (N_8151,N_7161,N_7499);
and U8152 (N_8152,N_7336,N_6940);
or U8153 (N_8153,N_6956,N_7025);
nor U8154 (N_8154,N_7128,N_6833);
and U8155 (N_8155,N_7337,N_7112);
and U8156 (N_8156,N_7438,N_6989);
or U8157 (N_8157,N_7107,N_6958);
and U8158 (N_8158,N_7238,N_7181);
and U8159 (N_8159,N_7124,N_7417);
and U8160 (N_8160,N_7068,N_6874);
xnor U8161 (N_8161,N_7444,N_7250);
or U8162 (N_8162,N_7396,N_7115);
nor U8163 (N_8163,N_7238,N_7077);
nor U8164 (N_8164,N_6888,N_6915);
nand U8165 (N_8165,N_7315,N_6834);
or U8166 (N_8166,N_7465,N_6784);
or U8167 (N_8167,N_7361,N_7133);
nor U8168 (N_8168,N_7018,N_6777);
nand U8169 (N_8169,N_7294,N_7295);
nand U8170 (N_8170,N_6928,N_6797);
and U8171 (N_8171,N_6990,N_7258);
and U8172 (N_8172,N_7422,N_7212);
or U8173 (N_8173,N_6894,N_6893);
and U8174 (N_8174,N_6759,N_7164);
xor U8175 (N_8175,N_7096,N_6792);
nor U8176 (N_8176,N_7093,N_6755);
nor U8177 (N_8177,N_6810,N_7049);
and U8178 (N_8178,N_7020,N_6813);
or U8179 (N_8179,N_7211,N_6852);
and U8180 (N_8180,N_6942,N_6774);
or U8181 (N_8181,N_6880,N_7288);
and U8182 (N_8182,N_7141,N_6836);
nor U8183 (N_8183,N_7142,N_7361);
and U8184 (N_8184,N_6827,N_7402);
nand U8185 (N_8185,N_7478,N_7161);
nand U8186 (N_8186,N_7150,N_6787);
and U8187 (N_8187,N_7225,N_6967);
nand U8188 (N_8188,N_6928,N_7316);
and U8189 (N_8189,N_7316,N_6910);
nand U8190 (N_8190,N_6974,N_7265);
or U8191 (N_8191,N_7355,N_7043);
nor U8192 (N_8192,N_7136,N_6983);
nand U8193 (N_8193,N_7343,N_7337);
and U8194 (N_8194,N_7061,N_6799);
nor U8195 (N_8195,N_7062,N_7164);
nor U8196 (N_8196,N_7066,N_7230);
nand U8197 (N_8197,N_7059,N_7291);
nor U8198 (N_8198,N_7284,N_7025);
nor U8199 (N_8199,N_7126,N_6981);
nor U8200 (N_8200,N_7435,N_7424);
nand U8201 (N_8201,N_6820,N_7431);
xor U8202 (N_8202,N_7091,N_6756);
nor U8203 (N_8203,N_7383,N_7112);
or U8204 (N_8204,N_7177,N_6975);
nor U8205 (N_8205,N_6763,N_7472);
and U8206 (N_8206,N_6961,N_7099);
nand U8207 (N_8207,N_7050,N_7498);
or U8208 (N_8208,N_7288,N_6831);
and U8209 (N_8209,N_7330,N_7037);
or U8210 (N_8210,N_7069,N_7437);
or U8211 (N_8211,N_7179,N_6922);
and U8212 (N_8212,N_7326,N_7248);
nand U8213 (N_8213,N_6965,N_7211);
and U8214 (N_8214,N_6919,N_7018);
nor U8215 (N_8215,N_6952,N_6921);
and U8216 (N_8216,N_7005,N_7304);
nor U8217 (N_8217,N_7411,N_6893);
nor U8218 (N_8218,N_6858,N_7013);
and U8219 (N_8219,N_7252,N_6931);
nor U8220 (N_8220,N_7003,N_7270);
and U8221 (N_8221,N_7377,N_7395);
nand U8222 (N_8222,N_6861,N_7211);
and U8223 (N_8223,N_6917,N_7357);
nand U8224 (N_8224,N_7232,N_6972);
and U8225 (N_8225,N_7374,N_7424);
or U8226 (N_8226,N_6825,N_7058);
nor U8227 (N_8227,N_7215,N_6872);
or U8228 (N_8228,N_7242,N_6860);
and U8229 (N_8229,N_7073,N_7492);
nor U8230 (N_8230,N_6855,N_6908);
nor U8231 (N_8231,N_7288,N_7473);
nand U8232 (N_8232,N_6978,N_6849);
and U8233 (N_8233,N_6957,N_7044);
nand U8234 (N_8234,N_7458,N_6950);
nor U8235 (N_8235,N_7201,N_7399);
nor U8236 (N_8236,N_7436,N_7413);
or U8237 (N_8237,N_7144,N_7483);
and U8238 (N_8238,N_6836,N_6956);
nand U8239 (N_8239,N_7362,N_6842);
and U8240 (N_8240,N_6820,N_6760);
nor U8241 (N_8241,N_7287,N_6927);
or U8242 (N_8242,N_7443,N_7341);
xnor U8243 (N_8243,N_7219,N_6906);
and U8244 (N_8244,N_7458,N_7449);
or U8245 (N_8245,N_7262,N_6809);
or U8246 (N_8246,N_7359,N_7409);
and U8247 (N_8247,N_6808,N_6841);
or U8248 (N_8248,N_7224,N_7468);
xnor U8249 (N_8249,N_7390,N_7477);
nor U8250 (N_8250,N_7666,N_7517);
nand U8251 (N_8251,N_7612,N_7539);
nand U8252 (N_8252,N_7778,N_7685);
nor U8253 (N_8253,N_7523,N_8023);
nor U8254 (N_8254,N_7691,N_7514);
nand U8255 (N_8255,N_8029,N_7821);
or U8256 (N_8256,N_7674,N_7746);
nor U8257 (N_8257,N_7684,N_8166);
nor U8258 (N_8258,N_8122,N_7926);
nor U8259 (N_8259,N_8139,N_7594);
and U8260 (N_8260,N_8054,N_7629);
and U8261 (N_8261,N_7942,N_7974);
nand U8262 (N_8262,N_7921,N_7797);
or U8263 (N_8263,N_7544,N_7824);
xnor U8264 (N_8264,N_8144,N_8039);
nor U8265 (N_8265,N_8151,N_7796);
xnor U8266 (N_8266,N_7568,N_7671);
xnor U8267 (N_8267,N_7502,N_8210);
nand U8268 (N_8268,N_7664,N_7991);
nand U8269 (N_8269,N_8174,N_7793);
and U8270 (N_8270,N_7970,N_7769);
nand U8271 (N_8271,N_8000,N_8061);
nand U8272 (N_8272,N_8068,N_7698);
nor U8273 (N_8273,N_7944,N_7534);
and U8274 (N_8274,N_7950,N_8069);
nand U8275 (N_8275,N_8045,N_7724);
nor U8276 (N_8276,N_7570,N_7853);
or U8277 (N_8277,N_8186,N_7747);
nor U8278 (N_8278,N_8176,N_7906);
and U8279 (N_8279,N_7736,N_8107);
xnor U8280 (N_8280,N_7865,N_7990);
xor U8281 (N_8281,N_7799,N_7764);
or U8282 (N_8282,N_7501,N_8226);
and U8283 (N_8283,N_7946,N_7598);
and U8284 (N_8284,N_8046,N_7784);
nand U8285 (N_8285,N_7655,N_7558);
or U8286 (N_8286,N_8077,N_8052);
and U8287 (N_8287,N_7533,N_7789);
nand U8288 (N_8288,N_8131,N_8175);
and U8289 (N_8289,N_8221,N_7994);
or U8290 (N_8290,N_7509,N_8106);
and U8291 (N_8291,N_8031,N_7927);
or U8292 (N_8292,N_7934,N_7776);
and U8293 (N_8293,N_7752,N_7914);
nor U8294 (N_8294,N_7549,N_7707);
nand U8295 (N_8295,N_8218,N_7722);
and U8296 (N_8296,N_8017,N_7965);
nand U8297 (N_8297,N_7762,N_8246);
xnor U8298 (N_8298,N_7713,N_7755);
nand U8299 (N_8299,N_8240,N_7840);
xor U8300 (N_8300,N_7739,N_8161);
nor U8301 (N_8301,N_8148,N_7567);
nor U8302 (N_8302,N_7624,N_8130);
nor U8303 (N_8303,N_8132,N_7938);
nor U8304 (N_8304,N_7611,N_7908);
nor U8305 (N_8305,N_7852,N_8105);
and U8306 (N_8306,N_7977,N_8116);
nor U8307 (N_8307,N_7667,N_7975);
nor U8308 (N_8308,N_8147,N_8158);
nor U8309 (N_8309,N_8173,N_8047);
nand U8310 (N_8310,N_8229,N_7876);
nand U8311 (N_8311,N_8187,N_7948);
nor U8312 (N_8312,N_7580,N_8193);
and U8313 (N_8313,N_7910,N_7719);
nor U8314 (N_8314,N_7550,N_7911);
or U8315 (N_8315,N_8050,N_7896);
and U8316 (N_8316,N_7727,N_8238);
and U8317 (N_8317,N_8108,N_8171);
or U8318 (N_8318,N_7937,N_7610);
nor U8319 (N_8319,N_8248,N_7553);
nor U8320 (N_8320,N_7602,N_8160);
nor U8321 (N_8321,N_7826,N_7618);
and U8322 (N_8322,N_7929,N_7642);
nand U8323 (N_8323,N_7895,N_7877);
and U8324 (N_8324,N_7725,N_7861);
xor U8325 (N_8325,N_7710,N_7781);
xor U8326 (N_8326,N_8201,N_7925);
or U8327 (N_8327,N_7639,N_8112);
or U8328 (N_8328,N_7662,N_7621);
or U8329 (N_8329,N_8236,N_8121);
and U8330 (N_8330,N_7585,N_8137);
nor U8331 (N_8331,N_7582,N_7772);
and U8332 (N_8332,N_8249,N_8198);
or U8333 (N_8333,N_8022,N_8033);
or U8334 (N_8334,N_8208,N_8037);
nor U8335 (N_8335,N_8007,N_7632);
or U8336 (N_8336,N_7613,N_7750);
xor U8337 (N_8337,N_7548,N_7716);
xnor U8338 (N_8338,N_7775,N_7694);
nand U8339 (N_8339,N_8034,N_8135);
xor U8340 (N_8340,N_8205,N_8183);
nor U8341 (N_8341,N_8111,N_7993);
and U8342 (N_8342,N_7633,N_8247);
xor U8343 (N_8343,N_7731,N_8170);
xor U8344 (N_8344,N_7907,N_7751);
or U8345 (N_8345,N_7783,N_7891);
and U8346 (N_8346,N_8098,N_7997);
nand U8347 (N_8347,N_8202,N_8097);
or U8348 (N_8348,N_7732,N_8220);
and U8349 (N_8349,N_7643,N_7590);
xnor U8350 (N_8350,N_8189,N_8060);
nand U8351 (N_8351,N_7500,N_8152);
and U8352 (N_8352,N_7924,N_7849);
and U8353 (N_8353,N_7868,N_8102);
nand U8354 (N_8354,N_7601,N_7768);
nor U8355 (N_8355,N_7996,N_7654);
nor U8356 (N_8356,N_7708,N_7972);
or U8357 (N_8357,N_7503,N_7960);
or U8358 (N_8358,N_7734,N_7545);
and U8359 (N_8359,N_7957,N_7803);
and U8360 (N_8360,N_8036,N_7804);
nand U8361 (N_8361,N_7663,N_8009);
and U8362 (N_8362,N_7827,N_8087);
xor U8363 (N_8363,N_7814,N_7984);
nand U8364 (N_8364,N_8213,N_7626);
nand U8365 (N_8365,N_8043,N_7519);
nand U8366 (N_8366,N_7536,N_7697);
or U8367 (N_8367,N_7717,N_8223);
or U8368 (N_8368,N_7761,N_8092);
nor U8369 (N_8369,N_7525,N_7980);
and U8370 (N_8370,N_7850,N_7763);
and U8371 (N_8371,N_7941,N_7588);
or U8372 (N_8372,N_7976,N_8203);
nand U8373 (N_8373,N_7528,N_7607);
nor U8374 (N_8374,N_8197,N_7681);
and U8375 (N_8375,N_8056,N_7730);
or U8376 (N_8376,N_7967,N_7933);
nand U8377 (N_8377,N_8094,N_8237);
nor U8378 (N_8378,N_7586,N_7506);
nor U8379 (N_8379,N_7843,N_7848);
or U8380 (N_8380,N_7873,N_8192);
and U8381 (N_8381,N_7640,N_7516);
nand U8382 (N_8382,N_7635,N_7617);
or U8383 (N_8383,N_8081,N_7985);
nor U8384 (N_8384,N_7883,N_7879);
nor U8385 (N_8385,N_7634,N_7801);
and U8386 (N_8386,N_7958,N_7530);
nand U8387 (N_8387,N_8071,N_7987);
or U8388 (N_8388,N_8101,N_7741);
or U8389 (N_8389,N_7859,N_7754);
xnor U8390 (N_8390,N_8028,N_7954);
nand U8391 (N_8391,N_8181,N_7882);
and U8392 (N_8392,N_7936,N_7524);
or U8393 (N_8393,N_7847,N_7505);
or U8394 (N_8394,N_8195,N_7805);
nor U8395 (N_8395,N_7718,N_8078);
and U8396 (N_8396,N_7543,N_8206);
and U8397 (N_8397,N_7862,N_7532);
and U8398 (N_8398,N_7964,N_8066);
nand U8399 (N_8399,N_7504,N_7949);
or U8400 (N_8400,N_8038,N_7904);
nor U8401 (N_8401,N_7627,N_7572);
or U8402 (N_8402,N_7540,N_7599);
nand U8403 (N_8403,N_7696,N_8011);
and U8404 (N_8404,N_7675,N_7798);
or U8405 (N_8405,N_7546,N_7899);
nand U8406 (N_8406,N_8041,N_7616);
xor U8407 (N_8407,N_7945,N_7609);
nand U8408 (N_8408,N_7756,N_7592);
nor U8409 (N_8409,N_7542,N_8055);
or U8410 (N_8410,N_7661,N_7705);
and U8411 (N_8411,N_7955,N_7777);
and U8412 (N_8412,N_7584,N_7813);
nor U8413 (N_8413,N_7575,N_7678);
or U8414 (N_8414,N_8233,N_7918);
or U8415 (N_8415,N_7641,N_7935);
nand U8416 (N_8416,N_7875,N_7828);
xnor U8417 (N_8417,N_7728,N_8190);
xor U8418 (N_8418,N_8244,N_8134);
and U8419 (N_8419,N_8180,N_7554);
and U8420 (N_8420,N_7983,N_8010);
xnor U8421 (N_8421,N_7759,N_8110);
nand U8422 (N_8422,N_7988,N_8128);
nor U8423 (N_8423,N_7952,N_7951);
nand U8424 (N_8424,N_8209,N_7704);
and U8425 (N_8425,N_7645,N_7874);
and U8426 (N_8426,N_7737,N_7846);
nand U8427 (N_8427,N_8235,N_7680);
and U8428 (N_8428,N_7650,N_8004);
or U8429 (N_8429,N_7529,N_7531);
nand U8430 (N_8430,N_7878,N_7829);
and U8431 (N_8431,N_7887,N_7552);
or U8432 (N_8432,N_8090,N_8120);
and U8433 (N_8433,N_8225,N_7712);
and U8434 (N_8434,N_7742,N_7686);
xor U8435 (N_8435,N_7526,N_7773);
nand U8436 (N_8436,N_8124,N_7884);
and U8437 (N_8437,N_8199,N_8172);
or U8438 (N_8438,N_7581,N_7587);
and U8439 (N_8439,N_8228,N_7864);
nor U8440 (N_8440,N_8005,N_7766);
and U8441 (N_8441,N_7919,N_8100);
nand U8442 (N_8442,N_8224,N_8242);
xnor U8443 (N_8443,N_7721,N_8014);
or U8444 (N_8444,N_7715,N_7792);
xor U8445 (N_8445,N_8217,N_7872);
or U8446 (N_8446,N_8065,N_8138);
and U8447 (N_8447,N_7981,N_7903);
nor U8448 (N_8448,N_7982,N_8035);
or U8449 (N_8449,N_7810,N_8018);
nand U8450 (N_8450,N_7902,N_7668);
nand U8451 (N_8451,N_7820,N_8048);
or U8452 (N_8452,N_8003,N_7656);
nor U8453 (N_8453,N_7753,N_7893);
nand U8454 (N_8454,N_7699,N_8200);
or U8455 (N_8455,N_7646,N_7782);
and U8456 (N_8456,N_7596,N_7961);
or U8457 (N_8457,N_7749,N_7744);
or U8458 (N_8458,N_7870,N_7867);
nand U8459 (N_8459,N_7513,N_8157);
nor U8460 (N_8460,N_7815,N_8089);
or U8461 (N_8461,N_7854,N_7771);
or U8462 (N_8462,N_7839,N_7669);
and U8463 (N_8463,N_7905,N_7931);
nor U8464 (N_8464,N_7703,N_7579);
nand U8465 (N_8465,N_7557,N_7986);
and U8466 (N_8466,N_7787,N_7807);
and U8467 (N_8467,N_8150,N_8133);
xor U8468 (N_8468,N_8093,N_8178);
or U8469 (N_8469,N_7665,N_7569);
or U8470 (N_8470,N_7830,N_8168);
or U8471 (N_8471,N_7962,N_8070);
xor U8472 (N_8472,N_7956,N_7690);
nand U8473 (N_8473,N_8136,N_8044);
nand U8474 (N_8474,N_8049,N_7600);
and U8475 (N_8475,N_7748,N_7559);
or U8476 (N_8476,N_7816,N_8064);
and U8477 (N_8477,N_7556,N_7998);
nor U8478 (N_8478,N_8164,N_7808);
and U8479 (N_8479,N_8013,N_7825);
and U8480 (N_8480,N_7615,N_7648);
nor U8481 (N_8481,N_7726,N_7989);
nand U8482 (N_8482,N_8146,N_7628);
or U8483 (N_8483,N_8002,N_8227);
or U8484 (N_8484,N_8230,N_7841);
xor U8485 (N_8485,N_7894,N_8154);
and U8486 (N_8486,N_8119,N_8159);
or U8487 (N_8487,N_7890,N_7880);
or U8488 (N_8488,N_7760,N_7818);
nor U8489 (N_8489,N_7765,N_7822);
or U8490 (N_8490,N_7966,N_7562);
and U8491 (N_8491,N_8073,N_7738);
and U8492 (N_8492,N_7591,N_7677);
and U8493 (N_8493,N_7711,N_7855);
nand U8494 (N_8494,N_7940,N_7670);
and U8495 (N_8495,N_7687,N_7623);
nor U8496 (N_8496,N_8169,N_7969);
nor U8497 (N_8497,N_7638,N_7537);
xor U8498 (N_8498,N_8058,N_7625);
or U8499 (N_8499,N_7885,N_7780);
xor U8500 (N_8500,N_7566,N_8001);
nand U8501 (N_8501,N_7794,N_7811);
nor U8502 (N_8502,N_8075,N_7953);
nor U8503 (N_8503,N_7920,N_8109);
or U8504 (N_8504,N_8232,N_8129);
nor U8505 (N_8505,N_7563,N_7620);
and U8506 (N_8506,N_7791,N_7963);
nor U8507 (N_8507,N_7743,N_7833);
or U8508 (N_8508,N_7909,N_8072);
nor U8509 (N_8509,N_8062,N_8162);
or U8510 (N_8510,N_7603,N_7578);
xnor U8511 (N_8511,N_7682,N_7923);
and U8512 (N_8512,N_7900,N_8207);
nor U8513 (N_8513,N_8113,N_7788);
nor U8514 (N_8514,N_8096,N_8239);
or U8515 (N_8515,N_8204,N_7832);
and U8516 (N_8516,N_8079,N_8245);
nand U8517 (N_8517,N_8088,N_7800);
nand U8518 (N_8518,N_7709,N_7604);
nand U8519 (N_8519,N_7614,N_8163);
or U8520 (N_8520,N_8053,N_8179);
nor U8521 (N_8521,N_8219,N_7812);
or U8522 (N_8522,N_7922,N_7672);
and U8523 (N_8523,N_7658,N_7720);
and U8524 (N_8524,N_8015,N_8012);
nor U8525 (N_8525,N_7683,N_7644);
xor U8526 (N_8526,N_7915,N_8243);
and U8527 (N_8527,N_7897,N_7995);
nor U8528 (N_8528,N_8241,N_7851);
nor U8529 (N_8529,N_7688,N_8184);
and U8530 (N_8530,N_7770,N_8188);
nand U8531 (N_8531,N_7706,N_7856);
or U8532 (N_8532,N_7871,N_7845);
and U8533 (N_8533,N_8051,N_7571);
or U8534 (N_8534,N_7866,N_7676);
nor U8535 (N_8535,N_7651,N_8222);
nor U8536 (N_8536,N_7999,N_7838);
and U8537 (N_8537,N_7573,N_7521);
or U8538 (N_8538,N_7745,N_7913);
or U8539 (N_8539,N_8006,N_7551);
xnor U8540 (N_8540,N_7973,N_7774);
nand U8541 (N_8541,N_7576,N_8085);
and U8542 (N_8542,N_7606,N_7930);
nor U8543 (N_8543,N_7510,N_7916);
or U8544 (N_8544,N_7595,N_7653);
and U8545 (N_8545,N_7535,N_7943);
nor U8546 (N_8546,N_7637,N_7857);
nand U8547 (N_8547,N_8076,N_8143);
or U8548 (N_8548,N_8084,N_8196);
and U8549 (N_8549,N_7979,N_7888);
nor U8550 (N_8550,N_7881,N_7947);
or U8551 (N_8551,N_8145,N_8234);
and U8552 (N_8552,N_8086,N_7858);
xnor U8553 (N_8553,N_8095,N_7608);
xnor U8554 (N_8554,N_7869,N_8099);
nor U8555 (N_8555,N_7844,N_7657);
nand U8556 (N_8556,N_7834,N_7842);
nand U8557 (N_8557,N_7836,N_8074);
and U8558 (N_8558,N_7837,N_8040);
nor U8559 (N_8559,N_8216,N_8117);
or U8560 (N_8560,N_8114,N_7589);
or U8561 (N_8561,N_7939,N_8125);
nor U8562 (N_8562,N_8021,N_8167);
nor U8563 (N_8563,N_8083,N_8019);
and U8564 (N_8564,N_7527,N_7898);
or U8565 (N_8565,N_8182,N_8020);
or U8566 (N_8566,N_8042,N_7819);
and U8567 (N_8567,N_8215,N_7740);
or U8568 (N_8568,N_8177,N_7806);
or U8569 (N_8569,N_8067,N_7515);
and U8570 (N_8570,N_7729,N_7522);
nor U8571 (N_8571,N_8016,N_7823);
nor U8572 (N_8572,N_7565,N_7652);
and U8573 (N_8573,N_8032,N_7802);
and U8574 (N_8574,N_7631,N_7647);
and U8575 (N_8575,N_7863,N_7917);
nor U8576 (N_8576,N_7673,N_7779);
or U8577 (N_8577,N_8025,N_7786);
or U8578 (N_8578,N_7860,N_8057);
and U8579 (N_8579,N_7689,N_7577);
or U8580 (N_8580,N_7912,N_8008);
nand U8581 (N_8581,N_7701,N_7636);
or U8582 (N_8582,N_7758,N_7520);
nor U8583 (N_8583,N_7649,N_8185);
nor U8584 (N_8584,N_7630,N_8026);
or U8585 (N_8585,N_7512,N_8194);
and U8586 (N_8586,N_7959,N_8059);
and U8587 (N_8587,N_7928,N_8126);
or U8588 (N_8588,N_7583,N_7889);
or U8589 (N_8589,N_7785,N_8156);
and U8590 (N_8590,N_7835,N_7619);
nor U8591 (N_8591,N_8211,N_7790);
nor U8592 (N_8592,N_8153,N_8231);
and U8593 (N_8593,N_7605,N_7555);
and U8594 (N_8594,N_7968,N_8141);
or U8595 (N_8595,N_7901,N_7735);
or U8596 (N_8596,N_7538,N_7932);
and U8597 (N_8597,N_7511,N_8115);
nor U8598 (N_8598,N_7560,N_7561);
and U8599 (N_8599,N_7622,N_8104);
and U8600 (N_8600,N_7679,N_8030);
nand U8601 (N_8601,N_7593,N_7978);
nor U8602 (N_8602,N_7817,N_8024);
and U8603 (N_8603,N_7597,N_8127);
or U8604 (N_8604,N_7886,N_8080);
nand U8605 (N_8605,N_7693,N_7992);
or U8606 (N_8606,N_8212,N_7659);
nor U8607 (N_8607,N_8123,N_7541);
nand U8608 (N_8608,N_8091,N_7757);
nor U8609 (N_8609,N_7700,N_7702);
nand U8610 (N_8610,N_7795,N_7547);
and U8611 (N_8611,N_7831,N_8063);
or U8612 (N_8612,N_8140,N_8027);
nor U8613 (N_8613,N_7733,N_7508);
and U8614 (N_8614,N_8214,N_8082);
and U8615 (N_8615,N_7809,N_7574);
and U8616 (N_8616,N_7714,N_8155);
and U8617 (N_8617,N_7518,N_7695);
nor U8618 (N_8618,N_7564,N_7971);
nand U8619 (N_8619,N_8142,N_7692);
nand U8620 (N_8620,N_8149,N_8103);
and U8621 (N_8621,N_7660,N_7507);
nand U8622 (N_8622,N_7892,N_7723);
xor U8623 (N_8623,N_8165,N_7767);
and U8624 (N_8624,N_8118,N_8191);
or U8625 (N_8625,N_7915,N_8206);
xnor U8626 (N_8626,N_8155,N_7837);
and U8627 (N_8627,N_7583,N_7840);
nor U8628 (N_8628,N_7992,N_7969);
and U8629 (N_8629,N_7769,N_7501);
and U8630 (N_8630,N_7663,N_7603);
and U8631 (N_8631,N_7722,N_8126);
and U8632 (N_8632,N_8111,N_7893);
nand U8633 (N_8633,N_8102,N_7508);
or U8634 (N_8634,N_7851,N_7858);
and U8635 (N_8635,N_7503,N_7716);
or U8636 (N_8636,N_8106,N_7924);
nand U8637 (N_8637,N_8075,N_7927);
and U8638 (N_8638,N_8174,N_8099);
or U8639 (N_8639,N_7856,N_8078);
nand U8640 (N_8640,N_7944,N_8182);
nand U8641 (N_8641,N_8147,N_7559);
nor U8642 (N_8642,N_7801,N_7707);
xnor U8643 (N_8643,N_7784,N_8091);
and U8644 (N_8644,N_7727,N_8048);
or U8645 (N_8645,N_8108,N_7976);
nor U8646 (N_8646,N_7707,N_8138);
and U8647 (N_8647,N_7600,N_8233);
nor U8648 (N_8648,N_8106,N_7796);
and U8649 (N_8649,N_7706,N_8178);
nand U8650 (N_8650,N_7653,N_7890);
or U8651 (N_8651,N_7518,N_7953);
xor U8652 (N_8652,N_8120,N_8175);
or U8653 (N_8653,N_8220,N_7972);
or U8654 (N_8654,N_8057,N_7668);
or U8655 (N_8655,N_7901,N_7836);
nor U8656 (N_8656,N_7760,N_7687);
nor U8657 (N_8657,N_8035,N_7768);
and U8658 (N_8658,N_7840,N_8106);
nand U8659 (N_8659,N_8200,N_7764);
nand U8660 (N_8660,N_8020,N_7755);
and U8661 (N_8661,N_8118,N_8210);
nor U8662 (N_8662,N_7974,N_7732);
nand U8663 (N_8663,N_8248,N_7902);
nand U8664 (N_8664,N_7505,N_7943);
and U8665 (N_8665,N_8234,N_7808);
xnor U8666 (N_8666,N_8160,N_7685);
nor U8667 (N_8667,N_7670,N_7772);
nor U8668 (N_8668,N_8025,N_7692);
nand U8669 (N_8669,N_8213,N_7802);
xnor U8670 (N_8670,N_7633,N_8232);
nor U8671 (N_8671,N_7561,N_7680);
nor U8672 (N_8672,N_7574,N_7620);
nand U8673 (N_8673,N_8032,N_7522);
and U8674 (N_8674,N_8029,N_7798);
xnor U8675 (N_8675,N_7543,N_7560);
xor U8676 (N_8676,N_7945,N_8139);
nor U8677 (N_8677,N_7816,N_8168);
or U8678 (N_8678,N_7598,N_7803);
nand U8679 (N_8679,N_7834,N_7677);
or U8680 (N_8680,N_7827,N_7554);
nor U8681 (N_8681,N_8098,N_7700);
and U8682 (N_8682,N_7964,N_8125);
and U8683 (N_8683,N_7958,N_7933);
and U8684 (N_8684,N_7626,N_7894);
and U8685 (N_8685,N_8209,N_8092);
or U8686 (N_8686,N_8141,N_7784);
or U8687 (N_8687,N_7931,N_7895);
nor U8688 (N_8688,N_7806,N_7634);
nand U8689 (N_8689,N_8125,N_7805);
xnor U8690 (N_8690,N_7546,N_7878);
nor U8691 (N_8691,N_8211,N_7993);
xnor U8692 (N_8692,N_8172,N_7941);
nand U8693 (N_8693,N_7927,N_7663);
nand U8694 (N_8694,N_7926,N_8130);
or U8695 (N_8695,N_7635,N_8035);
nand U8696 (N_8696,N_7531,N_7889);
or U8697 (N_8697,N_8154,N_7717);
xor U8698 (N_8698,N_8132,N_7513);
and U8699 (N_8699,N_7660,N_7610);
nor U8700 (N_8700,N_7953,N_8115);
nor U8701 (N_8701,N_8212,N_7606);
xor U8702 (N_8702,N_7974,N_7533);
xnor U8703 (N_8703,N_7935,N_7787);
nor U8704 (N_8704,N_7919,N_7660);
nor U8705 (N_8705,N_7793,N_7978);
nand U8706 (N_8706,N_7891,N_7809);
nor U8707 (N_8707,N_7713,N_8185);
and U8708 (N_8708,N_8080,N_8023);
nor U8709 (N_8709,N_7803,N_7790);
and U8710 (N_8710,N_7747,N_7576);
nor U8711 (N_8711,N_7685,N_7683);
and U8712 (N_8712,N_7625,N_7616);
and U8713 (N_8713,N_7827,N_7768);
nor U8714 (N_8714,N_7934,N_7553);
or U8715 (N_8715,N_7656,N_7565);
nand U8716 (N_8716,N_7618,N_7523);
or U8717 (N_8717,N_7728,N_7832);
and U8718 (N_8718,N_7844,N_8208);
nand U8719 (N_8719,N_8012,N_7623);
and U8720 (N_8720,N_8000,N_7531);
and U8721 (N_8721,N_7596,N_7774);
nor U8722 (N_8722,N_8048,N_7598);
nand U8723 (N_8723,N_8106,N_8158);
or U8724 (N_8724,N_7996,N_8209);
nor U8725 (N_8725,N_8149,N_7770);
and U8726 (N_8726,N_7692,N_8225);
or U8727 (N_8727,N_7864,N_7617);
and U8728 (N_8728,N_7586,N_7814);
nand U8729 (N_8729,N_7552,N_7632);
and U8730 (N_8730,N_7702,N_8209);
nor U8731 (N_8731,N_8091,N_8190);
or U8732 (N_8732,N_7562,N_7769);
nand U8733 (N_8733,N_7869,N_7884);
and U8734 (N_8734,N_7989,N_8125);
or U8735 (N_8735,N_7502,N_8078);
or U8736 (N_8736,N_7646,N_7549);
nand U8737 (N_8737,N_8172,N_7643);
and U8738 (N_8738,N_8045,N_7977);
nor U8739 (N_8739,N_7739,N_7928);
or U8740 (N_8740,N_7510,N_7602);
nand U8741 (N_8741,N_8017,N_8222);
and U8742 (N_8742,N_8241,N_7505);
nand U8743 (N_8743,N_7705,N_7749);
nor U8744 (N_8744,N_7953,N_7982);
or U8745 (N_8745,N_7686,N_7794);
xor U8746 (N_8746,N_7725,N_7631);
or U8747 (N_8747,N_7740,N_8164);
or U8748 (N_8748,N_8220,N_7787);
or U8749 (N_8749,N_7876,N_8207);
nor U8750 (N_8750,N_7688,N_7887);
nand U8751 (N_8751,N_7944,N_7516);
nand U8752 (N_8752,N_7545,N_8102);
and U8753 (N_8753,N_8011,N_7942);
nand U8754 (N_8754,N_8048,N_7953);
nor U8755 (N_8755,N_8012,N_8061);
or U8756 (N_8756,N_7688,N_8025);
nor U8757 (N_8757,N_7594,N_8213);
and U8758 (N_8758,N_7856,N_7854);
nor U8759 (N_8759,N_8166,N_8239);
nand U8760 (N_8760,N_8058,N_8155);
nand U8761 (N_8761,N_7670,N_8200);
nand U8762 (N_8762,N_7835,N_7768);
and U8763 (N_8763,N_8033,N_8134);
nand U8764 (N_8764,N_7505,N_7810);
nand U8765 (N_8765,N_7589,N_8159);
and U8766 (N_8766,N_8075,N_7783);
nor U8767 (N_8767,N_8201,N_7830);
nand U8768 (N_8768,N_8061,N_8084);
nor U8769 (N_8769,N_7746,N_7918);
nor U8770 (N_8770,N_7993,N_8165);
or U8771 (N_8771,N_7631,N_8135);
or U8772 (N_8772,N_7598,N_7638);
xnor U8773 (N_8773,N_7930,N_7993);
nand U8774 (N_8774,N_8123,N_7924);
nand U8775 (N_8775,N_8084,N_7681);
nand U8776 (N_8776,N_7718,N_8187);
nand U8777 (N_8777,N_8001,N_7972);
nand U8778 (N_8778,N_7756,N_7558);
or U8779 (N_8779,N_7532,N_7799);
nor U8780 (N_8780,N_7902,N_7726);
nand U8781 (N_8781,N_7794,N_8132);
nor U8782 (N_8782,N_7878,N_8039);
nand U8783 (N_8783,N_7687,N_8008);
and U8784 (N_8784,N_7822,N_7965);
nand U8785 (N_8785,N_7728,N_7646);
or U8786 (N_8786,N_7949,N_7545);
nand U8787 (N_8787,N_7865,N_7932);
or U8788 (N_8788,N_8198,N_7951);
nand U8789 (N_8789,N_7680,N_7594);
nor U8790 (N_8790,N_8006,N_7606);
and U8791 (N_8791,N_8154,N_8012);
nor U8792 (N_8792,N_8201,N_7970);
or U8793 (N_8793,N_8158,N_8175);
and U8794 (N_8794,N_8140,N_8105);
nand U8795 (N_8795,N_7797,N_7800);
nand U8796 (N_8796,N_7706,N_8080);
and U8797 (N_8797,N_7626,N_7909);
or U8798 (N_8798,N_8098,N_7978);
and U8799 (N_8799,N_7977,N_7837);
nor U8800 (N_8800,N_8181,N_7810);
or U8801 (N_8801,N_8079,N_7667);
or U8802 (N_8802,N_7828,N_7692);
nor U8803 (N_8803,N_7821,N_7539);
xor U8804 (N_8804,N_7967,N_7719);
or U8805 (N_8805,N_8166,N_7524);
nand U8806 (N_8806,N_8157,N_7579);
nor U8807 (N_8807,N_7886,N_7612);
and U8808 (N_8808,N_7642,N_8111);
nor U8809 (N_8809,N_7692,N_7628);
nor U8810 (N_8810,N_8088,N_7720);
or U8811 (N_8811,N_7835,N_8039);
or U8812 (N_8812,N_8003,N_7774);
nand U8813 (N_8813,N_8240,N_8221);
xnor U8814 (N_8814,N_7720,N_8233);
nor U8815 (N_8815,N_7836,N_7861);
nor U8816 (N_8816,N_8018,N_8055);
and U8817 (N_8817,N_7860,N_7547);
and U8818 (N_8818,N_7533,N_7897);
nor U8819 (N_8819,N_8240,N_8238);
xor U8820 (N_8820,N_8185,N_7554);
nand U8821 (N_8821,N_7813,N_7860);
or U8822 (N_8822,N_8155,N_7797);
nor U8823 (N_8823,N_8189,N_7995);
and U8824 (N_8824,N_8098,N_8229);
xor U8825 (N_8825,N_8043,N_7728);
and U8826 (N_8826,N_8006,N_8178);
or U8827 (N_8827,N_7631,N_7621);
nor U8828 (N_8828,N_7606,N_7514);
or U8829 (N_8829,N_7574,N_7682);
xnor U8830 (N_8830,N_7982,N_8057);
and U8831 (N_8831,N_7787,N_7665);
nand U8832 (N_8832,N_7802,N_8139);
nand U8833 (N_8833,N_8176,N_7735);
or U8834 (N_8834,N_7751,N_7586);
nand U8835 (N_8835,N_8161,N_8102);
nor U8836 (N_8836,N_8020,N_7575);
nand U8837 (N_8837,N_8224,N_7802);
nand U8838 (N_8838,N_8109,N_7941);
nand U8839 (N_8839,N_7845,N_8136);
and U8840 (N_8840,N_7693,N_8235);
nand U8841 (N_8841,N_7858,N_7890);
nand U8842 (N_8842,N_7964,N_7635);
nand U8843 (N_8843,N_8134,N_7553);
and U8844 (N_8844,N_7985,N_7560);
or U8845 (N_8845,N_7822,N_7823);
xor U8846 (N_8846,N_7710,N_7813);
or U8847 (N_8847,N_7915,N_7710);
nor U8848 (N_8848,N_7626,N_7818);
and U8849 (N_8849,N_8063,N_7973);
nand U8850 (N_8850,N_7799,N_7930);
or U8851 (N_8851,N_8177,N_8078);
xnor U8852 (N_8852,N_7750,N_7695);
or U8853 (N_8853,N_7578,N_8226);
and U8854 (N_8854,N_7656,N_8026);
nor U8855 (N_8855,N_7955,N_7603);
or U8856 (N_8856,N_7676,N_7656);
nor U8857 (N_8857,N_7957,N_8068);
and U8858 (N_8858,N_8127,N_8009);
and U8859 (N_8859,N_7930,N_8167);
nand U8860 (N_8860,N_7688,N_8093);
xor U8861 (N_8861,N_7506,N_7948);
and U8862 (N_8862,N_8103,N_7764);
or U8863 (N_8863,N_8011,N_8053);
nand U8864 (N_8864,N_7968,N_8088);
or U8865 (N_8865,N_8132,N_8194);
and U8866 (N_8866,N_7501,N_7742);
or U8867 (N_8867,N_7584,N_8165);
xnor U8868 (N_8868,N_8171,N_7796);
or U8869 (N_8869,N_7651,N_8183);
xnor U8870 (N_8870,N_8010,N_7669);
nand U8871 (N_8871,N_8215,N_7882);
and U8872 (N_8872,N_7539,N_7646);
nor U8873 (N_8873,N_7994,N_8116);
or U8874 (N_8874,N_7634,N_7568);
nand U8875 (N_8875,N_7904,N_7561);
and U8876 (N_8876,N_8130,N_7606);
nand U8877 (N_8877,N_8112,N_7601);
and U8878 (N_8878,N_8098,N_7643);
nand U8879 (N_8879,N_7916,N_7951);
nand U8880 (N_8880,N_7546,N_7996);
or U8881 (N_8881,N_8169,N_7994);
and U8882 (N_8882,N_8128,N_7628);
nand U8883 (N_8883,N_8090,N_7549);
or U8884 (N_8884,N_7863,N_7878);
nor U8885 (N_8885,N_8154,N_8075);
and U8886 (N_8886,N_7545,N_8009);
nor U8887 (N_8887,N_8222,N_7533);
and U8888 (N_8888,N_7715,N_8181);
xnor U8889 (N_8889,N_8192,N_7629);
nor U8890 (N_8890,N_7541,N_7900);
and U8891 (N_8891,N_7890,N_8023);
nand U8892 (N_8892,N_8116,N_8175);
or U8893 (N_8893,N_7623,N_8199);
nand U8894 (N_8894,N_7961,N_7537);
nor U8895 (N_8895,N_8216,N_7798);
and U8896 (N_8896,N_7699,N_8121);
or U8897 (N_8897,N_8133,N_7957);
xnor U8898 (N_8898,N_7914,N_7854);
or U8899 (N_8899,N_7633,N_8025);
xnor U8900 (N_8900,N_7531,N_7913);
nand U8901 (N_8901,N_7737,N_8089);
nor U8902 (N_8902,N_7942,N_8116);
and U8903 (N_8903,N_8055,N_7910);
xnor U8904 (N_8904,N_8011,N_7655);
nor U8905 (N_8905,N_8023,N_7910);
or U8906 (N_8906,N_8068,N_7912);
or U8907 (N_8907,N_7544,N_8105);
and U8908 (N_8908,N_7833,N_7531);
nor U8909 (N_8909,N_8065,N_7690);
xnor U8910 (N_8910,N_7706,N_8005);
nand U8911 (N_8911,N_7688,N_8018);
nand U8912 (N_8912,N_8071,N_8068);
and U8913 (N_8913,N_7886,N_7671);
and U8914 (N_8914,N_7954,N_8011);
nor U8915 (N_8915,N_8121,N_7698);
or U8916 (N_8916,N_7755,N_7571);
or U8917 (N_8917,N_8241,N_7987);
and U8918 (N_8918,N_7796,N_7701);
nor U8919 (N_8919,N_7883,N_7880);
or U8920 (N_8920,N_8123,N_8168);
or U8921 (N_8921,N_7803,N_7521);
and U8922 (N_8922,N_7704,N_8141);
or U8923 (N_8923,N_7959,N_7746);
and U8924 (N_8924,N_8188,N_7707);
nand U8925 (N_8925,N_7706,N_7808);
and U8926 (N_8926,N_7641,N_7561);
and U8927 (N_8927,N_7708,N_7867);
and U8928 (N_8928,N_7526,N_7606);
nand U8929 (N_8929,N_7767,N_7895);
nor U8930 (N_8930,N_7572,N_7754);
nor U8931 (N_8931,N_8189,N_7665);
nor U8932 (N_8932,N_7957,N_7551);
or U8933 (N_8933,N_7629,N_7801);
or U8934 (N_8934,N_7921,N_8151);
xnor U8935 (N_8935,N_7824,N_8039);
nand U8936 (N_8936,N_7623,N_8121);
nor U8937 (N_8937,N_7858,N_7771);
nand U8938 (N_8938,N_8030,N_7571);
nor U8939 (N_8939,N_7541,N_8167);
or U8940 (N_8940,N_7686,N_7831);
or U8941 (N_8941,N_7930,N_8115);
xnor U8942 (N_8942,N_7659,N_8078);
nand U8943 (N_8943,N_7633,N_7641);
and U8944 (N_8944,N_7663,N_7787);
or U8945 (N_8945,N_7627,N_7646);
nand U8946 (N_8946,N_7850,N_7852);
or U8947 (N_8947,N_7830,N_7591);
and U8948 (N_8948,N_7849,N_7788);
nor U8949 (N_8949,N_7584,N_7784);
or U8950 (N_8950,N_7643,N_7826);
nor U8951 (N_8951,N_7568,N_7843);
nor U8952 (N_8952,N_8154,N_7965);
nand U8953 (N_8953,N_7959,N_8184);
xor U8954 (N_8954,N_8225,N_8067);
and U8955 (N_8955,N_7639,N_7564);
nor U8956 (N_8956,N_7876,N_7655);
nand U8957 (N_8957,N_8188,N_7931);
nor U8958 (N_8958,N_7522,N_7539);
nor U8959 (N_8959,N_7970,N_7894);
nor U8960 (N_8960,N_7849,N_7870);
or U8961 (N_8961,N_7580,N_8050);
or U8962 (N_8962,N_7837,N_7793);
nor U8963 (N_8963,N_7923,N_8071);
or U8964 (N_8964,N_7506,N_7566);
and U8965 (N_8965,N_7770,N_7981);
xnor U8966 (N_8966,N_7831,N_7504);
xor U8967 (N_8967,N_7758,N_8091);
nor U8968 (N_8968,N_7764,N_7596);
nand U8969 (N_8969,N_8163,N_8111);
or U8970 (N_8970,N_8069,N_8108);
nor U8971 (N_8971,N_7512,N_7866);
nor U8972 (N_8972,N_8004,N_7800);
nand U8973 (N_8973,N_7725,N_7502);
nor U8974 (N_8974,N_7882,N_8039);
or U8975 (N_8975,N_7962,N_7749);
nand U8976 (N_8976,N_8186,N_7515);
nor U8977 (N_8977,N_7703,N_8118);
nor U8978 (N_8978,N_7926,N_8091);
and U8979 (N_8979,N_7634,N_7841);
and U8980 (N_8980,N_8048,N_7634);
and U8981 (N_8981,N_7885,N_7935);
nor U8982 (N_8982,N_8189,N_8061);
nand U8983 (N_8983,N_8050,N_7922);
and U8984 (N_8984,N_7671,N_7798);
nand U8985 (N_8985,N_7502,N_7579);
or U8986 (N_8986,N_8012,N_8038);
and U8987 (N_8987,N_7506,N_8192);
or U8988 (N_8988,N_7558,N_7521);
nand U8989 (N_8989,N_7543,N_8230);
xor U8990 (N_8990,N_8068,N_8044);
nor U8991 (N_8991,N_8043,N_7905);
xnor U8992 (N_8992,N_7501,N_8178);
nor U8993 (N_8993,N_7983,N_7874);
and U8994 (N_8994,N_7866,N_7989);
or U8995 (N_8995,N_7944,N_7871);
and U8996 (N_8996,N_7698,N_7934);
and U8997 (N_8997,N_8169,N_8073);
and U8998 (N_8998,N_7577,N_7666);
nand U8999 (N_8999,N_7816,N_7711);
nand U9000 (N_9000,N_8542,N_8272);
and U9001 (N_9001,N_8411,N_8787);
or U9002 (N_9002,N_8814,N_8559);
nor U9003 (N_9003,N_8502,N_8384);
nor U9004 (N_9004,N_8507,N_8983);
or U9005 (N_9005,N_8512,N_8882);
nand U9006 (N_9006,N_8344,N_8737);
and U9007 (N_9007,N_8899,N_8838);
or U9008 (N_9008,N_8661,N_8844);
and U9009 (N_9009,N_8812,N_8251);
or U9010 (N_9010,N_8354,N_8978);
nor U9011 (N_9011,N_8956,N_8475);
and U9012 (N_9012,N_8258,N_8527);
and U9013 (N_9013,N_8276,N_8607);
xnor U9014 (N_9014,N_8807,N_8491);
nor U9015 (N_9015,N_8995,N_8375);
xor U9016 (N_9016,N_8940,N_8690);
and U9017 (N_9017,N_8701,N_8855);
and U9018 (N_9018,N_8610,N_8526);
and U9019 (N_9019,N_8600,N_8890);
nand U9020 (N_9020,N_8285,N_8688);
nand U9021 (N_9021,N_8741,N_8565);
nor U9022 (N_9022,N_8457,N_8985);
and U9023 (N_9023,N_8637,N_8372);
and U9024 (N_9024,N_8413,N_8631);
and U9025 (N_9025,N_8823,N_8310);
or U9026 (N_9026,N_8874,N_8386);
and U9027 (N_9027,N_8443,N_8510);
or U9028 (N_9028,N_8558,N_8277);
or U9029 (N_9029,N_8324,N_8572);
nand U9030 (N_9030,N_8433,N_8820);
nand U9031 (N_9031,N_8795,N_8562);
nor U9032 (N_9032,N_8391,N_8529);
and U9033 (N_9033,N_8796,N_8392);
and U9034 (N_9034,N_8606,N_8545);
and U9035 (N_9035,N_8722,N_8909);
nor U9036 (N_9036,N_8912,N_8649);
and U9037 (N_9037,N_8412,N_8813);
nor U9038 (N_9038,N_8318,N_8366);
and U9039 (N_9039,N_8539,N_8908);
and U9040 (N_9040,N_8317,N_8867);
nand U9041 (N_9041,N_8346,N_8982);
or U9042 (N_9042,N_8699,N_8416);
nand U9043 (N_9043,N_8705,N_8902);
nor U9044 (N_9044,N_8835,N_8388);
nor U9045 (N_9045,N_8847,N_8656);
or U9046 (N_9046,N_8926,N_8733);
or U9047 (N_9047,N_8437,N_8967);
nor U9048 (N_9048,N_8336,N_8356);
xnor U9049 (N_9049,N_8691,N_8766);
and U9050 (N_9050,N_8948,N_8996);
nand U9051 (N_9051,N_8801,N_8553);
nor U9052 (N_9052,N_8773,N_8364);
nor U9053 (N_9053,N_8858,N_8765);
nor U9054 (N_9054,N_8357,N_8652);
nor U9055 (N_9055,N_8399,N_8341);
and U9056 (N_9056,N_8575,N_8824);
and U9057 (N_9057,N_8643,N_8464);
nand U9058 (N_9058,N_8450,N_8316);
or U9059 (N_9059,N_8551,N_8414);
nand U9060 (N_9060,N_8471,N_8634);
or U9061 (N_9061,N_8404,N_8546);
xnor U9062 (N_9062,N_8330,N_8642);
xor U9063 (N_9063,N_8872,N_8495);
xor U9064 (N_9064,N_8603,N_8467);
or U9065 (N_9065,N_8396,N_8877);
or U9066 (N_9066,N_8525,N_8776);
xnor U9067 (N_9067,N_8537,N_8334);
nor U9068 (N_9068,N_8370,N_8616);
and U9069 (N_9069,N_8530,N_8628);
nand U9070 (N_9070,N_8721,N_8683);
or U9071 (N_9071,N_8478,N_8786);
xor U9072 (N_9072,N_8481,N_8547);
nor U9073 (N_9073,N_8746,N_8793);
nand U9074 (N_9074,N_8816,N_8654);
nor U9075 (N_9075,N_8668,N_8720);
nand U9076 (N_9076,N_8968,N_8255);
and U9077 (N_9077,N_8871,N_8472);
or U9078 (N_9078,N_8454,N_8405);
nand U9079 (N_9079,N_8599,N_8687);
or U9080 (N_9080,N_8355,N_8659);
and U9081 (N_9081,N_8254,N_8830);
xnor U9082 (N_9082,N_8640,N_8923);
xor U9083 (N_9083,N_8928,N_8415);
nand U9084 (N_9084,N_8915,N_8750);
or U9085 (N_9085,N_8630,N_8887);
or U9086 (N_9086,N_8410,N_8358);
and U9087 (N_9087,N_8651,N_8519);
or U9088 (N_9088,N_8543,N_8518);
or U9089 (N_9089,N_8362,N_8712);
nand U9090 (N_9090,N_8431,N_8911);
nand U9091 (N_9091,N_8970,N_8740);
nor U9092 (N_9092,N_8520,N_8756);
and U9093 (N_9093,N_8647,N_8513);
nand U9094 (N_9094,N_8760,N_8323);
nand U9095 (N_9095,N_8440,N_8594);
nand U9096 (N_9096,N_8989,N_8291);
nand U9097 (N_9097,N_8508,N_8260);
nor U9098 (N_9098,N_8671,N_8639);
nand U9099 (N_9099,N_8762,N_8723);
and U9100 (N_9100,N_8865,N_8598);
or U9101 (N_9101,N_8955,N_8696);
nor U9102 (N_9102,N_8635,N_8252);
nand U9103 (N_9103,N_8307,N_8994);
nor U9104 (N_9104,N_8417,N_8658);
nand U9105 (N_9105,N_8966,N_8792);
or U9106 (N_9106,N_8663,N_8296);
and U9107 (N_9107,N_8282,N_8964);
nor U9108 (N_9108,N_8301,N_8257);
nor U9109 (N_9109,N_8477,N_8962);
nand U9110 (N_9110,N_8273,N_8314);
nand U9111 (N_9111,N_8561,N_8468);
or U9112 (N_9112,N_8275,N_8829);
nor U9113 (N_9113,N_8328,N_8303);
nor U9114 (N_9114,N_8430,N_8840);
nand U9115 (N_9115,N_8939,N_8425);
and U9116 (N_9116,N_8784,N_8724);
and U9117 (N_9117,N_8420,N_8706);
and U9118 (N_9118,N_8268,N_8798);
nand U9119 (N_9119,N_8408,N_8728);
and U9120 (N_9120,N_8866,N_8393);
nand U9121 (N_9121,N_8905,N_8832);
xor U9122 (N_9122,N_8574,N_8757);
nor U9123 (N_9123,N_8748,N_8903);
and U9124 (N_9124,N_8734,N_8483);
nor U9125 (N_9125,N_8624,N_8352);
xor U9126 (N_9126,N_8997,N_8522);
nor U9127 (N_9127,N_8774,N_8421);
or U9128 (N_9128,N_8505,N_8704);
and U9129 (N_9129,N_8782,N_8906);
and U9130 (N_9130,N_8917,N_8770);
or U9131 (N_9131,N_8515,N_8993);
or U9132 (N_9132,N_8895,N_8644);
nand U9133 (N_9133,N_8550,N_8571);
nor U9134 (N_9134,N_8609,N_8426);
nand U9135 (N_9135,N_8901,N_8359);
nor U9136 (N_9136,N_8287,N_8514);
and U9137 (N_9137,N_8921,N_8329);
nand U9138 (N_9138,N_8839,N_8753);
xor U9139 (N_9139,N_8579,N_8831);
nor U9140 (N_9140,N_8383,N_8294);
and U9141 (N_9141,N_8738,N_8933);
nand U9142 (N_9142,N_8290,N_8949);
nand U9143 (N_9143,N_8870,N_8886);
or U9144 (N_9144,N_8595,N_8367);
and U9145 (N_9145,N_8913,N_8567);
and U9146 (N_9146,N_8313,N_8374);
or U9147 (N_9147,N_8662,N_8938);
or U9148 (N_9148,N_8821,N_8988);
nand U9149 (N_9149,N_8946,N_8380);
nand U9150 (N_9150,N_8511,N_8509);
or U9151 (N_9151,N_8278,N_8250);
xor U9152 (N_9152,N_8263,N_8486);
xor U9153 (N_9153,N_8361,N_8685);
and U9154 (N_9154,N_8351,N_8907);
and U9155 (N_9155,N_8736,N_8369);
and U9156 (N_9156,N_8999,N_8689);
nand U9157 (N_9157,N_8944,N_8755);
nor U9158 (N_9158,N_8959,N_8629);
xnor U9159 (N_9159,N_8836,N_8854);
and U9160 (N_9160,N_8758,N_8549);
nand U9161 (N_9161,N_8934,N_8590);
and U9162 (N_9162,N_8343,N_8349);
nor U9163 (N_9163,N_8735,N_8397);
nor U9164 (N_9164,N_8779,N_8264);
nor U9165 (N_9165,N_8400,N_8672);
or U9166 (N_9166,N_8863,N_8697);
or U9167 (N_9167,N_8641,N_8969);
nand U9168 (N_9168,N_8802,N_8665);
nand U9169 (N_9169,N_8666,N_8764);
nor U9170 (N_9170,N_8568,N_8677);
nand U9171 (N_9171,N_8569,N_8407);
nand U9172 (N_9172,N_8675,N_8961);
and U9173 (N_9173,N_8267,N_8992);
or U9174 (N_9174,N_8381,N_8780);
nand U9175 (N_9175,N_8743,N_8794);
xnor U9176 (N_9176,N_8991,N_8850);
or U9177 (N_9177,N_8597,N_8494);
and U9178 (N_9178,N_8608,N_8853);
and U9179 (N_9179,N_8975,N_8582);
and U9180 (N_9180,N_8533,N_8876);
nor U9181 (N_9181,N_8914,N_8730);
nand U9182 (N_9182,N_8881,N_8726);
or U9183 (N_9183,N_8893,N_8935);
or U9184 (N_9184,N_8456,N_8604);
nor U9185 (N_9185,N_8521,N_8954);
and U9186 (N_9186,N_8419,N_8271);
and U9187 (N_9187,N_8427,N_8398);
nand U9188 (N_9188,N_8517,N_8432);
nand U9189 (N_9189,N_8327,N_8470);
or U9190 (N_9190,N_8605,N_8548);
nor U9191 (N_9191,N_8702,N_8304);
nand U9192 (N_9192,N_8958,N_8896);
nor U9193 (N_9193,N_8984,N_8971);
nand U9194 (N_9194,N_8990,N_8768);
or U9195 (N_9195,N_8857,N_8611);
nor U9196 (N_9196,N_8588,N_8274);
and U9197 (N_9197,N_8805,N_8645);
nor U9198 (N_9198,N_8418,N_8862);
nand U9199 (N_9199,N_8960,N_8297);
nor U9200 (N_9200,N_8373,N_8434);
nand U9201 (N_9201,N_8564,N_8972);
or U9202 (N_9202,N_8504,N_8700);
xor U9203 (N_9203,N_8657,N_8834);
xnor U9204 (N_9204,N_8761,N_8803);
xnor U9205 (N_9205,N_8843,N_8501);
and U9206 (N_9206,N_8583,N_8679);
or U9207 (N_9207,N_8406,N_8438);
and U9208 (N_9208,N_8286,N_8315);
nor U9209 (N_9209,N_8394,N_8910);
nor U9210 (N_9210,N_8566,N_8601);
nor U9211 (N_9211,N_8480,N_8487);
nand U9212 (N_9212,N_8833,N_8292);
nor U9213 (N_9213,N_8580,N_8321);
and U9214 (N_9214,N_8259,N_8473);
and U9215 (N_9215,N_8445,N_8716);
nand U9216 (N_9216,N_8459,N_8965);
and U9217 (N_9217,N_8632,N_8729);
nor U9218 (N_9218,N_8709,N_8469);
nor U9219 (N_9219,N_8573,N_8253);
and U9220 (N_9220,N_8621,N_8889);
and U9221 (N_9221,N_8749,N_8841);
nand U9222 (N_9222,N_8849,N_8810);
nor U9223 (N_9223,N_8422,N_8484);
nand U9224 (N_9224,N_8860,N_8325);
xor U9225 (N_9225,N_8602,N_8293);
or U9226 (N_9226,N_8261,N_8892);
nand U9227 (N_9227,N_8929,N_8648);
or U9228 (N_9228,N_8667,N_8952);
nand U9229 (N_9229,N_8528,N_8879);
or U9230 (N_9230,N_8458,N_8653);
nand U9231 (N_9231,N_8715,N_8937);
nor U9232 (N_9232,N_8342,N_8717);
nor U9233 (N_9233,N_8376,N_8680);
nor U9234 (N_9234,N_8806,N_8861);
xor U9235 (N_9235,N_8664,N_8489);
or U9236 (N_9236,N_8791,N_8300);
or U9237 (N_9237,N_8541,N_8320);
or U9238 (N_9238,N_8638,N_8739);
or U9239 (N_9239,N_8920,N_8326);
nand U9240 (N_9240,N_8353,N_8423);
nor U9241 (N_9241,N_8815,N_8845);
or U9242 (N_9242,N_8822,N_8591);
and U9243 (N_9243,N_8389,N_8347);
and U9244 (N_9244,N_8488,N_8873);
nor U9245 (N_9245,N_8676,N_8731);
and U9246 (N_9246,N_8693,N_8981);
nand U9247 (N_9247,N_8880,N_8950);
or U9248 (N_9248,N_8625,N_8851);
nand U9249 (N_9249,N_8500,N_8618);
nand U9250 (N_9250,N_8395,N_8837);
or U9251 (N_9251,N_8612,N_8744);
or U9252 (N_9252,N_8584,N_8544);
nand U9253 (N_9253,N_8563,N_8556);
xnor U9254 (N_9254,N_8345,N_8436);
nand U9255 (N_9255,N_8963,N_8852);
nand U9256 (N_9256,N_8589,N_8555);
nand U9257 (N_9257,N_8825,N_8875);
or U9258 (N_9258,N_8577,N_8581);
and U9259 (N_9259,N_8516,N_8614);
nand U9260 (N_9260,N_8789,N_8924);
or U9261 (N_9261,N_8987,N_8977);
and U9262 (N_9262,N_8681,N_8686);
nor U9263 (N_9263,N_8570,N_8884);
or U9264 (N_9264,N_8898,N_8781);
nand U9265 (N_9265,N_8695,N_8382);
or U9266 (N_9266,N_8769,N_8461);
nor U9267 (N_9267,N_8592,N_8348);
nor U9268 (N_9268,N_8897,N_8891);
nor U9269 (N_9269,N_8936,N_8312);
nor U9270 (N_9270,N_8465,N_8980);
or U9271 (N_9271,N_8280,N_8718);
nor U9272 (N_9272,N_8279,N_8623);
nor U9273 (N_9273,N_8435,N_8620);
or U9274 (N_9274,N_8868,N_8387);
or U9275 (N_9275,N_8335,N_8476);
nor U9276 (N_9276,N_8492,N_8650);
or U9277 (N_9277,N_8455,N_8298);
nor U9278 (N_9278,N_8811,N_8390);
nand U9279 (N_9279,N_8446,N_8503);
nand U9280 (N_9280,N_8797,N_8957);
or U9281 (N_9281,N_8826,N_8878);
nand U9282 (N_9282,N_8586,N_8560);
nand U9283 (N_9283,N_8775,N_8619);
nand U9284 (N_9284,N_8262,N_8692);
or U9285 (N_9285,N_8819,N_8943);
nand U9286 (N_9286,N_8827,N_8904);
or U9287 (N_9287,N_8885,N_8682);
and U9288 (N_9288,N_8622,N_8617);
nand U9289 (N_9289,N_8771,N_8540);
or U9290 (N_9290,N_8711,N_8684);
nor U9291 (N_9291,N_8385,N_8842);
nand U9292 (N_9292,N_8883,N_8447);
xnor U9293 (N_9293,N_8922,N_8284);
and U9294 (N_9294,N_8932,N_8670);
or U9295 (N_9295,N_8266,N_8256);
nand U9296 (N_9296,N_8295,N_8269);
nor U9297 (N_9297,N_8916,N_8674);
xnor U9298 (N_9298,N_8751,N_8485);
xor U9299 (N_9299,N_8747,N_8532);
nor U9300 (N_9300,N_8535,N_8424);
or U9301 (N_9301,N_8496,N_8919);
nor U9302 (N_9302,N_8332,N_8772);
nand U9303 (N_9303,N_8785,N_8808);
or U9304 (N_9304,N_8448,N_8360);
nand U9305 (N_9305,N_8429,N_8974);
nand U9306 (N_9306,N_8466,N_8451);
nand U9307 (N_9307,N_8463,N_8305);
and U9308 (N_9308,N_8322,N_8497);
and U9309 (N_9309,N_8698,N_8453);
and U9310 (N_9310,N_8350,N_8973);
and U9311 (N_9311,N_8462,N_8918);
nor U9312 (N_9312,N_8587,N_8333);
nand U9313 (N_9313,N_8552,N_8818);
nand U9314 (N_9314,N_8719,N_8615);
nor U9315 (N_9315,N_8319,N_8379);
and U9316 (N_9316,N_8809,N_8790);
nand U9317 (N_9317,N_8931,N_8627);
or U9318 (N_9318,N_8976,N_8763);
nor U9319 (N_9319,N_8678,N_8534);
nand U9320 (N_9320,N_8767,N_8311);
or U9321 (N_9321,N_8339,N_8646);
and U9322 (N_9322,N_8449,N_8506);
and U9323 (N_9323,N_8927,N_8554);
and U9324 (N_9324,N_8900,N_8368);
xor U9325 (N_9325,N_8925,N_8673);
nand U9326 (N_9326,N_8498,N_8864);
or U9327 (N_9327,N_8479,N_8947);
nor U9328 (N_9328,N_8777,N_8452);
xor U9329 (N_9329,N_8846,N_8371);
nor U9330 (N_9330,N_8804,N_8714);
xnor U9331 (N_9331,N_8593,N_8578);
nand U9332 (N_9332,N_8930,N_8270);
nand U9333 (N_9333,N_8669,N_8365);
and U9334 (N_9334,N_8759,N_8490);
nand U9335 (N_9335,N_8707,N_8538);
nor U9336 (N_9336,N_8283,N_8942);
or U9337 (N_9337,N_8660,N_8703);
nor U9338 (N_9338,N_8727,N_8265);
and U9339 (N_9339,N_8941,N_8289);
xor U9340 (N_9340,N_8713,N_8576);
nor U9341 (N_9341,N_8894,N_8331);
or U9342 (N_9342,N_8859,N_8708);
xnor U9343 (N_9343,N_8888,N_8482);
nand U9344 (N_9344,N_8636,N_8302);
or U9345 (N_9345,N_8402,N_8401);
or U9346 (N_9346,N_8378,N_8585);
or U9347 (N_9347,N_8856,N_8281);
and U9348 (N_9348,N_8444,N_8694);
and U9349 (N_9349,N_8800,N_8953);
nand U9350 (N_9350,N_8732,N_8523);
and U9351 (N_9351,N_8403,N_8945);
nor U9352 (N_9352,N_8409,N_8308);
or U9353 (N_9353,N_8428,N_8754);
and U9354 (N_9354,N_8557,N_8596);
and U9355 (N_9355,N_8363,N_8613);
and U9356 (N_9356,N_8869,N_8742);
xnor U9357 (N_9357,N_8848,N_8337);
or U9358 (N_9358,N_8986,N_8441);
and U9359 (N_9359,N_8309,N_8377);
nand U9360 (N_9360,N_8499,N_8626);
and U9361 (N_9361,N_8524,N_8745);
and U9362 (N_9362,N_8778,N_8783);
and U9363 (N_9363,N_8306,N_8655);
nor U9364 (N_9364,N_8998,N_8536);
or U9365 (N_9365,N_8338,N_8299);
xor U9366 (N_9366,N_8752,N_8633);
nor U9367 (N_9367,N_8460,N_8828);
nor U9368 (N_9368,N_8951,N_8799);
nand U9369 (N_9369,N_8788,N_8439);
or U9370 (N_9370,N_8725,N_8493);
and U9371 (N_9371,N_8531,N_8710);
nand U9372 (N_9372,N_8474,N_8817);
nor U9373 (N_9373,N_8340,N_8442);
and U9374 (N_9374,N_8979,N_8288);
and U9375 (N_9375,N_8273,N_8765);
nand U9376 (N_9376,N_8541,N_8962);
or U9377 (N_9377,N_8798,N_8900);
or U9378 (N_9378,N_8321,N_8454);
or U9379 (N_9379,N_8964,N_8694);
nand U9380 (N_9380,N_8734,N_8910);
nor U9381 (N_9381,N_8841,N_8260);
xor U9382 (N_9382,N_8623,N_8821);
xnor U9383 (N_9383,N_8864,N_8461);
nand U9384 (N_9384,N_8945,N_8383);
and U9385 (N_9385,N_8844,N_8404);
nand U9386 (N_9386,N_8393,N_8551);
xor U9387 (N_9387,N_8613,N_8813);
nand U9388 (N_9388,N_8606,N_8675);
or U9389 (N_9389,N_8650,N_8721);
and U9390 (N_9390,N_8532,N_8272);
nand U9391 (N_9391,N_8758,N_8969);
nor U9392 (N_9392,N_8868,N_8789);
and U9393 (N_9393,N_8819,N_8922);
or U9394 (N_9394,N_8602,N_8712);
or U9395 (N_9395,N_8341,N_8300);
nand U9396 (N_9396,N_8529,N_8723);
and U9397 (N_9397,N_8431,N_8780);
xnor U9398 (N_9398,N_8542,N_8262);
nand U9399 (N_9399,N_8352,N_8918);
or U9400 (N_9400,N_8708,N_8505);
nor U9401 (N_9401,N_8958,N_8759);
or U9402 (N_9402,N_8337,N_8272);
and U9403 (N_9403,N_8623,N_8609);
nor U9404 (N_9404,N_8338,N_8702);
and U9405 (N_9405,N_8979,N_8293);
nand U9406 (N_9406,N_8498,N_8669);
or U9407 (N_9407,N_8293,N_8552);
xnor U9408 (N_9408,N_8305,N_8993);
nor U9409 (N_9409,N_8682,N_8683);
or U9410 (N_9410,N_8330,N_8648);
or U9411 (N_9411,N_8746,N_8832);
or U9412 (N_9412,N_8514,N_8732);
nor U9413 (N_9413,N_8629,N_8588);
or U9414 (N_9414,N_8297,N_8453);
nor U9415 (N_9415,N_8478,N_8287);
and U9416 (N_9416,N_8388,N_8362);
nand U9417 (N_9417,N_8816,N_8303);
xnor U9418 (N_9418,N_8629,N_8388);
or U9419 (N_9419,N_8541,N_8619);
or U9420 (N_9420,N_8849,N_8373);
nor U9421 (N_9421,N_8352,N_8906);
nand U9422 (N_9422,N_8843,N_8873);
nand U9423 (N_9423,N_8316,N_8806);
nor U9424 (N_9424,N_8880,N_8638);
and U9425 (N_9425,N_8584,N_8916);
nand U9426 (N_9426,N_8941,N_8518);
and U9427 (N_9427,N_8637,N_8319);
or U9428 (N_9428,N_8408,N_8259);
nand U9429 (N_9429,N_8959,N_8265);
nor U9430 (N_9430,N_8767,N_8494);
nand U9431 (N_9431,N_8586,N_8613);
and U9432 (N_9432,N_8358,N_8791);
nand U9433 (N_9433,N_8790,N_8525);
nand U9434 (N_9434,N_8582,N_8390);
nor U9435 (N_9435,N_8471,N_8488);
xor U9436 (N_9436,N_8295,N_8517);
and U9437 (N_9437,N_8429,N_8257);
and U9438 (N_9438,N_8380,N_8900);
or U9439 (N_9439,N_8900,N_8450);
nor U9440 (N_9440,N_8927,N_8464);
and U9441 (N_9441,N_8914,N_8334);
nor U9442 (N_9442,N_8817,N_8313);
nand U9443 (N_9443,N_8876,N_8728);
nand U9444 (N_9444,N_8582,N_8261);
or U9445 (N_9445,N_8304,N_8870);
nor U9446 (N_9446,N_8822,N_8309);
xnor U9447 (N_9447,N_8470,N_8346);
and U9448 (N_9448,N_8939,N_8694);
or U9449 (N_9449,N_8668,N_8317);
nor U9450 (N_9450,N_8865,N_8651);
or U9451 (N_9451,N_8843,N_8877);
nand U9452 (N_9452,N_8259,N_8818);
nor U9453 (N_9453,N_8698,N_8783);
xnor U9454 (N_9454,N_8596,N_8299);
nor U9455 (N_9455,N_8766,N_8578);
nor U9456 (N_9456,N_8548,N_8763);
and U9457 (N_9457,N_8309,N_8414);
nor U9458 (N_9458,N_8467,N_8731);
and U9459 (N_9459,N_8406,N_8749);
and U9460 (N_9460,N_8813,N_8892);
or U9461 (N_9461,N_8780,N_8307);
or U9462 (N_9462,N_8312,N_8833);
nand U9463 (N_9463,N_8702,N_8704);
or U9464 (N_9464,N_8715,N_8540);
nor U9465 (N_9465,N_8902,N_8636);
nor U9466 (N_9466,N_8303,N_8645);
nor U9467 (N_9467,N_8909,N_8476);
and U9468 (N_9468,N_8941,N_8668);
nand U9469 (N_9469,N_8522,N_8382);
and U9470 (N_9470,N_8331,N_8684);
nand U9471 (N_9471,N_8916,N_8463);
nand U9472 (N_9472,N_8465,N_8978);
and U9473 (N_9473,N_8681,N_8383);
nand U9474 (N_9474,N_8728,N_8372);
and U9475 (N_9475,N_8907,N_8660);
or U9476 (N_9476,N_8936,N_8392);
nand U9477 (N_9477,N_8441,N_8391);
or U9478 (N_9478,N_8534,N_8711);
and U9479 (N_9479,N_8528,N_8275);
nor U9480 (N_9480,N_8267,N_8454);
nor U9481 (N_9481,N_8560,N_8421);
nand U9482 (N_9482,N_8667,N_8297);
nor U9483 (N_9483,N_8943,N_8759);
and U9484 (N_9484,N_8884,N_8675);
nor U9485 (N_9485,N_8405,N_8277);
or U9486 (N_9486,N_8305,N_8499);
nand U9487 (N_9487,N_8860,N_8746);
or U9488 (N_9488,N_8536,N_8792);
or U9489 (N_9489,N_8672,N_8340);
or U9490 (N_9490,N_8375,N_8617);
and U9491 (N_9491,N_8783,N_8285);
or U9492 (N_9492,N_8350,N_8533);
or U9493 (N_9493,N_8839,N_8897);
and U9494 (N_9494,N_8874,N_8770);
nor U9495 (N_9495,N_8555,N_8761);
nor U9496 (N_9496,N_8576,N_8333);
nor U9497 (N_9497,N_8914,N_8939);
xor U9498 (N_9498,N_8870,N_8468);
nor U9499 (N_9499,N_8890,N_8575);
or U9500 (N_9500,N_8924,N_8762);
xor U9501 (N_9501,N_8916,N_8331);
nand U9502 (N_9502,N_8842,N_8776);
and U9503 (N_9503,N_8675,N_8572);
or U9504 (N_9504,N_8600,N_8349);
nand U9505 (N_9505,N_8988,N_8341);
and U9506 (N_9506,N_8694,N_8758);
or U9507 (N_9507,N_8265,N_8606);
nor U9508 (N_9508,N_8985,N_8960);
or U9509 (N_9509,N_8953,N_8924);
or U9510 (N_9510,N_8333,N_8829);
nor U9511 (N_9511,N_8840,N_8414);
or U9512 (N_9512,N_8935,N_8426);
and U9513 (N_9513,N_8367,N_8629);
or U9514 (N_9514,N_8783,N_8946);
nor U9515 (N_9515,N_8376,N_8931);
or U9516 (N_9516,N_8686,N_8885);
nand U9517 (N_9517,N_8964,N_8789);
nand U9518 (N_9518,N_8403,N_8824);
nand U9519 (N_9519,N_8449,N_8743);
and U9520 (N_9520,N_8853,N_8583);
nor U9521 (N_9521,N_8709,N_8389);
or U9522 (N_9522,N_8666,N_8728);
or U9523 (N_9523,N_8770,N_8700);
and U9524 (N_9524,N_8701,N_8996);
nor U9525 (N_9525,N_8827,N_8954);
and U9526 (N_9526,N_8982,N_8882);
nor U9527 (N_9527,N_8883,N_8589);
and U9528 (N_9528,N_8443,N_8277);
or U9529 (N_9529,N_8763,N_8424);
nand U9530 (N_9530,N_8503,N_8944);
or U9531 (N_9531,N_8686,N_8997);
and U9532 (N_9532,N_8733,N_8540);
or U9533 (N_9533,N_8690,N_8586);
or U9534 (N_9534,N_8354,N_8660);
nor U9535 (N_9535,N_8987,N_8681);
xor U9536 (N_9536,N_8568,N_8792);
nand U9537 (N_9537,N_8520,N_8786);
or U9538 (N_9538,N_8552,N_8520);
xnor U9539 (N_9539,N_8626,N_8933);
nor U9540 (N_9540,N_8999,N_8842);
nand U9541 (N_9541,N_8413,N_8328);
and U9542 (N_9542,N_8992,N_8539);
or U9543 (N_9543,N_8921,N_8448);
and U9544 (N_9544,N_8478,N_8829);
or U9545 (N_9545,N_8654,N_8797);
nor U9546 (N_9546,N_8584,N_8619);
or U9547 (N_9547,N_8929,N_8253);
and U9548 (N_9548,N_8915,N_8514);
nand U9549 (N_9549,N_8616,N_8568);
or U9550 (N_9550,N_8501,N_8489);
and U9551 (N_9551,N_8749,N_8626);
nor U9552 (N_9552,N_8630,N_8859);
and U9553 (N_9553,N_8367,N_8335);
and U9554 (N_9554,N_8290,N_8606);
nor U9555 (N_9555,N_8516,N_8305);
or U9556 (N_9556,N_8956,N_8431);
and U9557 (N_9557,N_8256,N_8733);
xor U9558 (N_9558,N_8547,N_8718);
nand U9559 (N_9559,N_8299,N_8692);
nand U9560 (N_9560,N_8781,N_8619);
nand U9561 (N_9561,N_8810,N_8506);
and U9562 (N_9562,N_8993,N_8815);
or U9563 (N_9563,N_8347,N_8842);
and U9564 (N_9564,N_8627,N_8690);
and U9565 (N_9565,N_8873,N_8368);
xor U9566 (N_9566,N_8564,N_8785);
or U9567 (N_9567,N_8914,N_8645);
nor U9568 (N_9568,N_8381,N_8417);
and U9569 (N_9569,N_8388,N_8887);
and U9570 (N_9570,N_8520,N_8517);
and U9571 (N_9571,N_8775,N_8373);
xnor U9572 (N_9572,N_8640,N_8897);
nand U9573 (N_9573,N_8648,N_8705);
nor U9574 (N_9574,N_8402,N_8392);
and U9575 (N_9575,N_8764,N_8597);
nand U9576 (N_9576,N_8488,N_8696);
or U9577 (N_9577,N_8973,N_8932);
nor U9578 (N_9578,N_8680,N_8658);
nand U9579 (N_9579,N_8615,N_8815);
nor U9580 (N_9580,N_8640,N_8284);
and U9581 (N_9581,N_8770,N_8527);
and U9582 (N_9582,N_8412,N_8329);
nor U9583 (N_9583,N_8269,N_8375);
and U9584 (N_9584,N_8536,N_8396);
nor U9585 (N_9585,N_8997,N_8606);
and U9586 (N_9586,N_8800,N_8885);
and U9587 (N_9587,N_8971,N_8703);
or U9588 (N_9588,N_8995,N_8605);
or U9589 (N_9589,N_8749,N_8525);
or U9590 (N_9590,N_8432,N_8465);
nand U9591 (N_9591,N_8491,N_8487);
xor U9592 (N_9592,N_8419,N_8832);
xnor U9593 (N_9593,N_8605,N_8785);
and U9594 (N_9594,N_8698,N_8958);
nor U9595 (N_9595,N_8679,N_8497);
nor U9596 (N_9596,N_8254,N_8278);
nor U9597 (N_9597,N_8281,N_8713);
nand U9598 (N_9598,N_8251,N_8387);
and U9599 (N_9599,N_8667,N_8822);
or U9600 (N_9600,N_8764,N_8549);
and U9601 (N_9601,N_8911,N_8654);
nor U9602 (N_9602,N_8284,N_8894);
or U9603 (N_9603,N_8927,N_8751);
xnor U9604 (N_9604,N_8569,N_8635);
or U9605 (N_9605,N_8885,N_8483);
or U9606 (N_9606,N_8400,N_8343);
nor U9607 (N_9607,N_8586,N_8816);
and U9608 (N_9608,N_8272,N_8489);
nor U9609 (N_9609,N_8726,N_8380);
and U9610 (N_9610,N_8620,N_8859);
and U9611 (N_9611,N_8721,N_8567);
nor U9612 (N_9612,N_8620,N_8316);
xor U9613 (N_9613,N_8589,N_8353);
and U9614 (N_9614,N_8284,N_8836);
or U9615 (N_9615,N_8997,N_8521);
nand U9616 (N_9616,N_8845,N_8903);
or U9617 (N_9617,N_8738,N_8894);
and U9618 (N_9618,N_8981,N_8334);
nand U9619 (N_9619,N_8958,N_8616);
or U9620 (N_9620,N_8331,N_8635);
nand U9621 (N_9621,N_8543,N_8969);
xor U9622 (N_9622,N_8755,N_8371);
or U9623 (N_9623,N_8888,N_8742);
and U9624 (N_9624,N_8587,N_8579);
nor U9625 (N_9625,N_8455,N_8610);
and U9626 (N_9626,N_8398,N_8693);
nor U9627 (N_9627,N_8831,N_8443);
and U9628 (N_9628,N_8297,N_8581);
nand U9629 (N_9629,N_8277,N_8404);
nand U9630 (N_9630,N_8964,N_8313);
nand U9631 (N_9631,N_8774,N_8392);
nor U9632 (N_9632,N_8982,N_8408);
or U9633 (N_9633,N_8996,N_8399);
or U9634 (N_9634,N_8721,N_8363);
or U9635 (N_9635,N_8949,N_8586);
nor U9636 (N_9636,N_8420,N_8262);
nand U9637 (N_9637,N_8439,N_8407);
nor U9638 (N_9638,N_8574,N_8532);
xor U9639 (N_9639,N_8891,N_8780);
nand U9640 (N_9640,N_8754,N_8277);
and U9641 (N_9641,N_8451,N_8996);
nand U9642 (N_9642,N_8984,N_8929);
nand U9643 (N_9643,N_8942,N_8406);
nand U9644 (N_9644,N_8586,N_8557);
or U9645 (N_9645,N_8466,N_8410);
nor U9646 (N_9646,N_8473,N_8638);
or U9647 (N_9647,N_8576,N_8860);
nand U9648 (N_9648,N_8291,N_8439);
and U9649 (N_9649,N_8784,N_8996);
nor U9650 (N_9650,N_8250,N_8924);
nand U9651 (N_9651,N_8361,N_8468);
xor U9652 (N_9652,N_8669,N_8904);
and U9653 (N_9653,N_8277,N_8605);
xor U9654 (N_9654,N_8610,N_8268);
or U9655 (N_9655,N_8600,N_8383);
nor U9656 (N_9656,N_8790,N_8307);
nor U9657 (N_9657,N_8660,N_8783);
and U9658 (N_9658,N_8614,N_8857);
and U9659 (N_9659,N_8875,N_8423);
nand U9660 (N_9660,N_8962,N_8859);
nor U9661 (N_9661,N_8274,N_8726);
nand U9662 (N_9662,N_8850,N_8936);
nor U9663 (N_9663,N_8522,N_8940);
and U9664 (N_9664,N_8950,N_8926);
or U9665 (N_9665,N_8853,N_8793);
nand U9666 (N_9666,N_8287,N_8268);
nor U9667 (N_9667,N_8259,N_8760);
nand U9668 (N_9668,N_8444,N_8676);
nand U9669 (N_9669,N_8992,N_8332);
or U9670 (N_9670,N_8505,N_8801);
nand U9671 (N_9671,N_8552,N_8263);
nand U9672 (N_9672,N_8726,N_8613);
nor U9673 (N_9673,N_8559,N_8555);
nor U9674 (N_9674,N_8263,N_8797);
nor U9675 (N_9675,N_8682,N_8499);
nor U9676 (N_9676,N_8953,N_8550);
nor U9677 (N_9677,N_8867,N_8697);
and U9678 (N_9678,N_8656,N_8660);
and U9679 (N_9679,N_8887,N_8913);
nand U9680 (N_9680,N_8443,N_8992);
and U9681 (N_9681,N_8764,N_8297);
nand U9682 (N_9682,N_8726,N_8528);
and U9683 (N_9683,N_8794,N_8861);
nor U9684 (N_9684,N_8968,N_8979);
and U9685 (N_9685,N_8734,N_8501);
and U9686 (N_9686,N_8834,N_8909);
nand U9687 (N_9687,N_8912,N_8393);
nand U9688 (N_9688,N_8894,N_8636);
nand U9689 (N_9689,N_8808,N_8416);
nor U9690 (N_9690,N_8415,N_8396);
nand U9691 (N_9691,N_8976,N_8307);
and U9692 (N_9692,N_8735,N_8418);
or U9693 (N_9693,N_8988,N_8361);
and U9694 (N_9694,N_8865,N_8679);
and U9695 (N_9695,N_8617,N_8894);
or U9696 (N_9696,N_8820,N_8252);
or U9697 (N_9697,N_8489,N_8758);
or U9698 (N_9698,N_8355,N_8450);
or U9699 (N_9699,N_8542,N_8785);
xnor U9700 (N_9700,N_8536,N_8727);
nor U9701 (N_9701,N_8599,N_8415);
nand U9702 (N_9702,N_8974,N_8640);
nand U9703 (N_9703,N_8998,N_8899);
and U9704 (N_9704,N_8827,N_8869);
and U9705 (N_9705,N_8420,N_8433);
or U9706 (N_9706,N_8834,N_8898);
and U9707 (N_9707,N_8768,N_8988);
nor U9708 (N_9708,N_8353,N_8633);
nor U9709 (N_9709,N_8354,N_8840);
nor U9710 (N_9710,N_8699,N_8468);
or U9711 (N_9711,N_8766,N_8445);
and U9712 (N_9712,N_8576,N_8784);
nand U9713 (N_9713,N_8736,N_8818);
nor U9714 (N_9714,N_8362,N_8864);
nand U9715 (N_9715,N_8260,N_8654);
nor U9716 (N_9716,N_8392,N_8655);
nand U9717 (N_9717,N_8422,N_8498);
or U9718 (N_9718,N_8965,N_8476);
or U9719 (N_9719,N_8703,N_8478);
or U9720 (N_9720,N_8271,N_8794);
nand U9721 (N_9721,N_8701,N_8317);
and U9722 (N_9722,N_8816,N_8926);
or U9723 (N_9723,N_8529,N_8942);
nor U9724 (N_9724,N_8943,N_8938);
nor U9725 (N_9725,N_8614,N_8641);
xor U9726 (N_9726,N_8885,N_8998);
nor U9727 (N_9727,N_8838,N_8450);
nor U9728 (N_9728,N_8778,N_8839);
nor U9729 (N_9729,N_8605,N_8922);
nor U9730 (N_9730,N_8829,N_8952);
nor U9731 (N_9731,N_8920,N_8700);
and U9732 (N_9732,N_8715,N_8285);
and U9733 (N_9733,N_8932,N_8817);
or U9734 (N_9734,N_8804,N_8909);
or U9735 (N_9735,N_8515,N_8391);
and U9736 (N_9736,N_8308,N_8617);
nand U9737 (N_9737,N_8910,N_8609);
or U9738 (N_9738,N_8442,N_8307);
nor U9739 (N_9739,N_8947,N_8726);
or U9740 (N_9740,N_8722,N_8326);
or U9741 (N_9741,N_8911,N_8671);
and U9742 (N_9742,N_8355,N_8871);
xor U9743 (N_9743,N_8397,N_8981);
nor U9744 (N_9744,N_8938,N_8569);
xor U9745 (N_9745,N_8800,N_8792);
and U9746 (N_9746,N_8760,N_8607);
and U9747 (N_9747,N_8476,N_8488);
nand U9748 (N_9748,N_8822,N_8318);
and U9749 (N_9749,N_8280,N_8636);
nand U9750 (N_9750,N_9541,N_9409);
nor U9751 (N_9751,N_9280,N_9602);
or U9752 (N_9752,N_9289,N_9037);
xor U9753 (N_9753,N_9657,N_9012);
and U9754 (N_9754,N_9293,N_9006);
nand U9755 (N_9755,N_9318,N_9490);
or U9756 (N_9756,N_9587,N_9146);
nor U9757 (N_9757,N_9674,N_9390);
or U9758 (N_9758,N_9626,N_9458);
nor U9759 (N_9759,N_9089,N_9624);
nor U9760 (N_9760,N_9736,N_9655);
nand U9761 (N_9761,N_9447,N_9154);
or U9762 (N_9762,N_9034,N_9295);
xor U9763 (N_9763,N_9396,N_9322);
nor U9764 (N_9764,N_9005,N_9395);
or U9765 (N_9765,N_9579,N_9404);
nor U9766 (N_9766,N_9267,N_9671);
or U9767 (N_9767,N_9238,N_9584);
nor U9768 (N_9768,N_9177,N_9667);
and U9769 (N_9769,N_9506,N_9426);
nand U9770 (N_9770,N_9239,N_9328);
xor U9771 (N_9771,N_9697,N_9063);
or U9772 (N_9772,N_9670,N_9733);
and U9773 (N_9773,N_9611,N_9645);
xor U9774 (N_9774,N_9485,N_9469);
nand U9775 (N_9775,N_9100,N_9356);
nor U9776 (N_9776,N_9116,N_9616);
nor U9777 (N_9777,N_9140,N_9603);
xnor U9778 (N_9778,N_9588,N_9132);
xnor U9779 (N_9779,N_9539,N_9097);
and U9780 (N_9780,N_9263,N_9405);
nor U9781 (N_9781,N_9171,N_9118);
or U9782 (N_9782,N_9744,N_9481);
or U9783 (N_9783,N_9125,N_9323);
and U9784 (N_9784,N_9274,N_9149);
or U9785 (N_9785,N_9002,N_9739);
xor U9786 (N_9786,N_9462,N_9305);
nor U9787 (N_9787,N_9480,N_9716);
and U9788 (N_9788,N_9375,N_9082);
or U9789 (N_9789,N_9659,N_9373);
nand U9790 (N_9790,N_9186,N_9727);
nand U9791 (N_9791,N_9105,N_9438);
and U9792 (N_9792,N_9275,N_9181);
or U9793 (N_9793,N_9741,N_9261);
and U9794 (N_9794,N_9415,N_9158);
nor U9795 (N_9795,N_9530,N_9392);
nor U9796 (N_9796,N_9561,N_9141);
and U9797 (N_9797,N_9494,N_9211);
or U9798 (N_9798,N_9104,N_9350);
and U9799 (N_9799,N_9424,N_9368);
xnor U9800 (N_9800,N_9195,N_9291);
xor U9801 (N_9801,N_9669,N_9018);
or U9802 (N_9802,N_9151,N_9121);
nand U9803 (N_9803,N_9184,N_9115);
and U9804 (N_9804,N_9256,N_9362);
nand U9805 (N_9805,N_9507,N_9427);
xnor U9806 (N_9806,N_9203,N_9008);
and U9807 (N_9807,N_9155,N_9269);
and U9808 (N_9808,N_9348,N_9650);
nand U9809 (N_9809,N_9166,N_9060);
nor U9810 (N_9810,N_9529,N_9000);
nor U9811 (N_9811,N_9622,N_9287);
or U9812 (N_9812,N_9672,N_9712);
or U9813 (N_9813,N_9734,N_9600);
nand U9814 (N_9814,N_9509,N_9412);
and U9815 (N_9815,N_9482,N_9001);
and U9816 (N_9816,N_9586,N_9525);
xnor U9817 (N_9817,N_9505,N_9284);
nand U9818 (N_9818,N_9080,N_9581);
nor U9819 (N_9819,N_9229,N_9649);
nor U9820 (N_9820,N_9123,N_9208);
nor U9821 (N_9821,N_9073,N_9047);
nor U9822 (N_9822,N_9514,N_9519);
and U9823 (N_9823,N_9613,N_9064);
xor U9824 (N_9824,N_9095,N_9048);
nor U9825 (N_9825,N_9648,N_9457);
xnor U9826 (N_9826,N_9662,N_9283);
xnor U9827 (N_9827,N_9076,N_9567);
xnor U9828 (N_9828,N_9321,N_9425);
xnor U9829 (N_9829,N_9410,N_9596);
or U9830 (N_9830,N_9167,N_9190);
nor U9831 (N_9831,N_9407,N_9159);
nand U9832 (N_9832,N_9435,N_9175);
nand U9833 (N_9833,N_9306,N_9501);
xor U9834 (N_9834,N_9068,N_9109);
and U9835 (N_9835,N_9397,N_9017);
or U9836 (N_9836,N_9249,N_9067);
and U9837 (N_9837,N_9399,N_9465);
nor U9838 (N_9838,N_9666,N_9643);
nor U9839 (N_9839,N_9554,N_9294);
nand U9840 (N_9840,N_9244,N_9354);
nor U9841 (N_9841,N_9242,N_9710);
or U9842 (N_9842,N_9138,N_9575);
and U9843 (N_9843,N_9742,N_9654);
and U9844 (N_9844,N_9013,N_9271);
nand U9845 (N_9845,N_9041,N_9381);
nand U9846 (N_9846,N_9459,N_9349);
nand U9847 (N_9847,N_9248,N_9163);
and U9848 (N_9848,N_9050,N_9698);
xnor U9849 (N_9849,N_9147,N_9088);
nand U9850 (N_9850,N_9385,N_9593);
or U9851 (N_9851,N_9428,N_9389);
nor U9852 (N_9852,N_9487,N_9610);
or U9853 (N_9853,N_9168,N_9452);
nand U9854 (N_9854,N_9574,N_9464);
or U9855 (N_9855,N_9538,N_9056);
and U9856 (N_9856,N_9084,N_9338);
nor U9857 (N_9857,N_9236,N_9612);
nor U9858 (N_9858,N_9706,N_9441);
or U9859 (N_9859,N_9470,N_9502);
nand U9860 (N_9860,N_9433,N_9226);
or U9861 (N_9861,N_9548,N_9641);
nor U9862 (N_9862,N_9169,N_9255);
or U9863 (N_9863,N_9510,N_9573);
or U9864 (N_9864,N_9747,N_9339);
nor U9865 (N_9865,N_9374,N_9212);
nor U9866 (N_9866,N_9411,N_9165);
nand U9867 (N_9867,N_9652,N_9546);
nor U9868 (N_9868,N_9376,N_9243);
or U9869 (N_9869,N_9078,N_9679);
xor U9870 (N_9870,N_9331,N_9498);
nor U9871 (N_9871,N_9023,N_9137);
and U9872 (N_9872,N_9721,N_9044);
nand U9873 (N_9873,N_9194,N_9536);
nand U9874 (N_9874,N_9062,N_9454);
or U9875 (N_9875,N_9077,N_9150);
and U9876 (N_9876,N_9492,N_9673);
nor U9877 (N_9877,N_9199,N_9517);
nor U9878 (N_9878,N_9179,N_9352);
nand U9879 (N_9879,N_9206,N_9042);
and U9880 (N_9880,N_9552,N_9086);
or U9881 (N_9881,N_9631,N_9634);
or U9882 (N_9882,N_9038,N_9276);
and U9883 (N_9883,N_9508,N_9406);
and U9884 (N_9884,N_9033,N_9499);
nand U9885 (N_9885,N_9443,N_9707);
or U9886 (N_9886,N_9281,N_9491);
nand U9887 (N_9887,N_9401,N_9614);
or U9888 (N_9888,N_9647,N_9419);
or U9889 (N_9889,N_9156,N_9213);
nor U9890 (N_9890,N_9367,N_9134);
nor U9891 (N_9891,N_9442,N_9597);
and U9892 (N_9892,N_9675,N_9594);
or U9893 (N_9893,N_9282,N_9273);
xor U9894 (N_9894,N_9709,N_9545);
nor U9895 (N_9895,N_9504,N_9416);
nor U9896 (N_9896,N_9632,N_9639);
nor U9897 (N_9897,N_9476,N_9377);
nand U9898 (N_9898,N_9014,N_9730);
and U9899 (N_9899,N_9658,N_9052);
and U9900 (N_9900,N_9515,N_9093);
and U9901 (N_9901,N_9524,N_9319);
and U9902 (N_9902,N_9749,N_9025);
or U9903 (N_9903,N_9748,N_9101);
nor U9904 (N_9904,N_9259,N_9192);
nand U9905 (N_9905,N_9298,N_9430);
or U9906 (N_9906,N_9439,N_9345);
or U9907 (N_9907,N_9317,N_9364);
nand U9908 (N_9908,N_9591,N_9188);
and U9909 (N_9909,N_9043,N_9726);
nand U9910 (N_9910,N_9022,N_9224);
nand U9911 (N_9911,N_9534,N_9081);
nor U9912 (N_9912,N_9383,N_9260);
or U9913 (N_9913,N_9725,N_9153);
and U9914 (N_9914,N_9735,N_9031);
xnor U9915 (N_9915,N_9394,N_9526);
and U9916 (N_9916,N_9637,N_9705);
nor U9917 (N_9917,N_9531,N_9676);
xor U9918 (N_9918,N_9661,N_9329);
nor U9919 (N_9919,N_9098,N_9701);
nand U9920 (N_9920,N_9096,N_9182);
and U9921 (N_9921,N_9414,N_9142);
nor U9922 (N_9922,N_9562,N_9094);
or U9923 (N_9923,N_9262,N_9585);
nor U9924 (N_9924,N_9556,N_9286);
nand U9925 (N_9925,N_9209,N_9180);
nor U9926 (N_9926,N_9446,N_9173);
nand U9927 (N_9927,N_9126,N_9577);
nor U9928 (N_9928,N_9070,N_9051);
nor U9929 (N_9929,N_9359,N_9692);
nor U9930 (N_9930,N_9099,N_9592);
nor U9931 (N_9931,N_9049,N_9387);
and U9932 (N_9932,N_9265,N_9489);
and U9933 (N_9933,N_9161,N_9432);
nand U9934 (N_9934,N_9231,N_9344);
nor U9935 (N_9935,N_9668,N_9720);
nor U9936 (N_9936,N_9131,N_9440);
or U9937 (N_9937,N_9232,N_9589);
and U9938 (N_9938,N_9301,N_9746);
nor U9939 (N_9939,N_9120,N_9629);
nor U9940 (N_9940,N_9714,N_9472);
and U9941 (N_9941,N_9711,N_9638);
nand U9942 (N_9942,N_9028,N_9625);
nand U9943 (N_9943,N_9583,N_9431);
or U9944 (N_9944,N_9475,N_9054);
nor U9945 (N_9945,N_9026,N_9532);
and U9946 (N_9946,N_9136,N_9379);
nand U9947 (N_9947,N_9477,N_9691);
and U9948 (N_9948,N_9337,N_9633);
or U9949 (N_9949,N_9245,N_9237);
nand U9950 (N_9950,N_9145,N_9484);
nor U9951 (N_9951,N_9393,N_9718);
or U9952 (N_9952,N_9057,N_9066);
and U9953 (N_9953,N_9608,N_9087);
or U9954 (N_9954,N_9300,N_9421);
or U9955 (N_9955,N_9330,N_9324);
and U9956 (N_9956,N_9272,N_9467);
nand U9957 (N_9957,N_9170,N_9699);
nand U9958 (N_9958,N_9266,N_9664);
xnor U9959 (N_9959,N_9103,N_9320);
xor U9960 (N_9960,N_9717,N_9688);
xor U9961 (N_9961,N_9277,N_9240);
nand U9962 (N_9962,N_9576,N_9302);
and U9963 (N_9963,N_9113,N_9270);
or U9964 (N_9964,N_9032,N_9351);
nand U9965 (N_9965,N_9690,N_9370);
nand U9966 (N_9966,N_9106,N_9010);
and U9967 (N_9967,N_9299,N_9423);
or U9968 (N_9968,N_9055,N_9251);
nand U9969 (N_9969,N_9523,N_9656);
nand U9970 (N_9970,N_9011,N_9630);
nand U9971 (N_9971,N_9724,N_9450);
and U9972 (N_9972,N_9326,N_9559);
and U9973 (N_9973,N_9500,N_9316);
and U9974 (N_9974,N_9618,N_9537);
or U9975 (N_9975,N_9363,N_9029);
xnor U9976 (N_9976,N_9466,N_9285);
nand U9977 (N_9977,N_9402,N_9143);
nand U9978 (N_9978,N_9107,N_9478);
or U9979 (N_9979,N_9681,N_9111);
and U9980 (N_9980,N_9522,N_9495);
or U9981 (N_9981,N_9685,N_9388);
or U9982 (N_9982,N_9369,N_9327);
nor U9983 (N_9983,N_9564,N_9535);
nor U9984 (N_9984,N_9700,N_9148);
xor U9985 (N_9985,N_9549,N_9129);
nor U9986 (N_9986,N_9516,N_9292);
or U9987 (N_9987,N_9016,N_9391);
and U9988 (N_9988,N_9053,N_9024);
nor U9989 (N_9989,N_9743,N_9434);
or U9990 (N_9990,N_9448,N_9473);
nor U9991 (N_9991,N_9580,N_9468);
nand U9992 (N_9992,N_9220,N_9729);
or U9993 (N_9993,N_9197,N_9009);
nor U9994 (N_9994,N_9196,N_9738);
or U9995 (N_9995,N_9030,N_9160);
xnor U9996 (N_9996,N_9486,N_9451);
or U9997 (N_9997,N_9357,N_9644);
xnor U9998 (N_9998,N_9278,N_9418);
or U9999 (N_9999,N_9310,N_9740);
nor U10000 (N_10000,N_9663,N_9258);
and U10001 (N_10001,N_9544,N_9512);
and U10002 (N_10002,N_9214,N_9444);
nor U10003 (N_10003,N_9723,N_9533);
nand U10004 (N_10004,N_9039,N_9241);
nand U10005 (N_10005,N_9557,N_9445);
or U10006 (N_10006,N_9646,N_9193);
and U10007 (N_10007,N_9620,N_9313);
and U10008 (N_10008,N_9619,N_9378);
or U10009 (N_10009,N_9371,N_9615);
and U10010 (N_10010,N_9463,N_9071);
or U10011 (N_10011,N_9342,N_9550);
xnor U10012 (N_10012,N_9130,N_9069);
or U10013 (N_10013,N_9004,N_9380);
nand U10014 (N_10014,N_9595,N_9225);
and U10015 (N_10015,N_9527,N_9198);
or U10016 (N_10016,N_9413,N_9606);
or U10017 (N_10017,N_9221,N_9015);
nor U10018 (N_10018,N_9623,N_9601);
or U10019 (N_10019,N_9704,N_9483);
nor U10020 (N_10020,N_9164,N_9311);
nor U10021 (N_10021,N_9687,N_9127);
and U10022 (N_10022,N_9621,N_9046);
and U10023 (N_10023,N_9566,N_9400);
nor U10024 (N_10024,N_9021,N_9122);
or U10025 (N_10025,N_9112,N_9455);
nand U10026 (N_10026,N_9511,N_9636);
xnor U10027 (N_10027,N_9437,N_9335);
nor U10028 (N_10028,N_9117,N_9075);
or U10029 (N_10029,N_9230,N_9253);
nand U10030 (N_10030,N_9223,N_9449);
nor U10031 (N_10031,N_9341,N_9684);
nor U10032 (N_10032,N_9702,N_9040);
and U10033 (N_10033,N_9713,N_9560);
nor U10034 (N_10034,N_9366,N_9290);
xnor U10035 (N_10035,N_9653,N_9607);
nor U10036 (N_10036,N_9185,N_9569);
or U10037 (N_10037,N_9119,N_9540);
nor U10038 (N_10038,N_9635,N_9264);
and U10039 (N_10039,N_9547,N_9570);
nand U10040 (N_10040,N_9372,N_9058);
and U10041 (N_10041,N_9315,N_9382);
nand U10042 (N_10042,N_9157,N_9558);
or U10043 (N_10043,N_9235,N_9027);
or U10044 (N_10044,N_9139,N_9219);
nor U10045 (N_10045,N_9542,N_9346);
nor U10046 (N_10046,N_9496,N_9204);
and U10047 (N_10047,N_9355,N_9471);
and U10048 (N_10048,N_9628,N_9340);
xnor U10049 (N_10049,N_9128,N_9133);
or U10050 (N_10050,N_9202,N_9178);
nand U10051 (N_10051,N_9218,N_9110);
and U10052 (N_10052,N_9617,N_9360);
nand U10053 (N_10053,N_9719,N_9217);
xnor U10054 (N_10054,N_9144,N_9497);
nand U10055 (N_10055,N_9247,N_9246);
nand U10056 (N_10056,N_9061,N_9172);
nor U10057 (N_10057,N_9312,N_9257);
nor U10058 (N_10058,N_9090,N_9114);
or U10059 (N_10059,N_9677,N_9191);
nor U10060 (N_10060,N_9518,N_9083);
nand U10061 (N_10061,N_9553,N_9201);
or U10062 (N_10062,N_9059,N_9488);
and U10063 (N_10063,N_9200,N_9215);
xnor U10064 (N_10064,N_9461,N_9353);
nand U10065 (N_10065,N_9332,N_9436);
and U10066 (N_10066,N_9689,N_9660);
nor U10067 (N_10067,N_9722,N_9429);
or U10068 (N_10068,N_9309,N_9227);
xor U10069 (N_10069,N_9314,N_9715);
nor U10070 (N_10070,N_9108,N_9565);
nand U10071 (N_10071,N_9696,N_9403);
xor U10072 (N_10072,N_9543,N_9358);
xor U10073 (N_10073,N_9279,N_9693);
nor U10074 (N_10074,N_9325,N_9640);
xor U10075 (N_10075,N_9065,N_9187);
and U10076 (N_10076,N_9474,N_9605);
or U10077 (N_10077,N_9745,N_9604);
nand U10078 (N_10078,N_9555,N_9503);
nand U10079 (N_10079,N_9408,N_9453);
or U10080 (N_10080,N_9189,N_9420);
or U10081 (N_10081,N_9020,N_9079);
nand U10082 (N_10082,N_9695,N_9456);
nand U10083 (N_10083,N_9365,N_9520);
or U10084 (N_10084,N_9642,N_9683);
xnor U10085 (N_10085,N_9234,N_9091);
or U10086 (N_10086,N_9578,N_9678);
nand U10087 (N_10087,N_9609,N_9228);
xnor U10088 (N_10088,N_9651,N_9568);
nand U10089 (N_10089,N_9493,N_9124);
nor U10090 (N_10090,N_9398,N_9563);
nand U10091 (N_10091,N_9268,N_9361);
and U10092 (N_10092,N_9092,N_9422);
or U10093 (N_10093,N_9072,N_9176);
or U10094 (N_10094,N_9085,N_9333);
nor U10095 (N_10095,N_9207,N_9304);
and U10096 (N_10096,N_9035,N_9288);
nor U10097 (N_10097,N_9162,N_9135);
or U10098 (N_10098,N_9174,N_9731);
and U10099 (N_10099,N_9045,N_9551);
nor U10100 (N_10100,N_9074,N_9036);
nand U10101 (N_10101,N_9296,N_9152);
or U10102 (N_10102,N_9528,N_9708);
or U10103 (N_10103,N_9347,N_9205);
or U10104 (N_10104,N_9336,N_9007);
nor U10105 (N_10105,N_9665,N_9582);
or U10106 (N_10106,N_9216,N_9222);
nand U10107 (N_10107,N_9307,N_9694);
and U10108 (N_10108,N_9728,N_9384);
or U10109 (N_10109,N_9252,N_9460);
nor U10110 (N_10110,N_9003,N_9572);
and U10111 (N_10111,N_9417,N_9019);
or U10112 (N_10112,N_9571,N_9598);
nand U10113 (N_10113,N_9686,N_9513);
or U10114 (N_10114,N_9102,N_9308);
nor U10115 (N_10115,N_9343,N_9732);
xnor U10116 (N_10116,N_9479,N_9210);
xor U10117 (N_10117,N_9297,N_9680);
and U10118 (N_10118,N_9682,N_9737);
or U10119 (N_10119,N_9627,N_9254);
and U10120 (N_10120,N_9386,N_9703);
or U10121 (N_10121,N_9183,N_9334);
nand U10122 (N_10122,N_9250,N_9590);
and U10123 (N_10123,N_9303,N_9233);
or U10124 (N_10124,N_9599,N_9521);
nor U10125 (N_10125,N_9038,N_9125);
and U10126 (N_10126,N_9354,N_9613);
or U10127 (N_10127,N_9143,N_9211);
and U10128 (N_10128,N_9309,N_9423);
nand U10129 (N_10129,N_9607,N_9465);
and U10130 (N_10130,N_9428,N_9495);
xor U10131 (N_10131,N_9036,N_9522);
nor U10132 (N_10132,N_9715,N_9551);
nor U10133 (N_10133,N_9157,N_9364);
and U10134 (N_10134,N_9712,N_9182);
nand U10135 (N_10135,N_9276,N_9222);
or U10136 (N_10136,N_9556,N_9512);
and U10137 (N_10137,N_9737,N_9513);
nor U10138 (N_10138,N_9533,N_9177);
or U10139 (N_10139,N_9654,N_9020);
and U10140 (N_10140,N_9175,N_9038);
nand U10141 (N_10141,N_9143,N_9452);
nor U10142 (N_10142,N_9171,N_9085);
xor U10143 (N_10143,N_9059,N_9109);
or U10144 (N_10144,N_9183,N_9587);
or U10145 (N_10145,N_9042,N_9609);
nor U10146 (N_10146,N_9310,N_9518);
nand U10147 (N_10147,N_9073,N_9505);
nand U10148 (N_10148,N_9190,N_9427);
or U10149 (N_10149,N_9423,N_9378);
nor U10150 (N_10150,N_9485,N_9449);
nand U10151 (N_10151,N_9550,N_9302);
nand U10152 (N_10152,N_9506,N_9730);
nand U10153 (N_10153,N_9491,N_9684);
or U10154 (N_10154,N_9189,N_9563);
and U10155 (N_10155,N_9105,N_9240);
nor U10156 (N_10156,N_9749,N_9211);
or U10157 (N_10157,N_9309,N_9166);
and U10158 (N_10158,N_9287,N_9500);
nand U10159 (N_10159,N_9607,N_9308);
nor U10160 (N_10160,N_9341,N_9105);
or U10161 (N_10161,N_9697,N_9281);
nand U10162 (N_10162,N_9650,N_9123);
and U10163 (N_10163,N_9596,N_9715);
nand U10164 (N_10164,N_9396,N_9633);
or U10165 (N_10165,N_9219,N_9271);
and U10166 (N_10166,N_9387,N_9390);
xor U10167 (N_10167,N_9061,N_9446);
nor U10168 (N_10168,N_9059,N_9465);
nand U10169 (N_10169,N_9200,N_9174);
nor U10170 (N_10170,N_9432,N_9231);
nand U10171 (N_10171,N_9589,N_9678);
and U10172 (N_10172,N_9301,N_9254);
or U10173 (N_10173,N_9367,N_9515);
nor U10174 (N_10174,N_9700,N_9267);
and U10175 (N_10175,N_9390,N_9339);
and U10176 (N_10176,N_9584,N_9343);
nand U10177 (N_10177,N_9103,N_9264);
and U10178 (N_10178,N_9365,N_9284);
nand U10179 (N_10179,N_9596,N_9683);
and U10180 (N_10180,N_9289,N_9403);
and U10181 (N_10181,N_9601,N_9739);
nand U10182 (N_10182,N_9447,N_9238);
and U10183 (N_10183,N_9383,N_9495);
nor U10184 (N_10184,N_9468,N_9639);
and U10185 (N_10185,N_9609,N_9447);
nor U10186 (N_10186,N_9265,N_9107);
and U10187 (N_10187,N_9159,N_9094);
nor U10188 (N_10188,N_9186,N_9333);
nor U10189 (N_10189,N_9112,N_9647);
or U10190 (N_10190,N_9610,N_9179);
and U10191 (N_10191,N_9269,N_9120);
and U10192 (N_10192,N_9577,N_9018);
and U10193 (N_10193,N_9102,N_9035);
nand U10194 (N_10194,N_9529,N_9319);
xnor U10195 (N_10195,N_9260,N_9480);
and U10196 (N_10196,N_9069,N_9011);
nand U10197 (N_10197,N_9074,N_9461);
or U10198 (N_10198,N_9580,N_9022);
nand U10199 (N_10199,N_9091,N_9705);
and U10200 (N_10200,N_9156,N_9545);
xnor U10201 (N_10201,N_9498,N_9404);
nand U10202 (N_10202,N_9485,N_9197);
or U10203 (N_10203,N_9681,N_9045);
or U10204 (N_10204,N_9077,N_9535);
or U10205 (N_10205,N_9431,N_9204);
and U10206 (N_10206,N_9725,N_9618);
and U10207 (N_10207,N_9440,N_9062);
nand U10208 (N_10208,N_9028,N_9466);
xor U10209 (N_10209,N_9331,N_9547);
or U10210 (N_10210,N_9590,N_9075);
nor U10211 (N_10211,N_9642,N_9081);
and U10212 (N_10212,N_9427,N_9413);
nor U10213 (N_10213,N_9342,N_9637);
nand U10214 (N_10214,N_9600,N_9554);
or U10215 (N_10215,N_9748,N_9447);
xnor U10216 (N_10216,N_9239,N_9615);
nor U10217 (N_10217,N_9208,N_9302);
nor U10218 (N_10218,N_9273,N_9369);
nor U10219 (N_10219,N_9611,N_9017);
or U10220 (N_10220,N_9264,N_9709);
or U10221 (N_10221,N_9075,N_9173);
nand U10222 (N_10222,N_9257,N_9309);
or U10223 (N_10223,N_9728,N_9382);
nand U10224 (N_10224,N_9453,N_9387);
nor U10225 (N_10225,N_9077,N_9609);
nor U10226 (N_10226,N_9572,N_9339);
or U10227 (N_10227,N_9503,N_9648);
nand U10228 (N_10228,N_9012,N_9165);
and U10229 (N_10229,N_9542,N_9599);
and U10230 (N_10230,N_9725,N_9557);
nand U10231 (N_10231,N_9146,N_9404);
nand U10232 (N_10232,N_9013,N_9278);
and U10233 (N_10233,N_9251,N_9024);
or U10234 (N_10234,N_9162,N_9282);
nor U10235 (N_10235,N_9435,N_9656);
or U10236 (N_10236,N_9481,N_9537);
and U10237 (N_10237,N_9158,N_9510);
and U10238 (N_10238,N_9167,N_9501);
nor U10239 (N_10239,N_9062,N_9106);
nand U10240 (N_10240,N_9166,N_9451);
nand U10241 (N_10241,N_9339,N_9250);
xnor U10242 (N_10242,N_9281,N_9679);
and U10243 (N_10243,N_9035,N_9587);
nor U10244 (N_10244,N_9618,N_9527);
and U10245 (N_10245,N_9055,N_9573);
or U10246 (N_10246,N_9711,N_9636);
nor U10247 (N_10247,N_9467,N_9105);
or U10248 (N_10248,N_9168,N_9260);
and U10249 (N_10249,N_9034,N_9093);
nor U10250 (N_10250,N_9143,N_9413);
nor U10251 (N_10251,N_9613,N_9380);
and U10252 (N_10252,N_9213,N_9572);
nand U10253 (N_10253,N_9744,N_9377);
nor U10254 (N_10254,N_9054,N_9403);
or U10255 (N_10255,N_9740,N_9543);
and U10256 (N_10256,N_9358,N_9446);
nand U10257 (N_10257,N_9476,N_9570);
or U10258 (N_10258,N_9229,N_9109);
and U10259 (N_10259,N_9245,N_9100);
nor U10260 (N_10260,N_9494,N_9550);
nor U10261 (N_10261,N_9456,N_9235);
nand U10262 (N_10262,N_9242,N_9417);
or U10263 (N_10263,N_9314,N_9222);
or U10264 (N_10264,N_9614,N_9044);
and U10265 (N_10265,N_9147,N_9524);
nand U10266 (N_10266,N_9257,N_9283);
or U10267 (N_10267,N_9544,N_9345);
or U10268 (N_10268,N_9025,N_9623);
and U10269 (N_10269,N_9502,N_9523);
or U10270 (N_10270,N_9215,N_9408);
or U10271 (N_10271,N_9133,N_9188);
or U10272 (N_10272,N_9266,N_9611);
nor U10273 (N_10273,N_9273,N_9638);
and U10274 (N_10274,N_9231,N_9387);
xnor U10275 (N_10275,N_9572,N_9139);
nor U10276 (N_10276,N_9571,N_9005);
nor U10277 (N_10277,N_9265,N_9558);
or U10278 (N_10278,N_9034,N_9646);
nand U10279 (N_10279,N_9247,N_9507);
xnor U10280 (N_10280,N_9604,N_9500);
nor U10281 (N_10281,N_9300,N_9088);
nand U10282 (N_10282,N_9430,N_9123);
and U10283 (N_10283,N_9047,N_9125);
nor U10284 (N_10284,N_9451,N_9732);
and U10285 (N_10285,N_9676,N_9210);
and U10286 (N_10286,N_9221,N_9247);
and U10287 (N_10287,N_9317,N_9649);
xnor U10288 (N_10288,N_9309,N_9374);
or U10289 (N_10289,N_9447,N_9531);
and U10290 (N_10290,N_9514,N_9464);
nand U10291 (N_10291,N_9734,N_9133);
or U10292 (N_10292,N_9320,N_9156);
xnor U10293 (N_10293,N_9599,N_9420);
nor U10294 (N_10294,N_9615,N_9391);
and U10295 (N_10295,N_9194,N_9094);
or U10296 (N_10296,N_9047,N_9142);
nor U10297 (N_10297,N_9105,N_9741);
and U10298 (N_10298,N_9037,N_9658);
xnor U10299 (N_10299,N_9524,N_9037);
nor U10300 (N_10300,N_9226,N_9565);
nand U10301 (N_10301,N_9354,N_9071);
or U10302 (N_10302,N_9728,N_9639);
and U10303 (N_10303,N_9432,N_9110);
nand U10304 (N_10304,N_9545,N_9272);
or U10305 (N_10305,N_9411,N_9696);
or U10306 (N_10306,N_9368,N_9294);
xnor U10307 (N_10307,N_9329,N_9209);
nor U10308 (N_10308,N_9219,N_9493);
nor U10309 (N_10309,N_9348,N_9729);
xnor U10310 (N_10310,N_9057,N_9432);
and U10311 (N_10311,N_9046,N_9200);
or U10312 (N_10312,N_9381,N_9316);
nor U10313 (N_10313,N_9477,N_9148);
nor U10314 (N_10314,N_9532,N_9515);
and U10315 (N_10315,N_9003,N_9198);
and U10316 (N_10316,N_9222,N_9252);
or U10317 (N_10317,N_9426,N_9184);
nor U10318 (N_10318,N_9130,N_9247);
or U10319 (N_10319,N_9552,N_9429);
nand U10320 (N_10320,N_9348,N_9704);
and U10321 (N_10321,N_9395,N_9308);
or U10322 (N_10322,N_9350,N_9028);
or U10323 (N_10323,N_9188,N_9060);
or U10324 (N_10324,N_9192,N_9572);
nand U10325 (N_10325,N_9376,N_9017);
or U10326 (N_10326,N_9412,N_9575);
nand U10327 (N_10327,N_9619,N_9616);
nor U10328 (N_10328,N_9344,N_9025);
nand U10329 (N_10329,N_9078,N_9090);
or U10330 (N_10330,N_9068,N_9563);
and U10331 (N_10331,N_9227,N_9300);
or U10332 (N_10332,N_9633,N_9305);
nand U10333 (N_10333,N_9533,N_9463);
nand U10334 (N_10334,N_9715,N_9124);
xor U10335 (N_10335,N_9491,N_9159);
and U10336 (N_10336,N_9491,N_9487);
nand U10337 (N_10337,N_9207,N_9245);
nand U10338 (N_10338,N_9110,N_9728);
nand U10339 (N_10339,N_9190,N_9322);
nand U10340 (N_10340,N_9670,N_9714);
or U10341 (N_10341,N_9565,N_9554);
nor U10342 (N_10342,N_9284,N_9291);
nor U10343 (N_10343,N_9466,N_9404);
xnor U10344 (N_10344,N_9037,N_9261);
and U10345 (N_10345,N_9147,N_9391);
nand U10346 (N_10346,N_9134,N_9527);
and U10347 (N_10347,N_9172,N_9239);
nor U10348 (N_10348,N_9222,N_9251);
or U10349 (N_10349,N_9479,N_9143);
and U10350 (N_10350,N_9672,N_9420);
xnor U10351 (N_10351,N_9746,N_9076);
and U10352 (N_10352,N_9623,N_9161);
nand U10353 (N_10353,N_9136,N_9609);
and U10354 (N_10354,N_9389,N_9320);
xor U10355 (N_10355,N_9469,N_9664);
xnor U10356 (N_10356,N_9245,N_9471);
or U10357 (N_10357,N_9258,N_9105);
nand U10358 (N_10358,N_9193,N_9617);
xor U10359 (N_10359,N_9243,N_9304);
nor U10360 (N_10360,N_9447,N_9630);
nor U10361 (N_10361,N_9628,N_9305);
nand U10362 (N_10362,N_9339,N_9040);
and U10363 (N_10363,N_9407,N_9066);
nand U10364 (N_10364,N_9642,N_9400);
and U10365 (N_10365,N_9266,N_9219);
xnor U10366 (N_10366,N_9260,N_9616);
xor U10367 (N_10367,N_9324,N_9293);
nor U10368 (N_10368,N_9704,N_9411);
or U10369 (N_10369,N_9263,N_9516);
nand U10370 (N_10370,N_9293,N_9700);
or U10371 (N_10371,N_9606,N_9496);
nand U10372 (N_10372,N_9038,N_9192);
nor U10373 (N_10373,N_9147,N_9264);
and U10374 (N_10374,N_9093,N_9611);
nor U10375 (N_10375,N_9218,N_9183);
nor U10376 (N_10376,N_9356,N_9730);
nor U10377 (N_10377,N_9024,N_9073);
nand U10378 (N_10378,N_9682,N_9705);
xor U10379 (N_10379,N_9194,N_9236);
and U10380 (N_10380,N_9405,N_9077);
nand U10381 (N_10381,N_9727,N_9540);
nand U10382 (N_10382,N_9216,N_9619);
and U10383 (N_10383,N_9573,N_9644);
nor U10384 (N_10384,N_9269,N_9727);
nand U10385 (N_10385,N_9359,N_9025);
nand U10386 (N_10386,N_9518,N_9425);
nor U10387 (N_10387,N_9155,N_9663);
nand U10388 (N_10388,N_9314,N_9001);
and U10389 (N_10389,N_9322,N_9000);
and U10390 (N_10390,N_9516,N_9049);
or U10391 (N_10391,N_9248,N_9326);
and U10392 (N_10392,N_9150,N_9036);
nor U10393 (N_10393,N_9731,N_9655);
xnor U10394 (N_10394,N_9585,N_9244);
nand U10395 (N_10395,N_9473,N_9088);
nand U10396 (N_10396,N_9175,N_9717);
and U10397 (N_10397,N_9001,N_9709);
nor U10398 (N_10398,N_9724,N_9496);
nand U10399 (N_10399,N_9181,N_9043);
and U10400 (N_10400,N_9509,N_9145);
or U10401 (N_10401,N_9666,N_9316);
and U10402 (N_10402,N_9036,N_9255);
nor U10403 (N_10403,N_9208,N_9719);
nand U10404 (N_10404,N_9326,N_9563);
nand U10405 (N_10405,N_9074,N_9644);
and U10406 (N_10406,N_9194,N_9602);
nor U10407 (N_10407,N_9531,N_9359);
nor U10408 (N_10408,N_9653,N_9083);
nor U10409 (N_10409,N_9372,N_9666);
xnor U10410 (N_10410,N_9422,N_9588);
and U10411 (N_10411,N_9052,N_9170);
xnor U10412 (N_10412,N_9363,N_9043);
nor U10413 (N_10413,N_9189,N_9268);
nor U10414 (N_10414,N_9092,N_9435);
nand U10415 (N_10415,N_9644,N_9219);
or U10416 (N_10416,N_9286,N_9557);
and U10417 (N_10417,N_9276,N_9181);
nand U10418 (N_10418,N_9514,N_9477);
nor U10419 (N_10419,N_9420,N_9596);
nand U10420 (N_10420,N_9579,N_9232);
or U10421 (N_10421,N_9254,N_9256);
or U10422 (N_10422,N_9171,N_9377);
and U10423 (N_10423,N_9133,N_9599);
nand U10424 (N_10424,N_9419,N_9611);
nor U10425 (N_10425,N_9517,N_9612);
nand U10426 (N_10426,N_9637,N_9360);
nand U10427 (N_10427,N_9530,N_9421);
xnor U10428 (N_10428,N_9221,N_9405);
nor U10429 (N_10429,N_9137,N_9682);
and U10430 (N_10430,N_9016,N_9425);
nand U10431 (N_10431,N_9028,N_9299);
nor U10432 (N_10432,N_9196,N_9442);
nor U10433 (N_10433,N_9598,N_9103);
and U10434 (N_10434,N_9142,N_9256);
nand U10435 (N_10435,N_9083,N_9143);
nor U10436 (N_10436,N_9346,N_9242);
nand U10437 (N_10437,N_9614,N_9246);
xor U10438 (N_10438,N_9578,N_9533);
or U10439 (N_10439,N_9553,N_9575);
or U10440 (N_10440,N_9626,N_9635);
xnor U10441 (N_10441,N_9223,N_9550);
nand U10442 (N_10442,N_9156,N_9285);
nand U10443 (N_10443,N_9555,N_9551);
nor U10444 (N_10444,N_9314,N_9252);
nand U10445 (N_10445,N_9538,N_9646);
nor U10446 (N_10446,N_9136,N_9466);
nand U10447 (N_10447,N_9377,N_9430);
xnor U10448 (N_10448,N_9715,N_9627);
xnor U10449 (N_10449,N_9182,N_9347);
and U10450 (N_10450,N_9638,N_9698);
and U10451 (N_10451,N_9056,N_9591);
nor U10452 (N_10452,N_9239,N_9229);
xnor U10453 (N_10453,N_9468,N_9311);
or U10454 (N_10454,N_9625,N_9379);
or U10455 (N_10455,N_9151,N_9352);
nand U10456 (N_10456,N_9206,N_9460);
or U10457 (N_10457,N_9003,N_9511);
nand U10458 (N_10458,N_9421,N_9379);
or U10459 (N_10459,N_9313,N_9438);
nand U10460 (N_10460,N_9153,N_9733);
and U10461 (N_10461,N_9134,N_9465);
nand U10462 (N_10462,N_9711,N_9466);
or U10463 (N_10463,N_9159,N_9598);
or U10464 (N_10464,N_9290,N_9052);
nor U10465 (N_10465,N_9412,N_9242);
nor U10466 (N_10466,N_9575,N_9370);
nor U10467 (N_10467,N_9333,N_9609);
or U10468 (N_10468,N_9049,N_9532);
or U10469 (N_10469,N_9575,N_9161);
and U10470 (N_10470,N_9543,N_9452);
and U10471 (N_10471,N_9385,N_9117);
nor U10472 (N_10472,N_9125,N_9255);
or U10473 (N_10473,N_9350,N_9198);
nand U10474 (N_10474,N_9641,N_9382);
nand U10475 (N_10475,N_9563,N_9044);
nand U10476 (N_10476,N_9385,N_9686);
nor U10477 (N_10477,N_9696,N_9565);
and U10478 (N_10478,N_9484,N_9326);
nand U10479 (N_10479,N_9285,N_9266);
nand U10480 (N_10480,N_9332,N_9017);
or U10481 (N_10481,N_9121,N_9347);
nor U10482 (N_10482,N_9383,N_9225);
nor U10483 (N_10483,N_9175,N_9267);
xnor U10484 (N_10484,N_9483,N_9268);
xnor U10485 (N_10485,N_9081,N_9583);
nor U10486 (N_10486,N_9456,N_9458);
or U10487 (N_10487,N_9105,N_9127);
and U10488 (N_10488,N_9670,N_9661);
or U10489 (N_10489,N_9483,N_9337);
or U10490 (N_10490,N_9512,N_9245);
nor U10491 (N_10491,N_9733,N_9575);
and U10492 (N_10492,N_9530,N_9080);
and U10493 (N_10493,N_9709,N_9025);
and U10494 (N_10494,N_9246,N_9393);
and U10495 (N_10495,N_9195,N_9253);
or U10496 (N_10496,N_9106,N_9108);
nor U10497 (N_10497,N_9155,N_9456);
nor U10498 (N_10498,N_9704,N_9187);
xor U10499 (N_10499,N_9478,N_9149);
xnor U10500 (N_10500,N_9944,N_9955);
and U10501 (N_10501,N_10142,N_10462);
or U10502 (N_10502,N_10112,N_9770);
nand U10503 (N_10503,N_9997,N_10450);
nor U10504 (N_10504,N_10293,N_10147);
or U10505 (N_10505,N_10086,N_10113);
nand U10506 (N_10506,N_10138,N_10110);
or U10507 (N_10507,N_9882,N_10277);
nor U10508 (N_10508,N_10184,N_10245);
and U10509 (N_10509,N_10382,N_9918);
and U10510 (N_10510,N_10210,N_9848);
or U10511 (N_10511,N_9982,N_9755);
or U10512 (N_10512,N_10349,N_10451);
or U10513 (N_10513,N_10129,N_10287);
nor U10514 (N_10514,N_9990,N_10009);
and U10515 (N_10515,N_10188,N_10356);
nand U10516 (N_10516,N_10226,N_9920);
nor U10517 (N_10517,N_10411,N_10442);
or U10518 (N_10518,N_10056,N_9949);
or U10519 (N_10519,N_10099,N_10313);
nor U10520 (N_10520,N_10433,N_10047);
nand U10521 (N_10521,N_10141,N_10120);
nand U10522 (N_10522,N_10082,N_10085);
nor U10523 (N_10523,N_10397,N_9909);
or U10524 (N_10524,N_9901,N_10381);
and U10525 (N_10525,N_10385,N_10322);
or U10526 (N_10526,N_10211,N_10280);
and U10527 (N_10527,N_9912,N_10107);
and U10528 (N_10528,N_10027,N_10288);
nor U10529 (N_10529,N_10464,N_10380);
or U10530 (N_10530,N_9974,N_9972);
nand U10531 (N_10531,N_10285,N_10236);
and U10532 (N_10532,N_10209,N_10109);
and U10533 (N_10533,N_9831,N_9847);
or U10534 (N_10534,N_9753,N_10376);
xnor U10535 (N_10535,N_9858,N_10020);
and U10536 (N_10536,N_9813,N_10241);
or U10537 (N_10537,N_9981,N_9815);
or U10538 (N_10538,N_10488,N_10386);
or U10539 (N_10539,N_10067,N_10041);
and U10540 (N_10540,N_10190,N_9807);
nor U10541 (N_10541,N_9797,N_10263);
nor U10542 (N_10542,N_10365,N_10319);
and U10543 (N_10543,N_10444,N_10072);
or U10544 (N_10544,N_9766,N_10471);
nand U10545 (N_10545,N_10206,N_10203);
and U10546 (N_10546,N_10253,N_9934);
or U10547 (N_10547,N_10266,N_9860);
and U10548 (N_10548,N_9841,N_10205);
nand U10549 (N_10549,N_10435,N_9895);
nand U10550 (N_10550,N_10437,N_10182);
and U10551 (N_10551,N_9925,N_10183);
nand U10552 (N_10552,N_10102,N_9965);
xor U10553 (N_10553,N_10005,N_10428);
and U10554 (N_10554,N_10157,N_9854);
nand U10555 (N_10555,N_9919,N_10318);
nand U10556 (N_10556,N_10195,N_10219);
nand U10557 (N_10557,N_10048,N_10491);
nand U10558 (N_10558,N_9810,N_10031);
and U10559 (N_10559,N_10425,N_10060);
xor U10560 (N_10560,N_9796,N_10242);
nor U10561 (N_10561,N_10248,N_10191);
nor U10562 (N_10562,N_9889,N_9906);
nand U10563 (N_10563,N_10216,N_10459);
nand U10564 (N_10564,N_10101,N_10370);
or U10565 (N_10565,N_10057,N_10292);
or U10566 (N_10566,N_10323,N_10493);
nand U10567 (N_10567,N_10391,N_9885);
and U10568 (N_10568,N_10221,N_9870);
nand U10569 (N_10569,N_9768,N_10460);
nand U10570 (N_10570,N_10383,N_10126);
or U10571 (N_10571,N_9904,N_10273);
and U10572 (N_10572,N_9887,N_10472);
nor U10573 (N_10573,N_9838,N_10324);
nand U10574 (N_10574,N_10494,N_10423);
nand U10575 (N_10575,N_10247,N_9952);
xor U10576 (N_10576,N_10496,N_10125);
nand U10577 (N_10577,N_10390,N_9843);
or U10578 (N_10578,N_10244,N_10469);
xor U10579 (N_10579,N_9933,N_10497);
nand U10580 (N_10580,N_10062,N_9792);
or U10581 (N_10581,N_9794,N_9940);
nand U10582 (N_10582,N_10478,N_10044);
nand U10583 (N_10583,N_10164,N_9868);
nand U10584 (N_10584,N_9822,N_10064);
nor U10585 (N_10585,N_10095,N_10305);
nand U10586 (N_10586,N_10137,N_9855);
nor U10587 (N_10587,N_9964,N_10066);
and U10588 (N_10588,N_9975,N_10418);
nor U10589 (N_10589,N_10132,N_9908);
nor U10590 (N_10590,N_9902,N_10368);
nor U10591 (N_10591,N_9820,N_9899);
nor U10592 (N_10592,N_10345,N_10130);
and U10593 (N_10593,N_10202,N_9968);
nand U10594 (N_10594,N_10021,N_10022);
or U10595 (N_10595,N_10078,N_9872);
nand U10596 (N_10596,N_10140,N_9951);
xor U10597 (N_10597,N_9988,N_10363);
and U10598 (N_10598,N_10177,N_9754);
nand U10599 (N_10599,N_10414,N_9994);
or U10600 (N_10600,N_10467,N_10108);
xnor U10601 (N_10601,N_10269,N_10456);
xnor U10602 (N_10602,N_10474,N_9782);
nand U10603 (N_10603,N_9913,N_9845);
nor U10604 (N_10604,N_10149,N_10036);
or U10605 (N_10605,N_10260,N_9916);
nor U10606 (N_10606,N_10198,N_9957);
and U10607 (N_10607,N_9846,N_9978);
or U10608 (N_10608,N_10161,N_10420);
nand U10609 (N_10609,N_9874,N_10301);
and U10610 (N_10610,N_10134,N_9837);
nor U10611 (N_10611,N_10443,N_10025);
nor U10612 (N_10612,N_9996,N_10401);
or U10613 (N_10613,N_10194,N_10001);
nor U10614 (N_10614,N_10052,N_10336);
or U10615 (N_10615,N_10410,N_10295);
xnor U10616 (N_10616,N_10321,N_9926);
nor U10617 (N_10617,N_10393,N_10454);
and U10618 (N_10618,N_10002,N_10154);
nor U10619 (N_10619,N_10343,N_9824);
and U10620 (N_10620,N_9921,N_10333);
nor U10621 (N_10621,N_9928,N_9750);
and U10622 (N_10622,N_10360,N_9773);
nand U10623 (N_10623,N_9842,N_10495);
nand U10624 (N_10624,N_9938,N_10104);
and U10625 (N_10625,N_9900,N_10475);
and U10626 (N_10626,N_9832,N_9853);
nor U10627 (N_10627,N_10463,N_10042);
and U10628 (N_10628,N_9941,N_10215);
and U10629 (N_10629,N_10178,N_9776);
nor U10630 (N_10630,N_10094,N_10276);
xor U10631 (N_10631,N_10374,N_10071);
or U10632 (N_10632,N_10290,N_10254);
or U10633 (N_10633,N_9771,N_10186);
or U10634 (N_10634,N_10337,N_10417);
and U10635 (N_10635,N_10004,N_10372);
nand U10636 (N_10636,N_9799,N_10201);
nor U10637 (N_10637,N_10426,N_10235);
or U10638 (N_10638,N_9759,N_10026);
and U10639 (N_10639,N_10053,N_9775);
nor U10640 (N_10640,N_9945,N_10232);
nor U10641 (N_10641,N_10268,N_10144);
xor U10642 (N_10642,N_10421,N_10065);
nor U10643 (N_10643,N_9819,N_10077);
and U10644 (N_10644,N_9893,N_10334);
or U10645 (N_10645,N_10175,N_10058);
or U10646 (N_10646,N_9783,N_9953);
nor U10647 (N_10647,N_10388,N_10088);
nand U10648 (N_10648,N_10402,N_10106);
and U10649 (N_10649,N_10124,N_10220);
nor U10650 (N_10650,N_10392,N_10278);
nor U10651 (N_10651,N_9769,N_10430);
or U10652 (N_10652,N_9856,N_10196);
and U10653 (N_10653,N_9956,N_10006);
and U10654 (N_10654,N_9786,N_10274);
and U10655 (N_10655,N_9795,N_9939);
and U10656 (N_10656,N_9762,N_9894);
nor U10657 (N_10657,N_10424,N_9806);
nand U10658 (N_10658,N_9798,N_10340);
nor U10659 (N_10659,N_10013,N_10373);
or U10660 (N_10660,N_9781,N_9930);
nor U10661 (N_10661,N_10117,N_10146);
nand U10662 (N_10662,N_10148,N_10302);
nor U10663 (N_10663,N_10181,N_10468);
nor U10664 (N_10664,N_9986,N_10093);
or U10665 (N_10665,N_9836,N_10379);
or U10666 (N_10666,N_10347,N_10246);
nor U10667 (N_10667,N_10300,N_9816);
xnor U10668 (N_10668,N_10054,N_10311);
nand U10669 (N_10669,N_10080,N_9958);
or U10670 (N_10670,N_10039,N_9867);
nor U10671 (N_10671,N_9932,N_9777);
nand U10672 (N_10672,N_9821,N_10170);
nand U10673 (N_10673,N_10350,N_9863);
and U10674 (N_10674,N_10075,N_10335);
and U10675 (N_10675,N_10441,N_10485);
or U10676 (N_10676,N_10097,N_10408);
or U10677 (N_10677,N_10098,N_10355);
or U10678 (N_10678,N_10000,N_9802);
and U10679 (N_10679,N_10012,N_10312);
or U10680 (N_10680,N_9851,N_9970);
xnor U10681 (N_10681,N_10189,N_9774);
nor U10682 (N_10682,N_10476,N_9866);
nand U10683 (N_10683,N_9929,N_10121);
and U10684 (N_10684,N_10342,N_10331);
nor U10685 (N_10685,N_9973,N_9761);
or U10686 (N_10686,N_9803,N_10172);
nand U10687 (N_10687,N_9850,N_10229);
xnor U10688 (N_10688,N_10014,N_10413);
nand U10689 (N_10689,N_9977,N_9879);
and U10690 (N_10690,N_10084,N_10227);
or U10691 (N_10691,N_10256,N_9980);
nor U10692 (N_10692,N_9857,N_10482);
or U10693 (N_10693,N_9839,N_9825);
nand U10694 (N_10694,N_10291,N_10399);
or U10695 (N_10695,N_10330,N_10258);
nor U10696 (N_10696,N_10040,N_10050);
nand U10697 (N_10697,N_10087,N_10403);
or U10698 (N_10698,N_10017,N_10167);
and U10699 (N_10699,N_9892,N_10240);
or U10700 (N_10700,N_10296,N_9859);
nand U10701 (N_10701,N_9897,N_9995);
xnor U10702 (N_10702,N_9878,N_9873);
or U10703 (N_10703,N_9967,N_10139);
or U10704 (N_10704,N_9817,N_9765);
nor U10705 (N_10705,N_10090,N_10259);
nand U10706 (N_10706,N_9828,N_10152);
and U10707 (N_10707,N_9966,N_9942);
nor U10708 (N_10708,N_10328,N_10233);
or U10709 (N_10709,N_9772,N_10212);
and U10710 (N_10710,N_10489,N_10162);
nor U10711 (N_10711,N_10320,N_10314);
and U10712 (N_10712,N_9876,N_10466);
xor U10713 (N_10713,N_10486,N_10389);
and U10714 (N_10714,N_9862,N_10307);
nor U10715 (N_10715,N_10159,N_10264);
or U10716 (N_10716,N_10145,N_10270);
or U10717 (N_10717,N_10361,N_9804);
and U10718 (N_10718,N_9961,N_10452);
nand U10719 (N_10719,N_9883,N_9751);
nand U10720 (N_10720,N_10128,N_10116);
nor U10721 (N_10721,N_9946,N_10434);
nand U10722 (N_10722,N_10344,N_10275);
or U10723 (N_10723,N_10304,N_10282);
nand U10724 (N_10724,N_9785,N_9914);
and U10725 (N_10725,N_10208,N_9877);
xor U10726 (N_10726,N_10169,N_9789);
nor U10727 (N_10727,N_9969,N_10325);
or U10728 (N_10728,N_10310,N_10427);
nor U10729 (N_10729,N_9823,N_10338);
nor U10730 (N_10730,N_9752,N_10238);
and U10731 (N_10731,N_9959,N_10165);
and U10732 (N_10732,N_10429,N_9805);
and U10733 (N_10733,N_10457,N_10483);
or U10734 (N_10734,N_10272,N_9757);
nand U10735 (N_10735,N_9763,N_10028);
or U10736 (N_10736,N_10136,N_10412);
and U10737 (N_10737,N_10029,N_9787);
nand U10738 (N_10738,N_10378,N_9954);
nand U10739 (N_10739,N_10465,N_10123);
nand U10740 (N_10740,N_10228,N_10317);
nor U10741 (N_10741,N_10354,N_10431);
or U10742 (N_10742,N_10407,N_10237);
or U10743 (N_10743,N_10396,N_10449);
nand U10744 (N_10744,N_10173,N_9793);
or U10745 (N_10745,N_10166,N_10023);
xnor U10746 (N_10746,N_10114,N_9907);
or U10747 (N_10747,N_9888,N_9896);
and U10748 (N_10748,N_9779,N_10329);
and U10749 (N_10749,N_10447,N_9833);
nor U10750 (N_10750,N_10369,N_10153);
and U10751 (N_10751,N_10192,N_9801);
nand U10752 (N_10752,N_9764,N_10461);
nand U10753 (N_10753,N_9931,N_9903);
nor U10754 (N_10754,N_10315,N_10158);
and U10755 (N_10755,N_9987,N_10394);
or U10756 (N_10756,N_10257,N_10422);
nor U10757 (N_10757,N_10351,N_9835);
nor U10758 (N_10758,N_9998,N_10150);
nand U10759 (N_10759,N_10499,N_9947);
nor U10760 (N_10760,N_9780,N_10498);
xnor U10761 (N_10761,N_9963,N_10160);
or U10762 (N_10762,N_10286,N_10479);
and U10763 (N_10763,N_9971,N_10398);
and U10764 (N_10764,N_10332,N_9985);
nor U10765 (N_10765,N_10284,N_10079);
nor U10766 (N_10766,N_10359,N_9890);
or U10767 (N_10767,N_9791,N_9767);
nor U10768 (N_10768,N_10016,N_10439);
xor U10769 (N_10769,N_10119,N_9911);
nand U10770 (N_10770,N_10251,N_10366);
nor U10771 (N_10771,N_9844,N_10234);
nand U10772 (N_10772,N_10069,N_10448);
and U10773 (N_10773,N_10100,N_9915);
and U10774 (N_10774,N_9812,N_10316);
and U10775 (N_10775,N_9922,N_10289);
or U10776 (N_10776,N_9834,N_10339);
and U10777 (N_10777,N_10415,N_10416);
nor U10778 (N_10778,N_10387,N_9937);
or U10779 (N_10779,N_10409,N_10018);
xor U10780 (N_10780,N_10255,N_10364);
nor U10781 (N_10781,N_10358,N_10019);
nand U10782 (N_10782,N_10400,N_10405);
and U10783 (N_10783,N_10003,N_10281);
or U10784 (N_10784,N_10115,N_9917);
nand U10785 (N_10785,N_10033,N_10377);
xnor U10786 (N_10786,N_9875,N_10035);
nand U10787 (N_10787,N_10222,N_10156);
nor U10788 (N_10788,N_10207,N_9790);
nand U10789 (N_10789,N_10174,N_9818);
nor U10790 (N_10790,N_10271,N_10224);
or U10791 (N_10791,N_10279,N_9984);
and U10792 (N_10792,N_10225,N_10218);
xor U10793 (N_10793,N_10440,N_10046);
nor U10794 (N_10794,N_9784,N_10135);
and U10795 (N_10795,N_10105,N_10199);
nand U10796 (N_10796,N_10168,N_10239);
xnor U10797 (N_10797,N_10091,N_10083);
nand U10798 (N_10798,N_9861,N_10458);
xnor U10799 (N_10799,N_10143,N_10089);
nor U10800 (N_10800,N_10453,N_10074);
and U10801 (N_10801,N_9788,N_10308);
xor U10802 (N_10802,N_9991,N_10375);
or U10803 (N_10803,N_10055,N_10438);
and U10804 (N_10804,N_10133,N_10118);
and U10805 (N_10805,N_9869,N_10353);
nor U10806 (N_10806,N_10481,N_10024);
nand U10807 (N_10807,N_9808,N_10348);
nand U10808 (N_10808,N_10007,N_9989);
and U10809 (N_10809,N_10306,N_9936);
or U10810 (N_10810,N_10034,N_9864);
nor U10811 (N_10811,N_10231,N_10384);
nand U10812 (N_10812,N_9756,N_9905);
nor U10813 (N_10813,N_10477,N_10470);
or U10814 (N_10814,N_10473,N_10303);
and U10815 (N_10815,N_9760,N_9960);
nor U10816 (N_10816,N_9865,N_10419);
nor U10817 (N_10817,N_10371,N_10103);
nand U10818 (N_10818,N_9778,N_9976);
nand U10819 (N_10819,N_9849,N_10063);
nand U10820 (N_10820,N_10484,N_10294);
nand U10821 (N_10821,N_9924,N_10171);
xor U10822 (N_10822,N_9943,N_10045);
nor U10823 (N_10823,N_10032,N_10111);
nand U10824 (N_10824,N_10180,N_10395);
and U10825 (N_10825,N_9979,N_9992);
and U10826 (N_10826,N_10262,N_10092);
nand U10827 (N_10827,N_10179,N_10297);
or U10828 (N_10828,N_9935,N_10213);
and U10829 (N_10829,N_9827,N_10151);
xor U10830 (N_10830,N_10081,N_9948);
nor U10831 (N_10831,N_10185,N_10362);
nand U10832 (N_10832,N_9811,N_10030);
nand U10833 (N_10833,N_9881,N_10214);
nand U10834 (N_10834,N_9999,N_10436);
nor U10835 (N_10835,N_10265,N_10200);
xnor U10836 (N_10836,N_10073,N_9800);
nand U10837 (N_10837,N_10043,N_10008);
nor U10838 (N_10838,N_10076,N_10352);
nand U10839 (N_10839,N_10455,N_10243);
nand U10840 (N_10840,N_9927,N_10367);
xnor U10841 (N_10841,N_10406,N_10445);
nand U10842 (N_10842,N_10176,N_9830);
or U10843 (N_10843,N_9871,N_10122);
or U10844 (N_10844,N_10204,N_10230);
nand U10845 (N_10845,N_10283,N_10487);
and U10846 (N_10846,N_10326,N_10015);
nand U10847 (N_10847,N_9886,N_10261);
and U10848 (N_10848,N_10346,N_9758);
or U10849 (N_10849,N_9983,N_10309);
and U10850 (N_10850,N_9826,N_9840);
or U10851 (N_10851,N_10299,N_9923);
or U10852 (N_10852,N_10127,N_10432);
or U10853 (N_10853,N_10327,N_9809);
nand U10854 (N_10854,N_10252,N_10059);
nor U10855 (N_10855,N_10037,N_10480);
nand U10856 (N_10856,N_10051,N_10249);
nand U10857 (N_10857,N_10010,N_10217);
nand U10858 (N_10858,N_9884,N_9962);
or U10859 (N_10859,N_10492,N_10267);
xor U10860 (N_10860,N_9910,N_10341);
or U10861 (N_10861,N_10404,N_10197);
xor U10862 (N_10862,N_10357,N_9950);
nor U10863 (N_10863,N_10068,N_10011);
or U10864 (N_10864,N_9829,N_10061);
or U10865 (N_10865,N_10250,N_10298);
nor U10866 (N_10866,N_10490,N_10131);
nor U10867 (N_10867,N_10187,N_9993);
nor U10868 (N_10868,N_10096,N_9898);
xor U10869 (N_10869,N_10223,N_9891);
nor U10870 (N_10870,N_10446,N_10155);
nand U10871 (N_10871,N_10038,N_9852);
nand U10872 (N_10872,N_10049,N_9814);
nand U10873 (N_10873,N_10193,N_10163);
nor U10874 (N_10874,N_10070,N_9880);
or U10875 (N_10875,N_9844,N_10253);
nor U10876 (N_10876,N_9884,N_10118);
nand U10877 (N_10877,N_9914,N_9955);
or U10878 (N_10878,N_10139,N_10150);
nor U10879 (N_10879,N_10425,N_10110);
or U10880 (N_10880,N_10250,N_9884);
or U10881 (N_10881,N_10281,N_10039);
nand U10882 (N_10882,N_10309,N_10055);
and U10883 (N_10883,N_10243,N_9921);
nand U10884 (N_10884,N_9899,N_10129);
or U10885 (N_10885,N_10123,N_10236);
or U10886 (N_10886,N_10156,N_9963);
or U10887 (N_10887,N_10151,N_9921);
nand U10888 (N_10888,N_9879,N_10219);
nand U10889 (N_10889,N_10230,N_10086);
nand U10890 (N_10890,N_9778,N_9840);
nand U10891 (N_10891,N_10030,N_10191);
or U10892 (N_10892,N_9909,N_9964);
nand U10893 (N_10893,N_10162,N_10247);
nand U10894 (N_10894,N_10348,N_10163);
nor U10895 (N_10895,N_9755,N_10374);
and U10896 (N_10896,N_9876,N_10419);
or U10897 (N_10897,N_10426,N_9913);
xor U10898 (N_10898,N_10415,N_10357);
and U10899 (N_10899,N_9930,N_10103);
nand U10900 (N_10900,N_10139,N_10445);
and U10901 (N_10901,N_10391,N_10035);
or U10902 (N_10902,N_10091,N_10338);
or U10903 (N_10903,N_10255,N_10400);
xnor U10904 (N_10904,N_10460,N_9881);
nor U10905 (N_10905,N_10195,N_9750);
and U10906 (N_10906,N_9806,N_10052);
and U10907 (N_10907,N_10249,N_10208);
nand U10908 (N_10908,N_10240,N_10244);
nor U10909 (N_10909,N_10297,N_10316);
and U10910 (N_10910,N_10229,N_9993);
nand U10911 (N_10911,N_10310,N_10239);
or U10912 (N_10912,N_9993,N_10238);
xor U10913 (N_10913,N_9932,N_9900);
or U10914 (N_10914,N_10440,N_10350);
or U10915 (N_10915,N_10055,N_9868);
and U10916 (N_10916,N_10428,N_10457);
nor U10917 (N_10917,N_9892,N_10340);
nand U10918 (N_10918,N_9841,N_10401);
and U10919 (N_10919,N_10180,N_10312);
or U10920 (N_10920,N_10197,N_10097);
and U10921 (N_10921,N_9877,N_9967);
or U10922 (N_10922,N_10258,N_10332);
or U10923 (N_10923,N_10342,N_10264);
and U10924 (N_10924,N_10318,N_10326);
nor U10925 (N_10925,N_9952,N_10320);
nor U10926 (N_10926,N_10477,N_9862);
nor U10927 (N_10927,N_9880,N_9865);
and U10928 (N_10928,N_10287,N_10221);
nand U10929 (N_10929,N_10479,N_9884);
or U10930 (N_10930,N_10454,N_10229);
nand U10931 (N_10931,N_10164,N_10042);
or U10932 (N_10932,N_10453,N_10033);
nand U10933 (N_10933,N_10417,N_10154);
nor U10934 (N_10934,N_10162,N_10226);
nor U10935 (N_10935,N_10173,N_9808);
nor U10936 (N_10936,N_10201,N_10077);
nand U10937 (N_10937,N_10097,N_10019);
nand U10938 (N_10938,N_10318,N_10474);
or U10939 (N_10939,N_10254,N_9957);
and U10940 (N_10940,N_9964,N_9943);
nor U10941 (N_10941,N_9844,N_10147);
and U10942 (N_10942,N_9781,N_9807);
and U10943 (N_10943,N_10407,N_10203);
and U10944 (N_10944,N_10207,N_10367);
nand U10945 (N_10945,N_10220,N_10443);
nand U10946 (N_10946,N_10025,N_10238);
nor U10947 (N_10947,N_9783,N_9823);
and U10948 (N_10948,N_10134,N_10369);
or U10949 (N_10949,N_10347,N_9839);
nor U10950 (N_10950,N_10100,N_9954);
xor U10951 (N_10951,N_9816,N_10489);
xor U10952 (N_10952,N_9989,N_10329);
or U10953 (N_10953,N_9876,N_10407);
and U10954 (N_10954,N_10221,N_9918);
or U10955 (N_10955,N_9946,N_10177);
or U10956 (N_10956,N_10299,N_9951);
nand U10957 (N_10957,N_9761,N_10188);
or U10958 (N_10958,N_10351,N_9904);
nand U10959 (N_10959,N_10337,N_9923);
or U10960 (N_10960,N_10309,N_10133);
or U10961 (N_10961,N_10068,N_9941);
xnor U10962 (N_10962,N_9959,N_10366);
nand U10963 (N_10963,N_10351,N_9851);
nand U10964 (N_10964,N_9890,N_9964);
nand U10965 (N_10965,N_10496,N_10203);
nor U10966 (N_10966,N_10125,N_9792);
or U10967 (N_10967,N_10057,N_10321);
nand U10968 (N_10968,N_9797,N_9854);
nor U10969 (N_10969,N_9919,N_10223);
or U10970 (N_10970,N_9976,N_10054);
or U10971 (N_10971,N_9815,N_10165);
nor U10972 (N_10972,N_10330,N_10271);
or U10973 (N_10973,N_10017,N_10027);
or U10974 (N_10974,N_9816,N_10462);
nor U10975 (N_10975,N_10384,N_10280);
nand U10976 (N_10976,N_9788,N_9806);
nor U10977 (N_10977,N_9968,N_10472);
xor U10978 (N_10978,N_10296,N_10079);
or U10979 (N_10979,N_10295,N_10395);
nand U10980 (N_10980,N_9914,N_10088);
and U10981 (N_10981,N_9987,N_10299);
nor U10982 (N_10982,N_9925,N_10125);
nor U10983 (N_10983,N_9862,N_10185);
nor U10984 (N_10984,N_9776,N_9851);
nand U10985 (N_10985,N_10021,N_9990);
nor U10986 (N_10986,N_9786,N_9999);
nor U10987 (N_10987,N_9907,N_9882);
nand U10988 (N_10988,N_9929,N_10476);
and U10989 (N_10989,N_9930,N_10354);
and U10990 (N_10990,N_9791,N_10328);
or U10991 (N_10991,N_9931,N_10465);
or U10992 (N_10992,N_10109,N_10393);
nand U10993 (N_10993,N_10014,N_10417);
or U10994 (N_10994,N_10144,N_10034);
or U10995 (N_10995,N_9834,N_10088);
and U10996 (N_10996,N_10462,N_10485);
and U10997 (N_10997,N_9764,N_10251);
nand U10998 (N_10998,N_9782,N_9879);
nand U10999 (N_10999,N_9985,N_10485);
nand U11000 (N_11000,N_9869,N_10387);
xnor U11001 (N_11001,N_9773,N_10394);
nor U11002 (N_11002,N_10010,N_10356);
and U11003 (N_11003,N_10433,N_9962);
or U11004 (N_11004,N_10322,N_10267);
and U11005 (N_11005,N_10144,N_10383);
nor U11006 (N_11006,N_9969,N_9834);
and U11007 (N_11007,N_10291,N_10301);
nor U11008 (N_11008,N_10135,N_10298);
nand U11009 (N_11009,N_10056,N_10208);
and U11010 (N_11010,N_10255,N_10045);
and U11011 (N_11011,N_10022,N_9839);
nand U11012 (N_11012,N_9808,N_10282);
and U11013 (N_11013,N_10009,N_10379);
and U11014 (N_11014,N_10055,N_10468);
and U11015 (N_11015,N_10347,N_10483);
or U11016 (N_11016,N_10368,N_9884);
and U11017 (N_11017,N_9976,N_9770);
nand U11018 (N_11018,N_9937,N_10330);
or U11019 (N_11019,N_10053,N_9955);
or U11020 (N_11020,N_10152,N_10311);
or U11021 (N_11021,N_10204,N_9871);
or U11022 (N_11022,N_9923,N_10331);
and U11023 (N_11023,N_10226,N_10049);
and U11024 (N_11024,N_9924,N_10403);
or U11025 (N_11025,N_10126,N_9945);
or U11026 (N_11026,N_10293,N_10320);
nor U11027 (N_11027,N_10378,N_9986);
or U11028 (N_11028,N_10337,N_10182);
and U11029 (N_11029,N_9939,N_10294);
nand U11030 (N_11030,N_10287,N_10001);
or U11031 (N_11031,N_9825,N_10032);
nand U11032 (N_11032,N_9767,N_10493);
or U11033 (N_11033,N_10477,N_10155);
nand U11034 (N_11034,N_10078,N_10281);
and U11035 (N_11035,N_10457,N_10272);
nor U11036 (N_11036,N_10213,N_10336);
and U11037 (N_11037,N_10396,N_10359);
and U11038 (N_11038,N_9888,N_10353);
nor U11039 (N_11039,N_10123,N_9863);
or U11040 (N_11040,N_10258,N_9867);
nand U11041 (N_11041,N_10430,N_10493);
or U11042 (N_11042,N_9896,N_9761);
nor U11043 (N_11043,N_10391,N_10126);
nor U11044 (N_11044,N_10270,N_10348);
and U11045 (N_11045,N_10281,N_10067);
nand U11046 (N_11046,N_10488,N_10351);
nor U11047 (N_11047,N_10451,N_10017);
nand U11048 (N_11048,N_10029,N_10368);
and U11049 (N_11049,N_10043,N_10263);
or U11050 (N_11050,N_10037,N_9821);
nand U11051 (N_11051,N_10239,N_10498);
nand U11052 (N_11052,N_9781,N_10489);
nand U11053 (N_11053,N_10177,N_10222);
nand U11054 (N_11054,N_10303,N_10418);
nand U11055 (N_11055,N_10200,N_10354);
nor U11056 (N_11056,N_10103,N_10473);
nand U11057 (N_11057,N_9968,N_10158);
nor U11058 (N_11058,N_9979,N_10310);
and U11059 (N_11059,N_10386,N_10405);
nor U11060 (N_11060,N_9975,N_10491);
xor U11061 (N_11061,N_10104,N_10395);
nor U11062 (N_11062,N_10216,N_10011);
nor U11063 (N_11063,N_9778,N_10379);
and U11064 (N_11064,N_10295,N_9834);
nand U11065 (N_11065,N_9786,N_9857);
or U11066 (N_11066,N_9750,N_10337);
nor U11067 (N_11067,N_9779,N_10479);
xor U11068 (N_11068,N_10057,N_10399);
nor U11069 (N_11069,N_9756,N_10315);
nand U11070 (N_11070,N_10017,N_9942);
and U11071 (N_11071,N_9877,N_9868);
nand U11072 (N_11072,N_9978,N_9887);
or U11073 (N_11073,N_9772,N_9945);
or U11074 (N_11074,N_9991,N_10155);
nor U11075 (N_11075,N_9775,N_9753);
nor U11076 (N_11076,N_10416,N_10265);
nor U11077 (N_11077,N_10029,N_10482);
xnor U11078 (N_11078,N_9784,N_10087);
nand U11079 (N_11079,N_10406,N_10196);
nand U11080 (N_11080,N_10232,N_9885);
nor U11081 (N_11081,N_10186,N_10147);
and U11082 (N_11082,N_9838,N_10411);
nor U11083 (N_11083,N_10346,N_9849);
and U11084 (N_11084,N_10302,N_9994);
nand U11085 (N_11085,N_10426,N_10350);
nand U11086 (N_11086,N_10390,N_10209);
and U11087 (N_11087,N_10036,N_10381);
or U11088 (N_11088,N_10311,N_9795);
or U11089 (N_11089,N_10226,N_9848);
or U11090 (N_11090,N_10298,N_10202);
nand U11091 (N_11091,N_9843,N_9945);
and U11092 (N_11092,N_10365,N_9849);
xnor U11093 (N_11093,N_10105,N_9784);
xnor U11094 (N_11094,N_9805,N_9850);
or U11095 (N_11095,N_10038,N_10160);
and U11096 (N_11096,N_10235,N_9893);
or U11097 (N_11097,N_9829,N_10348);
or U11098 (N_11098,N_10019,N_9999);
or U11099 (N_11099,N_10000,N_9899);
xor U11100 (N_11100,N_10116,N_10451);
or U11101 (N_11101,N_10005,N_10217);
xnor U11102 (N_11102,N_10392,N_10444);
or U11103 (N_11103,N_9817,N_9751);
xnor U11104 (N_11104,N_10167,N_10040);
nor U11105 (N_11105,N_10358,N_9844);
nor U11106 (N_11106,N_9807,N_10186);
nor U11107 (N_11107,N_10421,N_10130);
nand U11108 (N_11108,N_9972,N_10338);
nand U11109 (N_11109,N_10019,N_9761);
and U11110 (N_11110,N_10038,N_10478);
nand U11111 (N_11111,N_9891,N_10094);
and U11112 (N_11112,N_10313,N_9846);
nand U11113 (N_11113,N_9917,N_10188);
nor U11114 (N_11114,N_10112,N_9937);
xor U11115 (N_11115,N_10158,N_9763);
nand U11116 (N_11116,N_9869,N_9943);
nor U11117 (N_11117,N_9895,N_10008);
and U11118 (N_11118,N_10203,N_10307);
xnor U11119 (N_11119,N_10436,N_9887);
or U11120 (N_11120,N_9870,N_10143);
nand U11121 (N_11121,N_10023,N_10003);
and U11122 (N_11122,N_9888,N_9893);
or U11123 (N_11123,N_10162,N_10378);
or U11124 (N_11124,N_10348,N_9798);
nand U11125 (N_11125,N_10247,N_10442);
nand U11126 (N_11126,N_10243,N_9966);
nor U11127 (N_11127,N_9900,N_10172);
nand U11128 (N_11128,N_10339,N_9829);
xor U11129 (N_11129,N_10244,N_9768);
xor U11130 (N_11130,N_10444,N_10069);
or U11131 (N_11131,N_9883,N_9810);
and U11132 (N_11132,N_10118,N_10087);
and U11133 (N_11133,N_9847,N_10408);
nor U11134 (N_11134,N_10261,N_9837);
nand U11135 (N_11135,N_10295,N_10272);
nor U11136 (N_11136,N_10319,N_9831);
nor U11137 (N_11137,N_10254,N_10347);
or U11138 (N_11138,N_10177,N_9855);
or U11139 (N_11139,N_9897,N_9876);
nand U11140 (N_11140,N_10265,N_10194);
nor U11141 (N_11141,N_9819,N_10260);
nor U11142 (N_11142,N_10339,N_10380);
xor U11143 (N_11143,N_10491,N_9841);
nor U11144 (N_11144,N_10124,N_9757);
xnor U11145 (N_11145,N_9821,N_9844);
nor U11146 (N_11146,N_9997,N_9884);
and U11147 (N_11147,N_10417,N_10439);
or U11148 (N_11148,N_10133,N_9841);
nand U11149 (N_11149,N_9829,N_10422);
xor U11150 (N_11150,N_10455,N_9906);
nor U11151 (N_11151,N_9771,N_9766);
nor U11152 (N_11152,N_10095,N_10285);
nand U11153 (N_11153,N_9899,N_10464);
nor U11154 (N_11154,N_10110,N_9960);
and U11155 (N_11155,N_10301,N_10342);
nand U11156 (N_11156,N_10415,N_10216);
and U11157 (N_11157,N_9936,N_10254);
nand U11158 (N_11158,N_10067,N_10331);
xnor U11159 (N_11159,N_9915,N_9822);
nor U11160 (N_11160,N_9918,N_9967);
nand U11161 (N_11161,N_10430,N_10110);
or U11162 (N_11162,N_10336,N_9750);
nor U11163 (N_11163,N_9774,N_10457);
nor U11164 (N_11164,N_10251,N_10309);
nor U11165 (N_11165,N_10124,N_10320);
nand U11166 (N_11166,N_9865,N_9810);
or U11167 (N_11167,N_10338,N_10402);
nand U11168 (N_11168,N_9978,N_10129);
nand U11169 (N_11169,N_10192,N_10262);
nor U11170 (N_11170,N_10003,N_10282);
and U11171 (N_11171,N_10123,N_10103);
xor U11172 (N_11172,N_10040,N_10382);
and U11173 (N_11173,N_10319,N_10448);
nand U11174 (N_11174,N_10209,N_9913);
nor U11175 (N_11175,N_10443,N_10214);
nand U11176 (N_11176,N_9875,N_10043);
nand U11177 (N_11177,N_10370,N_9948);
nand U11178 (N_11178,N_10333,N_10415);
and U11179 (N_11179,N_9949,N_10078);
or U11180 (N_11180,N_9771,N_9832);
nand U11181 (N_11181,N_10356,N_10497);
or U11182 (N_11182,N_9969,N_10494);
nor U11183 (N_11183,N_10160,N_10466);
xor U11184 (N_11184,N_10192,N_10275);
nand U11185 (N_11185,N_10443,N_10495);
xor U11186 (N_11186,N_10313,N_9927);
nor U11187 (N_11187,N_10194,N_9962);
nand U11188 (N_11188,N_10409,N_10195);
nand U11189 (N_11189,N_10305,N_10180);
or U11190 (N_11190,N_10079,N_10455);
nor U11191 (N_11191,N_9795,N_10091);
and U11192 (N_11192,N_10130,N_9903);
or U11193 (N_11193,N_10068,N_9775);
and U11194 (N_11194,N_10377,N_10430);
nand U11195 (N_11195,N_10173,N_9906);
nor U11196 (N_11196,N_10191,N_10129);
nand U11197 (N_11197,N_10433,N_9775);
nor U11198 (N_11198,N_9800,N_10289);
xor U11199 (N_11199,N_10094,N_9804);
and U11200 (N_11200,N_9973,N_10192);
nor U11201 (N_11201,N_10251,N_10142);
nand U11202 (N_11202,N_10157,N_10405);
nand U11203 (N_11203,N_10125,N_10493);
nor U11204 (N_11204,N_10034,N_10418);
nand U11205 (N_11205,N_10360,N_10160);
or U11206 (N_11206,N_10339,N_10376);
xor U11207 (N_11207,N_9826,N_10010);
and U11208 (N_11208,N_10474,N_10014);
xnor U11209 (N_11209,N_10017,N_9861);
nor U11210 (N_11210,N_9750,N_10470);
and U11211 (N_11211,N_10080,N_9906);
nor U11212 (N_11212,N_10369,N_10493);
or U11213 (N_11213,N_10497,N_10336);
nor U11214 (N_11214,N_10029,N_10008);
nor U11215 (N_11215,N_9916,N_9884);
and U11216 (N_11216,N_10250,N_9845);
xnor U11217 (N_11217,N_10374,N_9941);
nand U11218 (N_11218,N_9852,N_9992);
xnor U11219 (N_11219,N_10035,N_10359);
and U11220 (N_11220,N_9872,N_10414);
nor U11221 (N_11221,N_10430,N_10155);
nand U11222 (N_11222,N_9897,N_10404);
and U11223 (N_11223,N_10412,N_10151);
and U11224 (N_11224,N_10016,N_10069);
and U11225 (N_11225,N_10403,N_10073);
nand U11226 (N_11226,N_9820,N_9907);
nor U11227 (N_11227,N_10157,N_9866);
nand U11228 (N_11228,N_9961,N_10367);
nor U11229 (N_11229,N_10413,N_9781);
or U11230 (N_11230,N_9970,N_9965);
or U11231 (N_11231,N_10159,N_10445);
xnor U11232 (N_11232,N_10018,N_9836);
and U11233 (N_11233,N_10448,N_10068);
nor U11234 (N_11234,N_10471,N_10220);
or U11235 (N_11235,N_9862,N_10349);
nor U11236 (N_11236,N_10114,N_9816);
or U11237 (N_11237,N_10390,N_10450);
or U11238 (N_11238,N_9985,N_10148);
nand U11239 (N_11239,N_9828,N_10038);
and U11240 (N_11240,N_10010,N_9751);
or U11241 (N_11241,N_10097,N_10367);
and U11242 (N_11242,N_10038,N_9993);
and U11243 (N_11243,N_10110,N_9799);
or U11244 (N_11244,N_10324,N_10020);
nand U11245 (N_11245,N_9793,N_9827);
or U11246 (N_11246,N_9852,N_9920);
and U11247 (N_11247,N_10322,N_9929);
nand U11248 (N_11248,N_10191,N_10198);
or U11249 (N_11249,N_10282,N_10352);
and U11250 (N_11250,N_10921,N_10637);
and U11251 (N_11251,N_11139,N_10882);
and U11252 (N_11252,N_10655,N_10932);
or U11253 (N_11253,N_11090,N_11196);
or U11254 (N_11254,N_11080,N_11013);
nand U11255 (N_11255,N_10728,N_10792);
xor U11256 (N_11256,N_10591,N_10675);
xnor U11257 (N_11257,N_11143,N_10966);
and U11258 (N_11258,N_11040,N_11228);
or U11259 (N_11259,N_10880,N_11206);
and U11260 (N_11260,N_11066,N_10557);
nand U11261 (N_11261,N_10917,N_10944);
or U11262 (N_11262,N_10732,N_10963);
nor U11263 (N_11263,N_11144,N_11224);
nand U11264 (N_11264,N_10708,N_10746);
nor U11265 (N_11265,N_10945,N_10936);
nand U11266 (N_11266,N_10711,N_11106);
nor U11267 (N_11267,N_10807,N_10626);
or U11268 (N_11268,N_10687,N_10910);
xnor U11269 (N_11269,N_10791,N_10786);
nand U11270 (N_11270,N_11054,N_11010);
nor U11271 (N_11271,N_10766,N_10813);
nor U11272 (N_11272,N_11068,N_10794);
xor U11273 (N_11273,N_10605,N_10751);
and U11274 (N_11274,N_11022,N_10744);
and U11275 (N_11275,N_10552,N_11097);
or U11276 (N_11276,N_11023,N_10938);
nor U11277 (N_11277,N_10601,N_10901);
nor U11278 (N_11278,N_10610,N_10506);
nand U11279 (N_11279,N_11152,N_10509);
or U11280 (N_11280,N_10815,N_11035);
nand U11281 (N_11281,N_10510,N_10712);
nand U11282 (N_11282,N_10679,N_10600);
nor U11283 (N_11283,N_10707,N_10689);
nor U11284 (N_11284,N_10577,N_10690);
or U11285 (N_11285,N_11173,N_11094);
and U11286 (N_11286,N_11232,N_10926);
nor U11287 (N_11287,N_10832,N_11088);
or U11288 (N_11288,N_10902,N_10952);
nand U11289 (N_11289,N_11205,N_11081);
nand U11290 (N_11290,N_10940,N_10955);
nor U11291 (N_11291,N_10915,N_11132);
or U11292 (N_11292,N_10544,N_10602);
nor U11293 (N_11293,N_10623,N_11174);
or U11294 (N_11294,N_10671,N_10923);
nor U11295 (N_11295,N_10775,N_11154);
and U11296 (N_11296,N_10849,N_11103);
xnor U11297 (N_11297,N_10654,N_10759);
nand U11298 (N_11298,N_10918,N_10651);
or U11299 (N_11299,N_11243,N_10512);
nand U11300 (N_11300,N_10677,N_10907);
xnor U11301 (N_11301,N_11169,N_10593);
nor U11302 (N_11302,N_11133,N_10554);
nand U11303 (N_11303,N_10884,N_10505);
xnor U11304 (N_11304,N_11027,N_10795);
nand U11305 (N_11305,N_10906,N_11170);
or U11306 (N_11306,N_11158,N_10565);
and U11307 (N_11307,N_11202,N_10636);
and U11308 (N_11308,N_10978,N_10987);
and U11309 (N_11309,N_11070,N_10716);
xnor U11310 (N_11310,N_11122,N_11182);
and U11311 (N_11311,N_11234,N_11091);
nand U11312 (N_11312,N_10972,N_10925);
or U11313 (N_11313,N_11084,N_10586);
nand U11314 (N_11314,N_10549,N_10620);
or U11315 (N_11315,N_10953,N_10771);
or U11316 (N_11316,N_10782,N_11093);
nor U11317 (N_11317,N_10580,N_11037);
nand U11318 (N_11318,N_10912,N_10797);
nand U11319 (N_11319,N_10673,N_10665);
xor U11320 (N_11320,N_11180,N_10648);
or U11321 (N_11321,N_11026,N_11100);
and U11322 (N_11322,N_10919,N_10578);
nand U11323 (N_11323,N_11204,N_10559);
and U11324 (N_11324,N_10830,N_11108);
nand U11325 (N_11325,N_10543,N_11151);
or U11326 (N_11326,N_10958,N_11101);
and U11327 (N_11327,N_11160,N_10676);
nand U11328 (N_11328,N_11141,N_10803);
nand U11329 (N_11329,N_11059,N_11007);
or U11330 (N_11330,N_11045,N_11057);
or U11331 (N_11331,N_10800,N_11236);
and U11332 (N_11332,N_10762,N_11172);
nor U11333 (N_11333,N_10804,N_10866);
and U11334 (N_11334,N_11208,N_10717);
nor U11335 (N_11335,N_10860,N_10727);
or U11336 (N_11336,N_11120,N_10553);
or U11337 (N_11337,N_10533,N_10905);
or U11338 (N_11338,N_10599,N_10777);
and U11339 (N_11339,N_11183,N_10563);
nand U11340 (N_11340,N_11055,N_11166);
and U11341 (N_11341,N_10974,N_10962);
and U11342 (N_11342,N_10778,N_11248);
and U11343 (N_11343,N_10576,N_10574);
and U11344 (N_11344,N_10562,N_10625);
and U11345 (N_11345,N_11118,N_10761);
or U11346 (N_11346,N_10783,N_11213);
and U11347 (N_11347,N_11214,N_10501);
nand U11348 (N_11348,N_10756,N_10603);
and U11349 (N_11349,N_10887,N_11085);
xnor U11350 (N_11350,N_10556,N_11241);
and U11351 (N_11351,N_10725,N_10691);
or U11352 (N_11352,N_10993,N_10930);
or U11353 (N_11353,N_11074,N_11155);
and U11354 (N_11354,N_10518,N_10871);
nor U11355 (N_11355,N_11092,N_10808);
nand U11356 (N_11356,N_10839,N_11095);
and U11357 (N_11357,N_10942,N_11046);
and U11358 (N_11358,N_10848,N_11187);
nor U11359 (N_11359,N_10971,N_10816);
or U11360 (N_11360,N_10644,N_11192);
nand U11361 (N_11361,N_10522,N_11015);
nor U11362 (N_11362,N_11082,N_11159);
nor U11363 (N_11363,N_10841,N_11012);
or U11364 (N_11364,N_11038,N_11096);
and U11365 (N_11365,N_11107,N_10570);
nor U11366 (N_11366,N_10596,N_11000);
xnor U11367 (N_11367,N_11011,N_10519);
nand U11368 (N_11368,N_10566,N_10956);
nor U11369 (N_11369,N_11052,N_11203);
nand U11370 (N_11370,N_11005,N_10529);
or U11371 (N_11371,N_10667,N_11110);
xor U11372 (N_11372,N_10516,N_10703);
or U11373 (N_11373,N_10617,N_10560);
and U11374 (N_11374,N_10827,N_10640);
nand U11375 (N_11375,N_11147,N_10619);
xor U11376 (N_11376,N_10856,N_10730);
or U11377 (N_11377,N_11157,N_10545);
and U11378 (N_11378,N_10686,N_10838);
nand U11379 (N_11379,N_10948,N_10656);
or U11380 (N_11380,N_10634,N_10685);
nand U11381 (N_11381,N_10729,N_10503);
xnor U11382 (N_11382,N_10863,N_10535);
and U11383 (N_11383,N_10811,N_11226);
nand U11384 (N_11384,N_10997,N_10643);
nand U11385 (N_11385,N_10844,N_10742);
nand U11386 (N_11386,N_11211,N_11177);
nand U11387 (N_11387,N_10718,N_10755);
and U11388 (N_11388,N_10627,N_10810);
nand U11389 (N_11389,N_11197,N_10564);
nor U11390 (N_11390,N_10977,N_10579);
nor U11391 (N_11391,N_11140,N_11222);
nand U11392 (N_11392,N_11242,N_10957);
and U11393 (N_11393,N_11217,N_10969);
or U11394 (N_11394,N_10949,N_10779);
nand U11395 (N_11395,N_10852,N_10861);
xnor U11396 (N_11396,N_11077,N_10666);
or U11397 (N_11397,N_10678,N_10674);
nor U11398 (N_11398,N_11069,N_11239);
or U11399 (N_11399,N_10870,N_11064);
xnor U11400 (N_11400,N_10897,N_10511);
nand U11401 (N_11401,N_11089,N_11067);
nand U11402 (N_11402,N_11021,N_10749);
and U11403 (N_11403,N_10988,N_10622);
and U11404 (N_11404,N_11249,N_11071);
and U11405 (N_11405,N_10927,N_10959);
xor U11406 (N_11406,N_10735,N_10747);
nand U11407 (N_11407,N_11235,N_10547);
or U11408 (N_11408,N_10913,N_10753);
xnor U11409 (N_11409,N_11223,N_10594);
nand U11410 (N_11410,N_10572,N_10850);
nand U11411 (N_11411,N_10883,N_11171);
nor U11412 (N_11412,N_10701,N_10612);
and U11413 (N_11413,N_11207,N_10934);
nand U11414 (N_11414,N_10542,N_10822);
nand U11415 (N_11415,N_10981,N_11176);
nor U11416 (N_11416,N_11033,N_11009);
nor U11417 (N_11417,N_10967,N_10631);
or U11418 (N_11418,N_10774,N_10715);
nand U11419 (N_11419,N_11201,N_10688);
nand U11420 (N_11420,N_10878,N_10650);
or U11421 (N_11421,N_11185,N_11198);
or U11422 (N_11422,N_10515,N_10857);
or U11423 (N_11423,N_10968,N_11209);
nor U11424 (N_11424,N_10858,N_10891);
xor U11425 (N_11425,N_10788,N_11212);
nand U11426 (N_11426,N_10680,N_10639);
nor U11427 (N_11427,N_11104,N_10611);
nor U11428 (N_11428,N_10983,N_10911);
nor U11429 (N_11429,N_11028,N_11221);
or U11430 (N_11430,N_11238,N_11179);
and U11431 (N_11431,N_11246,N_11247);
nor U11432 (N_11432,N_11167,N_10820);
or U11433 (N_11433,N_10660,N_10581);
and U11434 (N_11434,N_10790,N_10835);
and U11435 (N_11435,N_11060,N_11244);
and U11436 (N_11436,N_10785,N_10796);
nor U11437 (N_11437,N_10693,N_10865);
and U11438 (N_11438,N_10597,N_10946);
or U11439 (N_11439,N_11076,N_11215);
nand U11440 (N_11440,N_10886,N_11014);
nand U11441 (N_11441,N_11137,N_10672);
or U11442 (N_11442,N_10824,N_10970);
and U11443 (N_11443,N_10741,N_11017);
nor U11444 (N_11444,N_10933,N_10931);
and U11445 (N_11445,N_10696,N_10895);
or U11446 (N_11446,N_10534,N_11138);
nand U11447 (N_11447,N_10659,N_10979);
nand U11448 (N_11448,N_10748,N_10538);
and U11449 (N_11449,N_10985,N_10641);
or U11450 (N_11450,N_10573,N_10984);
or U11451 (N_11451,N_11225,N_10645);
nand U11452 (N_11452,N_10699,N_10721);
nor U11453 (N_11453,N_11131,N_11124);
or U11454 (N_11454,N_11175,N_11061);
or U11455 (N_11455,N_10642,N_11079);
nand U11456 (N_11456,N_10604,N_11142);
nor U11457 (N_11457,N_10592,N_10828);
or U11458 (N_11458,N_11126,N_10881);
nand U11459 (N_11459,N_10561,N_10550);
xor U11460 (N_11460,N_10541,N_10507);
or U11461 (N_11461,N_11195,N_11109);
or U11462 (N_11462,N_11186,N_10776);
or U11463 (N_11463,N_10855,N_10525);
nand U11464 (N_11464,N_10750,N_10769);
or U11465 (N_11465,N_11168,N_10632);
nor U11466 (N_11466,N_10825,N_10836);
nand U11467 (N_11467,N_10664,N_11161);
nor U11468 (N_11468,N_11129,N_10722);
and U11469 (N_11469,N_11098,N_10862);
nand U11470 (N_11470,N_10874,N_10531);
and U11471 (N_11471,N_10812,N_11051);
nand U11472 (N_11472,N_10904,N_10767);
nand U11473 (N_11473,N_10684,N_10635);
or U11474 (N_11474,N_10532,N_10526);
or U11475 (N_11475,N_10873,N_11024);
and U11476 (N_11476,N_11008,N_11156);
or U11477 (N_11477,N_11164,N_11062);
nor U11478 (N_11478,N_10724,N_11034);
and U11479 (N_11479,N_10705,N_10896);
nand U11480 (N_11480,N_11127,N_10998);
or U11481 (N_11481,N_10859,N_11220);
or U11482 (N_11482,N_11117,N_10999);
nand U11483 (N_11483,N_10681,N_10787);
nor U11484 (N_11484,N_10698,N_11065);
xor U11485 (N_11485,N_10663,N_10657);
xnor U11486 (N_11486,N_10845,N_10840);
nor U11487 (N_11487,N_10924,N_11184);
nand U11488 (N_11488,N_11072,N_10521);
and U11489 (N_11489,N_10589,N_11042);
or U11490 (N_11490,N_11087,N_10613);
and U11491 (N_11491,N_11237,N_10991);
or U11492 (N_11492,N_11049,N_10714);
nand U11493 (N_11493,N_10670,N_10965);
nor U11494 (N_11494,N_10768,N_10540);
nor U11495 (N_11495,N_10615,N_10668);
or U11496 (N_11496,N_11149,N_11053);
or U11497 (N_11497,N_11146,N_10763);
and U11498 (N_11498,N_11114,N_10986);
or U11499 (N_11499,N_11189,N_11099);
nand U11500 (N_11500,N_10704,N_10834);
nor U11501 (N_11501,N_10809,N_11135);
or U11502 (N_11502,N_10647,N_11003);
or U11503 (N_11503,N_10894,N_10996);
nand U11504 (N_11504,N_11047,N_11004);
nor U11505 (N_11505,N_11163,N_10793);
and U11506 (N_11506,N_10502,N_10821);
nand U11507 (N_11507,N_11078,N_10853);
nor U11508 (N_11508,N_11229,N_10831);
nand U11509 (N_11509,N_10558,N_10843);
or U11510 (N_11510,N_10837,N_10598);
or U11511 (N_11511,N_10889,N_10713);
and U11512 (N_11512,N_10536,N_10964);
or U11513 (N_11513,N_10528,N_11200);
nand U11514 (N_11514,N_10903,N_11112);
or U11515 (N_11515,N_10630,N_11006);
and U11516 (N_11516,N_11086,N_11019);
xor U11517 (N_11517,N_10764,N_10618);
nor U11518 (N_11518,N_10569,N_10773);
nand U11519 (N_11519,N_11073,N_10826);
or U11520 (N_11520,N_11058,N_10738);
nand U11521 (N_11521,N_11111,N_10719);
nor U11522 (N_11522,N_11048,N_10819);
xor U11523 (N_11523,N_11199,N_10734);
nor U11524 (N_11524,N_10973,N_10624);
and U11525 (N_11525,N_10517,N_10607);
and U11526 (N_11526,N_10818,N_11136);
and U11527 (N_11527,N_11056,N_10802);
nor U11528 (N_11528,N_10723,N_10745);
nand U11529 (N_11529,N_11219,N_10928);
and U11530 (N_11530,N_11130,N_10954);
nand U11531 (N_11531,N_10683,N_11181);
nand U11532 (N_11532,N_10799,N_10575);
and U11533 (N_11533,N_10888,N_10854);
nor U11534 (N_11534,N_10548,N_11190);
and U11535 (N_11535,N_10752,N_11227);
nor U11536 (N_11536,N_10982,N_10899);
or U11537 (N_11537,N_11240,N_10770);
or U11538 (N_11538,N_10765,N_10833);
nor U11539 (N_11539,N_10514,N_11125);
nand U11540 (N_11540,N_10568,N_11001);
nor U11541 (N_11541,N_11018,N_10909);
and U11542 (N_11542,N_11153,N_10817);
nand U11543 (N_11543,N_10702,N_11233);
or U11544 (N_11544,N_11043,N_11032);
nand U11545 (N_11545,N_10806,N_10757);
xor U11546 (N_11546,N_10846,N_10629);
nor U11547 (N_11547,N_10885,N_10726);
or U11548 (N_11548,N_11039,N_10869);
and U11549 (N_11549,N_10585,N_10760);
and U11550 (N_11550,N_10864,N_11083);
nand U11551 (N_11551,N_10914,N_10916);
nor U11552 (N_11552,N_11188,N_11145);
and U11553 (N_11553,N_10571,N_10508);
or U11554 (N_11554,N_11210,N_10920);
xnor U11555 (N_11555,N_10975,N_10939);
nand U11556 (N_11556,N_10567,N_10520);
or U11557 (N_11557,N_10546,N_10587);
xnor U11558 (N_11558,N_10695,N_11115);
nand U11559 (N_11559,N_10976,N_10661);
or U11560 (N_11560,N_10737,N_10606);
and U11561 (N_11561,N_10851,N_10584);
and U11562 (N_11562,N_11016,N_10989);
or U11563 (N_11563,N_10710,N_10583);
or U11564 (N_11564,N_10937,N_10658);
xor U11565 (N_11565,N_10842,N_10980);
nand U11566 (N_11566,N_11025,N_11162);
and U11567 (N_11567,N_11116,N_11030);
and U11568 (N_11568,N_10898,N_10960);
nand U11569 (N_11569,N_10614,N_11123);
xor U11570 (N_11570,N_10633,N_10590);
and U11571 (N_11571,N_11050,N_10947);
nand U11572 (N_11572,N_11134,N_10609);
nand U11573 (N_11573,N_10582,N_10720);
and U11574 (N_11574,N_11031,N_10539);
nand U11575 (N_11575,N_10798,N_11194);
nand U11576 (N_11576,N_10879,N_11148);
and U11577 (N_11577,N_10743,N_10653);
nand U11578 (N_11578,N_11128,N_10995);
nand U11579 (N_11579,N_10537,N_10616);
nand U11580 (N_11580,N_10877,N_11063);
and U11581 (N_11581,N_11245,N_10513);
or U11582 (N_11582,N_11216,N_10908);
or U11583 (N_11583,N_10709,N_10551);
nor U11584 (N_11584,N_11150,N_10731);
nand U11585 (N_11585,N_10595,N_10867);
nor U11586 (N_11586,N_10524,N_10504);
nand U11587 (N_11587,N_10992,N_10628);
or U11588 (N_11588,N_10692,N_10500);
and U11589 (N_11589,N_11218,N_11041);
xor U11590 (N_11590,N_10740,N_10951);
xor U11591 (N_11591,N_10649,N_10994);
nand U11592 (N_11592,N_10805,N_11113);
nor U11593 (N_11593,N_10893,N_10943);
or U11594 (N_11594,N_10784,N_10868);
and U11595 (N_11595,N_10588,N_10700);
nor U11596 (N_11596,N_10814,N_10662);
xor U11597 (N_11597,N_11165,N_10781);
and U11598 (N_11598,N_10758,N_11020);
or U11599 (N_11599,N_10950,N_11191);
or U11600 (N_11600,N_10694,N_10527);
nand U11601 (N_11601,N_11075,N_10697);
nand U11602 (N_11602,N_10801,N_10608);
or U11603 (N_11603,N_10789,N_11178);
nand U11604 (N_11604,N_10875,N_10733);
nor U11605 (N_11605,N_10929,N_10530);
or U11606 (N_11606,N_11044,N_10739);
xnor U11607 (N_11607,N_10652,N_11121);
or U11608 (N_11608,N_10935,N_10892);
and U11609 (N_11609,N_11102,N_11119);
or U11610 (N_11610,N_11230,N_10990);
and U11611 (N_11611,N_10876,N_10823);
nor U11612 (N_11612,N_10669,N_10523);
nand U11613 (N_11613,N_10872,N_10780);
or U11614 (N_11614,N_10961,N_10646);
and U11615 (N_11615,N_10922,N_11231);
nand U11616 (N_11616,N_11029,N_11193);
or U11617 (N_11617,N_10847,N_10555);
xnor U11618 (N_11618,N_10772,N_11105);
and U11619 (N_11619,N_11002,N_11036);
or U11620 (N_11620,N_10890,N_10706);
nor U11621 (N_11621,N_10829,N_10900);
nor U11622 (N_11622,N_10736,N_10941);
nor U11623 (N_11623,N_10621,N_10754);
nor U11624 (N_11624,N_10682,N_10638);
or U11625 (N_11625,N_10797,N_10798);
nand U11626 (N_11626,N_10752,N_11189);
nand U11627 (N_11627,N_10835,N_11025);
nor U11628 (N_11628,N_10701,N_10890);
or U11629 (N_11629,N_10644,N_10734);
nor U11630 (N_11630,N_10737,N_10787);
nand U11631 (N_11631,N_10558,N_10594);
or U11632 (N_11632,N_10665,N_10715);
or U11633 (N_11633,N_10649,N_11016);
xnor U11634 (N_11634,N_10671,N_11192);
and U11635 (N_11635,N_10596,N_10804);
or U11636 (N_11636,N_10931,N_10824);
and U11637 (N_11637,N_11045,N_11170);
or U11638 (N_11638,N_10521,N_10840);
and U11639 (N_11639,N_11205,N_10591);
nand U11640 (N_11640,N_10838,N_10913);
nand U11641 (N_11641,N_10910,N_11041);
xnor U11642 (N_11642,N_10772,N_10978);
nand U11643 (N_11643,N_11045,N_10895);
and U11644 (N_11644,N_10793,N_11235);
and U11645 (N_11645,N_11132,N_11156);
nor U11646 (N_11646,N_10877,N_11074);
nand U11647 (N_11647,N_10600,N_10682);
nand U11648 (N_11648,N_10660,N_10975);
nor U11649 (N_11649,N_10831,N_10655);
or U11650 (N_11650,N_10866,N_11189);
nand U11651 (N_11651,N_11055,N_10747);
or U11652 (N_11652,N_10514,N_11103);
or U11653 (N_11653,N_10986,N_10592);
nor U11654 (N_11654,N_10692,N_10620);
xnor U11655 (N_11655,N_10684,N_11019);
nor U11656 (N_11656,N_10908,N_11246);
nand U11657 (N_11657,N_10753,N_11078);
xnor U11658 (N_11658,N_11199,N_11154);
nor U11659 (N_11659,N_10929,N_11060);
nor U11660 (N_11660,N_11005,N_10632);
and U11661 (N_11661,N_11024,N_10894);
nor U11662 (N_11662,N_10796,N_10952);
nand U11663 (N_11663,N_11070,N_10652);
and U11664 (N_11664,N_10581,N_10705);
or U11665 (N_11665,N_10818,N_10966);
and U11666 (N_11666,N_10524,N_10828);
and U11667 (N_11667,N_10960,N_10982);
nand U11668 (N_11668,N_10759,N_11069);
nand U11669 (N_11669,N_10795,N_10656);
or U11670 (N_11670,N_10584,N_10731);
nor U11671 (N_11671,N_11144,N_11043);
nand U11672 (N_11672,N_10698,N_11166);
nor U11673 (N_11673,N_10660,N_11135);
and U11674 (N_11674,N_10922,N_10701);
and U11675 (N_11675,N_10801,N_10536);
nor U11676 (N_11676,N_10844,N_10563);
nand U11677 (N_11677,N_11154,N_11057);
or U11678 (N_11678,N_10912,N_10748);
and U11679 (N_11679,N_10659,N_11017);
nand U11680 (N_11680,N_11130,N_10638);
nor U11681 (N_11681,N_11095,N_10673);
nand U11682 (N_11682,N_10978,N_11167);
or U11683 (N_11683,N_10826,N_11057);
nand U11684 (N_11684,N_10766,N_10697);
xnor U11685 (N_11685,N_10881,N_11040);
xor U11686 (N_11686,N_10579,N_10907);
and U11687 (N_11687,N_10994,N_10816);
nand U11688 (N_11688,N_11119,N_10620);
nor U11689 (N_11689,N_11223,N_10880);
xor U11690 (N_11690,N_11143,N_11056);
xnor U11691 (N_11691,N_10819,N_10988);
nor U11692 (N_11692,N_10720,N_10833);
xnor U11693 (N_11693,N_10698,N_10928);
xnor U11694 (N_11694,N_10707,N_11135);
nand U11695 (N_11695,N_11039,N_10929);
xor U11696 (N_11696,N_10527,N_11002);
and U11697 (N_11697,N_10771,N_10695);
nand U11698 (N_11698,N_10518,N_11178);
or U11699 (N_11699,N_10981,N_11174);
nor U11700 (N_11700,N_10603,N_11204);
and U11701 (N_11701,N_10797,N_11213);
xnor U11702 (N_11702,N_10981,N_10729);
nor U11703 (N_11703,N_10783,N_10823);
nand U11704 (N_11704,N_10581,N_11095);
and U11705 (N_11705,N_10581,N_10774);
nor U11706 (N_11706,N_11059,N_10865);
nor U11707 (N_11707,N_11017,N_10636);
nand U11708 (N_11708,N_10825,N_10662);
and U11709 (N_11709,N_10961,N_10655);
xor U11710 (N_11710,N_10857,N_10787);
xnor U11711 (N_11711,N_10605,N_10968);
nand U11712 (N_11712,N_10734,N_10571);
xnor U11713 (N_11713,N_10575,N_11114);
nor U11714 (N_11714,N_10876,N_11215);
nand U11715 (N_11715,N_10582,N_10809);
nor U11716 (N_11716,N_11053,N_10960);
or U11717 (N_11717,N_10608,N_11123);
nor U11718 (N_11718,N_10677,N_10582);
nor U11719 (N_11719,N_11072,N_10725);
xor U11720 (N_11720,N_10801,N_11144);
nor U11721 (N_11721,N_10801,N_10831);
and U11722 (N_11722,N_10836,N_10950);
or U11723 (N_11723,N_11113,N_10544);
nand U11724 (N_11724,N_10924,N_10844);
or U11725 (N_11725,N_10889,N_11123);
nor U11726 (N_11726,N_11165,N_11133);
nand U11727 (N_11727,N_10553,N_11068);
and U11728 (N_11728,N_10687,N_10756);
and U11729 (N_11729,N_11131,N_11092);
or U11730 (N_11730,N_10581,N_11150);
nand U11731 (N_11731,N_11092,N_11111);
xor U11732 (N_11732,N_10787,N_11077);
xor U11733 (N_11733,N_11183,N_10699);
or U11734 (N_11734,N_11104,N_10600);
nand U11735 (N_11735,N_11153,N_10899);
nor U11736 (N_11736,N_11128,N_10705);
xor U11737 (N_11737,N_11200,N_11142);
and U11738 (N_11738,N_10975,N_10600);
and U11739 (N_11739,N_10618,N_11041);
nand U11740 (N_11740,N_10970,N_11040);
and U11741 (N_11741,N_10964,N_10776);
and U11742 (N_11742,N_10579,N_11243);
xnor U11743 (N_11743,N_10821,N_10790);
nand U11744 (N_11744,N_11058,N_10783);
or U11745 (N_11745,N_11141,N_10639);
or U11746 (N_11746,N_10605,N_10971);
nand U11747 (N_11747,N_10541,N_10502);
and U11748 (N_11748,N_10785,N_10534);
and U11749 (N_11749,N_10848,N_10664);
nand U11750 (N_11750,N_10556,N_10513);
and U11751 (N_11751,N_11085,N_10627);
or U11752 (N_11752,N_10671,N_10916);
or U11753 (N_11753,N_10861,N_11206);
and U11754 (N_11754,N_10909,N_11221);
nor U11755 (N_11755,N_10574,N_11166);
nor U11756 (N_11756,N_10858,N_11094);
nand U11757 (N_11757,N_10548,N_10839);
and U11758 (N_11758,N_11073,N_11248);
xor U11759 (N_11759,N_11237,N_10826);
xnor U11760 (N_11760,N_11007,N_10906);
nor U11761 (N_11761,N_10873,N_11025);
and U11762 (N_11762,N_10755,N_10667);
or U11763 (N_11763,N_10788,N_10945);
xnor U11764 (N_11764,N_10664,N_11173);
and U11765 (N_11765,N_11002,N_10700);
or U11766 (N_11766,N_10538,N_10937);
and U11767 (N_11767,N_10672,N_10784);
xnor U11768 (N_11768,N_10608,N_11248);
or U11769 (N_11769,N_10934,N_10537);
nand U11770 (N_11770,N_11002,N_10550);
or U11771 (N_11771,N_10519,N_11140);
or U11772 (N_11772,N_10810,N_10956);
nor U11773 (N_11773,N_11126,N_10745);
nand U11774 (N_11774,N_11126,N_11243);
or U11775 (N_11775,N_10691,N_10681);
nand U11776 (N_11776,N_10995,N_11211);
xor U11777 (N_11777,N_10833,N_10520);
and U11778 (N_11778,N_10564,N_11115);
xnor U11779 (N_11779,N_10891,N_11210);
nor U11780 (N_11780,N_10952,N_10640);
nand U11781 (N_11781,N_10998,N_10664);
and U11782 (N_11782,N_10603,N_11001);
nand U11783 (N_11783,N_10584,N_11185);
xor U11784 (N_11784,N_10741,N_11099);
and U11785 (N_11785,N_11191,N_11000);
and U11786 (N_11786,N_10826,N_10808);
xor U11787 (N_11787,N_10640,N_10595);
nor U11788 (N_11788,N_10909,N_11186);
nand U11789 (N_11789,N_10978,N_10593);
xnor U11790 (N_11790,N_10749,N_10617);
and U11791 (N_11791,N_11163,N_11226);
or U11792 (N_11792,N_10865,N_10839);
nor U11793 (N_11793,N_10897,N_10543);
or U11794 (N_11794,N_10670,N_11128);
and U11795 (N_11795,N_10582,N_11045);
nand U11796 (N_11796,N_10938,N_11132);
or U11797 (N_11797,N_10912,N_10766);
and U11798 (N_11798,N_10956,N_10910);
nand U11799 (N_11799,N_10915,N_11133);
and U11800 (N_11800,N_10923,N_11052);
nor U11801 (N_11801,N_11078,N_11124);
nand U11802 (N_11802,N_10811,N_10965);
xnor U11803 (N_11803,N_11233,N_10930);
nor U11804 (N_11804,N_11005,N_11172);
or U11805 (N_11805,N_11067,N_11208);
nand U11806 (N_11806,N_11206,N_11185);
or U11807 (N_11807,N_11002,N_10725);
nor U11808 (N_11808,N_10775,N_11126);
and U11809 (N_11809,N_10510,N_10704);
xor U11810 (N_11810,N_10733,N_11194);
nor U11811 (N_11811,N_10619,N_10878);
nor U11812 (N_11812,N_10876,N_11094);
xor U11813 (N_11813,N_10629,N_10636);
nor U11814 (N_11814,N_11097,N_10991);
and U11815 (N_11815,N_10916,N_10918);
and U11816 (N_11816,N_10767,N_10751);
or U11817 (N_11817,N_11016,N_10603);
nand U11818 (N_11818,N_11086,N_11133);
or U11819 (N_11819,N_10938,N_10757);
nor U11820 (N_11820,N_10908,N_10586);
nor U11821 (N_11821,N_10689,N_10989);
nor U11822 (N_11822,N_10551,N_10956);
or U11823 (N_11823,N_11242,N_10924);
nand U11824 (N_11824,N_10562,N_10861);
nor U11825 (N_11825,N_11172,N_10920);
nor U11826 (N_11826,N_10510,N_10690);
nor U11827 (N_11827,N_10619,N_10589);
nor U11828 (N_11828,N_11147,N_10679);
xnor U11829 (N_11829,N_10754,N_11024);
and U11830 (N_11830,N_10789,N_11067);
or U11831 (N_11831,N_11204,N_11180);
or U11832 (N_11832,N_10519,N_11128);
or U11833 (N_11833,N_10651,N_10546);
nor U11834 (N_11834,N_11030,N_11039);
or U11835 (N_11835,N_10790,N_11237);
nor U11836 (N_11836,N_10706,N_10661);
or U11837 (N_11837,N_10619,N_10991);
or U11838 (N_11838,N_10850,N_11009);
xnor U11839 (N_11839,N_10734,N_10560);
or U11840 (N_11840,N_10873,N_11118);
nor U11841 (N_11841,N_11019,N_11212);
and U11842 (N_11842,N_10793,N_11025);
nor U11843 (N_11843,N_11228,N_10933);
or U11844 (N_11844,N_10692,N_10891);
nand U11845 (N_11845,N_10504,N_11027);
and U11846 (N_11846,N_10617,N_11033);
and U11847 (N_11847,N_11248,N_10639);
xnor U11848 (N_11848,N_11072,N_10862);
or U11849 (N_11849,N_11083,N_11205);
nor U11850 (N_11850,N_11178,N_10927);
or U11851 (N_11851,N_10731,N_11214);
or U11852 (N_11852,N_11113,N_11241);
or U11853 (N_11853,N_10776,N_11157);
nor U11854 (N_11854,N_10618,N_10841);
nand U11855 (N_11855,N_10721,N_11041);
xnor U11856 (N_11856,N_10880,N_10514);
or U11857 (N_11857,N_10785,N_11056);
and U11858 (N_11858,N_10682,N_10740);
and U11859 (N_11859,N_11013,N_11026);
or U11860 (N_11860,N_10747,N_10854);
and U11861 (N_11861,N_10943,N_11202);
nor U11862 (N_11862,N_10513,N_10572);
xor U11863 (N_11863,N_11096,N_10567);
and U11864 (N_11864,N_10662,N_11009);
nor U11865 (N_11865,N_11129,N_10676);
and U11866 (N_11866,N_10931,N_10728);
nand U11867 (N_11867,N_10967,N_10879);
and U11868 (N_11868,N_10948,N_11187);
xor U11869 (N_11869,N_10947,N_10859);
nand U11870 (N_11870,N_10975,N_10727);
nand U11871 (N_11871,N_10756,N_10706);
or U11872 (N_11872,N_11089,N_11069);
nor U11873 (N_11873,N_10642,N_10876);
nor U11874 (N_11874,N_11154,N_11068);
xor U11875 (N_11875,N_10991,N_10938);
nor U11876 (N_11876,N_10969,N_10694);
or U11877 (N_11877,N_10947,N_10794);
or U11878 (N_11878,N_10503,N_10779);
and U11879 (N_11879,N_10755,N_11096);
or U11880 (N_11880,N_10961,N_11112);
nand U11881 (N_11881,N_11062,N_10615);
and U11882 (N_11882,N_10707,N_11111);
and U11883 (N_11883,N_10766,N_10600);
xnor U11884 (N_11884,N_10922,N_11149);
nor U11885 (N_11885,N_11049,N_10587);
nor U11886 (N_11886,N_10989,N_11008);
nor U11887 (N_11887,N_10893,N_10844);
or U11888 (N_11888,N_10543,N_11153);
xor U11889 (N_11889,N_11241,N_11211);
and U11890 (N_11890,N_10725,N_11220);
nor U11891 (N_11891,N_11217,N_11238);
nand U11892 (N_11892,N_10697,N_11167);
nand U11893 (N_11893,N_11117,N_10749);
and U11894 (N_11894,N_10944,N_11140);
nor U11895 (N_11895,N_11024,N_10652);
nor U11896 (N_11896,N_10800,N_11000);
or U11897 (N_11897,N_10958,N_10943);
nand U11898 (N_11898,N_11076,N_10950);
and U11899 (N_11899,N_10939,N_10683);
nor U11900 (N_11900,N_11039,N_10936);
and U11901 (N_11901,N_10662,N_10927);
nor U11902 (N_11902,N_10833,N_10844);
and U11903 (N_11903,N_11075,N_10760);
xor U11904 (N_11904,N_10936,N_10882);
nand U11905 (N_11905,N_10681,N_10827);
and U11906 (N_11906,N_11103,N_10929);
nor U11907 (N_11907,N_10848,N_11001);
or U11908 (N_11908,N_10881,N_11231);
nand U11909 (N_11909,N_10507,N_10548);
and U11910 (N_11910,N_11030,N_10728);
or U11911 (N_11911,N_10715,N_11014);
and U11912 (N_11912,N_10931,N_10558);
nor U11913 (N_11913,N_10547,N_10869);
and U11914 (N_11914,N_10902,N_10964);
nand U11915 (N_11915,N_10910,N_10758);
nand U11916 (N_11916,N_10604,N_10587);
and U11917 (N_11917,N_10961,N_10690);
and U11918 (N_11918,N_10970,N_10636);
nand U11919 (N_11919,N_10852,N_10885);
nand U11920 (N_11920,N_10564,N_10599);
nor U11921 (N_11921,N_10881,N_11083);
and U11922 (N_11922,N_10970,N_10794);
or U11923 (N_11923,N_10548,N_10979);
nor U11924 (N_11924,N_11243,N_10733);
or U11925 (N_11925,N_10903,N_10815);
or U11926 (N_11926,N_10594,N_11195);
nor U11927 (N_11927,N_11023,N_10717);
nand U11928 (N_11928,N_10820,N_10672);
and U11929 (N_11929,N_10613,N_11215);
nand U11930 (N_11930,N_10906,N_11121);
xnor U11931 (N_11931,N_11123,N_10688);
xnor U11932 (N_11932,N_10666,N_11134);
nand U11933 (N_11933,N_10931,N_10661);
nor U11934 (N_11934,N_11146,N_10599);
and U11935 (N_11935,N_11061,N_10871);
or U11936 (N_11936,N_10569,N_10589);
and U11937 (N_11937,N_10713,N_10863);
xnor U11938 (N_11938,N_10764,N_10517);
nor U11939 (N_11939,N_10824,N_11017);
and U11940 (N_11940,N_11054,N_11139);
nor U11941 (N_11941,N_11195,N_11062);
and U11942 (N_11942,N_10882,N_11082);
and U11943 (N_11943,N_10799,N_10727);
or U11944 (N_11944,N_10571,N_10712);
or U11945 (N_11945,N_10926,N_10938);
nor U11946 (N_11946,N_10578,N_10880);
or U11947 (N_11947,N_11061,N_10815);
nor U11948 (N_11948,N_11170,N_10792);
nand U11949 (N_11949,N_10566,N_10927);
nand U11950 (N_11950,N_10636,N_11105);
nand U11951 (N_11951,N_10750,N_11028);
or U11952 (N_11952,N_10510,N_10706);
and U11953 (N_11953,N_10900,N_10574);
or U11954 (N_11954,N_10759,N_10503);
or U11955 (N_11955,N_10997,N_10674);
or U11956 (N_11956,N_10921,N_10704);
or U11957 (N_11957,N_10714,N_10607);
nand U11958 (N_11958,N_10715,N_10684);
nor U11959 (N_11959,N_10722,N_10503);
nand U11960 (N_11960,N_11150,N_11060);
and U11961 (N_11961,N_10975,N_11152);
nand U11962 (N_11962,N_10684,N_11210);
nor U11963 (N_11963,N_11237,N_10576);
and U11964 (N_11964,N_10992,N_11086);
and U11965 (N_11965,N_10723,N_10779);
or U11966 (N_11966,N_10633,N_11192);
nor U11967 (N_11967,N_11071,N_10640);
or U11968 (N_11968,N_10658,N_10765);
nor U11969 (N_11969,N_10562,N_10834);
nand U11970 (N_11970,N_10707,N_10923);
nand U11971 (N_11971,N_10864,N_11199);
and U11972 (N_11972,N_10904,N_10566);
nand U11973 (N_11973,N_10704,N_11088);
nand U11974 (N_11974,N_10960,N_10828);
or U11975 (N_11975,N_11037,N_10910);
and U11976 (N_11976,N_10808,N_11007);
and U11977 (N_11977,N_11115,N_10966);
or U11978 (N_11978,N_11161,N_10586);
nand U11979 (N_11979,N_10846,N_10641);
or U11980 (N_11980,N_10541,N_11002);
xor U11981 (N_11981,N_10909,N_10882);
nand U11982 (N_11982,N_10960,N_10954);
nor U11983 (N_11983,N_10767,N_10766);
and U11984 (N_11984,N_11171,N_11126);
and U11985 (N_11985,N_10749,N_10921);
nor U11986 (N_11986,N_10903,N_10650);
or U11987 (N_11987,N_11019,N_11011);
and U11988 (N_11988,N_11024,N_10688);
or U11989 (N_11989,N_11091,N_10937);
or U11990 (N_11990,N_11062,N_10502);
or U11991 (N_11991,N_11141,N_10969);
or U11992 (N_11992,N_10959,N_10889);
nor U11993 (N_11993,N_10765,N_10885);
and U11994 (N_11994,N_10864,N_10600);
nor U11995 (N_11995,N_10615,N_10832);
and U11996 (N_11996,N_11200,N_11042);
nand U11997 (N_11997,N_10761,N_10557);
nor U11998 (N_11998,N_10567,N_11020);
or U11999 (N_11999,N_10825,N_10549);
and U12000 (N_12000,N_11945,N_11693);
or U12001 (N_12001,N_11717,N_11975);
nand U12002 (N_12002,N_11325,N_11802);
nand U12003 (N_12003,N_11999,N_11702);
nand U12004 (N_12004,N_11437,N_11995);
and U12005 (N_12005,N_11668,N_11792);
or U12006 (N_12006,N_11314,N_11286);
and U12007 (N_12007,N_11615,N_11515);
and U12008 (N_12008,N_11973,N_11295);
nor U12009 (N_12009,N_11337,N_11559);
nor U12010 (N_12010,N_11639,N_11871);
nor U12011 (N_12011,N_11277,N_11330);
nor U12012 (N_12012,N_11591,N_11268);
nand U12013 (N_12013,N_11416,N_11952);
xor U12014 (N_12014,N_11569,N_11968);
nand U12015 (N_12015,N_11431,N_11393);
or U12016 (N_12016,N_11498,N_11819);
and U12017 (N_12017,N_11442,N_11827);
nand U12018 (N_12018,N_11430,N_11478);
nor U12019 (N_12019,N_11421,N_11598);
and U12020 (N_12020,N_11327,N_11950);
xnor U12021 (N_12021,N_11949,N_11824);
or U12022 (N_12022,N_11989,N_11537);
nand U12023 (N_12023,N_11705,N_11874);
nor U12024 (N_12024,N_11524,N_11374);
nand U12025 (N_12025,N_11879,N_11650);
nor U12026 (N_12026,N_11407,N_11508);
nor U12027 (N_12027,N_11788,N_11310);
and U12028 (N_12028,N_11730,N_11673);
nor U12029 (N_12029,N_11954,N_11993);
nand U12030 (N_12030,N_11371,N_11605);
nor U12031 (N_12031,N_11872,N_11542);
and U12032 (N_12032,N_11332,N_11358);
and U12033 (N_12033,N_11625,N_11721);
nand U12034 (N_12034,N_11386,N_11804);
nor U12035 (N_12035,N_11587,N_11632);
or U12036 (N_12036,N_11775,N_11379);
or U12037 (N_12037,N_11748,N_11820);
or U12038 (N_12038,N_11494,N_11613);
xor U12039 (N_12039,N_11671,N_11831);
nand U12040 (N_12040,N_11341,N_11397);
or U12041 (N_12041,N_11688,N_11758);
or U12042 (N_12042,N_11479,N_11271);
and U12043 (N_12043,N_11511,N_11724);
or U12044 (N_12044,N_11739,N_11510);
or U12045 (N_12045,N_11536,N_11331);
nand U12046 (N_12046,N_11847,N_11518);
xor U12047 (N_12047,N_11911,N_11500);
and U12048 (N_12048,N_11336,N_11453);
nand U12049 (N_12049,N_11828,N_11714);
or U12050 (N_12050,N_11311,N_11813);
nand U12051 (N_12051,N_11365,N_11880);
xor U12052 (N_12052,N_11313,N_11641);
nor U12053 (N_12053,N_11791,N_11335);
nor U12054 (N_12054,N_11990,N_11533);
and U12055 (N_12055,N_11571,N_11996);
nand U12056 (N_12056,N_11750,N_11502);
or U12057 (N_12057,N_11894,N_11535);
nor U12058 (N_12058,N_11596,N_11812);
nand U12059 (N_12059,N_11583,N_11710);
nor U12060 (N_12060,N_11390,N_11763);
nand U12061 (N_12061,N_11377,N_11556);
nand U12062 (N_12062,N_11944,N_11723);
nand U12063 (N_12063,N_11998,N_11823);
and U12064 (N_12064,N_11637,N_11910);
nor U12065 (N_12065,N_11577,N_11438);
or U12066 (N_12066,N_11662,N_11432);
nand U12067 (N_12067,N_11830,N_11617);
nand U12068 (N_12068,N_11261,N_11259);
and U12069 (N_12069,N_11741,N_11581);
nand U12070 (N_12070,N_11356,N_11713);
xnor U12071 (N_12071,N_11939,N_11808);
and U12072 (N_12072,N_11983,N_11903);
or U12073 (N_12073,N_11593,N_11987);
or U12074 (N_12074,N_11686,N_11833);
or U12075 (N_12075,N_11660,N_11285);
nor U12076 (N_12076,N_11404,N_11633);
and U12077 (N_12077,N_11951,N_11287);
and U12078 (N_12078,N_11980,N_11921);
or U12079 (N_12079,N_11564,N_11448);
nor U12080 (N_12080,N_11849,N_11561);
nand U12081 (N_12081,N_11289,N_11928);
nand U12082 (N_12082,N_11863,N_11842);
nand U12083 (N_12083,N_11636,N_11651);
nand U12084 (N_12084,N_11736,N_11489);
or U12085 (N_12085,N_11252,N_11811);
xnor U12086 (N_12086,N_11899,N_11405);
nand U12087 (N_12087,N_11452,N_11606);
or U12088 (N_12088,N_11882,N_11917);
nor U12089 (N_12089,N_11519,N_11909);
and U12090 (N_12090,N_11343,N_11659);
nand U12091 (N_12091,N_11580,N_11349);
nand U12092 (N_12092,N_11565,N_11434);
and U12093 (N_12093,N_11265,N_11395);
or U12094 (N_12094,N_11752,N_11915);
or U12095 (N_12095,N_11256,N_11982);
nand U12096 (N_12096,N_11316,N_11684);
and U12097 (N_12097,N_11406,N_11733);
or U12098 (N_12098,N_11756,N_11441);
nor U12099 (N_12099,N_11822,N_11677);
nor U12100 (N_12100,N_11608,N_11427);
and U12101 (N_12101,N_11992,N_11957);
and U12102 (N_12102,N_11366,N_11491);
or U12103 (N_12103,N_11937,N_11582);
and U12104 (N_12104,N_11844,N_11918);
xnor U12105 (N_12105,N_11906,N_11302);
nand U12106 (N_12106,N_11644,N_11679);
nor U12107 (N_12107,N_11279,N_11898);
nor U12108 (N_12108,N_11293,N_11925);
nor U12109 (N_12109,N_11454,N_11436);
nor U12110 (N_12110,N_11317,N_11887);
nand U12111 (N_12111,N_11435,N_11514);
nor U12112 (N_12112,N_11751,N_11594);
or U12113 (N_12113,N_11692,N_11720);
and U12114 (N_12114,N_11426,N_11482);
nand U12115 (N_12115,N_11548,N_11912);
nand U12116 (N_12116,N_11778,N_11428);
xnor U12117 (N_12117,N_11324,N_11509);
and U12118 (N_12118,N_11297,N_11661);
or U12119 (N_12119,N_11300,N_11786);
and U12120 (N_12120,N_11943,N_11584);
nor U12121 (N_12121,N_11487,N_11676);
nand U12122 (N_12122,N_11984,N_11450);
nor U12123 (N_12123,N_11318,N_11412);
or U12124 (N_12124,N_11866,N_11868);
xnor U12125 (N_12125,N_11744,N_11635);
and U12126 (N_12126,N_11706,N_11503);
nand U12127 (N_12127,N_11532,N_11303);
nand U12128 (N_12128,N_11653,N_11463);
or U12129 (N_12129,N_11781,N_11601);
nand U12130 (N_12130,N_11839,N_11718);
or U12131 (N_12131,N_11904,N_11762);
and U12132 (N_12132,N_11770,N_11609);
or U12133 (N_12133,N_11779,N_11628);
or U12134 (N_12134,N_11381,N_11892);
nand U12135 (N_12135,N_11607,N_11418);
xnor U12136 (N_12136,N_11339,N_11328);
nor U12137 (N_12137,N_11398,N_11563);
nor U12138 (N_12138,N_11321,N_11704);
or U12139 (N_12139,N_11576,N_11782);
nor U12140 (N_12140,N_11354,N_11664);
or U12141 (N_12141,N_11364,N_11629);
or U12142 (N_12142,N_11965,N_11308);
nor U12143 (N_12143,N_11930,N_11709);
nor U12144 (N_12144,N_11496,N_11986);
and U12145 (N_12145,N_11767,N_11886);
xor U12146 (N_12146,N_11976,N_11274);
and U12147 (N_12147,N_11391,N_11760);
nand U12148 (N_12148,N_11858,N_11807);
or U12149 (N_12149,N_11678,N_11864);
xor U12150 (N_12150,N_11806,N_11888);
xnor U12151 (N_12151,N_11440,N_11459);
or U12152 (N_12152,N_11852,N_11988);
nor U12153 (N_12153,N_11488,N_11712);
nor U12154 (N_12154,N_11857,N_11815);
or U12155 (N_12155,N_11549,N_11768);
nor U12156 (N_12156,N_11447,N_11838);
nand U12157 (N_12157,N_11455,N_11264);
nand U12158 (N_12158,N_11270,N_11350);
and U12159 (N_12159,N_11298,N_11338);
and U12160 (N_12160,N_11610,N_11665);
nand U12161 (N_12161,N_11408,N_11738);
nor U12162 (N_12162,N_11375,N_11497);
and U12163 (N_12163,N_11818,N_11296);
and U12164 (N_12164,N_11855,N_11357);
xor U12165 (N_12165,N_11588,N_11630);
nand U12166 (N_12166,N_11785,N_11516);
and U12167 (N_12167,N_11645,N_11716);
nand U12168 (N_12168,N_11443,N_11810);
and U12169 (N_12169,N_11936,N_11380);
nand U12170 (N_12170,N_11687,N_11616);
nor U12171 (N_12171,N_11470,N_11856);
nor U12172 (N_12172,N_11322,N_11618);
nor U12173 (N_12173,N_11970,N_11257);
xnor U12174 (N_12174,N_11955,N_11919);
xnor U12175 (N_12175,N_11326,N_11732);
nand U12176 (N_12176,N_11734,N_11423);
nand U12177 (N_12177,N_11929,N_11825);
nand U12178 (N_12178,N_11590,N_11425);
or U12179 (N_12179,N_11315,N_11280);
nand U12180 (N_12180,N_11319,N_11623);
and U12181 (N_12181,N_11586,N_11926);
or U12182 (N_12182,N_11603,N_11743);
nand U12183 (N_12183,N_11708,N_11520);
nor U12184 (N_12184,N_11773,N_11527);
nor U12185 (N_12185,N_11384,N_11490);
or U12186 (N_12186,N_11964,N_11776);
and U12187 (N_12187,N_11578,N_11460);
nor U12188 (N_12188,N_11541,N_11495);
nand U12189 (N_12189,N_11893,N_11790);
nand U12190 (N_12190,N_11814,N_11891);
nor U12191 (N_12191,N_11355,N_11877);
nand U12192 (N_12192,N_11931,N_11846);
and U12193 (N_12193,N_11994,N_11747);
and U12194 (N_12194,N_11753,N_11638);
and U12195 (N_12195,N_11534,N_11777);
and U12196 (N_12196,N_11640,N_11570);
or U12197 (N_12197,N_11251,N_11461);
nand U12198 (N_12198,N_11348,N_11344);
nand U12199 (N_12199,N_11938,N_11794);
and U12200 (N_12200,N_11648,N_11729);
nor U12201 (N_12201,N_11359,N_11560);
xnor U12202 (N_12202,N_11922,N_11622);
or U12203 (N_12203,N_11991,N_11263);
nor U12204 (N_12204,N_11544,N_11410);
and U12205 (N_12205,N_11961,N_11875);
nor U12206 (N_12206,N_11935,N_11283);
nand U12207 (N_12207,N_11740,N_11468);
and U12208 (N_12208,N_11558,N_11415);
nor U12209 (N_12209,N_11974,N_11419);
nor U12210 (N_12210,N_11731,N_11306);
and U12211 (N_12211,N_11481,N_11834);
or U12212 (N_12212,N_11553,N_11799);
and U12213 (N_12213,N_11985,N_11614);
and U12214 (N_12214,N_11837,N_11552);
and U12215 (N_12215,N_11663,N_11890);
xor U12216 (N_12216,N_11728,N_11977);
nand U12217 (N_12217,N_11528,N_11884);
nand U12218 (N_12218,N_11764,N_11387);
and U12219 (N_12219,N_11798,N_11826);
and U12220 (N_12220,N_11787,N_11870);
nor U12221 (N_12221,N_11626,N_11567);
and U12222 (N_12222,N_11631,N_11372);
nand U12223 (N_12223,N_11299,N_11531);
or U12224 (N_12224,N_11845,N_11550);
or U12225 (N_12225,N_11486,N_11557);
nand U12226 (N_12226,N_11471,N_11670);
or U12227 (N_12227,N_11889,N_11963);
nor U12228 (N_12228,N_11475,N_11255);
and U12229 (N_12229,N_11881,N_11462);
and U12230 (N_12230,N_11924,N_11682);
nand U12231 (N_12231,N_11554,N_11658);
and U12232 (N_12232,N_11476,N_11288);
and U12233 (N_12233,N_11953,N_11429);
and U12234 (N_12234,N_11967,N_11267);
xor U12235 (N_12235,N_11346,N_11843);
nand U12236 (N_12236,N_11755,N_11378);
nor U12237 (N_12237,N_11522,N_11969);
and U12238 (N_12238,N_11449,N_11273);
and U12239 (N_12239,N_11643,N_11342);
xor U12240 (N_12240,N_11269,N_11451);
xnor U12241 (N_12241,N_11484,N_11568);
or U12242 (N_12242,N_11897,N_11262);
xor U12243 (N_12243,N_11853,N_11333);
and U12244 (N_12244,N_11701,N_11759);
nand U12245 (N_12245,N_11941,N_11674);
and U12246 (N_12246,N_11766,N_11424);
nor U12247 (N_12247,N_11396,N_11546);
or U12248 (N_12248,N_11499,N_11652);
nand U12249 (N_12249,N_11281,N_11551);
xnor U12250 (N_12250,N_11654,N_11361);
nand U12251 (N_12251,N_11388,N_11477);
and U12252 (N_12252,N_11932,N_11507);
nor U12253 (N_12253,N_11320,N_11895);
and U12254 (N_12254,N_11352,N_11707);
nand U12255 (N_12255,N_11646,N_11727);
nand U12256 (N_12256,N_11681,N_11627);
or U12257 (N_12257,N_11885,N_11647);
and U12258 (N_12258,N_11504,N_11719);
nor U12259 (N_12259,N_11699,N_11749);
nand U12260 (N_12260,N_11848,N_11275);
nand U12261 (N_12261,N_11445,N_11526);
or U12262 (N_12262,N_11923,N_11278);
and U12263 (N_12263,N_11914,N_11685);
or U12264 (N_12264,N_11305,N_11392);
or U12265 (N_12265,N_11966,N_11666);
nand U12266 (N_12266,N_11840,N_11592);
nor U12267 (N_12267,N_11409,N_11363);
nor U12268 (N_12268,N_11385,N_11530);
xor U12269 (N_12269,N_11290,N_11611);
and U12270 (N_12270,N_11997,N_11927);
nor U12271 (N_12271,N_11574,N_11962);
and U12272 (N_12272,N_11940,N_11276);
nor U12273 (N_12273,N_11373,N_11523);
or U12274 (N_12274,N_11566,N_11735);
or U12275 (N_12275,N_11323,N_11382);
nand U12276 (N_12276,N_11521,N_11402);
nor U12277 (N_12277,N_11960,N_11422);
and U12278 (N_12278,N_11403,N_11309);
xor U12279 (N_12279,N_11292,N_11394);
or U12280 (N_12280,N_11800,N_11829);
or U12281 (N_12281,N_11793,N_11469);
or U12282 (N_12282,N_11439,N_11850);
xor U12283 (N_12283,N_11572,N_11555);
or U12284 (N_12284,N_11411,N_11517);
nor U12285 (N_12285,N_11399,N_11765);
or U12286 (N_12286,N_11876,N_11769);
xor U12287 (N_12287,N_11304,N_11745);
and U12288 (N_12288,N_11401,N_11284);
xnor U12289 (N_12289,N_11865,N_11370);
and U12290 (N_12290,N_11862,N_11465);
nor U12291 (N_12291,N_11691,N_11420);
nand U12292 (N_12292,N_11595,N_11389);
nor U12293 (N_12293,N_11902,N_11972);
and U12294 (N_12294,N_11913,N_11784);
nand U12295 (N_12295,N_11258,N_11347);
nand U12296 (N_12296,N_11345,N_11492);
nor U12297 (N_12297,N_11854,N_11312);
and U12298 (N_12298,N_11307,N_11417);
nand U12299 (N_12299,N_11900,N_11600);
or U12300 (N_12300,N_11947,N_11473);
and U12301 (N_12301,N_11620,N_11294);
nand U12302 (N_12302,N_11958,N_11485);
and U12303 (N_12303,N_11272,N_11667);
nor U12304 (N_12304,N_11851,N_11805);
and U12305 (N_12305,N_11979,N_11513);
nand U12306 (N_12306,N_11867,N_11400);
nor U12307 (N_12307,N_11506,N_11971);
and U12308 (N_12308,N_11860,N_11683);
nand U12309 (N_12309,N_11797,N_11675);
and U12310 (N_12310,N_11696,N_11841);
nor U12311 (N_12311,N_11783,N_11301);
or U12312 (N_12312,N_11757,N_11538);
or U12313 (N_12313,N_11780,N_11599);
or U12314 (N_12314,N_11353,N_11726);
nand U12315 (N_12315,N_11376,N_11254);
nor U12316 (N_12316,N_11529,N_11575);
or U12317 (N_12317,N_11367,N_11669);
nand U12318 (N_12318,N_11512,N_11446);
and U12319 (N_12319,N_11413,N_11589);
nand U12320 (N_12320,N_11501,N_11698);
and U12321 (N_12321,N_11383,N_11250);
nor U12322 (N_12322,N_11493,N_11444);
and U12323 (N_12323,N_11700,N_11883);
xor U12324 (N_12324,N_11959,N_11772);
xor U12325 (N_12325,N_11789,N_11573);
nor U12326 (N_12326,N_11474,N_11656);
or U12327 (N_12327,N_11690,N_11466);
nand U12328 (N_12328,N_11859,N_11472);
nor U12329 (N_12329,N_11956,N_11878);
and U12330 (N_12330,N_11579,N_11672);
nand U12331 (N_12331,N_11545,N_11624);
nand U12332 (N_12332,N_11803,N_11291);
nand U12333 (N_12333,N_11642,N_11414);
nand U12334 (N_12334,N_11896,N_11562);
nor U12335 (N_12335,N_11368,N_11505);
nand U12336 (N_12336,N_11948,N_11901);
or U12337 (N_12337,N_11649,N_11916);
xor U12338 (N_12338,N_11836,N_11360);
nor U12339 (N_12339,N_11260,N_11832);
or U12340 (N_12340,N_11540,N_11585);
nand U12341 (N_12341,N_11933,N_11483);
xor U12342 (N_12342,N_11771,N_11737);
or U12343 (N_12343,N_11774,N_11920);
and U12344 (N_12344,N_11547,N_11821);
and U12345 (N_12345,N_11981,N_11433);
nor U12346 (N_12346,N_11458,N_11467);
or U12347 (N_12347,N_11942,N_11266);
nor U12348 (N_12348,N_11978,N_11334);
nor U12349 (N_12349,N_11602,N_11725);
xor U12350 (N_12350,N_11861,N_11715);
nor U12351 (N_12351,N_11695,N_11934);
and U12352 (N_12352,N_11480,N_11796);
and U12353 (N_12353,N_11539,N_11680);
nor U12354 (N_12354,N_11612,N_11456);
or U12355 (N_12355,N_11282,N_11746);
nor U12356 (N_12356,N_11722,N_11457);
or U12357 (N_12357,N_11907,N_11689);
or U12358 (N_12358,N_11621,N_11761);
xor U12359 (N_12359,N_11809,N_11351);
or U12360 (N_12360,N_11543,N_11697);
or U12361 (N_12361,N_11817,N_11905);
and U12362 (N_12362,N_11946,N_11655);
nand U12363 (N_12363,N_11908,N_11703);
and U12364 (N_12364,N_11604,N_11873);
and U12365 (N_12365,N_11329,N_11597);
nor U12366 (N_12366,N_11816,N_11464);
xnor U12367 (N_12367,N_11795,N_11869);
nand U12368 (N_12368,N_11657,N_11253);
or U12369 (N_12369,N_11362,N_11801);
xnor U12370 (N_12370,N_11694,N_11619);
or U12371 (N_12371,N_11742,N_11835);
nand U12372 (N_12372,N_11340,N_11754);
or U12373 (N_12373,N_11369,N_11634);
xor U12374 (N_12374,N_11711,N_11525);
nor U12375 (N_12375,N_11651,N_11568);
xor U12376 (N_12376,N_11302,N_11252);
nor U12377 (N_12377,N_11583,N_11557);
and U12378 (N_12378,N_11822,N_11785);
nor U12379 (N_12379,N_11468,N_11381);
nand U12380 (N_12380,N_11614,N_11843);
and U12381 (N_12381,N_11811,N_11276);
and U12382 (N_12382,N_11506,N_11437);
and U12383 (N_12383,N_11346,N_11330);
nand U12384 (N_12384,N_11642,N_11353);
nor U12385 (N_12385,N_11483,N_11914);
and U12386 (N_12386,N_11668,N_11344);
or U12387 (N_12387,N_11658,N_11488);
nor U12388 (N_12388,N_11350,N_11714);
and U12389 (N_12389,N_11694,N_11859);
and U12390 (N_12390,N_11633,N_11794);
nor U12391 (N_12391,N_11399,N_11622);
nand U12392 (N_12392,N_11921,N_11305);
or U12393 (N_12393,N_11900,N_11321);
or U12394 (N_12394,N_11404,N_11376);
nor U12395 (N_12395,N_11737,N_11363);
nand U12396 (N_12396,N_11337,N_11777);
xor U12397 (N_12397,N_11963,N_11508);
and U12398 (N_12398,N_11367,N_11857);
and U12399 (N_12399,N_11723,N_11821);
nand U12400 (N_12400,N_11919,N_11415);
and U12401 (N_12401,N_11330,N_11502);
and U12402 (N_12402,N_11981,N_11984);
nand U12403 (N_12403,N_11870,N_11828);
xor U12404 (N_12404,N_11565,N_11994);
nand U12405 (N_12405,N_11565,N_11828);
nand U12406 (N_12406,N_11692,N_11634);
nand U12407 (N_12407,N_11611,N_11969);
nor U12408 (N_12408,N_11927,N_11510);
or U12409 (N_12409,N_11664,N_11591);
and U12410 (N_12410,N_11850,N_11908);
and U12411 (N_12411,N_11374,N_11297);
or U12412 (N_12412,N_11608,N_11556);
or U12413 (N_12413,N_11512,N_11779);
or U12414 (N_12414,N_11716,N_11743);
or U12415 (N_12415,N_11300,N_11928);
nor U12416 (N_12416,N_11742,N_11848);
or U12417 (N_12417,N_11550,N_11453);
nand U12418 (N_12418,N_11618,N_11670);
nand U12419 (N_12419,N_11727,N_11664);
nor U12420 (N_12420,N_11256,N_11713);
nor U12421 (N_12421,N_11686,N_11969);
or U12422 (N_12422,N_11604,N_11582);
nor U12423 (N_12423,N_11778,N_11707);
and U12424 (N_12424,N_11297,N_11904);
or U12425 (N_12425,N_11826,N_11494);
nand U12426 (N_12426,N_11988,N_11256);
nand U12427 (N_12427,N_11849,N_11973);
nor U12428 (N_12428,N_11515,N_11419);
or U12429 (N_12429,N_11713,N_11865);
xor U12430 (N_12430,N_11696,N_11952);
nand U12431 (N_12431,N_11668,N_11722);
nand U12432 (N_12432,N_11548,N_11559);
or U12433 (N_12433,N_11970,N_11475);
nor U12434 (N_12434,N_11696,N_11637);
nor U12435 (N_12435,N_11329,N_11807);
and U12436 (N_12436,N_11919,N_11471);
and U12437 (N_12437,N_11904,N_11412);
and U12438 (N_12438,N_11250,N_11691);
nor U12439 (N_12439,N_11599,N_11999);
and U12440 (N_12440,N_11512,N_11483);
nor U12441 (N_12441,N_11861,N_11900);
and U12442 (N_12442,N_11821,N_11359);
nor U12443 (N_12443,N_11338,N_11803);
nand U12444 (N_12444,N_11591,N_11447);
or U12445 (N_12445,N_11453,N_11622);
nor U12446 (N_12446,N_11558,N_11644);
nor U12447 (N_12447,N_11340,N_11409);
and U12448 (N_12448,N_11391,N_11279);
nor U12449 (N_12449,N_11612,N_11273);
and U12450 (N_12450,N_11260,N_11771);
nor U12451 (N_12451,N_11635,N_11261);
and U12452 (N_12452,N_11590,N_11654);
nor U12453 (N_12453,N_11639,N_11941);
or U12454 (N_12454,N_11451,N_11378);
nand U12455 (N_12455,N_11895,N_11809);
nor U12456 (N_12456,N_11524,N_11664);
xnor U12457 (N_12457,N_11782,N_11835);
xor U12458 (N_12458,N_11847,N_11477);
nand U12459 (N_12459,N_11715,N_11651);
and U12460 (N_12460,N_11760,N_11664);
and U12461 (N_12461,N_11446,N_11893);
or U12462 (N_12462,N_11974,N_11555);
and U12463 (N_12463,N_11252,N_11329);
nand U12464 (N_12464,N_11386,N_11482);
or U12465 (N_12465,N_11701,N_11772);
or U12466 (N_12466,N_11741,N_11864);
nor U12467 (N_12467,N_11692,N_11734);
and U12468 (N_12468,N_11582,N_11800);
and U12469 (N_12469,N_11518,N_11378);
or U12470 (N_12470,N_11343,N_11282);
or U12471 (N_12471,N_11748,N_11287);
or U12472 (N_12472,N_11991,N_11987);
xnor U12473 (N_12473,N_11989,N_11584);
and U12474 (N_12474,N_11599,N_11364);
and U12475 (N_12475,N_11484,N_11886);
nand U12476 (N_12476,N_11964,N_11699);
or U12477 (N_12477,N_11951,N_11524);
and U12478 (N_12478,N_11783,N_11429);
nor U12479 (N_12479,N_11437,N_11617);
and U12480 (N_12480,N_11935,N_11369);
nor U12481 (N_12481,N_11737,N_11654);
or U12482 (N_12482,N_11365,N_11587);
or U12483 (N_12483,N_11716,N_11516);
and U12484 (N_12484,N_11861,N_11965);
nand U12485 (N_12485,N_11550,N_11317);
nor U12486 (N_12486,N_11383,N_11632);
nand U12487 (N_12487,N_11568,N_11321);
and U12488 (N_12488,N_11637,N_11440);
or U12489 (N_12489,N_11953,N_11804);
nand U12490 (N_12490,N_11513,N_11546);
xnor U12491 (N_12491,N_11873,N_11911);
nor U12492 (N_12492,N_11815,N_11622);
or U12493 (N_12493,N_11447,N_11475);
nand U12494 (N_12494,N_11874,N_11529);
xnor U12495 (N_12495,N_11332,N_11745);
xnor U12496 (N_12496,N_11404,N_11553);
nor U12497 (N_12497,N_11870,N_11941);
or U12498 (N_12498,N_11508,N_11726);
nor U12499 (N_12499,N_11256,N_11330);
or U12500 (N_12500,N_11633,N_11250);
and U12501 (N_12501,N_11780,N_11758);
and U12502 (N_12502,N_11322,N_11308);
nand U12503 (N_12503,N_11661,N_11460);
nand U12504 (N_12504,N_11917,N_11521);
nand U12505 (N_12505,N_11400,N_11985);
or U12506 (N_12506,N_11456,N_11993);
or U12507 (N_12507,N_11771,N_11691);
nor U12508 (N_12508,N_11957,N_11667);
nor U12509 (N_12509,N_11835,N_11501);
and U12510 (N_12510,N_11612,N_11301);
nand U12511 (N_12511,N_11484,N_11260);
nor U12512 (N_12512,N_11491,N_11483);
xor U12513 (N_12513,N_11537,N_11922);
and U12514 (N_12514,N_11501,N_11772);
nor U12515 (N_12515,N_11828,N_11844);
or U12516 (N_12516,N_11751,N_11556);
and U12517 (N_12517,N_11879,N_11361);
nand U12518 (N_12518,N_11748,N_11455);
nand U12519 (N_12519,N_11399,N_11950);
nor U12520 (N_12520,N_11741,N_11527);
nand U12521 (N_12521,N_11751,N_11395);
or U12522 (N_12522,N_11425,N_11511);
nand U12523 (N_12523,N_11762,N_11519);
nand U12524 (N_12524,N_11751,N_11433);
nand U12525 (N_12525,N_11742,N_11259);
nand U12526 (N_12526,N_11647,N_11435);
or U12527 (N_12527,N_11554,N_11947);
xnor U12528 (N_12528,N_11994,N_11336);
xor U12529 (N_12529,N_11813,N_11814);
and U12530 (N_12530,N_11928,N_11499);
xor U12531 (N_12531,N_11520,N_11662);
nand U12532 (N_12532,N_11812,N_11823);
nor U12533 (N_12533,N_11927,N_11657);
nand U12534 (N_12534,N_11912,N_11477);
nand U12535 (N_12535,N_11941,N_11300);
or U12536 (N_12536,N_11736,N_11795);
nor U12537 (N_12537,N_11402,N_11868);
or U12538 (N_12538,N_11681,N_11408);
and U12539 (N_12539,N_11667,N_11328);
nand U12540 (N_12540,N_11559,N_11444);
xor U12541 (N_12541,N_11848,N_11871);
xor U12542 (N_12542,N_11904,N_11349);
and U12543 (N_12543,N_11286,N_11332);
and U12544 (N_12544,N_11740,N_11343);
and U12545 (N_12545,N_11503,N_11533);
xor U12546 (N_12546,N_11763,N_11516);
nor U12547 (N_12547,N_11778,N_11361);
nor U12548 (N_12548,N_11543,N_11901);
or U12549 (N_12549,N_11537,N_11908);
or U12550 (N_12550,N_11396,N_11500);
xnor U12551 (N_12551,N_11565,N_11548);
nor U12552 (N_12552,N_11917,N_11555);
nand U12553 (N_12553,N_11808,N_11611);
nor U12554 (N_12554,N_11848,N_11492);
xnor U12555 (N_12555,N_11653,N_11289);
or U12556 (N_12556,N_11332,N_11673);
and U12557 (N_12557,N_11254,N_11636);
nor U12558 (N_12558,N_11930,N_11600);
nor U12559 (N_12559,N_11522,N_11677);
nor U12560 (N_12560,N_11764,N_11862);
and U12561 (N_12561,N_11957,N_11345);
and U12562 (N_12562,N_11639,N_11935);
and U12563 (N_12563,N_11801,N_11827);
and U12564 (N_12564,N_11927,N_11595);
and U12565 (N_12565,N_11652,N_11955);
nand U12566 (N_12566,N_11572,N_11435);
nand U12567 (N_12567,N_11798,N_11569);
or U12568 (N_12568,N_11257,N_11907);
and U12569 (N_12569,N_11507,N_11673);
nand U12570 (N_12570,N_11566,N_11398);
nor U12571 (N_12571,N_11357,N_11782);
and U12572 (N_12572,N_11597,N_11836);
or U12573 (N_12573,N_11741,N_11615);
and U12574 (N_12574,N_11733,N_11269);
nand U12575 (N_12575,N_11528,N_11541);
nor U12576 (N_12576,N_11806,N_11956);
nor U12577 (N_12577,N_11796,N_11639);
nand U12578 (N_12578,N_11895,N_11270);
nor U12579 (N_12579,N_11637,N_11689);
and U12580 (N_12580,N_11653,N_11650);
and U12581 (N_12581,N_11545,N_11456);
and U12582 (N_12582,N_11419,N_11438);
nor U12583 (N_12583,N_11438,N_11591);
nand U12584 (N_12584,N_11438,N_11587);
and U12585 (N_12585,N_11488,N_11746);
and U12586 (N_12586,N_11915,N_11695);
or U12587 (N_12587,N_11858,N_11755);
xnor U12588 (N_12588,N_11792,N_11618);
nor U12589 (N_12589,N_11463,N_11992);
nor U12590 (N_12590,N_11980,N_11595);
or U12591 (N_12591,N_11698,N_11686);
xor U12592 (N_12592,N_11861,N_11393);
or U12593 (N_12593,N_11433,N_11736);
xnor U12594 (N_12594,N_11484,N_11544);
nand U12595 (N_12595,N_11255,N_11683);
or U12596 (N_12596,N_11250,N_11833);
nor U12597 (N_12597,N_11334,N_11900);
nor U12598 (N_12598,N_11444,N_11446);
or U12599 (N_12599,N_11840,N_11506);
nand U12600 (N_12600,N_11579,N_11875);
or U12601 (N_12601,N_11276,N_11930);
nor U12602 (N_12602,N_11531,N_11944);
nor U12603 (N_12603,N_11841,N_11264);
nand U12604 (N_12604,N_11368,N_11710);
nor U12605 (N_12605,N_11561,N_11474);
xnor U12606 (N_12606,N_11766,N_11914);
and U12607 (N_12607,N_11876,N_11380);
and U12608 (N_12608,N_11972,N_11564);
and U12609 (N_12609,N_11690,N_11768);
and U12610 (N_12610,N_11640,N_11930);
and U12611 (N_12611,N_11878,N_11515);
and U12612 (N_12612,N_11949,N_11989);
nor U12613 (N_12613,N_11986,N_11727);
xnor U12614 (N_12614,N_11541,N_11567);
nor U12615 (N_12615,N_11689,N_11896);
or U12616 (N_12616,N_11661,N_11816);
nor U12617 (N_12617,N_11342,N_11744);
and U12618 (N_12618,N_11488,N_11786);
or U12619 (N_12619,N_11333,N_11917);
or U12620 (N_12620,N_11853,N_11729);
and U12621 (N_12621,N_11757,N_11713);
or U12622 (N_12622,N_11836,N_11270);
nand U12623 (N_12623,N_11435,N_11770);
or U12624 (N_12624,N_11704,N_11899);
nor U12625 (N_12625,N_11935,N_11418);
or U12626 (N_12626,N_11321,N_11869);
and U12627 (N_12627,N_11655,N_11679);
nand U12628 (N_12628,N_11778,N_11262);
and U12629 (N_12629,N_11329,N_11581);
xnor U12630 (N_12630,N_11733,N_11522);
nand U12631 (N_12631,N_11960,N_11646);
nand U12632 (N_12632,N_11872,N_11893);
or U12633 (N_12633,N_11481,N_11504);
nand U12634 (N_12634,N_11386,N_11511);
or U12635 (N_12635,N_11515,N_11292);
or U12636 (N_12636,N_11900,N_11302);
or U12637 (N_12637,N_11562,N_11942);
and U12638 (N_12638,N_11747,N_11636);
or U12639 (N_12639,N_11372,N_11510);
or U12640 (N_12640,N_11674,N_11949);
or U12641 (N_12641,N_11807,N_11623);
xnor U12642 (N_12642,N_11941,N_11840);
xnor U12643 (N_12643,N_11666,N_11522);
xor U12644 (N_12644,N_11267,N_11619);
and U12645 (N_12645,N_11473,N_11446);
or U12646 (N_12646,N_11781,N_11622);
or U12647 (N_12647,N_11473,N_11255);
xor U12648 (N_12648,N_11300,N_11791);
nand U12649 (N_12649,N_11398,N_11866);
or U12650 (N_12650,N_11876,N_11967);
nor U12651 (N_12651,N_11844,N_11314);
or U12652 (N_12652,N_11880,N_11331);
or U12653 (N_12653,N_11831,N_11322);
or U12654 (N_12654,N_11651,N_11279);
nand U12655 (N_12655,N_11819,N_11802);
nor U12656 (N_12656,N_11276,N_11981);
nand U12657 (N_12657,N_11368,N_11609);
xnor U12658 (N_12658,N_11443,N_11871);
nor U12659 (N_12659,N_11876,N_11358);
and U12660 (N_12660,N_11769,N_11825);
or U12661 (N_12661,N_11376,N_11487);
or U12662 (N_12662,N_11480,N_11723);
xnor U12663 (N_12663,N_11897,N_11676);
nand U12664 (N_12664,N_11732,N_11345);
nor U12665 (N_12665,N_11586,N_11503);
nand U12666 (N_12666,N_11756,N_11642);
nor U12667 (N_12667,N_11646,N_11363);
or U12668 (N_12668,N_11735,N_11831);
or U12669 (N_12669,N_11656,N_11374);
nand U12670 (N_12670,N_11355,N_11399);
nor U12671 (N_12671,N_11828,N_11265);
nor U12672 (N_12672,N_11569,N_11883);
nor U12673 (N_12673,N_11654,N_11527);
nand U12674 (N_12674,N_11261,N_11996);
xnor U12675 (N_12675,N_11371,N_11476);
or U12676 (N_12676,N_11448,N_11273);
nor U12677 (N_12677,N_11398,N_11281);
or U12678 (N_12678,N_11785,N_11669);
nand U12679 (N_12679,N_11286,N_11658);
and U12680 (N_12680,N_11390,N_11607);
or U12681 (N_12681,N_11625,N_11845);
or U12682 (N_12682,N_11872,N_11292);
nor U12683 (N_12683,N_11466,N_11679);
nand U12684 (N_12684,N_11593,N_11369);
and U12685 (N_12685,N_11850,N_11517);
or U12686 (N_12686,N_11958,N_11567);
or U12687 (N_12687,N_11428,N_11590);
nor U12688 (N_12688,N_11888,N_11663);
nor U12689 (N_12689,N_11746,N_11798);
or U12690 (N_12690,N_11727,N_11600);
nand U12691 (N_12691,N_11649,N_11360);
and U12692 (N_12692,N_11378,N_11313);
nor U12693 (N_12693,N_11511,N_11330);
xor U12694 (N_12694,N_11383,N_11847);
xnor U12695 (N_12695,N_11653,N_11279);
nand U12696 (N_12696,N_11972,N_11962);
nand U12697 (N_12697,N_11696,N_11800);
and U12698 (N_12698,N_11924,N_11277);
or U12699 (N_12699,N_11607,N_11646);
nand U12700 (N_12700,N_11459,N_11308);
nor U12701 (N_12701,N_11458,N_11417);
or U12702 (N_12702,N_11457,N_11569);
nand U12703 (N_12703,N_11931,N_11824);
or U12704 (N_12704,N_11657,N_11535);
or U12705 (N_12705,N_11869,N_11716);
nor U12706 (N_12706,N_11469,N_11955);
and U12707 (N_12707,N_11637,N_11429);
xnor U12708 (N_12708,N_11334,N_11463);
or U12709 (N_12709,N_11303,N_11962);
nand U12710 (N_12710,N_11407,N_11860);
and U12711 (N_12711,N_11694,N_11986);
or U12712 (N_12712,N_11863,N_11763);
nand U12713 (N_12713,N_11848,N_11346);
and U12714 (N_12714,N_11368,N_11293);
nand U12715 (N_12715,N_11565,N_11481);
or U12716 (N_12716,N_11859,N_11521);
and U12717 (N_12717,N_11326,N_11978);
or U12718 (N_12718,N_11658,N_11597);
nand U12719 (N_12719,N_11486,N_11470);
nor U12720 (N_12720,N_11708,N_11657);
xnor U12721 (N_12721,N_11297,N_11539);
or U12722 (N_12722,N_11997,N_11902);
or U12723 (N_12723,N_11296,N_11573);
nand U12724 (N_12724,N_11923,N_11407);
nor U12725 (N_12725,N_11259,N_11904);
nor U12726 (N_12726,N_11909,N_11815);
and U12727 (N_12727,N_11423,N_11346);
nor U12728 (N_12728,N_11263,N_11284);
nand U12729 (N_12729,N_11551,N_11455);
and U12730 (N_12730,N_11401,N_11385);
or U12731 (N_12731,N_11682,N_11572);
or U12732 (N_12732,N_11542,N_11777);
and U12733 (N_12733,N_11549,N_11461);
or U12734 (N_12734,N_11255,N_11388);
and U12735 (N_12735,N_11395,N_11552);
xor U12736 (N_12736,N_11720,N_11580);
nand U12737 (N_12737,N_11398,N_11261);
xor U12738 (N_12738,N_11467,N_11831);
or U12739 (N_12739,N_11823,N_11650);
or U12740 (N_12740,N_11666,N_11406);
or U12741 (N_12741,N_11862,N_11714);
or U12742 (N_12742,N_11935,N_11890);
or U12743 (N_12743,N_11723,N_11815);
nand U12744 (N_12744,N_11883,N_11751);
nand U12745 (N_12745,N_11756,N_11565);
and U12746 (N_12746,N_11953,N_11960);
nor U12747 (N_12747,N_11291,N_11382);
nor U12748 (N_12748,N_11794,N_11922);
or U12749 (N_12749,N_11601,N_11423);
and U12750 (N_12750,N_12239,N_12344);
nor U12751 (N_12751,N_12224,N_12582);
xor U12752 (N_12752,N_12167,N_12022);
and U12753 (N_12753,N_12090,N_12185);
nor U12754 (N_12754,N_12035,N_12730);
nor U12755 (N_12755,N_12371,N_12101);
nand U12756 (N_12756,N_12277,N_12365);
or U12757 (N_12757,N_12233,N_12369);
nand U12758 (N_12758,N_12316,N_12472);
or U12759 (N_12759,N_12418,N_12123);
or U12760 (N_12760,N_12315,N_12205);
nor U12761 (N_12761,N_12640,N_12109);
nand U12762 (N_12762,N_12720,N_12478);
xor U12763 (N_12763,N_12197,N_12335);
and U12764 (N_12764,N_12641,N_12722);
or U12765 (N_12765,N_12531,N_12413);
and U12766 (N_12766,N_12324,N_12083);
nor U12767 (N_12767,N_12415,N_12565);
or U12768 (N_12768,N_12716,N_12334);
and U12769 (N_12769,N_12406,N_12164);
or U12770 (N_12770,N_12595,N_12557);
xor U12771 (N_12771,N_12085,N_12046);
nor U12772 (N_12772,N_12590,N_12102);
xnor U12773 (N_12773,N_12068,N_12520);
nand U12774 (N_12774,N_12354,N_12744);
xor U12775 (N_12775,N_12516,N_12537);
nor U12776 (N_12776,N_12691,N_12096);
and U12777 (N_12777,N_12281,N_12455);
and U12778 (N_12778,N_12223,N_12417);
nand U12779 (N_12779,N_12412,N_12597);
nor U12780 (N_12780,N_12631,N_12392);
nand U12781 (N_12781,N_12280,N_12298);
xnor U12782 (N_12782,N_12091,N_12303);
or U12783 (N_12783,N_12092,N_12456);
or U12784 (N_12784,N_12144,N_12048);
and U12785 (N_12785,N_12162,N_12591);
and U12786 (N_12786,N_12683,N_12705);
nor U12787 (N_12787,N_12555,N_12302);
nor U12788 (N_12788,N_12188,N_12178);
or U12789 (N_12789,N_12718,N_12559);
and U12790 (N_12790,N_12570,N_12427);
nor U12791 (N_12791,N_12607,N_12206);
nor U12792 (N_12792,N_12491,N_12146);
nor U12793 (N_12793,N_12604,N_12440);
nor U12794 (N_12794,N_12363,N_12558);
or U12795 (N_12795,N_12657,N_12171);
nor U12796 (N_12796,N_12402,N_12645);
nand U12797 (N_12797,N_12739,N_12275);
nor U12798 (N_12798,N_12485,N_12130);
nor U12799 (N_12799,N_12470,N_12457);
and U12800 (N_12800,N_12002,N_12122);
nor U12801 (N_12801,N_12195,N_12287);
nand U12802 (N_12802,N_12309,N_12284);
and U12803 (N_12803,N_12421,N_12600);
and U12804 (N_12804,N_12056,N_12310);
nor U12805 (N_12805,N_12719,N_12329);
nor U12806 (N_12806,N_12232,N_12211);
xor U12807 (N_12807,N_12115,N_12154);
nor U12808 (N_12808,N_12124,N_12285);
or U12809 (N_12809,N_12743,N_12082);
or U12810 (N_12810,N_12707,N_12658);
or U12811 (N_12811,N_12611,N_12688);
and U12812 (N_12812,N_12395,N_12243);
nand U12813 (N_12813,N_12042,N_12337);
nand U12814 (N_12814,N_12050,N_12345);
nor U12815 (N_12815,N_12529,N_12038);
nor U12816 (N_12816,N_12080,N_12397);
nand U12817 (N_12817,N_12240,N_12332);
or U12818 (N_12818,N_12074,N_12136);
nand U12819 (N_12819,N_12069,N_12461);
nand U12820 (N_12820,N_12339,N_12450);
and U12821 (N_12821,N_12312,N_12493);
or U12822 (N_12822,N_12453,N_12499);
nor U12823 (N_12823,N_12501,N_12588);
or U12824 (N_12824,N_12256,N_12294);
nor U12825 (N_12825,N_12479,N_12387);
nand U12826 (N_12826,N_12218,N_12267);
or U12827 (N_12827,N_12677,N_12268);
nor U12828 (N_12828,N_12532,N_12086);
and U12829 (N_12829,N_12204,N_12250);
nor U12830 (N_12830,N_12401,N_12319);
and U12831 (N_12831,N_12653,N_12053);
nand U12832 (N_12832,N_12741,N_12140);
nand U12833 (N_12833,N_12432,N_12465);
and U12834 (N_12834,N_12051,N_12473);
nor U12835 (N_12835,N_12362,N_12674);
or U12836 (N_12836,N_12684,N_12749);
nor U12837 (N_12837,N_12576,N_12687);
or U12838 (N_12838,N_12668,N_12721);
nor U12839 (N_12839,N_12650,N_12638);
nand U12840 (N_12840,N_12325,N_12575);
or U12841 (N_12841,N_12694,N_12198);
or U12842 (N_12842,N_12405,N_12732);
or U12843 (N_12843,N_12617,N_12648);
and U12844 (N_12844,N_12601,N_12420);
or U12845 (N_12845,N_12540,N_12679);
nor U12846 (N_12846,N_12746,N_12106);
and U12847 (N_12847,N_12409,N_12437);
and U12848 (N_12848,N_12213,N_12297);
nor U12849 (N_12849,N_12574,N_12311);
xnor U12850 (N_12850,N_12610,N_12227);
xor U12851 (N_12851,N_12208,N_12646);
or U12852 (N_12852,N_12076,N_12643);
nand U12853 (N_12853,N_12020,N_12702);
and U12854 (N_12854,N_12681,N_12169);
or U12855 (N_12855,N_12567,N_12100);
or U12856 (N_12856,N_12360,N_12293);
nor U12857 (N_12857,N_12723,N_12709);
or U12858 (N_12858,N_12655,N_12221);
or U12859 (N_12859,N_12644,N_12623);
nand U12860 (N_12860,N_12554,N_12117);
nor U12861 (N_12861,N_12449,N_12375);
and U12862 (N_12862,N_12241,N_12141);
and U12863 (N_12863,N_12000,N_12699);
xor U12864 (N_12864,N_12636,N_12477);
and U12865 (N_12865,N_12138,N_12306);
or U12866 (N_12866,N_12353,N_12422);
xnor U12867 (N_12867,N_12466,N_12112);
or U12868 (N_12868,N_12403,N_12592);
or U12869 (N_12869,N_12127,N_12013);
and U12870 (N_12870,N_12536,N_12246);
and U12871 (N_12871,N_12075,N_12627);
and U12872 (N_12872,N_12220,N_12236);
or U12873 (N_12873,N_12613,N_12318);
nand U12874 (N_12874,N_12672,N_12553);
nor U12875 (N_12875,N_12632,N_12028);
or U12876 (N_12876,N_12252,N_12475);
xnor U12877 (N_12877,N_12662,N_12729);
nand U12878 (N_12878,N_12301,N_12033);
nand U12879 (N_12879,N_12669,N_12094);
nand U12880 (N_12880,N_12111,N_12549);
nor U12881 (N_12881,N_12724,N_12510);
or U12882 (N_12882,N_12304,N_12314);
or U12883 (N_12883,N_12242,N_12533);
and U12884 (N_12884,N_12216,N_12398);
nor U12885 (N_12885,N_12482,N_12159);
nand U12886 (N_12886,N_12016,N_12045);
xor U12887 (N_12887,N_12511,N_12125);
and U12888 (N_12888,N_12099,N_12010);
nand U12889 (N_12889,N_12098,N_12199);
or U12890 (N_12890,N_12270,N_12380);
or U12891 (N_12891,N_12384,N_12061);
and U12892 (N_12892,N_12580,N_12690);
nor U12893 (N_12893,N_12264,N_12528);
and U12894 (N_12894,N_12291,N_12522);
or U12895 (N_12895,N_12134,N_12464);
nand U12896 (N_12896,N_12391,N_12150);
and U12897 (N_12897,N_12589,N_12370);
or U12898 (N_12898,N_12468,N_12740);
nor U12899 (N_12899,N_12172,N_12110);
and U12900 (N_12900,N_12341,N_12659);
nand U12901 (N_12901,N_12368,N_12139);
nand U12902 (N_12902,N_12462,N_12546);
nand U12903 (N_12903,N_12490,N_12151);
nand U12904 (N_12904,N_12733,N_12584);
or U12905 (N_12905,N_12487,N_12713);
xor U12906 (N_12906,N_12416,N_12697);
nor U12907 (N_12907,N_12547,N_12411);
nor U12908 (N_12908,N_12067,N_12399);
and U12909 (N_12909,N_12609,N_12348);
and U12910 (N_12910,N_12346,N_12700);
and U12911 (N_12911,N_12651,N_12133);
nor U12912 (N_12912,N_12625,N_12147);
and U12913 (N_12913,N_12505,N_12003);
or U12914 (N_12914,N_12571,N_12006);
nand U12915 (N_12915,N_12748,N_12551);
nor U12916 (N_12916,N_12515,N_12063);
xor U12917 (N_12917,N_12299,N_12606);
nor U12918 (N_12918,N_12143,N_12378);
and U12919 (N_12919,N_12018,N_12121);
or U12920 (N_12920,N_12120,N_12433);
xnor U12921 (N_12921,N_12229,N_12326);
and U12922 (N_12922,N_12525,N_12231);
or U12923 (N_12923,N_12087,N_12542);
and U12924 (N_12924,N_12503,N_12193);
and U12925 (N_12925,N_12212,N_12269);
nand U12926 (N_12926,N_12666,N_12444);
nor U12927 (N_12927,N_12561,N_12447);
nor U12928 (N_12928,N_12261,N_12071);
and U12929 (N_12929,N_12262,N_12254);
nand U12930 (N_12930,N_12317,N_12030);
nor U12931 (N_12931,N_12633,N_12394);
nor U12932 (N_12932,N_12234,N_12322);
nor U12933 (N_12933,N_12031,N_12634);
nand U12934 (N_12934,N_12512,N_12430);
or U12935 (N_12935,N_12701,N_12620);
xnor U12936 (N_12936,N_12129,N_12273);
and U12937 (N_12937,N_12043,N_12116);
xnor U12938 (N_12938,N_12596,N_12355);
nand U12939 (N_12939,N_12237,N_12564);
nand U12940 (N_12940,N_12726,N_12614);
nor U12941 (N_12941,N_12352,N_12019);
and U12942 (N_12942,N_12215,N_12340);
or U12943 (N_12943,N_12157,N_12507);
or U12944 (N_12944,N_12283,N_12084);
or U12945 (N_12945,N_12563,N_12272);
or U12946 (N_12946,N_12118,N_12598);
or U12947 (N_12947,N_12331,N_12602);
and U12948 (N_12948,N_12095,N_12014);
nor U12949 (N_12949,N_12621,N_12710);
nand U12950 (N_12950,N_12599,N_12446);
and U12951 (N_12951,N_12217,N_12523);
xor U12952 (N_12952,N_12058,N_12693);
xor U12953 (N_12953,N_12255,N_12165);
and U12954 (N_12954,N_12431,N_12715);
nand U12955 (N_12955,N_12593,N_12073);
nor U12956 (N_12956,N_12343,N_12448);
and U12957 (N_12957,N_12060,N_12305);
or U12958 (N_12958,N_12728,N_12498);
and U12959 (N_12959,N_12029,N_12044);
nand U12960 (N_12960,N_12383,N_12374);
and U12961 (N_12961,N_12400,N_12163);
nand U12962 (N_12962,N_12426,N_12637);
xnor U12963 (N_12963,N_12481,N_12647);
nand U12964 (N_12964,N_12635,N_12671);
nor U12965 (N_12965,N_12410,N_12509);
and U12966 (N_12966,N_12530,N_12495);
and U12967 (N_12967,N_12615,N_12451);
nand U12968 (N_12968,N_12725,N_12434);
nand U12969 (N_12969,N_12731,N_12257);
and U12970 (N_12970,N_12153,N_12747);
nand U12971 (N_12971,N_12059,N_12054);
nand U12972 (N_12972,N_12200,N_12156);
or U12973 (N_12973,N_12489,N_12560);
nand U12974 (N_12974,N_12292,N_12351);
nor U12975 (N_12975,N_12605,N_12568);
xnor U12976 (N_12976,N_12696,N_12458);
and U12977 (N_12977,N_12113,N_12097);
nor U12978 (N_12978,N_12286,N_12454);
and U12979 (N_12979,N_12271,N_12488);
nor U12980 (N_12980,N_12572,N_12712);
or U12981 (N_12981,N_12504,N_12049);
nor U12982 (N_12982,N_12502,N_12093);
nor U12983 (N_12983,N_12078,N_12745);
nand U12984 (N_12984,N_12618,N_12191);
and U12985 (N_12985,N_12196,N_12214);
and U12986 (N_12986,N_12258,N_12581);
nand U12987 (N_12987,N_12289,N_12333);
and U12988 (N_12988,N_12288,N_12180);
or U12989 (N_12989,N_12308,N_12009);
nand U12990 (N_12990,N_12587,N_12727);
nand U12991 (N_12991,N_12586,N_12145);
and U12992 (N_12992,N_12266,N_12443);
and U12993 (N_12993,N_12541,N_12535);
nor U12994 (N_12994,N_12170,N_12321);
nand U12995 (N_12995,N_12296,N_12320);
nand U12996 (N_12996,N_12245,N_12550);
or U12997 (N_12997,N_12577,N_12356);
xnor U12998 (N_12998,N_12072,N_12459);
and U12999 (N_12999,N_12717,N_12077);
nor U13000 (N_13000,N_12004,N_12137);
nor U13001 (N_13001,N_12247,N_12419);
nor U13002 (N_13002,N_12692,N_12460);
or U13003 (N_13003,N_12037,N_12177);
nor U13004 (N_13004,N_12492,N_12698);
or U13005 (N_13005,N_12055,N_12131);
and U13006 (N_13006,N_12181,N_12182);
nor U13007 (N_13007,N_12506,N_12665);
nor U13008 (N_13008,N_12689,N_12279);
nand U13009 (N_13009,N_12678,N_12439);
and U13010 (N_13010,N_12471,N_12396);
and U13011 (N_13011,N_12079,N_12148);
or U13012 (N_13012,N_12210,N_12508);
nand U13013 (N_13013,N_12630,N_12361);
nor U13014 (N_13014,N_12088,N_12379);
nand U13015 (N_13015,N_12128,N_12235);
or U13016 (N_13016,N_12738,N_12104);
xor U13017 (N_13017,N_12414,N_12480);
and U13018 (N_13018,N_12367,N_12173);
and U13019 (N_13019,N_12047,N_12336);
or U13020 (N_13020,N_12442,N_12359);
nor U13021 (N_13021,N_12377,N_12408);
or U13022 (N_13022,N_12518,N_12189);
or U13023 (N_13023,N_12347,N_12486);
and U13024 (N_13024,N_12389,N_12500);
nor U13025 (N_13025,N_12323,N_12132);
nor U13026 (N_13026,N_12583,N_12675);
or U13027 (N_13027,N_12024,N_12021);
nand U13028 (N_13028,N_12190,N_12194);
nand U13029 (N_13029,N_12695,N_12328);
nor U13030 (N_13030,N_12661,N_12249);
nor U13031 (N_13031,N_12062,N_12494);
nor U13032 (N_13032,N_12142,N_12742);
or U13033 (N_13033,N_12158,N_12517);
xnor U13034 (N_13034,N_12441,N_12603);
nand U13035 (N_13035,N_12276,N_12081);
xor U13036 (N_13036,N_12174,N_12032);
nand U13037 (N_13037,N_12160,N_12263);
nand U13038 (N_13038,N_12552,N_12386);
nor U13039 (N_13039,N_12007,N_12027);
nor U13040 (N_13040,N_12089,N_12187);
nor U13041 (N_13041,N_12103,N_12569);
xnor U13042 (N_13042,N_12736,N_12483);
or U13043 (N_13043,N_12436,N_12544);
nor U13044 (N_13044,N_12274,N_12070);
nor U13045 (N_13045,N_12040,N_12497);
or U13046 (N_13046,N_12654,N_12226);
xor U13047 (N_13047,N_12149,N_12545);
xnor U13048 (N_13048,N_12382,N_12251);
nor U13049 (N_13049,N_12682,N_12735);
nor U13050 (N_13050,N_12023,N_12425);
nor U13051 (N_13051,N_12521,N_12342);
nand U13052 (N_13052,N_12708,N_12057);
and U13053 (N_13053,N_12704,N_12628);
nor U13054 (N_13054,N_12225,N_12358);
or U13055 (N_13055,N_12642,N_12660);
or U13056 (N_13056,N_12649,N_12585);
nor U13057 (N_13057,N_12667,N_12543);
nand U13058 (N_13058,N_12155,N_12676);
nand U13059 (N_13059,N_12166,N_12179);
nand U13060 (N_13060,N_12664,N_12652);
xor U13061 (N_13061,N_12001,N_12015);
nor U13062 (N_13062,N_12126,N_12686);
xor U13063 (N_13063,N_12626,N_12680);
or U13064 (N_13064,N_12017,N_12519);
nand U13065 (N_13065,N_12364,N_12108);
nand U13066 (N_13066,N_12376,N_12207);
nor U13067 (N_13067,N_12608,N_12012);
and U13068 (N_13068,N_12105,N_12244);
or U13069 (N_13069,N_12639,N_12295);
or U13070 (N_13070,N_12573,N_12209);
or U13071 (N_13071,N_12228,N_12373);
or U13072 (N_13072,N_12248,N_12734);
nor U13073 (N_13073,N_12670,N_12467);
xor U13074 (N_13074,N_12527,N_12429);
xor U13075 (N_13075,N_12579,N_12330);
nand U13076 (N_13076,N_12039,N_12428);
nand U13077 (N_13077,N_12036,N_12496);
nand U13078 (N_13078,N_12578,N_12052);
nand U13079 (N_13079,N_12366,N_12445);
nand U13080 (N_13080,N_12175,N_12556);
nor U13081 (N_13081,N_12168,N_12152);
nor U13082 (N_13082,N_12183,N_12463);
and U13083 (N_13083,N_12025,N_12706);
nand U13084 (N_13084,N_12260,N_12407);
and U13085 (N_13085,N_12278,N_12259);
nor U13086 (N_13086,N_12476,N_12385);
nor U13087 (N_13087,N_12622,N_12566);
or U13088 (N_13088,N_12685,N_12065);
nand U13089 (N_13089,N_12524,N_12612);
nand U13090 (N_13090,N_12107,N_12135);
xnor U13091 (N_13091,N_12011,N_12381);
nand U13092 (N_13092,N_12265,N_12526);
xor U13093 (N_13093,N_12404,N_12539);
nor U13094 (N_13094,N_12202,N_12041);
or U13095 (N_13095,N_12338,N_12350);
xor U13096 (N_13096,N_12327,N_12624);
or U13097 (N_13097,N_12176,N_12184);
and U13098 (N_13098,N_12538,N_12238);
or U13099 (N_13099,N_12562,N_12663);
nand U13100 (N_13100,N_12514,N_12066);
nor U13101 (N_13101,N_12219,N_12034);
and U13102 (N_13102,N_12290,N_12119);
xnor U13103 (N_13103,N_12703,N_12513);
or U13104 (N_13104,N_12656,N_12372);
and U13105 (N_13105,N_12619,N_12673);
xnor U13106 (N_13106,N_12307,N_12064);
and U13107 (N_13107,N_12357,N_12253);
nand U13108 (N_13108,N_12192,N_12737);
and U13109 (N_13109,N_12201,N_12438);
or U13110 (N_13110,N_12313,N_12008);
or U13111 (N_13111,N_12393,N_12594);
nor U13112 (N_13112,N_12203,N_12714);
nand U13113 (N_13113,N_12423,N_12452);
xor U13114 (N_13114,N_12026,N_12469);
nand U13115 (N_13115,N_12230,N_12629);
or U13116 (N_13116,N_12114,N_12186);
nand U13117 (N_13117,N_12005,N_12161);
nor U13118 (N_13118,N_12300,N_12711);
nor U13119 (N_13119,N_12222,N_12424);
or U13120 (N_13120,N_12534,N_12484);
and U13121 (N_13121,N_12390,N_12616);
nor U13122 (N_13122,N_12349,N_12282);
nor U13123 (N_13123,N_12474,N_12435);
or U13124 (N_13124,N_12388,N_12548);
nor U13125 (N_13125,N_12471,N_12459);
and U13126 (N_13126,N_12058,N_12591);
nor U13127 (N_13127,N_12743,N_12605);
nand U13128 (N_13128,N_12706,N_12405);
or U13129 (N_13129,N_12461,N_12417);
nand U13130 (N_13130,N_12126,N_12009);
xnor U13131 (N_13131,N_12359,N_12084);
or U13132 (N_13132,N_12739,N_12142);
and U13133 (N_13133,N_12065,N_12381);
nand U13134 (N_13134,N_12711,N_12221);
xnor U13135 (N_13135,N_12421,N_12695);
nor U13136 (N_13136,N_12131,N_12318);
nor U13137 (N_13137,N_12443,N_12016);
nand U13138 (N_13138,N_12748,N_12044);
and U13139 (N_13139,N_12504,N_12102);
nand U13140 (N_13140,N_12397,N_12029);
and U13141 (N_13141,N_12683,N_12265);
nor U13142 (N_13142,N_12010,N_12014);
nor U13143 (N_13143,N_12417,N_12335);
nor U13144 (N_13144,N_12027,N_12509);
or U13145 (N_13145,N_12447,N_12148);
and U13146 (N_13146,N_12548,N_12509);
nor U13147 (N_13147,N_12357,N_12664);
and U13148 (N_13148,N_12087,N_12563);
or U13149 (N_13149,N_12232,N_12250);
nand U13150 (N_13150,N_12495,N_12453);
and U13151 (N_13151,N_12087,N_12493);
or U13152 (N_13152,N_12565,N_12026);
nand U13153 (N_13153,N_12348,N_12095);
nand U13154 (N_13154,N_12585,N_12463);
or U13155 (N_13155,N_12641,N_12490);
nor U13156 (N_13156,N_12353,N_12357);
or U13157 (N_13157,N_12368,N_12044);
or U13158 (N_13158,N_12745,N_12276);
nand U13159 (N_13159,N_12665,N_12447);
nand U13160 (N_13160,N_12498,N_12590);
xnor U13161 (N_13161,N_12076,N_12303);
nand U13162 (N_13162,N_12248,N_12091);
and U13163 (N_13163,N_12445,N_12022);
nor U13164 (N_13164,N_12061,N_12614);
and U13165 (N_13165,N_12003,N_12170);
and U13166 (N_13166,N_12505,N_12085);
nor U13167 (N_13167,N_12339,N_12099);
nand U13168 (N_13168,N_12489,N_12593);
or U13169 (N_13169,N_12555,N_12132);
or U13170 (N_13170,N_12328,N_12210);
nor U13171 (N_13171,N_12604,N_12611);
xor U13172 (N_13172,N_12583,N_12357);
nand U13173 (N_13173,N_12127,N_12038);
nand U13174 (N_13174,N_12342,N_12663);
or U13175 (N_13175,N_12524,N_12271);
nand U13176 (N_13176,N_12663,N_12115);
and U13177 (N_13177,N_12341,N_12239);
nor U13178 (N_13178,N_12720,N_12652);
nand U13179 (N_13179,N_12261,N_12619);
nor U13180 (N_13180,N_12649,N_12693);
nor U13181 (N_13181,N_12645,N_12138);
nand U13182 (N_13182,N_12023,N_12147);
or U13183 (N_13183,N_12215,N_12162);
nand U13184 (N_13184,N_12672,N_12132);
xor U13185 (N_13185,N_12623,N_12621);
nand U13186 (N_13186,N_12355,N_12212);
nor U13187 (N_13187,N_12737,N_12065);
and U13188 (N_13188,N_12074,N_12290);
nor U13189 (N_13189,N_12673,N_12736);
or U13190 (N_13190,N_12468,N_12420);
or U13191 (N_13191,N_12136,N_12540);
or U13192 (N_13192,N_12398,N_12314);
xnor U13193 (N_13193,N_12450,N_12128);
or U13194 (N_13194,N_12351,N_12727);
and U13195 (N_13195,N_12030,N_12722);
or U13196 (N_13196,N_12391,N_12322);
nand U13197 (N_13197,N_12286,N_12005);
and U13198 (N_13198,N_12463,N_12270);
or U13199 (N_13199,N_12572,N_12493);
xor U13200 (N_13200,N_12041,N_12050);
nand U13201 (N_13201,N_12349,N_12665);
or U13202 (N_13202,N_12596,N_12231);
nor U13203 (N_13203,N_12038,N_12434);
nor U13204 (N_13204,N_12152,N_12687);
nor U13205 (N_13205,N_12157,N_12713);
nand U13206 (N_13206,N_12029,N_12716);
and U13207 (N_13207,N_12151,N_12223);
or U13208 (N_13208,N_12485,N_12507);
nand U13209 (N_13209,N_12120,N_12344);
nor U13210 (N_13210,N_12704,N_12545);
or U13211 (N_13211,N_12189,N_12678);
nor U13212 (N_13212,N_12032,N_12186);
or U13213 (N_13213,N_12491,N_12131);
xor U13214 (N_13214,N_12250,N_12277);
xor U13215 (N_13215,N_12062,N_12603);
or U13216 (N_13216,N_12011,N_12012);
nor U13217 (N_13217,N_12448,N_12540);
nor U13218 (N_13218,N_12191,N_12275);
nor U13219 (N_13219,N_12486,N_12642);
nand U13220 (N_13220,N_12535,N_12505);
nor U13221 (N_13221,N_12458,N_12065);
and U13222 (N_13222,N_12194,N_12183);
xor U13223 (N_13223,N_12157,N_12034);
nand U13224 (N_13224,N_12089,N_12656);
xor U13225 (N_13225,N_12401,N_12313);
or U13226 (N_13226,N_12035,N_12022);
nand U13227 (N_13227,N_12211,N_12194);
nor U13228 (N_13228,N_12331,N_12441);
and U13229 (N_13229,N_12521,N_12153);
nor U13230 (N_13230,N_12390,N_12247);
or U13231 (N_13231,N_12518,N_12020);
and U13232 (N_13232,N_12152,N_12401);
nor U13233 (N_13233,N_12483,N_12039);
or U13234 (N_13234,N_12686,N_12511);
nor U13235 (N_13235,N_12248,N_12076);
nand U13236 (N_13236,N_12257,N_12314);
xor U13237 (N_13237,N_12352,N_12220);
nand U13238 (N_13238,N_12087,N_12508);
nand U13239 (N_13239,N_12467,N_12128);
or U13240 (N_13240,N_12589,N_12056);
nand U13241 (N_13241,N_12710,N_12434);
and U13242 (N_13242,N_12742,N_12296);
or U13243 (N_13243,N_12476,N_12434);
or U13244 (N_13244,N_12531,N_12541);
nand U13245 (N_13245,N_12164,N_12675);
and U13246 (N_13246,N_12084,N_12342);
or U13247 (N_13247,N_12418,N_12370);
and U13248 (N_13248,N_12652,N_12743);
and U13249 (N_13249,N_12320,N_12027);
xnor U13250 (N_13250,N_12641,N_12201);
nor U13251 (N_13251,N_12568,N_12132);
and U13252 (N_13252,N_12179,N_12058);
nand U13253 (N_13253,N_12735,N_12012);
nand U13254 (N_13254,N_12413,N_12149);
or U13255 (N_13255,N_12709,N_12544);
and U13256 (N_13256,N_12049,N_12180);
and U13257 (N_13257,N_12040,N_12718);
and U13258 (N_13258,N_12592,N_12461);
or U13259 (N_13259,N_12551,N_12532);
or U13260 (N_13260,N_12679,N_12003);
nor U13261 (N_13261,N_12252,N_12025);
nor U13262 (N_13262,N_12411,N_12708);
nand U13263 (N_13263,N_12646,N_12059);
or U13264 (N_13264,N_12006,N_12159);
or U13265 (N_13265,N_12311,N_12528);
nand U13266 (N_13266,N_12053,N_12570);
nand U13267 (N_13267,N_12358,N_12672);
and U13268 (N_13268,N_12715,N_12642);
or U13269 (N_13269,N_12036,N_12431);
nand U13270 (N_13270,N_12227,N_12366);
nand U13271 (N_13271,N_12407,N_12136);
nor U13272 (N_13272,N_12157,N_12401);
and U13273 (N_13273,N_12345,N_12567);
or U13274 (N_13274,N_12235,N_12525);
nand U13275 (N_13275,N_12485,N_12497);
nand U13276 (N_13276,N_12738,N_12580);
nand U13277 (N_13277,N_12414,N_12520);
nor U13278 (N_13278,N_12174,N_12092);
nor U13279 (N_13279,N_12174,N_12441);
nand U13280 (N_13280,N_12384,N_12010);
and U13281 (N_13281,N_12517,N_12139);
and U13282 (N_13282,N_12067,N_12616);
or U13283 (N_13283,N_12600,N_12126);
and U13284 (N_13284,N_12397,N_12486);
and U13285 (N_13285,N_12295,N_12104);
and U13286 (N_13286,N_12327,N_12406);
and U13287 (N_13287,N_12408,N_12562);
or U13288 (N_13288,N_12331,N_12614);
nor U13289 (N_13289,N_12170,N_12029);
or U13290 (N_13290,N_12581,N_12686);
xor U13291 (N_13291,N_12412,N_12177);
nand U13292 (N_13292,N_12742,N_12427);
or U13293 (N_13293,N_12622,N_12376);
and U13294 (N_13294,N_12076,N_12467);
or U13295 (N_13295,N_12278,N_12672);
or U13296 (N_13296,N_12632,N_12276);
nand U13297 (N_13297,N_12194,N_12346);
nor U13298 (N_13298,N_12010,N_12180);
and U13299 (N_13299,N_12365,N_12608);
and U13300 (N_13300,N_12518,N_12335);
or U13301 (N_13301,N_12203,N_12207);
and U13302 (N_13302,N_12675,N_12133);
nand U13303 (N_13303,N_12479,N_12329);
nand U13304 (N_13304,N_12664,N_12068);
or U13305 (N_13305,N_12026,N_12589);
nor U13306 (N_13306,N_12274,N_12163);
nor U13307 (N_13307,N_12363,N_12408);
xnor U13308 (N_13308,N_12385,N_12083);
nor U13309 (N_13309,N_12642,N_12474);
nand U13310 (N_13310,N_12451,N_12557);
and U13311 (N_13311,N_12574,N_12163);
nor U13312 (N_13312,N_12112,N_12080);
or U13313 (N_13313,N_12229,N_12468);
nand U13314 (N_13314,N_12132,N_12541);
nor U13315 (N_13315,N_12255,N_12641);
or U13316 (N_13316,N_12340,N_12400);
nor U13317 (N_13317,N_12259,N_12497);
xor U13318 (N_13318,N_12153,N_12039);
nor U13319 (N_13319,N_12145,N_12376);
or U13320 (N_13320,N_12387,N_12634);
nand U13321 (N_13321,N_12311,N_12183);
and U13322 (N_13322,N_12318,N_12171);
nor U13323 (N_13323,N_12655,N_12091);
or U13324 (N_13324,N_12048,N_12704);
xnor U13325 (N_13325,N_12381,N_12006);
nand U13326 (N_13326,N_12387,N_12683);
nor U13327 (N_13327,N_12674,N_12001);
xnor U13328 (N_13328,N_12542,N_12167);
and U13329 (N_13329,N_12147,N_12524);
nor U13330 (N_13330,N_12172,N_12554);
nor U13331 (N_13331,N_12329,N_12560);
or U13332 (N_13332,N_12308,N_12289);
and U13333 (N_13333,N_12506,N_12003);
and U13334 (N_13334,N_12346,N_12218);
nand U13335 (N_13335,N_12218,N_12537);
and U13336 (N_13336,N_12202,N_12236);
nand U13337 (N_13337,N_12681,N_12272);
and U13338 (N_13338,N_12469,N_12543);
nor U13339 (N_13339,N_12359,N_12095);
and U13340 (N_13340,N_12306,N_12281);
and U13341 (N_13341,N_12147,N_12327);
or U13342 (N_13342,N_12122,N_12145);
nand U13343 (N_13343,N_12086,N_12198);
nor U13344 (N_13344,N_12628,N_12595);
or U13345 (N_13345,N_12255,N_12458);
and U13346 (N_13346,N_12286,N_12639);
nor U13347 (N_13347,N_12629,N_12713);
and U13348 (N_13348,N_12247,N_12730);
or U13349 (N_13349,N_12446,N_12212);
nand U13350 (N_13350,N_12700,N_12349);
nor U13351 (N_13351,N_12718,N_12266);
nor U13352 (N_13352,N_12165,N_12419);
nand U13353 (N_13353,N_12696,N_12348);
and U13354 (N_13354,N_12325,N_12405);
nand U13355 (N_13355,N_12600,N_12405);
or U13356 (N_13356,N_12455,N_12342);
nor U13357 (N_13357,N_12253,N_12604);
and U13358 (N_13358,N_12201,N_12580);
nor U13359 (N_13359,N_12387,N_12116);
and U13360 (N_13360,N_12329,N_12111);
or U13361 (N_13361,N_12050,N_12427);
and U13362 (N_13362,N_12549,N_12391);
or U13363 (N_13363,N_12732,N_12336);
or U13364 (N_13364,N_12259,N_12307);
nand U13365 (N_13365,N_12433,N_12254);
or U13366 (N_13366,N_12300,N_12270);
and U13367 (N_13367,N_12466,N_12694);
nand U13368 (N_13368,N_12670,N_12667);
xnor U13369 (N_13369,N_12375,N_12237);
nor U13370 (N_13370,N_12744,N_12429);
nand U13371 (N_13371,N_12651,N_12737);
or U13372 (N_13372,N_12659,N_12407);
and U13373 (N_13373,N_12189,N_12351);
nand U13374 (N_13374,N_12549,N_12510);
and U13375 (N_13375,N_12277,N_12087);
or U13376 (N_13376,N_12704,N_12505);
nand U13377 (N_13377,N_12414,N_12483);
and U13378 (N_13378,N_12041,N_12419);
nor U13379 (N_13379,N_12329,N_12581);
or U13380 (N_13380,N_12400,N_12058);
nand U13381 (N_13381,N_12002,N_12703);
and U13382 (N_13382,N_12012,N_12357);
and U13383 (N_13383,N_12076,N_12402);
nor U13384 (N_13384,N_12670,N_12242);
and U13385 (N_13385,N_12529,N_12149);
xor U13386 (N_13386,N_12127,N_12494);
nand U13387 (N_13387,N_12507,N_12668);
nand U13388 (N_13388,N_12114,N_12523);
nand U13389 (N_13389,N_12259,N_12145);
nand U13390 (N_13390,N_12558,N_12022);
or U13391 (N_13391,N_12260,N_12513);
xnor U13392 (N_13392,N_12291,N_12603);
xor U13393 (N_13393,N_12556,N_12621);
nor U13394 (N_13394,N_12070,N_12535);
or U13395 (N_13395,N_12732,N_12537);
nor U13396 (N_13396,N_12694,N_12016);
nor U13397 (N_13397,N_12073,N_12605);
and U13398 (N_13398,N_12568,N_12626);
nor U13399 (N_13399,N_12318,N_12493);
nor U13400 (N_13400,N_12385,N_12600);
or U13401 (N_13401,N_12239,N_12444);
nand U13402 (N_13402,N_12169,N_12658);
and U13403 (N_13403,N_12607,N_12588);
xor U13404 (N_13404,N_12518,N_12346);
nor U13405 (N_13405,N_12534,N_12439);
and U13406 (N_13406,N_12606,N_12380);
or U13407 (N_13407,N_12264,N_12349);
nand U13408 (N_13408,N_12708,N_12046);
and U13409 (N_13409,N_12512,N_12006);
and U13410 (N_13410,N_12256,N_12255);
or U13411 (N_13411,N_12211,N_12538);
and U13412 (N_13412,N_12591,N_12148);
nand U13413 (N_13413,N_12033,N_12128);
nor U13414 (N_13414,N_12261,N_12454);
nor U13415 (N_13415,N_12394,N_12072);
xnor U13416 (N_13416,N_12101,N_12574);
nor U13417 (N_13417,N_12256,N_12509);
or U13418 (N_13418,N_12287,N_12597);
xor U13419 (N_13419,N_12490,N_12120);
or U13420 (N_13420,N_12277,N_12608);
nand U13421 (N_13421,N_12393,N_12425);
and U13422 (N_13422,N_12485,N_12079);
nand U13423 (N_13423,N_12303,N_12194);
nand U13424 (N_13424,N_12635,N_12565);
nand U13425 (N_13425,N_12668,N_12594);
and U13426 (N_13426,N_12649,N_12605);
xor U13427 (N_13427,N_12265,N_12115);
nand U13428 (N_13428,N_12319,N_12548);
or U13429 (N_13429,N_12433,N_12499);
nand U13430 (N_13430,N_12402,N_12479);
nor U13431 (N_13431,N_12534,N_12181);
nand U13432 (N_13432,N_12043,N_12185);
and U13433 (N_13433,N_12496,N_12636);
xor U13434 (N_13434,N_12464,N_12502);
nand U13435 (N_13435,N_12274,N_12637);
nand U13436 (N_13436,N_12433,N_12293);
or U13437 (N_13437,N_12664,N_12475);
xnor U13438 (N_13438,N_12532,N_12738);
and U13439 (N_13439,N_12237,N_12626);
nand U13440 (N_13440,N_12306,N_12518);
nor U13441 (N_13441,N_12126,N_12366);
nor U13442 (N_13442,N_12402,N_12284);
nand U13443 (N_13443,N_12546,N_12273);
and U13444 (N_13444,N_12235,N_12202);
nor U13445 (N_13445,N_12138,N_12132);
nand U13446 (N_13446,N_12409,N_12156);
or U13447 (N_13447,N_12711,N_12170);
nand U13448 (N_13448,N_12550,N_12393);
nand U13449 (N_13449,N_12719,N_12598);
nand U13450 (N_13450,N_12637,N_12124);
and U13451 (N_13451,N_12074,N_12625);
xor U13452 (N_13452,N_12723,N_12394);
or U13453 (N_13453,N_12697,N_12301);
and U13454 (N_13454,N_12595,N_12014);
nor U13455 (N_13455,N_12453,N_12233);
and U13456 (N_13456,N_12033,N_12546);
or U13457 (N_13457,N_12617,N_12222);
nor U13458 (N_13458,N_12414,N_12639);
nand U13459 (N_13459,N_12746,N_12702);
or U13460 (N_13460,N_12243,N_12377);
or U13461 (N_13461,N_12574,N_12024);
and U13462 (N_13462,N_12653,N_12338);
or U13463 (N_13463,N_12691,N_12603);
or U13464 (N_13464,N_12460,N_12248);
nand U13465 (N_13465,N_12459,N_12136);
nor U13466 (N_13466,N_12605,N_12680);
nor U13467 (N_13467,N_12113,N_12473);
nor U13468 (N_13468,N_12006,N_12741);
nand U13469 (N_13469,N_12017,N_12173);
or U13470 (N_13470,N_12217,N_12327);
xor U13471 (N_13471,N_12535,N_12130);
xor U13472 (N_13472,N_12594,N_12406);
nor U13473 (N_13473,N_12131,N_12641);
or U13474 (N_13474,N_12708,N_12079);
nor U13475 (N_13475,N_12288,N_12100);
nand U13476 (N_13476,N_12511,N_12645);
and U13477 (N_13477,N_12256,N_12177);
and U13478 (N_13478,N_12735,N_12409);
and U13479 (N_13479,N_12058,N_12185);
nand U13480 (N_13480,N_12100,N_12717);
and U13481 (N_13481,N_12333,N_12044);
or U13482 (N_13482,N_12145,N_12462);
and U13483 (N_13483,N_12054,N_12211);
or U13484 (N_13484,N_12536,N_12622);
nand U13485 (N_13485,N_12275,N_12591);
and U13486 (N_13486,N_12369,N_12527);
nor U13487 (N_13487,N_12022,N_12194);
or U13488 (N_13488,N_12308,N_12651);
and U13489 (N_13489,N_12076,N_12638);
nor U13490 (N_13490,N_12658,N_12585);
and U13491 (N_13491,N_12588,N_12507);
nor U13492 (N_13492,N_12650,N_12298);
nor U13493 (N_13493,N_12403,N_12641);
nand U13494 (N_13494,N_12195,N_12390);
nand U13495 (N_13495,N_12280,N_12534);
and U13496 (N_13496,N_12631,N_12304);
and U13497 (N_13497,N_12134,N_12146);
nor U13498 (N_13498,N_12435,N_12116);
and U13499 (N_13499,N_12746,N_12339);
xor U13500 (N_13500,N_13075,N_13144);
xnor U13501 (N_13501,N_12982,N_13440);
nand U13502 (N_13502,N_12991,N_13277);
xor U13503 (N_13503,N_12972,N_13251);
nand U13504 (N_13504,N_13206,N_12948);
nor U13505 (N_13505,N_12945,N_12808);
and U13506 (N_13506,N_12902,N_12762);
and U13507 (N_13507,N_12780,N_13096);
nor U13508 (N_13508,N_13309,N_13341);
nand U13509 (N_13509,N_12775,N_13246);
nand U13510 (N_13510,N_13190,N_12852);
nand U13511 (N_13511,N_12925,N_13221);
nor U13512 (N_13512,N_12949,N_13281);
nor U13513 (N_13513,N_12952,N_12854);
or U13514 (N_13514,N_13092,N_13237);
or U13515 (N_13515,N_13443,N_13116);
or U13516 (N_13516,N_12855,N_12897);
nand U13517 (N_13517,N_12773,N_13317);
or U13518 (N_13518,N_12983,N_12956);
and U13519 (N_13519,N_13106,N_13180);
or U13520 (N_13520,N_12878,N_13118);
or U13521 (N_13521,N_13271,N_13037);
nand U13522 (N_13522,N_13299,N_12950);
and U13523 (N_13523,N_12926,N_13257);
or U13524 (N_13524,N_13326,N_13377);
nor U13525 (N_13525,N_12896,N_13456);
or U13526 (N_13526,N_13016,N_12984);
nand U13527 (N_13527,N_13064,N_13031);
nand U13528 (N_13528,N_12874,N_12997);
xor U13529 (N_13529,N_12943,N_12848);
and U13530 (N_13530,N_12767,N_13437);
nor U13531 (N_13531,N_12790,N_13347);
nand U13532 (N_13532,N_12901,N_13025);
or U13533 (N_13533,N_13285,N_13234);
nand U13534 (N_13534,N_12799,N_13164);
nor U13535 (N_13535,N_13290,N_13272);
nor U13536 (N_13536,N_13141,N_12832);
or U13537 (N_13537,N_13335,N_12752);
nand U13538 (N_13538,N_12765,N_13266);
and U13539 (N_13539,N_12973,N_13273);
and U13540 (N_13540,N_13430,N_13426);
or U13541 (N_13541,N_13293,N_13094);
nor U13542 (N_13542,N_13315,N_12865);
and U13543 (N_13543,N_13449,N_13466);
or U13544 (N_13544,N_13302,N_13000);
and U13545 (N_13545,N_13334,N_13471);
nand U13546 (N_13546,N_12961,N_13475);
and U13547 (N_13547,N_13413,N_13279);
nor U13548 (N_13548,N_12760,N_13263);
nor U13549 (N_13549,N_13241,N_12922);
nor U13550 (N_13550,N_12846,N_12807);
nor U13551 (N_13551,N_12905,N_13482);
xnor U13552 (N_13552,N_13181,N_13342);
and U13553 (N_13553,N_13483,N_13311);
nor U13554 (N_13554,N_12927,N_12833);
nor U13555 (N_13555,N_13228,N_12797);
nand U13556 (N_13556,N_13052,N_12985);
nor U13557 (N_13557,N_12824,N_13245);
nor U13558 (N_13558,N_12994,N_13170);
nor U13559 (N_13559,N_13236,N_13161);
and U13560 (N_13560,N_13079,N_13336);
and U13561 (N_13561,N_12875,N_13187);
or U13562 (N_13562,N_13403,N_13023);
or U13563 (N_13563,N_12757,N_12754);
nor U13564 (N_13564,N_13287,N_13332);
nand U13565 (N_13565,N_13070,N_12931);
xor U13566 (N_13566,N_12835,N_13423);
and U13567 (N_13567,N_13425,N_13132);
and U13568 (N_13568,N_13200,N_12784);
nand U13569 (N_13569,N_12771,N_13254);
nand U13570 (N_13570,N_13419,N_12890);
nor U13571 (N_13571,N_13265,N_13465);
and U13572 (N_13572,N_13496,N_13422);
nand U13573 (N_13573,N_13223,N_13355);
or U13574 (N_13574,N_13433,N_13148);
and U13575 (N_13575,N_13391,N_12810);
or U13576 (N_13576,N_13091,N_13002);
or U13577 (N_13577,N_12796,N_13343);
nand U13578 (N_13578,N_13415,N_13264);
and U13579 (N_13579,N_13452,N_13358);
and U13580 (N_13580,N_13197,N_13340);
or U13581 (N_13581,N_12763,N_13244);
and U13582 (N_13582,N_13409,N_13369);
nor U13583 (N_13583,N_13169,N_13039);
nand U13584 (N_13584,N_12978,N_12989);
xnor U13585 (N_13585,N_13359,N_13421);
and U13586 (N_13586,N_12840,N_13416);
nand U13587 (N_13587,N_13215,N_13217);
nand U13588 (N_13588,N_13374,N_12960);
or U13589 (N_13589,N_13331,N_13414);
and U13590 (N_13590,N_13247,N_13112);
nand U13591 (N_13591,N_12786,N_13216);
xnor U13592 (N_13592,N_12861,N_13140);
nor U13593 (N_13593,N_12859,N_13153);
or U13594 (N_13594,N_12750,N_13276);
xnor U13595 (N_13595,N_13427,N_13082);
xor U13596 (N_13596,N_13199,N_12867);
nor U13597 (N_13597,N_13213,N_13283);
and U13598 (N_13598,N_13136,N_12766);
and U13599 (N_13599,N_13322,N_13121);
and U13600 (N_13600,N_12975,N_13151);
nor U13601 (N_13601,N_13142,N_13324);
xnor U13602 (N_13602,N_13072,N_12980);
nor U13603 (N_13603,N_13494,N_13020);
or U13604 (N_13604,N_13366,N_13189);
nand U13605 (N_13605,N_13368,N_13120);
and U13606 (N_13606,N_13371,N_12889);
nand U13607 (N_13607,N_13099,N_13435);
xnor U13608 (N_13608,N_12825,N_13364);
or U13609 (N_13609,N_12844,N_13104);
xor U13610 (N_13610,N_13476,N_12959);
or U13611 (N_13611,N_12779,N_12966);
nand U13612 (N_13612,N_12899,N_12849);
xnor U13613 (N_13613,N_12805,N_13387);
or U13614 (N_13614,N_13351,N_12820);
nor U13615 (N_13615,N_13018,N_13110);
nor U13616 (N_13616,N_13318,N_13249);
nand U13617 (N_13617,N_13350,N_13402);
nor U13618 (N_13618,N_13211,N_12962);
nand U13619 (N_13619,N_12774,N_12782);
nor U13620 (N_13620,N_12992,N_13145);
nand U13621 (N_13621,N_13128,N_12813);
or U13622 (N_13622,N_13220,N_13182);
or U13623 (N_13623,N_12898,N_13259);
or U13624 (N_13624,N_12895,N_12803);
nand U13625 (N_13625,N_12798,N_13165);
nand U13626 (N_13626,N_13487,N_13447);
xnor U13627 (N_13627,N_13134,N_13219);
nand U13628 (N_13628,N_13167,N_12804);
and U13629 (N_13629,N_12868,N_13294);
and U13630 (N_13630,N_13146,N_13300);
or U13631 (N_13631,N_13286,N_13485);
nand U13632 (N_13632,N_13231,N_12995);
and U13633 (N_13633,N_13306,N_12826);
or U13634 (N_13634,N_13036,N_12839);
or U13635 (N_13635,N_12955,N_13455);
and U13636 (N_13636,N_13381,N_13101);
nor U13637 (N_13637,N_13460,N_13235);
nand U13638 (N_13638,N_13479,N_12974);
xnor U13639 (N_13639,N_12822,N_12932);
nand U13640 (N_13640,N_13004,N_13090);
nand U13641 (N_13641,N_13394,N_13345);
or U13642 (N_13642,N_13208,N_13133);
and U13643 (N_13643,N_13308,N_13348);
nand U13644 (N_13644,N_13401,N_13115);
or U13645 (N_13645,N_13379,N_13207);
nor U13646 (N_13646,N_13323,N_13418);
nand U13647 (N_13647,N_12892,N_13178);
nand U13648 (N_13648,N_13086,N_12823);
or U13649 (N_13649,N_12977,N_13212);
nand U13650 (N_13650,N_12979,N_13360);
nor U13651 (N_13651,N_13058,N_12800);
nor U13652 (N_13652,N_13319,N_13149);
or U13653 (N_13653,N_13222,N_13367);
or U13654 (N_13654,N_13390,N_13399);
or U13655 (N_13655,N_12853,N_13174);
nor U13656 (N_13656,N_13473,N_13489);
nor U13657 (N_13657,N_13051,N_12887);
nor U13658 (N_13658,N_13453,N_13375);
or U13659 (N_13659,N_13188,N_13383);
nand U13660 (N_13660,N_13400,N_13396);
or U13661 (N_13661,N_12769,N_13233);
or U13662 (N_13662,N_12812,N_12930);
nor U13663 (N_13663,N_12764,N_13130);
or U13664 (N_13664,N_13119,N_13229);
nand U13665 (N_13665,N_13061,N_13314);
nand U13666 (N_13666,N_13410,N_12879);
nor U13667 (N_13667,N_12967,N_13108);
nor U13668 (N_13668,N_13327,N_13202);
and U13669 (N_13669,N_13370,N_13027);
and U13670 (N_13670,N_13258,N_13005);
xnor U13671 (N_13671,N_13050,N_12951);
and U13672 (N_13672,N_12888,N_12891);
and U13673 (N_13673,N_13313,N_13282);
nor U13674 (N_13674,N_13139,N_13382);
and U13675 (N_13675,N_12998,N_13491);
nor U13676 (N_13676,N_13441,N_12876);
and U13677 (N_13677,N_13068,N_13467);
nor U13678 (N_13678,N_13218,N_12870);
nor U13679 (N_13679,N_12776,N_13480);
and U13680 (N_13680,N_13166,N_13123);
nand U13681 (N_13681,N_13150,N_13495);
nor U13682 (N_13682,N_13095,N_12919);
nor U13683 (N_13683,N_13275,N_13038);
nor U13684 (N_13684,N_13284,N_13291);
xnor U13685 (N_13685,N_13474,N_13349);
and U13686 (N_13686,N_13261,N_12830);
nor U13687 (N_13687,N_13014,N_13227);
or U13688 (N_13688,N_12860,N_12828);
or U13689 (N_13689,N_13310,N_13298);
nand U13690 (N_13690,N_13124,N_13365);
or U13691 (N_13691,N_12903,N_13089);
and U13692 (N_13692,N_13262,N_13209);
nand U13693 (N_13693,N_13439,N_13172);
and U13694 (N_13694,N_12885,N_12871);
and U13695 (N_13695,N_12946,N_12916);
or U13696 (N_13696,N_12882,N_13238);
nor U13697 (N_13697,N_13003,N_13029);
and U13698 (N_13698,N_13183,N_13492);
and U13699 (N_13699,N_13446,N_13088);
nor U13700 (N_13700,N_13363,N_13329);
nand U13701 (N_13701,N_12827,N_12965);
and U13702 (N_13702,N_12912,N_13191);
or U13703 (N_13703,N_13067,N_13267);
xor U13704 (N_13704,N_13454,N_12829);
nor U13705 (N_13705,N_13010,N_13226);
or U13706 (N_13706,N_13295,N_13129);
nand U13707 (N_13707,N_13252,N_12838);
and U13708 (N_13708,N_13011,N_13021);
nor U13709 (N_13709,N_13076,N_13232);
nand U13710 (N_13710,N_13185,N_13472);
xor U13711 (N_13711,N_13389,N_12924);
nand U13712 (N_13712,N_12938,N_13077);
and U13713 (N_13713,N_12993,N_12850);
xnor U13714 (N_13714,N_13464,N_12866);
or U13715 (N_13715,N_13179,N_13204);
xnor U13716 (N_13716,N_12969,N_12893);
or U13717 (N_13717,N_13147,N_13040);
and U13718 (N_13718,N_13325,N_13434);
nand U13719 (N_13719,N_12759,N_13143);
or U13720 (N_13720,N_13160,N_12857);
or U13721 (N_13721,N_13429,N_12845);
and U13722 (N_13722,N_13488,N_12792);
and U13723 (N_13723,N_13321,N_13184);
or U13724 (N_13724,N_13412,N_13162);
or U13725 (N_13725,N_13111,N_13289);
or U13726 (N_13726,N_13156,N_12806);
and U13727 (N_13727,N_13013,N_13431);
or U13728 (N_13728,N_13035,N_13084);
and U13729 (N_13729,N_13034,N_13356);
nand U13730 (N_13730,N_13225,N_13346);
or U13731 (N_13731,N_13171,N_13044);
or U13732 (N_13732,N_13239,N_12751);
nor U13733 (N_13733,N_13097,N_13063);
and U13734 (N_13734,N_12939,N_13357);
and U13735 (N_13735,N_13354,N_13404);
or U13736 (N_13736,N_13320,N_12834);
nand U13737 (N_13737,N_13372,N_13192);
nor U13738 (N_13738,N_13380,N_13022);
or U13739 (N_13739,N_13378,N_13490);
or U13740 (N_13740,N_12787,N_12886);
or U13741 (N_13741,N_13296,N_12831);
xor U13742 (N_13742,N_13376,N_13292);
and U13743 (N_13743,N_13053,N_13468);
and U13744 (N_13744,N_13459,N_12957);
and U13745 (N_13745,N_12781,N_13457);
nand U13746 (N_13746,N_13493,N_13499);
nand U13747 (N_13747,N_13196,N_12947);
nor U13748 (N_13748,N_13138,N_12819);
or U13749 (N_13749,N_13337,N_13019);
and U13750 (N_13750,N_12909,N_13069);
and U13751 (N_13751,N_13477,N_13102);
nor U13752 (N_13752,N_13408,N_12811);
or U13753 (N_13753,N_13484,N_12772);
and U13754 (N_13754,N_13081,N_13428);
nor U13755 (N_13755,N_13385,N_13157);
or U13756 (N_13756,N_13195,N_13497);
xnor U13757 (N_13757,N_12758,N_12981);
and U13758 (N_13758,N_13352,N_13126);
nand U13759 (N_13759,N_12935,N_13339);
xor U13760 (N_13760,N_13248,N_13158);
nand U13761 (N_13761,N_13193,N_13398);
xor U13762 (N_13762,N_12785,N_12999);
xnor U13763 (N_13763,N_13127,N_13303);
or U13764 (N_13764,N_13333,N_13113);
nor U13765 (N_13765,N_12869,N_13280);
nor U13766 (N_13766,N_13451,N_12953);
xor U13767 (N_13767,N_13085,N_12964);
nor U13768 (N_13768,N_12988,N_13159);
and U13769 (N_13769,N_12880,N_13288);
nor U13770 (N_13770,N_12802,N_12937);
nand U13771 (N_13771,N_13201,N_12929);
nor U13772 (N_13772,N_12881,N_12788);
or U13773 (N_13773,N_13393,N_13442);
nand U13774 (N_13774,N_13463,N_13253);
xnor U13775 (N_13775,N_13330,N_13041);
or U13776 (N_13776,N_13436,N_13012);
and U13777 (N_13777,N_12917,N_13105);
and U13778 (N_13778,N_13131,N_13424);
and U13779 (N_13779,N_13344,N_12856);
xnor U13780 (N_13780,N_13045,N_13107);
nand U13781 (N_13781,N_13270,N_12971);
or U13782 (N_13782,N_12944,N_13186);
and U13783 (N_13783,N_12783,N_13420);
nor U13784 (N_13784,N_13312,N_12911);
or U13785 (N_13785,N_12816,N_13210);
or U13786 (N_13786,N_13194,N_13250);
xor U13787 (N_13787,N_12918,N_12941);
nand U13788 (N_13788,N_13224,N_13015);
nand U13789 (N_13789,N_13461,N_13498);
or U13790 (N_13790,N_13049,N_12873);
and U13791 (N_13791,N_13432,N_12864);
and U13792 (N_13792,N_12847,N_12913);
or U13793 (N_13793,N_12794,N_13009);
nand U13794 (N_13794,N_13033,N_13297);
and U13795 (N_13795,N_12791,N_13066);
xor U13796 (N_13796,N_12914,N_12778);
or U13797 (N_13797,N_13074,N_13243);
or U13798 (N_13798,N_12921,N_12795);
and U13799 (N_13799,N_13054,N_12801);
and U13800 (N_13800,N_12862,N_13163);
nor U13801 (N_13801,N_13080,N_13007);
nor U13802 (N_13802,N_12920,N_13417);
or U13803 (N_13803,N_13056,N_13278);
and U13804 (N_13804,N_12915,N_12894);
nand U13805 (N_13805,N_13205,N_13406);
or U13806 (N_13806,N_12936,N_13448);
nand U13807 (N_13807,N_13307,N_12877);
xor U13808 (N_13808,N_12817,N_12872);
and U13809 (N_13809,N_12933,N_12863);
or U13810 (N_13810,N_13316,N_13047);
or U13811 (N_13811,N_12923,N_13006);
nand U13812 (N_13812,N_13444,N_13438);
nand U13813 (N_13813,N_13135,N_13478);
nor U13814 (N_13814,N_13203,N_12841);
or U13815 (N_13815,N_13328,N_12768);
nand U13816 (N_13816,N_12907,N_13073);
or U13817 (N_13817,N_12908,N_13361);
nand U13818 (N_13818,N_13043,N_13030);
nor U13819 (N_13819,N_13304,N_13032);
or U13820 (N_13820,N_13230,N_12987);
and U13821 (N_13821,N_13268,N_13395);
and U13822 (N_13822,N_13042,N_13384);
and U13823 (N_13823,N_12793,N_13458);
nor U13824 (N_13824,N_13462,N_13411);
nand U13825 (N_13825,N_13173,N_13445);
and U13826 (N_13826,N_13198,N_13008);
and U13827 (N_13827,N_13386,N_12815);
xor U13828 (N_13828,N_12996,N_12954);
or U13829 (N_13829,N_12858,N_13175);
or U13830 (N_13830,N_12842,N_13117);
nand U13831 (N_13831,N_13305,N_13214);
and U13832 (N_13832,N_13098,N_13152);
or U13833 (N_13833,N_13071,N_12968);
nand U13834 (N_13834,N_13001,N_13450);
or U13835 (N_13835,N_13055,N_13155);
nor U13836 (N_13836,N_12836,N_13397);
nand U13837 (N_13837,N_13046,N_13114);
nor U13838 (N_13838,N_13122,N_13405);
and U13839 (N_13839,N_13059,N_13469);
and U13840 (N_13840,N_13256,N_12963);
nor U13841 (N_13841,N_13060,N_12934);
xor U13842 (N_13842,N_12789,N_12753);
nand U13843 (N_13843,N_12756,N_12777);
and U13844 (N_13844,N_12990,N_12986);
and U13845 (N_13845,N_13240,N_12970);
or U13846 (N_13846,N_12884,N_13176);
nor U13847 (N_13847,N_12904,N_13470);
or U13848 (N_13848,N_12942,N_13065);
nand U13849 (N_13849,N_13373,N_13362);
nand U13850 (N_13850,N_12851,N_13125);
and U13851 (N_13851,N_13026,N_12976);
nor U13852 (N_13852,N_12883,N_13338);
nand U13853 (N_13853,N_13083,N_12761);
nor U13854 (N_13854,N_13301,N_12818);
nor U13855 (N_13855,N_13260,N_12928);
or U13856 (N_13856,N_12843,N_13168);
or U13857 (N_13857,N_12814,N_12837);
or U13858 (N_13858,N_13017,N_13388);
and U13859 (N_13859,N_13100,N_12900);
nand U13860 (N_13860,N_13154,N_12958);
nand U13861 (N_13861,N_13078,N_12940);
nor U13862 (N_13862,N_12906,N_13274);
nor U13863 (N_13863,N_13087,N_12910);
xor U13864 (N_13864,N_13486,N_13177);
nor U13865 (N_13865,N_12755,N_13057);
xnor U13866 (N_13866,N_12809,N_13137);
and U13867 (N_13867,N_13109,N_13062);
and U13868 (N_13868,N_13481,N_13353);
and U13869 (N_13869,N_13093,N_13028);
nor U13870 (N_13870,N_13242,N_13048);
nor U13871 (N_13871,N_13255,N_13392);
and U13872 (N_13872,N_13407,N_12821);
xor U13873 (N_13873,N_13103,N_13024);
or U13874 (N_13874,N_13269,N_12770);
nor U13875 (N_13875,N_13192,N_13000);
or U13876 (N_13876,N_13094,N_12845);
nand U13877 (N_13877,N_13207,N_12753);
nor U13878 (N_13878,N_12816,N_13059);
or U13879 (N_13879,N_13334,N_13278);
and U13880 (N_13880,N_13313,N_12765);
xnor U13881 (N_13881,N_12936,N_13055);
or U13882 (N_13882,N_13172,N_13321);
or U13883 (N_13883,N_13200,N_13123);
nand U13884 (N_13884,N_13015,N_13148);
or U13885 (N_13885,N_13401,N_12967);
and U13886 (N_13886,N_13268,N_13338);
nand U13887 (N_13887,N_13175,N_12938);
nor U13888 (N_13888,N_13142,N_12817);
or U13889 (N_13889,N_13298,N_12764);
nor U13890 (N_13890,N_12850,N_13220);
xor U13891 (N_13891,N_12996,N_13442);
and U13892 (N_13892,N_13488,N_13229);
and U13893 (N_13893,N_12984,N_13475);
or U13894 (N_13894,N_13075,N_13457);
nand U13895 (N_13895,N_13266,N_13115);
and U13896 (N_13896,N_13107,N_13411);
and U13897 (N_13897,N_13202,N_12911);
xor U13898 (N_13898,N_12868,N_13009);
or U13899 (N_13899,N_13275,N_12885);
and U13900 (N_13900,N_12971,N_13475);
or U13901 (N_13901,N_13466,N_13362);
nand U13902 (N_13902,N_13422,N_13095);
or U13903 (N_13903,N_13120,N_13103);
or U13904 (N_13904,N_12900,N_13264);
xnor U13905 (N_13905,N_13286,N_13403);
and U13906 (N_13906,N_12922,N_13080);
nor U13907 (N_13907,N_12903,N_12975);
and U13908 (N_13908,N_12902,N_13204);
and U13909 (N_13909,N_13177,N_13325);
xor U13910 (N_13910,N_12761,N_12904);
and U13911 (N_13911,N_13428,N_13461);
nor U13912 (N_13912,N_13408,N_12789);
and U13913 (N_13913,N_13340,N_12901);
nor U13914 (N_13914,N_12940,N_13290);
xor U13915 (N_13915,N_13335,N_13132);
and U13916 (N_13916,N_12962,N_13131);
or U13917 (N_13917,N_13138,N_13239);
nand U13918 (N_13918,N_12980,N_12822);
or U13919 (N_13919,N_12935,N_13072);
nor U13920 (N_13920,N_13410,N_12834);
or U13921 (N_13921,N_13147,N_13245);
nor U13922 (N_13922,N_13277,N_13200);
nand U13923 (N_13923,N_13401,N_12822);
or U13924 (N_13924,N_12927,N_13258);
nand U13925 (N_13925,N_12804,N_13495);
nand U13926 (N_13926,N_12809,N_13134);
nor U13927 (N_13927,N_12963,N_12765);
and U13928 (N_13928,N_12790,N_13160);
nand U13929 (N_13929,N_13197,N_13055);
nor U13930 (N_13930,N_13135,N_13056);
and U13931 (N_13931,N_12868,N_13499);
nor U13932 (N_13932,N_13178,N_12784);
nand U13933 (N_13933,N_13474,N_13449);
nor U13934 (N_13934,N_13478,N_13452);
nand U13935 (N_13935,N_13394,N_13029);
nor U13936 (N_13936,N_13200,N_13311);
xor U13937 (N_13937,N_13464,N_13245);
nand U13938 (N_13938,N_13238,N_13233);
nand U13939 (N_13939,N_13062,N_12767);
nand U13940 (N_13940,N_12793,N_13405);
nand U13941 (N_13941,N_12824,N_13138);
and U13942 (N_13942,N_13256,N_12832);
xor U13943 (N_13943,N_13147,N_13095);
nand U13944 (N_13944,N_13038,N_13376);
nor U13945 (N_13945,N_13064,N_13282);
or U13946 (N_13946,N_13182,N_12776);
and U13947 (N_13947,N_13238,N_13414);
and U13948 (N_13948,N_12988,N_13080);
nor U13949 (N_13949,N_12887,N_13445);
nand U13950 (N_13950,N_12920,N_12822);
or U13951 (N_13951,N_12761,N_13170);
xor U13952 (N_13952,N_13265,N_13183);
or U13953 (N_13953,N_12880,N_12881);
and U13954 (N_13954,N_12773,N_12957);
xor U13955 (N_13955,N_13029,N_13229);
or U13956 (N_13956,N_13126,N_12994);
nor U13957 (N_13957,N_12887,N_13114);
nor U13958 (N_13958,N_12767,N_13229);
nand U13959 (N_13959,N_13185,N_13007);
or U13960 (N_13960,N_13113,N_13084);
nor U13961 (N_13961,N_13339,N_13079);
nor U13962 (N_13962,N_12857,N_13485);
nor U13963 (N_13963,N_13168,N_13222);
xnor U13964 (N_13964,N_13242,N_13169);
or U13965 (N_13965,N_12873,N_12800);
nor U13966 (N_13966,N_12915,N_12954);
nand U13967 (N_13967,N_13404,N_12835);
and U13968 (N_13968,N_12924,N_13371);
or U13969 (N_13969,N_12784,N_13480);
xnor U13970 (N_13970,N_13002,N_13266);
xnor U13971 (N_13971,N_13427,N_13285);
and U13972 (N_13972,N_13171,N_13079);
nand U13973 (N_13973,N_12915,N_13315);
nand U13974 (N_13974,N_13164,N_13406);
or U13975 (N_13975,N_12892,N_13077);
nand U13976 (N_13976,N_12876,N_13051);
xnor U13977 (N_13977,N_12948,N_13311);
xnor U13978 (N_13978,N_13325,N_13246);
or U13979 (N_13979,N_13408,N_12881);
or U13980 (N_13980,N_13342,N_13301);
or U13981 (N_13981,N_13372,N_13335);
nand U13982 (N_13982,N_12894,N_12948);
or U13983 (N_13983,N_12922,N_13224);
or U13984 (N_13984,N_13254,N_13251);
xnor U13985 (N_13985,N_13264,N_13261);
and U13986 (N_13986,N_13073,N_12919);
and U13987 (N_13987,N_13092,N_13456);
nor U13988 (N_13988,N_12754,N_13472);
xnor U13989 (N_13989,N_13133,N_13443);
nor U13990 (N_13990,N_13399,N_13322);
nor U13991 (N_13991,N_13227,N_13419);
xnor U13992 (N_13992,N_13218,N_13477);
nand U13993 (N_13993,N_13396,N_13476);
nor U13994 (N_13994,N_12836,N_12911);
nor U13995 (N_13995,N_13319,N_12846);
nor U13996 (N_13996,N_13078,N_12770);
xnor U13997 (N_13997,N_13261,N_12809);
nand U13998 (N_13998,N_13378,N_12864);
nor U13999 (N_13999,N_13030,N_13072);
and U14000 (N_14000,N_12891,N_13391);
and U14001 (N_14001,N_12905,N_13005);
or U14002 (N_14002,N_12887,N_13045);
nand U14003 (N_14003,N_13014,N_12995);
or U14004 (N_14004,N_13255,N_13251);
xnor U14005 (N_14005,N_12785,N_13100);
nor U14006 (N_14006,N_13401,N_13102);
or U14007 (N_14007,N_12911,N_12800);
nor U14008 (N_14008,N_13284,N_13160);
or U14009 (N_14009,N_12875,N_12987);
nand U14010 (N_14010,N_13367,N_12969);
and U14011 (N_14011,N_13129,N_12776);
nand U14012 (N_14012,N_13318,N_13313);
nor U14013 (N_14013,N_13082,N_12880);
xnor U14014 (N_14014,N_13426,N_12885);
or U14015 (N_14015,N_13244,N_12905);
or U14016 (N_14016,N_12936,N_12839);
or U14017 (N_14017,N_13234,N_12811);
nand U14018 (N_14018,N_13460,N_12805);
nand U14019 (N_14019,N_13047,N_13271);
nand U14020 (N_14020,N_12889,N_13315);
and U14021 (N_14021,N_12925,N_12899);
or U14022 (N_14022,N_13043,N_13177);
and U14023 (N_14023,N_13260,N_13094);
nor U14024 (N_14024,N_12767,N_12892);
and U14025 (N_14025,N_12950,N_12840);
nor U14026 (N_14026,N_12778,N_13432);
and U14027 (N_14027,N_13397,N_13469);
nand U14028 (N_14028,N_12804,N_13001);
and U14029 (N_14029,N_13317,N_13496);
or U14030 (N_14030,N_13288,N_13058);
nand U14031 (N_14031,N_13397,N_13210);
and U14032 (N_14032,N_13478,N_13436);
xor U14033 (N_14033,N_13090,N_12849);
and U14034 (N_14034,N_13346,N_12797);
and U14035 (N_14035,N_13369,N_12925);
or U14036 (N_14036,N_12884,N_13349);
or U14037 (N_14037,N_13341,N_13177);
or U14038 (N_14038,N_13243,N_13460);
nand U14039 (N_14039,N_13191,N_13440);
nor U14040 (N_14040,N_13069,N_12843);
and U14041 (N_14041,N_13333,N_12818);
xnor U14042 (N_14042,N_13449,N_13044);
or U14043 (N_14043,N_12765,N_13044);
and U14044 (N_14044,N_12906,N_12945);
nor U14045 (N_14045,N_12974,N_12835);
nand U14046 (N_14046,N_13271,N_12836);
nor U14047 (N_14047,N_13430,N_12953);
nand U14048 (N_14048,N_12769,N_12820);
or U14049 (N_14049,N_13491,N_13454);
xnor U14050 (N_14050,N_12967,N_12794);
nand U14051 (N_14051,N_13150,N_12891);
and U14052 (N_14052,N_13038,N_12764);
nor U14053 (N_14053,N_13183,N_13219);
and U14054 (N_14054,N_12893,N_13220);
nand U14055 (N_14055,N_13323,N_13336);
nor U14056 (N_14056,N_12893,N_12783);
nor U14057 (N_14057,N_12960,N_12789);
or U14058 (N_14058,N_13297,N_13177);
nand U14059 (N_14059,N_13377,N_13245);
nor U14060 (N_14060,N_13278,N_13282);
nor U14061 (N_14061,N_13031,N_13279);
nand U14062 (N_14062,N_13167,N_13285);
or U14063 (N_14063,N_12926,N_13140);
nand U14064 (N_14064,N_13002,N_13312);
and U14065 (N_14065,N_13412,N_13382);
or U14066 (N_14066,N_13131,N_13457);
nor U14067 (N_14067,N_13226,N_13328);
or U14068 (N_14068,N_13089,N_13286);
xnor U14069 (N_14069,N_13020,N_12864);
or U14070 (N_14070,N_12964,N_12776);
nor U14071 (N_14071,N_13335,N_13068);
nor U14072 (N_14072,N_13041,N_13074);
nor U14073 (N_14073,N_13344,N_12935);
and U14074 (N_14074,N_12758,N_13018);
and U14075 (N_14075,N_13391,N_12924);
nand U14076 (N_14076,N_12877,N_12944);
nand U14077 (N_14077,N_12974,N_13443);
and U14078 (N_14078,N_13486,N_13314);
and U14079 (N_14079,N_13131,N_13383);
and U14080 (N_14080,N_13373,N_12890);
nand U14081 (N_14081,N_13204,N_13221);
nor U14082 (N_14082,N_12894,N_12778);
nand U14083 (N_14083,N_13451,N_12896);
or U14084 (N_14084,N_13432,N_13268);
nand U14085 (N_14085,N_13395,N_13297);
or U14086 (N_14086,N_12754,N_13291);
xnor U14087 (N_14087,N_12814,N_13317);
and U14088 (N_14088,N_13407,N_13367);
nand U14089 (N_14089,N_12957,N_12997);
or U14090 (N_14090,N_12811,N_13452);
or U14091 (N_14091,N_13393,N_13444);
nor U14092 (N_14092,N_13471,N_12825);
and U14093 (N_14093,N_13245,N_12803);
or U14094 (N_14094,N_12913,N_13133);
and U14095 (N_14095,N_13425,N_13486);
nand U14096 (N_14096,N_13420,N_12897);
nand U14097 (N_14097,N_12818,N_13385);
nand U14098 (N_14098,N_12871,N_13370);
or U14099 (N_14099,N_13232,N_12890);
and U14100 (N_14100,N_13315,N_13217);
nand U14101 (N_14101,N_13017,N_13177);
xnor U14102 (N_14102,N_13388,N_13076);
and U14103 (N_14103,N_13234,N_12816);
xor U14104 (N_14104,N_13412,N_12758);
or U14105 (N_14105,N_13108,N_13260);
or U14106 (N_14106,N_13047,N_12841);
nor U14107 (N_14107,N_13269,N_13150);
and U14108 (N_14108,N_13230,N_13085);
nand U14109 (N_14109,N_13357,N_12874);
nor U14110 (N_14110,N_12901,N_12966);
and U14111 (N_14111,N_12786,N_12832);
or U14112 (N_14112,N_13463,N_12821);
nand U14113 (N_14113,N_12913,N_12905);
or U14114 (N_14114,N_12865,N_13204);
xor U14115 (N_14115,N_12792,N_12904);
nor U14116 (N_14116,N_13414,N_13408);
nand U14117 (N_14117,N_12940,N_12818);
nand U14118 (N_14118,N_13125,N_12823);
nor U14119 (N_14119,N_12771,N_13456);
nor U14120 (N_14120,N_13087,N_13045);
nor U14121 (N_14121,N_13212,N_12942);
or U14122 (N_14122,N_12867,N_13083);
or U14123 (N_14123,N_12915,N_12933);
nand U14124 (N_14124,N_12970,N_13018);
nor U14125 (N_14125,N_13459,N_13086);
or U14126 (N_14126,N_13275,N_12833);
or U14127 (N_14127,N_12988,N_13386);
nand U14128 (N_14128,N_12930,N_12927);
or U14129 (N_14129,N_13142,N_12989);
or U14130 (N_14130,N_13250,N_13229);
nor U14131 (N_14131,N_12790,N_13179);
or U14132 (N_14132,N_13171,N_13235);
nor U14133 (N_14133,N_13352,N_13006);
or U14134 (N_14134,N_13482,N_12985);
nor U14135 (N_14135,N_13081,N_13369);
or U14136 (N_14136,N_13110,N_13249);
and U14137 (N_14137,N_13337,N_13392);
and U14138 (N_14138,N_12808,N_13380);
or U14139 (N_14139,N_13397,N_13201);
or U14140 (N_14140,N_13345,N_13213);
nor U14141 (N_14141,N_12994,N_13287);
nor U14142 (N_14142,N_13262,N_13492);
nor U14143 (N_14143,N_13106,N_12953);
nand U14144 (N_14144,N_13084,N_13081);
nand U14145 (N_14145,N_13224,N_12983);
or U14146 (N_14146,N_13177,N_12946);
and U14147 (N_14147,N_13380,N_12963);
nor U14148 (N_14148,N_12769,N_13448);
xnor U14149 (N_14149,N_12861,N_13286);
nand U14150 (N_14150,N_13389,N_13271);
nand U14151 (N_14151,N_13372,N_13403);
or U14152 (N_14152,N_13006,N_12797);
nor U14153 (N_14153,N_13455,N_13367);
or U14154 (N_14154,N_13421,N_13458);
and U14155 (N_14155,N_13428,N_13356);
and U14156 (N_14156,N_13373,N_13458);
or U14157 (N_14157,N_13400,N_13475);
and U14158 (N_14158,N_13157,N_13052);
and U14159 (N_14159,N_13237,N_13219);
or U14160 (N_14160,N_13442,N_13255);
or U14161 (N_14161,N_12873,N_12903);
nand U14162 (N_14162,N_13061,N_12769);
nor U14163 (N_14163,N_13251,N_13340);
or U14164 (N_14164,N_13119,N_12853);
and U14165 (N_14165,N_12903,N_12806);
nor U14166 (N_14166,N_12862,N_13446);
xor U14167 (N_14167,N_13159,N_13331);
and U14168 (N_14168,N_12952,N_13272);
nor U14169 (N_14169,N_13114,N_13230);
or U14170 (N_14170,N_12975,N_13019);
nand U14171 (N_14171,N_13387,N_13459);
or U14172 (N_14172,N_12957,N_13081);
nor U14173 (N_14173,N_13039,N_13100);
xor U14174 (N_14174,N_13252,N_12962);
or U14175 (N_14175,N_12986,N_13424);
nor U14176 (N_14176,N_12766,N_12892);
and U14177 (N_14177,N_13484,N_13401);
or U14178 (N_14178,N_13304,N_12936);
and U14179 (N_14179,N_13426,N_13228);
nand U14180 (N_14180,N_13387,N_12920);
nor U14181 (N_14181,N_12899,N_13413);
xor U14182 (N_14182,N_13199,N_12892);
and U14183 (N_14183,N_13073,N_13146);
nor U14184 (N_14184,N_12943,N_13124);
xnor U14185 (N_14185,N_12914,N_13116);
nand U14186 (N_14186,N_12998,N_12762);
or U14187 (N_14187,N_13368,N_12837);
nor U14188 (N_14188,N_12765,N_13033);
nor U14189 (N_14189,N_12755,N_13102);
and U14190 (N_14190,N_13253,N_13353);
and U14191 (N_14191,N_13200,N_12797);
nand U14192 (N_14192,N_13149,N_13055);
and U14193 (N_14193,N_13365,N_13476);
nor U14194 (N_14194,N_12783,N_13025);
or U14195 (N_14195,N_13042,N_12882);
and U14196 (N_14196,N_12798,N_13379);
or U14197 (N_14197,N_13127,N_13464);
nor U14198 (N_14198,N_12975,N_13457);
and U14199 (N_14199,N_13252,N_13150);
or U14200 (N_14200,N_12884,N_13365);
and U14201 (N_14201,N_13457,N_13134);
nor U14202 (N_14202,N_13046,N_12783);
and U14203 (N_14203,N_12784,N_12976);
or U14204 (N_14204,N_13499,N_12928);
nor U14205 (N_14205,N_13127,N_13091);
and U14206 (N_14206,N_13327,N_12758);
or U14207 (N_14207,N_13114,N_12996);
or U14208 (N_14208,N_13162,N_13426);
nor U14209 (N_14209,N_13369,N_12938);
and U14210 (N_14210,N_12904,N_13281);
or U14211 (N_14211,N_12765,N_13375);
and U14212 (N_14212,N_12908,N_13012);
or U14213 (N_14213,N_13305,N_12870);
and U14214 (N_14214,N_13462,N_12957);
or U14215 (N_14215,N_12805,N_13473);
nor U14216 (N_14216,N_12900,N_13278);
nor U14217 (N_14217,N_13434,N_12778);
nand U14218 (N_14218,N_12842,N_13261);
and U14219 (N_14219,N_12760,N_13042);
and U14220 (N_14220,N_12820,N_13139);
and U14221 (N_14221,N_12818,N_13370);
or U14222 (N_14222,N_12871,N_12966);
or U14223 (N_14223,N_13182,N_12991);
and U14224 (N_14224,N_12908,N_12984);
and U14225 (N_14225,N_12878,N_12962);
nor U14226 (N_14226,N_13201,N_13323);
or U14227 (N_14227,N_13310,N_13394);
and U14228 (N_14228,N_12801,N_12943);
nor U14229 (N_14229,N_13075,N_13198);
nor U14230 (N_14230,N_13398,N_12938);
nand U14231 (N_14231,N_12806,N_13292);
nand U14232 (N_14232,N_12985,N_12774);
nand U14233 (N_14233,N_12857,N_13362);
and U14234 (N_14234,N_13490,N_12909);
or U14235 (N_14235,N_13217,N_13127);
and U14236 (N_14236,N_13205,N_13021);
nand U14237 (N_14237,N_13143,N_13323);
nand U14238 (N_14238,N_12983,N_13120);
nand U14239 (N_14239,N_12846,N_12852);
and U14240 (N_14240,N_13072,N_12879);
nand U14241 (N_14241,N_13184,N_12955);
nor U14242 (N_14242,N_13256,N_12946);
or U14243 (N_14243,N_13251,N_13352);
xnor U14244 (N_14244,N_12834,N_12938);
and U14245 (N_14245,N_13207,N_13398);
nor U14246 (N_14246,N_12834,N_13495);
and U14247 (N_14247,N_13144,N_13217);
nand U14248 (N_14248,N_13468,N_13457);
nor U14249 (N_14249,N_13445,N_13125);
nand U14250 (N_14250,N_13767,N_13817);
and U14251 (N_14251,N_13780,N_13657);
xor U14252 (N_14252,N_14177,N_13985);
xnor U14253 (N_14253,N_13892,N_13688);
and U14254 (N_14254,N_14139,N_13515);
nor U14255 (N_14255,N_13638,N_14002);
nand U14256 (N_14256,N_13570,N_14179);
or U14257 (N_14257,N_13874,N_13619);
and U14258 (N_14258,N_13875,N_13683);
xnor U14259 (N_14259,N_13805,N_13562);
nand U14260 (N_14260,N_13753,N_13860);
or U14261 (N_14261,N_14052,N_13856);
and U14262 (N_14262,N_13653,N_13741);
or U14263 (N_14263,N_13757,N_14186);
and U14264 (N_14264,N_14083,N_14201);
or U14265 (N_14265,N_13525,N_13876);
nand U14266 (N_14266,N_14023,N_13977);
nand U14267 (N_14267,N_13520,N_13691);
or U14268 (N_14268,N_14075,N_13821);
nor U14269 (N_14269,N_13703,N_14035);
and U14270 (N_14270,N_13877,N_13981);
nor U14271 (N_14271,N_14150,N_14209);
nand U14272 (N_14272,N_13640,N_13958);
nor U14273 (N_14273,N_13716,N_13695);
nor U14274 (N_14274,N_13844,N_13933);
nand U14275 (N_14275,N_14088,N_13715);
and U14276 (N_14276,N_13663,N_13778);
nor U14277 (N_14277,N_13847,N_13647);
nand U14278 (N_14278,N_14025,N_13689);
nand U14279 (N_14279,N_14232,N_14077);
nor U14280 (N_14280,N_13552,N_13983);
and U14281 (N_14281,N_13781,N_13554);
nor U14282 (N_14282,N_13928,N_13761);
xor U14283 (N_14283,N_14247,N_13807);
nand U14284 (N_14284,N_13600,N_13564);
or U14285 (N_14285,N_14159,N_14029);
nor U14286 (N_14286,N_13585,N_13690);
nor U14287 (N_14287,N_13698,N_14061);
nor U14288 (N_14288,N_13718,N_13998);
nand U14289 (N_14289,N_14093,N_13617);
and U14290 (N_14290,N_13541,N_14102);
and U14291 (N_14291,N_14234,N_14231);
and U14292 (N_14292,N_14095,N_13957);
xor U14293 (N_14293,N_13586,N_14031);
nor U14294 (N_14294,N_13924,N_14187);
and U14295 (N_14295,N_13526,N_14069);
nand U14296 (N_14296,N_13889,N_14239);
nand U14297 (N_14297,N_13976,N_14063);
nor U14298 (N_14298,N_14181,N_13575);
and U14299 (N_14299,N_13838,N_13758);
or U14300 (N_14300,N_14018,N_14017);
nand U14301 (N_14301,N_14005,N_14055);
or U14302 (N_14302,N_14195,N_13770);
nor U14303 (N_14303,N_13738,N_14078);
or U14304 (N_14304,N_13936,N_13929);
or U14305 (N_14305,N_13605,N_13872);
and U14306 (N_14306,N_13886,N_13862);
nor U14307 (N_14307,N_14240,N_14236);
or U14308 (N_14308,N_13722,N_13949);
nor U14309 (N_14309,N_13907,N_14176);
nor U14310 (N_14310,N_13991,N_13988);
nand U14311 (N_14311,N_13651,N_14051);
or U14312 (N_14312,N_14060,N_13595);
and U14313 (N_14313,N_14098,N_13662);
nand U14314 (N_14314,N_13978,N_13707);
nand U14315 (N_14315,N_13890,N_13545);
nor U14316 (N_14316,N_14110,N_13628);
nor U14317 (N_14317,N_13742,N_13669);
or U14318 (N_14318,N_13516,N_14070);
nand U14319 (N_14319,N_13547,N_13550);
and U14320 (N_14320,N_14114,N_13711);
and U14321 (N_14321,N_13896,N_13814);
xor U14322 (N_14322,N_14185,N_14022);
nor U14323 (N_14323,N_13897,N_14219);
nand U14324 (N_14324,N_13563,N_13580);
nand U14325 (N_14325,N_13645,N_14246);
or U14326 (N_14326,N_13732,N_13577);
nor U14327 (N_14327,N_13713,N_13754);
nand U14328 (N_14328,N_13675,N_13996);
and U14329 (N_14329,N_14109,N_13532);
nor U14330 (N_14330,N_13769,N_13756);
xor U14331 (N_14331,N_13646,N_14049);
and U14332 (N_14332,N_13658,N_13818);
xor U14333 (N_14333,N_14020,N_13836);
or U14334 (N_14334,N_13522,N_14132);
xor U14335 (N_14335,N_14221,N_13910);
nand U14336 (N_14336,N_13951,N_13939);
nand U14337 (N_14337,N_13944,N_14131);
nand U14338 (N_14338,N_13800,N_14226);
or U14339 (N_14339,N_14036,N_13829);
or U14340 (N_14340,N_13819,N_14238);
nor U14341 (N_14341,N_13825,N_13945);
nor U14342 (N_14342,N_13612,N_13955);
and U14343 (N_14343,N_13613,N_13553);
nor U14344 (N_14344,N_14237,N_13810);
nand U14345 (N_14345,N_13791,N_13654);
nand U14346 (N_14346,N_13863,N_14121);
and U14347 (N_14347,N_14107,N_13797);
nand U14348 (N_14348,N_14225,N_13503);
nor U14349 (N_14349,N_13519,N_13771);
or U14350 (N_14350,N_13834,N_13898);
nor U14351 (N_14351,N_13511,N_13630);
nor U14352 (N_14352,N_13636,N_13566);
nor U14353 (N_14353,N_14081,N_13569);
or U14354 (N_14354,N_13891,N_13915);
or U14355 (N_14355,N_13934,N_13704);
nand U14356 (N_14356,N_13543,N_13606);
and U14357 (N_14357,N_13815,N_14082);
or U14358 (N_14358,N_13973,N_13840);
and U14359 (N_14359,N_13787,N_14074);
nor U14360 (N_14360,N_14210,N_13942);
and U14361 (N_14361,N_13528,N_13887);
nand U14362 (N_14362,N_13782,N_13549);
nand U14363 (N_14363,N_13776,N_13544);
or U14364 (N_14364,N_13678,N_13557);
or U14365 (N_14365,N_13967,N_14161);
and U14366 (N_14366,N_14058,N_13894);
nor U14367 (N_14367,N_14206,N_13546);
nor U14368 (N_14368,N_14050,N_14111);
and U14369 (N_14369,N_13583,N_13947);
nor U14370 (N_14370,N_14175,N_13509);
xor U14371 (N_14371,N_14012,N_13812);
or U14372 (N_14372,N_14028,N_14090);
and U14373 (N_14373,N_13775,N_13670);
nand U14374 (N_14374,N_13765,N_13560);
xnor U14375 (N_14375,N_13846,N_13710);
nand U14376 (N_14376,N_13614,N_13885);
or U14377 (N_14377,N_13661,N_14188);
or U14378 (N_14378,N_14097,N_13932);
nand U14379 (N_14379,N_14189,N_14126);
nand U14380 (N_14380,N_14038,N_14019);
or U14381 (N_14381,N_13869,N_14096);
nand U14382 (N_14382,N_14080,N_13925);
and U14383 (N_14383,N_14101,N_14212);
or U14384 (N_14384,N_14091,N_13982);
nand U14385 (N_14385,N_14194,N_14072);
or U14386 (N_14386,N_14037,N_13620);
xnor U14387 (N_14387,N_14228,N_13609);
or U14388 (N_14388,N_14173,N_14146);
or U14389 (N_14389,N_14133,N_13622);
nand U14390 (N_14390,N_14085,N_13880);
and U14391 (N_14391,N_13652,N_14200);
and U14392 (N_14392,N_13687,N_13708);
and U14393 (N_14393,N_14208,N_13786);
nor U14394 (N_14394,N_13914,N_13843);
or U14395 (N_14395,N_13729,N_13591);
xor U14396 (N_14396,N_13668,N_14152);
nand U14397 (N_14397,N_13627,N_13510);
nand U14398 (N_14398,N_13531,N_13739);
xor U14399 (N_14399,N_13633,N_14135);
nand U14400 (N_14400,N_13584,N_13736);
or U14401 (N_14401,N_13558,N_14148);
xor U14402 (N_14402,N_13607,N_14244);
nor U14403 (N_14403,N_13868,N_13751);
and U14404 (N_14404,N_14073,N_13774);
nor U14405 (N_14405,N_13899,N_13799);
nand U14406 (N_14406,N_13625,N_14116);
nand U14407 (N_14407,N_13517,N_13824);
and U14408 (N_14408,N_13734,N_14129);
nor U14409 (N_14409,N_13851,N_13971);
and U14410 (N_14410,N_13895,N_13961);
or U14411 (N_14411,N_13608,N_13748);
nand U14412 (N_14412,N_13701,N_13615);
and U14413 (N_14413,N_13723,N_13634);
nor U14414 (N_14414,N_13788,N_13850);
and U14415 (N_14415,N_14157,N_13832);
xor U14416 (N_14416,N_13801,N_13696);
nor U14417 (N_14417,N_13624,N_13883);
or U14418 (N_14418,N_13822,N_14108);
nand U14419 (N_14419,N_14106,N_14138);
nand U14420 (N_14420,N_13952,N_13611);
nor U14421 (N_14421,N_13916,N_14071);
and U14422 (N_14422,N_13773,N_13946);
xnor U14423 (N_14423,N_14140,N_13731);
or U14424 (N_14424,N_14167,N_13793);
nor U14425 (N_14425,N_13559,N_13959);
or U14426 (N_14426,N_13699,N_14087);
nor U14427 (N_14427,N_13537,N_14143);
nand U14428 (N_14428,N_13980,N_13994);
or U14429 (N_14429,N_13621,N_13644);
nand U14430 (N_14430,N_13866,N_13763);
xor U14431 (N_14431,N_13764,N_13576);
xor U14432 (N_14432,N_13616,N_13920);
nor U14433 (N_14433,N_14100,N_14223);
nor U14434 (N_14434,N_14197,N_13592);
nor U14435 (N_14435,N_13759,N_14218);
and U14436 (N_14436,N_13903,N_13660);
or U14437 (N_14437,N_13830,N_13556);
and U14438 (N_14438,N_13902,N_13649);
and U14439 (N_14439,N_13969,N_13501);
nor U14440 (N_14440,N_14165,N_13623);
or U14441 (N_14441,N_13524,N_14103);
nand U14442 (N_14442,N_14044,N_14123);
or U14443 (N_14443,N_14006,N_14113);
xnor U14444 (N_14444,N_13857,N_14203);
or U14445 (N_14445,N_14154,N_13727);
and U14446 (N_14446,N_13984,N_13966);
or U14447 (N_14447,N_13940,N_13855);
nand U14448 (N_14448,N_14014,N_14119);
or U14449 (N_14449,N_13823,N_13637);
and U14450 (N_14450,N_14182,N_13849);
or U14451 (N_14451,N_14062,N_14163);
or U14452 (N_14452,N_13629,N_13518);
or U14453 (N_14453,N_14004,N_13602);
and U14454 (N_14454,N_14160,N_13953);
nor U14455 (N_14455,N_13746,N_14130);
and U14456 (N_14456,N_14158,N_13852);
and U14457 (N_14457,N_14117,N_13507);
xnor U14458 (N_14458,N_13725,N_14064);
and U14459 (N_14459,N_14193,N_13972);
and U14460 (N_14460,N_13755,N_13572);
xor U14461 (N_14461,N_13574,N_13567);
nand U14462 (N_14462,N_14086,N_13724);
nor U14463 (N_14463,N_13919,N_13642);
or U14464 (N_14464,N_13963,N_13785);
or U14465 (N_14465,N_14054,N_13534);
xor U14466 (N_14466,N_14147,N_13548);
xnor U14467 (N_14467,N_14166,N_13694);
and U14468 (N_14468,N_14204,N_13842);
or U14469 (N_14469,N_13726,N_13749);
and U14470 (N_14470,N_13536,N_14243);
or U14471 (N_14471,N_13697,N_14190);
and U14472 (N_14472,N_13950,N_13908);
nor U14473 (N_14473,N_13954,N_14222);
or U14474 (N_14474,N_13597,N_13937);
and U14475 (N_14475,N_13712,N_14003);
or U14476 (N_14476,N_13579,N_14015);
nor U14477 (N_14477,N_14178,N_13671);
nand U14478 (N_14478,N_13841,N_13747);
nor U14479 (N_14479,N_13760,N_14030);
or U14480 (N_14480,N_13508,N_13926);
nand U14481 (N_14481,N_14248,N_14042);
and U14482 (N_14482,N_14000,N_14043);
and U14483 (N_14483,N_13999,N_14205);
nor U14484 (N_14484,N_13672,N_14045);
and U14485 (N_14485,N_13828,N_13911);
nand U14486 (N_14486,N_14184,N_13700);
or U14487 (N_14487,N_13744,N_14048);
xnor U14488 (N_14488,N_13979,N_13667);
nor U14489 (N_14489,N_13809,N_13514);
or U14490 (N_14490,N_14149,N_13803);
and U14491 (N_14491,N_13831,N_13655);
or U14492 (N_14492,N_13673,N_13737);
nand U14493 (N_14493,N_13594,N_14220);
or U14494 (N_14494,N_13858,N_13581);
nor U14495 (N_14495,N_13884,N_13990);
nand U14496 (N_14496,N_13674,N_13768);
or U14497 (N_14497,N_14180,N_13873);
and U14498 (N_14498,N_13684,N_13505);
nand U14499 (N_14499,N_13551,N_13938);
nand U14500 (N_14500,N_14034,N_13992);
and U14501 (N_14501,N_13882,N_14235);
or U14502 (N_14502,N_14084,N_13752);
or U14503 (N_14503,N_13588,N_13735);
or U14504 (N_14504,N_13599,N_13590);
nand U14505 (N_14505,N_13648,N_13879);
and U14506 (N_14506,N_13705,N_14227);
and U14507 (N_14507,N_14242,N_14168);
and U14508 (N_14508,N_14011,N_13709);
and U14509 (N_14509,N_14192,N_14122);
and U14510 (N_14510,N_13593,N_14009);
nor U14511 (N_14511,N_13721,N_14039);
nand U14512 (N_14512,N_14155,N_13813);
or U14513 (N_14513,N_14169,N_14001);
nor U14514 (N_14514,N_13643,N_14196);
nor U14515 (N_14515,N_13539,N_13794);
nand U14516 (N_14516,N_14207,N_14245);
and U14517 (N_14517,N_13854,N_14156);
and U14518 (N_14518,N_13745,N_13530);
xnor U14519 (N_14519,N_14040,N_13626);
nor U14520 (N_14520,N_14215,N_13909);
nor U14521 (N_14521,N_14047,N_14056);
nor U14522 (N_14522,N_13582,N_13719);
nand U14523 (N_14523,N_13997,N_13968);
xnor U14524 (N_14524,N_13523,N_13974);
or U14525 (N_14525,N_14217,N_14027);
and U14526 (N_14526,N_13740,N_13783);
or U14527 (N_14527,N_13789,N_13601);
nor U14528 (N_14528,N_13604,N_14124);
and U14529 (N_14529,N_13792,N_13561);
and U14530 (N_14530,N_14059,N_14112);
and U14531 (N_14531,N_13806,N_13502);
and U14532 (N_14532,N_13512,N_13772);
nand U14533 (N_14533,N_13965,N_13811);
nor U14534 (N_14534,N_14115,N_13917);
nor U14535 (N_14535,N_14076,N_13666);
and U14536 (N_14536,N_14053,N_13513);
nor U14537 (N_14537,N_13527,N_14094);
nor U14538 (N_14538,N_13888,N_14067);
nor U14539 (N_14539,N_13573,N_13962);
nor U14540 (N_14540,N_13881,N_13970);
nor U14541 (N_14541,N_13720,N_14032);
xor U14542 (N_14542,N_13568,N_13964);
or U14543 (N_14543,N_13692,N_13665);
or U14544 (N_14544,N_14120,N_13598);
nand U14545 (N_14545,N_13714,N_13686);
or U14546 (N_14546,N_13766,N_14202);
nor U14547 (N_14547,N_13589,N_13798);
nand U14548 (N_14548,N_13779,N_14046);
and U14549 (N_14549,N_13871,N_14099);
nor U14550 (N_14550,N_13878,N_14127);
nor U14551 (N_14551,N_14041,N_13542);
or U14552 (N_14552,N_13927,N_14230);
nand U14553 (N_14553,N_14199,N_13618);
nor U14554 (N_14554,N_14198,N_13603);
or U14555 (N_14555,N_13650,N_13717);
and U14556 (N_14556,N_13901,N_13702);
and U14557 (N_14557,N_13845,N_13535);
nor U14558 (N_14558,N_14065,N_14007);
nor U14559 (N_14559,N_13795,N_14144);
nand U14560 (N_14560,N_13664,N_13682);
nor U14561 (N_14561,N_13635,N_13930);
xnor U14562 (N_14562,N_13922,N_13906);
nor U14563 (N_14563,N_13656,N_13555);
nor U14564 (N_14564,N_13864,N_13816);
and U14565 (N_14565,N_13538,N_13676);
and U14566 (N_14566,N_13960,N_14211);
xnor U14567 (N_14567,N_13500,N_13837);
nand U14568 (N_14568,N_13987,N_13993);
nor U14569 (N_14569,N_14118,N_13681);
nand U14570 (N_14570,N_13826,N_13750);
or U14571 (N_14571,N_13587,N_14136);
and U14572 (N_14572,N_13578,N_14092);
and U14573 (N_14573,N_13571,N_13802);
nor U14574 (N_14574,N_13905,N_14172);
nor U14575 (N_14575,N_13533,N_13913);
nand U14576 (N_14576,N_14066,N_13693);
and U14577 (N_14577,N_14249,N_13784);
or U14578 (N_14578,N_14224,N_13867);
nand U14579 (N_14579,N_14026,N_14164);
nor U14580 (N_14580,N_14170,N_13931);
nand U14581 (N_14581,N_13762,N_14142);
nor U14582 (N_14582,N_13853,N_14137);
or U14583 (N_14583,N_13808,N_14134);
xor U14584 (N_14584,N_13986,N_14104);
nand U14585 (N_14585,N_14183,N_13956);
nor U14586 (N_14586,N_14241,N_13679);
xor U14587 (N_14587,N_13790,N_13685);
and U14588 (N_14588,N_14171,N_14105);
or U14589 (N_14589,N_13521,N_13659);
and U14590 (N_14590,N_13989,N_14213);
nor U14591 (N_14591,N_13540,N_14128);
and U14592 (N_14592,N_13529,N_13923);
or U14593 (N_14593,N_14068,N_13631);
and U14594 (N_14594,N_13639,N_14151);
or U14595 (N_14595,N_13995,N_14089);
or U14596 (N_14596,N_13859,N_13861);
nand U14597 (N_14597,N_13870,N_13948);
nor U14598 (N_14598,N_13680,N_13743);
nand U14599 (N_14599,N_14079,N_13839);
nor U14600 (N_14600,N_14214,N_13893);
and U14601 (N_14601,N_13941,N_13943);
or U14602 (N_14602,N_13641,N_13632);
and U14603 (N_14603,N_13677,N_14174);
xor U14604 (N_14604,N_13565,N_13900);
and U14605 (N_14605,N_13596,N_14010);
xnor U14606 (N_14606,N_13504,N_14057);
or U14607 (N_14607,N_14125,N_13820);
or U14608 (N_14608,N_14021,N_13865);
nand U14609 (N_14609,N_13730,N_13706);
or U14610 (N_14610,N_14016,N_13835);
nand U14611 (N_14611,N_13833,N_13733);
and U14612 (N_14612,N_13728,N_13804);
or U14613 (N_14613,N_13827,N_13975);
and U14614 (N_14614,N_14024,N_13921);
nand U14615 (N_14615,N_13935,N_14153);
and U14616 (N_14616,N_14216,N_14141);
and U14617 (N_14617,N_13904,N_14229);
or U14618 (N_14618,N_14013,N_13610);
or U14619 (N_14619,N_13506,N_13777);
and U14620 (N_14620,N_13796,N_14191);
or U14621 (N_14621,N_14033,N_14008);
and U14622 (N_14622,N_13912,N_14145);
nand U14623 (N_14623,N_14233,N_13848);
nor U14624 (N_14624,N_14162,N_13918);
or U14625 (N_14625,N_14232,N_13765);
or U14626 (N_14626,N_13510,N_13554);
and U14627 (N_14627,N_14148,N_13780);
or U14628 (N_14628,N_14233,N_14054);
and U14629 (N_14629,N_13793,N_13505);
nor U14630 (N_14630,N_13824,N_14157);
or U14631 (N_14631,N_14074,N_13505);
nor U14632 (N_14632,N_13967,N_13515);
or U14633 (N_14633,N_13906,N_14198);
and U14634 (N_14634,N_13917,N_13688);
nand U14635 (N_14635,N_13640,N_13836);
or U14636 (N_14636,N_13839,N_13725);
or U14637 (N_14637,N_14139,N_13841);
and U14638 (N_14638,N_14136,N_13907);
or U14639 (N_14639,N_13714,N_13836);
nor U14640 (N_14640,N_14247,N_13681);
xor U14641 (N_14641,N_14212,N_14037);
nor U14642 (N_14642,N_13929,N_14062);
and U14643 (N_14643,N_13672,N_13872);
and U14644 (N_14644,N_14178,N_13553);
xnor U14645 (N_14645,N_13516,N_13562);
xnor U14646 (N_14646,N_13686,N_13991);
or U14647 (N_14647,N_14043,N_13934);
nor U14648 (N_14648,N_14097,N_13939);
or U14649 (N_14649,N_13831,N_14034);
nand U14650 (N_14650,N_13915,N_13587);
and U14651 (N_14651,N_13799,N_13939);
and U14652 (N_14652,N_13877,N_13640);
nor U14653 (N_14653,N_14059,N_14180);
or U14654 (N_14654,N_14000,N_14026);
and U14655 (N_14655,N_13991,N_13722);
or U14656 (N_14656,N_14214,N_14152);
nand U14657 (N_14657,N_13516,N_13587);
or U14658 (N_14658,N_13754,N_13955);
xnor U14659 (N_14659,N_14092,N_13733);
xor U14660 (N_14660,N_13719,N_14035);
and U14661 (N_14661,N_13546,N_13779);
nor U14662 (N_14662,N_14172,N_13958);
xnor U14663 (N_14663,N_13503,N_13879);
nand U14664 (N_14664,N_13893,N_13770);
or U14665 (N_14665,N_14140,N_13996);
or U14666 (N_14666,N_13804,N_13873);
nor U14667 (N_14667,N_14059,N_14073);
or U14668 (N_14668,N_13513,N_14044);
xor U14669 (N_14669,N_13799,N_13763);
and U14670 (N_14670,N_13730,N_14212);
nand U14671 (N_14671,N_14062,N_14229);
nor U14672 (N_14672,N_14026,N_13546);
nor U14673 (N_14673,N_14002,N_13507);
or U14674 (N_14674,N_14089,N_13926);
and U14675 (N_14675,N_13951,N_14107);
and U14676 (N_14676,N_14169,N_14010);
nand U14677 (N_14677,N_13668,N_14242);
nor U14678 (N_14678,N_13623,N_14172);
nor U14679 (N_14679,N_13521,N_13562);
xor U14680 (N_14680,N_14055,N_13876);
and U14681 (N_14681,N_13841,N_13561);
nor U14682 (N_14682,N_13888,N_13616);
and U14683 (N_14683,N_14051,N_14223);
nor U14684 (N_14684,N_14054,N_13943);
xnor U14685 (N_14685,N_13624,N_13821);
or U14686 (N_14686,N_13910,N_14034);
nor U14687 (N_14687,N_14131,N_13812);
or U14688 (N_14688,N_13744,N_13607);
xnor U14689 (N_14689,N_14069,N_13689);
nor U14690 (N_14690,N_13767,N_14109);
nand U14691 (N_14691,N_13854,N_14095);
xnor U14692 (N_14692,N_13549,N_13882);
nand U14693 (N_14693,N_14026,N_13839);
nand U14694 (N_14694,N_14140,N_13861);
nor U14695 (N_14695,N_13624,N_13760);
xnor U14696 (N_14696,N_13737,N_14105);
nand U14697 (N_14697,N_14151,N_14023);
nand U14698 (N_14698,N_14184,N_14140);
nor U14699 (N_14699,N_13841,N_13718);
nand U14700 (N_14700,N_14061,N_13604);
nor U14701 (N_14701,N_13957,N_13825);
or U14702 (N_14702,N_13547,N_13572);
nor U14703 (N_14703,N_13951,N_14106);
nand U14704 (N_14704,N_13931,N_14109);
nand U14705 (N_14705,N_14120,N_14085);
nor U14706 (N_14706,N_13770,N_13844);
xor U14707 (N_14707,N_13910,N_13750);
or U14708 (N_14708,N_13706,N_14185);
and U14709 (N_14709,N_13563,N_14152);
nand U14710 (N_14710,N_13524,N_14082);
nor U14711 (N_14711,N_14141,N_13918);
nand U14712 (N_14712,N_14002,N_13590);
nand U14713 (N_14713,N_14247,N_13532);
or U14714 (N_14714,N_13736,N_14076);
xnor U14715 (N_14715,N_13561,N_13922);
nor U14716 (N_14716,N_13589,N_13544);
and U14717 (N_14717,N_13532,N_13905);
nand U14718 (N_14718,N_13623,N_14232);
and U14719 (N_14719,N_13994,N_13748);
and U14720 (N_14720,N_14124,N_13806);
xor U14721 (N_14721,N_14123,N_13768);
or U14722 (N_14722,N_13999,N_13663);
nand U14723 (N_14723,N_14054,N_13780);
and U14724 (N_14724,N_13635,N_13600);
nor U14725 (N_14725,N_13747,N_14087);
nor U14726 (N_14726,N_13594,N_13795);
nand U14727 (N_14727,N_13516,N_14082);
and U14728 (N_14728,N_13918,N_14124);
nor U14729 (N_14729,N_14111,N_13944);
nand U14730 (N_14730,N_14118,N_13832);
nand U14731 (N_14731,N_14221,N_13669);
nor U14732 (N_14732,N_14189,N_14083);
nor U14733 (N_14733,N_13622,N_13968);
or U14734 (N_14734,N_13787,N_14009);
or U14735 (N_14735,N_13622,N_13730);
and U14736 (N_14736,N_13897,N_14159);
xnor U14737 (N_14737,N_13511,N_14155);
xnor U14738 (N_14738,N_13949,N_14015);
or U14739 (N_14739,N_14189,N_13960);
nor U14740 (N_14740,N_13670,N_13820);
and U14741 (N_14741,N_13964,N_13731);
or U14742 (N_14742,N_13860,N_13646);
or U14743 (N_14743,N_14059,N_13949);
nor U14744 (N_14744,N_13798,N_13636);
or U14745 (N_14745,N_14137,N_13789);
or U14746 (N_14746,N_13591,N_13857);
nand U14747 (N_14747,N_13587,N_13973);
and U14748 (N_14748,N_13834,N_14070);
nand U14749 (N_14749,N_14236,N_14102);
or U14750 (N_14750,N_14227,N_13849);
or U14751 (N_14751,N_13510,N_13658);
or U14752 (N_14752,N_13802,N_14062);
or U14753 (N_14753,N_14102,N_14097);
nor U14754 (N_14754,N_13748,N_14184);
nand U14755 (N_14755,N_13579,N_13709);
and U14756 (N_14756,N_13732,N_13801);
or U14757 (N_14757,N_13698,N_13538);
nor U14758 (N_14758,N_13993,N_13703);
nand U14759 (N_14759,N_13913,N_14147);
nor U14760 (N_14760,N_13601,N_13859);
and U14761 (N_14761,N_13727,N_14104);
nand U14762 (N_14762,N_13683,N_13626);
nor U14763 (N_14763,N_14044,N_13551);
nand U14764 (N_14764,N_14226,N_13644);
and U14765 (N_14765,N_14202,N_13732);
or U14766 (N_14766,N_13757,N_13824);
xnor U14767 (N_14767,N_13525,N_14153);
or U14768 (N_14768,N_14142,N_13711);
nor U14769 (N_14769,N_13909,N_13712);
and U14770 (N_14770,N_13912,N_13798);
or U14771 (N_14771,N_14194,N_14124);
xnor U14772 (N_14772,N_13964,N_14128);
nand U14773 (N_14773,N_14083,N_14159);
and U14774 (N_14774,N_14138,N_13958);
nor U14775 (N_14775,N_13562,N_13830);
or U14776 (N_14776,N_13709,N_13799);
and U14777 (N_14777,N_14136,N_13965);
xor U14778 (N_14778,N_13964,N_13630);
xnor U14779 (N_14779,N_14110,N_13549);
or U14780 (N_14780,N_14028,N_13513);
xnor U14781 (N_14781,N_13574,N_13865);
and U14782 (N_14782,N_13648,N_13972);
nor U14783 (N_14783,N_13819,N_14188);
nand U14784 (N_14784,N_14197,N_14066);
nor U14785 (N_14785,N_13841,N_13706);
or U14786 (N_14786,N_14145,N_14146);
and U14787 (N_14787,N_13999,N_14158);
nand U14788 (N_14788,N_13585,N_14029);
or U14789 (N_14789,N_13541,N_14089);
nor U14790 (N_14790,N_13943,N_13725);
and U14791 (N_14791,N_13878,N_14097);
or U14792 (N_14792,N_14219,N_13511);
and U14793 (N_14793,N_14174,N_14166);
xnor U14794 (N_14794,N_13845,N_13766);
and U14795 (N_14795,N_13977,N_13625);
or U14796 (N_14796,N_13849,N_13803);
nand U14797 (N_14797,N_13691,N_13746);
and U14798 (N_14798,N_13832,N_14068);
nor U14799 (N_14799,N_13743,N_13541);
nor U14800 (N_14800,N_14114,N_13978);
or U14801 (N_14801,N_14214,N_14127);
xnor U14802 (N_14802,N_13618,N_13664);
or U14803 (N_14803,N_14160,N_13934);
and U14804 (N_14804,N_13987,N_14192);
nand U14805 (N_14805,N_13584,N_13519);
nand U14806 (N_14806,N_13688,N_14047);
or U14807 (N_14807,N_13780,N_13765);
or U14808 (N_14808,N_13862,N_13935);
nand U14809 (N_14809,N_14233,N_14078);
xnor U14810 (N_14810,N_14145,N_13633);
and U14811 (N_14811,N_13789,N_13991);
and U14812 (N_14812,N_14124,N_14074);
nand U14813 (N_14813,N_13559,N_13900);
or U14814 (N_14814,N_14141,N_14061);
and U14815 (N_14815,N_14046,N_14192);
or U14816 (N_14816,N_13908,N_14101);
and U14817 (N_14817,N_13640,N_14036);
or U14818 (N_14818,N_13570,N_14236);
nand U14819 (N_14819,N_13627,N_13762);
nor U14820 (N_14820,N_13580,N_13679);
xnor U14821 (N_14821,N_14155,N_13540);
nor U14822 (N_14822,N_13991,N_13842);
or U14823 (N_14823,N_13721,N_13896);
or U14824 (N_14824,N_13671,N_14218);
or U14825 (N_14825,N_13976,N_13545);
nand U14826 (N_14826,N_13567,N_13965);
nand U14827 (N_14827,N_13856,N_13775);
and U14828 (N_14828,N_13627,N_14140);
nand U14829 (N_14829,N_13861,N_13993);
nand U14830 (N_14830,N_13601,N_14172);
nor U14831 (N_14831,N_13775,N_13628);
xor U14832 (N_14832,N_13553,N_13713);
xor U14833 (N_14833,N_13623,N_14238);
and U14834 (N_14834,N_13891,N_13764);
and U14835 (N_14835,N_13606,N_14110);
nand U14836 (N_14836,N_13932,N_14002);
nor U14837 (N_14837,N_13577,N_13850);
or U14838 (N_14838,N_14167,N_13870);
and U14839 (N_14839,N_13993,N_13948);
or U14840 (N_14840,N_13781,N_13646);
nor U14841 (N_14841,N_13662,N_13949);
or U14842 (N_14842,N_13556,N_14086);
nor U14843 (N_14843,N_13755,N_13650);
xor U14844 (N_14844,N_13911,N_14190);
and U14845 (N_14845,N_13958,N_13998);
and U14846 (N_14846,N_13865,N_13632);
and U14847 (N_14847,N_13521,N_13993);
and U14848 (N_14848,N_13536,N_13790);
or U14849 (N_14849,N_14248,N_14118);
or U14850 (N_14850,N_13793,N_13854);
and U14851 (N_14851,N_13546,N_13690);
xor U14852 (N_14852,N_13738,N_13974);
or U14853 (N_14853,N_13830,N_14098);
or U14854 (N_14854,N_13796,N_13595);
xor U14855 (N_14855,N_13868,N_13836);
and U14856 (N_14856,N_13738,N_13917);
nor U14857 (N_14857,N_13716,N_13908);
xor U14858 (N_14858,N_14083,N_13919);
or U14859 (N_14859,N_13836,N_14207);
and U14860 (N_14860,N_14205,N_14115);
and U14861 (N_14861,N_14243,N_14159);
and U14862 (N_14862,N_13531,N_14229);
nand U14863 (N_14863,N_13896,N_13984);
and U14864 (N_14864,N_13514,N_13980);
nand U14865 (N_14865,N_13598,N_14061);
nand U14866 (N_14866,N_13765,N_13743);
xor U14867 (N_14867,N_13831,N_14086);
nand U14868 (N_14868,N_13624,N_13673);
nand U14869 (N_14869,N_13883,N_14005);
nand U14870 (N_14870,N_13669,N_13561);
or U14871 (N_14871,N_14055,N_13868);
nand U14872 (N_14872,N_13888,N_13726);
nand U14873 (N_14873,N_13650,N_14110);
and U14874 (N_14874,N_13692,N_13827);
and U14875 (N_14875,N_13706,N_14189);
and U14876 (N_14876,N_13914,N_13909);
nor U14877 (N_14877,N_13717,N_14248);
and U14878 (N_14878,N_13774,N_13988);
nor U14879 (N_14879,N_14036,N_13527);
or U14880 (N_14880,N_13836,N_13826);
or U14881 (N_14881,N_13814,N_14207);
or U14882 (N_14882,N_13827,N_13889);
or U14883 (N_14883,N_14225,N_14024);
nor U14884 (N_14884,N_13890,N_14074);
nor U14885 (N_14885,N_14206,N_13821);
nand U14886 (N_14886,N_14132,N_14163);
or U14887 (N_14887,N_14112,N_13763);
and U14888 (N_14888,N_14154,N_13776);
or U14889 (N_14889,N_13934,N_14190);
nor U14890 (N_14890,N_13955,N_13984);
and U14891 (N_14891,N_13937,N_13714);
or U14892 (N_14892,N_14135,N_14125);
and U14893 (N_14893,N_14006,N_13880);
nor U14894 (N_14894,N_14233,N_13804);
nand U14895 (N_14895,N_13517,N_13631);
or U14896 (N_14896,N_13518,N_14185);
and U14897 (N_14897,N_13848,N_13974);
xor U14898 (N_14898,N_14100,N_14040);
or U14899 (N_14899,N_13832,N_14076);
nor U14900 (N_14900,N_13612,N_13739);
nor U14901 (N_14901,N_13604,N_14064);
and U14902 (N_14902,N_13902,N_13702);
xor U14903 (N_14903,N_13946,N_13790);
and U14904 (N_14904,N_14171,N_14019);
or U14905 (N_14905,N_14204,N_13658);
and U14906 (N_14906,N_13610,N_13573);
nand U14907 (N_14907,N_14169,N_13782);
nor U14908 (N_14908,N_13868,N_13846);
and U14909 (N_14909,N_13696,N_13948);
or U14910 (N_14910,N_13648,N_14223);
xnor U14911 (N_14911,N_13590,N_13760);
and U14912 (N_14912,N_14161,N_13872);
or U14913 (N_14913,N_13523,N_13893);
and U14914 (N_14914,N_13888,N_14123);
and U14915 (N_14915,N_14113,N_14020);
nand U14916 (N_14916,N_14228,N_13548);
nand U14917 (N_14917,N_14047,N_13858);
nor U14918 (N_14918,N_13605,N_13808);
xor U14919 (N_14919,N_13515,N_13500);
or U14920 (N_14920,N_13616,N_13705);
or U14921 (N_14921,N_14030,N_14081);
or U14922 (N_14922,N_13642,N_13807);
nor U14923 (N_14923,N_13703,N_13675);
or U14924 (N_14924,N_13726,N_13915);
or U14925 (N_14925,N_13570,N_13757);
and U14926 (N_14926,N_13617,N_13673);
nor U14927 (N_14927,N_14182,N_14158);
and U14928 (N_14928,N_14108,N_13837);
nand U14929 (N_14929,N_13663,N_13895);
nor U14930 (N_14930,N_13741,N_13542);
or U14931 (N_14931,N_13887,N_13612);
or U14932 (N_14932,N_13832,N_13663);
nand U14933 (N_14933,N_13636,N_13725);
xor U14934 (N_14934,N_13989,N_13554);
nor U14935 (N_14935,N_14204,N_13805);
nor U14936 (N_14936,N_14034,N_13908);
nor U14937 (N_14937,N_14077,N_13600);
nand U14938 (N_14938,N_13895,N_13686);
nor U14939 (N_14939,N_14021,N_13886);
and U14940 (N_14940,N_14010,N_13591);
nand U14941 (N_14941,N_13617,N_13949);
and U14942 (N_14942,N_13575,N_13963);
or U14943 (N_14943,N_13594,N_13729);
nand U14944 (N_14944,N_13757,N_13731);
or U14945 (N_14945,N_14074,N_14064);
xor U14946 (N_14946,N_14249,N_13992);
and U14947 (N_14947,N_13965,N_13846);
nor U14948 (N_14948,N_13636,N_13835);
nor U14949 (N_14949,N_13598,N_14128);
or U14950 (N_14950,N_13602,N_14084);
nor U14951 (N_14951,N_13970,N_14115);
nor U14952 (N_14952,N_13787,N_13644);
nor U14953 (N_14953,N_13788,N_14063);
or U14954 (N_14954,N_13743,N_14104);
or U14955 (N_14955,N_13903,N_13511);
nor U14956 (N_14956,N_13880,N_13956);
and U14957 (N_14957,N_14165,N_14192);
and U14958 (N_14958,N_13701,N_13538);
or U14959 (N_14959,N_14196,N_13608);
nand U14960 (N_14960,N_13702,N_13804);
nor U14961 (N_14961,N_13972,N_13525);
and U14962 (N_14962,N_13632,N_14092);
nand U14963 (N_14963,N_13688,N_14148);
nand U14964 (N_14964,N_13621,N_14033);
nand U14965 (N_14965,N_13893,N_13710);
nor U14966 (N_14966,N_13812,N_13736);
and U14967 (N_14967,N_13583,N_13978);
nor U14968 (N_14968,N_13577,N_13567);
nor U14969 (N_14969,N_13587,N_14076);
and U14970 (N_14970,N_13689,N_13707);
nor U14971 (N_14971,N_14173,N_13536);
nor U14972 (N_14972,N_13682,N_13948);
nor U14973 (N_14973,N_13588,N_13965);
nand U14974 (N_14974,N_13706,N_14241);
or U14975 (N_14975,N_14146,N_13927);
nor U14976 (N_14976,N_13839,N_13510);
or U14977 (N_14977,N_14097,N_14047);
nand U14978 (N_14978,N_13855,N_14165);
or U14979 (N_14979,N_14214,N_14227);
nor U14980 (N_14980,N_14118,N_14236);
xor U14981 (N_14981,N_13914,N_13707);
and U14982 (N_14982,N_14050,N_14136);
nor U14983 (N_14983,N_14086,N_13590);
nor U14984 (N_14984,N_13998,N_14029);
and U14985 (N_14985,N_13535,N_14193);
nand U14986 (N_14986,N_13796,N_13970);
xnor U14987 (N_14987,N_13907,N_13712);
or U14988 (N_14988,N_13970,N_13839);
nand U14989 (N_14989,N_13674,N_13684);
or U14990 (N_14990,N_13746,N_14014);
nand U14991 (N_14991,N_13927,N_13615);
and U14992 (N_14992,N_13528,N_13756);
nand U14993 (N_14993,N_13683,N_13717);
nand U14994 (N_14994,N_14116,N_14104);
and U14995 (N_14995,N_13810,N_14071);
nand U14996 (N_14996,N_13594,N_13585);
nor U14997 (N_14997,N_13559,N_14226);
or U14998 (N_14998,N_13814,N_13550);
or U14999 (N_14999,N_13746,N_14230);
nand UO_0 (O_0,N_14631,N_14708);
or UO_1 (O_1,N_14567,N_14494);
nand UO_2 (O_2,N_14646,N_14390);
nor UO_3 (O_3,N_14421,N_14408);
and UO_4 (O_4,N_14310,N_14900);
and UO_5 (O_5,N_14859,N_14937);
nor UO_6 (O_6,N_14958,N_14824);
nor UO_7 (O_7,N_14802,N_14771);
or UO_8 (O_8,N_14395,N_14487);
or UO_9 (O_9,N_14531,N_14645);
and UO_10 (O_10,N_14478,N_14878);
nand UO_11 (O_11,N_14558,N_14890);
and UO_12 (O_12,N_14983,N_14412);
or UO_13 (O_13,N_14587,N_14629);
nand UO_14 (O_14,N_14852,N_14435);
or UO_15 (O_15,N_14268,N_14843);
and UO_16 (O_16,N_14911,N_14807);
nor UO_17 (O_17,N_14944,N_14840);
and UO_18 (O_18,N_14952,N_14823);
nand UO_19 (O_19,N_14875,N_14790);
xor UO_20 (O_20,N_14598,N_14376);
nand UO_21 (O_21,N_14861,N_14902);
nor UO_22 (O_22,N_14438,N_14489);
xnor UO_23 (O_23,N_14672,N_14725);
and UO_24 (O_24,N_14447,N_14656);
nand UO_25 (O_25,N_14520,N_14806);
nand UO_26 (O_26,N_14626,N_14251);
xnor UO_27 (O_27,N_14668,N_14568);
nor UO_28 (O_28,N_14787,N_14681);
or UO_29 (O_29,N_14354,N_14866);
nand UO_30 (O_30,N_14292,N_14868);
and UO_31 (O_31,N_14924,N_14510);
and UO_32 (O_32,N_14953,N_14382);
and UO_33 (O_33,N_14456,N_14273);
or UO_34 (O_34,N_14916,N_14550);
nand UO_35 (O_35,N_14355,N_14608);
nand UO_36 (O_36,N_14921,N_14719);
and UO_37 (O_37,N_14315,N_14663);
or UO_38 (O_38,N_14403,N_14709);
nand UO_39 (O_39,N_14640,N_14563);
nand UO_40 (O_40,N_14285,N_14400);
nor UO_41 (O_41,N_14420,N_14695);
and UO_42 (O_42,N_14280,N_14387);
nor UO_43 (O_43,N_14737,N_14455);
and UO_44 (O_44,N_14989,N_14665);
nand UO_45 (O_45,N_14814,N_14688);
and UO_46 (O_46,N_14381,N_14618);
or UO_47 (O_47,N_14407,N_14961);
nand UO_48 (O_48,N_14459,N_14939);
nor UO_49 (O_49,N_14954,N_14877);
nor UO_50 (O_50,N_14615,N_14661);
and UO_51 (O_51,N_14516,N_14848);
or UO_52 (O_52,N_14312,N_14886);
xnor UO_53 (O_53,N_14345,N_14811);
or UO_54 (O_54,N_14850,N_14847);
and UO_55 (O_55,N_14366,N_14915);
xnor UO_56 (O_56,N_14658,N_14323);
and UO_57 (O_57,N_14981,N_14832);
nand UO_58 (O_58,N_14610,N_14584);
nand UO_59 (O_59,N_14577,N_14579);
xnor UO_60 (O_60,N_14503,N_14572);
nand UO_61 (O_61,N_14263,N_14675);
and UO_62 (O_62,N_14296,N_14769);
or UO_63 (O_63,N_14519,N_14842);
or UO_64 (O_64,N_14545,N_14255);
nand UO_65 (O_65,N_14976,N_14942);
nand UO_66 (O_66,N_14554,N_14405);
nand UO_67 (O_67,N_14964,N_14705);
nand UO_68 (O_68,N_14731,N_14909);
xnor UO_69 (O_69,N_14333,N_14397);
or UO_70 (O_70,N_14763,N_14884);
xor UO_71 (O_71,N_14517,N_14473);
or UO_72 (O_72,N_14349,N_14882);
nand UO_73 (O_73,N_14896,N_14327);
nand UO_74 (O_74,N_14913,N_14370);
nor UO_75 (O_75,N_14756,N_14690);
and UO_76 (O_76,N_14547,N_14476);
or UO_77 (O_77,N_14858,N_14367);
nand UO_78 (O_78,N_14325,N_14458);
and UO_79 (O_79,N_14962,N_14860);
or UO_80 (O_80,N_14997,N_14335);
nor UO_81 (O_81,N_14600,N_14922);
nor UO_82 (O_82,N_14780,N_14261);
nand UO_83 (O_83,N_14299,N_14301);
and UO_84 (O_84,N_14839,N_14704);
nand UO_85 (O_85,N_14630,N_14761);
or UO_86 (O_86,N_14256,N_14999);
and UO_87 (O_87,N_14609,N_14934);
nor UO_88 (O_88,N_14712,N_14309);
or UO_89 (O_89,N_14393,N_14791);
nor UO_90 (O_90,N_14298,N_14541);
or UO_91 (O_91,N_14744,N_14794);
nand UO_92 (O_92,N_14796,N_14970);
nor UO_93 (O_93,N_14360,N_14887);
xor UO_94 (O_94,N_14506,N_14923);
or UO_95 (O_95,N_14497,N_14339);
xor UO_96 (O_96,N_14904,N_14523);
or UO_97 (O_97,N_14930,N_14835);
nor UO_98 (O_98,N_14437,N_14827);
nor UO_99 (O_99,N_14689,N_14912);
nor UO_100 (O_100,N_14592,N_14575);
nor UO_101 (O_101,N_14966,N_14557);
nand UO_102 (O_102,N_14965,N_14485);
nor UO_103 (O_103,N_14736,N_14528);
xnor UO_104 (O_104,N_14957,N_14371);
nand UO_105 (O_105,N_14760,N_14926);
nand UO_106 (O_106,N_14936,N_14805);
nand UO_107 (O_107,N_14644,N_14483);
and UO_108 (O_108,N_14929,N_14594);
or UO_109 (O_109,N_14578,N_14873);
nand UO_110 (O_110,N_14809,N_14803);
or UO_111 (O_111,N_14318,N_14469);
nor UO_112 (O_112,N_14996,N_14450);
nor UO_113 (O_113,N_14259,N_14735);
nor UO_114 (O_114,N_14286,N_14767);
or UO_115 (O_115,N_14717,N_14582);
or UO_116 (O_116,N_14559,N_14826);
nand UO_117 (O_117,N_14862,N_14306);
xor UO_118 (O_118,N_14490,N_14738);
and UO_119 (O_119,N_14816,N_14642);
xor UO_120 (O_120,N_14625,N_14785);
and UO_121 (O_121,N_14655,N_14951);
and UO_122 (O_122,N_14270,N_14752);
nand UO_123 (O_123,N_14604,N_14423);
or UO_124 (O_124,N_14694,N_14938);
xnor UO_125 (O_125,N_14893,N_14632);
xor UO_126 (O_126,N_14978,N_14932);
xnor UO_127 (O_127,N_14566,N_14253);
nand UO_128 (O_128,N_14508,N_14369);
or UO_129 (O_129,N_14838,N_14673);
and UO_130 (O_130,N_14727,N_14649);
and UO_131 (O_131,N_14368,N_14386);
or UO_132 (O_132,N_14331,N_14856);
xor UO_133 (O_133,N_14328,N_14880);
nand UO_134 (O_134,N_14730,N_14553);
nor UO_135 (O_135,N_14274,N_14676);
xor UO_136 (O_136,N_14617,N_14419);
and UO_137 (O_137,N_14334,N_14549);
nor UO_138 (O_138,N_14363,N_14430);
nor UO_139 (O_139,N_14666,N_14425);
nand UO_140 (O_140,N_14889,N_14963);
nand UO_141 (O_141,N_14741,N_14431);
xnor UO_142 (O_142,N_14596,N_14851);
nand UO_143 (O_143,N_14797,N_14278);
nor UO_144 (O_144,N_14313,N_14406);
or UO_145 (O_145,N_14518,N_14910);
or UO_146 (O_146,N_14987,N_14466);
and UO_147 (O_147,N_14602,N_14303);
nand UO_148 (O_148,N_14792,N_14611);
nand UO_149 (O_149,N_14511,N_14664);
and UO_150 (O_150,N_14949,N_14603);
and UO_151 (O_151,N_14500,N_14831);
nor UO_152 (O_152,N_14317,N_14484);
and UO_153 (O_153,N_14678,N_14828);
or UO_154 (O_154,N_14975,N_14452);
nor UO_155 (O_155,N_14982,N_14540);
nand UO_156 (O_156,N_14322,N_14260);
and UO_157 (O_157,N_14765,N_14380);
or UO_158 (O_158,N_14706,N_14992);
nor UO_159 (O_159,N_14679,N_14434);
xnor UO_160 (O_160,N_14591,N_14994);
or UO_161 (O_161,N_14925,N_14496);
nand UO_162 (O_162,N_14837,N_14340);
nor UO_163 (O_163,N_14973,N_14683);
and UO_164 (O_164,N_14956,N_14977);
and UO_165 (O_165,N_14534,N_14304);
nor UO_166 (O_166,N_14290,N_14544);
or UO_167 (O_167,N_14674,N_14470);
nor UO_168 (O_168,N_14398,N_14457);
nor UO_169 (O_169,N_14394,N_14513);
or UO_170 (O_170,N_14462,N_14362);
or UO_171 (O_171,N_14635,N_14696);
nand UO_172 (O_172,N_14894,N_14819);
nand UO_173 (O_173,N_14772,N_14379);
nand UO_174 (O_174,N_14556,N_14501);
nor UO_175 (O_175,N_14507,N_14855);
or UO_176 (O_176,N_14372,N_14723);
or UO_177 (O_177,N_14770,N_14433);
or UO_178 (O_178,N_14897,N_14871);
xnor UO_179 (O_179,N_14745,N_14801);
and UO_180 (O_180,N_14492,N_14264);
xor UO_181 (O_181,N_14337,N_14959);
xnor UO_182 (O_182,N_14650,N_14338);
and UO_183 (O_183,N_14417,N_14758);
or UO_184 (O_184,N_14754,N_14378);
nand UO_185 (O_185,N_14968,N_14291);
nor UO_186 (O_186,N_14906,N_14931);
nor UO_187 (O_187,N_14616,N_14332);
nor UO_188 (O_188,N_14853,N_14308);
nor UO_189 (O_189,N_14491,N_14316);
or UO_190 (O_190,N_14588,N_14766);
or UO_191 (O_191,N_14972,N_14388);
and UO_192 (O_192,N_14895,N_14542);
and UO_193 (O_193,N_14746,N_14401);
and UO_194 (O_194,N_14637,N_14687);
xor UO_195 (O_195,N_14812,N_14933);
or UO_196 (O_196,N_14277,N_14391);
nor UO_197 (O_197,N_14980,N_14524);
xor UO_198 (O_198,N_14585,N_14947);
nand UO_199 (O_199,N_14446,N_14879);
nor UO_200 (O_200,N_14562,N_14699);
nor UO_201 (O_201,N_14702,N_14724);
nand UO_202 (O_202,N_14597,N_14351);
or UO_203 (O_203,N_14498,N_14636);
nor UO_204 (O_204,N_14624,N_14950);
nand UO_205 (O_205,N_14798,N_14595);
or UO_206 (O_206,N_14899,N_14872);
xnor UO_207 (O_207,N_14427,N_14782);
nand UO_208 (O_208,N_14905,N_14825);
xnor UO_209 (O_209,N_14716,N_14747);
or UO_210 (O_210,N_14935,N_14991);
nand UO_211 (O_211,N_14440,N_14444);
nor UO_212 (O_212,N_14845,N_14729);
nor UO_213 (O_213,N_14634,N_14776);
nor UO_214 (O_214,N_14365,N_14821);
and UO_215 (O_215,N_14710,N_14495);
nor UO_216 (O_216,N_14414,N_14888);
nand UO_217 (O_217,N_14881,N_14844);
nand UO_218 (O_218,N_14829,N_14804);
xnor UO_219 (O_219,N_14948,N_14432);
and UO_220 (O_220,N_14529,N_14521);
nand UO_221 (O_221,N_14527,N_14775);
nor UO_222 (O_222,N_14443,N_14293);
or UO_223 (O_223,N_14289,N_14472);
and UO_224 (O_224,N_14721,N_14336);
xnor UO_225 (O_225,N_14620,N_14530);
nand UO_226 (O_226,N_14750,N_14539);
nand UO_227 (O_227,N_14903,N_14413);
and UO_228 (O_228,N_14841,N_14422);
xnor UO_229 (O_229,N_14300,N_14555);
and UO_230 (O_230,N_14751,N_14789);
and UO_231 (O_231,N_14522,N_14686);
nor UO_232 (O_232,N_14918,N_14633);
and UO_233 (O_233,N_14471,N_14343);
nand UO_234 (O_234,N_14898,N_14374);
and UO_235 (O_235,N_14734,N_14416);
nor UO_236 (O_236,N_14670,N_14757);
or UO_237 (O_237,N_14580,N_14783);
or UO_238 (O_238,N_14396,N_14377);
and UO_239 (O_239,N_14574,N_14786);
nor UO_240 (O_240,N_14605,N_14593);
xor UO_241 (O_241,N_14799,N_14565);
or UO_242 (O_242,N_14319,N_14353);
nand UO_243 (O_243,N_14307,N_14891);
xor UO_244 (O_244,N_14774,N_14822);
xnor UO_245 (O_245,N_14691,N_14448);
xor UO_246 (O_246,N_14548,N_14287);
or UO_247 (O_247,N_14623,N_14711);
nor UO_248 (O_248,N_14692,N_14984);
nand UO_249 (O_249,N_14262,N_14945);
nand UO_250 (O_250,N_14546,N_14955);
and UO_251 (O_251,N_14614,N_14643);
or UO_252 (O_252,N_14795,N_14917);
or UO_253 (O_253,N_14275,N_14667);
and UO_254 (O_254,N_14607,N_14863);
and UO_255 (O_255,N_14677,N_14532);
nand UO_256 (O_256,N_14342,N_14453);
nand UO_257 (O_257,N_14647,N_14373);
nand UO_258 (O_258,N_14581,N_14463);
nor UO_259 (O_259,N_14254,N_14876);
and UO_260 (O_260,N_14265,N_14788);
or UO_261 (O_261,N_14883,N_14583);
nand UO_262 (O_262,N_14504,N_14324);
nor UO_263 (O_263,N_14467,N_14815);
or UO_264 (O_264,N_14907,N_14759);
and UO_265 (O_265,N_14482,N_14764);
and UO_266 (O_266,N_14714,N_14693);
or UO_267 (O_267,N_14514,N_14940);
or UO_268 (O_268,N_14943,N_14392);
nand UO_269 (O_269,N_14657,N_14281);
or UO_270 (O_270,N_14986,N_14864);
or UO_271 (O_271,N_14480,N_14869);
and UO_272 (O_272,N_14454,N_14680);
nor UO_273 (O_273,N_14908,N_14701);
and UO_274 (O_274,N_14326,N_14671);
nor UO_275 (O_275,N_14475,N_14748);
or UO_276 (O_276,N_14820,N_14707);
or UO_277 (O_277,N_14509,N_14384);
or UO_278 (O_278,N_14488,N_14653);
and UO_279 (O_279,N_14536,N_14276);
and UO_280 (O_280,N_14960,N_14314);
nor UO_281 (O_281,N_14266,N_14295);
nor UO_282 (O_282,N_14846,N_14571);
nor UO_283 (O_283,N_14621,N_14426);
nand UO_284 (O_284,N_14267,N_14589);
nand UO_285 (O_285,N_14773,N_14612);
xor UO_286 (O_286,N_14356,N_14874);
nor UO_287 (O_287,N_14271,N_14720);
nand UO_288 (O_288,N_14793,N_14329);
or UO_289 (O_289,N_14493,N_14993);
or UO_290 (O_290,N_14341,N_14662);
and UO_291 (O_291,N_14613,N_14305);
nand UO_292 (O_292,N_14512,N_14330);
or UO_293 (O_293,N_14870,N_14533);
or UO_294 (O_294,N_14375,N_14321);
nand UO_295 (O_295,N_14800,N_14619);
and UO_296 (O_296,N_14590,N_14346);
nor UO_297 (O_297,N_14415,N_14389);
or UO_298 (O_298,N_14728,N_14311);
or UO_299 (O_299,N_14867,N_14685);
nor UO_300 (O_300,N_14700,N_14552);
or UO_301 (O_301,N_14865,N_14352);
or UO_302 (O_302,N_14732,N_14399);
xnor UO_303 (O_303,N_14743,N_14543);
nor UO_304 (O_304,N_14358,N_14627);
nor UO_305 (O_305,N_14347,N_14830);
nor UO_306 (O_306,N_14817,N_14499);
or UO_307 (O_307,N_14998,N_14282);
nor UO_308 (O_308,N_14357,N_14928);
or UO_309 (O_309,N_14302,N_14713);
and UO_310 (O_310,N_14460,N_14854);
and UO_311 (O_311,N_14974,N_14857);
or UO_312 (O_312,N_14833,N_14697);
and UO_313 (O_313,N_14361,N_14272);
or UO_314 (O_314,N_14779,N_14990);
and UO_315 (O_315,N_14753,N_14526);
nand UO_316 (O_316,N_14402,N_14628);
or UO_317 (O_317,N_14525,N_14252);
and UO_318 (O_318,N_14439,N_14250);
or UO_319 (O_319,N_14269,N_14979);
and UO_320 (O_320,N_14988,N_14477);
or UO_321 (O_321,N_14660,N_14995);
nand UO_322 (O_322,N_14461,N_14465);
nand UO_323 (O_323,N_14652,N_14257);
nor UO_324 (O_324,N_14781,N_14502);
nand UO_325 (O_325,N_14564,N_14409);
nor UO_326 (O_326,N_14885,N_14320);
nor UO_327 (O_327,N_14777,N_14808);
and UO_328 (O_328,N_14570,N_14768);
nand UO_329 (O_329,N_14297,N_14969);
nor UO_330 (O_330,N_14505,N_14538);
or UO_331 (O_331,N_14429,N_14703);
nand UO_332 (O_332,N_14411,N_14364);
or UO_333 (O_333,N_14515,N_14599);
nand UO_334 (O_334,N_14718,N_14449);
nor UO_335 (O_335,N_14722,N_14383);
nor UO_336 (O_336,N_14573,N_14441);
or UO_337 (O_337,N_14849,N_14971);
nor UO_338 (O_338,N_14784,N_14698);
and UO_339 (O_339,N_14834,N_14919);
or UO_340 (O_340,N_14344,N_14920);
nor UO_341 (O_341,N_14901,N_14659);
nor UO_342 (O_342,N_14468,N_14424);
nand UO_343 (O_343,N_14586,N_14451);
xnor UO_344 (O_344,N_14622,N_14733);
or UO_345 (O_345,N_14258,N_14350);
and UO_346 (O_346,N_14479,N_14892);
nand UO_347 (O_347,N_14606,N_14669);
nand UO_348 (O_348,N_14639,N_14967);
and UO_349 (O_349,N_14385,N_14348);
nand UO_350 (O_350,N_14404,N_14294);
xor UO_351 (O_351,N_14561,N_14284);
or UO_352 (O_352,N_14927,N_14428);
or UO_353 (O_353,N_14715,N_14946);
nor UO_354 (O_354,N_14442,N_14537);
or UO_355 (O_355,N_14410,N_14418);
nand UO_356 (O_356,N_14359,N_14486);
nand UO_357 (O_357,N_14464,N_14560);
and UO_358 (O_358,N_14576,N_14836);
and UO_359 (O_359,N_14813,N_14641);
xnor UO_360 (O_360,N_14445,N_14638);
nand UO_361 (O_361,N_14654,N_14288);
nor UO_362 (O_362,N_14535,N_14684);
nand UO_363 (O_363,N_14283,N_14914);
or UO_364 (O_364,N_14481,N_14551);
nor UO_365 (O_365,N_14810,N_14818);
xnor UO_366 (O_366,N_14985,N_14742);
nor UO_367 (O_367,N_14436,N_14726);
and UO_368 (O_368,N_14755,N_14778);
and UO_369 (O_369,N_14601,N_14474);
and UO_370 (O_370,N_14762,N_14941);
or UO_371 (O_371,N_14651,N_14740);
and UO_372 (O_372,N_14749,N_14739);
nor UO_373 (O_373,N_14569,N_14648);
nor UO_374 (O_374,N_14682,N_14279);
or UO_375 (O_375,N_14590,N_14896);
or UO_376 (O_376,N_14654,N_14942);
nor UO_377 (O_377,N_14977,N_14289);
nand UO_378 (O_378,N_14733,N_14952);
and UO_379 (O_379,N_14691,N_14844);
and UO_380 (O_380,N_14480,N_14833);
nand UO_381 (O_381,N_14940,N_14664);
or UO_382 (O_382,N_14500,N_14400);
or UO_383 (O_383,N_14611,N_14703);
nor UO_384 (O_384,N_14885,N_14769);
and UO_385 (O_385,N_14750,N_14328);
nand UO_386 (O_386,N_14425,N_14344);
nand UO_387 (O_387,N_14673,N_14303);
nand UO_388 (O_388,N_14667,N_14289);
nor UO_389 (O_389,N_14763,N_14696);
nand UO_390 (O_390,N_14332,N_14283);
nor UO_391 (O_391,N_14503,N_14507);
nand UO_392 (O_392,N_14839,N_14903);
or UO_393 (O_393,N_14741,N_14335);
or UO_394 (O_394,N_14499,N_14805);
or UO_395 (O_395,N_14506,N_14690);
or UO_396 (O_396,N_14536,N_14842);
nand UO_397 (O_397,N_14460,N_14434);
nor UO_398 (O_398,N_14562,N_14893);
nand UO_399 (O_399,N_14518,N_14407);
and UO_400 (O_400,N_14320,N_14546);
nor UO_401 (O_401,N_14930,N_14927);
nand UO_402 (O_402,N_14434,N_14691);
or UO_403 (O_403,N_14786,N_14318);
or UO_404 (O_404,N_14770,N_14610);
nand UO_405 (O_405,N_14902,N_14324);
xnor UO_406 (O_406,N_14374,N_14828);
nor UO_407 (O_407,N_14609,N_14423);
nor UO_408 (O_408,N_14843,N_14312);
and UO_409 (O_409,N_14703,N_14980);
or UO_410 (O_410,N_14422,N_14773);
nand UO_411 (O_411,N_14260,N_14775);
nand UO_412 (O_412,N_14868,N_14731);
and UO_413 (O_413,N_14489,N_14862);
nor UO_414 (O_414,N_14556,N_14471);
nand UO_415 (O_415,N_14568,N_14326);
nand UO_416 (O_416,N_14572,N_14950);
or UO_417 (O_417,N_14693,N_14871);
xnor UO_418 (O_418,N_14687,N_14421);
nand UO_419 (O_419,N_14950,N_14877);
nand UO_420 (O_420,N_14410,N_14933);
and UO_421 (O_421,N_14318,N_14869);
nor UO_422 (O_422,N_14281,N_14351);
nand UO_423 (O_423,N_14958,N_14784);
nand UO_424 (O_424,N_14822,N_14733);
or UO_425 (O_425,N_14700,N_14257);
nor UO_426 (O_426,N_14646,N_14790);
and UO_427 (O_427,N_14825,N_14727);
or UO_428 (O_428,N_14974,N_14457);
and UO_429 (O_429,N_14417,N_14987);
nor UO_430 (O_430,N_14480,N_14380);
nand UO_431 (O_431,N_14852,N_14818);
or UO_432 (O_432,N_14330,N_14665);
and UO_433 (O_433,N_14696,N_14526);
xor UO_434 (O_434,N_14543,N_14909);
xnor UO_435 (O_435,N_14752,N_14862);
nand UO_436 (O_436,N_14959,N_14422);
nor UO_437 (O_437,N_14390,N_14911);
xnor UO_438 (O_438,N_14289,N_14714);
and UO_439 (O_439,N_14280,N_14818);
nand UO_440 (O_440,N_14992,N_14881);
or UO_441 (O_441,N_14777,N_14943);
nand UO_442 (O_442,N_14977,N_14678);
or UO_443 (O_443,N_14973,N_14931);
and UO_444 (O_444,N_14713,N_14915);
nor UO_445 (O_445,N_14404,N_14757);
and UO_446 (O_446,N_14857,N_14832);
nand UO_447 (O_447,N_14846,N_14623);
nand UO_448 (O_448,N_14592,N_14630);
nand UO_449 (O_449,N_14813,N_14505);
and UO_450 (O_450,N_14570,N_14954);
nor UO_451 (O_451,N_14324,N_14885);
nand UO_452 (O_452,N_14930,N_14536);
xnor UO_453 (O_453,N_14364,N_14260);
xnor UO_454 (O_454,N_14801,N_14418);
and UO_455 (O_455,N_14412,N_14784);
nand UO_456 (O_456,N_14424,N_14651);
xor UO_457 (O_457,N_14549,N_14817);
and UO_458 (O_458,N_14852,N_14346);
or UO_459 (O_459,N_14854,N_14297);
or UO_460 (O_460,N_14781,N_14709);
nor UO_461 (O_461,N_14757,N_14823);
and UO_462 (O_462,N_14616,N_14507);
and UO_463 (O_463,N_14518,N_14981);
or UO_464 (O_464,N_14860,N_14794);
nor UO_465 (O_465,N_14526,N_14372);
nor UO_466 (O_466,N_14926,N_14356);
nand UO_467 (O_467,N_14426,N_14563);
and UO_468 (O_468,N_14468,N_14843);
and UO_469 (O_469,N_14481,N_14705);
nor UO_470 (O_470,N_14775,N_14430);
nand UO_471 (O_471,N_14264,N_14911);
nor UO_472 (O_472,N_14439,N_14347);
xnor UO_473 (O_473,N_14326,N_14634);
nand UO_474 (O_474,N_14940,N_14300);
and UO_475 (O_475,N_14478,N_14808);
xnor UO_476 (O_476,N_14853,N_14302);
or UO_477 (O_477,N_14477,N_14343);
nor UO_478 (O_478,N_14766,N_14651);
nor UO_479 (O_479,N_14598,N_14631);
nand UO_480 (O_480,N_14422,N_14681);
nor UO_481 (O_481,N_14934,N_14497);
xor UO_482 (O_482,N_14866,N_14520);
and UO_483 (O_483,N_14744,N_14784);
or UO_484 (O_484,N_14608,N_14390);
xor UO_485 (O_485,N_14994,N_14909);
nand UO_486 (O_486,N_14519,N_14739);
xnor UO_487 (O_487,N_14478,N_14654);
xor UO_488 (O_488,N_14301,N_14808);
nor UO_489 (O_489,N_14547,N_14905);
nand UO_490 (O_490,N_14649,N_14532);
or UO_491 (O_491,N_14637,N_14833);
nand UO_492 (O_492,N_14780,N_14263);
nand UO_493 (O_493,N_14317,N_14837);
and UO_494 (O_494,N_14251,N_14296);
nand UO_495 (O_495,N_14756,N_14760);
nor UO_496 (O_496,N_14608,N_14269);
or UO_497 (O_497,N_14723,N_14563);
nor UO_498 (O_498,N_14423,N_14510);
and UO_499 (O_499,N_14990,N_14629);
nand UO_500 (O_500,N_14742,N_14278);
xor UO_501 (O_501,N_14922,N_14871);
nor UO_502 (O_502,N_14791,N_14418);
nand UO_503 (O_503,N_14634,N_14452);
and UO_504 (O_504,N_14277,N_14337);
or UO_505 (O_505,N_14876,N_14309);
or UO_506 (O_506,N_14789,N_14979);
nor UO_507 (O_507,N_14273,N_14962);
nor UO_508 (O_508,N_14369,N_14368);
nor UO_509 (O_509,N_14381,N_14554);
nand UO_510 (O_510,N_14783,N_14569);
or UO_511 (O_511,N_14614,N_14310);
nor UO_512 (O_512,N_14675,N_14802);
or UO_513 (O_513,N_14629,N_14679);
nor UO_514 (O_514,N_14361,N_14715);
and UO_515 (O_515,N_14804,N_14470);
or UO_516 (O_516,N_14853,N_14747);
and UO_517 (O_517,N_14950,N_14376);
and UO_518 (O_518,N_14995,N_14265);
nor UO_519 (O_519,N_14776,N_14477);
nand UO_520 (O_520,N_14522,N_14910);
nor UO_521 (O_521,N_14800,N_14759);
and UO_522 (O_522,N_14825,N_14265);
and UO_523 (O_523,N_14791,N_14378);
xnor UO_524 (O_524,N_14608,N_14420);
or UO_525 (O_525,N_14768,N_14461);
and UO_526 (O_526,N_14800,N_14344);
and UO_527 (O_527,N_14999,N_14522);
nand UO_528 (O_528,N_14925,N_14553);
and UO_529 (O_529,N_14952,N_14515);
or UO_530 (O_530,N_14657,N_14958);
or UO_531 (O_531,N_14913,N_14511);
and UO_532 (O_532,N_14485,N_14673);
nor UO_533 (O_533,N_14791,N_14547);
nand UO_534 (O_534,N_14856,N_14647);
nand UO_535 (O_535,N_14840,N_14829);
nand UO_536 (O_536,N_14842,N_14832);
or UO_537 (O_537,N_14848,N_14997);
and UO_538 (O_538,N_14288,N_14984);
and UO_539 (O_539,N_14648,N_14976);
nand UO_540 (O_540,N_14431,N_14538);
or UO_541 (O_541,N_14725,N_14933);
or UO_542 (O_542,N_14397,N_14506);
or UO_543 (O_543,N_14643,N_14988);
nor UO_544 (O_544,N_14501,N_14474);
nor UO_545 (O_545,N_14549,N_14704);
or UO_546 (O_546,N_14909,N_14758);
nand UO_547 (O_547,N_14391,N_14928);
nand UO_548 (O_548,N_14775,N_14364);
nor UO_549 (O_549,N_14695,N_14631);
or UO_550 (O_550,N_14703,N_14884);
nand UO_551 (O_551,N_14874,N_14931);
and UO_552 (O_552,N_14717,N_14691);
nand UO_553 (O_553,N_14712,N_14994);
nor UO_554 (O_554,N_14626,N_14818);
xor UO_555 (O_555,N_14709,N_14972);
nor UO_556 (O_556,N_14482,N_14354);
or UO_557 (O_557,N_14850,N_14757);
nor UO_558 (O_558,N_14810,N_14992);
nor UO_559 (O_559,N_14496,N_14305);
or UO_560 (O_560,N_14691,N_14532);
xor UO_561 (O_561,N_14580,N_14367);
xor UO_562 (O_562,N_14698,N_14367);
nand UO_563 (O_563,N_14950,N_14790);
and UO_564 (O_564,N_14738,N_14321);
nand UO_565 (O_565,N_14716,N_14672);
xnor UO_566 (O_566,N_14676,N_14358);
and UO_567 (O_567,N_14975,N_14321);
nand UO_568 (O_568,N_14276,N_14803);
nor UO_569 (O_569,N_14908,N_14650);
and UO_570 (O_570,N_14345,N_14683);
and UO_571 (O_571,N_14663,N_14492);
and UO_572 (O_572,N_14760,N_14672);
nand UO_573 (O_573,N_14723,N_14268);
or UO_574 (O_574,N_14421,N_14413);
and UO_575 (O_575,N_14332,N_14492);
and UO_576 (O_576,N_14395,N_14353);
xnor UO_577 (O_577,N_14573,N_14717);
nand UO_578 (O_578,N_14653,N_14479);
xnor UO_579 (O_579,N_14688,N_14323);
and UO_580 (O_580,N_14301,N_14743);
or UO_581 (O_581,N_14345,N_14251);
nand UO_582 (O_582,N_14901,N_14388);
and UO_583 (O_583,N_14626,N_14383);
nor UO_584 (O_584,N_14625,N_14888);
nor UO_585 (O_585,N_14512,N_14400);
or UO_586 (O_586,N_14394,N_14543);
or UO_587 (O_587,N_14325,N_14833);
or UO_588 (O_588,N_14396,N_14778);
and UO_589 (O_589,N_14673,N_14722);
or UO_590 (O_590,N_14366,N_14761);
nor UO_591 (O_591,N_14522,N_14503);
or UO_592 (O_592,N_14919,N_14983);
nand UO_593 (O_593,N_14838,N_14691);
and UO_594 (O_594,N_14272,N_14515);
or UO_595 (O_595,N_14781,N_14261);
or UO_596 (O_596,N_14432,N_14602);
nand UO_597 (O_597,N_14769,N_14435);
nand UO_598 (O_598,N_14648,N_14257);
nand UO_599 (O_599,N_14836,N_14838);
nand UO_600 (O_600,N_14670,N_14712);
nor UO_601 (O_601,N_14808,N_14585);
or UO_602 (O_602,N_14458,N_14322);
nor UO_603 (O_603,N_14290,N_14383);
nand UO_604 (O_604,N_14966,N_14810);
xnor UO_605 (O_605,N_14480,N_14259);
and UO_606 (O_606,N_14370,N_14353);
and UO_607 (O_607,N_14950,N_14906);
or UO_608 (O_608,N_14797,N_14647);
nand UO_609 (O_609,N_14733,N_14635);
or UO_610 (O_610,N_14980,N_14583);
xor UO_611 (O_611,N_14377,N_14432);
nor UO_612 (O_612,N_14276,N_14996);
and UO_613 (O_613,N_14632,N_14385);
nand UO_614 (O_614,N_14270,N_14506);
nand UO_615 (O_615,N_14634,N_14832);
or UO_616 (O_616,N_14330,N_14751);
or UO_617 (O_617,N_14281,N_14273);
nor UO_618 (O_618,N_14582,N_14727);
nor UO_619 (O_619,N_14749,N_14889);
xnor UO_620 (O_620,N_14572,N_14920);
and UO_621 (O_621,N_14456,N_14728);
and UO_622 (O_622,N_14631,N_14508);
or UO_623 (O_623,N_14424,N_14684);
and UO_624 (O_624,N_14592,N_14414);
and UO_625 (O_625,N_14502,N_14286);
nor UO_626 (O_626,N_14740,N_14284);
or UO_627 (O_627,N_14720,N_14309);
nand UO_628 (O_628,N_14537,N_14391);
nor UO_629 (O_629,N_14441,N_14284);
and UO_630 (O_630,N_14514,N_14859);
nor UO_631 (O_631,N_14516,N_14344);
xor UO_632 (O_632,N_14493,N_14448);
or UO_633 (O_633,N_14566,N_14859);
nand UO_634 (O_634,N_14631,N_14259);
or UO_635 (O_635,N_14752,N_14526);
and UO_636 (O_636,N_14559,N_14333);
xor UO_637 (O_637,N_14473,N_14820);
nand UO_638 (O_638,N_14538,N_14768);
xor UO_639 (O_639,N_14852,N_14825);
and UO_640 (O_640,N_14373,N_14685);
and UO_641 (O_641,N_14652,N_14778);
xor UO_642 (O_642,N_14781,N_14705);
nor UO_643 (O_643,N_14841,N_14958);
xor UO_644 (O_644,N_14957,N_14547);
xor UO_645 (O_645,N_14467,N_14729);
and UO_646 (O_646,N_14405,N_14917);
or UO_647 (O_647,N_14493,N_14807);
or UO_648 (O_648,N_14317,N_14871);
nor UO_649 (O_649,N_14468,N_14276);
xnor UO_650 (O_650,N_14677,N_14465);
nand UO_651 (O_651,N_14365,N_14419);
nand UO_652 (O_652,N_14527,N_14570);
and UO_653 (O_653,N_14536,N_14412);
nand UO_654 (O_654,N_14825,N_14592);
or UO_655 (O_655,N_14908,N_14655);
nand UO_656 (O_656,N_14733,N_14644);
nor UO_657 (O_657,N_14724,N_14642);
or UO_658 (O_658,N_14690,N_14507);
and UO_659 (O_659,N_14358,N_14397);
nand UO_660 (O_660,N_14526,N_14319);
nor UO_661 (O_661,N_14400,N_14323);
and UO_662 (O_662,N_14974,N_14287);
xnor UO_663 (O_663,N_14542,N_14305);
and UO_664 (O_664,N_14746,N_14397);
nand UO_665 (O_665,N_14439,N_14876);
nor UO_666 (O_666,N_14845,N_14723);
and UO_667 (O_667,N_14959,N_14976);
or UO_668 (O_668,N_14866,N_14813);
nor UO_669 (O_669,N_14967,N_14445);
or UO_670 (O_670,N_14807,N_14726);
nor UO_671 (O_671,N_14380,N_14753);
and UO_672 (O_672,N_14842,N_14592);
or UO_673 (O_673,N_14802,N_14888);
nand UO_674 (O_674,N_14994,N_14615);
or UO_675 (O_675,N_14864,N_14610);
nor UO_676 (O_676,N_14305,N_14447);
and UO_677 (O_677,N_14708,N_14896);
nor UO_678 (O_678,N_14405,N_14852);
or UO_679 (O_679,N_14917,N_14262);
nand UO_680 (O_680,N_14373,N_14446);
and UO_681 (O_681,N_14926,N_14427);
nand UO_682 (O_682,N_14822,N_14426);
nand UO_683 (O_683,N_14580,N_14345);
nand UO_684 (O_684,N_14511,N_14900);
nor UO_685 (O_685,N_14595,N_14465);
nand UO_686 (O_686,N_14870,N_14277);
and UO_687 (O_687,N_14591,N_14974);
and UO_688 (O_688,N_14466,N_14396);
nand UO_689 (O_689,N_14641,N_14990);
nor UO_690 (O_690,N_14956,N_14605);
or UO_691 (O_691,N_14527,N_14937);
and UO_692 (O_692,N_14571,N_14290);
xnor UO_693 (O_693,N_14373,N_14912);
and UO_694 (O_694,N_14425,N_14296);
or UO_695 (O_695,N_14919,N_14797);
nand UO_696 (O_696,N_14497,N_14479);
and UO_697 (O_697,N_14618,N_14558);
or UO_698 (O_698,N_14496,N_14294);
nand UO_699 (O_699,N_14391,N_14445);
nor UO_700 (O_700,N_14954,N_14382);
or UO_701 (O_701,N_14570,N_14390);
or UO_702 (O_702,N_14622,N_14761);
nand UO_703 (O_703,N_14394,N_14676);
nor UO_704 (O_704,N_14574,N_14699);
nor UO_705 (O_705,N_14680,N_14286);
nor UO_706 (O_706,N_14915,N_14491);
nand UO_707 (O_707,N_14577,N_14563);
and UO_708 (O_708,N_14907,N_14853);
xnor UO_709 (O_709,N_14966,N_14998);
and UO_710 (O_710,N_14812,N_14782);
and UO_711 (O_711,N_14265,N_14890);
nand UO_712 (O_712,N_14888,N_14754);
nand UO_713 (O_713,N_14268,N_14610);
nand UO_714 (O_714,N_14466,N_14292);
nor UO_715 (O_715,N_14713,N_14584);
nor UO_716 (O_716,N_14260,N_14499);
nor UO_717 (O_717,N_14499,N_14251);
nor UO_718 (O_718,N_14687,N_14778);
nor UO_719 (O_719,N_14802,N_14941);
nor UO_720 (O_720,N_14870,N_14312);
or UO_721 (O_721,N_14542,N_14911);
or UO_722 (O_722,N_14823,N_14688);
or UO_723 (O_723,N_14265,N_14803);
nor UO_724 (O_724,N_14746,N_14634);
and UO_725 (O_725,N_14411,N_14500);
or UO_726 (O_726,N_14808,N_14639);
or UO_727 (O_727,N_14498,N_14869);
nor UO_728 (O_728,N_14603,N_14499);
nor UO_729 (O_729,N_14695,N_14419);
and UO_730 (O_730,N_14414,N_14267);
and UO_731 (O_731,N_14892,N_14280);
nand UO_732 (O_732,N_14778,N_14668);
nand UO_733 (O_733,N_14367,N_14715);
or UO_734 (O_734,N_14739,N_14691);
xor UO_735 (O_735,N_14981,N_14524);
nor UO_736 (O_736,N_14934,N_14284);
nor UO_737 (O_737,N_14260,N_14890);
nand UO_738 (O_738,N_14544,N_14383);
xnor UO_739 (O_739,N_14711,N_14439);
xor UO_740 (O_740,N_14756,N_14781);
xor UO_741 (O_741,N_14402,N_14804);
xnor UO_742 (O_742,N_14922,N_14258);
and UO_743 (O_743,N_14286,N_14988);
and UO_744 (O_744,N_14908,N_14541);
and UO_745 (O_745,N_14307,N_14495);
or UO_746 (O_746,N_14665,N_14493);
and UO_747 (O_747,N_14584,N_14465);
xor UO_748 (O_748,N_14716,N_14985);
nor UO_749 (O_749,N_14580,N_14944);
nor UO_750 (O_750,N_14847,N_14465);
or UO_751 (O_751,N_14304,N_14716);
and UO_752 (O_752,N_14695,N_14700);
nor UO_753 (O_753,N_14486,N_14810);
nor UO_754 (O_754,N_14935,N_14405);
xnor UO_755 (O_755,N_14724,N_14647);
or UO_756 (O_756,N_14495,N_14921);
and UO_757 (O_757,N_14635,N_14801);
nand UO_758 (O_758,N_14446,N_14891);
nor UO_759 (O_759,N_14517,N_14315);
nand UO_760 (O_760,N_14821,N_14996);
or UO_761 (O_761,N_14908,N_14380);
or UO_762 (O_762,N_14862,N_14905);
nand UO_763 (O_763,N_14637,N_14365);
nand UO_764 (O_764,N_14271,N_14691);
nand UO_765 (O_765,N_14956,N_14625);
nor UO_766 (O_766,N_14648,N_14609);
xor UO_767 (O_767,N_14498,N_14294);
and UO_768 (O_768,N_14668,N_14674);
nand UO_769 (O_769,N_14770,N_14511);
xor UO_770 (O_770,N_14524,N_14339);
or UO_771 (O_771,N_14840,N_14591);
nor UO_772 (O_772,N_14809,N_14715);
and UO_773 (O_773,N_14778,N_14320);
and UO_774 (O_774,N_14348,N_14571);
or UO_775 (O_775,N_14393,N_14499);
xor UO_776 (O_776,N_14553,N_14499);
nor UO_777 (O_777,N_14845,N_14888);
nor UO_778 (O_778,N_14550,N_14899);
xnor UO_779 (O_779,N_14604,N_14559);
nand UO_780 (O_780,N_14873,N_14533);
nor UO_781 (O_781,N_14514,N_14707);
xnor UO_782 (O_782,N_14365,N_14559);
or UO_783 (O_783,N_14938,N_14382);
and UO_784 (O_784,N_14404,N_14925);
nand UO_785 (O_785,N_14333,N_14486);
xnor UO_786 (O_786,N_14316,N_14759);
or UO_787 (O_787,N_14658,N_14868);
nor UO_788 (O_788,N_14709,N_14814);
nor UO_789 (O_789,N_14434,N_14706);
nand UO_790 (O_790,N_14563,N_14284);
or UO_791 (O_791,N_14703,N_14914);
nand UO_792 (O_792,N_14948,N_14440);
nand UO_793 (O_793,N_14639,N_14898);
nand UO_794 (O_794,N_14774,N_14457);
nand UO_795 (O_795,N_14814,N_14863);
nor UO_796 (O_796,N_14737,N_14639);
xnor UO_797 (O_797,N_14292,N_14302);
or UO_798 (O_798,N_14804,N_14986);
nor UO_799 (O_799,N_14291,N_14371);
and UO_800 (O_800,N_14839,N_14567);
or UO_801 (O_801,N_14594,N_14970);
or UO_802 (O_802,N_14286,N_14501);
nor UO_803 (O_803,N_14933,N_14863);
or UO_804 (O_804,N_14790,N_14913);
or UO_805 (O_805,N_14855,N_14724);
and UO_806 (O_806,N_14808,N_14711);
nor UO_807 (O_807,N_14810,N_14950);
nor UO_808 (O_808,N_14668,N_14747);
or UO_809 (O_809,N_14956,N_14307);
nand UO_810 (O_810,N_14414,N_14754);
nor UO_811 (O_811,N_14481,N_14744);
or UO_812 (O_812,N_14719,N_14262);
nor UO_813 (O_813,N_14541,N_14832);
and UO_814 (O_814,N_14362,N_14373);
or UO_815 (O_815,N_14699,N_14871);
or UO_816 (O_816,N_14719,N_14798);
and UO_817 (O_817,N_14736,N_14454);
nor UO_818 (O_818,N_14349,N_14792);
nor UO_819 (O_819,N_14955,N_14353);
nor UO_820 (O_820,N_14438,N_14445);
or UO_821 (O_821,N_14927,N_14602);
or UO_822 (O_822,N_14547,N_14568);
nor UO_823 (O_823,N_14537,N_14652);
and UO_824 (O_824,N_14452,N_14968);
nand UO_825 (O_825,N_14529,N_14866);
or UO_826 (O_826,N_14320,N_14697);
or UO_827 (O_827,N_14400,N_14798);
nor UO_828 (O_828,N_14893,N_14368);
and UO_829 (O_829,N_14579,N_14607);
and UO_830 (O_830,N_14963,N_14316);
xor UO_831 (O_831,N_14353,N_14587);
or UO_832 (O_832,N_14905,N_14712);
or UO_833 (O_833,N_14882,N_14291);
nand UO_834 (O_834,N_14432,N_14284);
nand UO_835 (O_835,N_14806,N_14830);
nand UO_836 (O_836,N_14622,N_14602);
and UO_837 (O_837,N_14892,N_14291);
nand UO_838 (O_838,N_14265,N_14627);
nand UO_839 (O_839,N_14942,N_14617);
or UO_840 (O_840,N_14375,N_14474);
and UO_841 (O_841,N_14551,N_14766);
nand UO_842 (O_842,N_14608,N_14600);
nand UO_843 (O_843,N_14911,N_14308);
nand UO_844 (O_844,N_14784,N_14777);
nand UO_845 (O_845,N_14423,N_14638);
or UO_846 (O_846,N_14592,N_14975);
or UO_847 (O_847,N_14709,N_14554);
or UO_848 (O_848,N_14492,N_14260);
nor UO_849 (O_849,N_14394,N_14668);
nand UO_850 (O_850,N_14310,N_14404);
or UO_851 (O_851,N_14386,N_14590);
nand UO_852 (O_852,N_14382,N_14808);
xnor UO_853 (O_853,N_14699,N_14307);
nor UO_854 (O_854,N_14569,N_14340);
and UO_855 (O_855,N_14322,N_14981);
and UO_856 (O_856,N_14475,N_14904);
xor UO_857 (O_857,N_14495,N_14382);
or UO_858 (O_858,N_14340,N_14598);
and UO_859 (O_859,N_14464,N_14576);
or UO_860 (O_860,N_14467,N_14681);
and UO_861 (O_861,N_14394,N_14650);
nor UO_862 (O_862,N_14901,N_14424);
or UO_863 (O_863,N_14412,N_14522);
nor UO_864 (O_864,N_14305,N_14391);
nor UO_865 (O_865,N_14698,N_14285);
or UO_866 (O_866,N_14334,N_14871);
and UO_867 (O_867,N_14530,N_14381);
or UO_868 (O_868,N_14608,N_14286);
nand UO_869 (O_869,N_14991,N_14837);
and UO_870 (O_870,N_14920,N_14524);
nand UO_871 (O_871,N_14426,N_14393);
nand UO_872 (O_872,N_14329,N_14813);
nand UO_873 (O_873,N_14712,N_14522);
or UO_874 (O_874,N_14637,N_14677);
or UO_875 (O_875,N_14580,N_14656);
nor UO_876 (O_876,N_14649,N_14758);
or UO_877 (O_877,N_14351,N_14986);
or UO_878 (O_878,N_14691,N_14693);
and UO_879 (O_879,N_14783,N_14910);
and UO_880 (O_880,N_14352,N_14312);
or UO_881 (O_881,N_14972,N_14408);
and UO_882 (O_882,N_14332,N_14779);
or UO_883 (O_883,N_14359,N_14489);
or UO_884 (O_884,N_14838,N_14798);
and UO_885 (O_885,N_14992,N_14927);
or UO_886 (O_886,N_14887,N_14513);
or UO_887 (O_887,N_14958,N_14449);
xnor UO_888 (O_888,N_14342,N_14481);
nand UO_889 (O_889,N_14259,N_14918);
or UO_890 (O_890,N_14546,N_14914);
or UO_891 (O_891,N_14578,N_14957);
or UO_892 (O_892,N_14784,N_14362);
nand UO_893 (O_893,N_14436,N_14898);
nand UO_894 (O_894,N_14466,N_14619);
and UO_895 (O_895,N_14922,N_14611);
or UO_896 (O_896,N_14742,N_14505);
nand UO_897 (O_897,N_14995,N_14645);
nand UO_898 (O_898,N_14529,N_14705);
and UO_899 (O_899,N_14373,N_14563);
and UO_900 (O_900,N_14836,N_14627);
nand UO_901 (O_901,N_14773,N_14923);
xor UO_902 (O_902,N_14343,N_14684);
xnor UO_903 (O_903,N_14399,N_14729);
nor UO_904 (O_904,N_14462,N_14697);
and UO_905 (O_905,N_14977,N_14983);
and UO_906 (O_906,N_14999,N_14286);
nand UO_907 (O_907,N_14994,N_14930);
and UO_908 (O_908,N_14783,N_14679);
nor UO_909 (O_909,N_14587,N_14636);
and UO_910 (O_910,N_14406,N_14699);
nand UO_911 (O_911,N_14792,N_14453);
and UO_912 (O_912,N_14512,N_14810);
nor UO_913 (O_913,N_14319,N_14988);
nand UO_914 (O_914,N_14357,N_14793);
or UO_915 (O_915,N_14936,N_14307);
nor UO_916 (O_916,N_14382,N_14892);
or UO_917 (O_917,N_14423,N_14809);
or UO_918 (O_918,N_14669,N_14469);
nand UO_919 (O_919,N_14441,N_14961);
and UO_920 (O_920,N_14383,N_14584);
nand UO_921 (O_921,N_14779,N_14620);
nand UO_922 (O_922,N_14964,N_14853);
and UO_923 (O_923,N_14663,N_14799);
or UO_924 (O_924,N_14620,N_14896);
or UO_925 (O_925,N_14709,N_14930);
nand UO_926 (O_926,N_14592,N_14508);
and UO_927 (O_927,N_14340,N_14351);
nor UO_928 (O_928,N_14438,N_14555);
or UO_929 (O_929,N_14841,N_14395);
nand UO_930 (O_930,N_14940,N_14494);
and UO_931 (O_931,N_14903,N_14628);
or UO_932 (O_932,N_14396,N_14649);
nand UO_933 (O_933,N_14510,N_14348);
nand UO_934 (O_934,N_14792,N_14774);
and UO_935 (O_935,N_14779,N_14843);
or UO_936 (O_936,N_14539,N_14831);
xnor UO_937 (O_937,N_14633,N_14673);
nand UO_938 (O_938,N_14272,N_14443);
and UO_939 (O_939,N_14501,N_14405);
nor UO_940 (O_940,N_14570,N_14796);
nor UO_941 (O_941,N_14364,N_14603);
xor UO_942 (O_942,N_14995,N_14405);
nor UO_943 (O_943,N_14882,N_14631);
nand UO_944 (O_944,N_14635,N_14893);
nor UO_945 (O_945,N_14863,N_14328);
or UO_946 (O_946,N_14452,N_14661);
or UO_947 (O_947,N_14457,N_14898);
or UO_948 (O_948,N_14265,N_14782);
nand UO_949 (O_949,N_14753,N_14404);
nand UO_950 (O_950,N_14318,N_14438);
nand UO_951 (O_951,N_14947,N_14335);
nand UO_952 (O_952,N_14515,N_14868);
nand UO_953 (O_953,N_14868,N_14743);
xor UO_954 (O_954,N_14533,N_14766);
nand UO_955 (O_955,N_14969,N_14656);
nand UO_956 (O_956,N_14900,N_14749);
xor UO_957 (O_957,N_14267,N_14466);
nand UO_958 (O_958,N_14588,N_14683);
and UO_959 (O_959,N_14358,N_14927);
or UO_960 (O_960,N_14278,N_14934);
or UO_961 (O_961,N_14738,N_14330);
nand UO_962 (O_962,N_14946,N_14901);
nand UO_963 (O_963,N_14962,N_14876);
nand UO_964 (O_964,N_14492,N_14361);
and UO_965 (O_965,N_14279,N_14674);
nor UO_966 (O_966,N_14352,N_14500);
and UO_967 (O_967,N_14557,N_14484);
or UO_968 (O_968,N_14760,N_14680);
nand UO_969 (O_969,N_14658,N_14920);
nand UO_970 (O_970,N_14950,N_14816);
nand UO_971 (O_971,N_14311,N_14580);
xor UO_972 (O_972,N_14960,N_14796);
and UO_973 (O_973,N_14577,N_14730);
and UO_974 (O_974,N_14346,N_14585);
or UO_975 (O_975,N_14730,N_14264);
or UO_976 (O_976,N_14626,N_14949);
or UO_977 (O_977,N_14847,N_14506);
xnor UO_978 (O_978,N_14867,N_14460);
and UO_979 (O_979,N_14297,N_14917);
nand UO_980 (O_980,N_14263,N_14528);
nor UO_981 (O_981,N_14278,N_14823);
nor UO_982 (O_982,N_14812,N_14637);
nand UO_983 (O_983,N_14880,N_14277);
nand UO_984 (O_984,N_14985,N_14542);
nand UO_985 (O_985,N_14844,N_14531);
nor UO_986 (O_986,N_14308,N_14543);
nand UO_987 (O_987,N_14721,N_14581);
nand UO_988 (O_988,N_14606,N_14828);
nor UO_989 (O_989,N_14771,N_14649);
or UO_990 (O_990,N_14851,N_14583);
and UO_991 (O_991,N_14652,N_14829);
and UO_992 (O_992,N_14444,N_14421);
or UO_993 (O_993,N_14924,N_14272);
and UO_994 (O_994,N_14595,N_14446);
xor UO_995 (O_995,N_14443,N_14738);
and UO_996 (O_996,N_14777,N_14750);
and UO_997 (O_997,N_14351,N_14411);
and UO_998 (O_998,N_14736,N_14839);
xor UO_999 (O_999,N_14552,N_14672);
and UO_1000 (O_1000,N_14347,N_14892);
or UO_1001 (O_1001,N_14625,N_14879);
and UO_1002 (O_1002,N_14274,N_14889);
xnor UO_1003 (O_1003,N_14944,N_14417);
nand UO_1004 (O_1004,N_14685,N_14493);
nand UO_1005 (O_1005,N_14924,N_14823);
nand UO_1006 (O_1006,N_14647,N_14519);
or UO_1007 (O_1007,N_14653,N_14564);
nor UO_1008 (O_1008,N_14877,N_14782);
nor UO_1009 (O_1009,N_14339,N_14329);
nor UO_1010 (O_1010,N_14548,N_14635);
xnor UO_1011 (O_1011,N_14393,N_14763);
or UO_1012 (O_1012,N_14586,N_14967);
nor UO_1013 (O_1013,N_14491,N_14460);
nor UO_1014 (O_1014,N_14832,N_14906);
and UO_1015 (O_1015,N_14616,N_14589);
xnor UO_1016 (O_1016,N_14901,N_14466);
xnor UO_1017 (O_1017,N_14828,N_14323);
or UO_1018 (O_1018,N_14867,N_14654);
nand UO_1019 (O_1019,N_14944,N_14716);
xnor UO_1020 (O_1020,N_14938,N_14655);
nor UO_1021 (O_1021,N_14815,N_14430);
nand UO_1022 (O_1022,N_14684,N_14788);
or UO_1023 (O_1023,N_14613,N_14727);
or UO_1024 (O_1024,N_14933,N_14982);
and UO_1025 (O_1025,N_14418,N_14651);
nor UO_1026 (O_1026,N_14827,N_14868);
and UO_1027 (O_1027,N_14779,N_14972);
and UO_1028 (O_1028,N_14619,N_14865);
and UO_1029 (O_1029,N_14534,N_14959);
or UO_1030 (O_1030,N_14692,N_14483);
or UO_1031 (O_1031,N_14668,N_14331);
and UO_1032 (O_1032,N_14871,N_14599);
and UO_1033 (O_1033,N_14500,N_14779);
or UO_1034 (O_1034,N_14909,N_14732);
nand UO_1035 (O_1035,N_14515,N_14410);
or UO_1036 (O_1036,N_14894,N_14687);
nand UO_1037 (O_1037,N_14289,N_14261);
or UO_1038 (O_1038,N_14871,N_14608);
or UO_1039 (O_1039,N_14638,N_14896);
nor UO_1040 (O_1040,N_14518,N_14911);
and UO_1041 (O_1041,N_14788,N_14680);
or UO_1042 (O_1042,N_14557,N_14345);
nand UO_1043 (O_1043,N_14284,N_14682);
nor UO_1044 (O_1044,N_14286,N_14990);
nor UO_1045 (O_1045,N_14814,N_14897);
nor UO_1046 (O_1046,N_14719,N_14576);
and UO_1047 (O_1047,N_14773,N_14732);
nor UO_1048 (O_1048,N_14774,N_14587);
nand UO_1049 (O_1049,N_14878,N_14359);
or UO_1050 (O_1050,N_14808,N_14722);
or UO_1051 (O_1051,N_14966,N_14639);
xor UO_1052 (O_1052,N_14345,N_14784);
xnor UO_1053 (O_1053,N_14265,N_14967);
or UO_1054 (O_1054,N_14274,N_14942);
and UO_1055 (O_1055,N_14897,N_14483);
and UO_1056 (O_1056,N_14923,N_14432);
and UO_1057 (O_1057,N_14941,N_14400);
and UO_1058 (O_1058,N_14463,N_14292);
or UO_1059 (O_1059,N_14846,N_14878);
nand UO_1060 (O_1060,N_14772,N_14882);
and UO_1061 (O_1061,N_14516,N_14839);
nor UO_1062 (O_1062,N_14925,N_14509);
xnor UO_1063 (O_1063,N_14649,N_14992);
or UO_1064 (O_1064,N_14436,N_14733);
nor UO_1065 (O_1065,N_14862,N_14549);
nor UO_1066 (O_1066,N_14890,N_14775);
nand UO_1067 (O_1067,N_14701,N_14557);
nor UO_1068 (O_1068,N_14777,N_14363);
nor UO_1069 (O_1069,N_14642,N_14740);
nand UO_1070 (O_1070,N_14423,N_14417);
nor UO_1071 (O_1071,N_14267,N_14881);
nor UO_1072 (O_1072,N_14851,N_14319);
nor UO_1073 (O_1073,N_14463,N_14390);
or UO_1074 (O_1074,N_14617,N_14681);
nand UO_1075 (O_1075,N_14955,N_14705);
nor UO_1076 (O_1076,N_14653,N_14625);
nand UO_1077 (O_1077,N_14396,N_14356);
and UO_1078 (O_1078,N_14611,N_14843);
nor UO_1079 (O_1079,N_14412,N_14771);
xnor UO_1080 (O_1080,N_14553,N_14978);
and UO_1081 (O_1081,N_14678,N_14294);
and UO_1082 (O_1082,N_14363,N_14995);
nand UO_1083 (O_1083,N_14375,N_14760);
nand UO_1084 (O_1084,N_14480,N_14907);
nand UO_1085 (O_1085,N_14587,N_14506);
xnor UO_1086 (O_1086,N_14801,N_14455);
and UO_1087 (O_1087,N_14734,N_14368);
and UO_1088 (O_1088,N_14608,N_14442);
nor UO_1089 (O_1089,N_14459,N_14418);
or UO_1090 (O_1090,N_14857,N_14760);
nor UO_1091 (O_1091,N_14288,N_14508);
and UO_1092 (O_1092,N_14574,N_14896);
and UO_1093 (O_1093,N_14524,N_14802);
and UO_1094 (O_1094,N_14370,N_14577);
nand UO_1095 (O_1095,N_14519,N_14517);
nand UO_1096 (O_1096,N_14956,N_14800);
and UO_1097 (O_1097,N_14595,N_14906);
or UO_1098 (O_1098,N_14750,N_14415);
or UO_1099 (O_1099,N_14324,N_14400);
nand UO_1100 (O_1100,N_14921,N_14363);
nor UO_1101 (O_1101,N_14351,N_14857);
or UO_1102 (O_1102,N_14515,N_14490);
nand UO_1103 (O_1103,N_14846,N_14735);
and UO_1104 (O_1104,N_14609,N_14947);
and UO_1105 (O_1105,N_14953,N_14289);
and UO_1106 (O_1106,N_14762,N_14772);
nand UO_1107 (O_1107,N_14558,N_14677);
nand UO_1108 (O_1108,N_14953,N_14969);
or UO_1109 (O_1109,N_14899,N_14760);
or UO_1110 (O_1110,N_14963,N_14977);
nor UO_1111 (O_1111,N_14540,N_14291);
or UO_1112 (O_1112,N_14861,N_14671);
nor UO_1113 (O_1113,N_14962,N_14683);
nand UO_1114 (O_1114,N_14386,N_14550);
or UO_1115 (O_1115,N_14896,N_14973);
nand UO_1116 (O_1116,N_14332,N_14511);
or UO_1117 (O_1117,N_14261,N_14598);
or UO_1118 (O_1118,N_14278,N_14261);
and UO_1119 (O_1119,N_14400,N_14865);
and UO_1120 (O_1120,N_14753,N_14664);
or UO_1121 (O_1121,N_14957,N_14587);
or UO_1122 (O_1122,N_14315,N_14494);
nand UO_1123 (O_1123,N_14483,N_14676);
nand UO_1124 (O_1124,N_14424,N_14889);
nor UO_1125 (O_1125,N_14997,N_14257);
nand UO_1126 (O_1126,N_14789,N_14627);
nor UO_1127 (O_1127,N_14277,N_14886);
and UO_1128 (O_1128,N_14333,N_14459);
and UO_1129 (O_1129,N_14448,N_14518);
and UO_1130 (O_1130,N_14996,N_14760);
or UO_1131 (O_1131,N_14819,N_14837);
nor UO_1132 (O_1132,N_14928,N_14581);
and UO_1133 (O_1133,N_14924,N_14790);
or UO_1134 (O_1134,N_14931,N_14942);
and UO_1135 (O_1135,N_14371,N_14778);
or UO_1136 (O_1136,N_14523,N_14430);
nor UO_1137 (O_1137,N_14603,N_14987);
nor UO_1138 (O_1138,N_14811,N_14373);
nand UO_1139 (O_1139,N_14431,N_14489);
nand UO_1140 (O_1140,N_14723,N_14470);
xnor UO_1141 (O_1141,N_14372,N_14623);
or UO_1142 (O_1142,N_14954,N_14415);
or UO_1143 (O_1143,N_14397,N_14879);
nand UO_1144 (O_1144,N_14696,N_14747);
and UO_1145 (O_1145,N_14733,N_14966);
or UO_1146 (O_1146,N_14888,N_14706);
and UO_1147 (O_1147,N_14584,N_14578);
or UO_1148 (O_1148,N_14935,N_14327);
nor UO_1149 (O_1149,N_14522,N_14303);
and UO_1150 (O_1150,N_14831,N_14329);
nor UO_1151 (O_1151,N_14292,N_14358);
or UO_1152 (O_1152,N_14940,N_14688);
nand UO_1153 (O_1153,N_14978,N_14771);
or UO_1154 (O_1154,N_14436,N_14560);
nor UO_1155 (O_1155,N_14553,N_14514);
xor UO_1156 (O_1156,N_14536,N_14579);
or UO_1157 (O_1157,N_14807,N_14530);
nand UO_1158 (O_1158,N_14510,N_14551);
nand UO_1159 (O_1159,N_14717,N_14381);
nor UO_1160 (O_1160,N_14425,N_14311);
or UO_1161 (O_1161,N_14433,N_14480);
and UO_1162 (O_1162,N_14867,N_14849);
nor UO_1163 (O_1163,N_14332,N_14889);
and UO_1164 (O_1164,N_14416,N_14429);
nand UO_1165 (O_1165,N_14768,N_14640);
and UO_1166 (O_1166,N_14779,N_14368);
nor UO_1167 (O_1167,N_14872,N_14254);
nand UO_1168 (O_1168,N_14936,N_14653);
nand UO_1169 (O_1169,N_14527,N_14960);
xor UO_1170 (O_1170,N_14533,N_14825);
nor UO_1171 (O_1171,N_14729,N_14881);
nand UO_1172 (O_1172,N_14731,N_14490);
xnor UO_1173 (O_1173,N_14386,N_14894);
and UO_1174 (O_1174,N_14580,N_14368);
nand UO_1175 (O_1175,N_14610,N_14348);
or UO_1176 (O_1176,N_14461,N_14664);
and UO_1177 (O_1177,N_14576,N_14951);
nand UO_1178 (O_1178,N_14458,N_14413);
xor UO_1179 (O_1179,N_14475,N_14933);
nand UO_1180 (O_1180,N_14611,N_14988);
nor UO_1181 (O_1181,N_14973,N_14261);
xnor UO_1182 (O_1182,N_14532,N_14683);
nor UO_1183 (O_1183,N_14957,N_14671);
nand UO_1184 (O_1184,N_14463,N_14431);
nor UO_1185 (O_1185,N_14974,N_14773);
nor UO_1186 (O_1186,N_14916,N_14633);
or UO_1187 (O_1187,N_14978,N_14485);
nand UO_1188 (O_1188,N_14812,N_14931);
and UO_1189 (O_1189,N_14878,N_14879);
or UO_1190 (O_1190,N_14700,N_14262);
nand UO_1191 (O_1191,N_14729,N_14429);
or UO_1192 (O_1192,N_14330,N_14395);
or UO_1193 (O_1193,N_14783,N_14936);
nand UO_1194 (O_1194,N_14673,N_14312);
and UO_1195 (O_1195,N_14572,N_14536);
or UO_1196 (O_1196,N_14588,N_14895);
and UO_1197 (O_1197,N_14417,N_14366);
or UO_1198 (O_1198,N_14513,N_14461);
nand UO_1199 (O_1199,N_14895,N_14881);
and UO_1200 (O_1200,N_14351,N_14684);
nand UO_1201 (O_1201,N_14811,N_14605);
nor UO_1202 (O_1202,N_14704,N_14334);
nand UO_1203 (O_1203,N_14527,N_14342);
nor UO_1204 (O_1204,N_14868,N_14568);
and UO_1205 (O_1205,N_14320,N_14948);
nand UO_1206 (O_1206,N_14604,N_14642);
and UO_1207 (O_1207,N_14815,N_14647);
xor UO_1208 (O_1208,N_14288,N_14532);
and UO_1209 (O_1209,N_14681,N_14507);
xnor UO_1210 (O_1210,N_14411,N_14709);
nor UO_1211 (O_1211,N_14984,N_14675);
nor UO_1212 (O_1212,N_14410,N_14775);
and UO_1213 (O_1213,N_14978,N_14714);
and UO_1214 (O_1214,N_14479,N_14742);
nor UO_1215 (O_1215,N_14922,N_14953);
and UO_1216 (O_1216,N_14699,N_14463);
nor UO_1217 (O_1217,N_14261,N_14443);
and UO_1218 (O_1218,N_14306,N_14906);
or UO_1219 (O_1219,N_14537,N_14693);
nand UO_1220 (O_1220,N_14731,N_14265);
xor UO_1221 (O_1221,N_14681,N_14876);
and UO_1222 (O_1222,N_14325,N_14350);
or UO_1223 (O_1223,N_14527,N_14561);
nand UO_1224 (O_1224,N_14655,N_14974);
nor UO_1225 (O_1225,N_14458,N_14768);
nand UO_1226 (O_1226,N_14590,N_14489);
and UO_1227 (O_1227,N_14564,N_14956);
and UO_1228 (O_1228,N_14861,N_14552);
and UO_1229 (O_1229,N_14288,N_14556);
nand UO_1230 (O_1230,N_14930,N_14617);
and UO_1231 (O_1231,N_14308,N_14601);
and UO_1232 (O_1232,N_14987,N_14491);
and UO_1233 (O_1233,N_14687,N_14956);
xnor UO_1234 (O_1234,N_14537,N_14840);
nand UO_1235 (O_1235,N_14959,N_14321);
xor UO_1236 (O_1236,N_14541,N_14309);
and UO_1237 (O_1237,N_14665,N_14350);
or UO_1238 (O_1238,N_14822,N_14627);
nand UO_1239 (O_1239,N_14545,N_14322);
nand UO_1240 (O_1240,N_14804,N_14378);
or UO_1241 (O_1241,N_14307,N_14788);
or UO_1242 (O_1242,N_14281,N_14604);
or UO_1243 (O_1243,N_14615,N_14682);
nor UO_1244 (O_1244,N_14960,N_14681);
or UO_1245 (O_1245,N_14727,N_14777);
and UO_1246 (O_1246,N_14323,N_14329);
nand UO_1247 (O_1247,N_14448,N_14467);
and UO_1248 (O_1248,N_14401,N_14972);
and UO_1249 (O_1249,N_14503,N_14271);
and UO_1250 (O_1250,N_14542,N_14338);
or UO_1251 (O_1251,N_14931,N_14961);
and UO_1252 (O_1252,N_14327,N_14511);
nand UO_1253 (O_1253,N_14882,N_14888);
nand UO_1254 (O_1254,N_14352,N_14709);
xnor UO_1255 (O_1255,N_14354,N_14768);
nand UO_1256 (O_1256,N_14716,N_14800);
or UO_1257 (O_1257,N_14844,N_14985);
or UO_1258 (O_1258,N_14919,N_14986);
nand UO_1259 (O_1259,N_14803,N_14636);
and UO_1260 (O_1260,N_14535,N_14551);
and UO_1261 (O_1261,N_14489,N_14629);
and UO_1262 (O_1262,N_14644,N_14631);
nor UO_1263 (O_1263,N_14967,N_14883);
or UO_1264 (O_1264,N_14904,N_14562);
nor UO_1265 (O_1265,N_14382,N_14859);
nand UO_1266 (O_1266,N_14524,N_14632);
nand UO_1267 (O_1267,N_14342,N_14978);
or UO_1268 (O_1268,N_14659,N_14826);
xor UO_1269 (O_1269,N_14779,N_14964);
and UO_1270 (O_1270,N_14290,N_14298);
nand UO_1271 (O_1271,N_14337,N_14634);
nand UO_1272 (O_1272,N_14993,N_14994);
nand UO_1273 (O_1273,N_14612,N_14886);
or UO_1274 (O_1274,N_14608,N_14251);
nand UO_1275 (O_1275,N_14894,N_14279);
and UO_1276 (O_1276,N_14560,N_14395);
or UO_1277 (O_1277,N_14528,N_14362);
or UO_1278 (O_1278,N_14561,N_14701);
nand UO_1279 (O_1279,N_14703,N_14857);
nor UO_1280 (O_1280,N_14961,N_14992);
nor UO_1281 (O_1281,N_14530,N_14961);
nand UO_1282 (O_1282,N_14479,N_14985);
xnor UO_1283 (O_1283,N_14505,N_14397);
and UO_1284 (O_1284,N_14878,N_14925);
or UO_1285 (O_1285,N_14623,N_14803);
or UO_1286 (O_1286,N_14836,N_14944);
and UO_1287 (O_1287,N_14481,N_14269);
or UO_1288 (O_1288,N_14378,N_14345);
xor UO_1289 (O_1289,N_14430,N_14685);
and UO_1290 (O_1290,N_14462,N_14871);
nand UO_1291 (O_1291,N_14946,N_14543);
nand UO_1292 (O_1292,N_14308,N_14365);
nand UO_1293 (O_1293,N_14946,N_14762);
or UO_1294 (O_1294,N_14523,N_14807);
nor UO_1295 (O_1295,N_14794,N_14619);
nand UO_1296 (O_1296,N_14914,N_14387);
and UO_1297 (O_1297,N_14393,N_14623);
and UO_1298 (O_1298,N_14587,N_14634);
nor UO_1299 (O_1299,N_14624,N_14710);
or UO_1300 (O_1300,N_14569,N_14932);
xor UO_1301 (O_1301,N_14542,N_14883);
or UO_1302 (O_1302,N_14297,N_14812);
nand UO_1303 (O_1303,N_14566,N_14646);
or UO_1304 (O_1304,N_14702,N_14681);
and UO_1305 (O_1305,N_14337,N_14285);
and UO_1306 (O_1306,N_14419,N_14443);
nor UO_1307 (O_1307,N_14388,N_14502);
and UO_1308 (O_1308,N_14787,N_14297);
xnor UO_1309 (O_1309,N_14446,N_14526);
nor UO_1310 (O_1310,N_14562,N_14464);
nand UO_1311 (O_1311,N_14359,N_14539);
nand UO_1312 (O_1312,N_14409,N_14835);
nand UO_1313 (O_1313,N_14926,N_14765);
xor UO_1314 (O_1314,N_14771,N_14866);
and UO_1315 (O_1315,N_14633,N_14789);
nor UO_1316 (O_1316,N_14431,N_14680);
or UO_1317 (O_1317,N_14928,N_14361);
xnor UO_1318 (O_1318,N_14830,N_14887);
nand UO_1319 (O_1319,N_14434,N_14747);
nand UO_1320 (O_1320,N_14890,N_14294);
and UO_1321 (O_1321,N_14993,N_14478);
or UO_1322 (O_1322,N_14338,N_14356);
xor UO_1323 (O_1323,N_14495,N_14690);
xor UO_1324 (O_1324,N_14796,N_14394);
or UO_1325 (O_1325,N_14373,N_14370);
or UO_1326 (O_1326,N_14328,N_14950);
nor UO_1327 (O_1327,N_14348,N_14312);
nor UO_1328 (O_1328,N_14395,N_14772);
or UO_1329 (O_1329,N_14576,N_14830);
nand UO_1330 (O_1330,N_14625,N_14964);
or UO_1331 (O_1331,N_14817,N_14588);
nor UO_1332 (O_1332,N_14412,N_14826);
nand UO_1333 (O_1333,N_14298,N_14608);
nor UO_1334 (O_1334,N_14776,N_14397);
nor UO_1335 (O_1335,N_14707,N_14883);
or UO_1336 (O_1336,N_14871,N_14554);
nor UO_1337 (O_1337,N_14460,N_14681);
or UO_1338 (O_1338,N_14861,N_14960);
xnor UO_1339 (O_1339,N_14730,N_14268);
nor UO_1340 (O_1340,N_14414,N_14743);
or UO_1341 (O_1341,N_14706,N_14771);
nand UO_1342 (O_1342,N_14756,N_14832);
and UO_1343 (O_1343,N_14668,N_14350);
nor UO_1344 (O_1344,N_14404,N_14426);
and UO_1345 (O_1345,N_14932,N_14385);
nand UO_1346 (O_1346,N_14982,N_14980);
or UO_1347 (O_1347,N_14651,N_14593);
nand UO_1348 (O_1348,N_14281,N_14538);
xor UO_1349 (O_1349,N_14693,N_14531);
and UO_1350 (O_1350,N_14596,N_14573);
or UO_1351 (O_1351,N_14527,N_14994);
and UO_1352 (O_1352,N_14857,N_14935);
nand UO_1353 (O_1353,N_14823,N_14269);
nor UO_1354 (O_1354,N_14783,N_14764);
and UO_1355 (O_1355,N_14649,N_14563);
nor UO_1356 (O_1356,N_14893,N_14855);
nor UO_1357 (O_1357,N_14456,N_14756);
nand UO_1358 (O_1358,N_14420,N_14553);
nand UO_1359 (O_1359,N_14442,N_14392);
nand UO_1360 (O_1360,N_14829,N_14968);
nand UO_1361 (O_1361,N_14906,N_14298);
nor UO_1362 (O_1362,N_14923,N_14868);
and UO_1363 (O_1363,N_14366,N_14650);
or UO_1364 (O_1364,N_14796,N_14354);
nand UO_1365 (O_1365,N_14769,N_14278);
nand UO_1366 (O_1366,N_14546,N_14632);
and UO_1367 (O_1367,N_14739,N_14779);
nor UO_1368 (O_1368,N_14912,N_14584);
nand UO_1369 (O_1369,N_14479,N_14633);
or UO_1370 (O_1370,N_14303,N_14740);
or UO_1371 (O_1371,N_14411,N_14598);
xnor UO_1372 (O_1372,N_14581,N_14500);
and UO_1373 (O_1373,N_14736,N_14305);
xor UO_1374 (O_1374,N_14362,N_14705);
nand UO_1375 (O_1375,N_14742,N_14933);
and UO_1376 (O_1376,N_14914,N_14818);
and UO_1377 (O_1377,N_14419,N_14533);
nor UO_1378 (O_1378,N_14551,N_14865);
and UO_1379 (O_1379,N_14859,N_14434);
xor UO_1380 (O_1380,N_14486,N_14787);
and UO_1381 (O_1381,N_14478,N_14893);
and UO_1382 (O_1382,N_14521,N_14373);
and UO_1383 (O_1383,N_14790,N_14811);
nor UO_1384 (O_1384,N_14834,N_14920);
nor UO_1385 (O_1385,N_14730,N_14978);
nand UO_1386 (O_1386,N_14539,N_14420);
and UO_1387 (O_1387,N_14903,N_14660);
or UO_1388 (O_1388,N_14844,N_14903);
and UO_1389 (O_1389,N_14785,N_14681);
and UO_1390 (O_1390,N_14572,N_14433);
or UO_1391 (O_1391,N_14909,N_14530);
nand UO_1392 (O_1392,N_14263,N_14992);
and UO_1393 (O_1393,N_14340,N_14656);
or UO_1394 (O_1394,N_14532,N_14351);
nand UO_1395 (O_1395,N_14633,N_14963);
and UO_1396 (O_1396,N_14579,N_14841);
nand UO_1397 (O_1397,N_14401,N_14327);
nor UO_1398 (O_1398,N_14958,N_14370);
or UO_1399 (O_1399,N_14817,N_14979);
and UO_1400 (O_1400,N_14512,N_14940);
nor UO_1401 (O_1401,N_14617,N_14290);
and UO_1402 (O_1402,N_14823,N_14616);
or UO_1403 (O_1403,N_14454,N_14812);
nor UO_1404 (O_1404,N_14982,N_14856);
nand UO_1405 (O_1405,N_14462,N_14889);
or UO_1406 (O_1406,N_14708,N_14449);
nand UO_1407 (O_1407,N_14419,N_14753);
nand UO_1408 (O_1408,N_14430,N_14619);
or UO_1409 (O_1409,N_14769,N_14350);
nor UO_1410 (O_1410,N_14991,N_14606);
xnor UO_1411 (O_1411,N_14487,N_14699);
nand UO_1412 (O_1412,N_14802,N_14587);
nand UO_1413 (O_1413,N_14450,N_14517);
nand UO_1414 (O_1414,N_14920,N_14697);
and UO_1415 (O_1415,N_14325,N_14262);
nand UO_1416 (O_1416,N_14665,N_14564);
xnor UO_1417 (O_1417,N_14841,N_14668);
xor UO_1418 (O_1418,N_14833,N_14816);
nand UO_1419 (O_1419,N_14788,N_14797);
nor UO_1420 (O_1420,N_14478,N_14816);
nor UO_1421 (O_1421,N_14267,N_14907);
nand UO_1422 (O_1422,N_14583,N_14493);
or UO_1423 (O_1423,N_14377,N_14596);
nand UO_1424 (O_1424,N_14828,N_14863);
and UO_1425 (O_1425,N_14549,N_14547);
and UO_1426 (O_1426,N_14671,N_14533);
nor UO_1427 (O_1427,N_14712,N_14565);
nand UO_1428 (O_1428,N_14354,N_14647);
xor UO_1429 (O_1429,N_14414,N_14382);
and UO_1430 (O_1430,N_14685,N_14686);
and UO_1431 (O_1431,N_14802,N_14964);
nand UO_1432 (O_1432,N_14425,N_14356);
nand UO_1433 (O_1433,N_14323,N_14264);
or UO_1434 (O_1434,N_14532,N_14813);
xnor UO_1435 (O_1435,N_14299,N_14966);
and UO_1436 (O_1436,N_14262,N_14998);
nand UO_1437 (O_1437,N_14997,N_14779);
nand UO_1438 (O_1438,N_14962,N_14632);
nand UO_1439 (O_1439,N_14399,N_14686);
and UO_1440 (O_1440,N_14298,N_14653);
nor UO_1441 (O_1441,N_14323,N_14943);
or UO_1442 (O_1442,N_14961,N_14879);
nand UO_1443 (O_1443,N_14410,N_14809);
nor UO_1444 (O_1444,N_14374,N_14678);
nor UO_1445 (O_1445,N_14465,N_14503);
and UO_1446 (O_1446,N_14624,N_14436);
or UO_1447 (O_1447,N_14473,N_14692);
nand UO_1448 (O_1448,N_14703,N_14506);
nor UO_1449 (O_1449,N_14807,N_14608);
or UO_1450 (O_1450,N_14680,N_14742);
xor UO_1451 (O_1451,N_14786,N_14289);
nor UO_1452 (O_1452,N_14297,N_14423);
nand UO_1453 (O_1453,N_14981,N_14823);
nor UO_1454 (O_1454,N_14705,N_14884);
and UO_1455 (O_1455,N_14342,N_14534);
or UO_1456 (O_1456,N_14951,N_14876);
and UO_1457 (O_1457,N_14801,N_14617);
nand UO_1458 (O_1458,N_14976,N_14641);
or UO_1459 (O_1459,N_14826,N_14676);
and UO_1460 (O_1460,N_14321,N_14281);
nor UO_1461 (O_1461,N_14920,N_14760);
and UO_1462 (O_1462,N_14341,N_14363);
or UO_1463 (O_1463,N_14273,N_14975);
nor UO_1464 (O_1464,N_14621,N_14448);
nand UO_1465 (O_1465,N_14853,N_14482);
nand UO_1466 (O_1466,N_14688,N_14568);
nand UO_1467 (O_1467,N_14998,N_14520);
nand UO_1468 (O_1468,N_14699,N_14453);
xnor UO_1469 (O_1469,N_14556,N_14781);
xor UO_1470 (O_1470,N_14342,N_14688);
xor UO_1471 (O_1471,N_14629,N_14794);
nand UO_1472 (O_1472,N_14860,N_14527);
nand UO_1473 (O_1473,N_14869,N_14723);
nor UO_1474 (O_1474,N_14505,N_14306);
nor UO_1475 (O_1475,N_14374,N_14793);
and UO_1476 (O_1476,N_14517,N_14500);
and UO_1477 (O_1477,N_14904,N_14821);
and UO_1478 (O_1478,N_14826,N_14997);
and UO_1479 (O_1479,N_14760,N_14569);
nand UO_1480 (O_1480,N_14845,N_14273);
nor UO_1481 (O_1481,N_14693,N_14563);
nor UO_1482 (O_1482,N_14460,N_14612);
or UO_1483 (O_1483,N_14622,N_14434);
and UO_1484 (O_1484,N_14326,N_14488);
and UO_1485 (O_1485,N_14298,N_14780);
nand UO_1486 (O_1486,N_14905,N_14319);
and UO_1487 (O_1487,N_14891,N_14945);
nand UO_1488 (O_1488,N_14862,N_14497);
nand UO_1489 (O_1489,N_14741,N_14857);
nand UO_1490 (O_1490,N_14430,N_14576);
and UO_1491 (O_1491,N_14732,N_14498);
nand UO_1492 (O_1492,N_14767,N_14571);
nor UO_1493 (O_1493,N_14909,N_14586);
or UO_1494 (O_1494,N_14830,N_14403);
or UO_1495 (O_1495,N_14448,N_14514);
nand UO_1496 (O_1496,N_14288,N_14920);
nor UO_1497 (O_1497,N_14547,N_14741);
or UO_1498 (O_1498,N_14795,N_14977);
and UO_1499 (O_1499,N_14757,N_14541);
and UO_1500 (O_1500,N_14841,N_14989);
nand UO_1501 (O_1501,N_14361,N_14803);
nand UO_1502 (O_1502,N_14461,N_14287);
or UO_1503 (O_1503,N_14820,N_14341);
or UO_1504 (O_1504,N_14676,N_14817);
nor UO_1505 (O_1505,N_14557,N_14290);
nor UO_1506 (O_1506,N_14863,N_14836);
and UO_1507 (O_1507,N_14991,N_14494);
and UO_1508 (O_1508,N_14740,N_14616);
nand UO_1509 (O_1509,N_14366,N_14479);
and UO_1510 (O_1510,N_14577,N_14445);
xnor UO_1511 (O_1511,N_14319,N_14421);
or UO_1512 (O_1512,N_14960,N_14674);
nand UO_1513 (O_1513,N_14731,N_14586);
nand UO_1514 (O_1514,N_14626,N_14373);
or UO_1515 (O_1515,N_14560,N_14553);
nand UO_1516 (O_1516,N_14461,N_14304);
nand UO_1517 (O_1517,N_14615,N_14273);
or UO_1518 (O_1518,N_14384,N_14412);
and UO_1519 (O_1519,N_14999,N_14772);
or UO_1520 (O_1520,N_14671,N_14492);
or UO_1521 (O_1521,N_14699,N_14457);
nor UO_1522 (O_1522,N_14674,N_14503);
nor UO_1523 (O_1523,N_14401,N_14740);
or UO_1524 (O_1524,N_14831,N_14789);
or UO_1525 (O_1525,N_14456,N_14743);
or UO_1526 (O_1526,N_14629,N_14327);
or UO_1527 (O_1527,N_14741,N_14587);
nand UO_1528 (O_1528,N_14527,N_14484);
nand UO_1529 (O_1529,N_14386,N_14869);
nand UO_1530 (O_1530,N_14380,N_14754);
nand UO_1531 (O_1531,N_14345,N_14290);
nand UO_1532 (O_1532,N_14459,N_14350);
and UO_1533 (O_1533,N_14623,N_14802);
or UO_1534 (O_1534,N_14662,N_14771);
nand UO_1535 (O_1535,N_14833,N_14693);
nand UO_1536 (O_1536,N_14405,N_14402);
or UO_1537 (O_1537,N_14691,N_14270);
nor UO_1538 (O_1538,N_14721,N_14629);
xnor UO_1539 (O_1539,N_14788,N_14634);
nand UO_1540 (O_1540,N_14447,N_14974);
nand UO_1541 (O_1541,N_14349,N_14737);
or UO_1542 (O_1542,N_14428,N_14415);
nor UO_1543 (O_1543,N_14660,N_14339);
xnor UO_1544 (O_1544,N_14505,N_14482);
xor UO_1545 (O_1545,N_14386,N_14333);
xnor UO_1546 (O_1546,N_14923,N_14702);
xnor UO_1547 (O_1547,N_14476,N_14486);
and UO_1548 (O_1548,N_14891,N_14770);
and UO_1549 (O_1549,N_14333,N_14607);
nor UO_1550 (O_1550,N_14833,N_14985);
nor UO_1551 (O_1551,N_14789,N_14565);
or UO_1552 (O_1552,N_14376,N_14561);
xor UO_1553 (O_1553,N_14620,N_14710);
and UO_1554 (O_1554,N_14541,N_14430);
nand UO_1555 (O_1555,N_14296,N_14534);
or UO_1556 (O_1556,N_14890,N_14748);
nand UO_1557 (O_1557,N_14481,N_14630);
or UO_1558 (O_1558,N_14254,N_14609);
or UO_1559 (O_1559,N_14486,N_14675);
or UO_1560 (O_1560,N_14610,N_14707);
and UO_1561 (O_1561,N_14524,N_14569);
nor UO_1562 (O_1562,N_14417,N_14796);
or UO_1563 (O_1563,N_14332,N_14865);
nand UO_1564 (O_1564,N_14831,N_14878);
and UO_1565 (O_1565,N_14830,N_14634);
and UO_1566 (O_1566,N_14529,N_14389);
nor UO_1567 (O_1567,N_14848,N_14293);
nor UO_1568 (O_1568,N_14438,N_14540);
xor UO_1569 (O_1569,N_14482,N_14774);
nand UO_1570 (O_1570,N_14782,N_14928);
nand UO_1571 (O_1571,N_14563,N_14934);
nor UO_1572 (O_1572,N_14459,N_14759);
nand UO_1573 (O_1573,N_14637,N_14541);
nor UO_1574 (O_1574,N_14536,N_14997);
xnor UO_1575 (O_1575,N_14269,N_14835);
and UO_1576 (O_1576,N_14365,N_14899);
and UO_1577 (O_1577,N_14769,N_14996);
nand UO_1578 (O_1578,N_14725,N_14948);
and UO_1579 (O_1579,N_14342,N_14592);
and UO_1580 (O_1580,N_14969,N_14415);
or UO_1581 (O_1581,N_14573,N_14581);
and UO_1582 (O_1582,N_14650,N_14721);
nor UO_1583 (O_1583,N_14434,N_14641);
or UO_1584 (O_1584,N_14843,N_14768);
and UO_1585 (O_1585,N_14755,N_14332);
or UO_1586 (O_1586,N_14304,N_14603);
xnor UO_1587 (O_1587,N_14261,N_14927);
or UO_1588 (O_1588,N_14262,N_14577);
or UO_1589 (O_1589,N_14528,N_14393);
nand UO_1590 (O_1590,N_14537,N_14285);
nand UO_1591 (O_1591,N_14329,N_14613);
nand UO_1592 (O_1592,N_14483,N_14652);
nor UO_1593 (O_1593,N_14668,N_14938);
nand UO_1594 (O_1594,N_14949,N_14991);
and UO_1595 (O_1595,N_14965,N_14314);
and UO_1596 (O_1596,N_14571,N_14354);
or UO_1597 (O_1597,N_14503,N_14735);
nand UO_1598 (O_1598,N_14765,N_14662);
xnor UO_1599 (O_1599,N_14348,N_14845);
and UO_1600 (O_1600,N_14481,N_14951);
nand UO_1601 (O_1601,N_14800,N_14913);
nor UO_1602 (O_1602,N_14690,N_14878);
or UO_1603 (O_1603,N_14901,N_14914);
and UO_1604 (O_1604,N_14916,N_14703);
and UO_1605 (O_1605,N_14691,N_14412);
or UO_1606 (O_1606,N_14257,N_14333);
and UO_1607 (O_1607,N_14312,N_14687);
nor UO_1608 (O_1608,N_14870,N_14989);
xnor UO_1609 (O_1609,N_14903,N_14385);
nand UO_1610 (O_1610,N_14381,N_14395);
xor UO_1611 (O_1611,N_14431,N_14795);
and UO_1612 (O_1612,N_14832,N_14967);
nor UO_1613 (O_1613,N_14854,N_14948);
and UO_1614 (O_1614,N_14955,N_14255);
xnor UO_1615 (O_1615,N_14639,N_14806);
and UO_1616 (O_1616,N_14421,N_14392);
nand UO_1617 (O_1617,N_14833,N_14459);
nor UO_1618 (O_1618,N_14819,N_14547);
xnor UO_1619 (O_1619,N_14812,N_14943);
or UO_1620 (O_1620,N_14314,N_14719);
nand UO_1621 (O_1621,N_14346,N_14815);
nand UO_1622 (O_1622,N_14682,N_14820);
or UO_1623 (O_1623,N_14254,N_14610);
and UO_1624 (O_1624,N_14318,N_14989);
xnor UO_1625 (O_1625,N_14609,N_14805);
or UO_1626 (O_1626,N_14527,N_14334);
or UO_1627 (O_1627,N_14433,N_14674);
nor UO_1628 (O_1628,N_14609,N_14968);
and UO_1629 (O_1629,N_14340,N_14792);
nand UO_1630 (O_1630,N_14884,N_14392);
nand UO_1631 (O_1631,N_14891,N_14478);
or UO_1632 (O_1632,N_14255,N_14532);
or UO_1633 (O_1633,N_14376,N_14441);
nor UO_1634 (O_1634,N_14967,N_14539);
xor UO_1635 (O_1635,N_14347,N_14487);
nand UO_1636 (O_1636,N_14794,N_14953);
nand UO_1637 (O_1637,N_14522,N_14559);
nor UO_1638 (O_1638,N_14819,N_14579);
or UO_1639 (O_1639,N_14987,N_14824);
nand UO_1640 (O_1640,N_14449,N_14899);
xnor UO_1641 (O_1641,N_14357,N_14852);
xnor UO_1642 (O_1642,N_14772,N_14888);
and UO_1643 (O_1643,N_14440,N_14307);
nand UO_1644 (O_1644,N_14699,N_14630);
and UO_1645 (O_1645,N_14523,N_14824);
nor UO_1646 (O_1646,N_14847,N_14636);
xor UO_1647 (O_1647,N_14352,N_14411);
nand UO_1648 (O_1648,N_14617,N_14454);
nor UO_1649 (O_1649,N_14781,N_14523);
and UO_1650 (O_1650,N_14626,N_14416);
nor UO_1651 (O_1651,N_14955,N_14866);
or UO_1652 (O_1652,N_14654,N_14474);
nand UO_1653 (O_1653,N_14275,N_14726);
or UO_1654 (O_1654,N_14922,N_14859);
nor UO_1655 (O_1655,N_14362,N_14613);
nor UO_1656 (O_1656,N_14451,N_14392);
and UO_1657 (O_1657,N_14443,N_14683);
or UO_1658 (O_1658,N_14679,N_14803);
and UO_1659 (O_1659,N_14833,N_14979);
and UO_1660 (O_1660,N_14555,N_14790);
nor UO_1661 (O_1661,N_14650,N_14622);
and UO_1662 (O_1662,N_14477,N_14367);
nand UO_1663 (O_1663,N_14297,N_14759);
nand UO_1664 (O_1664,N_14296,N_14573);
nor UO_1665 (O_1665,N_14615,N_14953);
nor UO_1666 (O_1666,N_14829,N_14327);
or UO_1667 (O_1667,N_14489,N_14265);
nand UO_1668 (O_1668,N_14712,N_14587);
and UO_1669 (O_1669,N_14716,N_14317);
or UO_1670 (O_1670,N_14638,N_14738);
nor UO_1671 (O_1671,N_14935,N_14614);
or UO_1672 (O_1672,N_14745,N_14725);
and UO_1673 (O_1673,N_14397,N_14977);
and UO_1674 (O_1674,N_14671,N_14328);
or UO_1675 (O_1675,N_14826,N_14769);
and UO_1676 (O_1676,N_14755,N_14850);
and UO_1677 (O_1677,N_14732,N_14709);
nand UO_1678 (O_1678,N_14299,N_14821);
nand UO_1679 (O_1679,N_14332,N_14378);
xor UO_1680 (O_1680,N_14965,N_14460);
or UO_1681 (O_1681,N_14567,N_14302);
and UO_1682 (O_1682,N_14787,N_14312);
and UO_1683 (O_1683,N_14537,N_14878);
or UO_1684 (O_1684,N_14348,N_14597);
nand UO_1685 (O_1685,N_14654,N_14427);
nand UO_1686 (O_1686,N_14315,N_14459);
and UO_1687 (O_1687,N_14475,N_14728);
nor UO_1688 (O_1688,N_14453,N_14626);
nand UO_1689 (O_1689,N_14567,N_14381);
or UO_1690 (O_1690,N_14467,N_14358);
xor UO_1691 (O_1691,N_14336,N_14699);
and UO_1692 (O_1692,N_14515,N_14379);
nor UO_1693 (O_1693,N_14871,N_14400);
or UO_1694 (O_1694,N_14372,N_14884);
xor UO_1695 (O_1695,N_14502,N_14731);
or UO_1696 (O_1696,N_14486,N_14890);
and UO_1697 (O_1697,N_14757,N_14303);
nor UO_1698 (O_1698,N_14912,N_14430);
and UO_1699 (O_1699,N_14284,N_14890);
nor UO_1700 (O_1700,N_14330,N_14427);
and UO_1701 (O_1701,N_14474,N_14982);
or UO_1702 (O_1702,N_14381,N_14594);
nor UO_1703 (O_1703,N_14621,N_14874);
nor UO_1704 (O_1704,N_14364,N_14449);
nand UO_1705 (O_1705,N_14655,N_14877);
xor UO_1706 (O_1706,N_14263,N_14322);
nor UO_1707 (O_1707,N_14340,N_14624);
nor UO_1708 (O_1708,N_14865,N_14950);
xor UO_1709 (O_1709,N_14648,N_14647);
or UO_1710 (O_1710,N_14637,N_14847);
or UO_1711 (O_1711,N_14682,N_14579);
and UO_1712 (O_1712,N_14790,N_14749);
or UO_1713 (O_1713,N_14699,N_14840);
nor UO_1714 (O_1714,N_14250,N_14450);
and UO_1715 (O_1715,N_14712,N_14750);
xor UO_1716 (O_1716,N_14313,N_14674);
and UO_1717 (O_1717,N_14451,N_14591);
or UO_1718 (O_1718,N_14695,N_14665);
nor UO_1719 (O_1719,N_14953,N_14765);
and UO_1720 (O_1720,N_14843,N_14824);
nor UO_1721 (O_1721,N_14544,N_14740);
or UO_1722 (O_1722,N_14335,N_14569);
or UO_1723 (O_1723,N_14438,N_14713);
nor UO_1724 (O_1724,N_14612,N_14389);
nand UO_1725 (O_1725,N_14354,N_14336);
nor UO_1726 (O_1726,N_14872,N_14507);
nor UO_1727 (O_1727,N_14674,N_14522);
and UO_1728 (O_1728,N_14653,N_14942);
nand UO_1729 (O_1729,N_14809,N_14523);
xor UO_1730 (O_1730,N_14375,N_14927);
and UO_1731 (O_1731,N_14627,N_14385);
nor UO_1732 (O_1732,N_14431,N_14651);
and UO_1733 (O_1733,N_14659,N_14717);
or UO_1734 (O_1734,N_14728,N_14610);
nor UO_1735 (O_1735,N_14466,N_14525);
nor UO_1736 (O_1736,N_14438,N_14658);
nand UO_1737 (O_1737,N_14957,N_14303);
or UO_1738 (O_1738,N_14857,N_14737);
and UO_1739 (O_1739,N_14947,N_14563);
or UO_1740 (O_1740,N_14348,N_14756);
nor UO_1741 (O_1741,N_14548,N_14532);
xnor UO_1742 (O_1742,N_14976,N_14283);
nand UO_1743 (O_1743,N_14269,N_14875);
or UO_1744 (O_1744,N_14483,N_14411);
and UO_1745 (O_1745,N_14618,N_14595);
or UO_1746 (O_1746,N_14730,N_14362);
or UO_1747 (O_1747,N_14922,N_14331);
nor UO_1748 (O_1748,N_14339,N_14909);
nand UO_1749 (O_1749,N_14745,N_14923);
and UO_1750 (O_1750,N_14645,N_14530);
xnor UO_1751 (O_1751,N_14760,N_14964);
and UO_1752 (O_1752,N_14458,N_14796);
or UO_1753 (O_1753,N_14769,N_14815);
or UO_1754 (O_1754,N_14783,N_14448);
nand UO_1755 (O_1755,N_14538,N_14788);
nand UO_1756 (O_1756,N_14758,N_14686);
and UO_1757 (O_1757,N_14359,N_14644);
and UO_1758 (O_1758,N_14927,N_14493);
and UO_1759 (O_1759,N_14745,N_14440);
and UO_1760 (O_1760,N_14433,N_14560);
xor UO_1761 (O_1761,N_14760,N_14646);
nand UO_1762 (O_1762,N_14722,N_14986);
nor UO_1763 (O_1763,N_14737,N_14638);
nor UO_1764 (O_1764,N_14877,N_14907);
nand UO_1765 (O_1765,N_14920,N_14499);
nand UO_1766 (O_1766,N_14412,N_14367);
nand UO_1767 (O_1767,N_14678,N_14642);
and UO_1768 (O_1768,N_14406,N_14894);
or UO_1769 (O_1769,N_14814,N_14384);
and UO_1770 (O_1770,N_14645,N_14370);
or UO_1771 (O_1771,N_14445,N_14653);
or UO_1772 (O_1772,N_14745,N_14751);
or UO_1773 (O_1773,N_14865,N_14412);
or UO_1774 (O_1774,N_14984,N_14835);
xor UO_1775 (O_1775,N_14540,N_14437);
nand UO_1776 (O_1776,N_14581,N_14971);
nor UO_1777 (O_1777,N_14920,N_14474);
xor UO_1778 (O_1778,N_14395,N_14296);
xnor UO_1779 (O_1779,N_14424,N_14724);
nor UO_1780 (O_1780,N_14346,N_14870);
nor UO_1781 (O_1781,N_14896,N_14279);
nor UO_1782 (O_1782,N_14331,N_14927);
or UO_1783 (O_1783,N_14637,N_14921);
nand UO_1784 (O_1784,N_14613,N_14423);
nor UO_1785 (O_1785,N_14319,N_14766);
nand UO_1786 (O_1786,N_14281,N_14551);
xor UO_1787 (O_1787,N_14525,N_14842);
nor UO_1788 (O_1788,N_14992,N_14886);
and UO_1789 (O_1789,N_14524,N_14825);
nor UO_1790 (O_1790,N_14512,N_14647);
nand UO_1791 (O_1791,N_14952,N_14869);
xor UO_1792 (O_1792,N_14576,N_14497);
and UO_1793 (O_1793,N_14908,N_14512);
nor UO_1794 (O_1794,N_14473,N_14733);
nor UO_1795 (O_1795,N_14563,N_14924);
or UO_1796 (O_1796,N_14980,N_14646);
nor UO_1797 (O_1797,N_14487,N_14476);
nand UO_1798 (O_1798,N_14498,N_14938);
and UO_1799 (O_1799,N_14722,N_14299);
nand UO_1800 (O_1800,N_14847,N_14805);
or UO_1801 (O_1801,N_14509,N_14781);
and UO_1802 (O_1802,N_14868,N_14479);
xnor UO_1803 (O_1803,N_14984,N_14886);
nor UO_1804 (O_1804,N_14806,N_14894);
or UO_1805 (O_1805,N_14995,N_14572);
and UO_1806 (O_1806,N_14590,N_14635);
or UO_1807 (O_1807,N_14833,N_14814);
and UO_1808 (O_1808,N_14644,N_14500);
or UO_1809 (O_1809,N_14742,N_14463);
nand UO_1810 (O_1810,N_14919,N_14511);
and UO_1811 (O_1811,N_14666,N_14879);
or UO_1812 (O_1812,N_14622,N_14765);
nor UO_1813 (O_1813,N_14435,N_14716);
and UO_1814 (O_1814,N_14382,N_14934);
nand UO_1815 (O_1815,N_14603,N_14409);
nor UO_1816 (O_1816,N_14953,N_14362);
and UO_1817 (O_1817,N_14809,N_14573);
and UO_1818 (O_1818,N_14982,N_14650);
and UO_1819 (O_1819,N_14678,N_14810);
nand UO_1820 (O_1820,N_14923,N_14788);
or UO_1821 (O_1821,N_14515,N_14844);
or UO_1822 (O_1822,N_14761,N_14951);
and UO_1823 (O_1823,N_14743,N_14432);
nor UO_1824 (O_1824,N_14828,N_14763);
nand UO_1825 (O_1825,N_14303,N_14537);
nand UO_1826 (O_1826,N_14741,N_14804);
or UO_1827 (O_1827,N_14747,N_14899);
and UO_1828 (O_1828,N_14819,N_14277);
and UO_1829 (O_1829,N_14990,N_14963);
nand UO_1830 (O_1830,N_14905,N_14281);
nand UO_1831 (O_1831,N_14402,N_14721);
nand UO_1832 (O_1832,N_14877,N_14646);
xnor UO_1833 (O_1833,N_14432,N_14745);
or UO_1834 (O_1834,N_14560,N_14415);
or UO_1835 (O_1835,N_14686,N_14675);
nor UO_1836 (O_1836,N_14900,N_14449);
and UO_1837 (O_1837,N_14310,N_14903);
or UO_1838 (O_1838,N_14925,N_14346);
and UO_1839 (O_1839,N_14335,N_14713);
and UO_1840 (O_1840,N_14826,N_14525);
xnor UO_1841 (O_1841,N_14847,N_14298);
and UO_1842 (O_1842,N_14530,N_14923);
nand UO_1843 (O_1843,N_14985,N_14345);
xnor UO_1844 (O_1844,N_14972,N_14883);
and UO_1845 (O_1845,N_14411,N_14872);
nor UO_1846 (O_1846,N_14311,N_14736);
or UO_1847 (O_1847,N_14535,N_14576);
and UO_1848 (O_1848,N_14261,N_14849);
nand UO_1849 (O_1849,N_14449,N_14474);
xnor UO_1850 (O_1850,N_14693,N_14260);
nor UO_1851 (O_1851,N_14699,N_14818);
nand UO_1852 (O_1852,N_14926,N_14559);
nand UO_1853 (O_1853,N_14672,N_14366);
or UO_1854 (O_1854,N_14983,N_14641);
nand UO_1855 (O_1855,N_14277,N_14768);
and UO_1856 (O_1856,N_14351,N_14837);
nand UO_1857 (O_1857,N_14751,N_14970);
xor UO_1858 (O_1858,N_14630,N_14300);
and UO_1859 (O_1859,N_14620,N_14286);
or UO_1860 (O_1860,N_14575,N_14331);
or UO_1861 (O_1861,N_14897,N_14624);
xnor UO_1862 (O_1862,N_14752,N_14591);
nand UO_1863 (O_1863,N_14587,N_14646);
or UO_1864 (O_1864,N_14544,N_14975);
nand UO_1865 (O_1865,N_14362,N_14580);
or UO_1866 (O_1866,N_14558,N_14818);
nand UO_1867 (O_1867,N_14656,N_14781);
nor UO_1868 (O_1868,N_14383,N_14835);
and UO_1869 (O_1869,N_14581,N_14854);
nor UO_1870 (O_1870,N_14903,N_14695);
nor UO_1871 (O_1871,N_14259,N_14982);
nand UO_1872 (O_1872,N_14297,N_14472);
nand UO_1873 (O_1873,N_14334,N_14820);
or UO_1874 (O_1874,N_14374,N_14578);
nor UO_1875 (O_1875,N_14758,N_14308);
nand UO_1876 (O_1876,N_14616,N_14622);
xnor UO_1877 (O_1877,N_14439,N_14516);
nor UO_1878 (O_1878,N_14298,N_14792);
and UO_1879 (O_1879,N_14710,N_14576);
or UO_1880 (O_1880,N_14375,N_14971);
xor UO_1881 (O_1881,N_14467,N_14474);
and UO_1882 (O_1882,N_14761,N_14739);
or UO_1883 (O_1883,N_14563,N_14360);
or UO_1884 (O_1884,N_14318,N_14643);
nand UO_1885 (O_1885,N_14821,N_14549);
and UO_1886 (O_1886,N_14750,N_14738);
xor UO_1887 (O_1887,N_14433,N_14692);
nand UO_1888 (O_1888,N_14828,N_14856);
nand UO_1889 (O_1889,N_14908,N_14864);
nand UO_1890 (O_1890,N_14964,N_14943);
and UO_1891 (O_1891,N_14544,N_14552);
nand UO_1892 (O_1892,N_14757,N_14420);
xor UO_1893 (O_1893,N_14337,N_14635);
and UO_1894 (O_1894,N_14572,N_14589);
nand UO_1895 (O_1895,N_14621,N_14577);
nand UO_1896 (O_1896,N_14815,N_14520);
and UO_1897 (O_1897,N_14719,N_14982);
or UO_1898 (O_1898,N_14454,N_14320);
xor UO_1899 (O_1899,N_14421,N_14582);
and UO_1900 (O_1900,N_14784,N_14842);
or UO_1901 (O_1901,N_14981,N_14869);
nand UO_1902 (O_1902,N_14420,N_14599);
nand UO_1903 (O_1903,N_14406,N_14559);
nor UO_1904 (O_1904,N_14588,N_14353);
xnor UO_1905 (O_1905,N_14814,N_14658);
nor UO_1906 (O_1906,N_14531,N_14966);
nor UO_1907 (O_1907,N_14936,N_14573);
or UO_1908 (O_1908,N_14775,N_14994);
nand UO_1909 (O_1909,N_14754,N_14685);
nand UO_1910 (O_1910,N_14301,N_14362);
and UO_1911 (O_1911,N_14956,N_14598);
nand UO_1912 (O_1912,N_14755,N_14668);
nor UO_1913 (O_1913,N_14429,N_14912);
nor UO_1914 (O_1914,N_14255,N_14400);
nand UO_1915 (O_1915,N_14559,N_14635);
or UO_1916 (O_1916,N_14676,N_14619);
or UO_1917 (O_1917,N_14800,N_14934);
xor UO_1918 (O_1918,N_14986,N_14873);
nand UO_1919 (O_1919,N_14292,N_14981);
nand UO_1920 (O_1920,N_14392,N_14802);
nand UO_1921 (O_1921,N_14879,N_14276);
nor UO_1922 (O_1922,N_14703,N_14329);
or UO_1923 (O_1923,N_14379,N_14421);
or UO_1924 (O_1924,N_14561,N_14383);
nand UO_1925 (O_1925,N_14445,N_14704);
or UO_1926 (O_1926,N_14481,N_14712);
nor UO_1927 (O_1927,N_14498,N_14873);
nand UO_1928 (O_1928,N_14414,N_14943);
xnor UO_1929 (O_1929,N_14296,N_14550);
and UO_1930 (O_1930,N_14278,N_14556);
nand UO_1931 (O_1931,N_14486,N_14755);
and UO_1932 (O_1932,N_14679,N_14630);
nand UO_1933 (O_1933,N_14489,N_14698);
nand UO_1934 (O_1934,N_14390,N_14559);
nand UO_1935 (O_1935,N_14409,N_14255);
nand UO_1936 (O_1936,N_14638,N_14558);
or UO_1937 (O_1937,N_14796,N_14364);
xnor UO_1938 (O_1938,N_14936,N_14986);
nand UO_1939 (O_1939,N_14614,N_14378);
nand UO_1940 (O_1940,N_14446,N_14493);
xor UO_1941 (O_1941,N_14337,N_14783);
or UO_1942 (O_1942,N_14512,N_14502);
and UO_1943 (O_1943,N_14688,N_14826);
nor UO_1944 (O_1944,N_14499,N_14544);
nor UO_1945 (O_1945,N_14294,N_14313);
nand UO_1946 (O_1946,N_14610,N_14459);
nand UO_1947 (O_1947,N_14971,N_14673);
or UO_1948 (O_1948,N_14673,N_14436);
nand UO_1949 (O_1949,N_14265,N_14474);
or UO_1950 (O_1950,N_14746,N_14679);
nand UO_1951 (O_1951,N_14571,N_14994);
nand UO_1952 (O_1952,N_14490,N_14306);
and UO_1953 (O_1953,N_14771,N_14286);
nand UO_1954 (O_1954,N_14934,N_14826);
nand UO_1955 (O_1955,N_14853,N_14614);
nor UO_1956 (O_1956,N_14867,N_14367);
or UO_1957 (O_1957,N_14713,N_14542);
nand UO_1958 (O_1958,N_14478,N_14743);
and UO_1959 (O_1959,N_14398,N_14577);
xnor UO_1960 (O_1960,N_14317,N_14938);
and UO_1961 (O_1961,N_14407,N_14578);
nand UO_1962 (O_1962,N_14628,N_14526);
xor UO_1963 (O_1963,N_14337,N_14262);
nand UO_1964 (O_1964,N_14499,N_14314);
nor UO_1965 (O_1965,N_14939,N_14480);
nor UO_1966 (O_1966,N_14383,N_14834);
nand UO_1967 (O_1967,N_14301,N_14382);
xor UO_1968 (O_1968,N_14689,N_14859);
xnor UO_1969 (O_1969,N_14683,N_14914);
and UO_1970 (O_1970,N_14508,N_14359);
nor UO_1971 (O_1971,N_14602,N_14969);
nand UO_1972 (O_1972,N_14734,N_14340);
nand UO_1973 (O_1973,N_14437,N_14958);
or UO_1974 (O_1974,N_14407,N_14792);
or UO_1975 (O_1975,N_14723,N_14315);
nand UO_1976 (O_1976,N_14765,N_14346);
or UO_1977 (O_1977,N_14586,N_14305);
xnor UO_1978 (O_1978,N_14985,N_14618);
and UO_1979 (O_1979,N_14288,N_14401);
and UO_1980 (O_1980,N_14444,N_14926);
or UO_1981 (O_1981,N_14925,N_14549);
nor UO_1982 (O_1982,N_14689,N_14760);
nand UO_1983 (O_1983,N_14346,N_14435);
and UO_1984 (O_1984,N_14582,N_14611);
and UO_1985 (O_1985,N_14586,N_14494);
nor UO_1986 (O_1986,N_14770,N_14670);
nand UO_1987 (O_1987,N_14774,N_14513);
and UO_1988 (O_1988,N_14530,N_14732);
or UO_1989 (O_1989,N_14319,N_14389);
nand UO_1990 (O_1990,N_14351,N_14938);
nand UO_1991 (O_1991,N_14436,N_14483);
nand UO_1992 (O_1992,N_14822,N_14812);
nand UO_1993 (O_1993,N_14871,N_14256);
or UO_1994 (O_1994,N_14988,N_14779);
nand UO_1995 (O_1995,N_14460,N_14267);
and UO_1996 (O_1996,N_14965,N_14873);
nand UO_1997 (O_1997,N_14919,N_14450);
or UO_1998 (O_1998,N_14505,N_14503);
nor UO_1999 (O_1999,N_14558,N_14946);
endmodule