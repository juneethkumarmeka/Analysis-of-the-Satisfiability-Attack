module basic_2000_20000_2500_125_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
or U0 (N_0,In_1330,In_213);
xnor U1 (N_1,In_874,In_1371);
xnor U2 (N_2,In_1146,In_1586);
nand U3 (N_3,In_1410,In_47);
xnor U4 (N_4,In_236,In_442);
and U5 (N_5,In_1823,In_1312);
nand U6 (N_6,In_400,In_551);
or U7 (N_7,In_825,In_532);
xor U8 (N_8,In_307,In_1622);
nor U9 (N_9,In_416,In_877);
xnor U10 (N_10,In_61,In_564);
or U11 (N_11,In_107,In_1985);
nand U12 (N_12,In_305,In_1883);
nor U13 (N_13,In_722,In_1171);
xor U14 (N_14,In_872,In_1700);
xnor U15 (N_15,In_670,In_1188);
and U16 (N_16,In_1807,In_763);
xnor U17 (N_17,In_587,In_1096);
nor U18 (N_18,In_1671,In_46);
xnor U19 (N_19,In_477,In_113);
or U20 (N_20,In_707,In_569);
nand U21 (N_21,In_175,In_205);
nor U22 (N_22,In_1090,In_311);
xor U23 (N_23,In_1210,In_69);
and U24 (N_24,In_1655,In_382);
nor U25 (N_25,In_235,In_1944);
xor U26 (N_26,In_1429,In_507);
xor U27 (N_27,In_1556,In_94);
and U28 (N_28,In_1591,In_1157);
xnor U29 (N_29,In_162,In_263);
nor U30 (N_30,In_1027,In_844);
xnor U31 (N_31,In_278,In_942);
xor U32 (N_32,In_163,In_1943);
or U33 (N_33,In_192,In_1832);
nor U34 (N_34,In_196,In_1969);
or U35 (N_35,In_64,In_951);
xor U36 (N_36,In_464,In_1080);
nor U37 (N_37,In_989,In_1105);
nand U38 (N_38,In_1720,In_811);
xnor U39 (N_39,In_602,In_678);
nand U40 (N_40,In_1446,In_1820);
or U41 (N_41,In_1078,In_983);
and U42 (N_42,In_71,In_279);
and U43 (N_43,In_904,In_1924);
nor U44 (N_44,In_1863,In_625);
xor U45 (N_45,In_1341,In_186);
xnor U46 (N_46,In_1072,In_832);
or U47 (N_47,In_1786,In_1929);
nand U48 (N_48,In_1437,In_1136);
xor U49 (N_49,In_1884,In_1723);
and U50 (N_50,In_553,In_1672);
and U51 (N_51,In_821,In_1992);
and U52 (N_52,In_1834,In_215);
and U53 (N_53,In_1774,In_1523);
nand U54 (N_54,In_435,In_299);
or U55 (N_55,In_887,In_1397);
nor U56 (N_56,In_968,In_895);
nand U57 (N_57,In_62,In_1248);
xnor U58 (N_58,In_355,In_1558);
or U59 (N_59,In_1282,In_1030);
nor U60 (N_60,In_1901,In_706);
xnor U61 (N_61,In_1913,In_735);
and U62 (N_62,In_576,In_886);
nand U63 (N_63,In_1349,In_792);
xor U64 (N_64,In_1698,In_100);
and U65 (N_65,In_648,In_1760);
nor U66 (N_66,In_790,In_677);
nor U67 (N_67,In_1902,In_79);
nor U68 (N_68,In_1933,In_687);
nor U69 (N_69,In_1492,In_259);
nand U70 (N_70,In_1389,In_1277);
nand U71 (N_71,In_1460,In_1391);
or U72 (N_72,In_1604,In_519);
nand U73 (N_73,In_854,In_288);
and U74 (N_74,In_1579,In_191);
or U75 (N_75,In_1439,In_255);
nand U76 (N_76,In_588,In_1185);
nand U77 (N_77,In_1800,In_505);
xnor U78 (N_78,In_26,In_1721);
nand U79 (N_79,In_1173,In_549);
xor U80 (N_80,In_727,In_130);
xor U81 (N_81,In_1885,In_1704);
xnor U82 (N_82,In_1641,In_1369);
and U83 (N_83,In_53,In_1036);
or U84 (N_84,In_536,In_998);
xor U85 (N_85,In_118,In_1717);
and U86 (N_86,In_609,In_1008);
xor U87 (N_87,In_973,In_1117);
or U88 (N_88,In_33,In_226);
or U89 (N_89,In_1743,In_1051);
or U90 (N_90,In_1888,In_1861);
and U91 (N_91,In_1050,In_386);
nor U92 (N_92,In_710,In_247);
or U93 (N_93,In_1325,In_269);
xnor U94 (N_94,In_1935,In_1238);
nand U95 (N_95,In_1047,In_143);
and U96 (N_96,In_1311,In_499);
or U97 (N_97,In_1809,In_656);
xor U98 (N_98,In_1532,In_484);
nand U99 (N_99,In_132,In_1003);
nor U100 (N_100,In_672,In_27);
and U101 (N_101,In_1315,In_1142);
xnor U102 (N_102,In_1415,In_448);
nor U103 (N_103,In_622,In_1195);
xor U104 (N_104,In_744,In_879);
xnor U105 (N_105,In_1422,In_762);
nor U106 (N_106,In_662,In_1367);
nor U107 (N_107,In_1235,In_781);
nand U108 (N_108,In_227,In_104);
or U109 (N_109,In_693,In_1975);
nand U110 (N_110,In_1925,In_840);
nand U111 (N_111,In_761,In_1198);
or U112 (N_112,In_346,In_149);
nor U113 (N_113,In_356,In_675);
and U114 (N_114,In_1677,In_1320);
or U115 (N_115,In_1172,In_1515);
or U116 (N_116,In_718,In_455);
xor U117 (N_117,In_1247,In_785);
xor U118 (N_118,In_1660,In_975);
nand U119 (N_119,In_579,In_1250);
nand U120 (N_120,In_698,In_1085);
xor U121 (N_121,In_1139,In_909);
or U122 (N_122,In_1687,In_1833);
and U123 (N_123,In_1573,In_129);
nand U124 (N_124,In_1793,In_1331);
nand U125 (N_125,In_563,In_830);
or U126 (N_126,In_1756,In_1746);
xnor U127 (N_127,In_784,In_976);
and U128 (N_128,In_860,In_956);
nor U129 (N_129,In_1745,In_1890);
and U130 (N_130,In_1905,In_1652);
nor U131 (N_131,In_684,In_1847);
and U132 (N_132,In_1477,In_324);
nor U133 (N_133,In_1049,In_475);
and U134 (N_134,In_875,In_256);
xnor U135 (N_135,In_1587,In_1260);
nor U136 (N_136,In_1273,In_1919);
and U137 (N_137,In_1912,In_723);
or U138 (N_138,In_1202,In_1620);
or U139 (N_139,In_1664,In_161);
nor U140 (N_140,In_892,In_1201);
nand U141 (N_141,In_35,In_108);
or U142 (N_142,In_1358,In_804);
nor U143 (N_143,In_1264,In_908);
xnor U144 (N_144,In_521,In_266);
nand U145 (N_145,In_1661,In_1378);
or U146 (N_146,In_318,In_1827);
nor U147 (N_147,In_1728,In_1110);
nor U148 (N_148,In_1852,In_170);
nand U149 (N_149,In_357,In_506);
or U150 (N_150,In_1764,In_1947);
nand U151 (N_151,In_1091,In_1867);
nor U152 (N_152,In_1955,In_131);
and U153 (N_153,In_360,In_919);
xnor U154 (N_154,In_824,In_1896);
or U155 (N_155,In_606,In_1233);
nand U156 (N_156,In_645,In_1874);
or U157 (N_157,In_1963,In_1741);
or U158 (N_158,In_993,In_1444);
xor U159 (N_159,In_1819,In_1482);
nand U160 (N_160,In_20,N_117);
nor U161 (N_161,In_388,In_890);
or U162 (N_162,In_253,In_296);
or U163 (N_163,In_1420,N_31);
and U164 (N_164,In_485,In_1802);
nor U165 (N_165,In_1141,In_258);
nor U166 (N_166,In_316,In_831);
nor U167 (N_167,In_903,In_671);
nor U168 (N_168,N_65,In_1798);
or U169 (N_169,In_978,In_1032);
nor U170 (N_170,In_1249,In_1366);
xor U171 (N_171,In_1052,In_150);
xor U172 (N_172,In_932,In_611);
nor U173 (N_173,In_1013,In_1986);
and U174 (N_174,N_62,In_1624);
nand U175 (N_175,In_1526,N_33);
and U176 (N_176,In_1780,In_74);
nand U177 (N_177,In_425,N_30);
xnor U178 (N_178,In_565,N_113);
or U179 (N_179,N_85,In_1665);
or U180 (N_180,In_1137,In_971);
nand U181 (N_181,In_577,In_1508);
nor U182 (N_182,In_864,In_285);
xnor U183 (N_183,In_950,In_794);
xor U184 (N_184,In_1129,In_1143);
nand U185 (N_185,In_755,In_125);
nor U186 (N_186,In_812,In_1734);
and U187 (N_187,In_13,In_57);
and U188 (N_188,In_640,In_674);
and U189 (N_189,In_666,In_1594);
nand U190 (N_190,In_211,In_498);
nor U191 (N_191,In_1435,In_1528);
or U192 (N_192,In_1771,In_1368);
xor U193 (N_193,In_617,In_480);
xor U194 (N_194,In_38,In_1006);
nor U195 (N_195,In_1968,In_122);
xor U196 (N_196,In_408,In_852);
nand U197 (N_197,In_1927,In_925);
xnor U198 (N_198,In_516,In_1611);
nor U199 (N_199,In_1752,In_1855);
nand U200 (N_200,In_1033,In_148);
or U201 (N_201,In_1392,In_1295);
nand U202 (N_202,In_422,In_889);
xnor U203 (N_203,In_913,In_1064);
nand U204 (N_204,In_1633,In_51);
and U205 (N_205,N_68,In_835);
or U206 (N_206,In_1265,In_1253);
nor U207 (N_207,In_1803,In_935);
nor U208 (N_208,In_1982,N_63);
nand U209 (N_209,In_1213,In_1736);
nor U210 (N_210,In_1025,In_1093);
or U211 (N_211,In_1088,In_380);
or U212 (N_212,In_651,In_1044);
nand U213 (N_213,In_413,N_132);
nor U214 (N_214,In_1124,In_1726);
or U215 (N_215,In_1824,N_90);
and U216 (N_216,In_199,In_126);
and U217 (N_217,In_1840,In_829);
or U218 (N_218,In_598,In_1559);
nand U219 (N_219,In_1379,In_747);
xor U220 (N_220,In_1970,In_575);
and U221 (N_221,In_808,In_1191);
or U222 (N_222,N_81,In_972);
and U223 (N_223,In_1575,In_1769);
and U224 (N_224,In_847,In_702);
and U225 (N_225,In_152,N_28);
xnor U226 (N_226,N_127,In_1352);
nor U227 (N_227,In_290,N_17);
xnor U228 (N_228,In_1287,In_70);
nor U229 (N_229,In_733,In_1758);
or U230 (N_230,In_1237,In_194);
or U231 (N_231,In_1069,In_1877);
or U232 (N_232,In_159,In_451);
and U233 (N_233,In_1950,In_705);
and U234 (N_234,In_923,In_841);
nand U235 (N_235,In_749,In_1613);
xor U236 (N_236,In_271,In_433);
nor U237 (N_237,In_774,In_1267);
xor U238 (N_238,In_933,In_1791);
nand U239 (N_239,In_78,In_260);
nor U240 (N_240,In_352,In_1283);
and U241 (N_241,In_650,In_1285);
and U242 (N_242,In_1121,In_1393);
or U243 (N_243,In_1988,In_1563);
nand U244 (N_244,In_1154,In_43);
nand U245 (N_245,In_1548,N_46);
or U246 (N_246,In_1590,In_1147);
nand U247 (N_247,In_1270,In_1058);
nor U248 (N_248,In_773,In_142);
xnor U249 (N_249,In_1031,In_328);
and U250 (N_250,N_13,In_1286);
or U251 (N_251,In_655,In_696);
xnor U252 (N_252,In_466,In_428);
nor U253 (N_253,In_1015,In_1278);
xor U254 (N_254,In_751,In_766);
or U255 (N_255,In_1102,In_1386);
and U256 (N_256,In_412,In_91);
or U257 (N_257,In_396,In_503);
nor U258 (N_258,N_137,N_97);
nor U259 (N_259,In_1871,In_1469);
nand U260 (N_260,In_863,In_1513);
nand U261 (N_261,In_1406,N_22);
nor U262 (N_262,In_1221,In_1582);
xor U263 (N_263,In_1053,In_489);
nor U264 (N_264,In_341,In_1518);
xor U265 (N_265,In_1334,N_10);
xnor U266 (N_266,In_725,In_1306);
xnor U267 (N_267,In_534,In_362);
xor U268 (N_268,In_1540,In_1026);
nand U269 (N_269,In_1037,In_1327);
nand U270 (N_270,In_1070,In_504);
nor U271 (N_271,In_944,In_986);
xnor U272 (N_272,In_1068,In_712);
nor U273 (N_273,In_1075,In_293);
nor U274 (N_274,In_30,In_1243);
nand U275 (N_275,In_1360,N_26);
nor U276 (N_276,In_1848,In_1483);
nor U277 (N_277,In_742,In_239);
or U278 (N_278,In_929,In_764);
nand U279 (N_279,In_1984,In_741);
and U280 (N_280,In_1519,In_757);
or U281 (N_281,N_19,In_393);
xor U282 (N_282,N_79,In_1158);
nand U283 (N_283,In_1692,In_4);
or U284 (N_284,In_1599,In_492);
xnor U285 (N_285,N_153,In_1470);
or U286 (N_286,In_1461,In_1438);
xnor U287 (N_287,In_1502,In_1908);
and U288 (N_288,In_1733,In_560);
or U289 (N_289,In_1495,In_559);
nor U290 (N_290,In_254,In_344);
or U291 (N_291,In_658,In_850);
nand U292 (N_292,In_1667,In_780);
or U293 (N_293,In_1907,In_1380);
nor U294 (N_294,In_67,In_1066);
or U295 (N_295,In_513,In_1706);
nor U296 (N_296,In_56,In_1836);
xor U297 (N_297,In_483,In_796);
nand U298 (N_298,In_1546,In_7);
or U299 (N_299,In_488,In_421);
and U300 (N_300,In_312,In_1132);
nor U301 (N_301,In_1768,In_952);
nand U302 (N_302,In_680,In_600);
xnor U303 (N_303,In_1424,In_782);
xnor U304 (N_304,In_571,In_1356);
xor U305 (N_305,In_1845,In_189);
and U306 (N_306,In_277,In_1754);
and U307 (N_307,In_1472,In_1234);
nand U308 (N_308,In_371,In_372);
or U309 (N_309,In_714,In_691);
nand U310 (N_310,In_257,N_39);
nor U311 (N_311,In_1568,In_1281);
nand U312 (N_312,In_244,In_1595);
or U313 (N_313,In_164,In_462);
nand U314 (N_314,In_329,In_1826);
nor U315 (N_315,In_1714,In_682);
nand U316 (N_316,In_1544,N_128);
nor U317 (N_317,In_1958,In_1413);
xnor U318 (N_318,N_110,In_1615);
nor U319 (N_319,In_880,N_102);
nor U320 (N_320,In_1303,In_1092);
or U321 (N_321,In_1668,In_578);
and U322 (N_322,In_282,In_1022);
and U323 (N_323,In_898,In_1338);
xor U324 (N_324,In_144,In_326);
or U325 (N_325,N_286,In_945);
xnor U326 (N_326,In_810,In_478);
and U327 (N_327,In_430,N_266);
or U328 (N_328,In_1691,In_1453);
and U329 (N_329,In_709,In_572);
nand U330 (N_330,N_273,In_1456);
nor U331 (N_331,In_924,In_300);
xnor U332 (N_332,In_1207,In_212);
nand U333 (N_333,N_159,In_200);
xnor U334 (N_334,In_1550,In_893);
nor U335 (N_335,N_47,In_1061);
xor U336 (N_336,In_1227,In_1054);
and U337 (N_337,In_1817,In_1293);
xnor U338 (N_338,In_1416,In_1610);
or U339 (N_339,In_729,In_1631);
nand U340 (N_340,In_623,In_1099);
or U341 (N_341,N_139,In_392);
nor U342 (N_342,In_83,In_1844);
or U343 (N_343,N_61,In_1219);
nand U344 (N_344,In_1956,In_369);
xnor U345 (N_345,N_170,N_49);
nor U346 (N_346,In_121,In_1794);
or U347 (N_347,In_583,In_1294);
xnor U348 (N_348,In_268,In_1354);
or U349 (N_349,In_275,In_208);
nand U350 (N_350,In_262,In_353);
nand U351 (N_351,In_145,In_865);
nor U352 (N_352,In_988,In_97);
and U353 (N_353,In_1009,In_869);
and U354 (N_354,In_1583,In_348);
and U355 (N_355,N_167,In_866);
nor U356 (N_356,N_165,In_1875);
or U357 (N_357,N_4,In_1651);
nor U358 (N_358,In_699,In_1849);
or U359 (N_359,In_652,In_1375);
or U360 (N_360,N_299,In_1648);
nor U361 (N_361,N_29,N_250);
nor U362 (N_362,In_387,In_1108);
xnor U363 (N_363,In_1292,In_1187);
nand U364 (N_364,N_2,In_1405);
nand U365 (N_365,N_295,N_120);
and U366 (N_366,N_181,In_238);
xor U367 (N_367,In_1357,In_1384);
nand U368 (N_368,In_610,In_182);
nand U369 (N_369,In_283,N_74);
nand U370 (N_370,In_237,In_857);
or U371 (N_371,In_1814,N_230);
xor U372 (N_372,In_456,In_1178);
nor U373 (N_373,In_1252,N_80);
or U374 (N_374,N_198,In_214);
nor U375 (N_375,In_1019,In_527);
and U376 (N_376,In_814,N_103);
or U377 (N_377,In_1339,In_540);
nand U378 (N_378,N_160,In_1831);
nand U379 (N_379,In_721,N_130);
nand U380 (N_380,In_1321,In_891);
nor U381 (N_381,In_242,N_71);
xnor U382 (N_382,In_110,In_731);
xnor U383 (N_383,In_570,In_529);
and U384 (N_384,In_1788,In_1941);
nand U385 (N_385,In_302,In_246);
nor U386 (N_386,In_987,N_155);
nor U387 (N_387,In_1609,In_726);
nand U388 (N_388,In_759,In_1279);
and U389 (N_389,N_144,In_1225);
or U390 (N_390,In_541,In_29);
or U391 (N_391,In_1535,In_366);
xnor U392 (N_392,N_196,In_178);
xor U393 (N_393,In_1627,In_180);
or U394 (N_394,In_754,In_351);
and U395 (N_395,In_1347,In_1504);
or U396 (N_396,In_1906,In_1873);
and U397 (N_397,In_1464,In_3);
or U398 (N_398,In_1910,In_1634);
xnor U399 (N_399,N_253,In_470);
nand U400 (N_400,In_801,In_1696);
xor U401 (N_401,In_930,N_57);
nor U402 (N_402,In_1163,In_1936);
nand U403 (N_403,In_419,N_204);
nor U404 (N_404,In_55,In_1785);
nor U405 (N_405,In_1939,N_173);
or U406 (N_406,In_41,In_301);
and U407 (N_407,N_124,N_267);
xor U408 (N_408,In_332,In_954);
xnor U409 (N_409,In_1382,N_277);
and U410 (N_410,N_51,In_146);
xnor U411 (N_411,In_1777,N_162);
nand U412 (N_412,In_347,In_1454);
and U413 (N_413,N_177,In_1974);
xnor U414 (N_414,In_946,N_193);
and U415 (N_415,In_111,In_1792);
and U416 (N_416,In_537,In_1412);
nand U417 (N_417,In_1539,In_174);
or U418 (N_418,In_1398,In_1307);
nor U419 (N_419,In_1805,In_1928);
xnor U420 (N_420,In_1650,In_669);
nand U421 (N_421,In_660,In_1722);
and U422 (N_422,N_42,N_72);
xor U423 (N_423,In_1527,In_176);
nor U424 (N_424,In_914,In_1603);
or U425 (N_425,In_1576,In_1637);
nand U426 (N_426,In_806,In_1408);
nand U427 (N_427,In_1578,In_19);
xor U428 (N_428,In_601,In_635);
nor U429 (N_429,N_310,In_202);
nand U430 (N_430,In_123,In_1186);
xnor U431 (N_431,N_191,In_627);
xor U432 (N_432,In_1916,N_25);
nor U433 (N_433,In_1021,In_231);
nand U434 (N_434,In_719,N_43);
nand U435 (N_435,In_694,N_183);
and U436 (N_436,In_1463,In_331);
xnor U437 (N_437,In_676,In_443);
nand U438 (N_438,In_1656,In_966);
nand U439 (N_439,In_1709,In_493);
nand U440 (N_440,In_715,In_457);
or U441 (N_441,In_1783,In_1452);
and U442 (N_442,In_681,In_604);
nor U443 (N_443,In_839,In_1903);
nand U444 (N_444,In_304,In_802);
xor U445 (N_445,N_208,In_1055);
nor U446 (N_446,N_36,In_1635);
nor U447 (N_447,In_1261,In_1127);
nand U448 (N_448,In_955,In_1557);
or U449 (N_449,In_1245,N_247);
nand U450 (N_450,In_84,In_1571);
nor U451 (N_451,In_1177,In_1971);
nand U452 (N_452,In_686,In_1045);
nand U453 (N_453,N_52,In_1232);
xnor U454 (N_454,In_323,N_202);
xor U455 (N_455,In_1489,In_701);
and U456 (N_456,N_300,In_1781);
xor U457 (N_457,In_81,In_833);
and U458 (N_458,In_1640,In_964);
xor U459 (N_459,In_816,In_1776);
and U460 (N_460,In_89,In_298);
nor U461 (N_461,In_779,In_1166);
nor U462 (N_462,In_1713,In_1711);
nor U463 (N_463,N_56,In_1255);
or U464 (N_464,In_586,In_797);
nand U465 (N_465,In_151,In_1643);
nor U466 (N_466,In_1506,N_216);
and U467 (N_467,In_1256,N_206);
and U468 (N_468,In_287,In_8);
xnor U469 (N_469,In_1183,In_1160);
and U470 (N_470,In_95,In_379);
nor U471 (N_471,In_996,In_99);
nand U472 (N_472,In_1545,N_241);
nor U473 (N_473,In_1138,In_896);
nor U474 (N_474,In_697,In_700);
nand U475 (N_475,In_740,In_936);
xor U476 (N_476,In_1010,In_1301);
nand U477 (N_477,In_1481,In_902);
or U478 (N_478,In_1246,In_834);
xnor U479 (N_479,In_36,N_3);
nand U480 (N_480,In_728,In_447);
nand U481 (N_481,In_584,In_1894);
and U482 (N_482,In_1135,In_931);
and U483 (N_483,In_928,In_981);
xor U484 (N_484,In_689,In_1712);
or U485 (N_485,N_304,In_631);
xor U486 (N_486,In_272,In_1813);
nand U487 (N_487,In_858,N_218);
or U488 (N_488,In_418,N_477);
and U489 (N_489,N_303,N_399);
xor U490 (N_490,In_276,In_1104);
nand U491 (N_491,N_450,N_455);
or U492 (N_492,In_40,N_367);
nor U493 (N_493,In_1976,In_921);
or U494 (N_494,In_1866,In_730);
nor U495 (N_495,In_68,In_327);
xor U496 (N_496,In_1742,In_1296);
nor U497 (N_497,In_752,In_1612);
or U498 (N_498,In_1399,In_1123);
nand U499 (N_499,In_394,In_1980);
and U500 (N_500,In_1843,In_1617);
nor U501 (N_501,In_1772,In_1269);
nand U502 (N_502,In_668,In_1447);
nand U503 (N_503,In_1673,N_283);
nand U504 (N_504,In_1920,In_1747);
nor U505 (N_505,In_370,In_638);
xor U506 (N_506,N_444,In_1229);
nand U507 (N_507,N_265,In_1725);
and U508 (N_508,In_990,In_452);
nor U509 (N_509,In_1962,In_1216);
and U510 (N_510,In_1128,N_44);
nand U511 (N_511,In_1957,In_836);
xnor U512 (N_512,N_371,N_406);
and U513 (N_513,In_1647,In_1658);
nor U514 (N_514,In_345,N_413);
and U515 (N_515,In_753,In_112);
and U516 (N_516,In_358,In_795);
or U517 (N_517,N_0,In_9);
xor U518 (N_518,N_9,N_445);
nand U519 (N_519,N_420,In_402);
nand U520 (N_520,In_1775,N_462);
and U521 (N_521,In_1196,In_938);
nand U522 (N_522,N_306,In_1695);
and U523 (N_523,In_756,In_736);
nor U524 (N_524,In_767,N_467);
or U525 (N_525,In_1165,In_629);
or U526 (N_526,In_711,In_947);
and U527 (N_527,In_1681,In_1782);
xnor U528 (N_528,In_141,In_1948);
or U529 (N_529,In_1815,N_302);
nand U530 (N_530,N_232,In_1636);
nor U531 (N_531,In_1959,N_365);
nor U532 (N_532,In_1934,In_1194);
nand U533 (N_533,In_1459,In_1915);
nand U534 (N_534,In_1787,In_593);
nand U535 (N_535,In_1205,In_1676);
or U536 (N_536,In_1753,In_732);
nor U537 (N_537,In_411,N_293);
nand U538 (N_538,In_1383,In_1638);
or U539 (N_539,In_491,In_1870);
nor U540 (N_540,In_1395,In_218);
nand U541 (N_541,N_339,In_1914);
nand U542 (N_542,In_446,N_240);
xnor U543 (N_543,In_1520,In_39);
or U544 (N_544,In_1329,In_1569);
and U545 (N_545,In_1589,N_18);
nor U546 (N_546,N_15,In_770);
xnor U547 (N_547,In_167,In_241);
and U548 (N_548,N_425,In_11);
and U549 (N_549,In_1744,In_1895);
nor U550 (N_550,In_1176,In_1155);
xor U551 (N_551,In_1280,In_1811);
and U552 (N_552,N_332,N_386);
nand U553 (N_553,In_827,N_368);
or U554 (N_554,N_64,In_1474);
and U555 (N_555,N_145,In_1512);
and U556 (N_556,N_176,In_375);
and U557 (N_557,N_147,N_391);
xor U558 (N_558,In_1226,In_1494);
nand U559 (N_559,In_373,In_45);
xnor U560 (N_560,In_1621,In_1654);
nor U561 (N_561,N_14,In_1731);
nor U562 (N_562,In_1449,In_173);
nor U563 (N_563,In_878,In_403);
xor U564 (N_564,N_379,In_1841);
nand U565 (N_565,In_1039,N_190);
nor U566 (N_566,In_1868,In_166);
and U567 (N_567,In_15,In_1362);
nor U568 (N_568,In_384,In_1946);
or U569 (N_569,In_1973,In_934);
and U570 (N_570,In_140,In_1000);
xor U571 (N_571,In_1922,In_1266);
xnor U572 (N_572,In_22,In_1231);
nor U573 (N_573,In_616,In_1584);
xnor U574 (N_574,In_1659,In_1426);
and U575 (N_575,In_557,N_470);
nand U576 (N_576,In_1442,In_545);
and U577 (N_577,N_219,In_1680);
or U578 (N_578,In_482,In_859);
nand U579 (N_579,In_525,N_205);
nor U580 (N_580,N_284,In_90);
and U581 (N_581,N_308,In_817);
xor U582 (N_582,In_1263,In_171);
and U583 (N_583,N_393,In_1608);
or U584 (N_584,N_305,In_284);
nor U585 (N_585,In_1997,N_449);
xor U586 (N_586,In_995,In_1275);
nand U587 (N_587,N_93,In_800);
nand U588 (N_588,In_1799,In_605);
nand U589 (N_589,In_1904,N_272);
or U590 (N_590,In_1730,N_7);
nor U591 (N_591,In_1738,In_538);
nor U592 (N_592,In_280,In_376);
nand U593 (N_593,N_422,In_1041);
xnor U594 (N_594,In_1268,N_118);
nor U595 (N_595,N_149,In_391);
or U596 (N_596,In_937,In_87);
or U597 (N_597,In_1020,In_1309);
nand U598 (N_598,In_552,N_161);
xor U599 (N_599,In_1364,In_169);
or U600 (N_600,In_963,In_980);
nor U601 (N_601,N_236,In_303);
and U602 (N_602,In_1324,In_21);
or U603 (N_603,In_103,N_126);
xnor U604 (N_604,N_475,In_531);
nand U605 (N_605,N_148,In_905);
xor U606 (N_606,N_428,In_1450);
nand U607 (N_607,In_1467,In_426);
and U608 (N_608,In_190,In_984);
and U609 (N_609,In_1120,N_435);
and U610 (N_610,In_1373,In_1626);
and U611 (N_611,In_508,In_1350);
or U612 (N_612,In_630,In_580);
nor U613 (N_613,In_317,In_1242);
or U614 (N_614,In_297,In_1909);
xor U615 (N_615,In_618,In_1778);
and U616 (N_616,In_1476,In_322);
nor U617 (N_617,In_50,In_471);
and U618 (N_618,N_188,In_1345);
and U619 (N_619,In_820,In_962);
xor U620 (N_620,N_439,N_89);
or U621 (N_621,N_23,N_201);
nand U622 (N_622,In_803,In_1271);
nand U623 (N_623,In_1118,In_155);
and U624 (N_624,In_685,N_281);
xnor U625 (N_625,In_265,In_1486);
xor U626 (N_626,In_1153,N_20);
nand U627 (N_627,In_406,N_75);
and U628 (N_628,In_1887,In_1299);
or U629 (N_629,In_1067,N_382);
and U630 (N_630,In_1510,In_1812);
nor U631 (N_631,N_307,N_327);
nor U632 (N_632,N_83,N_217);
nand U633 (N_633,In_1522,In_1701);
nor U634 (N_634,N_98,In_224);
xnor U635 (N_635,In_556,In_168);
nor U636 (N_636,In_337,N_334);
nor U637 (N_637,In_308,In_1732);
xor U638 (N_638,N_134,In_615);
nor U639 (N_639,In_1175,In_562);
and U640 (N_640,N_12,N_336);
nor U641 (N_641,In_642,In_1821);
nor U642 (N_642,In_1200,In_867);
or U643 (N_643,In_294,In_459);
nor U644 (N_644,In_665,N_483);
or U645 (N_645,In_1942,N_199);
or U646 (N_646,In_926,N_572);
and U647 (N_647,In_1945,N_194);
xnor U648 (N_648,N_333,In_1179);
xor U649 (N_649,N_600,N_184);
nand U650 (N_650,In_743,In_1071);
and U651 (N_651,In_28,N_469);
and U652 (N_652,In_1086,N_164);
or U653 (N_653,In_1431,N_233);
xor U654 (N_654,In_1430,In_395);
nand U655 (N_655,In_894,In_1001);
and U656 (N_656,N_442,In_368);
nor U657 (N_657,N_260,N_40);
xnor U658 (N_658,N_41,In_815);
or U659 (N_659,N_583,N_588);
or U660 (N_660,In_734,In_1002);
and U661 (N_661,In_799,In_381);
and U662 (N_662,In_1115,In_982);
or U663 (N_663,In_185,N_541);
nor U664 (N_664,In_1872,In_1710);
or U665 (N_665,N_21,N_374);
and U666 (N_666,In_1018,N_11);
nand U667 (N_667,N_261,N_294);
nand U668 (N_668,N_639,In_476);
or U669 (N_669,In_1100,In_1122);
xor U670 (N_670,N_466,In_1116);
xnor U671 (N_671,In_1119,In_243);
nand U672 (N_672,In_1521,N_604);
xor U673 (N_673,In_568,In_1524);
xnor U674 (N_674,N_27,In_910);
nor U675 (N_675,In_1674,In_124);
xor U676 (N_676,In_1374,N_168);
and U677 (N_677,In_1663,N_625);
nand U678 (N_678,In_1983,In_941);
nor U679 (N_679,N_316,N_372);
nor U680 (N_680,In_1485,In_1062);
and U681 (N_681,In_528,In_1581);
nand U682 (N_682,In_1825,In_229);
or U683 (N_683,N_528,N_131);
nand U684 (N_684,N_481,N_389);
nand U685 (N_685,In_1588,In_885);
or U686 (N_686,In_1662,N_92);
xnor U687 (N_687,N_195,In_788);
nand U688 (N_688,In_92,In_210);
or U689 (N_689,N_141,In_250);
and U690 (N_690,N_387,In_916);
xor U691 (N_691,In_1425,N_395);
nand U692 (N_692,In_1496,In_509);
nor U693 (N_693,In_965,In_1387);
or U694 (N_694,N_585,N_511);
and U695 (N_695,N_624,In_1562);
xor U696 (N_696,N_494,In_901);
xor U697 (N_697,In_458,N_256);
nand U698 (N_698,N_359,In_1547);
xnor U699 (N_699,In_1770,In_1666);
or U700 (N_700,In_334,N_559);
nand U701 (N_701,In_991,In_1079);
nor U702 (N_702,In_1317,N_566);
nand U703 (N_703,N_239,N_419);
or U704 (N_704,N_486,In_1114);
xor U705 (N_705,N_433,N_58);
or U706 (N_706,In_819,N_325);
nor U707 (N_707,In_1083,In_523);
and U708 (N_708,In_807,N_319);
nor U709 (N_709,In_439,N_479);
xor U710 (N_710,N_610,In_1284);
or U711 (N_711,N_213,In_1365);
or U712 (N_712,N_321,N_275);
and U713 (N_713,In_849,N_622);
or U714 (N_714,In_106,In_1705);
or U715 (N_715,N_558,In_1288);
and U716 (N_716,In_1065,N_431);
or U717 (N_717,In_1029,N_353);
nor U718 (N_718,N_513,In_468);
nor U719 (N_719,N_109,N_104);
nor U720 (N_720,N_313,N_620);
xor U721 (N_721,In_1966,In_1407);
xnor U722 (N_722,In_884,N_457);
nand U723 (N_723,In_787,In_585);
nor U724 (N_724,N_381,In_116);
or U725 (N_725,In_659,In_1298);
nor U726 (N_726,In_851,In_1750);
or U727 (N_727,In_1319,In_82);
nor U728 (N_728,In_494,In_1762);
and U729 (N_729,N_492,In_1862);
and U730 (N_730,In_138,N_581);
nand U731 (N_731,In_1653,N_552);
xor U732 (N_732,In_1272,In_1333);
nor U733 (N_733,N_515,N_257);
or U734 (N_734,In_1343,In_1719);
xnor U735 (N_735,N_554,N_106);
nor U736 (N_736,N_326,N_289);
nor U737 (N_737,In_1503,In_628);
nor U738 (N_738,N_502,N_591);
or U739 (N_739,In_626,N_516);
and U740 (N_740,In_1223,N_209);
nor U741 (N_741,In_1103,In_1432);
nand U742 (N_742,In_354,N_557);
and U743 (N_743,N_115,In_1570);
nor U744 (N_744,N_478,In_1418);
and U745 (N_745,N_278,In_769);
nand U746 (N_746,In_1977,In_17);
nand U747 (N_747,N_448,In_1328);
and U748 (N_748,In_713,In_695);
nand U749 (N_749,In_473,In_1487);
and U750 (N_750,In_957,N_567);
or U751 (N_751,N_565,N_630);
xnor U752 (N_752,In_550,In_673);
or U753 (N_753,In_899,N_54);
xor U754 (N_754,N_322,In_1197);
and U755 (N_755,N_112,In_1965);
nand U756 (N_756,In_1505,In_646);
or U757 (N_757,In_1434,In_1657);
nor U758 (N_758,In_306,In_1276);
nor U759 (N_759,In_1490,N_551);
and U760 (N_760,In_637,In_592);
xnor U761 (N_761,N_50,N_225);
xor U762 (N_762,N_531,N_129);
and U763 (N_763,In_415,N_174);
nor U764 (N_764,In_1181,In_1297);
nor U765 (N_765,N_599,In_856);
xor U766 (N_766,N_519,In_1625);
or U767 (N_767,N_355,In_1729);
or U768 (N_768,In_643,N_618);
xor U769 (N_769,In_267,In_1209);
nor U770 (N_770,In_139,In_1332);
xor U771 (N_771,In_204,N_635);
or U772 (N_772,In_939,In_720);
or U773 (N_773,In_1801,In_1789);
and U774 (N_774,N_571,N_347);
nand U775 (N_775,In_1184,N_601);
nand U776 (N_776,In_157,In_1289);
nor U777 (N_777,N_520,N_311);
or U778 (N_778,In_1530,In_1308);
and U779 (N_779,In_1007,N_627);
xnor U780 (N_780,N_187,In_1372);
or U781 (N_781,In_460,N_345);
nand U782 (N_782,N_463,In_1411);
nor U783 (N_783,N_222,In_206);
and U784 (N_784,In_1865,N_53);
xor U785 (N_785,N_242,In_739);
nor U786 (N_786,In_1618,N_99);
xor U787 (N_787,In_1214,In_1538);
nor U788 (N_788,N_612,In_1552);
and U789 (N_789,N_621,In_209);
xor U790 (N_790,N_166,In_1856);
nand U791 (N_791,N_545,N_227);
and U792 (N_792,In_405,In_342);
and U793 (N_793,In_1323,In_343);
xnor U794 (N_794,N_221,In_154);
or U795 (N_795,In_1159,In_58);
or U796 (N_796,N_111,In_1854);
xor U797 (N_797,N_421,N_497);
and U798 (N_798,N_34,In_548);
nand U799 (N_799,In_1274,In_1930);
nor U800 (N_800,In_813,N_453);
and U801 (N_801,In_437,In_1314);
xor U802 (N_802,N_291,N_349);
xnor U803 (N_803,In_649,In_1107);
or U804 (N_804,In_216,In_1858);
nand U805 (N_805,In_1536,In_599);
or U806 (N_806,N_268,N_95);
and U807 (N_807,N_361,In_1466);
nor U808 (N_808,In_1757,In_883);
or U809 (N_809,N_154,N_417);
or U810 (N_810,In_313,N_487);
nand U811 (N_811,In_1224,In_1342);
xor U812 (N_812,N_203,In_1074);
or U813 (N_813,In_5,In_137);
or U814 (N_814,In_1755,In_561);
or U815 (N_815,N_763,In_1838);
xnor U816 (N_816,In_940,In_1012);
and U817 (N_817,N_683,N_269);
nand U818 (N_818,In_25,In_985);
or U819 (N_819,N_335,In_777);
nor U820 (N_820,N_650,In_248);
or U821 (N_821,In_1244,In_474);
xnor U822 (N_822,In_871,N_580);
nand U823 (N_823,In_1860,In_1685);
or U824 (N_824,N_197,N_726);
and U825 (N_825,N_136,In_1363);
or U826 (N_826,N_709,In_52);
nand U827 (N_827,N_358,In_805);
nor U828 (N_828,N_312,In_596);
and U829 (N_829,N_375,In_349);
or U830 (N_830,In_486,In_1468);
xor U831 (N_831,In_1839,In_1377);
or U832 (N_832,N_667,In_690);
nand U833 (N_833,In_1322,In_181);
nand U834 (N_834,In_264,In_310);
or U835 (N_835,N_180,N_443);
xor U836 (N_836,N_721,N_533);
nor U837 (N_837,In_245,In_73);
nor U838 (N_838,In_1999,In_1529);
xnor U839 (N_839,In_1642,In_708);
nand U840 (N_840,In_117,N_480);
nand U841 (N_841,In_862,In_1835);
xor U842 (N_842,N_186,In_431);
nand U843 (N_843,In_1125,N_171);
or U844 (N_844,In_911,In_249);
or U845 (N_845,N_1,N_649);
or U846 (N_846,In_518,In_786);
xor U847 (N_847,In_1126,N_351);
or U848 (N_848,In_85,N_276);
and U849 (N_849,In_63,In_1451);
nor U850 (N_850,N_671,In_1953);
nand U851 (N_851,In_158,N_514);
xnor U852 (N_852,N_179,In_160);
xor U853 (N_853,N_771,In_1702);
nand U854 (N_854,In_1669,N_737);
or U855 (N_855,N_799,In_399);
or U856 (N_856,In_321,In_1023);
nor U857 (N_857,In_1829,In_1427);
nor U858 (N_858,N_563,In_1967);
nor U859 (N_859,In_566,N_673);
nor U860 (N_860,In_1560,N_133);
or U861 (N_861,N_546,In_1869);
nor U862 (N_862,In_1131,N_77);
or U863 (N_863,In_1645,N_679);
or U864 (N_864,N_638,N_138);
and U865 (N_865,N_156,In_1979);
nand U866 (N_866,In_1580,N_681);
nand U867 (N_867,In_1215,N_632);
or U868 (N_868,In_724,N_343);
xnor U869 (N_869,In_490,N_754);
xnor U870 (N_870,In_661,In_1152);
and U871 (N_871,In_843,In_1212);
and U872 (N_872,N_765,N_452);
nor U873 (N_873,N_593,In_619);
nand U874 (N_874,In_539,N_398);
or U875 (N_875,In_1404,In_1751);
nand U876 (N_876,N_728,N_55);
or U877 (N_877,In_1340,In_1455);
or U878 (N_878,In_501,In_1300);
nor U879 (N_879,N_636,N_608);
or U880 (N_880,N_254,In_1735);
nor U881 (N_881,In_1850,N_529);
nor U882 (N_882,In_1952,N_730);
or U883 (N_883,In_512,In_1228);
nor U884 (N_884,N_86,N_676);
xnor U885 (N_885,In_1911,N_489);
nand U886 (N_886,In_1564,In_1779);
nor U887 (N_887,In_1940,In_918);
nor U888 (N_888,In_1938,In_543);
or U889 (N_889,In_1690,In_1304);
and U890 (N_890,N_175,In_594);
nand U891 (N_891,In_1222,N_5);
and U892 (N_892,In_1134,N_495);
and U893 (N_893,N_747,N_693);
nor U894 (N_894,N_716,In_1937);
and U895 (N_895,N_318,In_330);
xor U896 (N_896,In_65,N_748);
nor U897 (N_897,N_556,In_912);
and U898 (N_898,N_354,In_526);
or U899 (N_899,N_430,N_776);
or U900 (N_900,N_505,N_340);
nor U901 (N_901,N_555,N_611);
nand U902 (N_902,In_1818,N_701);
and U903 (N_903,N_69,In_1361);
nor U904 (N_904,In_1565,In_1168);
and U905 (N_905,N_647,N_568);
xnor U906 (N_906,N_424,N_248);
or U907 (N_907,In_228,N_666);
nor U908 (N_908,N_669,N_290);
or U909 (N_909,In_1057,N_587);
nand U910 (N_910,In_389,N_710);
and U911 (N_911,N_509,N_140);
or U912 (N_912,In_496,In_42);
or U913 (N_913,In_1491,In_1257);
nand U914 (N_914,N_508,In_1739);
nor U915 (N_915,N_677,N_562);
nand U916 (N_916,N_735,In_153);
nand U917 (N_917,In_1156,In_1898);
and U918 (N_918,In_1011,N_607);
and U919 (N_919,N_338,In_1891);
and U920 (N_920,N_782,In_949);
nand U921 (N_921,N_579,In_60);
and U922 (N_922,In_1795,In_1462);
and U923 (N_923,In_481,In_49);
or U924 (N_924,N_792,In_522);
nor U925 (N_925,In_1682,In_1727);
nand U926 (N_926,In_737,In_1089);
nand U927 (N_927,N_797,N_341);
nand U928 (N_928,In_289,N_569);
nor U929 (N_929,In_500,In_1436);
nand U930 (N_930,N_507,In_608);
xnor U931 (N_931,In_621,In_1593);
nand U932 (N_932,N_298,In_1414);
nor U933 (N_933,In_1063,N_76);
and U934 (N_934,In_1335,N_656);
nand U935 (N_935,N_643,In_434);
and U936 (N_936,N_369,In_1876);
xor U937 (N_937,N_252,N_576);
or U938 (N_938,In_365,In_93);
nor U939 (N_939,N_770,N_540);
nand U940 (N_940,N_691,In_1561);
and U941 (N_941,N_534,In_390);
xnor U942 (N_942,In_581,In_251);
or U943 (N_943,N_223,N_394);
or U944 (N_944,In_1443,In_633);
nand U945 (N_945,N_214,N_688);
and U946 (N_946,In_232,In_589);
and U947 (N_947,In_1402,N_228);
nor U948 (N_948,In_1501,N_758);
nor U949 (N_949,In_463,In_414);
and U950 (N_950,In_634,In_1497);
or U951 (N_951,In_1258,N_527);
nand U952 (N_952,In_967,In_445);
nor U953 (N_953,N_329,In_1989);
and U954 (N_954,In_992,In_80);
or U955 (N_955,N_207,N_518);
xnor U956 (N_956,N_561,N_397);
nand U957 (N_957,In_12,In_1081);
and U958 (N_958,In_1600,N_684);
or U959 (N_959,N_651,In_98);
xor U960 (N_960,In_240,In_424);
or U961 (N_961,In_1094,N_323);
and U962 (N_962,N_388,N_670);
xnor U963 (N_963,N_658,In_1864);
nor U964 (N_964,N_390,In_1098);
or U965 (N_965,In_1199,In_1889);
and U966 (N_966,N_408,N_919);
xnor U967 (N_967,In_1113,In_1511);
and U968 (N_968,In_1828,In_1993);
xor U969 (N_969,N_414,In_1555);
or U970 (N_970,N_504,N_654);
nand U971 (N_971,In_614,N_337);
and U972 (N_972,N_496,In_1886);
nand U973 (N_973,N_70,N_315);
xnor U974 (N_974,In_101,In_959);
or U975 (N_975,In_510,N_434);
or U976 (N_976,In_440,N_885);
nor U977 (N_977,In_1707,In_32);
nor U978 (N_978,N_659,In_544);
nand U979 (N_979,N_614,N_835);
or U980 (N_980,In_1797,In_647);
and U981 (N_981,In_1106,In_156);
and U982 (N_982,In_120,N_549);
nand U983 (N_983,In_1409,N_824);
nor U984 (N_984,N_853,N_48);
nand U985 (N_985,In_530,N_192);
or U986 (N_986,In_1290,In_1046);
nand U987 (N_987,N_59,N_617);
xnor U988 (N_988,N_766,N_949);
nand U989 (N_989,In_582,In_1773);
xnor U990 (N_990,N_476,N_818);
nand U991 (N_991,In_958,In_846);
xor U992 (N_992,N_957,In_1954);
or U993 (N_993,N_740,In_72);
and U994 (N_994,N_767,N_403);
nand U995 (N_995,N_350,N_953);
nor U996 (N_996,In_1087,N_88);
nand U997 (N_997,N_786,N_809);
nor U998 (N_998,In_745,In_542);
and U999 (N_999,In_1541,N_823);
and U1000 (N_1000,In_497,In_350);
and U1001 (N_1001,N_689,In_558);
xnor U1002 (N_1002,In_636,N_723);
nor U1003 (N_1003,In_320,N_764);
xnor U1004 (N_1004,N_734,N_530);
xnor U1005 (N_1005,In_1262,N_863);
nor U1006 (N_1006,N_887,N_959);
nand U1007 (N_1007,N_718,N_906);
nor U1008 (N_1008,N_742,N_143);
xnor U1009 (N_1009,N_852,In_404);
nand U1010 (N_1010,N_772,In_1370);
nand U1011 (N_1011,In_1167,In_193);
and U1012 (N_1012,N_928,In_823);
and U1013 (N_1013,In_1543,In_502);
xor U1014 (N_1014,N_682,In_1140);
and U1015 (N_1015,In_472,In_915);
nand U1016 (N_1016,In_664,N_785);
and U1017 (N_1017,In_997,N_623);
nor U1018 (N_1018,In_818,In_1310);
and U1019 (N_1019,N_804,N_897);
xnor U1020 (N_1020,In_778,In_1790);
nor U1021 (N_1021,N_930,In_385);
nor U1022 (N_1022,N_465,N_934);
and U1023 (N_1023,In_644,In_1471);
and U1024 (N_1024,In_667,N_182);
nand U1025 (N_1025,In_1597,N_761);
and U1026 (N_1026,N_810,N_921);
nor U1027 (N_1027,In_775,In_1017);
nand U1028 (N_1028,N_902,In_1241);
or U1029 (N_1029,N_157,In_333);
nor U1030 (N_1030,In_1084,N_285);
xnor U1031 (N_1031,In_603,N_814);
nor U1032 (N_1032,N_237,N_698);
and U1033 (N_1033,In_1348,N_699);
or U1034 (N_1034,N_947,In_1151);
and U1035 (N_1035,In_1689,N_523);
xor U1036 (N_1036,In_1457,N_401);
and U1037 (N_1037,In_1145,In_223);
nand U1038 (N_1038,In_1161,In_66);
and U1039 (N_1039,In_612,N_342);
and U1040 (N_1040,N_101,In_873);
and U1041 (N_1041,N_105,In_760);
xor U1042 (N_1042,N_447,N_842);
nand U1043 (N_1043,N_641,In_927);
or U1044 (N_1044,N_226,N_700);
and U1045 (N_1045,In_772,In_1390);
xor U1046 (N_1046,In_1484,N_648);
and U1047 (N_1047,N_8,In_1607);
nor U1048 (N_1048,In_922,In_172);
xor U1049 (N_1049,N_605,N_843);
nor U1050 (N_1050,In_1353,In_1337);
and U1051 (N_1051,N_107,N_499);
and U1052 (N_1052,N_731,N_665);
or U1053 (N_1053,N_330,In_1111);
nor U1054 (N_1054,In_273,N_883);
xnor U1055 (N_1055,N_526,In_1554);
and U1056 (N_1056,In_1077,In_1994);
xor U1057 (N_1057,N_596,N_352);
or U1058 (N_1058,In_688,N_759);
nand U1059 (N_1059,N_158,N_459);
or U1060 (N_1060,N_733,In_76);
nor U1061 (N_1061,N_871,In_274);
and U1062 (N_1062,In_1060,N_774);
and U1063 (N_1063,N_695,N_803);
nand U1064 (N_1064,In_1995,In_1480);
nand U1065 (N_1065,In_479,In_1897);
and U1066 (N_1066,N_172,N_813);
and U1067 (N_1067,In_683,In_1763);
nor U1068 (N_1068,In_515,In_219);
and U1069 (N_1069,In_1808,N_801);
and U1070 (N_1070,N_855,N_503);
nand U1071 (N_1071,N_745,N_441);
nor U1072 (N_1072,In_1169,N_660);
nor U1073 (N_1073,N_151,In_574);
or U1074 (N_1074,In_692,N_807);
nor U1075 (N_1075,N_901,N_907);
nor U1076 (N_1076,In_1949,N_829);
xor U1077 (N_1077,In_1619,In_1193);
and U1078 (N_1078,In_1981,N_595);
nand U1079 (N_1079,In_336,N_954);
nor U1080 (N_1080,N_60,In_401);
or U1081 (N_1081,N_380,N_616);
nand U1082 (N_1082,N_460,In_917);
nand U1083 (N_1083,N_560,N_750);
or U1084 (N_1084,N_410,N_923);
and U1085 (N_1085,In_292,In_377);
nand U1086 (N_1086,N_461,N_950);
xor U1087 (N_1087,In_14,In_1961);
xnor U1088 (N_1088,In_1623,In_135);
nor U1089 (N_1089,N_517,In_868);
nand U1090 (N_1090,N_35,N_736);
and U1091 (N_1091,In_1170,N_270);
nor U1092 (N_1092,N_933,In_102);
nand U1093 (N_1093,In_1693,In_1164);
and U1094 (N_1094,In_994,In_217);
nand U1095 (N_1095,In_1182,N_851);
or U1096 (N_1096,In_1498,N_899);
nand U1097 (N_1097,In_1240,In_1740);
nor U1098 (N_1098,N_697,N_224);
nand U1099 (N_1099,In_1388,In_1830);
nor U1100 (N_1100,N_500,N_784);
and U1101 (N_1101,In_567,N_762);
or U1102 (N_1102,N_790,N_836);
and U1103 (N_1103,In_876,N_672);
xnor U1104 (N_1104,N_416,N_909);
nand U1105 (N_1105,N_633,N_751);
nand U1106 (N_1106,In_465,N_246);
or U1107 (N_1107,In_1991,N_780);
nor U1108 (N_1108,In_663,N_932);
xor U1109 (N_1109,In_1880,In_1542);
or U1110 (N_1110,N_215,N_38);
or U1111 (N_1111,N_895,In_221);
xnor U1112 (N_1112,N_210,In_1109);
or U1113 (N_1113,In_136,In_639);
xnor U1114 (N_1114,In_1759,In_361);
xnor U1115 (N_1115,N_423,In_855);
nand U1116 (N_1116,In_1718,N_945);
nand U1117 (N_1117,N_429,N_749);
and U1118 (N_1118,In_595,In_953);
xor U1119 (N_1119,N_822,N_282);
and U1120 (N_1120,N_211,In_198);
or U1121 (N_1121,N_1037,N_411);
xnor U1122 (N_1122,N_314,N_637);
xnor U1123 (N_1123,In_1421,In_220);
xor U1124 (N_1124,N_402,N_521);
xnor U1125 (N_1125,In_1931,N_150);
nand U1126 (N_1126,In_363,N_910);
and U1127 (N_1127,N_816,N_722);
nand U1128 (N_1128,N_45,N_916);
and U1129 (N_1129,N_287,N_1115);
and U1130 (N_1130,N_490,In_1203);
nor U1131 (N_1131,N_839,In_590);
or U1132 (N_1132,N_493,N_831);
or U1133 (N_1133,In_1900,In_261);
xor U1134 (N_1134,In_960,In_776);
or U1135 (N_1135,In_340,N_244);
nor U1136 (N_1136,In_717,N_805);
xor U1137 (N_1137,N_685,In_1574);
nor U1138 (N_1138,In_1479,N_898);
nor U1139 (N_1139,In_613,In_828);
nand U1140 (N_1140,N_781,N_727);
nor U1141 (N_1141,N_1038,N_862);
and U1142 (N_1142,N_255,N_1021);
nand U1143 (N_1143,N_82,N_834);
nor U1144 (N_1144,In_838,N_1106);
or U1145 (N_1145,N_968,In_444);
nand U1146 (N_1146,N_32,In_554);
nand U1147 (N_1147,In_555,In_1796);
nor U1148 (N_1148,In_295,In_119);
nor U1149 (N_1149,N_1043,N_830);
or U1150 (N_1150,N_732,N_1109);
and U1151 (N_1151,N_264,N_1102);
nand U1152 (N_1152,N_777,In_1765);
and U1153 (N_1153,In_364,In_653);
and U1154 (N_1154,N_1119,In_378);
xor U1155 (N_1155,N_849,In_1646);
nand U1156 (N_1156,In_423,N_775);
nor U1157 (N_1157,N_436,N_598);
and U1158 (N_1158,N_119,In_1630);
or U1159 (N_1159,N_1009,N_259);
xor U1160 (N_1160,N_1057,In_1851);
and U1161 (N_1161,N_821,N_1066);
nand U1162 (N_1162,In_291,N_920);
nor U1163 (N_1163,N_857,N_1050);
xnor U1164 (N_1164,N_815,In_1206);
nor U1165 (N_1165,In_1493,In_374);
and U1166 (N_1166,N_861,In_771);
xnor U1167 (N_1167,N_543,In_1149);
or U1168 (N_1168,N_867,In_1822);
xor U1169 (N_1169,N_1061,N_426);
xor U1170 (N_1170,In_222,N_668);
and U1171 (N_1171,In_1708,In_1403);
or U1172 (N_1172,N_694,In_1893);
or U1173 (N_1173,N_796,In_6);
and U1174 (N_1174,N_584,In_438);
or U1175 (N_1175,N_602,N_753);
nor U1176 (N_1176,In_1217,N_1104);
nand U1177 (N_1177,In_1629,N_1041);
nor U1178 (N_1178,In_1401,N_1097);
nand U1179 (N_1179,In_1614,N_977);
and U1180 (N_1180,N_929,N_881);
nand U1181 (N_1181,N_966,N_802);
or U1182 (N_1182,In_716,N_793);
and U1183 (N_1183,In_1028,In_546);
or U1184 (N_1184,N_1067,N_661);
nand U1185 (N_1185,N_1079,N_931);
or U1186 (N_1186,In_31,N_438);
nor U1187 (N_1187,N_1010,In_1748);
and U1188 (N_1188,In_999,N_501);
and U1189 (N_1189,N_84,N_642);
nand U1190 (N_1190,N_37,In_16);
xnor U1191 (N_1191,In_0,N_696);
xnor U1192 (N_1192,N_1077,In_738);
nor U1193 (N_1193,N_975,In_1174);
and U1194 (N_1194,N_719,N_1060);
or U1195 (N_1195,N_873,N_980);
and U1196 (N_1196,N_951,N_714);
nand U1197 (N_1197,N_539,N_798);
or U1198 (N_1198,N_634,In_184);
nor U1199 (N_1199,N_1032,N_1028);
xor U1200 (N_1200,N_779,N_811);
xnor U1201 (N_1201,In_1688,N_989);
xor U1202 (N_1202,N_1030,In_1816);
xor U1203 (N_1203,In_1628,In_842);
and U1204 (N_1204,In_679,N_446);
xor U1205 (N_1205,N_1042,N_116);
nor U1206 (N_1206,N_258,N_870);
and U1207 (N_1207,In_319,N_400);
xnor U1208 (N_1208,N_1062,N_746);
and U1209 (N_1209,In_1926,N_912);
and U1210 (N_1210,In_1699,In_1531);
or U1211 (N_1211,N_946,N_993);
and U1212 (N_1212,N_789,N_364);
xnor U1213 (N_1213,N_245,N_1011);
and U1214 (N_1214,In_179,N_6);
nor U1215 (N_1215,N_905,In_165);
nor U1216 (N_1216,N_976,In_809);
xnor U1217 (N_1217,N_960,N_1029);
nor U1218 (N_1218,In_233,N_969);
nor U1219 (N_1219,In_461,In_848);
and U1220 (N_1220,In_1038,N_817);
xor U1221 (N_1221,N_309,In_203);
and U1222 (N_1222,N_346,In_252);
xnor U1223 (N_1223,N_922,N_231);
or U1224 (N_1224,N_1074,N_506);
or U1225 (N_1225,N_713,In_948);
nor U1226 (N_1226,N_664,N_738);
nand U1227 (N_1227,N_674,In_1749);
or U1228 (N_1228,N_570,In_1190);
nor U1229 (N_1229,N_657,N_756);
nor U1230 (N_1230,N_711,In_429);
or U1231 (N_1231,N_646,In_1566);
nor U1232 (N_1232,N_212,In_1879);
or U1233 (N_1233,N_844,In_335);
xor U1234 (N_1234,N_1019,N_1046);
nand U1235 (N_1235,N_1089,In_59);
or U1236 (N_1236,N_872,In_881);
nor U1237 (N_1237,In_1458,N_996);
and U1238 (N_1238,N_1070,N_729);
or U1239 (N_1239,N_91,N_769);
and U1240 (N_1240,In_1097,In_1180);
nor U1241 (N_1241,In_1602,N_952);
or U1242 (N_1242,In_974,N_135);
nand U1243 (N_1243,N_882,N_626);
or U1244 (N_1244,In_109,In_1236);
and U1245 (N_1245,N_609,N_686);
nor U1246 (N_1246,In_1514,N_537);
or U1247 (N_1247,In_487,N_854);
or U1248 (N_1248,In_77,N_971);
or U1249 (N_1249,N_456,In_837);
xor U1250 (N_1250,In_1678,N_708);
and U1251 (N_1251,In_24,N_808);
nor U1252 (N_1252,N_653,N_1090);
or U1253 (N_1253,N_229,In_1144);
nand U1254 (N_1254,In_1923,N_903);
nor U1255 (N_1255,In_535,N_344);
nor U1256 (N_1256,N_1099,N_1063);
nand U1257 (N_1257,In_1500,N_925);
or U1258 (N_1258,N_900,N_1026);
xor U1259 (N_1259,N_577,N_628);
or U1260 (N_1260,N_1072,In_1359);
xor U1261 (N_1261,In_573,N_983);
and U1262 (N_1262,In_888,N_1052);
nor U1263 (N_1263,In_758,N_986);
or U1264 (N_1264,N_220,N_864);
and U1265 (N_1265,N_1088,In_1302);
nor U1266 (N_1266,In_511,N_262);
xnor U1267 (N_1267,In_1553,N_146);
or U1268 (N_1268,In_1842,N_755);
xor U1269 (N_1269,N_1035,N_712);
xor U1270 (N_1270,N_956,N_962);
xnor U1271 (N_1271,N_869,N_373);
nor U1272 (N_1272,N_704,N_892);
and U1273 (N_1273,N_376,In_54);
nand U1274 (N_1274,N_915,N_243);
nand U1275 (N_1275,N_914,In_105);
and U1276 (N_1276,In_1724,N_982);
and U1277 (N_1277,In_420,N_468);
nand U1278 (N_1278,In_882,N_812);
or U1279 (N_1279,N_274,N_998);
nand U1280 (N_1280,N_94,N_1161);
and U1281 (N_1281,N_1216,In_1806);
nand U1282 (N_1282,In_1585,N_1178);
nor U1283 (N_1283,In_1899,N_1253);
nand U1284 (N_1284,N_948,N_850);
or U1285 (N_1285,N_1278,In_1336);
nor U1286 (N_1286,N_886,N_1196);
nand U1287 (N_1287,N_935,N_1233);
xnor U1288 (N_1288,N_1256,N_999);
xnor U1289 (N_1289,N_1175,N_24);
nand U1290 (N_1290,In_1048,N_655);
or U1291 (N_1291,In_1162,N_1173);
or U1292 (N_1292,N_185,In_1716);
nand U1293 (N_1293,In_1567,N_1267);
xor U1294 (N_1294,In_1517,N_251);
nor U1295 (N_1295,In_409,In_1150);
or U1296 (N_1296,In_826,N_640);
nand U1297 (N_1297,N_542,N_1181);
xnor U1298 (N_1298,In_397,N_819);
or U1299 (N_1299,N_1273,In_1670);
nor U1300 (N_1300,In_1259,N_1230);
nand U1301 (N_1301,In_133,N_958);
xnor U1302 (N_1302,N_482,In_1616);
xnor U1303 (N_1303,N_1264,In_1291);
xor U1304 (N_1304,N_590,N_200);
xor U1305 (N_1305,N_603,In_230);
and U1306 (N_1306,N_1122,N_1192);
or U1307 (N_1307,In_1761,N_1127);
or U1308 (N_1308,N_1242,In_1598);
xnor U1309 (N_1309,N_324,In_183);
xor U1310 (N_1310,N_744,N_997);
xnor U1311 (N_1311,In_114,N_87);
and U1312 (N_1312,In_1355,In_1918);
nor U1313 (N_1313,N_1201,In_783);
nor U1314 (N_1314,N_1059,N_553);
xnor U1315 (N_1315,In_281,N_123);
and U1316 (N_1316,N_1228,N_1075);
or U1317 (N_1317,N_1110,In_86);
and U1318 (N_1318,N_1246,N_1259);
or U1319 (N_1319,N_1190,In_2);
or U1320 (N_1320,N_1241,N_1215);
and U1321 (N_1321,N_378,In_1220);
and U1322 (N_1322,N_488,In_495);
or U1323 (N_1323,In_1572,In_1972);
xnor U1324 (N_1324,In_44,N_1205);
or U1325 (N_1325,N_348,In_1040);
nor U1326 (N_1326,N_1095,N_574);
or U1327 (N_1327,N_967,In_1551);
or U1328 (N_1328,In_1837,N_405);
nand U1329 (N_1329,N_1100,N_1135);
and U1330 (N_1330,In_1509,N_978);
or U1331 (N_1331,In_1533,In_514);
xnor U1332 (N_1332,N_1255,In_845);
nand U1333 (N_1333,In_632,N_1166);
nor U1334 (N_1334,N_1087,N_1249);
nor U1335 (N_1335,N_833,In_225);
nand U1336 (N_1336,In_607,N_874);
and U1337 (N_1337,In_1882,In_1346);
nand U1338 (N_1338,N_985,In_1208);
nor U1339 (N_1339,N_1204,N_613);
nand U1340 (N_1340,N_644,N_856);
xnor U1341 (N_1341,N_1048,N_1214);
or U1342 (N_1342,N_1000,N_794);
nand U1343 (N_1343,N_1206,N_890);
nand U1344 (N_1344,In_1499,N_385);
xor U1345 (N_1345,N_1217,In_1951);
nand U1346 (N_1346,N_249,N_360);
xnor U1347 (N_1347,In_469,In_10);
nor U1348 (N_1348,N_484,N_1156);
or U1349 (N_1349,N_678,N_1128);
xnor U1350 (N_1350,N_125,N_328);
xnor U1351 (N_1351,In_524,N_1084);
nor U1352 (N_1352,N_1193,N_235);
nand U1353 (N_1353,In_907,N_407);
nand U1354 (N_1354,N_943,N_924);
and U1355 (N_1355,N_1034,N_1134);
nand U1356 (N_1356,N_687,In_1996);
nor U1357 (N_1357,N_1047,In_1042);
nand U1358 (N_1358,N_1265,N_825);
nor U1359 (N_1359,N_1210,In_654);
nor U1360 (N_1360,N_1172,N_937);
or U1361 (N_1361,N_564,N_1116);
and U1362 (N_1362,N_720,N_331);
or U1363 (N_1363,N_1163,N_1221);
xnor U1364 (N_1364,N_988,N_1017);
nand U1365 (N_1365,In_789,In_979);
and U1366 (N_1366,N_1154,N_884);
xor U1367 (N_1367,N_1006,N_1112);
xor U1368 (N_1368,N_1237,N_1198);
or U1369 (N_1369,In_520,In_453);
and U1370 (N_1370,In_1251,N_942);
xnor U1371 (N_1371,In_1133,N_121);
nand U1372 (N_1372,N_1014,N_938);
xnor U1373 (N_1373,N_1008,N_1148);
nor U1374 (N_1374,N_1195,N_1081);
nor U1375 (N_1375,N_1202,In_1);
and U1376 (N_1376,N_981,N_1044);
or U1377 (N_1377,N_964,N_743);
xnor U1378 (N_1378,In_1964,In_1192);
or U1379 (N_1379,N_1153,N_1269);
nor U1380 (N_1380,N_877,N_645);
nand U1381 (N_1381,N_1194,N_498);
xor U1382 (N_1382,N_409,N_1262);
or U1383 (N_1383,N_894,In_1601);
nor U1384 (N_1384,N_752,N_783);
xor U1385 (N_1385,N_820,N_1054);
nor U1386 (N_1386,In_768,N_1151);
nand U1387 (N_1387,N_288,N_941);
xnor U1388 (N_1388,N_880,N_1222);
or U1389 (N_1389,In_1218,In_853);
nand U1390 (N_1390,In_1737,N_1113);
nand U1391 (N_1391,N_1212,In_1649);
and U1392 (N_1392,N_1263,In_1990);
nor U1393 (N_1393,N_1203,N_1053);
xnor U1394 (N_1394,N_1016,In_1978);
or U1395 (N_1395,N_875,N_827);
and U1396 (N_1396,N_837,In_533);
nor U1397 (N_1397,N_1138,In_197);
and U1398 (N_1398,N_1147,N_911);
xor U1399 (N_1399,N_280,N_702);
and U1400 (N_1400,N_578,In_1703);
or U1401 (N_1401,N_926,N_464);
nand U1402 (N_1402,N_1125,In_1230);
nor U1403 (N_1403,In_1998,N_363);
and U1404 (N_1404,N_1123,N_1094);
xor U1405 (N_1405,N_485,N_67);
and U1406 (N_1406,In_1428,N_597);
nor U1407 (N_1407,N_615,In_750);
xor U1408 (N_1408,N_631,In_870);
nand U1409 (N_1409,N_510,N_760);
nor U1410 (N_1410,In_1932,N_432);
and U1411 (N_1411,N_1150,N_832);
xor U1412 (N_1412,In_1148,N_1137);
xnor U1413 (N_1413,In_704,N_1238);
nand U1414 (N_1414,In_1095,N_1183);
and U1415 (N_1415,N_1189,N_474);
nand U1416 (N_1416,N_1003,N_1049);
or U1417 (N_1417,N_961,In_467);
nand U1418 (N_1418,N_1142,In_286);
nand U1419 (N_1419,N_301,N_845);
or U1420 (N_1420,N_1093,In_1073);
nand U1421 (N_1421,N_1223,In_793);
nand U1422 (N_1422,N_791,In_746);
nand U1423 (N_1423,In_75,N_1140);
nor U1424 (N_1424,In_1516,N_1023);
or U1425 (N_1425,N_544,N_955);
and U1426 (N_1426,N_418,N_1157);
xor U1427 (N_1427,N_1243,N_1180);
xnor U1428 (N_1428,N_1033,N_904);
nand U1429 (N_1429,N_896,N_415);
nand U1430 (N_1430,N_1164,N_994);
nor U1431 (N_1431,N_1001,In_338);
nand U1432 (N_1432,N_1174,N_1005);
nor U1433 (N_1433,N_1274,In_1881);
xor U1434 (N_1434,N_1058,N_1143);
or U1435 (N_1435,In_1606,N_1219);
xnor U1436 (N_1436,N_271,N_828);
or U1437 (N_1437,N_142,N_1101);
xor U1438 (N_1438,N_73,In_398);
nand U1439 (N_1439,In_1024,N_169);
nor U1440 (N_1440,N_1418,N_1159);
nor U1441 (N_1441,N_1275,N_940);
xor U1442 (N_1442,N_550,N_1076);
nor U1443 (N_1443,N_1260,In_1448);
nor U1444 (N_1444,N_1389,N_1425);
nor U1445 (N_1445,N_1428,N_703);
xnor U1446 (N_1446,N_739,N_1085);
nand U1447 (N_1447,In_1254,N_1131);
nor U1448 (N_1448,N_1211,N_1276);
nand U1449 (N_1449,In_18,N_1287);
nor U1450 (N_1450,N_768,In_1043);
xnor U1451 (N_1451,In_547,In_1878);
or U1452 (N_1452,N_1268,N_592);
nand U1453 (N_1453,In_449,N_535);
or U1454 (N_1454,N_848,N_1350);
or U1455 (N_1455,N_965,N_1218);
or U1456 (N_1456,In_657,N_936);
and U1457 (N_1457,In_427,N_1318);
or U1458 (N_1458,N_1412,N_1315);
xor U1459 (N_1459,N_662,N_1432);
xor U1460 (N_1460,In_1101,N_362);
and U1461 (N_1461,N_973,In_1394);
or U1462 (N_1462,N_1342,In_1592);
nand U1463 (N_1463,In_1694,N_1271);
or U1464 (N_1464,N_1340,N_1279);
and U1465 (N_1465,N_706,N_979);
xnor U1466 (N_1466,In_969,N_1435);
nand U1467 (N_1467,N_715,N_991);
nor U1468 (N_1468,N_1132,In_1679);
nand U1469 (N_1469,N_1083,N_1229);
nand U1470 (N_1470,N_1325,N_1024);
nor U1471 (N_1471,N_1313,N_1378);
and U1472 (N_1472,In_1697,N_573);
and U1473 (N_1473,N_296,N_1298);
xnor U1474 (N_1474,In_1605,In_1440);
xnor U1475 (N_1475,In_115,In_748);
xnor U1476 (N_1476,N_472,N_1169);
nand U1477 (N_1477,In_1056,N_1261);
nand U1478 (N_1478,N_974,N_1064);
or U1479 (N_1479,In_1035,N_1111);
nor U1480 (N_1480,N_725,N_437);
and U1481 (N_1481,N_1293,In_1014);
nand U1482 (N_1482,N_1405,N_1018);
and U1483 (N_1483,N_1092,In_339);
or U1484 (N_1484,N_1329,N_1406);
xnor U1485 (N_1485,In_1683,N_1117);
nand U1486 (N_1486,In_1396,N_990);
nor U1487 (N_1487,N_908,N_1007);
and U1488 (N_1488,N_1020,N_1022);
or U1489 (N_1489,N_357,In_1715);
xnor U1490 (N_1490,In_454,N_1068);
nand U1491 (N_1491,N_675,N_383);
xnor U1492 (N_1492,In_1537,N_1334);
and U1493 (N_1493,N_1141,In_195);
nand U1494 (N_1494,N_586,In_1475);
or U1495 (N_1495,N_1272,N_918);
and U1496 (N_1496,N_317,N_491);
nand U1497 (N_1497,N_1144,N_1319);
and U1498 (N_1498,N_1040,In_34);
or U1499 (N_1499,N_1086,N_1376);
xnor U1500 (N_1500,In_641,N_1277);
nand U1501 (N_1501,N_1096,N_893);
xor U1502 (N_1502,N_1179,N_1012);
and U1503 (N_1503,In_1684,N_522);
nand U1504 (N_1504,N_972,N_366);
and U1505 (N_1505,In_1381,N_458);
or U1506 (N_1506,In_1385,In_1112);
nor U1507 (N_1507,In_1784,N_122);
and U1508 (N_1508,N_1200,N_1254);
or U1509 (N_1509,N_876,In_270);
nor U1510 (N_1510,N_1158,N_1227);
xor U1511 (N_1511,In_315,N_1426);
or U1512 (N_1512,N_1300,N_1231);
or U1513 (N_1513,N_1208,N_538);
nor U1514 (N_1514,N_396,In_1465);
nand U1515 (N_1515,N_1236,N_1281);
nand U1516 (N_1516,N_1307,N_178);
xnor U1517 (N_1517,N_1355,N_1346);
nor U1518 (N_1518,N_1234,N_412);
xor U1519 (N_1519,In_407,In_1305);
nand U1520 (N_1520,N_1292,N_717);
or U1521 (N_1521,N_582,In_1853);
xnor U1522 (N_1522,N_1359,N_1283);
xnor U1523 (N_1523,In_591,N_1091);
or U1524 (N_1524,N_1295,N_1299);
or U1525 (N_1525,N_525,N_1069);
or U1526 (N_1526,N_987,N_1182);
and U1527 (N_1527,N_927,N_1078);
or U1528 (N_1528,N_663,In_367);
or U1529 (N_1529,N_847,N_1073);
or U1530 (N_1530,N_1411,N_1187);
nor U1531 (N_1531,In_48,N_1344);
nand U1532 (N_1532,N_1184,N_1289);
and U1533 (N_1533,N_1384,N_1129);
xnor U1534 (N_1534,N_1341,N_806);
and U1535 (N_1535,N_1266,N_524);
and U1536 (N_1536,N_1130,N_1419);
xnor U1537 (N_1537,N_1036,In_1987);
or U1538 (N_1538,In_177,N_1424);
nor U1539 (N_1539,N_1413,N_1331);
xnor U1540 (N_1540,N_866,N_1391);
or U1541 (N_1541,N_1280,N_1160);
nand U1542 (N_1542,N_1170,N_1240);
nand U1543 (N_1543,N_1270,In_897);
nor U1544 (N_1544,N_163,N_1377);
xnor U1545 (N_1545,N_1152,N_1400);
xnor U1546 (N_1546,N_1149,N_1408);
nor U1547 (N_1547,In_314,N_838);
and U1548 (N_1548,In_1433,In_1076);
nor U1549 (N_1549,In_201,N_1145);
nand U1550 (N_1550,N_1056,N_1423);
nor U1551 (N_1551,N_1321,N_1357);
xor U1552 (N_1552,N_1177,N_1328);
or U1553 (N_1553,N_1039,N_594);
and U1554 (N_1554,N_1403,N_1188);
and U1555 (N_1555,N_1250,N_1422);
xor U1556 (N_1556,N_741,N_1167);
or U1557 (N_1557,N_1248,N_860);
xnor U1558 (N_1558,In_900,N_1199);
and U1559 (N_1559,N_1133,In_1577);
xnor U1560 (N_1560,N_1343,In_1549);
and U1561 (N_1561,In_383,In_1960);
nand U1562 (N_1562,N_1322,N_1368);
nand U1563 (N_1563,N_532,N_1291);
xor U1564 (N_1564,N_800,N_995);
xnor U1565 (N_1565,In_88,N_1439);
or U1566 (N_1566,N_865,In_234);
nand U1567 (N_1567,In_1326,N_705);
or U1568 (N_1568,N_1312,N_606);
or U1569 (N_1569,In_798,N_1107);
and U1570 (N_1570,N_1375,In_1419);
or U1571 (N_1571,N_1335,N_1186);
and U1572 (N_1572,N_1191,N_1317);
or U1573 (N_1573,N_1392,In_134);
nand U1574 (N_1574,N_879,N_858);
nor U1575 (N_1575,N_370,N_826);
and U1576 (N_1576,N_680,N_1365);
or U1577 (N_1577,In_1596,N_1124);
nor U1578 (N_1578,N_1374,N_963);
nor U1579 (N_1579,N_1176,N_1120);
nand U1580 (N_1580,N_1332,N_1324);
xnor U1581 (N_1581,N_451,N_1168);
or U1582 (N_1582,In_1525,In_127);
or U1583 (N_1583,N_114,N_787);
xor U1584 (N_1584,N_1430,N_1361);
or U1585 (N_1585,N_473,In_920);
and U1586 (N_1586,In_1644,N_377);
or U1587 (N_1587,In_1376,N_1162);
nor U1588 (N_1588,In_96,N_1380);
and U1589 (N_1589,In_1767,N_1420);
nor U1590 (N_1590,N_1296,N_1326);
and U1591 (N_1591,N_1416,In_128);
nor U1592 (N_1592,In_187,In_147);
or U1593 (N_1593,N_189,In_1351);
or U1594 (N_1594,N_1013,N_1397);
xor U1595 (N_1595,In_1016,N_1302);
nand U1596 (N_1596,N_1239,N_1165);
nand U1597 (N_1597,N_788,N_868);
nor U1598 (N_1598,N_1294,N_440);
nor U1599 (N_1599,N_1257,N_292);
nand U1600 (N_1600,In_309,N_1410);
and U1601 (N_1601,N_1503,N_1471);
and U1602 (N_1602,In_325,N_1407);
nand U1603 (N_1603,In_1859,N_773);
and U1604 (N_1604,N_152,N_1209);
nand U1605 (N_1605,N_1414,N_1543);
nor U1606 (N_1606,N_1399,N_1055);
or U1607 (N_1607,N_1493,N_841);
and U1608 (N_1608,N_1515,N_1285);
nor U1609 (N_1609,N_1235,N_1510);
or U1610 (N_1610,N_1462,N_1108);
and U1611 (N_1611,N_1583,N_1347);
and U1612 (N_1612,In_1917,N_1449);
nor U1613 (N_1613,N_1105,In_1423);
nand U1614 (N_1614,N_1244,N_1385);
nor U1615 (N_1615,N_795,N_1504);
and U1616 (N_1616,N_1469,N_1593);
xnor U1617 (N_1617,N_1536,N_1478);
xnor U1618 (N_1618,N_1559,N_1458);
or U1619 (N_1619,N_1245,N_1457);
nand U1620 (N_1620,N_888,N_1598);
or U1621 (N_1621,N_1562,In_23);
xnor U1622 (N_1622,N_1103,In_1810);
xor U1623 (N_1623,In_1059,N_1305);
nor U1624 (N_1624,N_1303,N_1031);
or U1625 (N_1625,N_1538,In_597);
or U1626 (N_1626,N_1574,N_1596);
xor U1627 (N_1627,In_1921,N_1320);
nor U1628 (N_1628,N_1436,N_1118);
nor U1629 (N_1629,N_1529,N_1492);
nor U1630 (N_1630,N_944,N_1480);
xnor U1631 (N_1631,N_1589,N_1502);
nand U1632 (N_1632,N_1314,N_1025);
xnor U1633 (N_1633,N_1597,N_1065);
or U1634 (N_1634,N_1348,N_1585);
nand U1635 (N_1635,N_1468,In_517);
nand U1636 (N_1636,N_1496,N_1364);
nor U1637 (N_1637,In_1211,N_575);
and U1638 (N_1638,In_436,In_1189);
or U1639 (N_1639,In_1445,N_724);
or U1640 (N_1640,N_1485,N_1323);
xnor U1641 (N_1641,N_1136,N_1551);
xor U1642 (N_1642,N_1444,N_1587);
or U1643 (N_1643,N_100,N_1573);
and U1644 (N_1644,N_1434,N_512);
and U1645 (N_1645,N_1015,N_1508);
nor U1646 (N_1646,N_1467,In_1507);
or U1647 (N_1647,N_1518,N_384);
nor U1648 (N_1648,N_536,N_1316);
and U1649 (N_1649,N_1546,N_1288);
or U1650 (N_1650,N_1534,In_1130);
or U1651 (N_1651,N_1568,In_37);
nand U1652 (N_1652,N_320,N_1530);
xnor U1653 (N_1653,N_1345,In_970);
and U1654 (N_1654,In_1488,N_1522);
nand U1655 (N_1655,In_624,N_548);
nor U1656 (N_1656,N_1207,N_707);
and U1657 (N_1657,N_692,N_1388);
or U1658 (N_1658,N_1539,N_1080);
and U1659 (N_1659,N_1532,N_1396);
nand U1660 (N_1660,N_1045,N_1472);
or U1661 (N_1661,N_1284,N_1509);
nor U1662 (N_1662,N_1487,N_1398);
nand U1663 (N_1663,N_1486,N_454);
xor U1664 (N_1664,In_1313,N_1309);
nand U1665 (N_1665,N_1442,In_1766);
and U1666 (N_1666,In_961,N_757);
nor U1667 (N_1667,N_1448,N_1465);
and U1668 (N_1668,N_1500,N_1582);
nor U1669 (N_1669,In_906,N_891);
or U1670 (N_1670,N_1566,N_1521);
xnor U1671 (N_1671,N_1463,In_1639);
nand U1672 (N_1672,N_1258,N_1579);
and U1673 (N_1673,N_1584,N_1333);
or U1674 (N_1674,N_1501,N_1360);
and U1675 (N_1675,In_1082,N_778);
nor U1676 (N_1676,N_1577,N_1356);
nand U1677 (N_1677,N_1431,N_1476);
nand U1678 (N_1678,In_417,N_1451);
and U1679 (N_1679,In_620,N_1578);
nand U1680 (N_1680,N_984,In_943);
nand U1681 (N_1681,In_1318,In_1034);
nand U1682 (N_1682,In_1344,N_1595);
nand U1683 (N_1683,N_846,N_1126);
or U1684 (N_1684,N_1464,N_1560);
nor U1685 (N_1685,N_1443,N_1479);
and U1686 (N_1686,N_1488,N_1367);
xor U1687 (N_1687,N_1549,N_1417);
nand U1688 (N_1688,N_1513,N_1561);
nand U1689 (N_1689,N_1404,N_878);
or U1690 (N_1690,N_1226,N_1415);
nand U1691 (N_1691,N_1382,N_1494);
or U1692 (N_1692,N_1524,N_1514);
nand U1693 (N_1693,N_1220,N_1499);
nor U1694 (N_1694,In_1239,N_619);
and U1695 (N_1695,N_1051,N_1552);
xnor U1696 (N_1696,N_1592,N_1474);
or U1697 (N_1697,N_1252,N_589);
or U1698 (N_1698,N_1475,N_1580);
xnor U1699 (N_1699,N_1516,N_1507);
and U1700 (N_1700,N_992,N_889);
or U1701 (N_1701,In_1892,N_1466);
nor U1702 (N_1702,N_1527,N_1540);
xnor U1703 (N_1703,N_1330,N_1542);
nor U1704 (N_1704,N_279,N_1383);
nor U1705 (N_1705,In_441,N_1576);
or U1706 (N_1706,In_1632,N_1453);
xnor U1707 (N_1707,N_1563,N_1146);
xor U1708 (N_1708,N_1541,N_1071);
or U1709 (N_1709,N_1454,In_359);
nand U1710 (N_1710,N_1452,N_1590);
nand U1711 (N_1711,N_690,N_1371);
xor U1712 (N_1712,N_1353,N_297);
and U1713 (N_1713,N_1531,N_1481);
and U1714 (N_1714,N_1461,In_207);
nand U1715 (N_1715,N_108,N_1447);
nor U1716 (N_1716,N_1441,N_1525);
xor U1717 (N_1717,N_1520,N_1548);
nor U1718 (N_1718,N_1395,N_1114);
or U1719 (N_1719,N_1528,N_1297);
and U1720 (N_1720,N_1402,N_1438);
nor U1721 (N_1721,N_234,N_1387);
and U1722 (N_1722,N_1571,N_263);
xnor U1723 (N_1723,N_1470,N_1311);
or U1724 (N_1724,N_859,N_1506);
nor U1725 (N_1725,N_1517,N_1572);
and U1726 (N_1726,In_1004,N_1588);
or U1727 (N_1727,N_1004,N_1575);
nor U1728 (N_1728,N_1393,N_1247);
xor U1729 (N_1729,N_1338,N_1185);
nor U1730 (N_1730,N_392,N_1594);
or U1731 (N_1731,N_1490,N_1554);
xnor U1732 (N_1732,N_1491,N_1553);
or U1733 (N_1733,N_1484,N_1301);
or U1734 (N_1734,N_1369,N_1370);
xor U1735 (N_1735,N_1363,N_1390);
or U1736 (N_1736,N_1308,In_765);
nand U1737 (N_1737,N_1290,N_1366);
nand U1738 (N_1738,N_1460,N_1526);
or U1739 (N_1739,N_1450,N_1495);
nor U1740 (N_1740,In_1204,N_1306);
nor U1741 (N_1741,In_1804,N_1351);
nand U1742 (N_1742,N_1545,In_1316);
and U1743 (N_1743,N_1570,N_1421);
nand U1744 (N_1744,N_1567,In_1478);
nor U1745 (N_1745,In_977,N_1591);
and U1746 (N_1746,N_1394,N_16);
nand U1747 (N_1747,N_1171,N_1599);
or U1748 (N_1748,In_1005,N_1533);
xnor U1749 (N_1749,N_1337,N_1373);
xnor U1750 (N_1750,N_652,N_970);
or U1751 (N_1751,N_1445,In_1686);
xnor U1752 (N_1752,N_917,N_1121);
and U1753 (N_1753,N_1456,N_1225);
xnor U1754 (N_1754,N_1310,N_1550);
and U1755 (N_1755,N_1213,N_1556);
nand U1756 (N_1756,In_1846,N_1155);
nor U1757 (N_1757,N_1512,N_238);
xor U1758 (N_1758,N_1569,In_1675);
nand U1759 (N_1759,N_471,N_1523);
nand U1760 (N_1760,N_1557,N_1690);
xor U1761 (N_1761,N_1692,In_432);
xnor U1762 (N_1762,N_1139,N_1535);
nand U1763 (N_1763,N_1698,N_1723);
nand U1764 (N_1764,N_1718,N_1696);
and U1765 (N_1765,N_1282,N_1744);
or U1766 (N_1766,N_1645,N_1709);
or U1767 (N_1767,N_1615,N_1739);
xor U1768 (N_1768,N_1706,In_1473);
or U1769 (N_1769,N_1684,N_1612);
or U1770 (N_1770,N_1682,N_1633);
or U1771 (N_1771,N_1647,In_1417);
nor U1772 (N_1772,N_1734,N_1624);
nor U1773 (N_1773,N_1687,N_1637);
or U1774 (N_1774,N_629,N_1742);
nor U1775 (N_1775,N_1547,N_1565);
xor U1776 (N_1776,N_1610,N_1544);
and U1777 (N_1777,N_78,N_1603);
nor U1778 (N_1778,N_1477,In_1400);
or U1779 (N_1779,N_1605,N_1654);
xor U1780 (N_1780,N_1623,N_1620);
and U1781 (N_1781,N_1649,N_1746);
and U1782 (N_1782,N_1586,N_1663);
and U1783 (N_1783,N_1661,N_1497);
and U1784 (N_1784,N_1611,N_1648);
or U1785 (N_1785,N_1681,N_1651);
nor U1786 (N_1786,N_1286,N_1655);
nand U1787 (N_1787,N_1604,In_1857);
xor U1788 (N_1788,N_1702,N_1667);
and U1789 (N_1789,N_1745,N_1197);
nand U1790 (N_1790,N_1724,N_1354);
xor U1791 (N_1791,N_1673,N_1688);
nor U1792 (N_1792,N_1427,N_1082);
xor U1793 (N_1793,N_1429,N_1735);
and U1794 (N_1794,N_1641,N_1339);
or U1795 (N_1795,N_1511,N_1379);
and U1796 (N_1796,In_703,N_1741);
nand U1797 (N_1797,N_1607,N_66);
nand U1798 (N_1798,N_1634,N_1737);
xnor U1799 (N_1799,N_1644,In_188);
xnor U1800 (N_1800,N_1657,N_1440);
xnor U1801 (N_1801,N_1483,N_1733);
xor U1802 (N_1802,N_1618,N_1098);
nor U1803 (N_1803,N_1608,N_1665);
nand U1804 (N_1804,N_1712,N_1685);
and U1805 (N_1805,N_1704,N_1727);
nand U1806 (N_1806,N_1616,N_1757);
nor U1807 (N_1807,N_1631,N_1756);
or U1808 (N_1808,N_1433,N_1437);
nor U1809 (N_1809,N_1662,N_427);
or U1810 (N_1810,N_1636,N_1658);
or U1811 (N_1811,N_1666,N_1689);
or U1812 (N_1812,N_1482,N_1699);
and U1813 (N_1813,N_913,N_1711);
nand U1814 (N_1814,N_1659,In_1534);
or U1815 (N_1815,N_1738,N_1732);
nand U1816 (N_1816,N_1715,N_1498);
or U1817 (N_1817,N_939,N_1358);
or U1818 (N_1818,N_1725,N_1679);
or U1819 (N_1819,N_1002,N_1705);
nor U1820 (N_1820,N_1601,N_1650);
nor U1821 (N_1821,N_1747,N_1386);
and U1822 (N_1822,N_1251,N_1653);
or U1823 (N_1823,N_1752,N_1621);
nand U1824 (N_1824,N_1694,N_1642);
nand U1825 (N_1825,N_1668,In_410);
nor U1826 (N_1826,N_1677,N_1686);
nor U1827 (N_1827,N_96,N_1232);
xor U1828 (N_1828,N_1755,N_547);
xor U1829 (N_1829,N_1409,N_1697);
nor U1830 (N_1830,In_822,N_1675);
nor U1831 (N_1831,N_1672,N_1327);
or U1832 (N_1832,N_1646,N_1717);
or U1833 (N_1833,N_1707,N_1714);
nand U1834 (N_1834,N_1304,N_1736);
and U1835 (N_1835,N_1638,N_1750);
and U1836 (N_1836,N_1703,N_1669);
and U1837 (N_1837,N_1652,N_1740);
and U1838 (N_1838,N_1630,In_861);
nand U1839 (N_1839,N_1680,N_1695);
nand U1840 (N_1840,N_1505,N_1674);
and U1841 (N_1841,N_1729,N_1664);
nor U1842 (N_1842,N_1721,N_1489);
nor U1843 (N_1843,N_1629,N_1748);
or U1844 (N_1844,N_1352,N_1027);
nor U1845 (N_1845,In_791,N_1639);
nor U1846 (N_1846,N_1693,N_1606);
and U1847 (N_1847,N_404,N_1635);
nor U1848 (N_1848,N_1722,N_1632);
nor U1849 (N_1849,N_1678,N_1759);
or U1850 (N_1850,N_1720,N_1640);
nand U1851 (N_1851,N_840,N_1643);
xor U1852 (N_1852,N_1558,N_356);
xor U1853 (N_1853,N_1459,N_1670);
xor U1854 (N_1854,N_1602,N_1625);
or U1855 (N_1855,N_1701,N_1555);
and U1856 (N_1856,N_1613,N_1626);
and U1857 (N_1857,N_1381,N_1676);
nand U1858 (N_1858,N_1362,N_1401);
or U1859 (N_1859,N_1349,N_1719);
and U1860 (N_1860,N_1473,N_1716);
nor U1861 (N_1861,N_1728,N_1726);
and U1862 (N_1862,N_1743,N_1600);
or U1863 (N_1863,N_1614,N_1730);
nor U1864 (N_1864,N_1581,N_1691);
nor U1865 (N_1865,N_1617,N_1627);
and U1866 (N_1866,In_1441,N_1455);
and U1867 (N_1867,N_1619,N_1564);
nor U1868 (N_1868,N_1754,N_1519);
nand U1869 (N_1869,N_1671,N_1751);
xnor U1870 (N_1870,N_1708,N_1749);
or U1871 (N_1871,N_1700,N_1372);
xnor U1872 (N_1872,N_1713,N_1224);
and U1873 (N_1873,N_1622,N_1628);
or U1874 (N_1874,N_1758,In_450);
xnor U1875 (N_1875,N_1446,N_1656);
and U1876 (N_1876,N_1731,N_1537);
and U1877 (N_1877,N_1609,N_1660);
nor U1878 (N_1878,N_1753,N_1683);
nor U1879 (N_1879,N_1710,N_1336);
nand U1880 (N_1880,N_1650,N_1662);
nand U1881 (N_1881,N_1327,N_1630);
or U1882 (N_1882,N_1623,N_356);
nand U1883 (N_1883,N_1666,N_1304);
nand U1884 (N_1884,N_1354,N_840);
and U1885 (N_1885,N_1705,N_1427);
and U1886 (N_1886,N_1489,N_1654);
xnor U1887 (N_1887,N_1002,N_1618);
and U1888 (N_1888,N_1735,In_1400);
and U1889 (N_1889,N_1708,N_1082);
and U1890 (N_1890,N_1677,N_1700);
nand U1891 (N_1891,N_1713,N_1625);
or U1892 (N_1892,N_1642,N_1730);
nand U1893 (N_1893,N_1723,N_1741);
and U1894 (N_1894,N_1618,N_1644);
and U1895 (N_1895,N_1680,N_1718);
or U1896 (N_1896,N_1700,N_1743);
nor U1897 (N_1897,N_1662,N_1711);
nor U1898 (N_1898,N_1354,N_1657);
and U1899 (N_1899,N_1756,N_1732);
nor U1900 (N_1900,N_1752,N_1756);
xnor U1901 (N_1901,N_1645,N_1477);
or U1902 (N_1902,N_1693,N_1651);
nor U1903 (N_1903,N_1352,N_1740);
nand U1904 (N_1904,In_703,N_1637);
nand U1905 (N_1905,N_1680,N_1708);
nor U1906 (N_1906,N_1616,N_1649);
nand U1907 (N_1907,N_1681,N_1666);
nand U1908 (N_1908,N_1654,N_1098);
or U1909 (N_1909,N_1619,N_1688);
or U1910 (N_1910,N_1637,N_1027);
xor U1911 (N_1911,N_1586,N_1637);
and U1912 (N_1912,N_1707,N_1731);
nand U1913 (N_1913,N_1558,N_1658);
xor U1914 (N_1914,N_1717,N_1625);
xor U1915 (N_1915,N_1564,N_1642);
or U1916 (N_1916,N_1747,N_1696);
or U1917 (N_1917,In_1857,N_1674);
and U1918 (N_1918,N_1690,N_1647);
or U1919 (N_1919,N_1282,N_1251);
and U1920 (N_1920,N_1895,N_1803);
xor U1921 (N_1921,N_1871,N_1894);
or U1922 (N_1922,N_1771,N_1804);
nor U1923 (N_1923,N_1792,N_1886);
nand U1924 (N_1924,N_1866,N_1763);
and U1925 (N_1925,N_1761,N_1773);
or U1926 (N_1926,N_1917,N_1764);
and U1927 (N_1927,N_1860,N_1853);
xnor U1928 (N_1928,N_1760,N_1859);
nand U1929 (N_1929,N_1880,N_1887);
or U1930 (N_1930,N_1870,N_1893);
xor U1931 (N_1931,N_1903,N_1913);
xor U1932 (N_1932,N_1851,N_1772);
and U1933 (N_1933,N_1912,N_1826);
nor U1934 (N_1934,N_1831,N_1809);
or U1935 (N_1935,N_1915,N_1876);
nor U1936 (N_1936,N_1820,N_1815);
nor U1937 (N_1937,N_1786,N_1787);
nor U1938 (N_1938,N_1850,N_1885);
or U1939 (N_1939,N_1813,N_1841);
xor U1940 (N_1940,N_1856,N_1867);
xor U1941 (N_1941,N_1800,N_1794);
or U1942 (N_1942,N_1878,N_1762);
nor U1943 (N_1943,N_1846,N_1821);
or U1944 (N_1944,N_1905,N_1770);
xor U1945 (N_1945,N_1840,N_1843);
xor U1946 (N_1946,N_1896,N_1776);
and U1947 (N_1947,N_1814,N_1795);
nor U1948 (N_1948,N_1911,N_1863);
nor U1949 (N_1949,N_1779,N_1910);
and U1950 (N_1950,N_1799,N_1854);
and U1951 (N_1951,N_1852,N_1844);
xor U1952 (N_1952,N_1819,N_1857);
nor U1953 (N_1953,N_1883,N_1879);
nor U1954 (N_1954,N_1832,N_1918);
xnor U1955 (N_1955,N_1801,N_1909);
nor U1956 (N_1956,N_1884,N_1765);
and U1957 (N_1957,N_1899,N_1817);
or U1958 (N_1958,N_1872,N_1790);
and U1959 (N_1959,N_1825,N_1797);
or U1960 (N_1960,N_1902,N_1783);
nand U1961 (N_1961,N_1780,N_1836);
nor U1962 (N_1962,N_1833,N_1782);
and U1963 (N_1963,N_1789,N_1906);
or U1964 (N_1964,N_1769,N_1796);
and U1965 (N_1965,N_1808,N_1904);
nor U1966 (N_1966,N_1868,N_1805);
nand U1967 (N_1967,N_1914,N_1891);
xnor U1968 (N_1968,N_1807,N_1873);
nor U1969 (N_1969,N_1916,N_1861);
nand U1970 (N_1970,N_1818,N_1784);
and U1971 (N_1971,N_1806,N_1816);
nand U1972 (N_1972,N_1785,N_1855);
and U1973 (N_1973,N_1830,N_1791);
nor U1974 (N_1974,N_1824,N_1842);
xor U1975 (N_1975,N_1838,N_1862);
xor U1976 (N_1976,N_1828,N_1798);
xnor U1977 (N_1977,N_1901,N_1775);
xor U1978 (N_1978,N_1834,N_1835);
xnor U1979 (N_1979,N_1858,N_1907);
nor U1980 (N_1980,N_1888,N_1869);
or U1981 (N_1981,N_1889,N_1877);
xor U1982 (N_1982,N_1919,N_1766);
and U1983 (N_1983,N_1897,N_1829);
nand U1984 (N_1984,N_1812,N_1900);
and U1985 (N_1985,N_1822,N_1767);
nand U1986 (N_1986,N_1890,N_1793);
nand U1987 (N_1987,N_1802,N_1865);
or U1988 (N_1988,N_1874,N_1768);
nor U1989 (N_1989,N_1823,N_1810);
nand U1990 (N_1990,N_1908,N_1875);
nor U1991 (N_1991,N_1892,N_1827);
or U1992 (N_1992,N_1788,N_1811);
and U1993 (N_1993,N_1882,N_1848);
and U1994 (N_1994,N_1777,N_1864);
nor U1995 (N_1995,N_1837,N_1845);
nand U1996 (N_1996,N_1778,N_1774);
nand U1997 (N_1997,N_1839,N_1781);
or U1998 (N_1998,N_1881,N_1849);
and U1999 (N_1999,N_1898,N_1847);
or U2000 (N_2000,N_1800,N_1868);
xor U2001 (N_2001,N_1848,N_1764);
and U2002 (N_2002,N_1807,N_1825);
xor U2003 (N_2003,N_1859,N_1883);
xor U2004 (N_2004,N_1910,N_1879);
xnor U2005 (N_2005,N_1802,N_1898);
nor U2006 (N_2006,N_1771,N_1912);
xor U2007 (N_2007,N_1918,N_1883);
xor U2008 (N_2008,N_1917,N_1875);
and U2009 (N_2009,N_1906,N_1794);
nor U2010 (N_2010,N_1898,N_1911);
nor U2011 (N_2011,N_1809,N_1878);
nand U2012 (N_2012,N_1864,N_1819);
nand U2013 (N_2013,N_1830,N_1815);
nor U2014 (N_2014,N_1868,N_1891);
nand U2015 (N_2015,N_1902,N_1798);
nor U2016 (N_2016,N_1897,N_1775);
nor U2017 (N_2017,N_1815,N_1785);
nand U2018 (N_2018,N_1769,N_1912);
nand U2019 (N_2019,N_1816,N_1780);
and U2020 (N_2020,N_1847,N_1884);
or U2021 (N_2021,N_1896,N_1822);
and U2022 (N_2022,N_1810,N_1831);
nor U2023 (N_2023,N_1891,N_1895);
nand U2024 (N_2024,N_1838,N_1857);
or U2025 (N_2025,N_1800,N_1809);
nor U2026 (N_2026,N_1890,N_1888);
nand U2027 (N_2027,N_1805,N_1875);
and U2028 (N_2028,N_1857,N_1911);
or U2029 (N_2029,N_1866,N_1889);
or U2030 (N_2030,N_1764,N_1775);
or U2031 (N_2031,N_1817,N_1915);
nand U2032 (N_2032,N_1772,N_1872);
nor U2033 (N_2033,N_1868,N_1841);
nand U2034 (N_2034,N_1879,N_1876);
and U2035 (N_2035,N_1776,N_1835);
xor U2036 (N_2036,N_1902,N_1866);
nor U2037 (N_2037,N_1779,N_1909);
and U2038 (N_2038,N_1904,N_1803);
or U2039 (N_2039,N_1760,N_1808);
xnor U2040 (N_2040,N_1825,N_1873);
and U2041 (N_2041,N_1899,N_1847);
nand U2042 (N_2042,N_1780,N_1831);
or U2043 (N_2043,N_1792,N_1770);
xor U2044 (N_2044,N_1812,N_1766);
and U2045 (N_2045,N_1805,N_1870);
nor U2046 (N_2046,N_1843,N_1794);
or U2047 (N_2047,N_1792,N_1841);
nand U2048 (N_2048,N_1818,N_1908);
and U2049 (N_2049,N_1831,N_1908);
nand U2050 (N_2050,N_1849,N_1790);
or U2051 (N_2051,N_1885,N_1847);
nand U2052 (N_2052,N_1839,N_1842);
and U2053 (N_2053,N_1909,N_1894);
xnor U2054 (N_2054,N_1769,N_1905);
or U2055 (N_2055,N_1863,N_1876);
xor U2056 (N_2056,N_1774,N_1801);
or U2057 (N_2057,N_1844,N_1808);
nor U2058 (N_2058,N_1840,N_1821);
xor U2059 (N_2059,N_1910,N_1891);
or U2060 (N_2060,N_1821,N_1837);
nor U2061 (N_2061,N_1854,N_1791);
nand U2062 (N_2062,N_1818,N_1918);
and U2063 (N_2063,N_1820,N_1773);
nand U2064 (N_2064,N_1890,N_1858);
and U2065 (N_2065,N_1883,N_1836);
xor U2066 (N_2066,N_1882,N_1896);
xnor U2067 (N_2067,N_1903,N_1854);
nor U2068 (N_2068,N_1831,N_1915);
nand U2069 (N_2069,N_1855,N_1823);
nand U2070 (N_2070,N_1792,N_1879);
or U2071 (N_2071,N_1769,N_1833);
and U2072 (N_2072,N_1782,N_1769);
and U2073 (N_2073,N_1889,N_1835);
nor U2074 (N_2074,N_1784,N_1879);
nor U2075 (N_2075,N_1883,N_1890);
nand U2076 (N_2076,N_1873,N_1762);
and U2077 (N_2077,N_1913,N_1839);
xnor U2078 (N_2078,N_1842,N_1872);
or U2079 (N_2079,N_1817,N_1785);
xor U2080 (N_2080,N_1948,N_2010);
and U2081 (N_2081,N_1921,N_2066);
xnor U2082 (N_2082,N_1951,N_2007);
xnor U2083 (N_2083,N_1980,N_1992);
xnor U2084 (N_2084,N_2055,N_1976);
and U2085 (N_2085,N_2025,N_2064);
or U2086 (N_2086,N_1929,N_1968);
and U2087 (N_2087,N_1945,N_2071);
or U2088 (N_2088,N_1935,N_1972);
and U2089 (N_2089,N_2046,N_1970);
and U2090 (N_2090,N_1938,N_1933);
nand U2091 (N_2091,N_2056,N_2019);
or U2092 (N_2092,N_2040,N_2042);
xnor U2093 (N_2093,N_1996,N_2054);
nor U2094 (N_2094,N_2001,N_2022);
and U2095 (N_2095,N_1956,N_2045);
xor U2096 (N_2096,N_1947,N_1942);
nor U2097 (N_2097,N_1937,N_2038);
xnor U2098 (N_2098,N_1961,N_1959);
nor U2099 (N_2099,N_2049,N_2048);
or U2100 (N_2100,N_2012,N_1967);
nand U2101 (N_2101,N_2004,N_2053);
nand U2102 (N_2102,N_2047,N_1999);
nor U2103 (N_2103,N_2073,N_2075);
and U2104 (N_2104,N_1986,N_1983);
and U2105 (N_2105,N_1994,N_2060);
and U2106 (N_2106,N_2015,N_1931);
nor U2107 (N_2107,N_1982,N_2070);
and U2108 (N_2108,N_2062,N_1988);
nor U2109 (N_2109,N_1925,N_1997);
nand U2110 (N_2110,N_2039,N_2020);
and U2111 (N_2111,N_2069,N_1985);
xor U2112 (N_2112,N_2065,N_2074);
and U2113 (N_2113,N_2051,N_2063);
xor U2114 (N_2114,N_2072,N_1940);
or U2115 (N_2115,N_2006,N_1964);
xnor U2116 (N_2116,N_2021,N_1941);
and U2117 (N_2117,N_2059,N_2052);
xor U2118 (N_2118,N_1990,N_1963);
nor U2119 (N_2119,N_2011,N_1950);
and U2120 (N_2120,N_2032,N_1966);
and U2121 (N_2121,N_1946,N_2033);
nor U2122 (N_2122,N_1939,N_2068);
nand U2123 (N_2123,N_1930,N_2000);
nand U2124 (N_2124,N_2061,N_2041);
and U2125 (N_2125,N_1971,N_1974);
nand U2126 (N_2126,N_2077,N_1998);
and U2127 (N_2127,N_1952,N_2009);
or U2128 (N_2128,N_2037,N_1977);
and U2129 (N_2129,N_1920,N_2058);
or U2130 (N_2130,N_1922,N_2031);
xor U2131 (N_2131,N_1989,N_2014);
or U2132 (N_2132,N_2023,N_2028);
or U2133 (N_2133,N_1973,N_1965);
and U2134 (N_2134,N_1924,N_1944);
nor U2135 (N_2135,N_2044,N_2067);
or U2136 (N_2136,N_1955,N_1979);
nand U2137 (N_2137,N_1934,N_1958);
and U2138 (N_2138,N_2030,N_2050);
or U2139 (N_2139,N_1984,N_2003);
and U2140 (N_2140,N_2029,N_1943);
xnor U2141 (N_2141,N_1954,N_2078);
nand U2142 (N_2142,N_1960,N_1991);
xor U2143 (N_2143,N_1923,N_2034);
and U2144 (N_2144,N_2013,N_2005);
and U2145 (N_2145,N_2008,N_1957);
or U2146 (N_2146,N_1949,N_2035);
xor U2147 (N_2147,N_2017,N_1953);
nor U2148 (N_2148,N_1969,N_1927);
or U2149 (N_2149,N_2036,N_1975);
nand U2150 (N_2150,N_1987,N_1995);
or U2151 (N_2151,N_1928,N_1981);
nor U2152 (N_2152,N_1962,N_2024);
nor U2153 (N_2153,N_2043,N_1932);
and U2154 (N_2154,N_2002,N_1978);
nand U2155 (N_2155,N_1926,N_2057);
or U2156 (N_2156,N_2027,N_1936);
nand U2157 (N_2157,N_2018,N_2016);
xnor U2158 (N_2158,N_2026,N_1993);
xnor U2159 (N_2159,N_2076,N_2079);
nand U2160 (N_2160,N_1950,N_1970);
nor U2161 (N_2161,N_2018,N_2019);
xnor U2162 (N_2162,N_1944,N_2070);
nand U2163 (N_2163,N_2008,N_1989);
or U2164 (N_2164,N_1985,N_2047);
xnor U2165 (N_2165,N_2014,N_1962);
nor U2166 (N_2166,N_2045,N_1949);
and U2167 (N_2167,N_2014,N_1982);
xor U2168 (N_2168,N_1923,N_1957);
nor U2169 (N_2169,N_2055,N_1934);
nor U2170 (N_2170,N_2015,N_1954);
xor U2171 (N_2171,N_1999,N_2042);
xnor U2172 (N_2172,N_1965,N_1926);
nor U2173 (N_2173,N_1958,N_2035);
xor U2174 (N_2174,N_1951,N_2014);
xnor U2175 (N_2175,N_2042,N_1988);
xor U2176 (N_2176,N_2036,N_1983);
or U2177 (N_2177,N_1924,N_2006);
and U2178 (N_2178,N_1947,N_2065);
nand U2179 (N_2179,N_2030,N_1931);
and U2180 (N_2180,N_1960,N_2050);
nand U2181 (N_2181,N_2024,N_2021);
and U2182 (N_2182,N_1983,N_2064);
or U2183 (N_2183,N_1956,N_2030);
and U2184 (N_2184,N_1955,N_1984);
or U2185 (N_2185,N_1949,N_2036);
nand U2186 (N_2186,N_1977,N_1932);
xnor U2187 (N_2187,N_1964,N_1998);
xnor U2188 (N_2188,N_2051,N_1959);
nor U2189 (N_2189,N_1964,N_1983);
or U2190 (N_2190,N_2052,N_1999);
nor U2191 (N_2191,N_2056,N_1939);
and U2192 (N_2192,N_1967,N_1981);
and U2193 (N_2193,N_1927,N_1975);
xor U2194 (N_2194,N_1993,N_2033);
and U2195 (N_2195,N_2058,N_2053);
and U2196 (N_2196,N_1946,N_2059);
or U2197 (N_2197,N_2078,N_2072);
nand U2198 (N_2198,N_2071,N_2056);
nor U2199 (N_2199,N_2062,N_2053);
and U2200 (N_2200,N_2044,N_1935);
nand U2201 (N_2201,N_1957,N_1944);
and U2202 (N_2202,N_1976,N_2010);
and U2203 (N_2203,N_2070,N_2012);
and U2204 (N_2204,N_1986,N_1958);
nor U2205 (N_2205,N_1954,N_2019);
nand U2206 (N_2206,N_1939,N_2012);
or U2207 (N_2207,N_2019,N_2021);
and U2208 (N_2208,N_1922,N_1971);
nor U2209 (N_2209,N_1932,N_1927);
and U2210 (N_2210,N_2017,N_1980);
or U2211 (N_2211,N_2052,N_1945);
or U2212 (N_2212,N_1995,N_2070);
nand U2213 (N_2213,N_1941,N_2030);
nand U2214 (N_2214,N_1957,N_2020);
xor U2215 (N_2215,N_1946,N_2069);
and U2216 (N_2216,N_1958,N_2061);
or U2217 (N_2217,N_2047,N_1960);
xnor U2218 (N_2218,N_2055,N_2075);
and U2219 (N_2219,N_1998,N_2012);
xnor U2220 (N_2220,N_2033,N_1962);
xor U2221 (N_2221,N_2053,N_1971);
and U2222 (N_2222,N_2061,N_2004);
and U2223 (N_2223,N_1996,N_1941);
nor U2224 (N_2224,N_2009,N_2040);
and U2225 (N_2225,N_2008,N_1932);
nand U2226 (N_2226,N_2030,N_1943);
and U2227 (N_2227,N_2001,N_1932);
or U2228 (N_2228,N_1975,N_2053);
and U2229 (N_2229,N_1959,N_1927);
xnor U2230 (N_2230,N_1964,N_2019);
or U2231 (N_2231,N_1963,N_1954);
nor U2232 (N_2232,N_2000,N_2047);
or U2233 (N_2233,N_1972,N_1953);
nor U2234 (N_2234,N_2075,N_1961);
nor U2235 (N_2235,N_2068,N_2028);
or U2236 (N_2236,N_2025,N_2061);
nor U2237 (N_2237,N_1963,N_2039);
xnor U2238 (N_2238,N_1994,N_2034);
and U2239 (N_2239,N_2058,N_1977);
nor U2240 (N_2240,N_2154,N_2223);
and U2241 (N_2241,N_2215,N_2186);
xnor U2242 (N_2242,N_2220,N_2172);
xor U2243 (N_2243,N_2132,N_2127);
nand U2244 (N_2244,N_2135,N_2123);
nand U2245 (N_2245,N_2221,N_2149);
nand U2246 (N_2246,N_2128,N_2145);
nor U2247 (N_2247,N_2179,N_2089);
or U2248 (N_2248,N_2110,N_2239);
or U2249 (N_2249,N_2126,N_2093);
nand U2250 (N_2250,N_2109,N_2140);
nand U2251 (N_2251,N_2171,N_2102);
nand U2252 (N_2252,N_2119,N_2105);
nand U2253 (N_2253,N_2118,N_2111);
xor U2254 (N_2254,N_2116,N_2174);
nor U2255 (N_2255,N_2104,N_2133);
or U2256 (N_2256,N_2196,N_2148);
and U2257 (N_2257,N_2086,N_2081);
and U2258 (N_2258,N_2165,N_2184);
or U2259 (N_2259,N_2107,N_2214);
nor U2260 (N_2260,N_2122,N_2146);
nand U2261 (N_2261,N_2235,N_2182);
nand U2262 (N_2262,N_2142,N_2189);
nor U2263 (N_2263,N_2230,N_2229);
and U2264 (N_2264,N_2178,N_2129);
or U2265 (N_2265,N_2151,N_2117);
nand U2266 (N_2266,N_2156,N_2167);
or U2267 (N_2267,N_2098,N_2091);
xor U2268 (N_2268,N_2159,N_2187);
and U2269 (N_2269,N_2198,N_2180);
and U2270 (N_2270,N_2108,N_2099);
and U2271 (N_2271,N_2203,N_2100);
and U2272 (N_2272,N_2193,N_2088);
nor U2273 (N_2273,N_2124,N_2188);
or U2274 (N_2274,N_2197,N_2219);
nand U2275 (N_2275,N_2202,N_2094);
nor U2276 (N_2276,N_2103,N_2101);
or U2277 (N_2277,N_2225,N_2087);
or U2278 (N_2278,N_2194,N_2080);
nand U2279 (N_2279,N_2169,N_2224);
and U2280 (N_2280,N_2195,N_2160);
xor U2281 (N_2281,N_2238,N_2209);
nand U2282 (N_2282,N_2113,N_2084);
and U2283 (N_2283,N_2192,N_2125);
nor U2284 (N_2284,N_2153,N_2161);
nand U2285 (N_2285,N_2207,N_2152);
and U2286 (N_2286,N_2232,N_2106);
nor U2287 (N_2287,N_2082,N_2211);
xor U2288 (N_2288,N_2096,N_2085);
xor U2289 (N_2289,N_2181,N_2204);
or U2290 (N_2290,N_2206,N_2095);
and U2291 (N_2291,N_2175,N_2083);
or U2292 (N_2292,N_2176,N_2114);
nand U2293 (N_2293,N_2158,N_2183);
nand U2294 (N_2294,N_2228,N_2139);
xor U2295 (N_2295,N_2130,N_2155);
or U2296 (N_2296,N_2097,N_2164);
nor U2297 (N_2297,N_2162,N_2138);
xor U2298 (N_2298,N_2210,N_2163);
or U2299 (N_2299,N_2143,N_2137);
nand U2300 (N_2300,N_2136,N_2121);
or U2301 (N_2301,N_2157,N_2191);
nand U2302 (N_2302,N_2205,N_2234);
xor U2303 (N_2303,N_2199,N_2190);
nor U2304 (N_2304,N_2227,N_2144);
xor U2305 (N_2305,N_2201,N_2115);
nor U2306 (N_2306,N_2173,N_2185);
nor U2307 (N_2307,N_2231,N_2131);
and U2308 (N_2308,N_2208,N_2150);
or U2309 (N_2309,N_2236,N_2177);
and U2310 (N_2310,N_2213,N_2168);
and U2311 (N_2311,N_2090,N_2134);
xnor U2312 (N_2312,N_2222,N_2237);
nand U2313 (N_2313,N_2120,N_2217);
nor U2314 (N_2314,N_2112,N_2233);
nor U2315 (N_2315,N_2218,N_2147);
nor U2316 (N_2316,N_2226,N_2166);
or U2317 (N_2317,N_2092,N_2141);
and U2318 (N_2318,N_2216,N_2170);
and U2319 (N_2319,N_2212,N_2200);
nor U2320 (N_2320,N_2188,N_2081);
xnor U2321 (N_2321,N_2152,N_2119);
or U2322 (N_2322,N_2128,N_2104);
nor U2323 (N_2323,N_2116,N_2080);
or U2324 (N_2324,N_2236,N_2110);
nor U2325 (N_2325,N_2184,N_2147);
and U2326 (N_2326,N_2167,N_2160);
nand U2327 (N_2327,N_2189,N_2201);
xor U2328 (N_2328,N_2142,N_2195);
xnor U2329 (N_2329,N_2165,N_2210);
or U2330 (N_2330,N_2183,N_2106);
xnor U2331 (N_2331,N_2104,N_2210);
xnor U2332 (N_2332,N_2214,N_2090);
or U2333 (N_2333,N_2203,N_2157);
and U2334 (N_2334,N_2149,N_2224);
xnor U2335 (N_2335,N_2209,N_2196);
or U2336 (N_2336,N_2148,N_2080);
nand U2337 (N_2337,N_2222,N_2155);
or U2338 (N_2338,N_2103,N_2132);
nand U2339 (N_2339,N_2232,N_2172);
nand U2340 (N_2340,N_2101,N_2210);
or U2341 (N_2341,N_2211,N_2197);
nor U2342 (N_2342,N_2184,N_2188);
nor U2343 (N_2343,N_2171,N_2117);
nand U2344 (N_2344,N_2202,N_2088);
nor U2345 (N_2345,N_2230,N_2191);
nor U2346 (N_2346,N_2108,N_2237);
nor U2347 (N_2347,N_2161,N_2172);
or U2348 (N_2348,N_2216,N_2148);
and U2349 (N_2349,N_2130,N_2235);
and U2350 (N_2350,N_2132,N_2128);
nand U2351 (N_2351,N_2119,N_2229);
nand U2352 (N_2352,N_2140,N_2112);
nand U2353 (N_2353,N_2196,N_2150);
xnor U2354 (N_2354,N_2136,N_2084);
nand U2355 (N_2355,N_2093,N_2217);
and U2356 (N_2356,N_2140,N_2199);
nand U2357 (N_2357,N_2082,N_2180);
and U2358 (N_2358,N_2157,N_2171);
xnor U2359 (N_2359,N_2170,N_2212);
xor U2360 (N_2360,N_2155,N_2146);
nand U2361 (N_2361,N_2157,N_2094);
and U2362 (N_2362,N_2235,N_2080);
nor U2363 (N_2363,N_2212,N_2173);
nand U2364 (N_2364,N_2136,N_2207);
nor U2365 (N_2365,N_2086,N_2106);
nand U2366 (N_2366,N_2210,N_2167);
or U2367 (N_2367,N_2112,N_2094);
nor U2368 (N_2368,N_2149,N_2198);
or U2369 (N_2369,N_2174,N_2092);
and U2370 (N_2370,N_2235,N_2232);
and U2371 (N_2371,N_2210,N_2214);
xor U2372 (N_2372,N_2193,N_2084);
nand U2373 (N_2373,N_2215,N_2183);
and U2374 (N_2374,N_2080,N_2085);
xnor U2375 (N_2375,N_2144,N_2205);
and U2376 (N_2376,N_2188,N_2117);
and U2377 (N_2377,N_2152,N_2159);
nand U2378 (N_2378,N_2127,N_2161);
nand U2379 (N_2379,N_2121,N_2087);
xnor U2380 (N_2380,N_2130,N_2126);
and U2381 (N_2381,N_2139,N_2165);
xor U2382 (N_2382,N_2185,N_2202);
xnor U2383 (N_2383,N_2217,N_2094);
nand U2384 (N_2384,N_2236,N_2134);
nor U2385 (N_2385,N_2167,N_2180);
xnor U2386 (N_2386,N_2106,N_2142);
and U2387 (N_2387,N_2084,N_2094);
nor U2388 (N_2388,N_2082,N_2090);
xor U2389 (N_2389,N_2229,N_2215);
or U2390 (N_2390,N_2143,N_2161);
nand U2391 (N_2391,N_2174,N_2096);
and U2392 (N_2392,N_2122,N_2152);
xor U2393 (N_2393,N_2110,N_2170);
xor U2394 (N_2394,N_2096,N_2234);
nor U2395 (N_2395,N_2117,N_2217);
xor U2396 (N_2396,N_2211,N_2080);
or U2397 (N_2397,N_2155,N_2166);
nor U2398 (N_2398,N_2120,N_2140);
and U2399 (N_2399,N_2095,N_2168);
or U2400 (N_2400,N_2242,N_2260);
and U2401 (N_2401,N_2286,N_2377);
nand U2402 (N_2402,N_2290,N_2271);
and U2403 (N_2403,N_2259,N_2375);
nor U2404 (N_2404,N_2305,N_2276);
xnor U2405 (N_2405,N_2319,N_2398);
nor U2406 (N_2406,N_2334,N_2399);
nand U2407 (N_2407,N_2279,N_2310);
and U2408 (N_2408,N_2243,N_2254);
nor U2409 (N_2409,N_2397,N_2292);
or U2410 (N_2410,N_2371,N_2385);
nor U2411 (N_2411,N_2341,N_2318);
or U2412 (N_2412,N_2252,N_2246);
and U2413 (N_2413,N_2258,N_2280);
or U2414 (N_2414,N_2308,N_2351);
and U2415 (N_2415,N_2265,N_2391);
or U2416 (N_2416,N_2241,N_2342);
xor U2417 (N_2417,N_2302,N_2326);
nand U2418 (N_2418,N_2277,N_2272);
and U2419 (N_2419,N_2379,N_2285);
nand U2420 (N_2420,N_2328,N_2329);
nand U2421 (N_2421,N_2366,N_2293);
or U2422 (N_2422,N_2360,N_2386);
and U2423 (N_2423,N_2274,N_2257);
xor U2424 (N_2424,N_2253,N_2313);
and U2425 (N_2425,N_2343,N_2336);
and U2426 (N_2426,N_2381,N_2300);
and U2427 (N_2427,N_2370,N_2352);
nand U2428 (N_2428,N_2369,N_2340);
xnor U2429 (N_2429,N_2382,N_2393);
or U2430 (N_2430,N_2345,N_2387);
xnor U2431 (N_2431,N_2291,N_2301);
and U2432 (N_2432,N_2284,N_2298);
nand U2433 (N_2433,N_2354,N_2268);
nand U2434 (N_2434,N_2347,N_2339);
nor U2435 (N_2435,N_2270,N_2294);
nand U2436 (N_2436,N_2383,N_2333);
nor U2437 (N_2437,N_2250,N_2309);
nand U2438 (N_2438,N_2365,N_2349);
or U2439 (N_2439,N_2299,N_2262);
or U2440 (N_2440,N_2251,N_2395);
and U2441 (N_2441,N_2282,N_2331);
nand U2442 (N_2442,N_2353,N_2304);
xnor U2443 (N_2443,N_2364,N_2368);
xnor U2444 (N_2444,N_2337,N_2323);
xor U2445 (N_2445,N_2330,N_2240);
nor U2446 (N_2446,N_2255,N_2267);
nand U2447 (N_2447,N_2357,N_2263);
xnor U2448 (N_2448,N_2380,N_2346);
or U2449 (N_2449,N_2269,N_2356);
and U2450 (N_2450,N_2332,N_2278);
nand U2451 (N_2451,N_2317,N_2358);
and U2452 (N_2452,N_2256,N_2350);
or U2453 (N_2453,N_2359,N_2314);
xnor U2454 (N_2454,N_2245,N_2281);
nand U2455 (N_2455,N_2361,N_2322);
or U2456 (N_2456,N_2372,N_2320);
or U2457 (N_2457,N_2376,N_2311);
and U2458 (N_2458,N_2249,N_2384);
nor U2459 (N_2459,N_2344,N_2287);
and U2460 (N_2460,N_2355,N_2325);
and U2461 (N_2461,N_2348,N_2316);
or U2462 (N_2462,N_2266,N_2321);
nand U2463 (N_2463,N_2362,N_2283);
nand U2464 (N_2464,N_2288,N_2275);
nor U2465 (N_2465,N_2295,N_2248);
and U2466 (N_2466,N_2367,N_2307);
nand U2467 (N_2467,N_2327,N_2303);
xnor U2468 (N_2468,N_2273,N_2389);
or U2469 (N_2469,N_2264,N_2374);
and U2470 (N_2470,N_2388,N_2363);
nand U2471 (N_2471,N_2244,N_2289);
nand U2472 (N_2472,N_2306,N_2392);
or U2473 (N_2473,N_2247,N_2394);
xor U2474 (N_2474,N_2261,N_2312);
nand U2475 (N_2475,N_2378,N_2335);
or U2476 (N_2476,N_2324,N_2297);
nand U2477 (N_2477,N_2373,N_2396);
nor U2478 (N_2478,N_2296,N_2338);
or U2479 (N_2479,N_2390,N_2315);
nor U2480 (N_2480,N_2312,N_2308);
and U2481 (N_2481,N_2254,N_2291);
nor U2482 (N_2482,N_2288,N_2357);
nor U2483 (N_2483,N_2267,N_2294);
or U2484 (N_2484,N_2282,N_2340);
nor U2485 (N_2485,N_2312,N_2272);
and U2486 (N_2486,N_2306,N_2280);
nor U2487 (N_2487,N_2354,N_2263);
xnor U2488 (N_2488,N_2334,N_2307);
xor U2489 (N_2489,N_2397,N_2333);
nor U2490 (N_2490,N_2308,N_2288);
nor U2491 (N_2491,N_2379,N_2393);
xnor U2492 (N_2492,N_2311,N_2352);
and U2493 (N_2493,N_2333,N_2325);
xnor U2494 (N_2494,N_2295,N_2328);
or U2495 (N_2495,N_2335,N_2368);
xnor U2496 (N_2496,N_2399,N_2327);
nand U2497 (N_2497,N_2292,N_2312);
nand U2498 (N_2498,N_2331,N_2295);
nor U2499 (N_2499,N_2255,N_2328);
nor U2500 (N_2500,N_2301,N_2388);
nor U2501 (N_2501,N_2255,N_2341);
nand U2502 (N_2502,N_2290,N_2339);
nor U2503 (N_2503,N_2289,N_2364);
or U2504 (N_2504,N_2357,N_2338);
and U2505 (N_2505,N_2292,N_2346);
xor U2506 (N_2506,N_2257,N_2381);
or U2507 (N_2507,N_2364,N_2247);
xnor U2508 (N_2508,N_2247,N_2256);
and U2509 (N_2509,N_2359,N_2291);
nand U2510 (N_2510,N_2367,N_2365);
nor U2511 (N_2511,N_2367,N_2318);
or U2512 (N_2512,N_2357,N_2351);
xnor U2513 (N_2513,N_2333,N_2240);
and U2514 (N_2514,N_2263,N_2313);
and U2515 (N_2515,N_2266,N_2350);
xor U2516 (N_2516,N_2263,N_2267);
or U2517 (N_2517,N_2261,N_2393);
xor U2518 (N_2518,N_2334,N_2367);
and U2519 (N_2519,N_2333,N_2329);
xnor U2520 (N_2520,N_2357,N_2253);
or U2521 (N_2521,N_2240,N_2385);
nand U2522 (N_2522,N_2272,N_2354);
or U2523 (N_2523,N_2330,N_2374);
nor U2524 (N_2524,N_2338,N_2275);
nor U2525 (N_2525,N_2292,N_2386);
nor U2526 (N_2526,N_2330,N_2287);
or U2527 (N_2527,N_2269,N_2363);
nor U2528 (N_2528,N_2308,N_2343);
xnor U2529 (N_2529,N_2242,N_2328);
nand U2530 (N_2530,N_2266,N_2338);
xnor U2531 (N_2531,N_2323,N_2352);
and U2532 (N_2532,N_2243,N_2295);
and U2533 (N_2533,N_2278,N_2341);
nand U2534 (N_2534,N_2245,N_2250);
and U2535 (N_2535,N_2324,N_2274);
nor U2536 (N_2536,N_2261,N_2337);
nand U2537 (N_2537,N_2385,N_2364);
nor U2538 (N_2538,N_2282,N_2380);
nand U2539 (N_2539,N_2312,N_2252);
xnor U2540 (N_2540,N_2292,N_2302);
or U2541 (N_2541,N_2386,N_2334);
nor U2542 (N_2542,N_2246,N_2350);
nand U2543 (N_2543,N_2305,N_2300);
nor U2544 (N_2544,N_2268,N_2253);
nand U2545 (N_2545,N_2329,N_2294);
or U2546 (N_2546,N_2278,N_2319);
nand U2547 (N_2547,N_2281,N_2390);
xor U2548 (N_2548,N_2386,N_2284);
or U2549 (N_2549,N_2344,N_2378);
nand U2550 (N_2550,N_2393,N_2244);
xor U2551 (N_2551,N_2352,N_2328);
or U2552 (N_2552,N_2386,N_2315);
or U2553 (N_2553,N_2280,N_2345);
and U2554 (N_2554,N_2286,N_2297);
or U2555 (N_2555,N_2274,N_2353);
nor U2556 (N_2556,N_2378,N_2377);
or U2557 (N_2557,N_2329,N_2318);
nor U2558 (N_2558,N_2242,N_2283);
and U2559 (N_2559,N_2279,N_2265);
and U2560 (N_2560,N_2466,N_2504);
nor U2561 (N_2561,N_2403,N_2489);
nand U2562 (N_2562,N_2427,N_2496);
xnor U2563 (N_2563,N_2513,N_2495);
xor U2564 (N_2564,N_2436,N_2490);
nor U2565 (N_2565,N_2525,N_2470);
and U2566 (N_2566,N_2408,N_2558);
nand U2567 (N_2567,N_2528,N_2500);
and U2568 (N_2568,N_2417,N_2531);
xnor U2569 (N_2569,N_2477,N_2523);
xnor U2570 (N_2570,N_2412,N_2518);
nor U2571 (N_2571,N_2454,N_2494);
and U2572 (N_2572,N_2406,N_2467);
xor U2573 (N_2573,N_2509,N_2450);
xor U2574 (N_2574,N_2468,N_2459);
nor U2575 (N_2575,N_2542,N_2510);
or U2576 (N_2576,N_2448,N_2441);
nor U2577 (N_2577,N_2455,N_2514);
nand U2578 (N_2578,N_2550,N_2551);
and U2579 (N_2579,N_2407,N_2533);
nor U2580 (N_2580,N_2405,N_2473);
xor U2581 (N_2581,N_2440,N_2430);
nor U2582 (N_2582,N_2486,N_2425);
nor U2583 (N_2583,N_2458,N_2487);
xor U2584 (N_2584,N_2520,N_2445);
nand U2585 (N_2585,N_2439,N_2535);
or U2586 (N_2586,N_2422,N_2534);
xnor U2587 (N_2587,N_2540,N_2492);
xor U2588 (N_2588,N_2442,N_2471);
nor U2589 (N_2589,N_2474,N_2546);
xor U2590 (N_2590,N_2443,N_2512);
and U2591 (N_2591,N_2508,N_2544);
xnor U2592 (N_2592,N_2482,N_2515);
or U2593 (N_2593,N_2507,N_2538);
nor U2594 (N_2594,N_2400,N_2497);
xnor U2595 (N_2595,N_2451,N_2553);
nor U2596 (N_2596,N_2556,N_2522);
nand U2597 (N_2597,N_2545,N_2456);
or U2598 (N_2598,N_2438,N_2462);
xor U2599 (N_2599,N_2472,N_2409);
or U2600 (N_2600,N_2429,N_2552);
nand U2601 (N_2601,N_2418,N_2463);
and U2602 (N_2602,N_2452,N_2447);
nor U2603 (N_2603,N_2461,N_2506);
nor U2604 (N_2604,N_2457,N_2464);
and U2605 (N_2605,N_2401,N_2435);
nor U2606 (N_2606,N_2413,N_2559);
xnor U2607 (N_2607,N_2505,N_2499);
nand U2608 (N_2608,N_2475,N_2502);
and U2609 (N_2609,N_2530,N_2532);
nor U2610 (N_2610,N_2449,N_2537);
nor U2611 (N_2611,N_2423,N_2410);
xnor U2612 (N_2612,N_2503,N_2516);
and U2613 (N_2613,N_2453,N_2424);
and U2614 (N_2614,N_2543,N_2488);
nor U2615 (N_2615,N_2541,N_2517);
and U2616 (N_2616,N_2511,N_2527);
and U2617 (N_2617,N_2444,N_2493);
xnor U2618 (N_2618,N_2557,N_2549);
xnor U2619 (N_2619,N_2555,N_2434);
xnor U2620 (N_2620,N_2481,N_2469);
and U2621 (N_2621,N_2433,N_2524);
and U2622 (N_2622,N_2491,N_2404);
and U2623 (N_2623,N_2446,N_2547);
or U2624 (N_2624,N_2411,N_2414);
nand U2625 (N_2625,N_2465,N_2519);
nand U2626 (N_2626,N_2501,N_2526);
or U2627 (N_2627,N_2478,N_2480);
nor U2628 (N_2628,N_2416,N_2432);
nor U2629 (N_2629,N_2419,N_2415);
nor U2630 (N_2630,N_2421,N_2521);
xnor U2631 (N_2631,N_2437,N_2548);
nor U2632 (N_2632,N_2420,N_2426);
nand U2633 (N_2633,N_2402,N_2460);
or U2634 (N_2634,N_2536,N_2554);
and U2635 (N_2635,N_2539,N_2483);
nor U2636 (N_2636,N_2484,N_2529);
and U2637 (N_2637,N_2428,N_2498);
and U2638 (N_2638,N_2476,N_2431);
and U2639 (N_2639,N_2485,N_2479);
or U2640 (N_2640,N_2539,N_2442);
and U2641 (N_2641,N_2419,N_2542);
nor U2642 (N_2642,N_2530,N_2559);
and U2643 (N_2643,N_2454,N_2530);
xnor U2644 (N_2644,N_2476,N_2411);
nand U2645 (N_2645,N_2544,N_2423);
or U2646 (N_2646,N_2502,N_2555);
or U2647 (N_2647,N_2547,N_2542);
nand U2648 (N_2648,N_2483,N_2428);
nor U2649 (N_2649,N_2491,N_2437);
nand U2650 (N_2650,N_2528,N_2557);
xor U2651 (N_2651,N_2452,N_2411);
nor U2652 (N_2652,N_2522,N_2488);
or U2653 (N_2653,N_2473,N_2541);
and U2654 (N_2654,N_2533,N_2418);
or U2655 (N_2655,N_2437,N_2458);
and U2656 (N_2656,N_2510,N_2545);
nor U2657 (N_2657,N_2441,N_2462);
nor U2658 (N_2658,N_2538,N_2452);
nor U2659 (N_2659,N_2506,N_2416);
and U2660 (N_2660,N_2443,N_2414);
xnor U2661 (N_2661,N_2536,N_2499);
or U2662 (N_2662,N_2533,N_2401);
or U2663 (N_2663,N_2550,N_2485);
and U2664 (N_2664,N_2461,N_2415);
or U2665 (N_2665,N_2512,N_2450);
nand U2666 (N_2666,N_2496,N_2500);
and U2667 (N_2667,N_2463,N_2491);
and U2668 (N_2668,N_2415,N_2474);
and U2669 (N_2669,N_2516,N_2531);
or U2670 (N_2670,N_2511,N_2521);
and U2671 (N_2671,N_2455,N_2445);
nor U2672 (N_2672,N_2402,N_2438);
and U2673 (N_2673,N_2457,N_2499);
or U2674 (N_2674,N_2466,N_2464);
and U2675 (N_2675,N_2523,N_2411);
xnor U2676 (N_2676,N_2529,N_2462);
nor U2677 (N_2677,N_2553,N_2472);
xnor U2678 (N_2678,N_2473,N_2467);
or U2679 (N_2679,N_2440,N_2456);
and U2680 (N_2680,N_2496,N_2514);
and U2681 (N_2681,N_2491,N_2511);
nor U2682 (N_2682,N_2455,N_2463);
or U2683 (N_2683,N_2420,N_2492);
and U2684 (N_2684,N_2508,N_2550);
or U2685 (N_2685,N_2468,N_2508);
nor U2686 (N_2686,N_2551,N_2517);
or U2687 (N_2687,N_2494,N_2469);
and U2688 (N_2688,N_2528,N_2427);
and U2689 (N_2689,N_2458,N_2454);
or U2690 (N_2690,N_2452,N_2454);
xnor U2691 (N_2691,N_2454,N_2401);
nand U2692 (N_2692,N_2443,N_2473);
xnor U2693 (N_2693,N_2507,N_2546);
nand U2694 (N_2694,N_2477,N_2508);
xnor U2695 (N_2695,N_2499,N_2557);
or U2696 (N_2696,N_2497,N_2493);
and U2697 (N_2697,N_2494,N_2401);
and U2698 (N_2698,N_2409,N_2408);
or U2699 (N_2699,N_2503,N_2471);
or U2700 (N_2700,N_2504,N_2423);
nor U2701 (N_2701,N_2522,N_2448);
xor U2702 (N_2702,N_2556,N_2401);
and U2703 (N_2703,N_2484,N_2421);
and U2704 (N_2704,N_2471,N_2454);
nor U2705 (N_2705,N_2460,N_2499);
nand U2706 (N_2706,N_2425,N_2532);
nor U2707 (N_2707,N_2448,N_2515);
nand U2708 (N_2708,N_2478,N_2485);
or U2709 (N_2709,N_2551,N_2487);
nand U2710 (N_2710,N_2465,N_2495);
nor U2711 (N_2711,N_2428,N_2456);
and U2712 (N_2712,N_2524,N_2499);
nor U2713 (N_2713,N_2458,N_2476);
and U2714 (N_2714,N_2423,N_2456);
nor U2715 (N_2715,N_2427,N_2553);
xor U2716 (N_2716,N_2486,N_2439);
xor U2717 (N_2717,N_2480,N_2499);
nor U2718 (N_2718,N_2465,N_2445);
nand U2719 (N_2719,N_2540,N_2526);
or U2720 (N_2720,N_2642,N_2638);
nand U2721 (N_2721,N_2565,N_2719);
nand U2722 (N_2722,N_2589,N_2692);
or U2723 (N_2723,N_2569,N_2698);
and U2724 (N_2724,N_2583,N_2593);
nor U2725 (N_2725,N_2597,N_2570);
nor U2726 (N_2726,N_2685,N_2607);
or U2727 (N_2727,N_2680,N_2691);
nand U2728 (N_2728,N_2668,N_2681);
nor U2729 (N_2729,N_2711,N_2659);
or U2730 (N_2730,N_2623,N_2660);
xnor U2731 (N_2731,N_2651,N_2714);
xor U2732 (N_2732,N_2599,N_2580);
or U2733 (N_2733,N_2696,N_2641);
nand U2734 (N_2734,N_2703,N_2613);
or U2735 (N_2735,N_2713,N_2629);
xnor U2736 (N_2736,N_2591,N_2704);
and U2737 (N_2737,N_2648,N_2653);
or U2738 (N_2738,N_2602,N_2621);
or U2739 (N_2739,N_2575,N_2603);
and U2740 (N_2740,N_2630,N_2567);
and U2741 (N_2741,N_2631,N_2608);
or U2742 (N_2742,N_2665,N_2661);
nand U2743 (N_2743,N_2640,N_2586);
nand U2744 (N_2744,N_2646,N_2625);
or U2745 (N_2745,N_2611,N_2633);
nand U2746 (N_2746,N_2581,N_2652);
nor U2747 (N_2747,N_2654,N_2617);
xor U2748 (N_2748,N_2635,N_2624);
or U2749 (N_2749,N_2592,N_2715);
and U2750 (N_2750,N_2673,N_2687);
xor U2751 (N_2751,N_2573,N_2574);
nand U2752 (N_2752,N_2560,N_2644);
or U2753 (N_2753,N_2595,N_2561);
or U2754 (N_2754,N_2667,N_2582);
xor U2755 (N_2755,N_2676,N_2647);
or U2756 (N_2756,N_2701,N_2679);
nor U2757 (N_2757,N_2632,N_2643);
and U2758 (N_2758,N_2639,N_2600);
xnor U2759 (N_2759,N_2709,N_2699);
or U2760 (N_2760,N_2587,N_2578);
xor U2761 (N_2761,N_2590,N_2695);
nand U2762 (N_2762,N_2664,N_2585);
nand U2763 (N_2763,N_2666,N_2572);
nor U2764 (N_2764,N_2615,N_2628);
nand U2765 (N_2765,N_2675,N_2563);
or U2766 (N_2766,N_2707,N_2622);
nor U2767 (N_2767,N_2694,N_2657);
xor U2768 (N_2768,N_2606,N_2674);
nand U2769 (N_2769,N_2700,N_2683);
nor U2770 (N_2770,N_2618,N_2634);
and U2771 (N_2771,N_2619,N_2604);
or U2772 (N_2772,N_2568,N_2614);
nand U2773 (N_2773,N_2576,N_2658);
xnor U2774 (N_2774,N_2564,N_2690);
nand U2775 (N_2775,N_2669,N_2688);
xnor U2776 (N_2776,N_2717,N_2598);
or U2777 (N_2777,N_2571,N_2705);
nand U2778 (N_2778,N_2588,N_2689);
nor U2779 (N_2779,N_2616,N_2649);
or U2780 (N_2780,N_2718,N_2670);
nor U2781 (N_2781,N_2712,N_2702);
nand U2782 (N_2782,N_2663,N_2637);
and U2783 (N_2783,N_2636,N_2655);
or U2784 (N_2784,N_2693,N_2605);
nor U2785 (N_2785,N_2566,N_2656);
or U2786 (N_2786,N_2562,N_2682);
xor U2787 (N_2787,N_2686,N_2684);
and U2788 (N_2788,N_2672,N_2620);
and U2789 (N_2789,N_2626,N_2610);
or U2790 (N_2790,N_2671,N_2612);
nor U2791 (N_2791,N_2596,N_2645);
nand U2792 (N_2792,N_2627,N_2677);
xor U2793 (N_2793,N_2697,N_2650);
and U2794 (N_2794,N_2678,N_2577);
xnor U2795 (N_2795,N_2601,N_2662);
nor U2796 (N_2796,N_2708,N_2584);
and U2797 (N_2797,N_2706,N_2716);
or U2798 (N_2798,N_2710,N_2594);
xor U2799 (N_2799,N_2579,N_2609);
and U2800 (N_2800,N_2645,N_2586);
nor U2801 (N_2801,N_2687,N_2597);
nor U2802 (N_2802,N_2699,N_2666);
and U2803 (N_2803,N_2633,N_2592);
xor U2804 (N_2804,N_2562,N_2568);
and U2805 (N_2805,N_2648,N_2717);
or U2806 (N_2806,N_2610,N_2659);
and U2807 (N_2807,N_2602,N_2585);
nor U2808 (N_2808,N_2573,N_2640);
and U2809 (N_2809,N_2591,N_2602);
nand U2810 (N_2810,N_2707,N_2708);
nand U2811 (N_2811,N_2688,N_2693);
nand U2812 (N_2812,N_2687,N_2563);
and U2813 (N_2813,N_2710,N_2590);
and U2814 (N_2814,N_2589,N_2574);
nand U2815 (N_2815,N_2624,N_2636);
xnor U2816 (N_2816,N_2710,N_2617);
nand U2817 (N_2817,N_2677,N_2622);
and U2818 (N_2818,N_2705,N_2620);
nand U2819 (N_2819,N_2702,N_2633);
or U2820 (N_2820,N_2565,N_2716);
or U2821 (N_2821,N_2624,N_2585);
xor U2822 (N_2822,N_2673,N_2597);
or U2823 (N_2823,N_2591,N_2626);
xnor U2824 (N_2824,N_2578,N_2598);
or U2825 (N_2825,N_2599,N_2604);
or U2826 (N_2826,N_2641,N_2671);
nor U2827 (N_2827,N_2691,N_2577);
nand U2828 (N_2828,N_2604,N_2661);
and U2829 (N_2829,N_2659,N_2565);
and U2830 (N_2830,N_2561,N_2618);
and U2831 (N_2831,N_2617,N_2638);
nor U2832 (N_2832,N_2663,N_2575);
or U2833 (N_2833,N_2669,N_2576);
and U2834 (N_2834,N_2666,N_2684);
nor U2835 (N_2835,N_2618,N_2628);
xnor U2836 (N_2836,N_2642,N_2608);
nand U2837 (N_2837,N_2715,N_2634);
or U2838 (N_2838,N_2636,N_2576);
or U2839 (N_2839,N_2685,N_2719);
nand U2840 (N_2840,N_2701,N_2599);
xnor U2841 (N_2841,N_2705,N_2609);
or U2842 (N_2842,N_2658,N_2651);
nand U2843 (N_2843,N_2697,N_2717);
or U2844 (N_2844,N_2621,N_2641);
or U2845 (N_2845,N_2574,N_2575);
nand U2846 (N_2846,N_2631,N_2670);
or U2847 (N_2847,N_2597,N_2663);
nor U2848 (N_2848,N_2627,N_2669);
nand U2849 (N_2849,N_2708,N_2709);
nand U2850 (N_2850,N_2590,N_2616);
nor U2851 (N_2851,N_2560,N_2584);
nor U2852 (N_2852,N_2585,N_2593);
xor U2853 (N_2853,N_2710,N_2589);
and U2854 (N_2854,N_2590,N_2673);
nand U2855 (N_2855,N_2678,N_2560);
and U2856 (N_2856,N_2567,N_2660);
and U2857 (N_2857,N_2574,N_2692);
or U2858 (N_2858,N_2615,N_2708);
or U2859 (N_2859,N_2702,N_2660);
nand U2860 (N_2860,N_2716,N_2677);
xor U2861 (N_2861,N_2643,N_2703);
nor U2862 (N_2862,N_2686,N_2651);
or U2863 (N_2863,N_2617,N_2653);
xnor U2864 (N_2864,N_2594,N_2591);
xnor U2865 (N_2865,N_2684,N_2623);
xor U2866 (N_2866,N_2596,N_2708);
or U2867 (N_2867,N_2628,N_2704);
nand U2868 (N_2868,N_2613,N_2607);
and U2869 (N_2869,N_2632,N_2574);
nand U2870 (N_2870,N_2671,N_2650);
nor U2871 (N_2871,N_2688,N_2615);
and U2872 (N_2872,N_2664,N_2619);
xor U2873 (N_2873,N_2712,N_2629);
or U2874 (N_2874,N_2564,N_2688);
nand U2875 (N_2875,N_2696,N_2645);
nor U2876 (N_2876,N_2681,N_2606);
or U2877 (N_2877,N_2639,N_2701);
or U2878 (N_2878,N_2565,N_2569);
xor U2879 (N_2879,N_2701,N_2611);
and U2880 (N_2880,N_2770,N_2769);
xor U2881 (N_2881,N_2836,N_2730);
nand U2882 (N_2882,N_2849,N_2796);
xor U2883 (N_2883,N_2826,N_2794);
and U2884 (N_2884,N_2743,N_2788);
nand U2885 (N_2885,N_2821,N_2773);
nand U2886 (N_2886,N_2808,N_2732);
xnor U2887 (N_2887,N_2729,N_2725);
nand U2888 (N_2888,N_2823,N_2860);
xor U2889 (N_2889,N_2723,N_2771);
xnor U2890 (N_2890,N_2816,N_2843);
xor U2891 (N_2891,N_2840,N_2807);
nand U2892 (N_2892,N_2878,N_2870);
nor U2893 (N_2893,N_2760,N_2813);
and U2894 (N_2894,N_2797,N_2750);
or U2895 (N_2895,N_2798,N_2863);
or U2896 (N_2896,N_2765,N_2842);
nor U2897 (N_2897,N_2805,N_2772);
xor U2898 (N_2898,N_2873,N_2817);
and U2899 (N_2899,N_2833,N_2753);
and U2900 (N_2900,N_2846,N_2787);
and U2901 (N_2901,N_2825,N_2757);
nand U2902 (N_2902,N_2847,N_2830);
or U2903 (N_2903,N_2856,N_2828);
and U2904 (N_2904,N_2774,N_2800);
xnor U2905 (N_2905,N_2793,N_2744);
and U2906 (N_2906,N_2726,N_2755);
nor U2907 (N_2907,N_2754,N_2876);
nand U2908 (N_2908,N_2865,N_2792);
xor U2909 (N_2909,N_2851,N_2752);
xnor U2910 (N_2910,N_2740,N_2789);
or U2911 (N_2911,N_2837,N_2855);
or U2912 (N_2912,N_2814,N_2779);
xor U2913 (N_2913,N_2832,N_2812);
nor U2914 (N_2914,N_2791,N_2733);
or U2915 (N_2915,N_2742,N_2835);
nor U2916 (N_2916,N_2864,N_2848);
xor U2917 (N_2917,N_2766,N_2745);
nand U2918 (N_2918,N_2806,N_2871);
and U2919 (N_2919,N_2738,N_2841);
nor U2920 (N_2920,N_2721,N_2861);
and U2921 (N_2921,N_2875,N_2868);
nor U2922 (N_2922,N_2804,N_2756);
nor U2923 (N_2923,N_2751,N_2727);
and U2924 (N_2924,N_2785,N_2799);
nor U2925 (N_2925,N_2746,N_2810);
and U2926 (N_2926,N_2759,N_2831);
nand U2927 (N_2927,N_2819,N_2728);
and U2928 (N_2928,N_2786,N_2780);
or U2929 (N_2929,N_2844,N_2763);
nand U2930 (N_2930,N_2741,N_2762);
nor U2931 (N_2931,N_2839,N_2775);
and U2932 (N_2932,N_2768,N_2790);
xor U2933 (N_2933,N_2801,N_2829);
or U2934 (N_2934,N_2867,N_2777);
or U2935 (N_2935,N_2784,N_2737);
xor U2936 (N_2936,N_2815,N_2866);
nand U2937 (N_2937,N_2879,N_2852);
nand U2938 (N_2938,N_2724,N_2874);
nor U2939 (N_2939,N_2736,N_2749);
nor U2940 (N_2940,N_2822,N_2767);
and U2941 (N_2941,N_2845,N_2720);
xor U2942 (N_2942,N_2781,N_2783);
and U2943 (N_2943,N_2869,N_2758);
nand U2944 (N_2944,N_2877,N_2802);
nand U2945 (N_2945,N_2827,N_2834);
or U2946 (N_2946,N_2778,N_2818);
or U2947 (N_2947,N_2748,N_2820);
xor U2948 (N_2948,N_2853,N_2862);
nand U2949 (N_2949,N_2734,N_2859);
nand U2950 (N_2950,N_2722,N_2857);
xor U2951 (N_2951,N_2776,N_2854);
and U2952 (N_2952,N_2803,N_2731);
or U2953 (N_2953,N_2824,N_2764);
or U2954 (N_2954,N_2735,N_2739);
nor U2955 (N_2955,N_2761,N_2858);
nor U2956 (N_2956,N_2811,N_2809);
and U2957 (N_2957,N_2838,N_2872);
nor U2958 (N_2958,N_2747,N_2782);
nand U2959 (N_2959,N_2795,N_2850);
nor U2960 (N_2960,N_2851,N_2740);
nor U2961 (N_2961,N_2787,N_2775);
or U2962 (N_2962,N_2775,N_2845);
xor U2963 (N_2963,N_2780,N_2810);
xnor U2964 (N_2964,N_2817,N_2854);
xnor U2965 (N_2965,N_2858,N_2758);
xor U2966 (N_2966,N_2787,N_2743);
and U2967 (N_2967,N_2783,N_2830);
nand U2968 (N_2968,N_2765,N_2722);
or U2969 (N_2969,N_2803,N_2781);
or U2970 (N_2970,N_2805,N_2878);
xnor U2971 (N_2971,N_2758,N_2839);
or U2972 (N_2972,N_2768,N_2758);
nor U2973 (N_2973,N_2743,N_2752);
and U2974 (N_2974,N_2749,N_2823);
nor U2975 (N_2975,N_2834,N_2739);
or U2976 (N_2976,N_2721,N_2736);
or U2977 (N_2977,N_2812,N_2868);
nand U2978 (N_2978,N_2852,N_2878);
and U2979 (N_2979,N_2794,N_2761);
nor U2980 (N_2980,N_2799,N_2873);
xor U2981 (N_2981,N_2788,N_2777);
or U2982 (N_2982,N_2798,N_2828);
nor U2983 (N_2983,N_2824,N_2808);
or U2984 (N_2984,N_2741,N_2790);
or U2985 (N_2985,N_2824,N_2730);
and U2986 (N_2986,N_2813,N_2735);
xor U2987 (N_2987,N_2855,N_2865);
or U2988 (N_2988,N_2805,N_2754);
or U2989 (N_2989,N_2795,N_2838);
nand U2990 (N_2990,N_2761,N_2738);
nor U2991 (N_2991,N_2782,N_2734);
nor U2992 (N_2992,N_2745,N_2821);
or U2993 (N_2993,N_2767,N_2874);
xor U2994 (N_2994,N_2869,N_2865);
and U2995 (N_2995,N_2769,N_2816);
or U2996 (N_2996,N_2866,N_2816);
nand U2997 (N_2997,N_2865,N_2734);
nand U2998 (N_2998,N_2763,N_2789);
nand U2999 (N_2999,N_2840,N_2797);
and U3000 (N_3000,N_2765,N_2864);
nor U3001 (N_3001,N_2753,N_2761);
nand U3002 (N_3002,N_2802,N_2748);
xor U3003 (N_3003,N_2827,N_2868);
nor U3004 (N_3004,N_2773,N_2833);
and U3005 (N_3005,N_2732,N_2753);
xnor U3006 (N_3006,N_2796,N_2844);
or U3007 (N_3007,N_2877,N_2876);
nand U3008 (N_3008,N_2836,N_2824);
xor U3009 (N_3009,N_2759,N_2861);
and U3010 (N_3010,N_2806,N_2720);
nor U3011 (N_3011,N_2759,N_2811);
or U3012 (N_3012,N_2780,N_2871);
and U3013 (N_3013,N_2729,N_2764);
xor U3014 (N_3014,N_2737,N_2726);
or U3015 (N_3015,N_2742,N_2735);
xnor U3016 (N_3016,N_2785,N_2750);
and U3017 (N_3017,N_2844,N_2824);
and U3018 (N_3018,N_2833,N_2730);
and U3019 (N_3019,N_2758,N_2729);
and U3020 (N_3020,N_2786,N_2839);
xnor U3021 (N_3021,N_2797,N_2862);
and U3022 (N_3022,N_2757,N_2809);
nor U3023 (N_3023,N_2763,N_2876);
or U3024 (N_3024,N_2743,N_2775);
or U3025 (N_3025,N_2845,N_2810);
nor U3026 (N_3026,N_2802,N_2815);
nand U3027 (N_3027,N_2871,N_2861);
and U3028 (N_3028,N_2744,N_2769);
xnor U3029 (N_3029,N_2802,N_2791);
xor U3030 (N_3030,N_2755,N_2795);
xor U3031 (N_3031,N_2862,N_2851);
nand U3032 (N_3032,N_2725,N_2747);
nor U3033 (N_3033,N_2753,N_2842);
xnor U3034 (N_3034,N_2755,N_2824);
or U3035 (N_3035,N_2734,N_2863);
nand U3036 (N_3036,N_2795,N_2798);
or U3037 (N_3037,N_2801,N_2820);
or U3038 (N_3038,N_2779,N_2824);
and U3039 (N_3039,N_2797,N_2859);
nor U3040 (N_3040,N_2897,N_3024);
or U3041 (N_3041,N_3004,N_2934);
or U3042 (N_3042,N_2901,N_2899);
or U3043 (N_3043,N_2969,N_2959);
or U3044 (N_3044,N_2929,N_2990);
nor U3045 (N_3045,N_2997,N_2960);
nor U3046 (N_3046,N_2905,N_3036);
or U3047 (N_3047,N_3006,N_2946);
or U3048 (N_3048,N_2940,N_3014);
and U3049 (N_3049,N_2956,N_3022);
nand U3050 (N_3050,N_2936,N_2916);
xnor U3051 (N_3051,N_2998,N_2935);
and U3052 (N_3052,N_3032,N_3026);
nand U3053 (N_3053,N_3016,N_2925);
xnor U3054 (N_3054,N_2895,N_2971);
nor U3055 (N_3055,N_2970,N_2930);
and U3056 (N_3056,N_2993,N_3003);
xor U3057 (N_3057,N_2915,N_2989);
nor U3058 (N_3058,N_2954,N_3000);
xor U3059 (N_3059,N_2903,N_2928);
nor U3060 (N_3060,N_2986,N_2952);
or U3061 (N_3061,N_2923,N_2947);
nor U3062 (N_3062,N_2885,N_2988);
or U3063 (N_3063,N_2898,N_2942);
nand U3064 (N_3064,N_2908,N_2918);
nor U3065 (N_3065,N_3030,N_3001);
and U3066 (N_3066,N_2964,N_2995);
and U3067 (N_3067,N_3011,N_2991);
nor U3068 (N_3068,N_3035,N_2881);
and U3069 (N_3069,N_3029,N_2891);
or U3070 (N_3070,N_2987,N_2893);
xnor U3071 (N_3071,N_2883,N_3020);
xor U3072 (N_3072,N_2961,N_3031);
nand U3073 (N_3073,N_3009,N_2910);
nor U3074 (N_3074,N_3037,N_2913);
xnor U3075 (N_3075,N_2973,N_2963);
and U3076 (N_3076,N_3013,N_3034);
nand U3077 (N_3077,N_3019,N_2965);
nor U3078 (N_3078,N_2902,N_3012);
xor U3079 (N_3079,N_2886,N_3015);
nor U3080 (N_3080,N_2882,N_3023);
or U3081 (N_3081,N_3017,N_2887);
and U3082 (N_3082,N_2978,N_2984);
xor U3083 (N_3083,N_2950,N_2957);
and U3084 (N_3084,N_2938,N_2979);
xnor U3085 (N_3085,N_2975,N_2944);
xnor U3086 (N_3086,N_2953,N_2907);
and U3087 (N_3087,N_2958,N_3008);
xnor U3088 (N_3088,N_2888,N_2976);
nor U3089 (N_3089,N_2931,N_2906);
or U3090 (N_3090,N_2922,N_2912);
or U3091 (N_3091,N_3018,N_2983);
and U3092 (N_3092,N_3039,N_3002);
nor U3093 (N_3093,N_2939,N_2992);
nor U3094 (N_3094,N_2974,N_3028);
and U3095 (N_3095,N_2977,N_3010);
nor U3096 (N_3096,N_2889,N_2982);
nor U3097 (N_3097,N_3025,N_2951);
xnor U3098 (N_3098,N_2932,N_2948);
xnor U3099 (N_3099,N_3021,N_2937);
nand U3100 (N_3100,N_2892,N_3005);
xnor U3101 (N_3101,N_2884,N_2926);
and U3102 (N_3102,N_2994,N_2999);
or U3103 (N_3103,N_2967,N_2924);
or U3104 (N_3104,N_2919,N_2955);
or U3105 (N_3105,N_3007,N_2904);
nor U3106 (N_3106,N_2896,N_2921);
and U3107 (N_3107,N_2996,N_2909);
nor U3108 (N_3108,N_2981,N_2972);
nand U3109 (N_3109,N_2900,N_3033);
nand U3110 (N_3110,N_2920,N_2917);
nand U3111 (N_3111,N_2941,N_2985);
and U3112 (N_3112,N_2933,N_2966);
nand U3113 (N_3113,N_3027,N_2927);
nand U3114 (N_3114,N_2949,N_3038);
nand U3115 (N_3115,N_2943,N_2890);
or U3116 (N_3116,N_2968,N_2980);
and U3117 (N_3117,N_2962,N_2945);
or U3118 (N_3118,N_2911,N_2914);
xnor U3119 (N_3119,N_2880,N_2894);
or U3120 (N_3120,N_3009,N_3039);
nor U3121 (N_3121,N_2941,N_2897);
and U3122 (N_3122,N_3022,N_2970);
nand U3123 (N_3123,N_2904,N_2958);
nor U3124 (N_3124,N_3001,N_3007);
nand U3125 (N_3125,N_2964,N_3028);
or U3126 (N_3126,N_2907,N_2962);
or U3127 (N_3127,N_2972,N_2975);
and U3128 (N_3128,N_2953,N_2914);
and U3129 (N_3129,N_2988,N_2965);
and U3130 (N_3130,N_2969,N_2994);
nor U3131 (N_3131,N_3037,N_3000);
xnor U3132 (N_3132,N_3012,N_2978);
nand U3133 (N_3133,N_2975,N_2942);
or U3134 (N_3134,N_2973,N_2923);
nor U3135 (N_3135,N_2890,N_2958);
and U3136 (N_3136,N_2969,N_2940);
or U3137 (N_3137,N_2997,N_2956);
nand U3138 (N_3138,N_2902,N_2882);
and U3139 (N_3139,N_2948,N_2954);
or U3140 (N_3140,N_2949,N_2956);
nand U3141 (N_3141,N_3016,N_2898);
nor U3142 (N_3142,N_3018,N_2880);
xnor U3143 (N_3143,N_2962,N_2934);
or U3144 (N_3144,N_2997,N_2961);
nor U3145 (N_3145,N_2979,N_3019);
and U3146 (N_3146,N_2929,N_2946);
or U3147 (N_3147,N_2973,N_2938);
and U3148 (N_3148,N_2948,N_2980);
and U3149 (N_3149,N_3036,N_2956);
and U3150 (N_3150,N_2948,N_2886);
nand U3151 (N_3151,N_2984,N_3029);
or U3152 (N_3152,N_2939,N_2901);
and U3153 (N_3153,N_3002,N_2892);
nor U3154 (N_3154,N_3010,N_3016);
nand U3155 (N_3155,N_2977,N_2939);
nand U3156 (N_3156,N_2951,N_2962);
nand U3157 (N_3157,N_2967,N_2906);
and U3158 (N_3158,N_2893,N_2968);
and U3159 (N_3159,N_2975,N_3023);
xor U3160 (N_3160,N_2908,N_3032);
nand U3161 (N_3161,N_2901,N_2998);
xor U3162 (N_3162,N_2912,N_2938);
and U3163 (N_3163,N_2981,N_2998);
or U3164 (N_3164,N_3005,N_2910);
xor U3165 (N_3165,N_2901,N_2897);
nor U3166 (N_3166,N_2915,N_2935);
or U3167 (N_3167,N_2901,N_2908);
nand U3168 (N_3168,N_2881,N_2927);
and U3169 (N_3169,N_3015,N_2972);
and U3170 (N_3170,N_2940,N_3017);
and U3171 (N_3171,N_2941,N_2986);
nor U3172 (N_3172,N_2950,N_3000);
and U3173 (N_3173,N_2946,N_2991);
or U3174 (N_3174,N_2915,N_2930);
nor U3175 (N_3175,N_2998,N_2951);
and U3176 (N_3176,N_2968,N_2882);
xnor U3177 (N_3177,N_3032,N_2937);
nor U3178 (N_3178,N_2997,N_2988);
nor U3179 (N_3179,N_3030,N_2937);
nand U3180 (N_3180,N_2985,N_2911);
nand U3181 (N_3181,N_2953,N_2946);
xnor U3182 (N_3182,N_2939,N_2955);
nand U3183 (N_3183,N_2990,N_2899);
and U3184 (N_3184,N_3014,N_3024);
nor U3185 (N_3185,N_3002,N_2891);
nand U3186 (N_3186,N_2890,N_2947);
xnor U3187 (N_3187,N_2884,N_2935);
and U3188 (N_3188,N_3009,N_2973);
xor U3189 (N_3189,N_2968,N_2944);
nand U3190 (N_3190,N_2881,N_3028);
and U3191 (N_3191,N_3004,N_3006);
xnor U3192 (N_3192,N_2972,N_2916);
and U3193 (N_3193,N_2959,N_2908);
nand U3194 (N_3194,N_2946,N_2963);
or U3195 (N_3195,N_2996,N_3002);
or U3196 (N_3196,N_2938,N_2900);
and U3197 (N_3197,N_2885,N_2933);
or U3198 (N_3198,N_2913,N_2967);
xor U3199 (N_3199,N_2959,N_2904);
nor U3200 (N_3200,N_3060,N_3094);
nor U3201 (N_3201,N_3180,N_3044);
nand U3202 (N_3202,N_3108,N_3156);
or U3203 (N_3203,N_3067,N_3051);
xnor U3204 (N_3204,N_3074,N_3148);
or U3205 (N_3205,N_3198,N_3158);
nand U3206 (N_3206,N_3053,N_3045);
xor U3207 (N_3207,N_3114,N_3185);
xnor U3208 (N_3208,N_3162,N_3055);
and U3209 (N_3209,N_3189,N_3079);
nand U3210 (N_3210,N_3059,N_3177);
nand U3211 (N_3211,N_3166,N_3154);
and U3212 (N_3212,N_3122,N_3139);
nand U3213 (N_3213,N_3197,N_3173);
and U3214 (N_3214,N_3179,N_3088);
nand U3215 (N_3215,N_3110,N_3111);
nand U3216 (N_3216,N_3047,N_3116);
nand U3217 (N_3217,N_3090,N_3068);
or U3218 (N_3218,N_3048,N_3123);
and U3219 (N_3219,N_3167,N_3147);
nor U3220 (N_3220,N_3109,N_3112);
nor U3221 (N_3221,N_3155,N_3153);
xnor U3222 (N_3222,N_3195,N_3042);
nor U3223 (N_3223,N_3191,N_3190);
nand U3224 (N_3224,N_3165,N_3152);
nand U3225 (N_3225,N_3159,N_3086);
nor U3226 (N_3226,N_3193,N_3138);
nand U3227 (N_3227,N_3163,N_3084);
xnor U3228 (N_3228,N_3085,N_3157);
and U3229 (N_3229,N_3066,N_3121);
xor U3230 (N_3230,N_3174,N_3171);
and U3231 (N_3231,N_3081,N_3199);
or U3232 (N_3232,N_3149,N_3056);
nand U3233 (N_3233,N_3102,N_3129);
and U3234 (N_3234,N_3145,N_3130);
or U3235 (N_3235,N_3098,N_3097);
xnor U3236 (N_3236,N_3101,N_3140);
nor U3237 (N_3237,N_3192,N_3172);
or U3238 (N_3238,N_3141,N_3120);
xor U3239 (N_3239,N_3196,N_3040);
nand U3240 (N_3240,N_3063,N_3099);
nand U3241 (N_3241,N_3057,N_3076);
nor U3242 (N_3242,N_3150,N_3164);
and U3243 (N_3243,N_3126,N_3103);
nand U3244 (N_3244,N_3151,N_3096);
and U3245 (N_3245,N_3069,N_3064);
nor U3246 (N_3246,N_3071,N_3049);
xnor U3247 (N_3247,N_3107,N_3161);
or U3248 (N_3248,N_3117,N_3089);
or U3249 (N_3249,N_3182,N_3183);
nand U3250 (N_3250,N_3077,N_3124);
nand U3251 (N_3251,N_3115,N_3087);
nand U3252 (N_3252,N_3061,N_3132);
or U3253 (N_3253,N_3128,N_3058);
nor U3254 (N_3254,N_3186,N_3136);
and U3255 (N_3255,N_3176,N_3082);
and U3256 (N_3256,N_3072,N_3160);
or U3257 (N_3257,N_3083,N_3118);
or U3258 (N_3258,N_3070,N_3178);
nor U3259 (N_3259,N_3043,N_3135);
nand U3260 (N_3260,N_3146,N_3142);
nor U3261 (N_3261,N_3187,N_3075);
nand U3262 (N_3262,N_3170,N_3050);
nand U3263 (N_3263,N_3052,N_3137);
xnor U3264 (N_3264,N_3080,N_3092);
and U3265 (N_3265,N_3133,N_3046);
or U3266 (N_3266,N_3188,N_3144);
and U3267 (N_3267,N_3131,N_3134);
nor U3268 (N_3268,N_3073,N_3181);
nor U3269 (N_3269,N_3106,N_3105);
nand U3270 (N_3270,N_3100,N_3062);
or U3271 (N_3271,N_3175,N_3168);
nand U3272 (N_3272,N_3127,N_3194);
or U3273 (N_3273,N_3184,N_3125);
or U3274 (N_3274,N_3041,N_3113);
or U3275 (N_3275,N_3065,N_3093);
or U3276 (N_3276,N_3104,N_3119);
nand U3277 (N_3277,N_3095,N_3078);
nor U3278 (N_3278,N_3091,N_3169);
or U3279 (N_3279,N_3143,N_3054);
and U3280 (N_3280,N_3041,N_3180);
or U3281 (N_3281,N_3185,N_3097);
or U3282 (N_3282,N_3191,N_3091);
or U3283 (N_3283,N_3197,N_3121);
xor U3284 (N_3284,N_3071,N_3194);
nand U3285 (N_3285,N_3121,N_3078);
nand U3286 (N_3286,N_3112,N_3183);
xnor U3287 (N_3287,N_3057,N_3050);
nand U3288 (N_3288,N_3180,N_3127);
nand U3289 (N_3289,N_3139,N_3130);
nand U3290 (N_3290,N_3062,N_3175);
and U3291 (N_3291,N_3053,N_3100);
or U3292 (N_3292,N_3074,N_3144);
nand U3293 (N_3293,N_3075,N_3136);
and U3294 (N_3294,N_3043,N_3095);
nor U3295 (N_3295,N_3069,N_3104);
nor U3296 (N_3296,N_3055,N_3149);
or U3297 (N_3297,N_3180,N_3099);
xor U3298 (N_3298,N_3128,N_3074);
xnor U3299 (N_3299,N_3100,N_3103);
nor U3300 (N_3300,N_3068,N_3098);
or U3301 (N_3301,N_3154,N_3099);
nand U3302 (N_3302,N_3095,N_3042);
xor U3303 (N_3303,N_3157,N_3140);
or U3304 (N_3304,N_3142,N_3058);
and U3305 (N_3305,N_3126,N_3188);
nand U3306 (N_3306,N_3174,N_3185);
nand U3307 (N_3307,N_3133,N_3107);
or U3308 (N_3308,N_3099,N_3055);
nand U3309 (N_3309,N_3124,N_3103);
xnor U3310 (N_3310,N_3155,N_3137);
nand U3311 (N_3311,N_3042,N_3193);
nor U3312 (N_3312,N_3121,N_3041);
nand U3313 (N_3313,N_3152,N_3181);
or U3314 (N_3314,N_3174,N_3048);
and U3315 (N_3315,N_3066,N_3181);
or U3316 (N_3316,N_3134,N_3099);
and U3317 (N_3317,N_3170,N_3072);
and U3318 (N_3318,N_3185,N_3179);
nor U3319 (N_3319,N_3075,N_3061);
nand U3320 (N_3320,N_3181,N_3199);
and U3321 (N_3321,N_3133,N_3116);
or U3322 (N_3322,N_3169,N_3122);
or U3323 (N_3323,N_3112,N_3093);
nor U3324 (N_3324,N_3116,N_3163);
nand U3325 (N_3325,N_3166,N_3192);
or U3326 (N_3326,N_3124,N_3191);
or U3327 (N_3327,N_3063,N_3115);
or U3328 (N_3328,N_3079,N_3087);
and U3329 (N_3329,N_3193,N_3199);
and U3330 (N_3330,N_3131,N_3193);
nor U3331 (N_3331,N_3131,N_3075);
nor U3332 (N_3332,N_3056,N_3060);
and U3333 (N_3333,N_3143,N_3074);
nor U3334 (N_3334,N_3057,N_3075);
and U3335 (N_3335,N_3122,N_3179);
xor U3336 (N_3336,N_3060,N_3148);
xor U3337 (N_3337,N_3062,N_3069);
nor U3338 (N_3338,N_3184,N_3147);
or U3339 (N_3339,N_3134,N_3142);
xor U3340 (N_3340,N_3196,N_3047);
xnor U3341 (N_3341,N_3058,N_3107);
nor U3342 (N_3342,N_3191,N_3149);
or U3343 (N_3343,N_3180,N_3101);
nand U3344 (N_3344,N_3059,N_3118);
xor U3345 (N_3345,N_3183,N_3095);
and U3346 (N_3346,N_3113,N_3177);
xor U3347 (N_3347,N_3073,N_3108);
nor U3348 (N_3348,N_3184,N_3199);
xor U3349 (N_3349,N_3091,N_3157);
nor U3350 (N_3350,N_3174,N_3085);
xor U3351 (N_3351,N_3149,N_3045);
xor U3352 (N_3352,N_3070,N_3119);
or U3353 (N_3353,N_3123,N_3089);
and U3354 (N_3354,N_3065,N_3155);
and U3355 (N_3355,N_3134,N_3080);
nor U3356 (N_3356,N_3047,N_3084);
or U3357 (N_3357,N_3098,N_3045);
nand U3358 (N_3358,N_3197,N_3109);
and U3359 (N_3359,N_3144,N_3071);
and U3360 (N_3360,N_3204,N_3302);
or U3361 (N_3361,N_3220,N_3286);
xnor U3362 (N_3362,N_3303,N_3267);
or U3363 (N_3363,N_3277,N_3338);
and U3364 (N_3364,N_3297,N_3240);
or U3365 (N_3365,N_3254,N_3263);
xnor U3366 (N_3366,N_3351,N_3335);
xnor U3367 (N_3367,N_3246,N_3315);
and U3368 (N_3368,N_3317,N_3299);
xnor U3369 (N_3369,N_3225,N_3260);
xnor U3370 (N_3370,N_3331,N_3336);
and U3371 (N_3371,N_3208,N_3308);
nand U3372 (N_3372,N_3262,N_3249);
and U3373 (N_3373,N_3236,N_3322);
or U3374 (N_3374,N_3233,N_3268);
and U3375 (N_3375,N_3227,N_3347);
or U3376 (N_3376,N_3304,N_3242);
xor U3377 (N_3377,N_3241,N_3329);
nor U3378 (N_3378,N_3340,N_3327);
nand U3379 (N_3379,N_3265,N_3206);
and U3380 (N_3380,N_3276,N_3324);
or U3381 (N_3381,N_3257,N_3200);
and U3382 (N_3382,N_3235,N_3224);
nor U3383 (N_3383,N_3339,N_3203);
nand U3384 (N_3384,N_3313,N_3239);
nor U3385 (N_3385,N_3215,N_3216);
and U3386 (N_3386,N_3231,N_3284);
nand U3387 (N_3387,N_3358,N_3345);
xnor U3388 (N_3388,N_3346,N_3258);
xnor U3389 (N_3389,N_3274,N_3323);
nand U3390 (N_3390,N_3292,N_3234);
or U3391 (N_3391,N_3333,N_3226);
nand U3392 (N_3392,N_3328,N_3282);
nand U3393 (N_3393,N_3355,N_3210);
nand U3394 (N_3394,N_3205,N_3269);
nor U3395 (N_3395,N_3311,N_3237);
or U3396 (N_3396,N_3309,N_3341);
nor U3397 (N_3397,N_3261,N_3252);
or U3398 (N_3398,N_3306,N_3279);
or U3399 (N_3399,N_3348,N_3207);
xor U3400 (N_3400,N_3310,N_3273);
xor U3401 (N_3401,N_3217,N_3283);
nand U3402 (N_3402,N_3320,N_3352);
nand U3403 (N_3403,N_3314,N_3305);
or U3404 (N_3404,N_3287,N_3218);
nand U3405 (N_3405,N_3298,N_3238);
nor U3406 (N_3406,N_3290,N_3295);
or U3407 (N_3407,N_3278,N_3357);
xor U3408 (N_3408,N_3281,N_3250);
nor U3409 (N_3409,N_3244,N_3266);
nor U3410 (N_3410,N_3321,N_3243);
nand U3411 (N_3411,N_3296,N_3256);
or U3412 (N_3412,N_3221,N_3280);
nand U3413 (N_3413,N_3228,N_3300);
or U3414 (N_3414,N_3293,N_3350);
xnor U3415 (N_3415,N_3201,N_3223);
xor U3416 (N_3416,N_3354,N_3209);
nor U3417 (N_3417,N_3285,N_3222);
or U3418 (N_3418,N_3343,N_3270);
or U3419 (N_3419,N_3289,N_3316);
xor U3420 (N_3420,N_3326,N_3271);
nor U3421 (N_3421,N_3214,N_3275);
nand U3422 (N_3422,N_3248,N_3330);
or U3423 (N_3423,N_3294,N_3245);
xor U3424 (N_3424,N_3251,N_3312);
xnor U3425 (N_3425,N_3213,N_3353);
nor U3426 (N_3426,N_3301,N_3337);
or U3427 (N_3427,N_3359,N_3229);
nand U3428 (N_3428,N_3344,N_3356);
nand U3429 (N_3429,N_3232,N_3325);
or U3430 (N_3430,N_3307,N_3253);
xor U3431 (N_3431,N_3318,N_3288);
and U3432 (N_3432,N_3255,N_3230);
and U3433 (N_3433,N_3349,N_3342);
xor U3434 (N_3434,N_3334,N_3264);
xor U3435 (N_3435,N_3247,N_3211);
nor U3436 (N_3436,N_3291,N_3319);
and U3437 (N_3437,N_3219,N_3202);
and U3438 (N_3438,N_3272,N_3212);
nand U3439 (N_3439,N_3259,N_3332);
xnor U3440 (N_3440,N_3207,N_3218);
nor U3441 (N_3441,N_3210,N_3230);
nor U3442 (N_3442,N_3241,N_3276);
or U3443 (N_3443,N_3330,N_3275);
nor U3444 (N_3444,N_3311,N_3286);
nor U3445 (N_3445,N_3282,N_3290);
and U3446 (N_3446,N_3216,N_3312);
xor U3447 (N_3447,N_3289,N_3267);
xnor U3448 (N_3448,N_3292,N_3273);
xnor U3449 (N_3449,N_3269,N_3317);
nor U3450 (N_3450,N_3273,N_3290);
or U3451 (N_3451,N_3225,N_3273);
or U3452 (N_3452,N_3232,N_3251);
nand U3453 (N_3453,N_3304,N_3213);
xnor U3454 (N_3454,N_3203,N_3223);
or U3455 (N_3455,N_3340,N_3215);
nor U3456 (N_3456,N_3200,N_3327);
and U3457 (N_3457,N_3304,N_3350);
and U3458 (N_3458,N_3292,N_3263);
or U3459 (N_3459,N_3334,N_3332);
xnor U3460 (N_3460,N_3336,N_3323);
nand U3461 (N_3461,N_3344,N_3275);
nand U3462 (N_3462,N_3208,N_3304);
xor U3463 (N_3463,N_3254,N_3238);
and U3464 (N_3464,N_3285,N_3270);
nor U3465 (N_3465,N_3223,N_3249);
and U3466 (N_3466,N_3230,N_3267);
or U3467 (N_3467,N_3305,N_3321);
nand U3468 (N_3468,N_3343,N_3206);
or U3469 (N_3469,N_3286,N_3235);
nand U3470 (N_3470,N_3280,N_3347);
or U3471 (N_3471,N_3258,N_3287);
and U3472 (N_3472,N_3295,N_3318);
and U3473 (N_3473,N_3299,N_3234);
or U3474 (N_3474,N_3203,N_3238);
xor U3475 (N_3475,N_3277,N_3335);
nand U3476 (N_3476,N_3207,N_3212);
and U3477 (N_3477,N_3321,N_3358);
and U3478 (N_3478,N_3350,N_3207);
nand U3479 (N_3479,N_3282,N_3331);
nor U3480 (N_3480,N_3274,N_3269);
and U3481 (N_3481,N_3259,N_3336);
or U3482 (N_3482,N_3329,N_3214);
and U3483 (N_3483,N_3287,N_3290);
nor U3484 (N_3484,N_3314,N_3217);
nor U3485 (N_3485,N_3332,N_3225);
or U3486 (N_3486,N_3335,N_3320);
nand U3487 (N_3487,N_3226,N_3319);
nand U3488 (N_3488,N_3219,N_3247);
or U3489 (N_3489,N_3259,N_3258);
nor U3490 (N_3490,N_3253,N_3306);
or U3491 (N_3491,N_3332,N_3287);
and U3492 (N_3492,N_3278,N_3294);
xor U3493 (N_3493,N_3329,N_3358);
and U3494 (N_3494,N_3226,N_3281);
xnor U3495 (N_3495,N_3343,N_3337);
xor U3496 (N_3496,N_3210,N_3253);
or U3497 (N_3497,N_3230,N_3319);
xnor U3498 (N_3498,N_3258,N_3342);
nand U3499 (N_3499,N_3250,N_3253);
nor U3500 (N_3500,N_3290,N_3247);
or U3501 (N_3501,N_3244,N_3262);
nand U3502 (N_3502,N_3314,N_3229);
or U3503 (N_3503,N_3334,N_3239);
or U3504 (N_3504,N_3292,N_3304);
nand U3505 (N_3505,N_3348,N_3329);
xnor U3506 (N_3506,N_3214,N_3322);
nand U3507 (N_3507,N_3316,N_3247);
or U3508 (N_3508,N_3241,N_3330);
nor U3509 (N_3509,N_3220,N_3359);
xnor U3510 (N_3510,N_3346,N_3250);
or U3511 (N_3511,N_3200,N_3273);
and U3512 (N_3512,N_3325,N_3239);
and U3513 (N_3513,N_3238,N_3207);
nand U3514 (N_3514,N_3333,N_3260);
or U3515 (N_3515,N_3223,N_3318);
nand U3516 (N_3516,N_3265,N_3218);
or U3517 (N_3517,N_3298,N_3227);
xnor U3518 (N_3518,N_3313,N_3231);
nor U3519 (N_3519,N_3301,N_3341);
nor U3520 (N_3520,N_3366,N_3460);
and U3521 (N_3521,N_3453,N_3484);
or U3522 (N_3522,N_3426,N_3401);
xnor U3523 (N_3523,N_3385,N_3428);
nand U3524 (N_3524,N_3506,N_3384);
nor U3525 (N_3525,N_3382,N_3371);
xor U3526 (N_3526,N_3509,N_3363);
nor U3527 (N_3527,N_3431,N_3501);
or U3528 (N_3528,N_3397,N_3422);
xnor U3529 (N_3529,N_3380,N_3416);
and U3530 (N_3530,N_3446,N_3452);
nor U3531 (N_3531,N_3441,N_3487);
and U3532 (N_3532,N_3394,N_3498);
xor U3533 (N_3533,N_3507,N_3482);
and U3534 (N_3534,N_3468,N_3456);
and U3535 (N_3535,N_3517,N_3479);
or U3536 (N_3536,N_3373,N_3407);
and U3537 (N_3537,N_3418,N_3383);
nor U3538 (N_3538,N_3424,N_3374);
xnor U3539 (N_3539,N_3449,N_3387);
nor U3540 (N_3540,N_3378,N_3483);
or U3541 (N_3541,N_3417,N_3425);
and U3542 (N_3542,N_3473,N_3457);
nor U3543 (N_3543,N_3388,N_3377);
nor U3544 (N_3544,N_3386,N_3365);
xnor U3545 (N_3545,N_3376,N_3361);
nand U3546 (N_3546,N_3475,N_3375);
nand U3547 (N_3547,N_3519,N_3467);
and U3548 (N_3548,N_3493,N_3458);
or U3549 (N_3549,N_3502,N_3423);
and U3550 (N_3550,N_3360,N_3412);
nor U3551 (N_3551,N_3490,N_3372);
nor U3552 (N_3552,N_3445,N_3516);
xor U3553 (N_3553,N_3430,N_3393);
nand U3554 (N_3554,N_3362,N_3433);
nor U3555 (N_3555,N_3368,N_3503);
nor U3556 (N_3556,N_3451,N_3450);
nor U3557 (N_3557,N_3515,N_3472);
or U3558 (N_3558,N_3494,N_3391);
or U3559 (N_3559,N_3398,N_3455);
nor U3560 (N_3560,N_3403,N_3404);
or U3561 (N_3561,N_3512,N_3415);
nor U3562 (N_3562,N_3478,N_3514);
xor U3563 (N_3563,N_3486,N_3496);
or U3564 (N_3564,N_3461,N_3471);
or U3565 (N_3565,N_3406,N_3419);
nand U3566 (N_3566,N_3447,N_3409);
and U3567 (N_3567,N_3370,N_3476);
xnor U3568 (N_3568,N_3392,N_3504);
or U3569 (N_3569,N_3414,N_3491);
and U3570 (N_3570,N_3389,N_3480);
xnor U3571 (N_3571,N_3367,N_3364);
and U3572 (N_3572,N_3443,N_3465);
or U3573 (N_3573,N_3489,N_3405);
nand U3574 (N_3574,N_3505,N_3474);
nand U3575 (N_3575,N_3454,N_3379);
nand U3576 (N_3576,N_3518,N_3436);
nor U3577 (N_3577,N_3495,N_3485);
nor U3578 (N_3578,N_3395,N_3466);
xor U3579 (N_3579,N_3459,N_3508);
nand U3580 (N_3580,N_3440,N_3477);
nand U3581 (N_3581,N_3488,N_3463);
or U3582 (N_3582,N_3481,N_3437);
nor U3583 (N_3583,N_3381,N_3402);
xnor U3584 (N_3584,N_3511,N_3497);
or U3585 (N_3585,N_3411,N_3510);
nand U3586 (N_3586,N_3399,N_3420);
or U3587 (N_3587,N_3369,N_3439);
xnor U3588 (N_3588,N_3499,N_3421);
or U3589 (N_3589,N_3408,N_3432);
nand U3590 (N_3590,N_3435,N_3427);
xnor U3591 (N_3591,N_3492,N_3444);
and U3592 (N_3592,N_3470,N_3429);
nor U3593 (N_3593,N_3462,N_3396);
nand U3594 (N_3594,N_3469,N_3400);
xnor U3595 (N_3595,N_3448,N_3464);
and U3596 (N_3596,N_3438,N_3390);
xnor U3597 (N_3597,N_3442,N_3410);
or U3598 (N_3598,N_3413,N_3513);
xor U3599 (N_3599,N_3434,N_3500);
and U3600 (N_3600,N_3408,N_3388);
and U3601 (N_3601,N_3495,N_3383);
or U3602 (N_3602,N_3427,N_3476);
nor U3603 (N_3603,N_3395,N_3392);
or U3604 (N_3604,N_3432,N_3507);
xor U3605 (N_3605,N_3377,N_3471);
xor U3606 (N_3606,N_3416,N_3371);
and U3607 (N_3607,N_3408,N_3461);
or U3608 (N_3608,N_3435,N_3499);
or U3609 (N_3609,N_3460,N_3403);
or U3610 (N_3610,N_3422,N_3511);
and U3611 (N_3611,N_3430,N_3482);
nand U3612 (N_3612,N_3475,N_3492);
or U3613 (N_3613,N_3457,N_3481);
or U3614 (N_3614,N_3380,N_3417);
or U3615 (N_3615,N_3431,N_3371);
and U3616 (N_3616,N_3360,N_3463);
and U3617 (N_3617,N_3392,N_3480);
xor U3618 (N_3618,N_3442,N_3515);
nor U3619 (N_3619,N_3449,N_3412);
and U3620 (N_3620,N_3488,N_3408);
nand U3621 (N_3621,N_3483,N_3361);
and U3622 (N_3622,N_3448,N_3460);
nor U3623 (N_3623,N_3427,N_3407);
xor U3624 (N_3624,N_3421,N_3445);
xnor U3625 (N_3625,N_3442,N_3516);
xnor U3626 (N_3626,N_3503,N_3391);
and U3627 (N_3627,N_3506,N_3388);
xor U3628 (N_3628,N_3498,N_3518);
and U3629 (N_3629,N_3480,N_3396);
xor U3630 (N_3630,N_3439,N_3385);
nand U3631 (N_3631,N_3500,N_3501);
or U3632 (N_3632,N_3397,N_3374);
or U3633 (N_3633,N_3481,N_3409);
nand U3634 (N_3634,N_3488,N_3395);
nand U3635 (N_3635,N_3430,N_3493);
or U3636 (N_3636,N_3503,N_3467);
xnor U3637 (N_3637,N_3518,N_3409);
nand U3638 (N_3638,N_3492,N_3453);
and U3639 (N_3639,N_3453,N_3511);
or U3640 (N_3640,N_3385,N_3384);
nand U3641 (N_3641,N_3387,N_3494);
xor U3642 (N_3642,N_3431,N_3363);
xor U3643 (N_3643,N_3420,N_3391);
nand U3644 (N_3644,N_3375,N_3518);
xor U3645 (N_3645,N_3495,N_3417);
xnor U3646 (N_3646,N_3504,N_3484);
and U3647 (N_3647,N_3499,N_3412);
xnor U3648 (N_3648,N_3472,N_3489);
and U3649 (N_3649,N_3497,N_3402);
or U3650 (N_3650,N_3400,N_3418);
or U3651 (N_3651,N_3498,N_3423);
nand U3652 (N_3652,N_3361,N_3487);
or U3653 (N_3653,N_3465,N_3479);
or U3654 (N_3654,N_3475,N_3514);
nand U3655 (N_3655,N_3409,N_3384);
xor U3656 (N_3656,N_3469,N_3489);
nor U3657 (N_3657,N_3365,N_3417);
or U3658 (N_3658,N_3393,N_3363);
and U3659 (N_3659,N_3403,N_3484);
xnor U3660 (N_3660,N_3481,N_3375);
or U3661 (N_3661,N_3400,N_3454);
nor U3662 (N_3662,N_3424,N_3373);
and U3663 (N_3663,N_3479,N_3511);
xnor U3664 (N_3664,N_3474,N_3387);
nor U3665 (N_3665,N_3420,N_3372);
nand U3666 (N_3666,N_3488,N_3492);
or U3667 (N_3667,N_3435,N_3360);
and U3668 (N_3668,N_3493,N_3365);
xnor U3669 (N_3669,N_3483,N_3379);
or U3670 (N_3670,N_3515,N_3454);
or U3671 (N_3671,N_3424,N_3496);
and U3672 (N_3672,N_3513,N_3478);
nor U3673 (N_3673,N_3509,N_3469);
and U3674 (N_3674,N_3470,N_3373);
nand U3675 (N_3675,N_3454,N_3394);
and U3676 (N_3676,N_3375,N_3424);
xnor U3677 (N_3677,N_3492,N_3365);
nor U3678 (N_3678,N_3364,N_3368);
xnor U3679 (N_3679,N_3490,N_3448);
or U3680 (N_3680,N_3537,N_3558);
and U3681 (N_3681,N_3671,N_3599);
or U3682 (N_3682,N_3568,N_3592);
xnor U3683 (N_3683,N_3634,N_3647);
nand U3684 (N_3684,N_3641,N_3541);
and U3685 (N_3685,N_3528,N_3672);
nor U3686 (N_3686,N_3535,N_3608);
nor U3687 (N_3687,N_3676,N_3637);
nand U3688 (N_3688,N_3563,N_3602);
nor U3689 (N_3689,N_3649,N_3555);
xnor U3690 (N_3690,N_3566,N_3668);
nor U3691 (N_3691,N_3648,N_3674);
and U3692 (N_3692,N_3533,N_3589);
nor U3693 (N_3693,N_3636,N_3594);
nor U3694 (N_3694,N_3605,N_3584);
nor U3695 (N_3695,N_3585,N_3583);
xor U3696 (N_3696,N_3570,N_3652);
and U3697 (N_3697,N_3580,N_3653);
or U3698 (N_3698,N_3581,N_3679);
and U3699 (N_3699,N_3593,N_3530);
nor U3700 (N_3700,N_3678,N_3625);
xnor U3701 (N_3701,N_3538,N_3643);
or U3702 (N_3702,N_3632,N_3574);
or U3703 (N_3703,N_3656,N_3567);
nand U3704 (N_3704,N_3638,N_3630);
nor U3705 (N_3705,N_3640,N_3655);
xnor U3706 (N_3706,N_3559,N_3600);
or U3707 (N_3707,N_3669,N_3557);
nand U3708 (N_3708,N_3662,N_3522);
or U3709 (N_3709,N_3610,N_3635);
nor U3710 (N_3710,N_3551,N_3616);
and U3711 (N_3711,N_3546,N_3601);
xnor U3712 (N_3712,N_3545,N_3663);
nand U3713 (N_3713,N_3572,N_3520);
and U3714 (N_3714,N_3664,N_3523);
nor U3715 (N_3715,N_3590,N_3573);
or U3716 (N_3716,N_3524,N_3606);
xnor U3717 (N_3717,N_3654,N_3526);
nor U3718 (N_3718,N_3677,N_3639);
xnor U3719 (N_3719,N_3521,N_3661);
or U3720 (N_3720,N_3614,N_3666);
and U3721 (N_3721,N_3673,N_3650);
nand U3722 (N_3722,N_3595,N_3613);
xor U3723 (N_3723,N_3531,N_3534);
nand U3724 (N_3724,N_3633,N_3626);
nor U3725 (N_3725,N_3611,N_3548);
xor U3726 (N_3726,N_3642,N_3619);
or U3727 (N_3727,N_3586,N_3644);
and U3728 (N_3728,N_3556,N_3620);
nand U3729 (N_3729,N_3598,N_3646);
xnor U3730 (N_3730,N_3542,N_3587);
and U3731 (N_3731,N_3547,N_3627);
nor U3732 (N_3732,N_3554,N_3561);
and U3733 (N_3733,N_3575,N_3645);
or U3734 (N_3734,N_3604,N_3527);
and U3735 (N_3735,N_3657,N_3628);
and U3736 (N_3736,N_3549,N_3670);
nor U3737 (N_3737,N_3536,N_3569);
or U3738 (N_3738,N_3579,N_3597);
or U3739 (N_3739,N_3631,N_3582);
or U3740 (N_3740,N_3615,N_3564);
nand U3741 (N_3741,N_3576,N_3571);
and U3742 (N_3742,N_3603,N_3529);
xor U3743 (N_3743,N_3532,N_3591);
nand U3744 (N_3744,N_3596,N_3623);
or U3745 (N_3745,N_3659,N_3560);
or U3746 (N_3746,N_3612,N_3651);
nor U3747 (N_3747,N_3552,N_3544);
or U3748 (N_3748,N_3675,N_3588);
and U3749 (N_3749,N_3622,N_3624);
nand U3750 (N_3750,N_3550,N_3609);
nand U3751 (N_3751,N_3578,N_3667);
nand U3752 (N_3752,N_3617,N_3618);
or U3753 (N_3753,N_3621,N_3553);
and U3754 (N_3754,N_3565,N_3658);
xor U3755 (N_3755,N_3665,N_3562);
or U3756 (N_3756,N_3577,N_3539);
or U3757 (N_3757,N_3607,N_3543);
nor U3758 (N_3758,N_3629,N_3540);
nand U3759 (N_3759,N_3660,N_3525);
xor U3760 (N_3760,N_3669,N_3603);
xnor U3761 (N_3761,N_3668,N_3606);
nor U3762 (N_3762,N_3591,N_3561);
and U3763 (N_3763,N_3574,N_3588);
nand U3764 (N_3764,N_3591,N_3623);
and U3765 (N_3765,N_3585,N_3604);
and U3766 (N_3766,N_3598,N_3557);
or U3767 (N_3767,N_3536,N_3594);
nand U3768 (N_3768,N_3585,N_3580);
nand U3769 (N_3769,N_3520,N_3575);
or U3770 (N_3770,N_3643,N_3526);
nand U3771 (N_3771,N_3672,N_3602);
and U3772 (N_3772,N_3639,N_3573);
xor U3773 (N_3773,N_3592,N_3560);
nand U3774 (N_3774,N_3607,N_3656);
nor U3775 (N_3775,N_3544,N_3614);
xor U3776 (N_3776,N_3655,N_3650);
or U3777 (N_3777,N_3591,N_3530);
nor U3778 (N_3778,N_3593,N_3576);
or U3779 (N_3779,N_3544,N_3538);
and U3780 (N_3780,N_3581,N_3659);
and U3781 (N_3781,N_3644,N_3598);
nand U3782 (N_3782,N_3617,N_3534);
or U3783 (N_3783,N_3610,N_3546);
and U3784 (N_3784,N_3655,N_3665);
nand U3785 (N_3785,N_3615,N_3619);
nor U3786 (N_3786,N_3592,N_3674);
nand U3787 (N_3787,N_3630,N_3566);
xnor U3788 (N_3788,N_3557,N_3533);
or U3789 (N_3789,N_3657,N_3642);
or U3790 (N_3790,N_3676,N_3674);
nor U3791 (N_3791,N_3537,N_3611);
xor U3792 (N_3792,N_3645,N_3571);
nor U3793 (N_3793,N_3645,N_3530);
or U3794 (N_3794,N_3590,N_3540);
xnor U3795 (N_3795,N_3632,N_3525);
or U3796 (N_3796,N_3634,N_3672);
or U3797 (N_3797,N_3613,N_3563);
nor U3798 (N_3798,N_3651,N_3630);
xnor U3799 (N_3799,N_3611,N_3662);
xor U3800 (N_3800,N_3667,N_3634);
or U3801 (N_3801,N_3641,N_3664);
or U3802 (N_3802,N_3523,N_3520);
xnor U3803 (N_3803,N_3674,N_3568);
nor U3804 (N_3804,N_3532,N_3540);
xor U3805 (N_3805,N_3642,N_3589);
xor U3806 (N_3806,N_3679,N_3583);
xor U3807 (N_3807,N_3609,N_3613);
nand U3808 (N_3808,N_3660,N_3528);
and U3809 (N_3809,N_3568,N_3679);
xor U3810 (N_3810,N_3637,N_3638);
nand U3811 (N_3811,N_3640,N_3630);
nor U3812 (N_3812,N_3544,N_3533);
xor U3813 (N_3813,N_3550,N_3597);
nor U3814 (N_3814,N_3583,N_3591);
nor U3815 (N_3815,N_3637,N_3644);
nand U3816 (N_3816,N_3558,N_3588);
nand U3817 (N_3817,N_3580,N_3613);
nand U3818 (N_3818,N_3651,N_3602);
and U3819 (N_3819,N_3539,N_3559);
xor U3820 (N_3820,N_3545,N_3559);
xnor U3821 (N_3821,N_3669,N_3590);
and U3822 (N_3822,N_3559,N_3640);
nand U3823 (N_3823,N_3661,N_3655);
nand U3824 (N_3824,N_3657,N_3609);
nor U3825 (N_3825,N_3586,N_3528);
nand U3826 (N_3826,N_3679,N_3521);
or U3827 (N_3827,N_3540,N_3543);
and U3828 (N_3828,N_3541,N_3606);
nand U3829 (N_3829,N_3678,N_3568);
nand U3830 (N_3830,N_3574,N_3665);
nand U3831 (N_3831,N_3559,N_3583);
or U3832 (N_3832,N_3656,N_3634);
or U3833 (N_3833,N_3650,N_3647);
nor U3834 (N_3834,N_3535,N_3651);
or U3835 (N_3835,N_3543,N_3655);
and U3836 (N_3836,N_3656,N_3653);
and U3837 (N_3837,N_3624,N_3564);
or U3838 (N_3838,N_3544,N_3547);
nor U3839 (N_3839,N_3621,N_3525);
nor U3840 (N_3840,N_3695,N_3777);
and U3841 (N_3841,N_3802,N_3771);
xnor U3842 (N_3842,N_3758,N_3747);
nand U3843 (N_3843,N_3746,N_3733);
nor U3844 (N_3844,N_3828,N_3725);
and U3845 (N_3845,N_3702,N_3682);
nor U3846 (N_3846,N_3683,N_3740);
nand U3847 (N_3847,N_3691,N_3750);
xor U3848 (N_3848,N_3693,N_3749);
xor U3849 (N_3849,N_3811,N_3738);
xor U3850 (N_3850,N_3745,N_3761);
nor U3851 (N_3851,N_3796,N_3769);
nor U3852 (N_3852,N_3705,N_3760);
or U3853 (N_3853,N_3770,N_3786);
or U3854 (N_3854,N_3696,N_3717);
or U3855 (N_3855,N_3780,N_3719);
nor U3856 (N_3856,N_3751,N_3793);
and U3857 (N_3857,N_3783,N_3795);
or U3858 (N_3858,N_3806,N_3797);
or U3859 (N_3859,N_3823,N_3778);
or U3860 (N_3860,N_3812,N_3831);
nor U3861 (N_3861,N_3768,N_3779);
nor U3862 (N_3862,N_3726,N_3834);
nor U3863 (N_3863,N_3788,N_3699);
or U3864 (N_3864,N_3814,N_3785);
nor U3865 (N_3865,N_3731,N_3718);
and U3866 (N_3866,N_3715,N_3694);
nand U3867 (N_3867,N_3689,N_3722);
or U3868 (N_3868,N_3775,N_3791);
and U3869 (N_3869,N_3784,N_3728);
and U3870 (N_3870,N_3735,N_3794);
or U3871 (N_3871,N_3776,N_3743);
nand U3872 (N_3872,N_3692,N_3804);
and U3873 (N_3873,N_3686,N_3707);
nand U3874 (N_3874,N_3822,N_3716);
xor U3875 (N_3875,N_3690,N_3836);
nand U3876 (N_3876,N_3826,N_3720);
and U3877 (N_3877,N_3782,N_3799);
nand U3878 (N_3878,N_3781,N_3727);
nor U3879 (N_3879,N_3704,N_3741);
nor U3880 (N_3880,N_3837,N_3698);
xnor U3881 (N_3881,N_3713,N_3734);
or U3882 (N_3882,N_3766,N_3681);
xnor U3883 (N_3883,N_3838,N_3832);
nand U3884 (N_3884,N_3712,N_3813);
and U3885 (N_3885,N_3801,N_3808);
nor U3886 (N_3886,N_3816,N_3772);
and U3887 (N_3887,N_3774,N_3724);
and U3888 (N_3888,N_3787,N_3697);
xor U3889 (N_3889,N_3764,N_3798);
or U3890 (N_3890,N_3737,N_3752);
nand U3891 (N_3891,N_3739,N_3824);
nor U3892 (N_3892,N_3807,N_3762);
and U3893 (N_3893,N_3835,N_3789);
nand U3894 (N_3894,N_3730,N_3790);
and U3895 (N_3895,N_3754,N_3708);
xnor U3896 (N_3896,N_3815,N_3688);
nand U3897 (N_3897,N_3744,N_3714);
or U3898 (N_3898,N_3703,N_3765);
nor U3899 (N_3899,N_3792,N_3710);
xnor U3900 (N_3900,N_3700,N_3800);
and U3901 (N_3901,N_3721,N_3732);
and U3902 (N_3902,N_3757,N_3759);
nor U3903 (N_3903,N_3742,N_3723);
and U3904 (N_3904,N_3825,N_3687);
or U3905 (N_3905,N_3763,N_3706);
nor U3906 (N_3906,N_3805,N_3817);
or U3907 (N_3907,N_3701,N_3684);
nor U3908 (N_3908,N_3755,N_3809);
and U3909 (N_3909,N_3680,N_3736);
xnor U3910 (N_3910,N_3803,N_3753);
or U3911 (N_3911,N_3819,N_3818);
xor U3912 (N_3912,N_3827,N_3821);
and U3913 (N_3913,N_3729,N_3830);
or U3914 (N_3914,N_3709,N_3767);
xnor U3915 (N_3915,N_3773,N_3839);
or U3916 (N_3916,N_3756,N_3829);
nor U3917 (N_3917,N_3820,N_3748);
xnor U3918 (N_3918,N_3685,N_3711);
and U3919 (N_3919,N_3833,N_3810);
xor U3920 (N_3920,N_3758,N_3761);
nand U3921 (N_3921,N_3814,N_3734);
nand U3922 (N_3922,N_3804,N_3682);
xnor U3923 (N_3923,N_3749,N_3761);
nand U3924 (N_3924,N_3760,N_3817);
nor U3925 (N_3925,N_3797,N_3775);
xor U3926 (N_3926,N_3735,N_3827);
nand U3927 (N_3927,N_3839,N_3777);
nor U3928 (N_3928,N_3835,N_3729);
nand U3929 (N_3929,N_3753,N_3794);
and U3930 (N_3930,N_3775,N_3725);
xnor U3931 (N_3931,N_3810,N_3705);
and U3932 (N_3932,N_3837,N_3745);
xnor U3933 (N_3933,N_3753,N_3831);
nor U3934 (N_3934,N_3784,N_3832);
xor U3935 (N_3935,N_3712,N_3760);
xor U3936 (N_3936,N_3745,N_3729);
nor U3937 (N_3937,N_3714,N_3687);
nand U3938 (N_3938,N_3700,N_3810);
nor U3939 (N_3939,N_3680,N_3752);
or U3940 (N_3940,N_3762,N_3741);
and U3941 (N_3941,N_3815,N_3750);
nand U3942 (N_3942,N_3827,N_3786);
or U3943 (N_3943,N_3739,N_3815);
nand U3944 (N_3944,N_3709,N_3700);
xnor U3945 (N_3945,N_3693,N_3682);
nor U3946 (N_3946,N_3696,N_3824);
or U3947 (N_3947,N_3718,N_3785);
or U3948 (N_3948,N_3730,N_3760);
and U3949 (N_3949,N_3780,N_3699);
xor U3950 (N_3950,N_3798,N_3775);
xor U3951 (N_3951,N_3807,N_3759);
or U3952 (N_3952,N_3763,N_3837);
nor U3953 (N_3953,N_3812,N_3733);
xor U3954 (N_3954,N_3709,N_3730);
and U3955 (N_3955,N_3746,N_3712);
nor U3956 (N_3956,N_3738,N_3809);
and U3957 (N_3957,N_3704,N_3773);
and U3958 (N_3958,N_3766,N_3742);
and U3959 (N_3959,N_3743,N_3683);
nor U3960 (N_3960,N_3709,N_3729);
nor U3961 (N_3961,N_3706,N_3762);
xor U3962 (N_3962,N_3810,N_3698);
nor U3963 (N_3963,N_3828,N_3685);
nor U3964 (N_3964,N_3810,N_3689);
xor U3965 (N_3965,N_3832,N_3684);
or U3966 (N_3966,N_3774,N_3836);
xnor U3967 (N_3967,N_3802,N_3786);
nor U3968 (N_3968,N_3689,N_3765);
nor U3969 (N_3969,N_3721,N_3813);
nor U3970 (N_3970,N_3709,N_3715);
xnor U3971 (N_3971,N_3745,N_3712);
xnor U3972 (N_3972,N_3828,N_3785);
nand U3973 (N_3973,N_3834,N_3801);
nor U3974 (N_3974,N_3781,N_3691);
xnor U3975 (N_3975,N_3803,N_3687);
and U3976 (N_3976,N_3709,N_3687);
xnor U3977 (N_3977,N_3706,N_3764);
xor U3978 (N_3978,N_3703,N_3808);
xnor U3979 (N_3979,N_3764,N_3715);
and U3980 (N_3980,N_3703,N_3830);
or U3981 (N_3981,N_3783,N_3720);
or U3982 (N_3982,N_3732,N_3769);
nor U3983 (N_3983,N_3829,N_3776);
xnor U3984 (N_3984,N_3825,N_3748);
and U3985 (N_3985,N_3738,N_3768);
and U3986 (N_3986,N_3739,N_3691);
or U3987 (N_3987,N_3757,N_3684);
xor U3988 (N_3988,N_3732,N_3812);
and U3989 (N_3989,N_3744,N_3719);
or U3990 (N_3990,N_3838,N_3685);
xnor U3991 (N_3991,N_3704,N_3686);
and U3992 (N_3992,N_3779,N_3774);
or U3993 (N_3993,N_3830,N_3792);
nand U3994 (N_3994,N_3838,N_3760);
xnor U3995 (N_3995,N_3732,N_3705);
or U3996 (N_3996,N_3754,N_3801);
nand U3997 (N_3997,N_3780,N_3747);
xnor U3998 (N_3998,N_3783,N_3797);
nand U3999 (N_3999,N_3730,N_3824);
nor U4000 (N_4000,N_3963,N_3858);
and U4001 (N_4001,N_3931,N_3846);
or U4002 (N_4002,N_3960,N_3987);
nand U4003 (N_4003,N_3887,N_3978);
nor U4004 (N_4004,N_3943,N_3955);
nand U4005 (N_4005,N_3967,N_3995);
or U4006 (N_4006,N_3906,N_3958);
nor U4007 (N_4007,N_3916,N_3965);
nand U4008 (N_4008,N_3927,N_3882);
xor U4009 (N_4009,N_3855,N_3971);
nor U4010 (N_4010,N_3873,N_3870);
nor U4011 (N_4011,N_3899,N_3973);
or U4012 (N_4012,N_3940,N_3966);
xnor U4013 (N_4013,N_3881,N_3984);
and U4014 (N_4014,N_3935,N_3879);
nand U4015 (N_4015,N_3944,N_3889);
nor U4016 (N_4016,N_3853,N_3996);
nor U4017 (N_4017,N_3864,N_3908);
nor U4018 (N_4018,N_3917,N_3945);
nand U4019 (N_4019,N_3961,N_3932);
nand U4020 (N_4020,N_3861,N_3918);
xnor U4021 (N_4021,N_3980,N_3901);
nand U4022 (N_4022,N_3957,N_3883);
nor U4023 (N_4023,N_3854,N_3851);
or U4024 (N_4024,N_3841,N_3868);
and U4025 (N_4025,N_3909,N_3856);
nand U4026 (N_4026,N_3869,N_3922);
nand U4027 (N_4027,N_3840,N_3900);
xnor U4028 (N_4028,N_3974,N_3952);
or U4029 (N_4029,N_3992,N_3976);
xnor U4030 (N_4030,N_3907,N_3885);
nor U4031 (N_4031,N_3993,N_3956);
nor U4032 (N_4032,N_3913,N_3894);
nand U4033 (N_4033,N_3937,N_3939);
nor U4034 (N_4034,N_3852,N_3949);
nor U4035 (N_4035,N_3941,N_3897);
xor U4036 (N_4036,N_3857,N_3994);
nor U4037 (N_4037,N_3926,N_3878);
or U4038 (N_4038,N_3863,N_3884);
nor U4039 (N_4039,N_3871,N_3847);
and U4040 (N_4040,N_3942,N_3982);
nor U4041 (N_4041,N_3876,N_3977);
nor U4042 (N_4042,N_3979,N_3880);
or U4043 (N_4043,N_3999,N_3891);
or U4044 (N_4044,N_3997,N_3924);
nand U4045 (N_4045,N_3842,N_3890);
xnor U4046 (N_4046,N_3972,N_3865);
or U4047 (N_4047,N_3872,N_3920);
and U4048 (N_4048,N_3948,N_3923);
nand U4049 (N_4049,N_3929,N_3866);
or U4050 (N_4050,N_3962,N_3896);
and U4051 (N_4051,N_3975,N_3990);
or U4052 (N_4052,N_3911,N_3875);
and U4053 (N_4053,N_3985,N_3933);
nor U4054 (N_4054,N_3969,N_3968);
and U4055 (N_4055,N_3910,N_3951);
nand U4056 (N_4056,N_3893,N_3859);
xnor U4057 (N_4057,N_3845,N_3848);
nor U4058 (N_4058,N_3874,N_3912);
and U4059 (N_4059,N_3928,N_3895);
nor U4060 (N_4060,N_3877,N_3862);
or U4061 (N_4061,N_3914,N_3970);
xor U4062 (N_4062,N_3954,N_3938);
xnor U4063 (N_4063,N_3892,N_3843);
nand U4064 (N_4064,N_3860,N_3867);
nor U4065 (N_4065,N_3959,N_3844);
xor U4066 (N_4066,N_3981,N_3915);
nand U4067 (N_4067,N_3898,N_3919);
nand U4068 (N_4068,N_3936,N_3930);
nand U4069 (N_4069,N_3888,N_3983);
or U4070 (N_4070,N_3886,N_3989);
and U4071 (N_4071,N_3998,N_3964);
xor U4072 (N_4072,N_3905,N_3947);
and U4073 (N_4073,N_3902,N_3849);
and U4074 (N_4074,N_3850,N_3991);
xor U4075 (N_4075,N_3950,N_3925);
nand U4076 (N_4076,N_3904,N_3953);
xnor U4077 (N_4077,N_3988,N_3946);
nor U4078 (N_4078,N_3903,N_3934);
xnor U4079 (N_4079,N_3986,N_3921);
nand U4080 (N_4080,N_3953,N_3998);
nor U4081 (N_4081,N_3896,N_3978);
nor U4082 (N_4082,N_3992,N_3912);
or U4083 (N_4083,N_3914,N_3878);
nor U4084 (N_4084,N_3952,N_3879);
nand U4085 (N_4085,N_3955,N_3950);
and U4086 (N_4086,N_3974,N_3972);
or U4087 (N_4087,N_3923,N_3853);
nor U4088 (N_4088,N_3954,N_3953);
or U4089 (N_4089,N_3868,N_3918);
and U4090 (N_4090,N_3880,N_3861);
xor U4091 (N_4091,N_3874,N_3986);
nand U4092 (N_4092,N_3905,N_3918);
and U4093 (N_4093,N_3995,N_3900);
and U4094 (N_4094,N_3922,N_3881);
or U4095 (N_4095,N_3873,N_3954);
and U4096 (N_4096,N_3968,N_3998);
nand U4097 (N_4097,N_3884,N_3996);
nor U4098 (N_4098,N_3883,N_3972);
nand U4099 (N_4099,N_3971,N_3967);
nor U4100 (N_4100,N_3984,N_3914);
nand U4101 (N_4101,N_3860,N_3858);
nand U4102 (N_4102,N_3960,N_3936);
xnor U4103 (N_4103,N_3950,N_3958);
nand U4104 (N_4104,N_3865,N_3937);
and U4105 (N_4105,N_3898,N_3883);
and U4106 (N_4106,N_3958,N_3886);
nor U4107 (N_4107,N_3849,N_3973);
and U4108 (N_4108,N_3970,N_3847);
xor U4109 (N_4109,N_3854,N_3968);
nand U4110 (N_4110,N_3846,N_3948);
and U4111 (N_4111,N_3876,N_3852);
xnor U4112 (N_4112,N_3885,N_3864);
or U4113 (N_4113,N_3935,N_3918);
or U4114 (N_4114,N_3873,N_3894);
nor U4115 (N_4115,N_3886,N_3955);
and U4116 (N_4116,N_3880,N_3892);
xor U4117 (N_4117,N_3961,N_3928);
or U4118 (N_4118,N_3926,N_3856);
xor U4119 (N_4119,N_3922,N_3987);
nor U4120 (N_4120,N_3887,N_3969);
xnor U4121 (N_4121,N_3845,N_3909);
nor U4122 (N_4122,N_3957,N_3911);
and U4123 (N_4123,N_3933,N_3894);
nand U4124 (N_4124,N_3937,N_3978);
nor U4125 (N_4125,N_3985,N_3909);
nand U4126 (N_4126,N_3909,N_3866);
and U4127 (N_4127,N_3944,N_3908);
or U4128 (N_4128,N_3937,N_3987);
and U4129 (N_4129,N_3875,N_3918);
xor U4130 (N_4130,N_3927,N_3944);
nand U4131 (N_4131,N_3881,N_3854);
nor U4132 (N_4132,N_3961,N_3924);
and U4133 (N_4133,N_3904,N_3847);
and U4134 (N_4134,N_3996,N_3874);
nand U4135 (N_4135,N_3893,N_3953);
xor U4136 (N_4136,N_3993,N_3962);
nand U4137 (N_4137,N_3977,N_3972);
or U4138 (N_4138,N_3954,N_3872);
xor U4139 (N_4139,N_3883,N_3977);
nand U4140 (N_4140,N_3925,N_3937);
or U4141 (N_4141,N_3911,N_3964);
or U4142 (N_4142,N_3998,N_3980);
nor U4143 (N_4143,N_3868,N_3905);
nand U4144 (N_4144,N_3906,N_3909);
nor U4145 (N_4145,N_3856,N_3878);
nand U4146 (N_4146,N_3912,N_3842);
xor U4147 (N_4147,N_3998,N_3948);
and U4148 (N_4148,N_3902,N_3933);
nor U4149 (N_4149,N_3842,N_3847);
or U4150 (N_4150,N_3957,N_3931);
and U4151 (N_4151,N_3969,N_3966);
and U4152 (N_4152,N_3889,N_3947);
xnor U4153 (N_4153,N_3935,N_3967);
nor U4154 (N_4154,N_3945,N_3908);
and U4155 (N_4155,N_3883,N_3856);
nor U4156 (N_4156,N_3931,N_3858);
xnor U4157 (N_4157,N_3964,N_3899);
nor U4158 (N_4158,N_3941,N_3867);
xor U4159 (N_4159,N_3976,N_3921);
nand U4160 (N_4160,N_4019,N_4077);
nor U4161 (N_4161,N_4099,N_4010);
and U4162 (N_4162,N_4082,N_4123);
xor U4163 (N_4163,N_4156,N_4104);
nand U4164 (N_4164,N_4141,N_4017);
xor U4165 (N_4165,N_4086,N_4041);
xnor U4166 (N_4166,N_4130,N_4052);
or U4167 (N_4167,N_4028,N_4014);
and U4168 (N_4168,N_4092,N_4125);
nand U4169 (N_4169,N_4039,N_4040);
nor U4170 (N_4170,N_4036,N_4091);
nor U4171 (N_4171,N_4064,N_4023);
nand U4172 (N_4172,N_4047,N_4158);
or U4173 (N_4173,N_4100,N_4006);
and U4174 (N_4174,N_4000,N_4081);
or U4175 (N_4175,N_4089,N_4129);
and U4176 (N_4176,N_4011,N_4002);
nor U4177 (N_4177,N_4085,N_4094);
xnor U4178 (N_4178,N_4061,N_4070);
and U4179 (N_4179,N_4003,N_4018);
xnor U4180 (N_4180,N_4118,N_4119);
nor U4181 (N_4181,N_4049,N_4053);
nand U4182 (N_4182,N_4126,N_4078);
nor U4183 (N_4183,N_4150,N_4080);
xor U4184 (N_4184,N_4043,N_4140);
nand U4185 (N_4185,N_4020,N_4009);
nor U4186 (N_4186,N_4055,N_4005);
nand U4187 (N_4187,N_4046,N_4026);
xnor U4188 (N_4188,N_4157,N_4124);
or U4189 (N_4189,N_4012,N_4074);
nand U4190 (N_4190,N_4030,N_4110);
and U4191 (N_4191,N_4044,N_4144);
xnor U4192 (N_4192,N_4122,N_4108);
nor U4193 (N_4193,N_4071,N_4143);
nor U4194 (N_4194,N_4051,N_4131);
nor U4195 (N_4195,N_4146,N_4058);
nand U4196 (N_4196,N_4139,N_4084);
nor U4197 (N_4197,N_4145,N_4107);
or U4198 (N_4198,N_4112,N_4135);
nor U4199 (N_4199,N_4022,N_4132);
nor U4200 (N_4200,N_4054,N_4062);
and U4201 (N_4201,N_4027,N_4034);
xnor U4202 (N_4202,N_4095,N_4153);
nand U4203 (N_4203,N_4117,N_4016);
or U4204 (N_4204,N_4083,N_4024);
nand U4205 (N_4205,N_4076,N_4103);
and U4206 (N_4206,N_4008,N_4015);
nor U4207 (N_4207,N_4148,N_4045);
xor U4208 (N_4208,N_4075,N_4121);
nand U4209 (N_4209,N_4134,N_4115);
and U4210 (N_4210,N_4072,N_4066);
and U4211 (N_4211,N_4065,N_4127);
and U4212 (N_4212,N_4098,N_4021);
and U4213 (N_4213,N_4013,N_4067);
nand U4214 (N_4214,N_4059,N_4001);
or U4215 (N_4215,N_4137,N_4154);
xor U4216 (N_4216,N_4031,N_4048);
xor U4217 (N_4217,N_4057,N_4079);
xor U4218 (N_4218,N_4090,N_4063);
nor U4219 (N_4219,N_4152,N_4136);
and U4220 (N_4220,N_4105,N_4147);
xnor U4221 (N_4221,N_4068,N_4138);
or U4222 (N_4222,N_4142,N_4056);
xor U4223 (N_4223,N_4106,N_4042);
nor U4224 (N_4224,N_4101,N_4037);
xnor U4225 (N_4225,N_4073,N_4109);
xnor U4226 (N_4226,N_4032,N_4113);
nand U4227 (N_4227,N_4060,N_4133);
xnor U4228 (N_4228,N_4007,N_4111);
nor U4229 (N_4229,N_4093,N_4151);
or U4230 (N_4230,N_4159,N_4116);
and U4231 (N_4231,N_4035,N_4155);
nor U4232 (N_4232,N_4114,N_4050);
nor U4233 (N_4233,N_4004,N_4088);
and U4234 (N_4234,N_4033,N_4038);
nor U4235 (N_4235,N_4149,N_4097);
nor U4236 (N_4236,N_4096,N_4128);
xnor U4237 (N_4237,N_4120,N_4069);
nand U4238 (N_4238,N_4025,N_4029);
or U4239 (N_4239,N_4102,N_4087);
nand U4240 (N_4240,N_4037,N_4151);
nor U4241 (N_4241,N_4155,N_4053);
xor U4242 (N_4242,N_4041,N_4050);
and U4243 (N_4243,N_4012,N_4150);
and U4244 (N_4244,N_4099,N_4117);
nor U4245 (N_4245,N_4108,N_4042);
and U4246 (N_4246,N_4068,N_4022);
and U4247 (N_4247,N_4134,N_4015);
xnor U4248 (N_4248,N_4051,N_4017);
and U4249 (N_4249,N_4002,N_4114);
xor U4250 (N_4250,N_4152,N_4146);
xor U4251 (N_4251,N_4144,N_4085);
xnor U4252 (N_4252,N_4112,N_4155);
xor U4253 (N_4253,N_4085,N_4153);
nand U4254 (N_4254,N_4057,N_4027);
xnor U4255 (N_4255,N_4102,N_4024);
and U4256 (N_4256,N_4113,N_4076);
and U4257 (N_4257,N_4151,N_4148);
nor U4258 (N_4258,N_4082,N_4020);
nor U4259 (N_4259,N_4008,N_4076);
nor U4260 (N_4260,N_4025,N_4014);
nand U4261 (N_4261,N_4096,N_4056);
and U4262 (N_4262,N_4041,N_4084);
nor U4263 (N_4263,N_4141,N_4143);
nand U4264 (N_4264,N_4140,N_4024);
xor U4265 (N_4265,N_4153,N_4096);
xnor U4266 (N_4266,N_4107,N_4069);
and U4267 (N_4267,N_4005,N_4069);
and U4268 (N_4268,N_4131,N_4092);
or U4269 (N_4269,N_4043,N_4014);
nand U4270 (N_4270,N_4025,N_4115);
xor U4271 (N_4271,N_4128,N_4111);
nor U4272 (N_4272,N_4127,N_4154);
or U4273 (N_4273,N_4143,N_4035);
and U4274 (N_4274,N_4019,N_4001);
nor U4275 (N_4275,N_4044,N_4091);
or U4276 (N_4276,N_4037,N_4018);
or U4277 (N_4277,N_4108,N_4086);
nand U4278 (N_4278,N_4044,N_4063);
or U4279 (N_4279,N_4025,N_4137);
xnor U4280 (N_4280,N_4096,N_4084);
nor U4281 (N_4281,N_4140,N_4070);
or U4282 (N_4282,N_4035,N_4043);
and U4283 (N_4283,N_4127,N_4133);
nand U4284 (N_4284,N_4129,N_4143);
nand U4285 (N_4285,N_4060,N_4146);
nor U4286 (N_4286,N_4020,N_4084);
nand U4287 (N_4287,N_4044,N_4155);
xnor U4288 (N_4288,N_4142,N_4123);
or U4289 (N_4289,N_4159,N_4095);
and U4290 (N_4290,N_4114,N_4023);
or U4291 (N_4291,N_4157,N_4099);
and U4292 (N_4292,N_4022,N_4156);
or U4293 (N_4293,N_4017,N_4132);
nand U4294 (N_4294,N_4104,N_4055);
nand U4295 (N_4295,N_4154,N_4054);
nor U4296 (N_4296,N_4120,N_4136);
and U4297 (N_4297,N_4067,N_4027);
nand U4298 (N_4298,N_4103,N_4037);
or U4299 (N_4299,N_4036,N_4008);
nand U4300 (N_4300,N_4081,N_4118);
nand U4301 (N_4301,N_4073,N_4136);
nand U4302 (N_4302,N_4099,N_4142);
nor U4303 (N_4303,N_4115,N_4139);
or U4304 (N_4304,N_4057,N_4149);
or U4305 (N_4305,N_4156,N_4038);
or U4306 (N_4306,N_4060,N_4043);
xnor U4307 (N_4307,N_4133,N_4023);
and U4308 (N_4308,N_4029,N_4022);
or U4309 (N_4309,N_4052,N_4136);
nor U4310 (N_4310,N_4128,N_4030);
nor U4311 (N_4311,N_4008,N_4096);
xnor U4312 (N_4312,N_4085,N_4156);
nor U4313 (N_4313,N_4148,N_4063);
and U4314 (N_4314,N_4101,N_4128);
xnor U4315 (N_4315,N_4110,N_4141);
and U4316 (N_4316,N_4026,N_4019);
xor U4317 (N_4317,N_4082,N_4147);
nand U4318 (N_4318,N_4001,N_4061);
or U4319 (N_4319,N_4124,N_4097);
nor U4320 (N_4320,N_4177,N_4223);
nand U4321 (N_4321,N_4275,N_4227);
nand U4322 (N_4322,N_4285,N_4311);
nand U4323 (N_4323,N_4234,N_4165);
nor U4324 (N_4324,N_4233,N_4307);
nand U4325 (N_4325,N_4281,N_4312);
nand U4326 (N_4326,N_4197,N_4248);
xor U4327 (N_4327,N_4259,N_4161);
and U4328 (N_4328,N_4215,N_4310);
xor U4329 (N_4329,N_4237,N_4218);
or U4330 (N_4330,N_4195,N_4246);
xnor U4331 (N_4331,N_4306,N_4256);
or U4332 (N_4332,N_4305,N_4203);
nor U4333 (N_4333,N_4180,N_4304);
or U4334 (N_4334,N_4172,N_4198);
nand U4335 (N_4335,N_4302,N_4283);
nor U4336 (N_4336,N_4219,N_4191);
nor U4337 (N_4337,N_4228,N_4258);
and U4338 (N_4338,N_4287,N_4313);
xnor U4339 (N_4339,N_4202,N_4231);
and U4340 (N_4340,N_4178,N_4199);
xor U4341 (N_4341,N_4261,N_4254);
xor U4342 (N_4342,N_4221,N_4235);
nand U4343 (N_4343,N_4297,N_4303);
or U4344 (N_4344,N_4170,N_4249);
and U4345 (N_4345,N_4205,N_4189);
nand U4346 (N_4346,N_4296,N_4271);
and U4347 (N_4347,N_4225,N_4187);
or U4348 (N_4348,N_4182,N_4222);
nor U4349 (N_4349,N_4168,N_4290);
nor U4350 (N_4350,N_4266,N_4282);
or U4351 (N_4351,N_4192,N_4267);
xnor U4352 (N_4352,N_4298,N_4299);
or U4353 (N_4353,N_4229,N_4272);
or U4354 (N_4354,N_4263,N_4174);
or U4355 (N_4355,N_4244,N_4179);
and U4356 (N_4356,N_4190,N_4232);
nor U4357 (N_4357,N_4318,N_4279);
nor U4358 (N_4358,N_4242,N_4186);
or U4359 (N_4359,N_4276,N_4300);
nand U4360 (N_4360,N_4280,N_4269);
nand U4361 (N_4361,N_4288,N_4204);
xnor U4362 (N_4362,N_4220,N_4257);
or U4363 (N_4363,N_4243,N_4175);
or U4364 (N_4364,N_4314,N_4260);
or U4365 (N_4365,N_4309,N_4301);
xnor U4366 (N_4366,N_4316,N_4274);
nand U4367 (N_4367,N_4210,N_4163);
nor U4368 (N_4368,N_4265,N_4245);
nand U4369 (N_4369,N_4238,N_4201);
nor U4370 (N_4370,N_4188,N_4236);
and U4371 (N_4371,N_4185,N_4286);
xor U4372 (N_4372,N_4268,N_4241);
xor U4373 (N_4373,N_4291,N_4240);
and U4374 (N_4374,N_4169,N_4193);
nand U4375 (N_4375,N_4171,N_4270);
xnor U4376 (N_4376,N_4184,N_4176);
nor U4377 (N_4377,N_4200,N_4289);
nand U4378 (N_4378,N_4181,N_4224);
nor U4379 (N_4379,N_4213,N_4253);
xnor U4380 (N_4380,N_4217,N_4255);
or U4381 (N_4381,N_4206,N_4208);
nand U4382 (N_4382,N_4214,N_4292);
or U4383 (N_4383,N_4293,N_4284);
nor U4384 (N_4384,N_4194,N_4226);
and U4385 (N_4385,N_4162,N_4230);
xnor U4386 (N_4386,N_4315,N_4211);
and U4387 (N_4387,N_4209,N_4183);
xor U4388 (N_4388,N_4308,N_4294);
xor U4389 (N_4389,N_4239,N_4319);
nand U4390 (N_4390,N_4216,N_4196);
and U4391 (N_4391,N_4167,N_4160);
or U4392 (N_4392,N_4273,N_4247);
nand U4393 (N_4393,N_4264,N_4212);
xor U4394 (N_4394,N_4166,N_4317);
or U4395 (N_4395,N_4173,N_4295);
or U4396 (N_4396,N_4262,N_4251);
nand U4397 (N_4397,N_4250,N_4252);
nor U4398 (N_4398,N_4277,N_4164);
and U4399 (N_4399,N_4278,N_4207);
or U4400 (N_4400,N_4318,N_4237);
xnor U4401 (N_4401,N_4179,N_4197);
or U4402 (N_4402,N_4205,N_4281);
and U4403 (N_4403,N_4288,N_4227);
nand U4404 (N_4404,N_4251,N_4263);
or U4405 (N_4405,N_4260,N_4223);
nand U4406 (N_4406,N_4271,N_4231);
xor U4407 (N_4407,N_4304,N_4189);
nand U4408 (N_4408,N_4297,N_4196);
and U4409 (N_4409,N_4279,N_4273);
nor U4410 (N_4410,N_4305,N_4295);
nand U4411 (N_4411,N_4301,N_4183);
nor U4412 (N_4412,N_4171,N_4185);
nand U4413 (N_4413,N_4273,N_4301);
or U4414 (N_4414,N_4192,N_4234);
and U4415 (N_4415,N_4268,N_4174);
nor U4416 (N_4416,N_4161,N_4265);
nand U4417 (N_4417,N_4298,N_4291);
and U4418 (N_4418,N_4270,N_4261);
xnor U4419 (N_4419,N_4165,N_4204);
or U4420 (N_4420,N_4228,N_4197);
nor U4421 (N_4421,N_4309,N_4219);
or U4422 (N_4422,N_4279,N_4252);
nor U4423 (N_4423,N_4299,N_4224);
xnor U4424 (N_4424,N_4269,N_4299);
xor U4425 (N_4425,N_4291,N_4249);
nand U4426 (N_4426,N_4219,N_4222);
xnor U4427 (N_4427,N_4268,N_4180);
nor U4428 (N_4428,N_4267,N_4304);
or U4429 (N_4429,N_4176,N_4164);
and U4430 (N_4430,N_4311,N_4199);
nand U4431 (N_4431,N_4178,N_4280);
nor U4432 (N_4432,N_4199,N_4235);
or U4433 (N_4433,N_4257,N_4248);
nor U4434 (N_4434,N_4274,N_4259);
xor U4435 (N_4435,N_4287,N_4209);
nor U4436 (N_4436,N_4276,N_4266);
nor U4437 (N_4437,N_4260,N_4301);
xnor U4438 (N_4438,N_4229,N_4225);
or U4439 (N_4439,N_4251,N_4315);
xnor U4440 (N_4440,N_4250,N_4259);
or U4441 (N_4441,N_4180,N_4253);
and U4442 (N_4442,N_4269,N_4163);
nand U4443 (N_4443,N_4253,N_4287);
nor U4444 (N_4444,N_4268,N_4312);
or U4445 (N_4445,N_4213,N_4173);
nor U4446 (N_4446,N_4229,N_4223);
and U4447 (N_4447,N_4179,N_4237);
nor U4448 (N_4448,N_4270,N_4291);
nor U4449 (N_4449,N_4303,N_4288);
xnor U4450 (N_4450,N_4236,N_4303);
nor U4451 (N_4451,N_4279,N_4172);
and U4452 (N_4452,N_4266,N_4300);
nor U4453 (N_4453,N_4181,N_4205);
and U4454 (N_4454,N_4194,N_4310);
and U4455 (N_4455,N_4265,N_4232);
or U4456 (N_4456,N_4286,N_4190);
or U4457 (N_4457,N_4174,N_4210);
or U4458 (N_4458,N_4179,N_4165);
nor U4459 (N_4459,N_4271,N_4246);
nor U4460 (N_4460,N_4183,N_4281);
and U4461 (N_4461,N_4185,N_4179);
and U4462 (N_4462,N_4191,N_4278);
nor U4463 (N_4463,N_4180,N_4314);
and U4464 (N_4464,N_4312,N_4244);
nor U4465 (N_4465,N_4162,N_4220);
and U4466 (N_4466,N_4161,N_4221);
nor U4467 (N_4467,N_4161,N_4179);
nor U4468 (N_4468,N_4230,N_4225);
or U4469 (N_4469,N_4197,N_4287);
or U4470 (N_4470,N_4201,N_4248);
nand U4471 (N_4471,N_4211,N_4172);
xor U4472 (N_4472,N_4277,N_4300);
xnor U4473 (N_4473,N_4232,N_4222);
nor U4474 (N_4474,N_4301,N_4261);
or U4475 (N_4475,N_4222,N_4304);
or U4476 (N_4476,N_4211,N_4170);
nor U4477 (N_4477,N_4187,N_4238);
or U4478 (N_4478,N_4175,N_4318);
xor U4479 (N_4479,N_4232,N_4295);
or U4480 (N_4480,N_4435,N_4441);
xnor U4481 (N_4481,N_4360,N_4427);
and U4482 (N_4482,N_4364,N_4424);
or U4483 (N_4483,N_4358,N_4450);
xor U4484 (N_4484,N_4451,N_4438);
xnor U4485 (N_4485,N_4468,N_4334);
or U4486 (N_4486,N_4385,N_4343);
or U4487 (N_4487,N_4473,N_4446);
xnor U4488 (N_4488,N_4325,N_4444);
xor U4489 (N_4489,N_4331,N_4398);
or U4490 (N_4490,N_4426,N_4432);
xor U4491 (N_4491,N_4423,N_4390);
nand U4492 (N_4492,N_4357,N_4340);
or U4493 (N_4493,N_4412,N_4453);
nand U4494 (N_4494,N_4346,N_4365);
nand U4495 (N_4495,N_4342,N_4338);
nand U4496 (N_4496,N_4369,N_4479);
and U4497 (N_4497,N_4328,N_4387);
and U4498 (N_4498,N_4456,N_4406);
and U4499 (N_4499,N_4344,N_4367);
and U4500 (N_4500,N_4478,N_4349);
nand U4501 (N_4501,N_4467,N_4404);
nor U4502 (N_4502,N_4347,N_4341);
nor U4503 (N_4503,N_4442,N_4366);
and U4504 (N_4504,N_4335,N_4419);
xnor U4505 (N_4505,N_4322,N_4382);
xor U4506 (N_4506,N_4401,N_4374);
nor U4507 (N_4507,N_4437,N_4454);
or U4508 (N_4508,N_4397,N_4448);
nor U4509 (N_4509,N_4443,N_4372);
xnor U4510 (N_4510,N_4380,N_4428);
nand U4511 (N_4511,N_4420,N_4383);
nand U4512 (N_4512,N_4466,N_4355);
nor U4513 (N_4513,N_4330,N_4323);
xor U4514 (N_4514,N_4421,N_4471);
nand U4515 (N_4515,N_4407,N_4327);
nand U4516 (N_4516,N_4425,N_4470);
xnor U4517 (N_4517,N_4445,N_4408);
and U4518 (N_4518,N_4352,N_4475);
nand U4519 (N_4519,N_4395,N_4363);
or U4520 (N_4520,N_4458,N_4403);
xnor U4521 (N_4521,N_4461,N_4464);
nor U4522 (N_4522,N_4411,N_4400);
or U4523 (N_4523,N_4339,N_4359);
nand U4524 (N_4524,N_4459,N_4329);
xor U4525 (N_4525,N_4477,N_4351);
and U4526 (N_4526,N_4410,N_4345);
nand U4527 (N_4527,N_4409,N_4361);
and U4528 (N_4528,N_4350,N_4455);
xnor U4529 (N_4529,N_4353,N_4433);
and U4530 (N_4530,N_4393,N_4386);
or U4531 (N_4531,N_4326,N_4348);
nand U4532 (N_4532,N_4368,N_4447);
and U4533 (N_4533,N_4381,N_4333);
nor U4534 (N_4534,N_4431,N_4457);
nand U4535 (N_4535,N_4405,N_4388);
xor U4536 (N_4536,N_4414,N_4379);
nor U4537 (N_4537,N_4384,N_4332);
and U4538 (N_4538,N_4356,N_4416);
and U4539 (N_4539,N_4370,N_4371);
or U4540 (N_4540,N_4378,N_4440);
nand U4541 (N_4541,N_4429,N_4376);
or U4542 (N_4542,N_4465,N_4474);
xnor U4543 (N_4543,N_4321,N_4324);
xnor U4544 (N_4544,N_4422,N_4396);
and U4545 (N_4545,N_4430,N_4391);
and U4546 (N_4546,N_4462,N_4392);
nor U4547 (N_4547,N_4463,N_4362);
and U4548 (N_4548,N_4320,N_4399);
and U4549 (N_4549,N_4394,N_4434);
and U4550 (N_4550,N_4439,N_4402);
nor U4551 (N_4551,N_4452,N_4415);
xor U4552 (N_4552,N_4377,N_4460);
xor U4553 (N_4553,N_4354,N_4449);
and U4554 (N_4554,N_4389,N_4472);
xor U4555 (N_4555,N_4469,N_4337);
and U4556 (N_4556,N_4476,N_4418);
nor U4557 (N_4557,N_4417,N_4336);
or U4558 (N_4558,N_4373,N_4413);
or U4559 (N_4559,N_4436,N_4375);
and U4560 (N_4560,N_4454,N_4339);
nor U4561 (N_4561,N_4413,N_4472);
nor U4562 (N_4562,N_4350,N_4445);
nand U4563 (N_4563,N_4365,N_4428);
nor U4564 (N_4564,N_4432,N_4398);
or U4565 (N_4565,N_4451,N_4355);
xnor U4566 (N_4566,N_4454,N_4330);
and U4567 (N_4567,N_4420,N_4333);
xor U4568 (N_4568,N_4479,N_4323);
nor U4569 (N_4569,N_4421,N_4475);
or U4570 (N_4570,N_4407,N_4463);
and U4571 (N_4571,N_4388,N_4422);
or U4572 (N_4572,N_4378,N_4394);
or U4573 (N_4573,N_4387,N_4395);
nor U4574 (N_4574,N_4331,N_4435);
xnor U4575 (N_4575,N_4449,N_4468);
xnor U4576 (N_4576,N_4476,N_4375);
nand U4577 (N_4577,N_4470,N_4386);
and U4578 (N_4578,N_4447,N_4413);
nand U4579 (N_4579,N_4479,N_4356);
or U4580 (N_4580,N_4395,N_4477);
and U4581 (N_4581,N_4426,N_4404);
and U4582 (N_4582,N_4443,N_4396);
xor U4583 (N_4583,N_4327,N_4383);
xor U4584 (N_4584,N_4378,N_4448);
nor U4585 (N_4585,N_4432,N_4397);
nand U4586 (N_4586,N_4447,N_4326);
or U4587 (N_4587,N_4443,N_4354);
xnor U4588 (N_4588,N_4393,N_4392);
and U4589 (N_4589,N_4346,N_4429);
and U4590 (N_4590,N_4427,N_4378);
nor U4591 (N_4591,N_4467,N_4380);
nor U4592 (N_4592,N_4339,N_4336);
or U4593 (N_4593,N_4395,N_4353);
xnor U4594 (N_4594,N_4402,N_4394);
xnor U4595 (N_4595,N_4339,N_4390);
xor U4596 (N_4596,N_4366,N_4470);
or U4597 (N_4597,N_4423,N_4444);
xor U4598 (N_4598,N_4475,N_4383);
nor U4599 (N_4599,N_4379,N_4356);
and U4600 (N_4600,N_4420,N_4419);
or U4601 (N_4601,N_4414,N_4396);
and U4602 (N_4602,N_4447,N_4346);
nor U4603 (N_4603,N_4407,N_4359);
nand U4604 (N_4604,N_4360,N_4420);
or U4605 (N_4605,N_4324,N_4326);
nor U4606 (N_4606,N_4355,N_4348);
nor U4607 (N_4607,N_4354,N_4321);
and U4608 (N_4608,N_4396,N_4463);
or U4609 (N_4609,N_4343,N_4452);
or U4610 (N_4610,N_4385,N_4388);
or U4611 (N_4611,N_4392,N_4442);
nor U4612 (N_4612,N_4414,N_4441);
or U4613 (N_4613,N_4434,N_4350);
or U4614 (N_4614,N_4370,N_4383);
nand U4615 (N_4615,N_4425,N_4446);
nor U4616 (N_4616,N_4416,N_4377);
and U4617 (N_4617,N_4468,N_4433);
xnor U4618 (N_4618,N_4343,N_4437);
nor U4619 (N_4619,N_4358,N_4353);
nor U4620 (N_4620,N_4350,N_4337);
xnor U4621 (N_4621,N_4411,N_4354);
or U4622 (N_4622,N_4454,N_4379);
and U4623 (N_4623,N_4327,N_4324);
and U4624 (N_4624,N_4391,N_4372);
nand U4625 (N_4625,N_4357,N_4331);
nand U4626 (N_4626,N_4334,N_4406);
nand U4627 (N_4627,N_4455,N_4409);
nor U4628 (N_4628,N_4397,N_4361);
and U4629 (N_4629,N_4378,N_4339);
or U4630 (N_4630,N_4329,N_4392);
or U4631 (N_4631,N_4337,N_4415);
xor U4632 (N_4632,N_4439,N_4438);
and U4633 (N_4633,N_4349,N_4419);
nor U4634 (N_4634,N_4468,N_4329);
nor U4635 (N_4635,N_4339,N_4346);
nand U4636 (N_4636,N_4443,N_4412);
and U4637 (N_4637,N_4382,N_4337);
nand U4638 (N_4638,N_4363,N_4436);
nor U4639 (N_4639,N_4446,N_4378);
nand U4640 (N_4640,N_4506,N_4582);
xor U4641 (N_4641,N_4619,N_4508);
xnor U4642 (N_4642,N_4530,N_4614);
xnor U4643 (N_4643,N_4586,N_4529);
nor U4644 (N_4644,N_4537,N_4617);
and U4645 (N_4645,N_4494,N_4588);
or U4646 (N_4646,N_4516,N_4553);
xor U4647 (N_4647,N_4594,N_4579);
and U4648 (N_4648,N_4603,N_4633);
or U4649 (N_4649,N_4544,N_4499);
nor U4650 (N_4650,N_4576,N_4597);
nand U4651 (N_4651,N_4492,N_4543);
or U4652 (N_4652,N_4518,N_4638);
xnor U4653 (N_4653,N_4622,N_4480);
nand U4654 (N_4654,N_4482,N_4496);
or U4655 (N_4655,N_4570,N_4564);
or U4656 (N_4656,N_4495,N_4573);
or U4657 (N_4657,N_4637,N_4624);
xor U4658 (N_4658,N_4599,N_4629);
and U4659 (N_4659,N_4571,N_4558);
nand U4660 (N_4660,N_4528,N_4612);
nand U4661 (N_4661,N_4504,N_4590);
nor U4662 (N_4662,N_4627,N_4519);
xnor U4663 (N_4663,N_4541,N_4538);
nand U4664 (N_4664,N_4595,N_4623);
nor U4665 (N_4665,N_4636,N_4490);
or U4666 (N_4666,N_4567,N_4610);
xnor U4667 (N_4667,N_4531,N_4565);
nand U4668 (N_4668,N_4539,N_4502);
nand U4669 (N_4669,N_4505,N_4489);
and U4670 (N_4670,N_4555,N_4549);
nand U4671 (N_4671,N_4632,N_4561);
xor U4672 (N_4672,N_4596,N_4601);
nor U4673 (N_4673,N_4551,N_4552);
or U4674 (N_4674,N_4536,N_4493);
xor U4675 (N_4675,N_4540,N_4483);
nand U4676 (N_4676,N_4510,N_4584);
nand U4677 (N_4677,N_4542,N_4498);
nor U4678 (N_4678,N_4592,N_4611);
and U4679 (N_4679,N_4522,N_4556);
and U4680 (N_4680,N_4618,N_4525);
nand U4681 (N_4681,N_4589,N_4604);
nor U4682 (N_4682,N_4574,N_4503);
xnor U4683 (N_4683,N_4545,N_4491);
nor U4684 (N_4684,N_4534,N_4608);
or U4685 (N_4685,N_4520,N_4524);
xnor U4686 (N_4686,N_4560,N_4548);
nor U4687 (N_4687,N_4513,N_4606);
nand U4688 (N_4688,N_4569,N_4587);
and U4689 (N_4689,N_4550,N_4484);
xor U4690 (N_4690,N_4581,N_4532);
or U4691 (N_4691,N_4523,N_4501);
xnor U4692 (N_4692,N_4563,N_4607);
or U4693 (N_4693,N_4631,N_4580);
nor U4694 (N_4694,N_4613,N_4527);
xor U4695 (N_4695,N_4609,N_4511);
and U4696 (N_4696,N_4562,N_4533);
or U4697 (N_4697,N_4507,N_4547);
xnor U4698 (N_4698,N_4616,N_4514);
and U4699 (N_4699,N_4605,N_4521);
and U4700 (N_4700,N_4535,N_4630);
nor U4701 (N_4701,N_4600,N_4578);
nand U4702 (N_4702,N_4639,N_4487);
xnor U4703 (N_4703,N_4585,N_4512);
nor U4704 (N_4704,N_4509,N_4628);
nor U4705 (N_4705,N_4488,N_4626);
and U4706 (N_4706,N_4577,N_4583);
nand U4707 (N_4707,N_4568,N_4602);
or U4708 (N_4708,N_4481,N_4615);
and U4709 (N_4709,N_4486,N_4515);
nand U4710 (N_4710,N_4485,N_4526);
or U4711 (N_4711,N_4635,N_4554);
and U4712 (N_4712,N_4572,N_4634);
xnor U4713 (N_4713,N_4566,N_4557);
nand U4714 (N_4714,N_4517,N_4625);
nand U4715 (N_4715,N_4500,N_4598);
nand U4716 (N_4716,N_4620,N_4591);
xor U4717 (N_4717,N_4546,N_4575);
nor U4718 (N_4718,N_4497,N_4559);
nand U4719 (N_4719,N_4621,N_4593);
or U4720 (N_4720,N_4494,N_4582);
nand U4721 (N_4721,N_4532,N_4612);
nor U4722 (N_4722,N_4541,N_4575);
xor U4723 (N_4723,N_4522,N_4551);
or U4724 (N_4724,N_4570,N_4595);
or U4725 (N_4725,N_4526,N_4518);
and U4726 (N_4726,N_4590,N_4522);
or U4727 (N_4727,N_4622,N_4549);
and U4728 (N_4728,N_4510,N_4530);
nand U4729 (N_4729,N_4592,N_4511);
nand U4730 (N_4730,N_4539,N_4630);
or U4731 (N_4731,N_4537,N_4573);
or U4732 (N_4732,N_4627,N_4597);
nor U4733 (N_4733,N_4608,N_4582);
nand U4734 (N_4734,N_4545,N_4586);
nand U4735 (N_4735,N_4517,N_4552);
nor U4736 (N_4736,N_4542,N_4484);
xnor U4737 (N_4737,N_4481,N_4523);
nor U4738 (N_4738,N_4554,N_4615);
or U4739 (N_4739,N_4566,N_4515);
nor U4740 (N_4740,N_4520,N_4495);
nor U4741 (N_4741,N_4503,N_4567);
nand U4742 (N_4742,N_4508,N_4572);
nor U4743 (N_4743,N_4491,N_4565);
or U4744 (N_4744,N_4618,N_4518);
nand U4745 (N_4745,N_4482,N_4639);
xor U4746 (N_4746,N_4541,N_4486);
or U4747 (N_4747,N_4521,N_4494);
or U4748 (N_4748,N_4504,N_4495);
or U4749 (N_4749,N_4598,N_4566);
nor U4750 (N_4750,N_4562,N_4565);
and U4751 (N_4751,N_4581,N_4515);
nor U4752 (N_4752,N_4510,N_4497);
nor U4753 (N_4753,N_4523,N_4613);
and U4754 (N_4754,N_4564,N_4501);
and U4755 (N_4755,N_4595,N_4504);
nand U4756 (N_4756,N_4527,N_4524);
nor U4757 (N_4757,N_4604,N_4480);
and U4758 (N_4758,N_4523,N_4510);
nand U4759 (N_4759,N_4628,N_4603);
or U4760 (N_4760,N_4553,N_4590);
or U4761 (N_4761,N_4591,N_4631);
nor U4762 (N_4762,N_4548,N_4580);
nand U4763 (N_4763,N_4614,N_4592);
nand U4764 (N_4764,N_4556,N_4614);
or U4765 (N_4765,N_4527,N_4616);
nor U4766 (N_4766,N_4530,N_4483);
and U4767 (N_4767,N_4629,N_4577);
or U4768 (N_4768,N_4574,N_4587);
nand U4769 (N_4769,N_4551,N_4515);
or U4770 (N_4770,N_4486,N_4554);
or U4771 (N_4771,N_4550,N_4492);
xnor U4772 (N_4772,N_4539,N_4497);
xnor U4773 (N_4773,N_4485,N_4579);
and U4774 (N_4774,N_4557,N_4518);
and U4775 (N_4775,N_4585,N_4545);
xnor U4776 (N_4776,N_4494,N_4600);
xor U4777 (N_4777,N_4544,N_4525);
or U4778 (N_4778,N_4568,N_4576);
and U4779 (N_4779,N_4491,N_4537);
xnor U4780 (N_4780,N_4492,N_4616);
or U4781 (N_4781,N_4493,N_4639);
nor U4782 (N_4782,N_4486,N_4587);
nor U4783 (N_4783,N_4542,N_4628);
nand U4784 (N_4784,N_4485,N_4482);
nand U4785 (N_4785,N_4570,N_4485);
and U4786 (N_4786,N_4575,N_4484);
and U4787 (N_4787,N_4589,N_4538);
xnor U4788 (N_4788,N_4541,N_4529);
or U4789 (N_4789,N_4519,N_4577);
xnor U4790 (N_4790,N_4625,N_4516);
and U4791 (N_4791,N_4560,N_4611);
nand U4792 (N_4792,N_4628,N_4579);
and U4793 (N_4793,N_4551,N_4532);
or U4794 (N_4794,N_4510,N_4594);
and U4795 (N_4795,N_4557,N_4487);
xor U4796 (N_4796,N_4573,N_4545);
and U4797 (N_4797,N_4560,N_4519);
nor U4798 (N_4798,N_4571,N_4615);
nor U4799 (N_4799,N_4595,N_4531);
or U4800 (N_4800,N_4737,N_4731);
nand U4801 (N_4801,N_4677,N_4797);
nor U4802 (N_4802,N_4670,N_4735);
nand U4803 (N_4803,N_4772,N_4722);
and U4804 (N_4804,N_4668,N_4712);
nor U4805 (N_4805,N_4643,N_4658);
nor U4806 (N_4806,N_4651,N_4657);
nand U4807 (N_4807,N_4793,N_4784);
or U4808 (N_4808,N_4669,N_4761);
xnor U4809 (N_4809,N_4650,N_4687);
or U4810 (N_4810,N_4771,N_4713);
nor U4811 (N_4811,N_4705,N_4799);
xnor U4812 (N_4812,N_4727,N_4640);
nand U4813 (N_4813,N_4641,N_4714);
nand U4814 (N_4814,N_4649,N_4773);
xor U4815 (N_4815,N_4752,N_4763);
and U4816 (N_4816,N_4749,N_4769);
and U4817 (N_4817,N_4718,N_4739);
and U4818 (N_4818,N_4674,N_4666);
xor U4819 (N_4819,N_4760,N_4715);
nand U4820 (N_4820,N_4787,N_4686);
xnor U4821 (N_4821,N_4711,N_4729);
or U4822 (N_4822,N_4781,N_4794);
and U4823 (N_4823,N_4779,N_4757);
xnor U4824 (N_4824,N_4782,N_4653);
xnor U4825 (N_4825,N_4768,N_4732);
xor U4826 (N_4826,N_4740,N_4764);
and U4827 (N_4827,N_4699,N_4770);
xor U4828 (N_4828,N_4742,N_4741);
or U4829 (N_4829,N_4788,N_4758);
nand U4830 (N_4830,N_4751,N_4673);
xor U4831 (N_4831,N_4746,N_4765);
and U4832 (N_4832,N_4682,N_4672);
xnor U4833 (N_4833,N_4691,N_4778);
nor U4834 (N_4834,N_4685,N_4780);
and U4835 (N_4835,N_4716,N_4690);
and U4836 (N_4836,N_4756,N_4744);
or U4837 (N_4837,N_4642,N_4681);
nand U4838 (N_4838,N_4725,N_4647);
xor U4839 (N_4839,N_4721,N_4717);
and U4840 (N_4840,N_4652,N_4697);
nor U4841 (N_4841,N_4724,N_4790);
and U4842 (N_4842,N_4707,N_4762);
nand U4843 (N_4843,N_4745,N_4678);
and U4844 (N_4844,N_4783,N_4703);
xnor U4845 (N_4845,N_4654,N_4750);
nor U4846 (N_4846,N_4700,N_4777);
nand U4847 (N_4847,N_4719,N_4680);
and U4848 (N_4848,N_4759,N_4648);
or U4849 (N_4849,N_4693,N_4734);
nor U4850 (N_4850,N_4694,N_4748);
xor U4851 (N_4851,N_4738,N_4692);
nor U4852 (N_4852,N_4710,N_4796);
or U4853 (N_4853,N_4706,N_4755);
nor U4854 (N_4854,N_4683,N_4730);
nor U4855 (N_4855,N_4728,N_4753);
nor U4856 (N_4856,N_4646,N_4667);
or U4857 (N_4857,N_4720,N_4688);
and U4858 (N_4858,N_4675,N_4655);
or U4859 (N_4859,N_4754,N_4665);
nand U4860 (N_4860,N_4791,N_4736);
or U4861 (N_4861,N_4659,N_4645);
and U4862 (N_4862,N_4695,N_4786);
nand U4863 (N_4863,N_4701,N_4774);
or U4864 (N_4864,N_4709,N_4671);
nor U4865 (N_4865,N_4776,N_4708);
nor U4866 (N_4866,N_4644,N_4789);
xnor U4867 (N_4867,N_4679,N_4733);
or U4868 (N_4868,N_4723,N_4702);
or U4869 (N_4869,N_4696,N_4798);
and U4870 (N_4870,N_4698,N_4743);
or U4871 (N_4871,N_4656,N_4662);
xnor U4872 (N_4872,N_4664,N_4747);
or U4873 (N_4873,N_4661,N_4689);
nor U4874 (N_4874,N_4726,N_4775);
nand U4875 (N_4875,N_4684,N_4660);
nor U4876 (N_4876,N_4704,N_4663);
and U4877 (N_4877,N_4792,N_4766);
and U4878 (N_4878,N_4795,N_4785);
nor U4879 (N_4879,N_4676,N_4767);
nor U4880 (N_4880,N_4651,N_4794);
xnor U4881 (N_4881,N_4758,N_4715);
nor U4882 (N_4882,N_4659,N_4795);
xor U4883 (N_4883,N_4786,N_4765);
and U4884 (N_4884,N_4789,N_4750);
nor U4885 (N_4885,N_4797,N_4757);
nor U4886 (N_4886,N_4725,N_4731);
and U4887 (N_4887,N_4690,N_4685);
and U4888 (N_4888,N_4772,N_4797);
xnor U4889 (N_4889,N_4736,N_4664);
and U4890 (N_4890,N_4751,N_4649);
or U4891 (N_4891,N_4749,N_4766);
nand U4892 (N_4892,N_4648,N_4771);
xnor U4893 (N_4893,N_4791,N_4747);
or U4894 (N_4894,N_4737,N_4701);
nor U4895 (N_4895,N_4671,N_4667);
xnor U4896 (N_4896,N_4774,N_4683);
xor U4897 (N_4897,N_4646,N_4687);
and U4898 (N_4898,N_4685,N_4734);
and U4899 (N_4899,N_4706,N_4719);
or U4900 (N_4900,N_4705,N_4741);
nor U4901 (N_4901,N_4640,N_4767);
and U4902 (N_4902,N_4683,N_4694);
nor U4903 (N_4903,N_4735,N_4742);
xnor U4904 (N_4904,N_4788,N_4780);
nor U4905 (N_4905,N_4771,N_4777);
nor U4906 (N_4906,N_4658,N_4770);
xor U4907 (N_4907,N_4712,N_4797);
and U4908 (N_4908,N_4733,N_4699);
xnor U4909 (N_4909,N_4733,N_4753);
or U4910 (N_4910,N_4674,N_4762);
nor U4911 (N_4911,N_4739,N_4728);
nor U4912 (N_4912,N_4739,N_4752);
xnor U4913 (N_4913,N_4773,N_4644);
nor U4914 (N_4914,N_4788,N_4658);
or U4915 (N_4915,N_4724,N_4683);
nand U4916 (N_4916,N_4680,N_4733);
xor U4917 (N_4917,N_4648,N_4691);
xor U4918 (N_4918,N_4641,N_4658);
nor U4919 (N_4919,N_4751,N_4718);
nor U4920 (N_4920,N_4700,N_4668);
or U4921 (N_4921,N_4772,N_4695);
or U4922 (N_4922,N_4765,N_4745);
nand U4923 (N_4923,N_4738,N_4761);
and U4924 (N_4924,N_4651,N_4707);
nand U4925 (N_4925,N_4702,N_4666);
xnor U4926 (N_4926,N_4752,N_4698);
nand U4927 (N_4927,N_4665,N_4755);
and U4928 (N_4928,N_4725,N_4799);
xor U4929 (N_4929,N_4708,N_4652);
nand U4930 (N_4930,N_4774,N_4730);
and U4931 (N_4931,N_4667,N_4651);
nand U4932 (N_4932,N_4717,N_4720);
or U4933 (N_4933,N_4717,N_4723);
and U4934 (N_4934,N_4726,N_4735);
nand U4935 (N_4935,N_4721,N_4760);
xnor U4936 (N_4936,N_4645,N_4748);
and U4937 (N_4937,N_4780,N_4669);
or U4938 (N_4938,N_4778,N_4713);
nor U4939 (N_4939,N_4781,N_4733);
and U4940 (N_4940,N_4774,N_4658);
nor U4941 (N_4941,N_4711,N_4660);
or U4942 (N_4942,N_4665,N_4685);
nor U4943 (N_4943,N_4753,N_4678);
and U4944 (N_4944,N_4727,N_4721);
xnor U4945 (N_4945,N_4754,N_4698);
xnor U4946 (N_4946,N_4674,N_4768);
nand U4947 (N_4947,N_4667,N_4645);
nor U4948 (N_4948,N_4700,N_4681);
xnor U4949 (N_4949,N_4649,N_4792);
nor U4950 (N_4950,N_4786,N_4665);
xor U4951 (N_4951,N_4752,N_4783);
nand U4952 (N_4952,N_4699,N_4674);
and U4953 (N_4953,N_4705,N_4678);
or U4954 (N_4954,N_4751,N_4736);
nor U4955 (N_4955,N_4652,N_4780);
nor U4956 (N_4956,N_4661,N_4731);
and U4957 (N_4957,N_4773,N_4770);
and U4958 (N_4958,N_4685,N_4688);
nand U4959 (N_4959,N_4717,N_4707);
xor U4960 (N_4960,N_4895,N_4832);
xor U4961 (N_4961,N_4877,N_4867);
and U4962 (N_4962,N_4901,N_4856);
xnor U4963 (N_4963,N_4853,N_4959);
nor U4964 (N_4964,N_4933,N_4891);
or U4965 (N_4965,N_4882,N_4879);
xnor U4966 (N_4966,N_4940,N_4814);
and U4967 (N_4967,N_4834,N_4905);
nor U4968 (N_4968,N_4805,N_4911);
nor U4969 (N_4969,N_4852,N_4806);
or U4970 (N_4970,N_4862,N_4836);
nand U4971 (N_4971,N_4843,N_4916);
nand U4972 (N_4972,N_4918,N_4939);
and U4973 (N_4973,N_4944,N_4954);
and U4974 (N_4974,N_4864,N_4909);
and U4975 (N_4975,N_4870,N_4899);
and U4976 (N_4976,N_4829,N_4898);
or U4977 (N_4977,N_4874,N_4889);
nor U4978 (N_4978,N_4925,N_4955);
and U4979 (N_4979,N_4854,N_4897);
xnor U4980 (N_4980,N_4850,N_4912);
and U4981 (N_4981,N_4841,N_4887);
nor U4982 (N_4982,N_4941,N_4845);
or U4983 (N_4983,N_4849,N_4902);
xor U4984 (N_4984,N_4858,N_4831);
nor U4985 (N_4985,N_4866,N_4908);
xor U4986 (N_4986,N_4943,N_4809);
nand U4987 (N_4987,N_4848,N_4921);
xnor U4988 (N_4988,N_4932,N_4930);
nor U4989 (N_4989,N_4885,N_4840);
xnor U4990 (N_4990,N_4802,N_4825);
and U4991 (N_4991,N_4817,N_4934);
nand U4992 (N_4992,N_4924,N_4839);
and U4993 (N_4993,N_4833,N_4926);
nand U4994 (N_4994,N_4938,N_4952);
or U4995 (N_4995,N_4903,N_4893);
and U4996 (N_4996,N_4824,N_4935);
and U4997 (N_4997,N_4917,N_4813);
nor U4998 (N_4998,N_4869,N_4865);
nor U4999 (N_4999,N_4804,N_4838);
nand U5000 (N_5000,N_4872,N_4931);
nand U5001 (N_5001,N_4950,N_4851);
nor U5002 (N_5002,N_4942,N_4894);
nand U5003 (N_5003,N_4880,N_4881);
or U5004 (N_5004,N_4807,N_4947);
xnor U5005 (N_5005,N_4928,N_4871);
nor U5006 (N_5006,N_4937,N_4949);
nor U5007 (N_5007,N_4946,N_4815);
or U5008 (N_5008,N_4810,N_4847);
nor U5009 (N_5009,N_4800,N_4886);
or U5010 (N_5010,N_4811,N_4922);
and U5011 (N_5011,N_4830,N_4859);
or U5012 (N_5012,N_4958,N_4868);
xor U5013 (N_5013,N_4883,N_4861);
and U5014 (N_5014,N_4822,N_4842);
xnor U5015 (N_5015,N_4803,N_4948);
xor U5016 (N_5016,N_4904,N_4808);
nand U5017 (N_5017,N_4857,N_4823);
and U5018 (N_5018,N_4827,N_4913);
xnor U5019 (N_5019,N_4855,N_4837);
and U5020 (N_5020,N_4884,N_4900);
or U5021 (N_5021,N_4863,N_4956);
and U5022 (N_5022,N_4860,N_4828);
xnor U5023 (N_5023,N_4910,N_4951);
or U5024 (N_5024,N_4945,N_4820);
or U5025 (N_5025,N_4927,N_4844);
nor U5026 (N_5026,N_4914,N_4801);
and U5027 (N_5027,N_4953,N_4907);
nand U5028 (N_5028,N_4920,N_4818);
xnor U5029 (N_5029,N_4957,N_4812);
xnor U5030 (N_5030,N_4906,N_4826);
and U5031 (N_5031,N_4876,N_4873);
xor U5032 (N_5032,N_4875,N_4915);
xor U5033 (N_5033,N_4816,N_4821);
or U5034 (N_5034,N_4896,N_4892);
nor U5035 (N_5035,N_4846,N_4919);
and U5036 (N_5036,N_4878,N_4819);
nor U5037 (N_5037,N_4890,N_4936);
nor U5038 (N_5038,N_4835,N_4923);
or U5039 (N_5039,N_4929,N_4888);
nand U5040 (N_5040,N_4856,N_4951);
nor U5041 (N_5041,N_4943,N_4893);
and U5042 (N_5042,N_4951,N_4881);
xor U5043 (N_5043,N_4953,N_4958);
and U5044 (N_5044,N_4896,N_4936);
xor U5045 (N_5045,N_4861,N_4806);
and U5046 (N_5046,N_4896,N_4822);
and U5047 (N_5047,N_4855,N_4819);
xor U5048 (N_5048,N_4817,N_4859);
and U5049 (N_5049,N_4894,N_4828);
xnor U5050 (N_5050,N_4939,N_4896);
and U5051 (N_5051,N_4882,N_4954);
nor U5052 (N_5052,N_4901,N_4937);
nand U5053 (N_5053,N_4890,N_4816);
nand U5054 (N_5054,N_4921,N_4955);
and U5055 (N_5055,N_4936,N_4893);
or U5056 (N_5056,N_4924,N_4957);
or U5057 (N_5057,N_4823,N_4848);
or U5058 (N_5058,N_4923,N_4921);
and U5059 (N_5059,N_4872,N_4899);
and U5060 (N_5060,N_4801,N_4802);
and U5061 (N_5061,N_4878,N_4814);
and U5062 (N_5062,N_4837,N_4880);
nand U5063 (N_5063,N_4886,N_4874);
or U5064 (N_5064,N_4815,N_4886);
nor U5065 (N_5065,N_4888,N_4937);
xor U5066 (N_5066,N_4881,N_4959);
or U5067 (N_5067,N_4948,N_4932);
nand U5068 (N_5068,N_4920,N_4820);
nand U5069 (N_5069,N_4897,N_4819);
or U5070 (N_5070,N_4852,N_4939);
and U5071 (N_5071,N_4901,N_4836);
nor U5072 (N_5072,N_4950,N_4878);
nor U5073 (N_5073,N_4883,N_4959);
or U5074 (N_5074,N_4939,N_4931);
or U5075 (N_5075,N_4808,N_4838);
nor U5076 (N_5076,N_4895,N_4843);
xnor U5077 (N_5077,N_4818,N_4844);
or U5078 (N_5078,N_4959,N_4843);
nor U5079 (N_5079,N_4922,N_4905);
nand U5080 (N_5080,N_4884,N_4806);
xor U5081 (N_5081,N_4833,N_4923);
or U5082 (N_5082,N_4950,N_4829);
xor U5083 (N_5083,N_4948,N_4849);
xnor U5084 (N_5084,N_4838,N_4858);
nor U5085 (N_5085,N_4903,N_4905);
or U5086 (N_5086,N_4957,N_4865);
or U5087 (N_5087,N_4834,N_4888);
or U5088 (N_5088,N_4902,N_4861);
and U5089 (N_5089,N_4838,N_4818);
nand U5090 (N_5090,N_4849,N_4884);
and U5091 (N_5091,N_4895,N_4824);
or U5092 (N_5092,N_4883,N_4934);
or U5093 (N_5093,N_4933,N_4881);
xnor U5094 (N_5094,N_4903,N_4912);
and U5095 (N_5095,N_4934,N_4816);
nor U5096 (N_5096,N_4888,N_4833);
or U5097 (N_5097,N_4829,N_4954);
and U5098 (N_5098,N_4906,N_4854);
xor U5099 (N_5099,N_4865,N_4896);
xor U5100 (N_5100,N_4873,N_4891);
nor U5101 (N_5101,N_4824,N_4920);
nand U5102 (N_5102,N_4837,N_4919);
or U5103 (N_5103,N_4811,N_4849);
and U5104 (N_5104,N_4899,N_4821);
or U5105 (N_5105,N_4848,N_4833);
or U5106 (N_5106,N_4943,N_4884);
or U5107 (N_5107,N_4809,N_4876);
xnor U5108 (N_5108,N_4839,N_4860);
or U5109 (N_5109,N_4954,N_4820);
nand U5110 (N_5110,N_4891,N_4838);
nor U5111 (N_5111,N_4800,N_4837);
xnor U5112 (N_5112,N_4805,N_4862);
and U5113 (N_5113,N_4892,N_4800);
or U5114 (N_5114,N_4879,N_4880);
nand U5115 (N_5115,N_4822,N_4893);
xnor U5116 (N_5116,N_4809,N_4840);
or U5117 (N_5117,N_4875,N_4841);
nand U5118 (N_5118,N_4840,N_4859);
xnor U5119 (N_5119,N_4871,N_4902);
xnor U5120 (N_5120,N_5082,N_5112);
nand U5121 (N_5121,N_5035,N_5015);
nor U5122 (N_5122,N_5044,N_4977);
or U5123 (N_5123,N_5024,N_5069);
nand U5124 (N_5124,N_5039,N_5116);
nor U5125 (N_5125,N_5048,N_4990);
xnor U5126 (N_5126,N_5041,N_5117);
nand U5127 (N_5127,N_5052,N_4995);
xor U5128 (N_5128,N_5088,N_5071);
nor U5129 (N_5129,N_4981,N_4999);
and U5130 (N_5130,N_5098,N_5103);
nor U5131 (N_5131,N_5115,N_5018);
and U5132 (N_5132,N_5000,N_4998);
nand U5133 (N_5133,N_5047,N_5080);
or U5134 (N_5134,N_4976,N_4963);
xor U5135 (N_5135,N_5101,N_5081);
and U5136 (N_5136,N_5066,N_5089);
nor U5137 (N_5137,N_5105,N_5063);
and U5138 (N_5138,N_5040,N_5085);
nor U5139 (N_5139,N_5006,N_5064);
nand U5140 (N_5140,N_5017,N_5072);
xor U5141 (N_5141,N_5097,N_4988);
or U5142 (N_5142,N_5113,N_5059);
nor U5143 (N_5143,N_5012,N_5104);
and U5144 (N_5144,N_5074,N_4989);
or U5145 (N_5145,N_5036,N_4997);
xnor U5146 (N_5146,N_5099,N_4994);
xnor U5147 (N_5147,N_4992,N_4965);
or U5148 (N_5148,N_5010,N_5013);
and U5149 (N_5149,N_5079,N_5026);
and U5150 (N_5150,N_5023,N_5030);
nor U5151 (N_5151,N_4969,N_5025);
nand U5152 (N_5152,N_4967,N_5095);
nor U5153 (N_5153,N_4960,N_4975);
or U5154 (N_5154,N_5092,N_5021);
xor U5155 (N_5155,N_5007,N_4985);
and U5156 (N_5156,N_5016,N_5019);
and U5157 (N_5157,N_5114,N_4964);
nand U5158 (N_5158,N_4974,N_5055);
nor U5159 (N_5159,N_5062,N_5093);
nand U5160 (N_5160,N_5091,N_5073);
nor U5161 (N_5161,N_5110,N_5083);
nor U5162 (N_5162,N_5054,N_5111);
nor U5163 (N_5163,N_5009,N_5086);
xnor U5164 (N_5164,N_5109,N_5100);
or U5165 (N_5165,N_5053,N_4986);
and U5166 (N_5166,N_5027,N_4983);
nor U5167 (N_5167,N_4972,N_5050);
xnor U5168 (N_5168,N_5102,N_5107);
nor U5169 (N_5169,N_4970,N_5042);
nand U5170 (N_5170,N_5078,N_5067);
and U5171 (N_5171,N_5051,N_5108);
nor U5172 (N_5172,N_5058,N_5032);
nor U5173 (N_5173,N_4979,N_4966);
xor U5174 (N_5174,N_5106,N_5029);
and U5175 (N_5175,N_5090,N_5119);
nand U5176 (N_5176,N_5094,N_4962);
nand U5177 (N_5177,N_5011,N_5031);
nand U5178 (N_5178,N_4973,N_5049);
nor U5179 (N_5179,N_5075,N_5056);
nand U5180 (N_5180,N_5005,N_5068);
or U5181 (N_5181,N_5034,N_4987);
or U5182 (N_5182,N_5038,N_4978);
or U5183 (N_5183,N_4968,N_5118);
or U5184 (N_5184,N_5004,N_5060);
xnor U5185 (N_5185,N_5077,N_4993);
or U5186 (N_5186,N_5076,N_4982);
nor U5187 (N_5187,N_5003,N_4971);
nor U5188 (N_5188,N_5022,N_5087);
or U5189 (N_5189,N_5037,N_5084);
xor U5190 (N_5190,N_4991,N_5045);
xnor U5191 (N_5191,N_5046,N_5043);
and U5192 (N_5192,N_5033,N_5070);
or U5193 (N_5193,N_4980,N_4961);
and U5194 (N_5194,N_5061,N_5002);
or U5195 (N_5195,N_4996,N_5028);
nand U5196 (N_5196,N_5096,N_5065);
or U5197 (N_5197,N_4984,N_5020);
nand U5198 (N_5198,N_5001,N_5057);
or U5199 (N_5199,N_5008,N_5014);
nand U5200 (N_5200,N_5092,N_4979);
and U5201 (N_5201,N_5013,N_5044);
nor U5202 (N_5202,N_5002,N_5041);
or U5203 (N_5203,N_5108,N_4966);
and U5204 (N_5204,N_5016,N_5117);
or U5205 (N_5205,N_4987,N_4985);
xor U5206 (N_5206,N_4985,N_5056);
nor U5207 (N_5207,N_5005,N_5080);
xor U5208 (N_5208,N_4996,N_5010);
xnor U5209 (N_5209,N_4960,N_5077);
and U5210 (N_5210,N_5081,N_4982);
or U5211 (N_5211,N_5045,N_5089);
or U5212 (N_5212,N_4969,N_5116);
nand U5213 (N_5213,N_5085,N_5053);
or U5214 (N_5214,N_5095,N_5003);
xnor U5215 (N_5215,N_5064,N_5020);
and U5216 (N_5216,N_5047,N_4998);
nor U5217 (N_5217,N_5082,N_4968);
or U5218 (N_5218,N_4968,N_5036);
or U5219 (N_5219,N_5088,N_5043);
xor U5220 (N_5220,N_4970,N_5044);
and U5221 (N_5221,N_4978,N_5048);
nand U5222 (N_5222,N_5064,N_5039);
xnor U5223 (N_5223,N_5088,N_5117);
or U5224 (N_5224,N_4972,N_5025);
or U5225 (N_5225,N_5096,N_4977);
and U5226 (N_5226,N_4964,N_4984);
nand U5227 (N_5227,N_4985,N_4995);
or U5228 (N_5228,N_5057,N_5117);
nor U5229 (N_5229,N_5007,N_5042);
and U5230 (N_5230,N_5018,N_4982);
nand U5231 (N_5231,N_5048,N_5040);
nand U5232 (N_5232,N_4967,N_5001);
nor U5233 (N_5233,N_5075,N_5033);
xnor U5234 (N_5234,N_4989,N_5103);
xnor U5235 (N_5235,N_5095,N_5097);
nor U5236 (N_5236,N_5007,N_5096);
or U5237 (N_5237,N_5029,N_5057);
nor U5238 (N_5238,N_5020,N_5085);
or U5239 (N_5239,N_4967,N_5028);
nand U5240 (N_5240,N_5101,N_4969);
nand U5241 (N_5241,N_5054,N_5035);
nor U5242 (N_5242,N_5110,N_4966);
or U5243 (N_5243,N_5062,N_4972);
nor U5244 (N_5244,N_5018,N_5042);
or U5245 (N_5245,N_5015,N_5045);
nand U5246 (N_5246,N_5031,N_5014);
xnor U5247 (N_5247,N_5060,N_5090);
nor U5248 (N_5248,N_4968,N_5051);
nand U5249 (N_5249,N_5046,N_5110);
or U5250 (N_5250,N_5115,N_5101);
or U5251 (N_5251,N_5102,N_5030);
xnor U5252 (N_5252,N_5118,N_4967);
nor U5253 (N_5253,N_5056,N_4969);
and U5254 (N_5254,N_5106,N_5075);
nor U5255 (N_5255,N_5078,N_5094);
xnor U5256 (N_5256,N_5065,N_5072);
nand U5257 (N_5257,N_5112,N_4970);
or U5258 (N_5258,N_4977,N_4976);
nand U5259 (N_5259,N_5104,N_5097);
or U5260 (N_5260,N_5062,N_5058);
nand U5261 (N_5261,N_4986,N_4967);
xnor U5262 (N_5262,N_5047,N_5028);
nand U5263 (N_5263,N_5056,N_4993);
and U5264 (N_5264,N_5094,N_5087);
xor U5265 (N_5265,N_5060,N_4970);
and U5266 (N_5266,N_5105,N_4969);
and U5267 (N_5267,N_4989,N_4965);
nand U5268 (N_5268,N_4968,N_5103);
xor U5269 (N_5269,N_5023,N_5115);
xor U5270 (N_5270,N_4971,N_4986);
nor U5271 (N_5271,N_5032,N_5021);
xor U5272 (N_5272,N_5073,N_4976);
nor U5273 (N_5273,N_5019,N_4997);
or U5274 (N_5274,N_5099,N_5026);
or U5275 (N_5275,N_5059,N_5023);
nand U5276 (N_5276,N_5107,N_5003);
or U5277 (N_5277,N_5111,N_4976);
and U5278 (N_5278,N_5029,N_5117);
xnor U5279 (N_5279,N_4965,N_5013);
and U5280 (N_5280,N_5148,N_5272);
nor U5281 (N_5281,N_5248,N_5277);
nand U5282 (N_5282,N_5208,N_5215);
xnor U5283 (N_5283,N_5226,N_5163);
or U5284 (N_5284,N_5120,N_5278);
nand U5285 (N_5285,N_5271,N_5142);
or U5286 (N_5286,N_5157,N_5188);
nor U5287 (N_5287,N_5230,N_5177);
xor U5288 (N_5288,N_5179,N_5165);
xor U5289 (N_5289,N_5256,N_5241);
nand U5290 (N_5290,N_5210,N_5178);
and U5291 (N_5291,N_5199,N_5161);
xor U5292 (N_5292,N_5133,N_5267);
and U5293 (N_5293,N_5218,N_5192);
xnor U5294 (N_5294,N_5213,N_5202);
nor U5295 (N_5295,N_5227,N_5275);
nor U5296 (N_5296,N_5261,N_5198);
xor U5297 (N_5297,N_5242,N_5222);
and U5298 (N_5298,N_5138,N_5122);
nand U5299 (N_5299,N_5257,N_5173);
and U5300 (N_5300,N_5187,N_5209);
and U5301 (N_5301,N_5132,N_5180);
or U5302 (N_5302,N_5212,N_5244);
xnor U5303 (N_5303,N_5124,N_5128);
nand U5304 (N_5304,N_5200,N_5146);
and U5305 (N_5305,N_5139,N_5154);
nand U5306 (N_5306,N_5254,N_5259);
and U5307 (N_5307,N_5220,N_5166);
nand U5308 (N_5308,N_5264,N_5206);
nor U5309 (N_5309,N_5262,N_5247);
nor U5310 (N_5310,N_5172,N_5145);
nand U5311 (N_5311,N_5135,N_5214);
and U5312 (N_5312,N_5223,N_5234);
and U5313 (N_5313,N_5194,N_5169);
and U5314 (N_5314,N_5253,N_5201);
xor U5315 (N_5315,N_5228,N_5164);
or U5316 (N_5316,N_5246,N_5204);
nand U5317 (N_5317,N_5252,N_5134);
xnor U5318 (N_5318,N_5184,N_5183);
nor U5319 (N_5319,N_5159,N_5121);
or U5320 (N_5320,N_5123,N_5224);
xor U5321 (N_5321,N_5266,N_5229);
nand U5322 (N_5322,N_5258,N_5176);
or U5323 (N_5323,N_5125,N_5182);
and U5324 (N_5324,N_5189,N_5131);
nor U5325 (N_5325,N_5197,N_5150);
nand U5326 (N_5326,N_5160,N_5207);
and U5327 (N_5327,N_5263,N_5250);
nand U5328 (N_5328,N_5130,N_5269);
or U5329 (N_5329,N_5153,N_5185);
nand U5330 (N_5330,N_5129,N_5219);
xnor U5331 (N_5331,N_5233,N_5195);
and U5332 (N_5332,N_5221,N_5136);
and U5333 (N_5333,N_5270,N_5143);
and U5334 (N_5334,N_5274,N_5151);
and U5335 (N_5335,N_5147,N_5255);
or U5336 (N_5336,N_5175,N_5260);
xnor U5337 (N_5337,N_5186,N_5190);
nor U5338 (N_5338,N_5170,N_5240);
or U5339 (N_5339,N_5162,N_5239);
nand U5340 (N_5340,N_5144,N_5171);
nor U5341 (N_5341,N_5141,N_5268);
or U5342 (N_5342,N_5237,N_5235);
or U5343 (N_5343,N_5152,N_5174);
nand U5344 (N_5344,N_5276,N_5205);
nor U5345 (N_5345,N_5127,N_5191);
xnor U5346 (N_5346,N_5243,N_5273);
xnor U5347 (N_5347,N_5193,N_5137);
and U5348 (N_5348,N_5249,N_5149);
nand U5349 (N_5349,N_5265,N_5211);
nor U5350 (N_5350,N_5251,N_5238);
or U5351 (N_5351,N_5217,N_5203);
or U5352 (N_5352,N_5167,N_5225);
xnor U5353 (N_5353,N_5232,N_5126);
nand U5354 (N_5354,N_5181,N_5216);
xor U5355 (N_5355,N_5140,N_5158);
nand U5356 (N_5356,N_5156,N_5279);
nor U5357 (N_5357,N_5155,N_5168);
or U5358 (N_5358,N_5196,N_5245);
nor U5359 (N_5359,N_5231,N_5236);
nand U5360 (N_5360,N_5138,N_5275);
or U5361 (N_5361,N_5229,N_5210);
or U5362 (N_5362,N_5191,N_5192);
xnor U5363 (N_5363,N_5188,N_5273);
or U5364 (N_5364,N_5166,N_5170);
nand U5365 (N_5365,N_5149,N_5222);
nor U5366 (N_5366,N_5170,N_5122);
nor U5367 (N_5367,N_5185,N_5120);
or U5368 (N_5368,N_5235,N_5274);
and U5369 (N_5369,N_5128,N_5144);
and U5370 (N_5370,N_5249,N_5152);
xnor U5371 (N_5371,N_5214,N_5208);
and U5372 (N_5372,N_5173,N_5150);
xnor U5373 (N_5373,N_5263,N_5157);
nand U5374 (N_5374,N_5146,N_5191);
and U5375 (N_5375,N_5212,N_5233);
nor U5376 (N_5376,N_5120,N_5258);
nand U5377 (N_5377,N_5271,N_5130);
nand U5378 (N_5378,N_5232,N_5226);
and U5379 (N_5379,N_5264,N_5201);
and U5380 (N_5380,N_5124,N_5161);
and U5381 (N_5381,N_5166,N_5173);
nand U5382 (N_5382,N_5218,N_5185);
nor U5383 (N_5383,N_5145,N_5258);
nor U5384 (N_5384,N_5267,N_5123);
xor U5385 (N_5385,N_5168,N_5183);
and U5386 (N_5386,N_5157,N_5140);
xor U5387 (N_5387,N_5204,N_5199);
or U5388 (N_5388,N_5150,N_5198);
and U5389 (N_5389,N_5169,N_5173);
xor U5390 (N_5390,N_5145,N_5271);
xnor U5391 (N_5391,N_5162,N_5179);
and U5392 (N_5392,N_5254,N_5149);
nand U5393 (N_5393,N_5130,N_5170);
nand U5394 (N_5394,N_5173,N_5187);
nor U5395 (N_5395,N_5253,N_5149);
xor U5396 (N_5396,N_5144,N_5273);
nor U5397 (N_5397,N_5265,N_5177);
xnor U5398 (N_5398,N_5185,N_5205);
or U5399 (N_5399,N_5137,N_5179);
nor U5400 (N_5400,N_5144,N_5254);
xnor U5401 (N_5401,N_5135,N_5248);
xor U5402 (N_5402,N_5155,N_5205);
xor U5403 (N_5403,N_5270,N_5202);
nor U5404 (N_5404,N_5256,N_5191);
and U5405 (N_5405,N_5261,N_5275);
or U5406 (N_5406,N_5270,N_5218);
nor U5407 (N_5407,N_5275,N_5125);
xor U5408 (N_5408,N_5172,N_5180);
nor U5409 (N_5409,N_5261,N_5129);
nor U5410 (N_5410,N_5227,N_5148);
nor U5411 (N_5411,N_5185,N_5170);
and U5412 (N_5412,N_5210,N_5238);
nor U5413 (N_5413,N_5218,N_5251);
xnor U5414 (N_5414,N_5248,N_5134);
or U5415 (N_5415,N_5158,N_5168);
nand U5416 (N_5416,N_5227,N_5179);
nand U5417 (N_5417,N_5249,N_5141);
nor U5418 (N_5418,N_5126,N_5260);
or U5419 (N_5419,N_5183,N_5154);
xor U5420 (N_5420,N_5142,N_5274);
or U5421 (N_5421,N_5244,N_5140);
or U5422 (N_5422,N_5188,N_5150);
and U5423 (N_5423,N_5132,N_5231);
nand U5424 (N_5424,N_5219,N_5167);
nand U5425 (N_5425,N_5160,N_5150);
nand U5426 (N_5426,N_5252,N_5256);
nand U5427 (N_5427,N_5143,N_5179);
or U5428 (N_5428,N_5256,N_5155);
nand U5429 (N_5429,N_5197,N_5144);
nand U5430 (N_5430,N_5134,N_5148);
xnor U5431 (N_5431,N_5127,N_5250);
xor U5432 (N_5432,N_5201,N_5182);
or U5433 (N_5433,N_5233,N_5258);
nand U5434 (N_5434,N_5153,N_5251);
and U5435 (N_5435,N_5146,N_5156);
nand U5436 (N_5436,N_5248,N_5200);
xor U5437 (N_5437,N_5211,N_5171);
nor U5438 (N_5438,N_5217,N_5169);
and U5439 (N_5439,N_5151,N_5153);
nor U5440 (N_5440,N_5435,N_5352);
nor U5441 (N_5441,N_5312,N_5382);
or U5442 (N_5442,N_5400,N_5353);
and U5443 (N_5443,N_5367,N_5315);
and U5444 (N_5444,N_5329,N_5281);
xnor U5445 (N_5445,N_5334,N_5320);
nand U5446 (N_5446,N_5330,N_5337);
or U5447 (N_5447,N_5380,N_5335);
or U5448 (N_5448,N_5328,N_5339);
and U5449 (N_5449,N_5381,N_5363);
and U5450 (N_5450,N_5387,N_5433);
xnor U5451 (N_5451,N_5421,N_5338);
nand U5452 (N_5452,N_5344,N_5431);
nand U5453 (N_5453,N_5358,N_5345);
nand U5454 (N_5454,N_5341,N_5299);
and U5455 (N_5455,N_5415,N_5384);
xor U5456 (N_5456,N_5340,N_5401);
xor U5457 (N_5457,N_5437,N_5294);
nand U5458 (N_5458,N_5280,N_5404);
or U5459 (N_5459,N_5418,N_5297);
and U5460 (N_5460,N_5306,N_5365);
nor U5461 (N_5461,N_5402,N_5285);
or U5462 (N_5462,N_5322,N_5364);
nand U5463 (N_5463,N_5287,N_5290);
or U5464 (N_5464,N_5347,N_5346);
xor U5465 (N_5465,N_5430,N_5385);
or U5466 (N_5466,N_5313,N_5283);
nand U5467 (N_5467,N_5325,N_5432);
nor U5468 (N_5468,N_5286,N_5439);
or U5469 (N_5469,N_5410,N_5311);
nand U5470 (N_5470,N_5407,N_5296);
nor U5471 (N_5471,N_5414,N_5291);
xnor U5472 (N_5472,N_5428,N_5323);
and U5473 (N_5473,N_5303,N_5282);
nor U5474 (N_5474,N_5292,N_5429);
or U5475 (N_5475,N_5343,N_5289);
or U5476 (N_5476,N_5436,N_5307);
or U5477 (N_5477,N_5390,N_5373);
nor U5478 (N_5478,N_5359,N_5305);
nand U5479 (N_5479,N_5394,N_5354);
nor U5480 (N_5480,N_5378,N_5420);
nor U5481 (N_5481,N_5379,N_5350);
or U5482 (N_5482,N_5369,N_5293);
and U5483 (N_5483,N_5308,N_5403);
xor U5484 (N_5484,N_5406,N_5309);
nor U5485 (N_5485,N_5409,N_5424);
xor U5486 (N_5486,N_5361,N_5408);
nand U5487 (N_5487,N_5371,N_5349);
nor U5488 (N_5488,N_5304,N_5356);
nor U5489 (N_5489,N_5405,N_5368);
or U5490 (N_5490,N_5366,N_5422);
or U5491 (N_5491,N_5362,N_5351);
or U5492 (N_5492,N_5393,N_5426);
nand U5493 (N_5493,N_5427,N_5417);
or U5494 (N_5494,N_5288,N_5327);
and U5495 (N_5495,N_5333,N_5372);
nor U5496 (N_5496,N_5316,N_5310);
xor U5497 (N_5497,N_5412,N_5397);
nor U5498 (N_5498,N_5355,N_5317);
and U5499 (N_5499,N_5391,N_5331);
xor U5500 (N_5500,N_5318,N_5419);
or U5501 (N_5501,N_5321,N_5388);
or U5502 (N_5502,N_5301,N_5398);
nand U5503 (N_5503,N_5438,N_5336);
nor U5504 (N_5504,N_5298,N_5375);
or U5505 (N_5505,N_5425,N_5302);
nor U5506 (N_5506,N_5360,N_5295);
and U5507 (N_5507,N_5314,N_5376);
nor U5508 (N_5508,N_5332,N_5348);
nand U5509 (N_5509,N_5399,N_5324);
or U5510 (N_5510,N_5413,N_5357);
nor U5511 (N_5511,N_5392,N_5383);
and U5512 (N_5512,N_5374,N_5395);
nor U5513 (N_5513,N_5423,N_5386);
and U5514 (N_5514,N_5300,N_5342);
and U5515 (N_5515,N_5319,N_5411);
or U5516 (N_5516,N_5389,N_5396);
nand U5517 (N_5517,N_5416,N_5434);
nor U5518 (N_5518,N_5326,N_5370);
or U5519 (N_5519,N_5284,N_5377);
or U5520 (N_5520,N_5417,N_5369);
or U5521 (N_5521,N_5299,N_5374);
nor U5522 (N_5522,N_5345,N_5319);
or U5523 (N_5523,N_5353,N_5377);
nand U5524 (N_5524,N_5324,N_5311);
and U5525 (N_5525,N_5287,N_5294);
nor U5526 (N_5526,N_5410,N_5343);
xnor U5527 (N_5527,N_5351,N_5422);
xor U5528 (N_5528,N_5324,N_5427);
nand U5529 (N_5529,N_5313,N_5370);
and U5530 (N_5530,N_5322,N_5409);
or U5531 (N_5531,N_5338,N_5344);
nor U5532 (N_5532,N_5327,N_5294);
nor U5533 (N_5533,N_5410,N_5438);
or U5534 (N_5534,N_5337,N_5339);
nand U5535 (N_5535,N_5377,N_5335);
nand U5536 (N_5536,N_5339,N_5296);
and U5537 (N_5537,N_5431,N_5361);
nor U5538 (N_5538,N_5292,N_5321);
or U5539 (N_5539,N_5432,N_5319);
and U5540 (N_5540,N_5299,N_5305);
xnor U5541 (N_5541,N_5377,N_5379);
xnor U5542 (N_5542,N_5403,N_5376);
nor U5543 (N_5543,N_5317,N_5387);
xor U5544 (N_5544,N_5309,N_5331);
and U5545 (N_5545,N_5314,N_5291);
nand U5546 (N_5546,N_5337,N_5297);
or U5547 (N_5547,N_5420,N_5363);
nand U5548 (N_5548,N_5328,N_5426);
or U5549 (N_5549,N_5364,N_5320);
nand U5550 (N_5550,N_5319,N_5416);
or U5551 (N_5551,N_5395,N_5328);
xnor U5552 (N_5552,N_5380,N_5311);
nand U5553 (N_5553,N_5351,N_5326);
and U5554 (N_5554,N_5345,N_5380);
nor U5555 (N_5555,N_5327,N_5423);
nand U5556 (N_5556,N_5426,N_5383);
xor U5557 (N_5557,N_5376,N_5431);
nand U5558 (N_5558,N_5298,N_5396);
nor U5559 (N_5559,N_5381,N_5434);
nand U5560 (N_5560,N_5411,N_5308);
xor U5561 (N_5561,N_5418,N_5428);
xnor U5562 (N_5562,N_5371,N_5411);
and U5563 (N_5563,N_5420,N_5288);
and U5564 (N_5564,N_5418,N_5292);
or U5565 (N_5565,N_5422,N_5344);
xor U5566 (N_5566,N_5327,N_5332);
or U5567 (N_5567,N_5316,N_5285);
and U5568 (N_5568,N_5283,N_5430);
nor U5569 (N_5569,N_5358,N_5371);
and U5570 (N_5570,N_5306,N_5397);
nand U5571 (N_5571,N_5403,N_5397);
nor U5572 (N_5572,N_5309,N_5417);
and U5573 (N_5573,N_5430,N_5346);
xnor U5574 (N_5574,N_5346,N_5401);
xor U5575 (N_5575,N_5430,N_5371);
xor U5576 (N_5576,N_5315,N_5382);
xnor U5577 (N_5577,N_5387,N_5319);
nand U5578 (N_5578,N_5402,N_5366);
nor U5579 (N_5579,N_5397,N_5361);
or U5580 (N_5580,N_5300,N_5328);
nand U5581 (N_5581,N_5328,N_5286);
xor U5582 (N_5582,N_5362,N_5313);
or U5583 (N_5583,N_5425,N_5393);
nand U5584 (N_5584,N_5410,N_5368);
nand U5585 (N_5585,N_5301,N_5321);
or U5586 (N_5586,N_5391,N_5369);
nor U5587 (N_5587,N_5307,N_5395);
or U5588 (N_5588,N_5383,N_5386);
nor U5589 (N_5589,N_5372,N_5285);
nor U5590 (N_5590,N_5380,N_5352);
xnor U5591 (N_5591,N_5411,N_5374);
and U5592 (N_5592,N_5340,N_5297);
nor U5593 (N_5593,N_5399,N_5435);
nand U5594 (N_5594,N_5344,N_5307);
and U5595 (N_5595,N_5290,N_5368);
or U5596 (N_5596,N_5319,N_5378);
nand U5597 (N_5597,N_5402,N_5363);
and U5598 (N_5598,N_5379,N_5365);
nand U5599 (N_5599,N_5366,N_5323);
and U5600 (N_5600,N_5484,N_5465);
xor U5601 (N_5601,N_5493,N_5504);
or U5602 (N_5602,N_5468,N_5511);
or U5603 (N_5603,N_5446,N_5521);
and U5604 (N_5604,N_5597,N_5578);
nand U5605 (N_5605,N_5515,N_5585);
and U5606 (N_5606,N_5588,N_5523);
nor U5607 (N_5607,N_5575,N_5576);
nand U5608 (N_5608,N_5563,N_5461);
nand U5609 (N_5609,N_5564,N_5481);
xor U5610 (N_5610,N_5551,N_5544);
and U5611 (N_5611,N_5556,N_5463);
and U5612 (N_5612,N_5513,N_5547);
and U5613 (N_5613,N_5571,N_5441);
nor U5614 (N_5614,N_5561,N_5459);
or U5615 (N_5615,N_5462,N_5533);
or U5616 (N_5616,N_5454,N_5443);
or U5617 (N_5617,N_5500,N_5593);
or U5618 (N_5618,N_5577,N_5573);
or U5619 (N_5619,N_5501,N_5472);
nand U5620 (N_5620,N_5505,N_5557);
nand U5621 (N_5621,N_5506,N_5509);
nor U5622 (N_5622,N_5540,N_5476);
nand U5623 (N_5623,N_5485,N_5589);
or U5624 (N_5624,N_5594,N_5494);
or U5625 (N_5625,N_5448,N_5497);
nand U5626 (N_5626,N_5545,N_5542);
nand U5627 (N_5627,N_5442,N_5479);
xnor U5628 (N_5628,N_5455,N_5487);
or U5629 (N_5629,N_5517,N_5591);
xnor U5630 (N_5630,N_5525,N_5586);
or U5631 (N_5631,N_5567,N_5580);
nor U5632 (N_5632,N_5512,N_5480);
nor U5633 (N_5633,N_5581,N_5469);
xor U5634 (N_5634,N_5473,N_5503);
nor U5635 (N_5635,N_5458,N_5535);
nand U5636 (N_5636,N_5452,N_5555);
nor U5637 (N_5637,N_5596,N_5447);
xor U5638 (N_5638,N_5543,N_5530);
and U5639 (N_5639,N_5536,N_5518);
and U5640 (N_5640,N_5519,N_5550);
nor U5641 (N_5641,N_5534,N_5532);
or U5642 (N_5642,N_5456,N_5531);
nor U5643 (N_5643,N_5548,N_5552);
xor U5644 (N_5644,N_5520,N_5507);
nand U5645 (N_5645,N_5527,N_5491);
and U5646 (N_5646,N_5558,N_5477);
and U5647 (N_5647,N_5508,N_5599);
and U5648 (N_5648,N_5470,N_5526);
nor U5649 (N_5649,N_5592,N_5549);
and U5650 (N_5650,N_5554,N_5475);
or U5651 (N_5651,N_5489,N_5574);
nor U5652 (N_5652,N_5565,N_5474);
and U5653 (N_5653,N_5502,N_5460);
nor U5654 (N_5654,N_5492,N_5449);
nor U5655 (N_5655,N_5464,N_5546);
or U5656 (N_5656,N_5450,N_5496);
nor U5657 (N_5657,N_5583,N_5566);
nor U5658 (N_5658,N_5582,N_5529);
nor U5659 (N_5659,N_5524,N_5483);
xor U5660 (N_5660,N_5587,N_5444);
nand U5661 (N_5661,N_5498,N_5539);
xor U5662 (N_5662,N_5490,N_5569);
and U5663 (N_5663,N_5579,N_5553);
nand U5664 (N_5664,N_5595,N_5560);
xnor U5665 (N_5665,N_5445,N_5538);
nand U5666 (N_5666,N_5453,N_5570);
nor U5667 (N_5667,N_5528,N_5451);
nor U5668 (N_5668,N_5510,N_5499);
xnor U5669 (N_5669,N_5572,N_5568);
nor U5670 (N_5670,N_5516,N_5467);
nor U5671 (N_5671,N_5541,N_5537);
nand U5672 (N_5672,N_5488,N_5466);
nor U5673 (N_5673,N_5590,N_5522);
and U5674 (N_5674,N_5471,N_5514);
or U5675 (N_5675,N_5598,N_5486);
or U5676 (N_5676,N_5440,N_5562);
xor U5677 (N_5677,N_5482,N_5584);
nand U5678 (N_5678,N_5457,N_5478);
xnor U5679 (N_5679,N_5495,N_5559);
nor U5680 (N_5680,N_5597,N_5564);
or U5681 (N_5681,N_5545,N_5551);
or U5682 (N_5682,N_5465,N_5453);
and U5683 (N_5683,N_5513,N_5481);
or U5684 (N_5684,N_5487,N_5480);
nand U5685 (N_5685,N_5526,N_5577);
and U5686 (N_5686,N_5448,N_5485);
and U5687 (N_5687,N_5588,N_5548);
or U5688 (N_5688,N_5598,N_5485);
xor U5689 (N_5689,N_5472,N_5592);
nor U5690 (N_5690,N_5479,N_5582);
xnor U5691 (N_5691,N_5590,N_5520);
nand U5692 (N_5692,N_5505,N_5507);
nand U5693 (N_5693,N_5487,N_5570);
and U5694 (N_5694,N_5493,N_5564);
nand U5695 (N_5695,N_5504,N_5537);
xnor U5696 (N_5696,N_5578,N_5507);
and U5697 (N_5697,N_5483,N_5442);
or U5698 (N_5698,N_5576,N_5545);
nand U5699 (N_5699,N_5586,N_5560);
or U5700 (N_5700,N_5591,N_5560);
or U5701 (N_5701,N_5513,N_5506);
nor U5702 (N_5702,N_5491,N_5464);
xor U5703 (N_5703,N_5521,N_5477);
xnor U5704 (N_5704,N_5501,N_5449);
nand U5705 (N_5705,N_5499,N_5554);
and U5706 (N_5706,N_5554,N_5483);
xor U5707 (N_5707,N_5446,N_5513);
or U5708 (N_5708,N_5573,N_5502);
and U5709 (N_5709,N_5541,N_5449);
xor U5710 (N_5710,N_5547,N_5509);
nor U5711 (N_5711,N_5508,N_5452);
nand U5712 (N_5712,N_5442,N_5481);
nand U5713 (N_5713,N_5597,N_5550);
xnor U5714 (N_5714,N_5565,N_5562);
nor U5715 (N_5715,N_5580,N_5508);
nand U5716 (N_5716,N_5453,N_5519);
or U5717 (N_5717,N_5548,N_5497);
xor U5718 (N_5718,N_5467,N_5578);
xor U5719 (N_5719,N_5480,N_5554);
or U5720 (N_5720,N_5578,N_5447);
nor U5721 (N_5721,N_5485,N_5593);
and U5722 (N_5722,N_5509,N_5581);
or U5723 (N_5723,N_5531,N_5540);
or U5724 (N_5724,N_5489,N_5550);
nor U5725 (N_5725,N_5594,N_5531);
nor U5726 (N_5726,N_5533,N_5547);
nor U5727 (N_5727,N_5487,N_5495);
nor U5728 (N_5728,N_5530,N_5497);
or U5729 (N_5729,N_5569,N_5487);
and U5730 (N_5730,N_5475,N_5587);
or U5731 (N_5731,N_5468,N_5530);
nor U5732 (N_5732,N_5440,N_5475);
or U5733 (N_5733,N_5572,N_5537);
nand U5734 (N_5734,N_5475,N_5503);
or U5735 (N_5735,N_5507,N_5538);
and U5736 (N_5736,N_5490,N_5579);
or U5737 (N_5737,N_5472,N_5467);
xor U5738 (N_5738,N_5451,N_5542);
nand U5739 (N_5739,N_5492,N_5524);
and U5740 (N_5740,N_5474,N_5533);
and U5741 (N_5741,N_5584,N_5529);
xor U5742 (N_5742,N_5591,N_5559);
nor U5743 (N_5743,N_5529,N_5448);
or U5744 (N_5744,N_5456,N_5567);
and U5745 (N_5745,N_5594,N_5518);
xnor U5746 (N_5746,N_5450,N_5571);
or U5747 (N_5747,N_5481,N_5521);
nand U5748 (N_5748,N_5555,N_5502);
nor U5749 (N_5749,N_5591,N_5495);
nor U5750 (N_5750,N_5599,N_5554);
nor U5751 (N_5751,N_5519,N_5462);
xnor U5752 (N_5752,N_5535,N_5517);
or U5753 (N_5753,N_5441,N_5516);
xor U5754 (N_5754,N_5543,N_5548);
xnor U5755 (N_5755,N_5521,N_5522);
xnor U5756 (N_5756,N_5495,N_5506);
nand U5757 (N_5757,N_5564,N_5558);
nor U5758 (N_5758,N_5455,N_5581);
nand U5759 (N_5759,N_5486,N_5479);
or U5760 (N_5760,N_5725,N_5685);
xor U5761 (N_5761,N_5635,N_5683);
or U5762 (N_5762,N_5653,N_5732);
nand U5763 (N_5763,N_5728,N_5707);
nor U5764 (N_5764,N_5745,N_5604);
nand U5765 (N_5765,N_5729,N_5715);
nand U5766 (N_5766,N_5724,N_5716);
and U5767 (N_5767,N_5608,N_5610);
nand U5768 (N_5768,N_5709,N_5670);
and U5769 (N_5769,N_5684,N_5679);
xor U5770 (N_5770,N_5634,N_5677);
xnor U5771 (N_5771,N_5721,N_5696);
xor U5772 (N_5772,N_5730,N_5713);
or U5773 (N_5773,N_5609,N_5743);
xor U5774 (N_5774,N_5629,N_5620);
and U5775 (N_5775,N_5739,N_5733);
or U5776 (N_5776,N_5686,N_5742);
or U5777 (N_5777,N_5680,N_5611);
nor U5778 (N_5778,N_5752,N_5669);
xnor U5779 (N_5779,N_5655,N_5665);
nand U5780 (N_5780,N_5623,N_5744);
xnor U5781 (N_5781,N_5642,N_5741);
nor U5782 (N_5782,N_5627,N_5628);
xnor U5783 (N_5783,N_5706,N_5617);
and U5784 (N_5784,N_5636,N_5632);
or U5785 (N_5785,N_5692,N_5671);
or U5786 (N_5786,N_5754,N_5690);
and U5787 (N_5787,N_5626,N_5606);
nand U5788 (N_5788,N_5693,N_5641);
nor U5789 (N_5789,N_5666,N_5664);
or U5790 (N_5790,N_5613,N_5746);
or U5791 (N_5791,N_5631,N_5735);
and U5792 (N_5792,N_5698,N_5749);
or U5793 (N_5793,N_5656,N_5649);
nand U5794 (N_5794,N_5748,N_5633);
nor U5795 (N_5795,N_5645,N_5672);
nand U5796 (N_5796,N_5704,N_5740);
or U5797 (N_5797,N_5614,N_5647);
and U5798 (N_5798,N_5619,N_5702);
nor U5799 (N_5799,N_5694,N_5750);
nor U5800 (N_5800,N_5691,N_5711);
xnor U5801 (N_5801,N_5757,N_5624);
or U5802 (N_5802,N_5687,N_5755);
nor U5803 (N_5803,N_5726,N_5618);
nand U5804 (N_5804,N_5637,N_5650);
and U5805 (N_5805,N_5737,N_5688);
or U5806 (N_5806,N_5731,N_5657);
nand U5807 (N_5807,N_5602,N_5605);
nor U5808 (N_5808,N_5612,N_5678);
nor U5809 (N_5809,N_5621,N_5630);
xor U5810 (N_5810,N_5663,N_5747);
nor U5811 (N_5811,N_5695,N_5753);
xor U5812 (N_5812,N_5660,N_5722);
nor U5813 (N_5813,N_5640,N_5699);
xnor U5814 (N_5814,N_5758,N_5654);
or U5815 (N_5815,N_5751,N_5700);
and U5816 (N_5816,N_5738,N_5600);
or U5817 (N_5817,N_5644,N_5718);
nand U5818 (N_5818,N_5734,N_5648);
xor U5819 (N_5819,N_5710,N_5736);
and U5820 (N_5820,N_5759,N_5651);
nand U5821 (N_5821,N_5607,N_5727);
nand U5822 (N_5822,N_5643,N_5689);
and U5823 (N_5823,N_5703,N_5659);
xnor U5824 (N_5824,N_5603,N_5662);
or U5825 (N_5825,N_5658,N_5616);
nor U5826 (N_5826,N_5682,N_5625);
nand U5827 (N_5827,N_5601,N_5674);
xnor U5828 (N_5828,N_5756,N_5717);
nand U5829 (N_5829,N_5646,N_5701);
nor U5830 (N_5830,N_5661,N_5705);
nor U5831 (N_5831,N_5720,N_5714);
xnor U5832 (N_5832,N_5719,N_5675);
xor U5833 (N_5833,N_5723,N_5676);
or U5834 (N_5834,N_5615,N_5622);
nand U5835 (N_5835,N_5668,N_5712);
xnor U5836 (N_5836,N_5697,N_5667);
and U5837 (N_5837,N_5652,N_5681);
xnor U5838 (N_5838,N_5638,N_5639);
or U5839 (N_5839,N_5708,N_5673);
xor U5840 (N_5840,N_5712,N_5699);
and U5841 (N_5841,N_5679,N_5731);
xnor U5842 (N_5842,N_5624,N_5644);
and U5843 (N_5843,N_5736,N_5624);
and U5844 (N_5844,N_5698,N_5680);
and U5845 (N_5845,N_5706,N_5675);
nand U5846 (N_5846,N_5720,N_5708);
nor U5847 (N_5847,N_5609,N_5600);
xor U5848 (N_5848,N_5669,N_5619);
nand U5849 (N_5849,N_5755,N_5669);
or U5850 (N_5850,N_5609,N_5683);
nand U5851 (N_5851,N_5678,N_5720);
nor U5852 (N_5852,N_5736,N_5614);
nor U5853 (N_5853,N_5693,N_5748);
or U5854 (N_5854,N_5644,N_5695);
nor U5855 (N_5855,N_5723,N_5635);
and U5856 (N_5856,N_5618,N_5688);
nand U5857 (N_5857,N_5672,N_5659);
or U5858 (N_5858,N_5655,N_5647);
and U5859 (N_5859,N_5629,N_5706);
and U5860 (N_5860,N_5728,N_5744);
nor U5861 (N_5861,N_5737,N_5668);
nor U5862 (N_5862,N_5607,N_5619);
or U5863 (N_5863,N_5726,N_5606);
nand U5864 (N_5864,N_5665,N_5602);
and U5865 (N_5865,N_5735,N_5730);
and U5866 (N_5866,N_5600,N_5684);
and U5867 (N_5867,N_5640,N_5701);
and U5868 (N_5868,N_5607,N_5646);
and U5869 (N_5869,N_5743,N_5621);
nor U5870 (N_5870,N_5608,N_5676);
and U5871 (N_5871,N_5739,N_5604);
nand U5872 (N_5872,N_5656,N_5727);
and U5873 (N_5873,N_5613,N_5610);
or U5874 (N_5874,N_5618,N_5622);
xnor U5875 (N_5875,N_5710,N_5687);
and U5876 (N_5876,N_5756,N_5667);
and U5877 (N_5877,N_5713,N_5719);
or U5878 (N_5878,N_5632,N_5622);
xor U5879 (N_5879,N_5718,N_5651);
xor U5880 (N_5880,N_5715,N_5700);
and U5881 (N_5881,N_5690,N_5609);
nand U5882 (N_5882,N_5731,N_5743);
and U5883 (N_5883,N_5692,N_5701);
or U5884 (N_5884,N_5624,N_5718);
nor U5885 (N_5885,N_5654,N_5643);
nor U5886 (N_5886,N_5740,N_5649);
and U5887 (N_5887,N_5608,N_5674);
nand U5888 (N_5888,N_5615,N_5706);
nor U5889 (N_5889,N_5668,N_5608);
nand U5890 (N_5890,N_5613,N_5712);
nor U5891 (N_5891,N_5602,N_5725);
nor U5892 (N_5892,N_5619,N_5723);
nor U5893 (N_5893,N_5728,N_5686);
xor U5894 (N_5894,N_5635,N_5707);
and U5895 (N_5895,N_5708,N_5700);
nand U5896 (N_5896,N_5691,N_5687);
nor U5897 (N_5897,N_5651,N_5606);
nor U5898 (N_5898,N_5673,N_5655);
or U5899 (N_5899,N_5661,N_5674);
or U5900 (N_5900,N_5677,N_5650);
xor U5901 (N_5901,N_5759,N_5745);
xor U5902 (N_5902,N_5707,N_5604);
and U5903 (N_5903,N_5726,N_5671);
or U5904 (N_5904,N_5663,N_5636);
nor U5905 (N_5905,N_5638,N_5614);
xor U5906 (N_5906,N_5732,N_5639);
nor U5907 (N_5907,N_5691,N_5681);
nor U5908 (N_5908,N_5708,N_5715);
nand U5909 (N_5909,N_5602,N_5684);
nor U5910 (N_5910,N_5608,N_5739);
nand U5911 (N_5911,N_5693,N_5686);
or U5912 (N_5912,N_5655,N_5658);
nand U5913 (N_5913,N_5647,N_5685);
nor U5914 (N_5914,N_5654,N_5722);
nand U5915 (N_5915,N_5680,N_5609);
nand U5916 (N_5916,N_5669,N_5625);
xor U5917 (N_5917,N_5703,N_5637);
nor U5918 (N_5918,N_5681,N_5712);
or U5919 (N_5919,N_5754,N_5678);
and U5920 (N_5920,N_5868,N_5891);
nand U5921 (N_5921,N_5794,N_5799);
nand U5922 (N_5922,N_5912,N_5863);
or U5923 (N_5923,N_5872,N_5904);
and U5924 (N_5924,N_5833,N_5903);
or U5925 (N_5925,N_5878,N_5839);
xor U5926 (N_5926,N_5781,N_5780);
and U5927 (N_5927,N_5814,N_5877);
nor U5928 (N_5928,N_5797,N_5854);
nand U5929 (N_5929,N_5834,N_5919);
or U5930 (N_5930,N_5767,N_5876);
nor U5931 (N_5931,N_5784,N_5793);
and U5932 (N_5932,N_5864,N_5860);
and U5933 (N_5933,N_5880,N_5769);
nor U5934 (N_5934,N_5875,N_5821);
nand U5935 (N_5935,N_5830,N_5853);
xor U5936 (N_5936,N_5867,N_5890);
and U5937 (N_5937,N_5847,N_5858);
nand U5938 (N_5938,N_5770,N_5832);
nor U5939 (N_5939,N_5851,N_5813);
nor U5940 (N_5940,N_5782,N_5888);
and U5941 (N_5941,N_5881,N_5911);
nor U5942 (N_5942,N_5862,N_5820);
nand U5943 (N_5943,N_5801,N_5789);
nand U5944 (N_5944,N_5764,N_5899);
nor U5945 (N_5945,N_5809,N_5776);
nor U5946 (N_5946,N_5802,N_5772);
xor U5947 (N_5947,N_5856,N_5783);
nor U5948 (N_5948,N_5791,N_5889);
or U5949 (N_5949,N_5822,N_5917);
nor U5950 (N_5950,N_5895,N_5805);
xor U5951 (N_5951,N_5913,N_5907);
or U5952 (N_5952,N_5779,N_5902);
xor U5953 (N_5953,N_5806,N_5892);
xor U5954 (N_5954,N_5788,N_5884);
nand U5955 (N_5955,N_5905,N_5798);
nand U5956 (N_5956,N_5855,N_5829);
xor U5957 (N_5957,N_5790,N_5827);
xor U5958 (N_5958,N_5819,N_5873);
nand U5959 (N_5959,N_5852,N_5909);
nand U5960 (N_5960,N_5894,N_5900);
nand U5961 (N_5961,N_5840,N_5774);
nand U5962 (N_5962,N_5850,N_5882);
and U5963 (N_5963,N_5844,N_5871);
nor U5964 (N_5964,N_5837,N_5896);
nor U5965 (N_5965,N_5804,N_5812);
nor U5966 (N_5966,N_5918,N_5762);
xnor U5967 (N_5967,N_5874,N_5796);
and U5968 (N_5968,N_5823,N_5810);
xor U5969 (N_5969,N_5828,N_5857);
or U5970 (N_5970,N_5897,N_5887);
nor U5971 (N_5971,N_5879,N_5778);
nand U5972 (N_5972,N_5777,N_5815);
and U5973 (N_5973,N_5775,N_5785);
nor U5974 (N_5974,N_5915,N_5845);
or U5975 (N_5975,N_5901,N_5787);
nand U5976 (N_5976,N_5766,N_5803);
or U5977 (N_5977,N_5825,N_5771);
nand U5978 (N_5978,N_5910,N_5893);
xnor U5979 (N_5979,N_5908,N_5898);
nor U5980 (N_5980,N_5886,N_5773);
and U5981 (N_5981,N_5786,N_5914);
and U5982 (N_5982,N_5836,N_5885);
xnor U5983 (N_5983,N_5870,N_5824);
nand U5984 (N_5984,N_5859,N_5768);
xor U5985 (N_5985,N_5841,N_5843);
nor U5986 (N_5986,N_5869,N_5861);
xnor U5987 (N_5987,N_5800,N_5842);
and U5988 (N_5988,N_5826,N_5846);
nor U5989 (N_5989,N_5916,N_5906);
and U5990 (N_5990,N_5838,N_5792);
or U5991 (N_5991,N_5849,N_5761);
nand U5992 (N_5992,N_5883,N_5866);
nand U5993 (N_5993,N_5816,N_5763);
nand U5994 (N_5994,N_5865,N_5817);
xor U5995 (N_5995,N_5831,N_5760);
or U5996 (N_5996,N_5808,N_5811);
xnor U5997 (N_5997,N_5848,N_5795);
or U5998 (N_5998,N_5818,N_5835);
or U5999 (N_5999,N_5807,N_5765);
nor U6000 (N_6000,N_5760,N_5868);
xor U6001 (N_6001,N_5913,N_5797);
xnor U6002 (N_6002,N_5852,N_5786);
or U6003 (N_6003,N_5891,N_5874);
or U6004 (N_6004,N_5814,N_5813);
and U6005 (N_6005,N_5880,N_5810);
and U6006 (N_6006,N_5822,N_5888);
nor U6007 (N_6007,N_5793,N_5892);
nor U6008 (N_6008,N_5775,N_5881);
and U6009 (N_6009,N_5830,N_5796);
nor U6010 (N_6010,N_5901,N_5902);
nor U6011 (N_6011,N_5818,N_5918);
and U6012 (N_6012,N_5834,N_5876);
and U6013 (N_6013,N_5819,N_5880);
or U6014 (N_6014,N_5780,N_5893);
nor U6015 (N_6015,N_5894,N_5799);
nor U6016 (N_6016,N_5786,N_5822);
and U6017 (N_6017,N_5816,N_5775);
xor U6018 (N_6018,N_5793,N_5788);
xnor U6019 (N_6019,N_5889,N_5786);
xor U6020 (N_6020,N_5766,N_5835);
xor U6021 (N_6021,N_5870,N_5887);
nor U6022 (N_6022,N_5860,N_5867);
nor U6023 (N_6023,N_5898,N_5808);
nand U6024 (N_6024,N_5903,N_5825);
and U6025 (N_6025,N_5918,N_5778);
xor U6026 (N_6026,N_5800,N_5872);
and U6027 (N_6027,N_5790,N_5777);
xnor U6028 (N_6028,N_5898,N_5802);
and U6029 (N_6029,N_5791,N_5918);
and U6030 (N_6030,N_5764,N_5870);
nand U6031 (N_6031,N_5798,N_5765);
or U6032 (N_6032,N_5841,N_5794);
nor U6033 (N_6033,N_5822,N_5800);
nand U6034 (N_6034,N_5810,N_5865);
or U6035 (N_6035,N_5775,N_5787);
nand U6036 (N_6036,N_5919,N_5855);
nor U6037 (N_6037,N_5796,N_5800);
xnor U6038 (N_6038,N_5915,N_5810);
nand U6039 (N_6039,N_5817,N_5792);
and U6040 (N_6040,N_5838,N_5797);
or U6041 (N_6041,N_5806,N_5918);
nor U6042 (N_6042,N_5893,N_5869);
or U6043 (N_6043,N_5869,N_5895);
and U6044 (N_6044,N_5849,N_5786);
or U6045 (N_6045,N_5860,N_5775);
or U6046 (N_6046,N_5875,N_5916);
or U6047 (N_6047,N_5854,N_5777);
or U6048 (N_6048,N_5839,N_5764);
and U6049 (N_6049,N_5791,N_5888);
xor U6050 (N_6050,N_5823,N_5767);
xnor U6051 (N_6051,N_5857,N_5909);
nand U6052 (N_6052,N_5770,N_5794);
xor U6053 (N_6053,N_5768,N_5916);
or U6054 (N_6054,N_5828,N_5872);
and U6055 (N_6055,N_5826,N_5847);
nor U6056 (N_6056,N_5915,N_5904);
xnor U6057 (N_6057,N_5780,N_5802);
xor U6058 (N_6058,N_5917,N_5826);
and U6059 (N_6059,N_5837,N_5795);
xor U6060 (N_6060,N_5897,N_5917);
nand U6061 (N_6061,N_5863,N_5898);
nor U6062 (N_6062,N_5788,N_5791);
nand U6063 (N_6063,N_5781,N_5909);
or U6064 (N_6064,N_5892,N_5770);
nor U6065 (N_6065,N_5903,N_5906);
and U6066 (N_6066,N_5900,N_5896);
and U6067 (N_6067,N_5792,N_5839);
or U6068 (N_6068,N_5760,N_5855);
nor U6069 (N_6069,N_5853,N_5880);
or U6070 (N_6070,N_5810,N_5877);
nor U6071 (N_6071,N_5905,N_5797);
or U6072 (N_6072,N_5832,N_5881);
and U6073 (N_6073,N_5890,N_5780);
or U6074 (N_6074,N_5834,N_5797);
or U6075 (N_6075,N_5859,N_5808);
nand U6076 (N_6076,N_5882,N_5871);
nand U6077 (N_6077,N_5806,N_5767);
nand U6078 (N_6078,N_5780,N_5794);
or U6079 (N_6079,N_5850,N_5819);
nand U6080 (N_6080,N_6074,N_6006);
or U6081 (N_6081,N_5944,N_6056);
xor U6082 (N_6082,N_5972,N_6061);
xor U6083 (N_6083,N_6028,N_5979);
and U6084 (N_6084,N_5971,N_5955);
and U6085 (N_6085,N_6001,N_6000);
nand U6086 (N_6086,N_5960,N_5969);
or U6087 (N_6087,N_5976,N_6063);
or U6088 (N_6088,N_6038,N_5941);
nor U6089 (N_6089,N_5929,N_6005);
and U6090 (N_6090,N_5964,N_5974);
xor U6091 (N_6091,N_6017,N_5952);
nand U6092 (N_6092,N_5966,N_6076);
xor U6093 (N_6093,N_5926,N_6071);
nand U6094 (N_6094,N_5998,N_6069);
nor U6095 (N_6095,N_6072,N_6058);
nor U6096 (N_6096,N_5993,N_6040);
xor U6097 (N_6097,N_6011,N_5936);
nor U6098 (N_6098,N_6019,N_5947);
or U6099 (N_6099,N_5996,N_5985);
nor U6100 (N_6100,N_6007,N_5942);
or U6101 (N_6101,N_5988,N_6016);
or U6102 (N_6102,N_5921,N_5967);
nand U6103 (N_6103,N_6012,N_6044);
or U6104 (N_6104,N_5968,N_6059);
nand U6105 (N_6105,N_5924,N_6025);
and U6106 (N_6106,N_6030,N_6041);
nand U6107 (N_6107,N_6047,N_6021);
nand U6108 (N_6108,N_6043,N_5932);
nor U6109 (N_6109,N_6004,N_5943);
or U6110 (N_6110,N_6008,N_5937);
xor U6111 (N_6111,N_6024,N_5928);
nand U6112 (N_6112,N_5982,N_5925);
nor U6113 (N_6113,N_5997,N_5946);
or U6114 (N_6114,N_5951,N_6050);
nand U6115 (N_6115,N_5975,N_5959);
nand U6116 (N_6116,N_6051,N_5953);
or U6117 (N_6117,N_5950,N_5938);
nor U6118 (N_6118,N_6026,N_5989);
nand U6119 (N_6119,N_6033,N_6075);
or U6120 (N_6120,N_6067,N_6077);
xnor U6121 (N_6121,N_5984,N_6068);
or U6122 (N_6122,N_5931,N_6010);
nand U6123 (N_6123,N_6064,N_6032);
and U6124 (N_6124,N_5954,N_5940);
nand U6125 (N_6125,N_6048,N_6039);
xor U6126 (N_6126,N_5927,N_6018);
or U6127 (N_6127,N_5962,N_6002);
nand U6128 (N_6128,N_5961,N_6065);
nand U6129 (N_6129,N_5987,N_5994);
xnor U6130 (N_6130,N_5999,N_6060);
and U6131 (N_6131,N_5973,N_5935);
and U6132 (N_6132,N_6029,N_6027);
nor U6133 (N_6133,N_5991,N_5990);
nor U6134 (N_6134,N_5980,N_5948);
xor U6135 (N_6135,N_6022,N_5983);
or U6136 (N_6136,N_5963,N_6053);
or U6137 (N_6137,N_5986,N_5920);
xnor U6138 (N_6138,N_5958,N_6009);
nor U6139 (N_6139,N_5945,N_5957);
or U6140 (N_6140,N_5965,N_6045);
nand U6141 (N_6141,N_6013,N_6062);
and U6142 (N_6142,N_5956,N_6055);
nor U6143 (N_6143,N_5949,N_5922);
xnor U6144 (N_6144,N_5981,N_6037);
xnor U6145 (N_6145,N_6073,N_5934);
nand U6146 (N_6146,N_6057,N_6054);
or U6147 (N_6147,N_5978,N_6031);
and U6148 (N_6148,N_6003,N_6015);
nor U6149 (N_6149,N_6014,N_6049);
xor U6150 (N_6150,N_6078,N_6066);
nor U6151 (N_6151,N_5992,N_6020);
and U6152 (N_6152,N_5933,N_5970);
nand U6153 (N_6153,N_6042,N_5930);
xor U6154 (N_6154,N_6035,N_6034);
nor U6155 (N_6155,N_5995,N_5939);
nand U6156 (N_6156,N_6036,N_6046);
or U6157 (N_6157,N_6070,N_5977);
or U6158 (N_6158,N_6023,N_6052);
nor U6159 (N_6159,N_6079,N_5923);
xor U6160 (N_6160,N_5965,N_6077);
nand U6161 (N_6161,N_5957,N_6027);
nor U6162 (N_6162,N_6025,N_6008);
and U6163 (N_6163,N_5946,N_6076);
xor U6164 (N_6164,N_6051,N_5937);
or U6165 (N_6165,N_6020,N_5973);
nor U6166 (N_6166,N_5956,N_5972);
nor U6167 (N_6167,N_6028,N_5971);
nand U6168 (N_6168,N_5971,N_5926);
or U6169 (N_6169,N_6045,N_5937);
nand U6170 (N_6170,N_5925,N_6062);
nor U6171 (N_6171,N_5990,N_5982);
xor U6172 (N_6172,N_6015,N_6002);
nor U6173 (N_6173,N_5956,N_5929);
or U6174 (N_6174,N_5979,N_5932);
nand U6175 (N_6175,N_5949,N_5933);
or U6176 (N_6176,N_6008,N_5967);
nor U6177 (N_6177,N_5958,N_6010);
and U6178 (N_6178,N_6070,N_6038);
nand U6179 (N_6179,N_5949,N_5998);
nor U6180 (N_6180,N_5999,N_5986);
and U6181 (N_6181,N_6006,N_5956);
and U6182 (N_6182,N_6007,N_6026);
xnor U6183 (N_6183,N_5979,N_5968);
xnor U6184 (N_6184,N_5948,N_6032);
xnor U6185 (N_6185,N_5958,N_6038);
nor U6186 (N_6186,N_5937,N_6049);
nor U6187 (N_6187,N_5973,N_5988);
nand U6188 (N_6188,N_6001,N_5945);
or U6189 (N_6189,N_5995,N_6028);
and U6190 (N_6190,N_6066,N_6023);
or U6191 (N_6191,N_5927,N_6061);
nand U6192 (N_6192,N_6046,N_5923);
nor U6193 (N_6193,N_5988,N_6032);
xnor U6194 (N_6194,N_5992,N_6057);
nor U6195 (N_6195,N_5976,N_6002);
xor U6196 (N_6196,N_6071,N_6050);
xnor U6197 (N_6197,N_6055,N_5946);
nor U6198 (N_6198,N_6004,N_6036);
nand U6199 (N_6199,N_6078,N_5936);
or U6200 (N_6200,N_5921,N_6066);
xnor U6201 (N_6201,N_6079,N_5966);
nand U6202 (N_6202,N_5973,N_5949);
nor U6203 (N_6203,N_5992,N_5953);
and U6204 (N_6204,N_6021,N_5936);
and U6205 (N_6205,N_5925,N_5949);
nor U6206 (N_6206,N_5994,N_6018);
and U6207 (N_6207,N_6050,N_6062);
and U6208 (N_6208,N_5939,N_6020);
xor U6209 (N_6209,N_5973,N_6041);
xor U6210 (N_6210,N_5930,N_5931);
or U6211 (N_6211,N_6018,N_5998);
xor U6212 (N_6212,N_5923,N_5946);
and U6213 (N_6213,N_6003,N_6046);
nand U6214 (N_6214,N_5944,N_6026);
and U6215 (N_6215,N_5941,N_5959);
nand U6216 (N_6216,N_6043,N_5992);
xnor U6217 (N_6217,N_5929,N_5933);
and U6218 (N_6218,N_6004,N_6008);
and U6219 (N_6219,N_6016,N_6071);
nor U6220 (N_6220,N_5978,N_6042);
nor U6221 (N_6221,N_5930,N_6008);
nor U6222 (N_6222,N_6053,N_5984);
nor U6223 (N_6223,N_6028,N_6070);
nand U6224 (N_6224,N_5927,N_5988);
nand U6225 (N_6225,N_6013,N_6018);
or U6226 (N_6226,N_6034,N_6033);
or U6227 (N_6227,N_6062,N_6012);
nand U6228 (N_6228,N_5934,N_5999);
or U6229 (N_6229,N_5928,N_6004);
and U6230 (N_6230,N_6047,N_6017);
nor U6231 (N_6231,N_6007,N_5991);
nand U6232 (N_6232,N_5938,N_6057);
nand U6233 (N_6233,N_5973,N_5974);
and U6234 (N_6234,N_6045,N_6067);
or U6235 (N_6235,N_6064,N_6009);
and U6236 (N_6236,N_5939,N_6035);
xnor U6237 (N_6237,N_6055,N_5942);
or U6238 (N_6238,N_5964,N_6029);
or U6239 (N_6239,N_6071,N_5966);
xnor U6240 (N_6240,N_6191,N_6173);
or U6241 (N_6241,N_6128,N_6195);
and U6242 (N_6242,N_6157,N_6132);
nor U6243 (N_6243,N_6108,N_6081);
or U6244 (N_6244,N_6158,N_6156);
xnor U6245 (N_6245,N_6089,N_6091);
and U6246 (N_6246,N_6144,N_6224);
nor U6247 (N_6247,N_6206,N_6117);
or U6248 (N_6248,N_6112,N_6134);
or U6249 (N_6249,N_6237,N_6119);
nor U6250 (N_6250,N_6236,N_6129);
and U6251 (N_6251,N_6087,N_6109);
or U6252 (N_6252,N_6226,N_6232);
xnor U6253 (N_6253,N_6127,N_6203);
nor U6254 (N_6254,N_6110,N_6220);
nand U6255 (N_6255,N_6212,N_6204);
nor U6256 (N_6256,N_6186,N_6178);
nand U6257 (N_6257,N_6163,N_6107);
xor U6258 (N_6258,N_6187,N_6114);
nor U6259 (N_6259,N_6205,N_6227);
and U6260 (N_6260,N_6124,N_6126);
xnor U6261 (N_6261,N_6214,N_6201);
and U6262 (N_6262,N_6218,N_6153);
xor U6263 (N_6263,N_6170,N_6202);
and U6264 (N_6264,N_6105,N_6100);
nand U6265 (N_6265,N_6184,N_6139);
and U6266 (N_6266,N_6185,N_6164);
nor U6267 (N_6267,N_6116,N_6149);
or U6268 (N_6268,N_6094,N_6123);
nor U6269 (N_6269,N_6148,N_6145);
nand U6270 (N_6270,N_6097,N_6189);
xor U6271 (N_6271,N_6172,N_6138);
xnor U6272 (N_6272,N_6221,N_6130);
and U6273 (N_6273,N_6135,N_6179);
nand U6274 (N_6274,N_6235,N_6151);
xor U6275 (N_6275,N_6154,N_6175);
nor U6276 (N_6276,N_6150,N_6161);
nor U6277 (N_6277,N_6181,N_6152);
and U6278 (N_6278,N_6197,N_6222);
and U6279 (N_6279,N_6136,N_6106);
and U6280 (N_6280,N_6193,N_6217);
nand U6281 (N_6281,N_6162,N_6099);
nor U6282 (N_6282,N_6141,N_6165);
nand U6283 (N_6283,N_6121,N_6103);
nor U6284 (N_6284,N_6190,N_6223);
or U6285 (N_6285,N_6102,N_6115);
xor U6286 (N_6286,N_6207,N_6200);
nand U6287 (N_6287,N_6167,N_6233);
nor U6288 (N_6288,N_6092,N_6182);
or U6289 (N_6289,N_6155,N_6096);
nor U6290 (N_6290,N_6180,N_6090);
nand U6291 (N_6291,N_6111,N_6176);
and U6292 (N_6292,N_6125,N_6146);
and U6293 (N_6293,N_6209,N_6082);
or U6294 (N_6294,N_6085,N_6215);
nand U6295 (N_6295,N_6228,N_6143);
nand U6296 (N_6296,N_6171,N_6086);
nor U6297 (N_6297,N_6160,N_6198);
xor U6298 (N_6298,N_6177,N_6140);
nor U6299 (N_6299,N_6196,N_6210);
and U6300 (N_6300,N_6213,N_6238);
and U6301 (N_6301,N_6231,N_6120);
and U6302 (N_6302,N_6118,N_6183);
nor U6303 (N_6303,N_6122,N_6083);
xnor U6304 (N_6304,N_6093,N_6239);
nor U6305 (N_6305,N_6188,N_6159);
xnor U6306 (N_6306,N_6234,N_6095);
xnor U6307 (N_6307,N_6219,N_6230);
and U6308 (N_6308,N_6133,N_6208);
or U6309 (N_6309,N_6147,N_6169);
nand U6310 (N_6310,N_6131,N_6216);
or U6311 (N_6311,N_6194,N_6084);
nor U6312 (N_6312,N_6192,N_6080);
nand U6313 (N_6313,N_6113,N_6174);
nand U6314 (N_6314,N_6088,N_6104);
nor U6315 (N_6315,N_6137,N_6166);
or U6316 (N_6316,N_6225,N_6199);
and U6317 (N_6317,N_6229,N_6168);
or U6318 (N_6318,N_6142,N_6211);
xnor U6319 (N_6319,N_6098,N_6101);
or U6320 (N_6320,N_6225,N_6202);
xnor U6321 (N_6321,N_6110,N_6145);
and U6322 (N_6322,N_6147,N_6209);
and U6323 (N_6323,N_6237,N_6127);
or U6324 (N_6324,N_6215,N_6115);
xor U6325 (N_6325,N_6085,N_6140);
xnor U6326 (N_6326,N_6127,N_6105);
and U6327 (N_6327,N_6108,N_6182);
nor U6328 (N_6328,N_6170,N_6131);
nor U6329 (N_6329,N_6207,N_6177);
nor U6330 (N_6330,N_6223,N_6099);
nor U6331 (N_6331,N_6086,N_6203);
xor U6332 (N_6332,N_6221,N_6186);
nor U6333 (N_6333,N_6195,N_6096);
and U6334 (N_6334,N_6197,N_6108);
xnor U6335 (N_6335,N_6155,N_6207);
nor U6336 (N_6336,N_6190,N_6174);
xor U6337 (N_6337,N_6106,N_6156);
and U6338 (N_6338,N_6142,N_6095);
xor U6339 (N_6339,N_6192,N_6138);
xor U6340 (N_6340,N_6228,N_6144);
or U6341 (N_6341,N_6084,N_6232);
xnor U6342 (N_6342,N_6105,N_6083);
and U6343 (N_6343,N_6190,N_6213);
nor U6344 (N_6344,N_6146,N_6194);
nand U6345 (N_6345,N_6094,N_6204);
or U6346 (N_6346,N_6159,N_6231);
or U6347 (N_6347,N_6126,N_6129);
or U6348 (N_6348,N_6163,N_6223);
and U6349 (N_6349,N_6083,N_6148);
and U6350 (N_6350,N_6114,N_6204);
nor U6351 (N_6351,N_6213,N_6156);
nor U6352 (N_6352,N_6108,N_6146);
nor U6353 (N_6353,N_6097,N_6088);
xor U6354 (N_6354,N_6218,N_6217);
nand U6355 (N_6355,N_6111,N_6110);
nor U6356 (N_6356,N_6087,N_6104);
nor U6357 (N_6357,N_6193,N_6151);
and U6358 (N_6358,N_6148,N_6190);
xor U6359 (N_6359,N_6093,N_6205);
and U6360 (N_6360,N_6131,N_6166);
or U6361 (N_6361,N_6166,N_6176);
nand U6362 (N_6362,N_6097,N_6126);
nand U6363 (N_6363,N_6205,N_6163);
nor U6364 (N_6364,N_6212,N_6180);
nor U6365 (N_6365,N_6161,N_6218);
nor U6366 (N_6366,N_6116,N_6174);
nor U6367 (N_6367,N_6160,N_6215);
nand U6368 (N_6368,N_6194,N_6136);
and U6369 (N_6369,N_6231,N_6147);
or U6370 (N_6370,N_6142,N_6221);
nor U6371 (N_6371,N_6105,N_6158);
nand U6372 (N_6372,N_6132,N_6206);
xor U6373 (N_6373,N_6216,N_6223);
xnor U6374 (N_6374,N_6231,N_6224);
and U6375 (N_6375,N_6144,N_6214);
and U6376 (N_6376,N_6232,N_6119);
xnor U6377 (N_6377,N_6151,N_6102);
xnor U6378 (N_6378,N_6082,N_6213);
nand U6379 (N_6379,N_6154,N_6156);
nor U6380 (N_6380,N_6116,N_6102);
nor U6381 (N_6381,N_6122,N_6081);
nor U6382 (N_6382,N_6100,N_6200);
xnor U6383 (N_6383,N_6111,N_6131);
nand U6384 (N_6384,N_6081,N_6121);
or U6385 (N_6385,N_6231,N_6083);
and U6386 (N_6386,N_6216,N_6193);
and U6387 (N_6387,N_6209,N_6206);
and U6388 (N_6388,N_6234,N_6181);
or U6389 (N_6389,N_6215,N_6128);
nor U6390 (N_6390,N_6166,N_6183);
and U6391 (N_6391,N_6108,N_6227);
nand U6392 (N_6392,N_6106,N_6161);
xnor U6393 (N_6393,N_6090,N_6154);
and U6394 (N_6394,N_6230,N_6192);
nand U6395 (N_6395,N_6224,N_6123);
xor U6396 (N_6396,N_6094,N_6151);
or U6397 (N_6397,N_6169,N_6090);
nand U6398 (N_6398,N_6095,N_6184);
xnor U6399 (N_6399,N_6183,N_6192);
xnor U6400 (N_6400,N_6380,N_6370);
and U6401 (N_6401,N_6361,N_6285);
xnor U6402 (N_6402,N_6310,N_6265);
and U6403 (N_6403,N_6271,N_6297);
nand U6404 (N_6404,N_6303,N_6321);
nand U6405 (N_6405,N_6358,N_6248);
xor U6406 (N_6406,N_6338,N_6342);
nor U6407 (N_6407,N_6278,N_6392);
nand U6408 (N_6408,N_6389,N_6391);
nor U6409 (N_6409,N_6256,N_6262);
and U6410 (N_6410,N_6384,N_6245);
nand U6411 (N_6411,N_6327,N_6296);
nand U6412 (N_6412,N_6330,N_6251);
nand U6413 (N_6413,N_6300,N_6311);
or U6414 (N_6414,N_6255,N_6395);
and U6415 (N_6415,N_6275,N_6366);
nand U6416 (N_6416,N_6242,N_6376);
and U6417 (N_6417,N_6273,N_6383);
and U6418 (N_6418,N_6346,N_6332);
and U6419 (N_6419,N_6249,N_6362);
and U6420 (N_6420,N_6369,N_6257);
and U6421 (N_6421,N_6315,N_6337);
or U6422 (N_6422,N_6368,N_6295);
nor U6423 (N_6423,N_6335,N_6250);
nor U6424 (N_6424,N_6339,N_6356);
xor U6425 (N_6425,N_6393,N_6287);
nand U6426 (N_6426,N_6318,N_6294);
xor U6427 (N_6427,N_6354,N_6390);
nor U6428 (N_6428,N_6373,N_6350);
or U6429 (N_6429,N_6279,N_6382);
or U6430 (N_6430,N_6284,N_6386);
xnor U6431 (N_6431,N_6398,N_6240);
nand U6432 (N_6432,N_6290,N_6241);
and U6433 (N_6433,N_6324,N_6293);
nand U6434 (N_6434,N_6291,N_6314);
or U6435 (N_6435,N_6276,N_6288);
or U6436 (N_6436,N_6349,N_6281);
and U6437 (N_6437,N_6360,N_6357);
nor U6438 (N_6438,N_6364,N_6266);
xor U6439 (N_6439,N_6283,N_6301);
and U6440 (N_6440,N_6286,N_6304);
xor U6441 (N_6441,N_6319,N_6308);
or U6442 (N_6442,N_6322,N_6329);
nor U6443 (N_6443,N_6313,N_6372);
or U6444 (N_6444,N_6307,N_6374);
nor U6445 (N_6445,N_6298,N_6359);
and U6446 (N_6446,N_6258,N_6247);
and U6447 (N_6447,N_6399,N_6254);
and U6448 (N_6448,N_6379,N_6306);
nand U6449 (N_6449,N_6312,N_6309);
nor U6450 (N_6450,N_6345,N_6347);
nand U6451 (N_6451,N_6326,N_6316);
and U6452 (N_6452,N_6394,N_6280);
or U6453 (N_6453,N_6269,N_6282);
or U6454 (N_6454,N_6253,N_6260);
nand U6455 (N_6455,N_6371,N_6352);
and U6456 (N_6456,N_6268,N_6317);
nand U6457 (N_6457,N_6387,N_6331);
and U6458 (N_6458,N_6377,N_6323);
nand U6459 (N_6459,N_6397,N_6320);
xor U6460 (N_6460,N_6375,N_6385);
nand U6461 (N_6461,N_6348,N_6270);
and U6462 (N_6462,N_6302,N_6344);
or U6463 (N_6463,N_6272,N_6334);
or U6464 (N_6464,N_6365,N_6259);
nor U6465 (N_6465,N_6267,N_6396);
or U6466 (N_6466,N_6340,N_6244);
nor U6467 (N_6467,N_6263,N_6305);
and U6468 (N_6468,N_6243,N_6299);
xnor U6469 (N_6469,N_6252,N_6363);
xor U6470 (N_6470,N_6336,N_6367);
xor U6471 (N_6471,N_6277,N_6355);
or U6472 (N_6472,N_6343,N_6246);
nor U6473 (N_6473,N_6378,N_6292);
or U6474 (N_6474,N_6333,N_6328);
or U6475 (N_6475,N_6289,N_6325);
xor U6476 (N_6476,N_6274,N_6261);
or U6477 (N_6477,N_6353,N_6388);
and U6478 (N_6478,N_6351,N_6341);
nor U6479 (N_6479,N_6381,N_6264);
nor U6480 (N_6480,N_6330,N_6388);
or U6481 (N_6481,N_6281,N_6367);
and U6482 (N_6482,N_6312,N_6364);
or U6483 (N_6483,N_6364,N_6321);
nand U6484 (N_6484,N_6350,N_6302);
xnor U6485 (N_6485,N_6384,N_6386);
nand U6486 (N_6486,N_6372,N_6267);
nand U6487 (N_6487,N_6398,N_6336);
xnor U6488 (N_6488,N_6281,N_6365);
or U6489 (N_6489,N_6380,N_6327);
xnor U6490 (N_6490,N_6323,N_6367);
xnor U6491 (N_6491,N_6344,N_6397);
and U6492 (N_6492,N_6299,N_6366);
xor U6493 (N_6493,N_6256,N_6279);
and U6494 (N_6494,N_6289,N_6368);
or U6495 (N_6495,N_6395,N_6314);
xnor U6496 (N_6496,N_6283,N_6297);
xnor U6497 (N_6497,N_6381,N_6376);
and U6498 (N_6498,N_6300,N_6266);
xor U6499 (N_6499,N_6371,N_6363);
nor U6500 (N_6500,N_6343,N_6300);
and U6501 (N_6501,N_6345,N_6308);
xor U6502 (N_6502,N_6344,N_6274);
nor U6503 (N_6503,N_6309,N_6299);
nand U6504 (N_6504,N_6268,N_6253);
xnor U6505 (N_6505,N_6263,N_6372);
xor U6506 (N_6506,N_6271,N_6248);
nor U6507 (N_6507,N_6313,N_6290);
or U6508 (N_6508,N_6323,N_6349);
or U6509 (N_6509,N_6245,N_6378);
nor U6510 (N_6510,N_6390,N_6291);
and U6511 (N_6511,N_6388,N_6247);
xor U6512 (N_6512,N_6276,N_6250);
xor U6513 (N_6513,N_6353,N_6244);
and U6514 (N_6514,N_6279,N_6350);
nand U6515 (N_6515,N_6387,N_6322);
or U6516 (N_6516,N_6339,N_6384);
and U6517 (N_6517,N_6256,N_6316);
xnor U6518 (N_6518,N_6244,N_6312);
nand U6519 (N_6519,N_6351,N_6288);
xnor U6520 (N_6520,N_6339,N_6245);
nor U6521 (N_6521,N_6397,N_6387);
or U6522 (N_6522,N_6362,N_6307);
xor U6523 (N_6523,N_6382,N_6398);
or U6524 (N_6524,N_6301,N_6338);
or U6525 (N_6525,N_6391,N_6276);
and U6526 (N_6526,N_6394,N_6266);
and U6527 (N_6527,N_6373,N_6381);
nand U6528 (N_6528,N_6259,N_6338);
or U6529 (N_6529,N_6354,N_6309);
nor U6530 (N_6530,N_6364,N_6294);
nand U6531 (N_6531,N_6349,N_6301);
nand U6532 (N_6532,N_6367,N_6291);
nand U6533 (N_6533,N_6336,N_6284);
nand U6534 (N_6534,N_6300,N_6354);
or U6535 (N_6535,N_6399,N_6344);
nand U6536 (N_6536,N_6248,N_6360);
xnor U6537 (N_6537,N_6284,N_6246);
or U6538 (N_6538,N_6248,N_6311);
and U6539 (N_6539,N_6354,N_6357);
nor U6540 (N_6540,N_6363,N_6253);
xor U6541 (N_6541,N_6274,N_6378);
xor U6542 (N_6542,N_6248,N_6362);
and U6543 (N_6543,N_6281,N_6370);
or U6544 (N_6544,N_6250,N_6371);
xnor U6545 (N_6545,N_6365,N_6323);
or U6546 (N_6546,N_6334,N_6275);
xor U6547 (N_6547,N_6391,N_6270);
and U6548 (N_6548,N_6245,N_6362);
nor U6549 (N_6549,N_6317,N_6388);
or U6550 (N_6550,N_6356,N_6247);
or U6551 (N_6551,N_6389,N_6272);
nor U6552 (N_6552,N_6391,N_6315);
nor U6553 (N_6553,N_6350,N_6390);
nand U6554 (N_6554,N_6278,N_6367);
and U6555 (N_6555,N_6304,N_6301);
xnor U6556 (N_6556,N_6383,N_6367);
xor U6557 (N_6557,N_6308,N_6260);
xnor U6558 (N_6558,N_6390,N_6376);
or U6559 (N_6559,N_6368,N_6288);
nand U6560 (N_6560,N_6533,N_6527);
or U6561 (N_6561,N_6546,N_6525);
nand U6562 (N_6562,N_6521,N_6534);
nor U6563 (N_6563,N_6410,N_6436);
xor U6564 (N_6564,N_6460,N_6452);
or U6565 (N_6565,N_6441,N_6400);
nand U6566 (N_6566,N_6494,N_6541);
or U6567 (N_6567,N_6538,N_6415);
nand U6568 (N_6568,N_6505,N_6475);
xor U6569 (N_6569,N_6483,N_6522);
nand U6570 (N_6570,N_6515,N_6555);
and U6571 (N_6571,N_6486,N_6556);
xnor U6572 (N_6572,N_6422,N_6518);
nor U6573 (N_6573,N_6401,N_6550);
or U6574 (N_6574,N_6524,N_6531);
nor U6575 (N_6575,N_6451,N_6544);
nor U6576 (N_6576,N_6434,N_6517);
or U6577 (N_6577,N_6498,N_6514);
nand U6578 (N_6578,N_6423,N_6501);
or U6579 (N_6579,N_6411,N_6542);
nor U6580 (N_6580,N_6419,N_6462);
xor U6581 (N_6581,N_6406,N_6511);
nor U6582 (N_6582,N_6520,N_6408);
nand U6583 (N_6583,N_6444,N_6543);
nor U6584 (N_6584,N_6450,N_6438);
or U6585 (N_6585,N_6548,N_6413);
nor U6586 (N_6586,N_6496,N_6536);
and U6587 (N_6587,N_6489,N_6557);
nand U6588 (N_6588,N_6491,N_6559);
or U6589 (N_6589,N_6487,N_6468);
nor U6590 (N_6590,N_6509,N_6537);
xnor U6591 (N_6591,N_6480,N_6429);
and U6592 (N_6592,N_6530,N_6549);
and U6593 (N_6593,N_6495,N_6448);
or U6594 (N_6594,N_6492,N_6507);
nor U6595 (N_6595,N_6532,N_6463);
nand U6596 (N_6596,N_6461,N_6516);
and U6597 (N_6597,N_6512,N_6403);
and U6598 (N_6598,N_6528,N_6523);
and U6599 (N_6599,N_6412,N_6407);
or U6600 (N_6600,N_6519,N_6497);
or U6601 (N_6601,N_6437,N_6464);
nor U6602 (N_6602,N_6470,N_6425);
xnor U6603 (N_6603,N_6535,N_6459);
xor U6604 (N_6604,N_6551,N_6427);
xor U6605 (N_6605,N_6502,N_6504);
nor U6606 (N_6606,N_6449,N_6402);
nand U6607 (N_6607,N_6446,N_6539);
nor U6608 (N_6608,N_6424,N_6405);
nor U6609 (N_6609,N_6490,N_6478);
xnor U6610 (N_6610,N_6529,N_6455);
nand U6611 (N_6611,N_6440,N_6477);
nand U6612 (N_6612,N_6474,N_6476);
and U6613 (N_6613,N_6493,N_6430);
or U6614 (N_6614,N_6552,N_6558);
and U6615 (N_6615,N_6445,N_6500);
xor U6616 (N_6616,N_6466,N_6442);
and U6617 (N_6617,N_6457,N_6417);
nand U6618 (N_6618,N_6472,N_6508);
nor U6619 (N_6619,N_6467,N_6488);
and U6620 (N_6620,N_6484,N_6447);
nor U6621 (N_6621,N_6547,N_6454);
nand U6622 (N_6622,N_6526,N_6431);
or U6623 (N_6623,N_6540,N_6414);
and U6624 (N_6624,N_6453,N_6510);
or U6625 (N_6625,N_6469,N_6421);
and U6626 (N_6626,N_6433,N_6485);
xor U6627 (N_6627,N_6428,N_6554);
nor U6628 (N_6628,N_6432,N_6439);
nor U6629 (N_6629,N_6545,N_6426);
nor U6630 (N_6630,N_6553,N_6473);
xor U6631 (N_6631,N_6456,N_6471);
nand U6632 (N_6632,N_6513,N_6479);
nand U6633 (N_6633,N_6416,N_6404);
nand U6634 (N_6634,N_6503,N_6482);
xnor U6635 (N_6635,N_6481,N_6420);
nor U6636 (N_6636,N_6499,N_6506);
and U6637 (N_6637,N_6418,N_6443);
or U6638 (N_6638,N_6435,N_6409);
nand U6639 (N_6639,N_6458,N_6465);
nand U6640 (N_6640,N_6430,N_6495);
xor U6641 (N_6641,N_6446,N_6524);
or U6642 (N_6642,N_6470,N_6473);
or U6643 (N_6643,N_6470,N_6558);
nand U6644 (N_6644,N_6534,N_6416);
or U6645 (N_6645,N_6516,N_6465);
nand U6646 (N_6646,N_6451,N_6480);
or U6647 (N_6647,N_6449,N_6508);
and U6648 (N_6648,N_6453,N_6444);
xor U6649 (N_6649,N_6532,N_6544);
xor U6650 (N_6650,N_6544,N_6411);
and U6651 (N_6651,N_6459,N_6479);
and U6652 (N_6652,N_6426,N_6469);
or U6653 (N_6653,N_6436,N_6475);
nor U6654 (N_6654,N_6455,N_6449);
and U6655 (N_6655,N_6557,N_6408);
and U6656 (N_6656,N_6472,N_6435);
nor U6657 (N_6657,N_6556,N_6495);
and U6658 (N_6658,N_6527,N_6548);
nor U6659 (N_6659,N_6539,N_6489);
or U6660 (N_6660,N_6456,N_6499);
and U6661 (N_6661,N_6518,N_6542);
nor U6662 (N_6662,N_6459,N_6468);
and U6663 (N_6663,N_6456,N_6451);
and U6664 (N_6664,N_6536,N_6526);
and U6665 (N_6665,N_6413,N_6426);
nor U6666 (N_6666,N_6428,N_6526);
xnor U6667 (N_6667,N_6471,N_6503);
and U6668 (N_6668,N_6437,N_6504);
nor U6669 (N_6669,N_6514,N_6546);
nand U6670 (N_6670,N_6449,N_6475);
xnor U6671 (N_6671,N_6506,N_6538);
nor U6672 (N_6672,N_6457,N_6473);
nor U6673 (N_6673,N_6401,N_6470);
xnor U6674 (N_6674,N_6507,N_6529);
and U6675 (N_6675,N_6483,N_6457);
nand U6676 (N_6676,N_6549,N_6468);
and U6677 (N_6677,N_6456,N_6466);
or U6678 (N_6678,N_6414,N_6551);
nor U6679 (N_6679,N_6448,N_6416);
nor U6680 (N_6680,N_6519,N_6413);
and U6681 (N_6681,N_6556,N_6446);
or U6682 (N_6682,N_6534,N_6497);
nor U6683 (N_6683,N_6406,N_6474);
nand U6684 (N_6684,N_6436,N_6422);
or U6685 (N_6685,N_6442,N_6417);
or U6686 (N_6686,N_6437,N_6541);
nand U6687 (N_6687,N_6509,N_6525);
and U6688 (N_6688,N_6448,N_6430);
xnor U6689 (N_6689,N_6508,N_6455);
nand U6690 (N_6690,N_6533,N_6522);
or U6691 (N_6691,N_6423,N_6518);
xnor U6692 (N_6692,N_6439,N_6534);
or U6693 (N_6693,N_6444,N_6509);
or U6694 (N_6694,N_6493,N_6428);
and U6695 (N_6695,N_6407,N_6430);
nand U6696 (N_6696,N_6550,N_6540);
xor U6697 (N_6697,N_6505,N_6519);
nor U6698 (N_6698,N_6517,N_6487);
nand U6699 (N_6699,N_6430,N_6429);
or U6700 (N_6700,N_6465,N_6544);
nor U6701 (N_6701,N_6449,N_6515);
xnor U6702 (N_6702,N_6538,N_6455);
and U6703 (N_6703,N_6557,N_6498);
nand U6704 (N_6704,N_6519,N_6465);
or U6705 (N_6705,N_6486,N_6542);
xor U6706 (N_6706,N_6488,N_6513);
nand U6707 (N_6707,N_6532,N_6540);
and U6708 (N_6708,N_6481,N_6437);
or U6709 (N_6709,N_6462,N_6416);
nand U6710 (N_6710,N_6557,N_6539);
nand U6711 (N_6711,N_6454,N_6499);
and U6712 (N_6712,N_6425,N_6525);
nor U6713 (N_6713,N_6425,N_6473);
xor U6714 (N_6714,N_6532,N_6516);
xor U6715 (N_6715,N_6529,N_6539);
nor U6716 (N_6716,N_6469,N_6452);
and U6717 (N_6717,N_6409,N_6424);
or U6718 (N_6718,N_6435,N_6444);
xnor U6719 (N_6719,N_6428,N_6445);
nor U6720 (N_6720,N_6621,N_6583);
nand U6721 (N_6721,N_6714,N_6612);
and U6722 (N_6722,N_6708,N_6588);
and U6723 (N_6723,N_6581,N_6620);
xnor U6724 (N_6724,N_6691,N_6683);
or U6725 (N_6725,N_6649,N_6654);
nand U6726 (N_6726,N_6681,N_6604);
nand U6727 (N_6727,N_6578,N_6693);
or U6728 (N_6728,N_6664,N_6695);
nor U6729 (N_6729,N_6670,N_6719);
nand U6730 (N_6730,N_6579,N_6584);
nor U6731 (N_6731,N_6647,N_6685);
and U6732 (N_6732,N_6630,N_6585);
nor U6733 (N_6733,N_6669,N_6663);
and U6734 (N_6734,N_6640,N_6700);
nor U6735 (N_6735,N_6594,N_6682);
nand U6736 (N_6736,N_6701,N_6635);
and U6737 (N_6737,N_6710,N_6570);
xnor U6738 (N_6738,N_6618,N_6602);
and U6739 (N_6739,N_6706,N_6629);
xnor U6740 (N_6740,N_6697,N_6613);
or U6741 (N_6741,N_6687,N_6605);
nand U6742 (N_6742,N_6597,N_6591);
or U6743 (N_6743,N_6600,N_6567);
and U6744 (N_6744,N_6679,N_6673);
or U6745 (N_6745,N_6653,N_6580);
xnor U6746 (N_6746,N_6672,N_6717);
nand U6747 (N_6747,N_6582,N_6641);
nor U6748 (N_6748,N_6587,N_6686);
and U6749 (N_6749,N_6575,N_6611);
or U6750 (N_6750,N_6662,N_6638);
or U6751 (N_6751,N_6655,N_6651);
or U6752 (N_6752,N_6625,N_6631);
xor U6753 (N_6753,N_6711,N_6639);
xnor U6754 (N_6754,N_6565,N_6633);
xor U6755 (N_6755,N_6696,N_6632);
or U6756 (N_6756,N_6688,N_6610);
nor U6757 (N_6757,N_6677,N_6576);
nand U6758 (N_6758,N_6657,N_6590);
and U6759 (N_6759,N_6628,N_6692);
nor U6760 (N_6760,N_6564,N_6569);
nor U6761 (N_6761,N_6577,N_6595);
xor U6762 (N_6762,N_6699,N_6703);
nand U6763 (N_6763,N_6680,N_6665);
or U6764 (N_6764,N_6603,N_6656);
or U6765 (N_6765,N_6676,N_6709);
or U6766 (N_6766,N_6593,N_6599);
or U6767 (N_6767,N_6619,N_6623);
nand U6768 (N_6768,N_6586,N_6626);
nor U6769 (N_6769,N_6560,N_6608);
and U6770 (N_6770,N_6689,N_6667);
and U6771 (N_6771,N_6616,N_6715);
and U6772 (N_6772,N_6648,N_6675);
or U6773 (N_6773,N_6661,N_6637);
nand U6774 (N_6774,N_6596,N_6573);
nor U6775 (N_6775,N_6592,N_6694);
nor U6776 (N_6776,N_6666,N_6615);
and U6777 (N_6777,N_6622,N_6617);
and U6778 (N_6778,N_6624,N_6643);
or U6779 (N_6779,N_6601,N_6644);
nor U6780 (N_6780,N_6659,N_6652);
or U6781 (N_6781,N_6713,N_6634);
or U6782 (N_6782,N_6606,N_6716);
nand U6783 (N_6783,N_6650,N_6646);
nor U6784 (N_6784,N_6568,N_6561);
or U6785 (N_6785,N_6678,N_6566);
or U6786 (N_6786,N_6712,N_6574);
xor U6787 (N_6787,N_6627,N_6589);
and U6788 (N_6788,N_6607,N_6671);
or U6789 (N_6789,N_6668,N_6642);
xor U6790 (N_6790,N_6690,N_6684);
or U6791 (N_6791,N_6702,N_6705);
nand U6792 (N_6792,N_6562,N_6698);
and U6793 (N_6793,N_6563,N_6609);
nor U6794 (N_6794,N_6645,N_6674);
nor U6795 (N_6795,N_6572,N_6636);
nand U6796 (N_6796,N_6571,N_6707);
and U6797 (N_6797,N_6614,N_6718);
and U6798 (N_6798,N_6598,N_6658);
or U6799 (N_6799,N_6660,N_6704);
xnor U6800 (N_6800,N_6691,N_6690);
or U6801 (N_6801,N_6599,N_6581);
or U6802 (N_6802,N_6590,N_6610);
nor U6803 (N_6803,N_6698,N_6585);
and U6804 (N_6804,N_6655,N_6611);
xnor U6805 (N_6805,N_6695,N_6713);
nand U6806 (N_6806,N_6667,N_6681);
and U6807 (N_6807,N_6605,N_6702);
nand U6808 (N_6808,N_6590,N_6686);
or U6809 (N_6809,N_6634,N_6578);
or U6810 (N_6810,N_6614,N_6699);
xnor U6811 (N_6811,N_6678,N_6709);
and U6812 (N_6812,N_6694,N_6633);
xnor U6813 (N_6813,N_6686,N_6647);
and U6814 (N_6814,N_6697,N_6666);
or U6815 (N_6815,N_6627,N_6638);
xnor U6816 (N_6816,N_6598,N_6573);
and U6817 (N_6817,N_6663,N_6662);
nand U6818 (N_6818,N_6673,N_6562);
xor U6819 (N_6819,N_6593,N_6654);
nor U6820 (N_6820,N_6641,N_6609);
and U6821 (N_6821,N_6569,N_6620);
nor U6822 (N_6822,N_6682,N_6609);
nand U6823 (N_6823,N_6646,N_6662);
xnor U6824 (N_6824,N_6567,N_6718);
nor U6825 (N_6825,N_6625,N_6695);
nor U6826 (N_6826,N_6667,N_6673);
nor U6827 (N_6827,N_6704,N_6587);
nand U6828 (N_6828,N_6703,N_6576);
xor U6829 (N_6829,N_6623,N_6685);
nor U6830 (N_6830,N_6572,N_6713);
and U6831 (N_6831,N_6658,N_6660);
nand U6832 (N_6832,N_6610,N_6616);
or U6833 (N_6833,N_6645,N_6683);
or U6834 (N_6834,N_6611,N_6619);
nand U6835 (N_6835,N_6619,N_6590);
xor U6836 (N_6836,N_6594,N_6593);
or U6837 (N_6837,N_6646,N_6587);
nand U6838 (N_6838,N_6575,N_6662);
xnor U6839 (N_6839,N_6640,N_6676);
nand U6840 (N_6840,N_6633,N_6579);
and U6841 (N_6841,N_6713,N_6647);
nand U6842 (N_6842,N_6567,N_6649);
xnor U6843 (N_6843,N_6641,N_6683);
nand U6844 (N_6844,N_6625,N_6620);
xnor U6845 (N_6845,N_6601,N_6604);
nand U6846 (N_6846,N_6702,N_6679);
or U6847 (N_6847,N_6690,N_6694);
nand U6848 (N_6848,N_6700,N_6608);
nand U6849 (N_6849,N_6701,N_6618);
or U6850 (N_6850,N_6614,N_6637);
and U6851 (N_6851,N_6562,N_6667);
nand U6852 (N_6852,N_6588,N_6638);
nand U6853 (N_6853,N_6566,N_6671);
and U6854 (N_6854,N_6675,N_6576);
xnor U6855 (N_6855,N_6706,N_6593);
and U6856 (N_6856,N_6695,N_6680);
xor U6857 (N_6857,N_6568,N_6700);
and U6858 (N_6858,N_6628,N_6719);
nand U6859 (N_6859,N_6617,N_6645);
nor U6860 (N_6860,N_6581,N_6679);
xor U6861 (N_6861,N_6581,N_6685);
nand U6862 (N_6862,N_6570,N_6567);
nor U6863 (N_6863,N_6656,N_6692);
nand U6864 (N_6864,N_6597,N_6696);
nand U6865 (N_6865,N_6581,N_6624);
nor U6866 (N_6866,N_6560,N_6630);
or U6867 (N_6867,N_6586,N_6627);
nand U6868 (N_6868,N_6596,N_6589);
or U6869 (N_6869,N_6681,N_6714);
and U6870 (N_6870,N_6592,N_6667);
xor U6871 (N_6871,N_6595,N_6623);
and U6872 (N_6872,N_6700,N_6697);
or U6873 (N_6873,N_6644,N_6608);
xor U6874 (N_6874,N_6667,N_6573);
nor U6875 (N_6875,N_6680,N_6596);
nand U6876 (N_6876,N_6685,N_6718);
or U6877 (N_6877,N_6713,N_6628);
and U6878 (N_6878,N_6706,N_6573);
or U6879 (N_6879,N_6656,N_6615);
xnor U6880 (N_6880,N_6825,N_6739);
nor U6881 (N_6881,N_6755,N_6868);
or U6882 (N_6882,N_6775,N_6758);
nor U6883 (N_6883,N_6753,N_6879);
or U6884 (N_6884,N_6781,N_6770);
and U6885 (N_6885,N_6807,N_6851);
nor U6886 (N_6886,N_6859,N_6789);
or U6887 (N_6887,N_6741,N_6757);
nor U6888 (N_6888,N_6801,N_6843);
nor U6889 (N_6889,N_6737,N_6805);
nor U6890 (N_6890,N_6867,N_6814);
nand U6891 (N_6891,N_6839,N_6724);
and U6892 (N_6892,N_6720,N_6762);
nand U6893 (N_6893,N_6874,N_6840);
nand U6894 (N_6894,N_6854,N_6733);
nand U6895 (N_6895,N_6742,N_6817);
nand U6896 (N_6896,N_6799,N_6873);
or U6897 (N_6897,N_6858,N_6752);
xnor U6898 (N_6898,N_6862,N_6782);
or U6899 (N_6899,N_6852,N_6878);
nor U6900 (N_6900,N_6783,N_6842);
nand U6901 (N_6901,N_6767,N_6725);
or U6902 (N_6902,N_6820,N_6802);
and U6903 (N_6903,N_6723,N_6750);
nor U6904 (N_6904,N_6732,N_6826);
nor U6905 (N_6905,N_6743,N_6827);
and U6906 (N_6906,N_6749,N_6777);
xnor U6907 (N_6907,N_6721,N_6822);
nor U6908 (N_6908,N_6809,N_6846);
nor U6909 (N_6909,N_6772,N_6808);
xor U6910 (N_6910,N_6869,N_6759);
nor U6911 (N_6911,N_6788,N_6857);
xnor U6912 (N_6912,N_6797,N_6790);
xor U6913 (N_6913,N_6727,N_6824);
nor U6914 (N_6914,N_6796,N_6779);
nand U6915 (N_6915,N_6804,N_6738);
nor U6916 (N_6916,N_6860,N_6792);
and U6917 (N_6917,N_6844,N_6751);
xor U6918 (N_6918,N_6806,N_6819);
nand U6919 (N_6919,N_6744,N_6847);
or U6920 (N_6920,N_6877,N_6754);
xor U6921 (N_6921,N_6821,N_6871);
and U6922 (N_6922,N_6803,N_6866);
xor U6923 (N_6923,N_6828,N_6810);
or U6924 (N_6924,N_6823,N_6766);
nand U6925 (N_6925,N_6769,N_6785);
or U6926 (N_6926,N_6756,N_6872);
xor U6927 (N_6927,N_6793,N_6748);
nand U6928 (N_6928,N_6856,N_6731);
nand U6929 (N_6929,N_6729,N_6816);
or U6930 (N_6930,N_6875,N_6787);
nand U6931 (N_6931,N_6855,N_6813);
or U6932 (N_6932,N_6849,N_6876);
and U6933 (N_6933,N_6726,N_6845);
nor U6934 (N_6934,N_6734,N_6761);
and U6935 (N_6935,N_6835,N_6773);
nand U6936 (N_6936,N_6776,N_6763);
and U6937 (N_6937,N_6746,N_6747);
or U6938 (N_6938,N_6836,N_6861);
nand U6939 (N_6939,N_6829,N_6853);
and U6940 (N_6940,N_6798,N_6864);
or U6941 (N_6941,N_6768,N_6794);
xnor U6942 (N_6942,N_6831,N_6736);
or U6943 (N_6943,N_6730,N_6786);
nand U6944 (N_6944,N_6780,N_6815);
nor U6945 (N_6945,N_6811,N_6838);
and U6946 (N_6946,N_6870,N_6795);
xor U6947 (N_6947,N_6735,N_6760);
nor U6948 (N_6948,N_6771,N_6745);
nand U6949 (N_6949,N_6800,N_6774);
or U6950 (N_6950,N_6818,N_6722);
xor U6951 (N_6951,N_6812,N_6830);
nor U6952 (N_6952,N_6765,N_6848);
or U6953 (N_6953,N_6833,N_6740);
or U6954 (N_6954,N_6728,N_6865);
nand U6955 (N_6955,N_6832,N_6850);
and U6956 (N_6956,N_6834,N_6837);
nand U6957 (N_6957,N_6841,N_6791);
nand U6958 (N_6958,N_6778,N_6764);
and U6959 (N_6959,N_6784,N_6863);
nor U6960 (N_6960,N_6759,N_6729);
and U6961 (N_6961,N_6865,N_6812);
or U6962 (N_6962,N_6843,N_6790);
or U6963 (N_6963,N_6756,N_6823);
xnor U6964 (N_6964,N_6800,N_6830);
and U6965 (N_6965,N_6773,N_6864);
or U6966 (N_6966,N_6865,N_6769);
nand U6967 (N_6967,N_6809,N_6822);
nor U6968 (N_6968,N_6837,N_6745);
nand U6969 (N_6969,N_6831,N_6873);
nand U6970 (N_6970,N_6798,N_6824);
nand U6971 (N_6971,N_6810,N_6856);
and U6972 (N_6972,N_6817,N_6802);
nand U6973 (N_6973,N_6804,N_6747);
nand U6974 (N_6974,N_6800,N_6759);
and U6975 (N_6975,N_6838,N_6829);
xnor U6976 (N_6976,N_6850,N_6847);
xor U6977 (N_6977,N_6794,N_6769);
xor U6978 (N_6978,N_6811,N_6820);
or U6979 (N_6979,N_6831,N_6742);
and U6980 (N_6980,N_6863,N_6749);
xnor U6981 (N_6981,N_6811,N_6816);
nand U6982 (N_6982,N_6801,N_6837);
nor U6983 (N_6983,N_6722,N_6732);
or U6984 (N_6984,N_6765,N_6779);
nor U6985 (N_6985,N_6768,N_6855);
nand U6986 (N_6986,N_6736,N_6789);
xnor U6987 (N_6987,N_6804,N_6877);
nand U6988 (N_6988,N_6763,N_6858);
or U6989 (N_6989,N_6750,N_6864);
xnor U6990 (N_6990,N_6804,N_6782);
nor U6991 (N_6991,N_6820,N_6736);
xnor U6992 (N_6992,N_6822,N_6837);
and U6993 (N_6993,N_6807,N_6744);
nor U6994 (N_6994,N_6879,N_6858);
nor U6995 (N_6995,N_6775,N_6749);
or U6996 (N_6996,N_6797,N_6840);
nand U6997 (N_6997,N_6742,N_6815);
or U6998 (N_6998,N_6864,N_6737);
nand U6999 (N_6999,N_6809,N_6849);
or U7000 (N_7000,N_6877,N_6766);
xor U7001 (N_7001,N_6804,N_6789);
nand U7002 (N_7002,N_6786,N_6875);
nand U7003 (N_7003,N_6827,N_6842);
and U7004 (N_7004,N_6747,N_6740);
nand U7005 (N_7005,N_6738,N_6729);
or U7006 (N_7006,N_6764,N_6829);
nor U7007 (N_7007,N_6751,N_6747);
and U7008 (N_7008,N_6801,N_6836);
nand U7009 (N_7009,N_6828,N_6833);
xnor U7010 (N_7010,N_6847,N_6830);
or U7011 (N_7011,N_6768,N_6806);
xor U7012 (N_7012,N_6782,N_6847);
nand U7013 (N_7013,N_6764,N_6869);
and U7014 (N_7014,N_6837,N_6871);
nor U7015 (N_7015,N_6822,N_6779);
or U7016 (N_7016,N_6805,N_6760);
nand U7017 (N_7017,N_6865,N_6851);
or U7018 (N_7018,N_6864,N_6863);
and U7019 (N_7019,N_6775,N_6767);
or U7020 (N_7020,N_6878,N_6822);
xnor U7021 (N_7021,N_6826,N_6763);
or U7022 (N_7022,N_6777,N_6780);
nor U7023 (N_7023,N_6743,N_6844);
or U7024 (N_7024,N_6767,N_6805);
nand U7025 (N_7025,N_6840,N_6753);
xor U7026 (N_7026,N_6831,N_6791);
and U7027 (N_7027,N_6767,N_6758);
or U7028 (N_7028,N_6817,N_6777);
nor U7029 (N_7029,N_6869,N_6815);
nor U7030 (N_7030,N_6793,N_6874);
or U7031 (N_7031,N_6864,N_6729);
or U7032 (N_7032,N_6866,N_6765);
xnor U7033 (N_7033,N_6858,N_6847);
xor U7034 (N_7034,N_6825,N_6749);
or U7035 (N_7035,N_6729,N_6774);
nor U7036 (N_7036,N_6793,N_6805);
xor U7037 (N_7037,N_6837,N_6774);
nor U7038 (N_7038,N_6865,N_6775);
nand U7039 (N_7039,N_6812,N_6854);
xnor U7040 (N_7040,N_6884,N_6968);
or U7041 (N_7041,N_7024,N_7013);
and U7042 (N_7042,N_7038,N_6944);
and U7043 (N_7043,N_6967,N_6986);
or U7044 (N_7044,N_7037,N_6909);
or U7045 (N_7045,N_6906,N_6932);
nand U7046 (N_7046,N_6960,N_6907);
nand U7047 (N_7047,N_6969,N_7019);
nor U7048 (N_7048,N_6953,N_6928);
or U7049 (N_7049,N_6898,N_7018);
nor U7050 (N_7050,N_6970,N_6983);
and U7051 (N_7051,N_6938,N_6995);
or U7052 (N_7052,N_6966,N_6971);
and U7053 (N_7053,N_6993,N_6905);
or U7054 (N_7054,N_6977,N_6998);
or U7055 (N_7055,N_6888,N_6997);
or U7056 (N_7056,N_6955,N_6891);
nand U7057 (N_7057,N_7000,N_7023);
nor U7058 (N_7058,N_7014,N_6918);
xnor U7059 (N_7059,N_7026,N_6881);
nor U7060 (N_7060,N_6999,N_7010);
nor U7061 (N_7061,N_6902,N_6889);
nor U7062 (N_7062,N_6931,N_7015);
xnor U7063 (N_7063,N_6935,N_7017);
nand U7064 (N_7064,N_6919,N_6947);
nand U7065 (N_7065,N_7009,N_7030);
nand U7066 (N_7066,N_6943,N_7008);
nor U7067 (N_7067,N_7001,N_6912);
or U7068 (N_7068,N_6886,N_7004);
xnor U7069 (N_7069,N_6990,N_6926);
nand U7070 (N_7070,N_7031,N_6894);
nand U7071 (N_7071,N_6946,N_6893);
xnor U7072 (N_7072,N_7022,N_6930);
nor U7073 (N_7073,N_6896,N_7006);
or U7074 (N_7074,N_6937,N_7028);
or U7075 (N_7075,N_6929,N_6957);
and U7076 (N_7076,N_6923,N_7002);
or U7077 (N_7077,N_6976,N_6948);
xor U7078 (N_7078,N_6897,N_6892);
or U7079 (N_7079,N_6965,N_6958);
nand U7080 (N_7080,N_6924,N_6887);
xnor U7081 (N_7081,N_7003,N_6964);
or U7082 (N_7082,N_6915,N_7007);
and U7083 (N_7083,N_6994,N_6921);
xnor U7084 (N_7084,N_7036,N_6934);
nand U7085 (N_7085,N_6883,N_6982);
nor U7086 (N_7086,N_7016,N_6959);
or U7087 (N_7087,N_6916,N_6899);
nand U7088 (N_7088,N_6922,N_7029);
nand U7089 (N_7089,N_6908,N_7012);
or U7090 (N_7090,N_7033,N_6941);
and U7091 (N_7091,N_6996,N_6917);
xor U7092 (N_7092,N_7025,N_7021);
and U7093 (N_7093,N_6913,N_6911);
nor U7094 (N_7094,N_6975,N_6985);
xnor U7095 (N_7095,N_6890,N_6962);
or U7096 (N_7096,N_6895,N_6882);
or U7097 (N_7097,N_6973,N_7032);
nor U7098 (N_7098,N_6980,N_6989);
nand U7099 (N_7099,N_6961,N_6901);
xnor U7100 (N_7100,N_6903,N_6940);
nor U7101 (N_7101,N_6974,N_7027);
or U7102 (N_7102,N_6978,N_6972);
xnor U7103 (N_7103,N_6951,N_6963);
nand U7104 (N_7104,N_6880,N_6979);
and U7105 (N_7105,N_7035,N_6914);
xor U7106 (N_7106,N_6984,N_7005);
nand U7107 (N_7107,N_6925,N_7011);
nor U7108 (N_7108,N_7039,N_6987);
xnor U7109 (N_7109,N_6991,N_6910);
xor U7110 (N_7110,N_6988,N_6936);
nor U7111 (N_7111,N_6933,N_7034);
or U7112 (N_7112,N_6981,N_6956);
nor U7113 (N_7113,N_6900,N_6920);
xnor U7114 (N_7114,N_6927,N_6885);
xnor U7115 (N_7115,N_6949,N_6939);
nor U7116 (N_7116,N_6952,N_6950);
nand U7117 (N_7117,N_7020,N_6942);
and U7118 (N_7118,N_6904,N_6945);
or U7119 (N_7119,N_6992,N_6954);
nor U7120 (N_7120,N_7035,N_6909);
xnor U7121 (N_7121,N_7014,N_6997);
nor U7122 (N_7122,N_6905,N_7032);
and U7123 (N_7123,N_6954,N_6900);
nor U7124 (N_7124,N_7016,N_6918);
nor U7125 (N_7125,N_7015,N_6881);
xor U7126 (N_7126,N_6919,N_6913);
xor U7127 (N_7127,N_7008,N_6973);
xnor U7128 (N_7128,N_6919,N_6895);
or U7129 (N_7129,N_6904,N_7020);
nand U7130 (N_7130,N_6923,N_6901);
xor U7131 (N_7131,N_6927,N_6979);
nor U7132 (N_7132,N_6982,N_6993);
xnor U7133 (N_7133,N_6911,N_6977);
nor U7134 (N_7134,N_6941,N_6984);
nand U7135 (N_7135,N_6979,N_6973);
xnor U7136 (N_7136,N_6939,N_7014);
or U7137 (N_7137,N_6936,N_6922);
xor U7138 (N_7138,N_6934,N_7027);
or U7139 (N_7139,N_6895,N_6980);
xnor U7140 (N_7140,N_7034,N_6939);
or U7141 (N_7141,N_6918,N_6922);
nor U7142 (N_7142,N_6985,N_6951);
nor U7143 (N_7143,N_7031,N_6901);
or U7144 (N_7144,N_6978,N_7013);
xnor U7145 (N_7145,N_6888,N_7021);
or U7146 (N_7146,N_6980,N_6887);
and U7147 (N_7147,N_6924,N_6902);
nand U7148 (N_7148,N_6913,N_7030);
xnor U7149 (N_7149,N_6973,N_6995);
or U7150 (N_7150,N_6939,N_6989);
nand U7151 (N_7151,N_6899,N_6895);
nor U7152 (N_7152,N_6975,N_6894);
xor U7153 (N_7153,N_6951,N_6924);
nand U7154 (N_7154,N_6931,N_7021);
nand U7155 (N_7155,N_7039,N_6977);
xnor U7156 (N_7156,N_6975,N_6908);
and U7157 (N_7157,N_7020,N_6946);
nand U7158 (N_7158,N_6891,N_6895);
nand U7159 (N_7159,N_7004,N_6947);
and U7160 (N_7160,N_6912,N_7033);
nor U7161 (N_7161,N_6930,N_6906);
or U7162 (N_7162,N_6884,N_6927);
and U7163 (N_7163,N_6895,N_7027);
xor U7164 (N_7164,N_6886,N_6893);
and U7165 (N_7165,N_7004,N_6917);
nand U7166 (N_7166,N_6933,N_6997);
nor U7167 (N_7167,N_7005,N_6968);
nor U7168 (N_7168,N_6946,N_6965);
or U7169 (N_7169,N_6894,N_6919);
nand U7170 (N_7170,N_6903,N_6966);
xnor U7171 (N_7171,N_7039,N_6971);
or U7172 (N_7172,N_6905,N_6931);
nand U7173 (N_7173,N_6970,N_6917);
nor U7174 (N_7174,N_6962,N_6968);
and U7175 (N_7175,N_6934,N_6991);
nand U7176 (N_7176,N_6885,N_6992);
and U7177 (N_7177,N_6924,N_7022);
and U7178 (N_7178,N_6894,N_6986);
and U7179 (N_7179,N_6991,N_6976);
xnor U7180 (N_7180,N_7001,N_6951);
and U7181 (N_7181,N_6888,N_7029);
nand U7182 (N_7182,N_6977,N_7003);
nand U7183 (N_7183,N_6984,N_6983);
and U7184 (N_7184,N_7001,N_6931);
nand U7185 (N_7185,N_7018,N_6880);
nand U7186 (N_7186,N_6896,N_6997);
and U7187 (N_7187,N_6910,N_6938);
nand U7188 (N_7188,N_6902,N_7035);
nand U7189 (N_7189,N_6890,N_7009);
or U7190 (N_7190,N_7016,N_6953);
nor U7191 (N_7191,N_6960,N_6972);
nand U7192 (N_7192,N_6894,N_7030);
nand U7193 (N_7193,N_6957,N_7033);
xor U7194 (N_7194,N_6959,N_6916);
nand U7195 (N_7195,N_6961,N_6988);
or U7196 (N_7196,N_6994,N_6965);
and U7197 (N_7197,N_6912,N_6993);
nor U7198 (N_7198,N_6973,N_6976);
xor U7199 (N_7199,N_6886,N_6966);
xnor U7200 (N_7200,N_7047,N_7192);
xnor U7201 (N_7201,N_7165,N_7116);
nand U7202 (N_7202,N_7119,N_7118);
nor U7203 (N_7203,N_7058,N_7050);
or U7204 (N_7204,N_7042,N_7114);
or U7205 (N_7205,N_7115,N_7189);
nor U7206 (N_7206,N_7158,N_7105);
and U7207 (N_7207,N_7187,N_7132);
and U7208 (N_7208,N_7057,N_7078);
and U7209 (N_7209,N_7134,N_7153);
nor U7210 (N_7210,N_7081,N_7088);
xor U7211 (N_7211,N_7087,N_7100);
nor U7212 (N_7212,N_7083,N_7131);
or U7213 (N_7213,N_7113,N_7090);
nand U7214 (N_7214,N_7043,N_7107);
and U7215 (N_7215,N_7154,N_7091);
xnor U7216 (N_7216,N_7164,N_7161);
xor U7217 (N_7217,N_7190,N_7052);
nor U7218 (N_7218,N_7186,N_7085);
and U7219 (N_7219,N_7102,N_7096);
nand U7220 (N_7220,N_7146,N_7097);
nand U7221 (N_7221,N_7143,N_7059);
and U7222 (N_7222,N_7053,N_7129);
nor U7223 (N_7223,N_7137,N_7159);
nor U7224 (N_7224,N_7140,N_7147);
and U7225 (N_7225,N_7193,N_7183);
nand U7226 (N_7226,N_7169,N_7051);
nor U7227 (N_7227,N_7124,N_7080);
nand U7228 (N_7228,N_7125,N_7196);
or U7229 (N_7229,N_7150,N_7139);
xor U7230 (N_7230,N_7086,N_7198);
or U7231 (N_7231,N_7064,N_7110);
or U7232 (N_7232,N_7095,N_7151);
xnor U7233 (N_7233,N_7055,N_7197);
and U7234 (N_7234,N_7104,N_7041);
nor U7235 (N_7235,N_7121,N_7166);
or U7236 (N_7236,N_7077,N_7112);
xnor U7237 (N_7237,N_7123,N_7120);
and U7238 (N_7238,N_7070,N_7176);
and U7239 (N_7239,N_7101,N_7093);
nor U7240 (N_7240,N_7054,N_7109);
xnor U7241 (N_7241,N_7149,N_7184);
nand U7242 (N_7242,N_7128,N_7069);
and U7243 (N_7243,N_7049,N_7062);
nand U7244 (N_7244,N_7170,N_7127);
nand U7245 (N_7245,N_7060,N_7067);
and U7246 (N_7246,N_7180,N_7122);
and U7247 (N_7247,N_7181,N_7136);
nand U7248 (N_7248,N_7163,N_7174);
nor U7249 (N_7249,N_7156,N_7108);
and U7250 (N_7250,N_7065,N_7084);
nor U7251 (N_7251,N_7040,N_7175);
xor U7252 (N_7252,N_7182,N_7160);
and U7253 (N_7253,N_7076,N_7074);
and U7254 (N_7254,N_7138,N_7117);
or U7255 (N_7255,N_7194,N_7191);
and U7256 (N_7256,N_7092,N_7098);
or U7257 (N_7257,N_7073,N_7148);
and U7258 (N_7258,N_7168,N_7066);
nand U7259 (N_7259,N_7071,N_7142);
and U7260 (N_7260,N_7171,N_7172);
and U7261 (N_7261,N_7173,N_7144);
nor U7262 (N_7262,N_7167,N_7046);
and U7263 (N_7263,N_7068,N_7135);
or U7264 (N_7264,N_7126,N_7195);
nand U7265 (N_7265,N_7082,N_7072);
or U7266 (N_7266,N_7079,N_7188);
xnor U7267 (N_7267,N_7177,N_7179);
xnor U7268 (N_7268,N_7152,N_7162);
nand U7269 (N_7269,N_7048,N_7061);
or U7270 (N_7270,N_7178,N_7106);
and U7271 (N_7271,N_7044,N_7063);
xnor U7272 (N_7272,N_7133,N_7045);
and U7273 (N_7273,N_7094,N_7075);
and U7274 (N_7274,N_7056,N_7089);
nand U7275 (N_7275,N_7199,N_7185);
nor U7276 (N_7276,N_7145,N_7130);
xnor U7277 (N_7277,N_7155,N_7103);
xor U7278 (N_7278,N_7099,N_7141);
and U7279 (N_7279,N_7157,N_7111);
or U7280 (N_7280,N_7114,N_7173);
nand U7281 (N_7281,N_7144,N_7107);
and U7282 (N_7282,N_7112,N_7080);
or U7283 (N_7283,N_7126,N_7159);
nor U7284 (N_7284,N_7124,N_7197);
nor U7285 (N_7285,N_7066,N_7079);
nand U7286 (N_7286,N_7178,N_7046);
and U7287 (N_7287,N_7154,N_7069);
nor U7288 (N_7288,N_7131,N_7087);
or U7289 (N_7289,N_7161,N_7146);
or U7290 (N_7290,N_7106,N_7088);
and U7291 (N_7291,N_7151,N_7108);
nand U7292 (N_7292,N_7185,N_7195);
or U7293 (N_7293,N_7129,N_7185);
or U7294 (N_7294,N_7099,N_7086);
and U7295 (N_7295,N_7065,N_7154);
or U7296 (N_7296,N_7097,N_7193);
nor U7297 (N_7297,N_7068,N_7107);
xor U7298 (N_7298,N_7055,N_7109);
and U7299 (N_7299,N_7189,N_7093);
nand U7300 (N_7300,N_7100,N_7102);
or U7301 (N_7301,N_7093,N_7120);
xor U7302 (N_7302,N_7108,N_7123);
nor U7303 (N_7303,N_7140,N_7093);
or U7304 (N_7304,N_7129,N_7158);
xor U7305 (N_7305,N_7106,N_7167);
and U7306 (N_7306,N_7115,N_7050);
or U7307 (N_7307,N_7111,N_7112);
xor U7308 (N_7308,N_7094,N_7141);
or U7309 (N_7309,N_7190,N_7108);
or U7310 (N_7310,N_7064,N_7087);
xor U7311 (N_7311,N_7156,N_7078);
nand U7312 (N_7312,N_7140,N_7179);
and U7313 (N_7313,N_7067,N_7109);
and U7314 (N_7314,N_7186,N_7105);
and U7315 (N_7315,N_7105,N_7174);
nor U7316 (N_7316,N_7117,N_7104);
and U7317 (N_7317,N_7069,N_7111);
and U7318 (N_7318,N_7194,N_7066);
or U7319 (N_7319,N_7123,N_7073);
xnor U7320 (N_7320,N_7095,N_7058);
nor U7321 (N_7321,N_7061,N_7153);
or U7322 (N_7322,N_7071,N_7083);
xor U7323 (N_7323,N_7188,N_7150);
xor U7324 (N_7324,N_7187,N_7182);
xnor U7325 (N_7325,N_7052,N_7130);
nor U7326 (N_7326,N_7150,N_7192);
nand U7327 (N_7327,N_7187,N_7103);
xor U7328 (N_7328,N_7095,N_7176);
nor U7329 (N_7329,N_7053,N_7052);
nor U7330 (N_7330,N_7101,N_7196);
and U7331 (N_7331,N_7180,N_7189);
or U7332 (N_7332,N_7192,N_7054);
nor U7333 (N_7333,N_7198,N_7110);
xnor U7334 (N_7334,N_7187,N_7129);
and U7335 (N_7335,N_7178,N_7056);
and U7336 (N_7336,N_7145,N_7183);
xor U7337 (N_7337,N_7142,N_7093);
xor U7338 (N_7338,N_7137,N_7108);
or U7339 (N_7339,N_7110,N_7196);
xnor U7340 (N_7340,N_7171,N_7084);
xor U7341 (N_7341,N_7109,N_7121);
nand U7342 (N_7342,N_7171,N_7071);
nand U7343 (N_7343,N_7195,N_7081);
nand U7344 (N_7344,N_7082,N_7073);
or U7345 (N_7345,N_7100,N_7086);
xnor U7346 (N_7346,N_7040,N_7188);
xnor U7347 (N_7347,N_7049,N_7055);
nand U7348 (N_7348,N_7192,N_7120);
and U7349 (N_7349,N_7176,N_7197);
and U7350 (N_7350,N_7076,N_7160);
nand U7351 (N_7351,N_7179,N_7185);
nand U7352 (N_7352,N_7124,N_7061);
or U7353 (N_7353,N_7172,N_7083);
nor U7354 (N_7354,N_7198,N_7126);
nand U7355 (N_7355,N_7091,N_7114);
or U7356 (N_7356,N_7064,N_7080);
nor U7357 (N_7357,N_7113,N_7083);
or U7358 (N_7358,N_7189,N_7083);
nor U7359 (N_7359,N_7184,N_7138);
nor U7360 (N_7360,N_7200,N_7274);
nand U7361 (N_7361,N_7245,N_7356);
xor U7362 (N_7362,N_7268,N_7244);
xnor U7363 (N_7363,N_7202,N_7340);
or U7364 (N_7364,N_7270,N_7276);
xnor U7365 (N_7365,N_7309,N_7290);
xnor U7366 (N_7366,N_7346,N_7288);
xor U7367 (N_7367,N_7249,N_7242);
or U7368 (N_7368,N_7211,N_7329);
and U7369 (N_7369,N_7218,N_7205);
nand U7370 (N_7370,N_7206,N_7338);
nor U7371 (N_7371,N_7286,N_7332);
or U7372 (N_7372,N_7252,N_7303);
and U7373 (N_7373,N_7267,N_7330);
and U7374 (N_7374,N_7289,N_7231);
xnor U7375 (N_7375,N_7307,N_7259);
and U7376 (N_7376,N_7347,N_7285);
xor U7377 (N_7377,N_7335,N_7209);
and U7378 (N_7378,N_7357,N_7263);
nor U7379 (N_7379,N_7339,N_7327);
and U7380 (N_7380,N_7217,N_7308);
nor U7381 (N_7381,N_7243,N_7254);
nand U7382 (N_7382,N_7251,N_7240);
or U7383 (N_7383,N_7279,N_7241);
nand U7384 (N_7384,N_7260,N_7219);
or U7385 (N_7385,N_7345,N_7204);
and U7386 (N_7386,N_7287,N_7325);
xnor U7387 (N_7387,N_7220,N_7277);
nand U7388 (N_7388,N_7355,N_7300);
or U7389 (N_7389,N_7296,N_7248);
xnor U7390 (N_7390,N_7358,N_7229);
xor U7391 (N_7391,N_7269,N_7341);
xor U7392 (N_7392,N_7232,N_7225);
xor U7393 (N_7393,N_7328,N_7237);
nand U7394 (N_7394,N_7230,N_7273);
nor U7395 (N_7395,N_7224,N_7250);
nand U7396 (N_7396,N_7344,N_7334);
or U7397 (N_7397,N_7236,N_7313);
or U7398 (N_7398,N_7283,N_7320);
and U7399 (N_7399,N_7226,N_7203);
or U7400 (N_7400,N_7350,N_7256);
xor U7401 (N_7401,N_7323,N_7280);
nand U7402 (N_7402,N_7297,N_7216);
or U7403 (N_7403,N_7312,N_7291);
or U7404 (N_7404,N_7352,N_7266);
xnor U7405 (N_7405,N_7223,N_7299);
or U7406 (N_7406,N_7333,N_7239);
and U7407 (N_7407,N_7318,N_7302);
or U7408 (N_7408,N_7305,N_7306);
and U7409 (N_7409,N_7262,N_7301);
nor U7410 (N_7410,N_7258,N_7348);
nor U7411 (N_7411,N_7214,N_7233);
nor U7412 (N_7412,N_7342,N_7343);
or U7413 (N_7413,N_7227,N_7351);
or U7414 (N_7414,N_7294,N_7261);
nand U7415 (N_7415,N_7264,N_7278);
xor U7416 (N_7416,N_7271,N_7293);
and U7417 (N_7417,N_7322,N_7272);
xor U7418 (N_7418,N_7235,N_7215);
nand U7419 (N_7419,N_7321,N_7295);
and U7420 (N_7420,N_7255,N_7228);
nand U7421 (N_7421,N_7292,N_7221);
or U7422 (N_7422,N_7238,N_7275);
xnor U7423 (N_7423,N_7208,N_7284);
and U7424 (N_7424,N_7311,N_7201);
nand U7425 (N_7425,N_7310,N_7212);
nor U7426 (N_7426,N_7317,N_7349);
and U7427 (N_7427,N_7304,N_7234);
and U7428 (N_7428,N_7210,N_7265);
nand U7429 (N_7429,N_7281,N_7316);
or U7430 (N_7430,N_7337,N_7319);
xor U7431 (N_7431,N_7326,N_7298);
nand U7432 (N_7432,N_7314,N_7331);
nand U7433 (N_7433,N_7246,N_7207);
xnor U7434 (N_7434,N_7247,N_7282);
and U7435 (N_7435,N_7222,N_7253);
nand U7436 (N_7436,N_7213,N_7257);
nand U7437 (N_7437,N_7324,N_7353);
or U7438 (N_7438,N_7359,N_7315);
xnor U7439 (N_7439,N_7354,N_7336);
or U7440 (N_7440,N_7230,N_7291);
and U7441 (N_7441,N_7233,N_7242);
nand U7442 (N_7442,N_7248,N_7285);
or U7443 (N_7443,N_7245,N_7255);
and U7444 (N_7444,N_7329,N_7241);
and U7445 (N_7445,N_7323,N_7213);
nor U7446 (N_7446,N_7295,N_7269);
or U7447 (N_7447,N_7227,N_7225);
nor U7448 (N_7448,N_7310,N_7341);
xor U7449 (N_7449,N_7325,N_7294);
nor U7450 (N_7450,N_7308,N_7303);
and U7451 (N_7451,N_7294,N_7300);
nor U7452 (N_7452,N_7254,N_7342);
xor U7453 (N_7453,N_7275,N_7256);
xor U7454 (N_7454,N_7355,N_7330);
and U7455 (N_7455,N_7274,N_7222);
nor U7456 (N_7456,N_7209,N_7306);
nor U7457 (N_7457,N_7359,N_7231);
xnor U7458 (N_7458,N_7247,N_7356);
xor U7459 (N_7459,N_7310,N_7269);
xor U7460 (N_7460,N_7282,N_7201);
xnor U7461 (N_7461,N_7315,N_7218);
or U7462 (N_7462,N_7354,N_7207);
xnor U7463 (N_7463,N_7333,N_7220);
or U7464 (N_7464,N_7287,N_7241);
nand U7465 (N_7465,N_7320,N_7227);
xnor U7466 (N_7466,N_7230,N_7298);
xnor U7467 (N_7467,N_7270,N_7213);
or U7468 (N_7468,N_7341,N_7318);
or U7469 (N_7469,N_7346,N_7314);
nor U7470 (N_7470,N_7242,N_7317);
xnor U7471 (N_7471,N_7357,N_7281);
nor U7472 (N_7472,N_7334,N_7217);
or U7473 (N_7473,N_7220,N_7219);
and U7474 (N_7474,N_7341,N_7257);
xnor U7475 (N_7475,N_7235,N_7308);
xor U7476 (N_7476,N_7265,N_7204);
or U7477 (N_7477,N_7282,N_7333);
xnor U7478 (N_7478,N_7306,N_7217);
or U7479 (N_7479,N_7284,N_7297);
or U7480 (N_7480,N_7215,N_7357);
nand U7481 (N_7481,N_7256,N_7228);
nand U7482 (N_7482,N_7313,N_7327);
nor U7483 (N_7483,N_7346,N_7204);
nand U7484 (N_7484,N_7331,N_7240);
and U7485 (N_7485,N_7319,N_7244);
nor U7486 (N_7486,N_7290,N_7231);
and U7487 (N_7487,N_7300,N_7323);
or U7488 (N_7488,N_7304,N_7239);
and U7489 (N_7489,N_7229,N_7200);
nand U7490 (N_7490,N_7304,N_7337);
or U7491 (N_7491,N_7256,N_7322);
and U7492 (N_7492,N_7317,N_7215);
and U7493 (N_7493,N_7349,N_7355);
xor U7494 (N_7494,N_7207,N_7333);
nor U7495 (N_7495,N_7239,N_7237);
xnor U7496 (N_7496,N_7279,N_7218);
xor U7497 (N_7497,N_7345,N_7258);
or U7498 (N_7498,N_7248,N_7244);
nand U7499 (N_7499,N_7267,N_7247);
or U7500 (N_7500,N_7203,N_7349);
or U7501 (N_7501,N_7305,N_7238);
nand U7502 (N_7502,N_7277,N_7263);
nand U7503 (N_7503,N_7251,N_7215);
xnor U7504 (N_7504,N_7213,N_7214);
or U7505 (N_7505,N_7263,N_7354);
xnor U7506 (N_7506,N_7210,N_7216);
nand U7507 (N_7507,N_7247,N_7309);
nor U7508 (N_7508,N_7234,N_7204);
or U7509 (N_7509,N_7295,N_7207);
nor U7510 (N_7510,N_7321,N_7244);
xnor U7511 (N_7511,N_7271,N_7315);
nand U7512 (N_7512,N_7340,N_7244);
xnor U7513 (N_7513,N_7226,N_7281);
nor U7514 (N_7514,N_7287,N_7229);
nand U7515 (N_7515,N_7312,N_7304);
and U7516 (N_7516,N_7357,N_7312);
or U7517 (N_7517,N_7345,N_7237);
and U7518 (N_7518,N_7250,N_7267);
nand U7519 (N_7519,N_7314,N_7309);
nand U7520 (N_7520,N_7441,N_7493);
nand U7521 (N_7521,N_7404,N_7508);
nand U7522 (N_7522,N_7382,N_7462);
or U7523 (N_7523,N_7423,N_7427);
and U7524 (N_7524,N_7385,N_7371);
xnor U7525 (N_7525,N_7367,N_7391);
xnor U7526 (N_7526,N_7512,N_7454);
nor U7527 (N_7527,N_7417,N_7504);
nand U7528 (N_7528,N_7510,N_7463);
xor U7529 (N_7529,N_7437,N_7414);
nand U7530 (N_7530,N_7482,N_7401);
and U7531 (N_7531,N_7449,N_7383);
xor U7532 (N_7532,N_7519,N_7509);
and U7533 (N_7533,N_7489,N_7416);
and U7534 (N_7534,N_7459,N_7502);
nor U7535 (N_7535,N_7490,N_7472);
and U7536 (N_7536,N_7430,N_7448);
xnor U7537 (N_7537,N_7458,N_7363);
nor U7538 (N_7538,N_7403,N_7365);
nand U7539 (N_7539,N_7439,N_7473);
or U7540 (N_7540,N_7484,N_7507);
or U7541 (N_7541,N_7491,N_7506);
nand U7542 (N_7542,N_7480,N_7460);
nand U7543 (N_7543,N_7488,N_7372);
and U7544 (N_7544,N_7445,N_7466);
or U7545 (N_7545,N_7438,N_7501);
nor U7546 (N_7546,N_7399,N_7373);
and U7547 (N_7547,N_7440,N_7486);
or U7548 (N_7548,N_7494,N_7408);
nor U7549 (N_7549,N_7377,N_7413);
nand U7550 (N_7550,N_7431,N_7406);
nand U7551 (N_7551,N_7456,N_7511);
nand U7552 (N_7552,N_7468,N_7495);
and U7553 (N_7553,N_7360,N_7361);
and U7554 (N_7554,N_7478,N_7443);
or U7555 (N_7555,N_7470,N_7422);
nor U7556 (N_7556,N_7464,N_7487);
xor U7557 (N_7557,N_7492,N_7398);
xnor U7558 (N_7558,N_7496,N_7387);
nor U7559 (N_7559,N_7412,N_7469);
and U7560 (N_7560,N_7393,N_7379);
xnor U7561 (N_7561,N_7499,N_7410);
nand U7562 (N_7562,N_7479,N_7375);
and U7563 (N_7563,N_7447,N_7369);
nand U7564 (N_7564,N_7515,N_7518);
xnor U7565 (N_7565,N_7517,N_7436);
or U7566 (N_7566,N_7368,N_7514);
nor U7567 (N_7567,N_7396,N_7505);
and U7568 (N_7568,N_7381,N_7394);
nand U7569 (N_7569,N_7389,N_7402);
nand U7570 (N_7570,N_7435,N_7446);
nand U7571 (N_7571,N_7380,N_7429);
or U7572 (N_7572,N_7444,N_7420);
nand U7573 (N_7573,N_7467,N_7366);
and U7574 (N_7574,N_7451,N_7483);
nand U7575 (N_7575,N_7400,N_7453);
or U7576 (N_7576,N_7485,N_7471);
and U7577 (N_7577,N_7418,N_7513);
nor U7578 (N_7578,N_7409,N_7461);
nor U7579 (N_7579,N_7407,N_7474);
nand U7580 (N_7580,N_7364,N_7498);
or U7581 (N_7581,N_7397,N_7433);
nand U7582 (N_7582,N_7450,N_7421);
nor U7583 (N_7583,N_7476,N_7386);
nor U7584 (N_7584,N_7475,N_7442);
or U7585 (N_7585,N_7395,N_7411);
xor U7586 (N_7586,N_7415,N_7434);
or U7587 (N_7587,N_7465,N_7384);
nand U7588 (N_7588,N_7405,N_7500);
nor U7589 (N_7589,N_7497,N_7362);
xor U7590 (N_7590,N_7392,N_7455);
and U7591 (N_7591,N_7426,N_7378);
and U7592 (N_7592,N_7370,N_7390);
xor U7593 (N_7593,N_7457,N_7516);
nor U7594 (N_7594,N_7419,N_7503);
nor U7595 (N_7595,N_7376,N_7432);
xnor U7596 (N_7596,N_7428,N_7374);
xor U7597 (N_7597,N_7388,N_7477);
nor U7598 (N_7598,N_7424,N_7425);
nand U7599 (N_7599,N_7481,N_7452);
or U7600 (N_7600,N_7390,N_7360);
nor U7601 (N_7601,N_7424,N_7518);
xor U7602 (N_7602,N_7448,N_7420);
or U7603 (N_7603,N_7507,N_7467);
nand U7604 (N_7604,N_7484,N_7491);
nor U7605 (N_7605,N_7361,N_7403);
or U7606 (N_7606,N_7452,N_7482);
nand U7607 (N_7607,N_7419,N_7440);
or U7608 (N_7608,N_7422,N_7455);
nand U7609 (N_7609,N_7453,N_7491);
nand U7610 (N_7610,N_7511,N_7487);
or U7611 (N_7611,N_7510,N_7365);
and U7612 (N_7612,N_7419,N_7505);
or U7613 (N_7613,N_7408,N_7389);
nor U7614 (N_7614,N_7513,N_7482);
and U7615 (N_7615,N_7487,N_7417);
nor U7616 (N_7616,N_7502,N_7449);
and U7617 (N_7617,N_7416,N_7498);
nor U7618 (N_7618,N_7409,N_7440);
nand U7619 (N_7619,N_7405,N_7404);
nand U7620 (N_7620,N_7455,N_7402);
xnor U7621 (N_7621,N_7502,N_7446);
nor U7622 (N_7622,N_7472,N_7503);
nor U7623 (N_7623,N_7377,N_7373);
xor U7624 (N_7624,N_7506,N_7379);
nor U7625 (N_7625,N_7424,N_7396);
nand U7626 (N_7626,N_7469,N_7363);
nand U7627 (N_7627,N_7500,N_7415);
xnor U7628 (N_7628,N_7489,N_7444);
nand U7629 (N_7629,N_7386,N_7498);
nor U7630 (N_7630,N_7372,N_7367);
and U7631 (N_7631,N_7381,N_7453);
nor U7632 (N_7632,N_7481,N_7416);
and U7633 (N_7633,N_7476,N_7465);
nor U7634 (N_7634,N_7517,N_7495);
or U7635 (N_7635,N_7400,N_7478);
and U7636 (N_7636,N_7474,N_7367);
nor U7637 (N_7637,N_7399,N_7409);
or U7638 (N_7638,N_7496,N_7367);
xor U7639 (N_7639,N_7428,N_7507);
xor U7640 (N_7640,N_7492,N_7455);
nor U7641 (N_7641,N_7415,N_7423);
nand U7642 (N_7642,N_7384,N_7397);
nand U7643 (N_7643,N_7514,N_7510);
nand U7644 (N_7644,N_7372,N_7407);
and U7645 (N_7645,N_7494,N_7418);
xnor U7646 (N_7646,N_7481,N_7379);
nor U7647 (N_7647,N_7511,N_7378);
nand U7648 (N_7648,N_7373,N_7364);
or U7649 (N_7649,N_7498,N_7508);
and U7650 (N_7650,N_7466,N_7483);
xnor U7651 (N_7651,N_7405,N_7481);
or U7652 (N_7652,N_7444,N_7495);
nand U7653 (N_7653,N_7485,N_7500);
and U7654 (N_7654,N_7385,N_7475);
xnor U7655 (N_7655,N_7505,N_7479);
xor U7656 (N_7656,N_7395,N_7469);
nor U7657 (N_7657,N_7389,N_7426);
xnor U7658 (N_7658,N_7477,N_7515);
nand U7659 (N_7659,N_7438,N_7389);
nand U7660 (N_7660,N_7393,N_7362);
and U7661 (N_7661,N_7451,N_7492);
and U7662 (N_7662,N_7474,N_7511);
nor U7663 (N_7663,N_7430,N_7489);
nor U7664 (N_7664,N_7435,N_7388);
xor U7665 (N_7665,N_7479,N_7460);
nor U7666 (N_7666,N_7450,N_7514);
nor U7667 (N_7667,N_7471,N_7370);
nor U7668 (N_7668,N_7419,N_7513);
xor U7669 (N_7669,N_7506,N_7512);
xor U7670 (N_7670,N_7374,N_7481);
and U7671 (N_7671,N_7388,N_7395);
nand U7672 (N_7672,N_7364,N_7454);
nand U7673 (N_7673,N_7413,N_7428);
nor U7674 (N_7674,N_7413,N_7448);
or U7675 (N_7675,N_7392,N_7441);
xnor U7676 (N_7676,N_7459,N_7460);
xor U7677 (N_7677,N_7474,N_7433);
nand U7678 (N_7678,N_7421,N_7395);
xnor U7679 (N_7679,N_7497,N_7405);
and U7680 (N_7680,N_7617,N_7586);
nor U7681 (N_7681,N_7592,N_7608);
xor U7682 (N_7682,N_7645,N_7593);
nand U7683 (N_7683,N_7648,N_7647);
nor U7684 (N_7684,N_7570,N_7659);
xor U7685 (N_7685,N_7676,N_7611);
and U7686 (N_7686,N_7587,N_7563);
or U7687 (N_7687,N_7523,N_7591);
xor U7688 (N_7688,N_7534,N_7664);
nor U7689 (N_7689,N_7636,N_7671);
xor U7690 (N_7690,N_7546,N_7521);
and U7691 (N_7691,N_7656,N_7569);
and U7692 (N_7692,N_7652,N_7595);
nand U7693 (N_7693,N_7579,N_7522);
or U7694 (N_7694,N_7643,N_7633);
or U7695 (N_7695,N_7594,N_7582);
and U7696 (N_7696,N_7529,N_7638);
and U7697 (N_7697,N_7547,N_7675);
and U7698 (N_7698,N_7628,N_7631);
nand U7699 (N_7699,N_7604,N_7666);
and U7700 (N_7700,N_7558,N_7613);
xnor U7701 (N_7701,N_7630,N_7574);
or U7702 (N_7702,N_7646,N_7642);
xor U7703 (N_7703,N_7560,N_7590);
and U7704 (N_7704,N_7549,N_7596);
and U7705 (N_7705,N_7532,N_7559);
and U7706 (N_7706,N_7557,N_7635);
or U7707 (N_7707,N_7620,N_7657);
nand U7708 (N_7708,N_7623,N_7577);
and U7709 (N_7709,N_7669,N_7580);
or U7710 (N_7710,N_7553,N_7562);
and U7711 (N_7711,N_7555,N_7545);
and U7712 (N_7712,N_7665,N_7629);
and U7713 (N_7713,N_7632,N_7542);
or U7714 (N_7714,N_7640,N_7539);
xor U7715 (N_7715,N_7637,N_7622);
nand U7716 (N_7716,N_7588,N_7520);
nand U7717 (N_7717,N_7634,N_7650);
nand U7718 (N_7718,N_7644,N_7544);
nand U7719 (N_7719,N_7653,N_7610);
nor U7720 (N_7720,N_7585,N_7679);
and U7721 (N_7721,N_7548,N_7605);
xnor U7722 (N_7722,N_7606,N_7609);
nand U7723 (N_7723,N_7537,N_7556);
nor U7724 (N_7724,N_7589,N_7526);
or U7725 (N_7725,N_7575,N_7552);
nor U7726 (N_7726,N_7541,N_7571);
xor U7727 (N_7727,N_7602,N_7576);
nor U7728 (N_7728,N_7619,N_7672);
nor U7729 (N_7729,N_7568,N_7538);
and U7730 (N_7730,N_7550,N_7627);
or U7731 (N_7731,N_7655,N_7599);
nor U7732 (N_7732,N_7658,N_7603);
nand U7733 (N_7733,N_7543,N_7615);
and U7734 (N_7734,N_7567,N_7662);
nand U7735 (N_7735,N_7535,N_7625);
and U7736 (N_7736,N_7536,N_7673);
nand U7737 (N_7737,N_7524,N_7601);
xor U7738 (N_7738,N_7573,N_7584);
nand U7739 (N_7739,N_7531,N_7641);
or U7740 (N_7740,N_7624,N_7581);
or U7741 (N_7741,N_7583,N_7614);
xor U7742 (N_7742,N_7572,N_7578);
nor U7743 (N_7743,N_7626,N_7551);
nand U7744 (N_7744,N_7660,N_7561);
and U7745 (N_7745,N_7663,N_7678);
xor U7746 (N_7746,N_7670,N_7667);
and U7747 (N_7747,N_7668,N_7533);
or U7748 (N_7748,N_7530,N_7618);
or U7749 (N_7749,N_7525,N_7528);
nor U7750 (N_7750,N_7564,N_7651);
nand U7751 (N_7751,N_7527,N_7621);
nor U7752 (N_7752,N_7639,N_7607);
or U7753 (N_7753,N_7661,N_7566);
or U7754 (N_7754,N_7674,N_7654);
and U7755 (N_7755,N_7540,N_7598);
or U7756 (N_7756,N_7597,N_7565);
xor U7757 (N_7757,N_7616,N_7649);
xor U7758 (N_7758,N_7600,N_7677);
nand U7759 (N_7759,N_7554,N_7612);
xnor U7760 (N_7760,N_7655,N_7583);
nand U7761 (N_7761,N_7536,N_7560);
xor U7762 (N_7762,N_7569,N_7595);
nand U7763 (N_7763,N_7602,N_7591);
and U7764 (N_7764,N_7628,N_7669);
nor U7765 (N_7765,N_7521,N_7566);
xnor U7766 (N_7766,N_7539,N_7563);
xor U7767 (N_7767,N_7621,N_7598);
and U7768 (N_7768,N_7666,N_7570);
and U7769 (N_7769,N_7629,N_7649);
or U7770 (N_7770,N_7565,N_7585);
xor U7771 (N_7771,N_7637,N_7671);
nand U7772 (N_7772,N_7571,N_7596);
nor U7773 (N_7773,N_7671,N_7583);
or U7774 (N_7774,N_7647,N_7623);
nor U7775 (N_7775,N_7628,N_7592);
nor U7776 (N_7776,N_7575,N_7678);
or U7777 (N_7777,N_7618,N_7562);
xor U7778 (N_7778,N_7551,N_7621);
or U7779 (N_7779,N_7582,N_7540);
and U7780 (N_7780,N_7672,N_7557);
nand U7781 (N_7781,N_7615,N_7535);
and U7782 (N_7782,N_7643,N_7525);
or U7783 (N_7783,N_7609,N_7654);
xnor U7784 (N_7784,N_7590,N_7624);
nor U7785 (N_7785,N_7532,N_7531);
and U7786 (N_7786,N_7537,N_7676);
nand U7787 (N_7787,N_7587,N_7637);
or U7788 (N_7788,N_7652,N_7614);
xnor U7789 (N_7789,N_7662,N_7590);
or U7790 (N_7790,N_7675,N_7539);
and U7791 (N_7791,N_7654,N_7636);
or U7792 (N_7792,N_7585,N_7560);
or U7793 (N_7793,N_7627,N_7596);
and U7794 (N_7794,N_7661,N_7574);
nand U7795 (N_7795,N_7654,N_7611);
or U7796 (N_7796,N_7593,N_7609);
and U7797 (N_7797,N_7573,N_7567);
nand U7798 (N_7798,N_7589,N_7670);
xor U7799 (N_7799,N_7525,N_7527);
nand U7800 (N_7800,N_7583,N_7600);
nor U7801 (N_7801,N_7662,N_7545);
or U7802 (N_7802,N_7625,N_7574);
nand U7803 (N_7803,N_7583,N_7650);
or U7804 (N_7804,N_7622,N_7607);
xor U7805 (N_7805,N_7586,N_7566);
nand U7806 (N_7806,N_7536,N_7579);
and U7807 (N_7807,N_7662,N_7633);
xnor U7808 (N_7808,N_7644,N_7584);
nand U7809 (N_7809,N_7578,N_7567);
nand U7810 (N_7810,N_7606,N_7627);
nor U7811 (N_7811,N_7576,N_7590);
or U7812 (N_7812,N_7642,N_7603);
xor U7813 (N_7813,N_7541,N_7624);
nor U7814 (N_7814,N_7603,N_7547);
nand U7815 (N_7815,N_7668,N_7576);
nand U7816 (N_7816,N_7552,N_7609);
and U7817 (N_7817,N_7645,N_7625);
nor U7818 (N_7818,N_7549,N_7644);
xor U7819 (N_7819,N_7599,N_7636);
nor U7820 (N_7820,N_7639,N_7621);
nand U7821 (N_7821,N_7577,N_7594);
or U7822 (N_7822,N_7566,N_7571);
and U7823 (N_7823,N_7625,N_7652);
nand U7824 (N_7824,N_7555,N_7534);
nand U7825 (N_7825,N_7591,N_7566);
nor U7826 (N_7826,N_7654,N_7638);
and U7827 (N_7827,N_7639,N_7622);
and U7828 (N_7828,N_7616,N_7544);
xnor U7829 (N_7829,N_7643,N_7553);
or U7830 (N_7830,N_7537,N_7580);
or U7831 (N_7831,N_7620,N_7582);
or U7832 (N_7832,N_7521,N_7589);
xor U7833 (N_7833,N_7526,N_7657);
nor U7834 (N_7834,N_7546,N_7602);
and U7835 (N_7835,N_7665,N_7569);
and U7836 (N_7836,N_7575,N_7606);
and U7837 (N_7837,N_7653,N_7580);
nand U7838 (N_7838,N_7547,N_7520);
nor U7839 (N_7839,N_7677,N_7542);
nand U7840 (N_7840,N_7720,N_7776);
and U7841 (N_7841,N_7725,N_7773);
nor U7842 (N_7842,N_7838,N_7811);
xor U7843 (N_7843,N_7692,N_7802);
and U7844 (N_7844,N_7785,N_7793);
or U7845 (N_7845,N_7835,N_7784);
or U7846 (N_7846,N_7822,N_7751);
nor U7847 (N_7847,N_7832,N_7742);
xor U7848 (N_7848,N_7775,N_7695);
xor U7849 (N_7849,N_7735,N_7709);
nor U7850 (N_7850,N_7801,N_7794);
xnor U7851 (N_7851,N_7824,N_7748);
nand U7852 (N_7852,N_7762,N_7791);
xnor U7853 (N_7853,N_7829,N_7701);
nor U7854 (N_7854,N_7781,N_7714);
xnor U7855 (N_7855,N_7739,N_7819);
and U7856 (N_7856,N_7733,N_7708);
xnor U7857 (N_7857,N_7715,N_7799);
nand U7858 (N_7858,N_7792,N_7753);
or U7859 (N_7859,N_7749,N_7833);
nor U7860 (N_7860,N_7731,N_7795);
and U7861 (N_7861,N_7745,N_7790);
xnor U7862 (N_7862,N_7780,N_7704);
and U7863 (N_7863,N_7828,N_7721);
nand U7864 (N_7864,N_7685,N_7681);
xor U7865 (N_7865,N_7724,N_7726);
xor U7866 (N_7866,N_7830,N_7746);
nor U7867 (N_7867,N_7750,N_7787);
and U7868 (N_7868,N_7728,N_7718);
nor U7869 (N_7869,N_7736,N_7688);
xnor U7870 (N_7870,N_7786,N_7820);
nor U7871 (N_7871,N_7810,N_7756);
nor U7872 (N_7872,N_7764,N_7823);
nor U7873 (N_7873,N_7686,N_7734);
and U7874 (N_7874,N_7818,N_7696);
or U7875 (N_7875,N_7796,N_7729);
nor U7876 (N_7876,N_7769,N_7767);
nor U7877 (N_7877,N_7682,N_7722);
xor U7878 (N_7878,N_7710,N_7763);
nor U7879 (N_7879,N_7683,N_7798);
xnor U7880 (N_7880,N_7740,N_7817);
nor U7881 (N_7881,N_7839,N_7768);
nor U7882 (N_7882,N_7737,N_7789);
nand U7883 (N_7883,N_7808,N_7698);
nand U7884 (N_7884,N_7788,N_7813);
and U7885 (N_7885,N_7706,N_7827);
nand U7886 (N_7886,N_7759,N_7691);
nand U7887 (N_7887,N_7754,N_7713);
and U7888 (N_7888,N_7719,N_7693);
and U7889 (N_7889,N_7804,N_7711);
nor U7890 (N_7890,N_7797,N_7752);
nor U7891 (N_7891,N_7765,N_7800);
nor U7892 (N_7892,N_7702,N_7717);
nand U7893 (N_7893,N_7744,N_7812);
xnor U7894 (N_7894,N_7803,N_7757);
xnor U7895 (N_7895,N_7684,N_7805);
nand U7896 (N_7896,N_7712,N_7747);
or U7897 (N_7897,N_7814,N_7716);
and U7898 (N_7898,N_7834,N_7816);
or U7899 (N_7899,N_7700,N_7727);
and U7900 (N_7900,N_7723,N_7836);
and U7901 (N_7901,N_7705,N_7831);
xnor U7902 (N_7902,N_7809,N_7821);
nor U7903 (N_7903,N_7690,N_7707);
or U7904 (N_7904,N_7783,N_7738);
nor U7905 (N_7905,N_7777,N_7779);
or U7906 (N_7906,N_7730,N_7699);
nand U7907 (N_7907,N_7770,N_7806);
or U7908 (N_7908,N_7703,N_7755);
or U7909 (N_7909,N_7778,N_7760);
and U7910 (N_7910,N_7732,N_7758);
xnor U7911 (N_7911,N_7694,N_7772);
xnor U7912 (N_7912,N_7697,N_7826);
and U7913 (N_7913,N_7782,N_7680);
or U7914 (N_7914,N_7689,N_7766);
or U7915 (N_7915,N_7807,N_7774);
nor U7916 (N_7916,N_7741,N_7743);
nor U7917 (N_7917,N_7687,N_7771);
xor U7918 (N_7918,N_7761,N_7837);
xnor U7919 (N_7919,N_7825,N_7815);
nand U7920 (N_7920,N_7757,N_7701);
and U7921 (N_7921,N_7705,N_7818);
nor U7922 (N_7922,N_7692,N_7768);
xnor U7923 (N_7923,N_7752,N_7760);
and U7924 (N_7924,N_7716,N_7746);
nor U7925 (N_7925,N_7767,N_7756);
nand U7926 (N_7926,N_7820,N_7739);
or U7927 (N_7927,N_7784,N_7786);
and U7928 (N_7928,N_7773,N_7805);
nor U7929 (N_7929,N_7692,N_7835);
or U7930 (N_7930,N_7767,N_7781);
nand U7931 (N_7931,N_7757,N_7795);
and U7932 (N_7932,N_7706,N_7715);
or U7933 (N_7933,N_7708,N_7830);
or U7934 (N_7934,N_7789,N_7837);
nor U7935 (N_7935,N_7684,N_7812);
nand U7936 (N_7936,N_7754,N_7727);
xnor U7937 (N_7937,N_7829,N_7762);
and U7938 (N_7938,N_7775,N_7764);
and U7939 (N_7939,N_7806,N_7813);
and U7940 (N_7940,N_7700,N_7760);
and U7941 (N_7941,N_7823,N_7711);
xor U7942 (N_7942,N_7736,N_7828);
and U7943 (N_7943,N_7811,N_7741);
nand U7944 (N_7944,N_7791,N_7782);
xnor U7945 (N_7945,N_7693,N_7755);
and U7946 (N_7946,N_7772,N_7711);
xnor U7947 (N_7947,N_7815,N_7726);
nand U7948 (N_7948,N_7763,N_7784);
xnor U7949 (N_7949,N_7708,N_7836);
nand U7950 (N_7950,N_7836,N_7817);
nand U7951 (N_7951,N_7754,N_7757);
and U7952 (N_7952,N_7756,N_7763);
nor U7953 (N_7953,N_7776,N_7696);
and U7954 (N_7954,N_7733,N_7692);
or U7955 (N_7955,N_7741,N_7824);
nand U7956 (N_7956,N_7785,N_7715);
or U7957 (N_7957,N_7796,N_7712);
nor U7958 (N_7958,N_7712,N_7691);
xor U7959 (N_7959,N_7773,N_7726);
nor U7960 (N_7960,N_7833,N_7781);
and U7961 (N_7961,N_7690,N_7836);
or U7962 (N_7962,N_7822,N_7746);
or U7963 (N_7963,N_7726,N_7781);
nand U7964 (N_7964,N_7703,N_7814);
nand U7965 (N_7965,N_7806,N_7753);
nor U7966 (N_7966,N_7781,N_7725);
xnor U7967 (N_7967,N_7706,N_7684);
or U7968 (N_7968,N_7783,N_7761);
nor U7969 (N_7969,N_7798,N_7772);
and U7970 (N_7970,N_7808,N_7791);
and U7971 (N_7971,N_7837,N_7749);
and U7972 (N_7972,N_7698,N_7701);
and U7973 (N_7973,N_7837,N_7685);
nor U7974 (N_7974,N_7749,N_7797);
and U7975 (N_7975,N_7730,N_7749);
nor U7976 (N_7976,N_7715,N_7729);
xor U7977 (N_7977,N_7794,N_7711);
or U7978 (N_7978,N_7825,N_7800);
or U7979 (N_7979,N_7720,N_7701);
and U7980 (N_7980,N_7828,N_7743);
and U7981 (N_7981,N_7767,N_7819);
or U7982 (N_7982,N_7824,N_7792);
and U7983 (N_7983,N_7702,N_7786);
or U7984 (N_7984,N_7802,N_7723);
xor U7985 (N_7985,N_7805,N_7807);
xnor U7986 (N_7986,N_7806,N_7757);
or U7987 (N_7987,N_7754,N_7735);
xnor U7988 (N_7988,N_7680,N_7730);
xnor U7989 (N_7989,N_7736,N_7723);
xor U7990 (N_7990,N_7752,N_7685);
nor U7991 (N_7991,N_7742,N_7758);
xor U7992 (N_7992,N_7801,N_7807);
or U7993 (N_7993,N_7792,N_7746);
xor U7994 (N_7994,N_7680,N_7733);
nand U7995 (N_7995,N_7732,N_7765);
or U7996 (N_7996,N_7737,N_7768);
or U7997 (N_7997,N_7790,N_7696);
nand U7998 (N_7998,N_7825,N_7799);
or U7999 (N_7999,N_7812,N_7816);
and U8000 (N_8000,N_7999,N_7994);
nor U8001 (N_8001,N_7908,N_7867);
nor U8002 (N_8002,N_7960,N_7866);
or U8003 (N_8003,N_7945,N_7876);
and U8004 (N_8004,N_7976,N_7861);
nand U8005 (N_8005,N_7844,N_7973);
or U8006 (N_8006,N_7899,N_7933);
or U8007 (N_8007,N_7874,N_7943);
and U8008 (N_8008,N_7845,N_7875);
nand U8009 (N_8009,N_7924,N_7935);
or U8010 (N_8010,N_7991,N_7920);
or U8011 (N_8011,N_7870,N_7891);
nor U8012 (N_8012,N_7909,N_7842);
nor U8013 (N_8013,N_7841,N_7941);
nor U8014 (N_8014,N_7938,N_7995);
and U8015 (N_8015,N_7864,N_7912);
nand U8016 (N_8016,N_7879,N_7902);
or U8017 (N_8017,N_7863,N_7982);
and U8018 (N_8018,N_7906,N_7974);
nor U8019 (N_8019,N_7884,N_7946);
xor U8020 (N_8020,N_7892,N_7926);
xor U8021 (N_8021,N_7948,N_7868);
or U8022 (N_8022,N_7860,N_7989);
and U8023 (N_8023,N_7971,N_7872);
nand U8024 (N_8024,N_7901,N_7966);
xor U8025 (N_8025,N_7852,N_7896);
nor U8026 (N_8026,N_7894,N_7882);
nor U8027 (N_8027,N_7987,N_7862);
and U8028 (N_8028,N_7956,N_7871);
xor U8029 (N_8029,N_7984,N_7880);
or U8030 (N_8030,N_7919,N_7877);
and U8031 (N_8031,N_7962,N_7923);
and U8032 (N_8032,N_7983,N_7903);
nor U8033 (N_8033,N_7859,N_7917);
nor U8034 (N_8034,N_7922,N_7843);
or U8035 (N_8035,N_7865,N_7972);
and U8036 (N_8036,N_7934,N_7889);
nor U8037 (N_8037,N_7952,N_7940);
or U8038 (N_8038,N_7975,N_7848);
nor U8039 (N_8039,N_7913,N_7890);
and U8040 (N_8040,N_7886,N_7961);
nand U8041 (N_8041,N_7929,N_7907);
xnor U8042 (N_8042,N_7897,N_7858);
or U8043 (N_8043,N_7905,N_7910);
nand U8044 (N_8044,N_7951,N_7996);
nor U8045 (N_8045,N_7887,N_7881);
and U8046 (N_8046,N_7992,N_7968);
xor U8047 (N_8047,N_7955,N_7979);
nand U8048 (N_8048,N_7965,N_7993);
nand U8049 (N_8049,N_7900,N_7853);
nand U8050 (N_8050,N_7854,N_7954);
nand U8051 (N_8051,N_7985,N_7883);
and U8052 (N_8052,N_7980,N_7998);
and U8053 (N_8053,N_7893,N_7847);
and U8054 (N_8054,N_7930,N_7953);
nor U8055 (N_8055,N_7914,N_7888);
nor U8056 (N_8056,N_7846,N_7958);
xor U8057 (N_8057,N_7895,N_7932);
xor U8058 (N_8058,N_7957,N_7925);
nand U8059 (N_8059,N_7851,N_7921);
nand U8060 (N_8060,N_7849,N_7850);
xor U8061 (N_8061,N_7970,N_7856);
and U8062 (N_8062,N_7857,N_7959);
nand U8063 (N_8063,N_7936,N_7931);
nor U8064 (N_8064,N_7918,N_7977);
nor U8065 (N_8065,N_7988,N_7916);
nand U8066 (N_8066,N_7878,N_7944);
or U8067 (N_8067,N_7942,N_7869);
nor U8068 (N_8068,N_7964,N_7840);
xnor U8069 (N_8069,N_7981,N_7997);
and U8070 (N_8070,N_7904,N_7963);
xnor U8071 (N_8071,N_7915,N_7947);
xor U8072 (N_8072,N_7990,N_7950);
xor U8073 (N_8073,N_7885,N_7986);
nand U8074 (N_8074,N_7949,N_7898);
nor U8075 (N_8075,N_7927,N_7978);
nand U8076 (N_8076,N_7939,N_7928);
nor U8077 (N_8077,N_7911,N_7873);
or U8078 (N_8078,N_7855,N_7969);
and U8079 (N_8079,N_7967,N_7937);
or U8080 (N_8080,N_7964,N_7963);
nor U8081 (N_8081,N_7977,N_7936);
and U8082 (N_8082,N_7867,N_7909);
and U8083 (N_8083,N_7846,N_7919);
nand U8084 (N_8084,N_7998,N_7863);
or U8085 (N_8085,N_7948,N_7917);
and U8086 (N_8086,N_7947,N_7908);
or U8087 (N_8087,N_7850,N_7947);
nor U8088 (N_8088,N_7914,N_7882);
and U8089 (N_8089,N_7847,N_7898);
xnor U8090 (N_8090,N_7853,N_7893);
or U8091 (N_8091,N_7947,N_7899);
xnor U8092 (N_8092,N_7941,N_7848);
nand U8093 (N_8093,N_7885,N_7891);
xor U8094 (N_8094,N_7908,N_7920);
nor U8095 (N_8095,N_7905,N_7901);
nor U8096 (N_8096,N_7872,N_7897);
xnor U8097 (N_8097,N_7956,N_7861);
xor U8098 (N_8098,N_7953,N_7869);
nor U8099 (N_8099,N_7956,N_7869);
or U8100 (N_8100,N_7995,N_7908);
and U8101 (N_8101,N_7880,N_7922);
nor U8102 (N_8102,N_7849,N_7994);
xnor U8103 (N_8103,N_7969,N_7938);
and U8104 (N_8104,N_7893,N_7915);
xnor U8105 (N_8105,N_7852,N_7875);
and U8106 (N_8106,N_7923,N_7898);
nand U8107 (N_8107,N_7841,N_7991);
xor U8108 (N_8108,N_7916,N_7871);
nand U8109 (N_8109,N_7907,N_7861);
or U8110 (N_8110,N_7873,N_7854);
nand U8111 (N_8111,N_7976,N_7975);
nand U8112 (N_8112,N_7845,N_7955);
xor U8113 (N_8113,N_7981,N_7973);
nor U8114 (N_8114,N_7846,N_7856);
nor U8115 (N_8115,N_7979,N_7922);
or U8116 (N_8116,N_7885,N_7949);
and U8117 (N_8117,N_7877,N_7889);
and U8118 (N_8118,N_7873,N_7993);
or U8119 (N_8119,N_7889,N_7896);
nor U8120 (N_8120,N_7877,N_7999);
nor U8121 (N_8121,N_7903,N_7948);
and U8122 (N_8122,N_7886,N_7872);
xor U8123 (N_8123,N_7987,N_7911);
xor U8124 (N_8124,N_7991,N_7936);
xor U8125 (N_8125,N_7969,N_7993);
xnor U8126 (N_8126,N_7907,N_7987);
and U8127 (N_8127,N_7931,N_7952);
or U8128 (N_8128,N_7970,N_7848);
xor U8129 (N_8129,N_7907,N_7968);
nor U8130 (N_8130,N_7941,N_7844);
nand U8131 (N_8131,N_7914,N_7873);
and U8132 (N_8132,N_7851,N_7955);
nand U8133 (N_8133,N_7933,N_7927);
nand U8134 (N_8134,N_7962,N_7885);
or U8135 (N_8135,N_7891,N_7889);
xnor U8136 (N_8136,N_7998,N_7958);
nor U8137 (N_8137,N_7944,N_7896);
xor U8138 (N_8138,N_7860,N_7842);
nand U8139 (N_8139,N_7907,N_7862);
nand U8140 (N_8140,N_7897,N_7876);
xor U8141 (N_8141,N_7877,N_7978);
xnor U8142 (N_8142,N_7855,N_7905);
or U8143 (N_8143,N_7974,N_7892);
and U8144 (N_8144,N_7986,N_7914);
or U8145 (N_8145,N_7856,N_7894);
xnor U8146 (N_8146,N_7969,N_7915);
nand U8147 (N_8147,N_7879,N_7993);
nor U8148 (N_8148,N_7950,N_7893);
nor U8149 (N_8149,N_7984,N_7907);
xnor U8150 (N_8150,N_7884,N_7931);
and U8151 (N_8151,N_7971,N_7912);
xnor U8152 (N_8152,N_7884,N_7844);
or U8153 (N_8153,N_7879,N_7884);
nor U8154 (N_8154,N_7922,N_7874);
or U8155 (N_8155,N_7911,N_7958);
nor U8156 (N_8156,N_7861,N_7997);
xnor U8157 (N_8157,N_7850,N_7846);
xnor U8158 (N_8158,N_7847,N_7950);
nand U8159 (N_8159,N_7940,N_7888);
and U8160 (N_8160,N_8125,N_8135);
or U8161 (N_8161,N_8049,N_8048);
xor U8162 (N_8162,N_8077,N_8067);
or U8163 (N_8163,N_8123,N_8073);
nand U8164 (N_8164,N_8013,N_8026);
nor U8165 (N_8165,N_8156,N_8037);
nor U8166 (N_8166,N_8101,N_8150);
and U8167 (N_8167,N_8021,N_8019);
and U8168 (N_8168,N_8116,N_8106);
or U8169 (N_8169,N_8153,N_8031);
nor U8170 (N_8170,N_8058,N_8043);
and U8171 (N_8171,N_8011,N_8079);
or U8172 (N_8172,N_8154,N_8007);
and U8173 (N_8173,N_8134,N_8059);
nor U8174 (N_8174,N_8017,N_8083);
nor U8175 (N_8175,N_8038,N_8143);
nand U8176 (N_8176,N_8062,N_8066);
nand U8177 (N_8177,N_8078,N_8088);
or U8178 (N_8178,N_8136,N_8130);
nand U8179 (N_8179,N_8052,N_8127);
xor U8180 (N_8180,N_8053,N_8029);
or U8181 (N_8181,N_8118,N_8045);
nand U8182 (N_8182,N_8041,N_8034);
or U8183 (N_8183,N_8039,N_8109);
and U8184 (N_8184,N_8144,N_8149);
or U8185 (N_8185,N_8155,N_8132);
and U8186 (N_8186,N_8159,N_8025);
or U8187 (N_8187,N_8003,N_8050);
and U8188 (N_8188,N_8090,N_8032);
nand U8189 (N_8189,N_8131,N_8044);
or U8190 (N_8190,N_8051,N_8068);
nand U8191 (N_8191,N_8028,N_8145);
and U8192 (N_8192,N_8057,N_8086);
xor U8193 (N_8193,N_8015,N_8110);
or U8194 (N_8194,N_8146,N_8107);
and U8195 (N_8195,N_8001,N_8103);
xnor U8196 (N_8196,N_8070,N_8085);
xor U8197 (N_8197,N_8033,N_8012);
or U8198 (N_8198,N_8138,N_8100);
nor U8199 (N_8199,N_8075,N_8124);
nand U8200 (N_8200,N_8102,N_8010);
or U8201 (N_8201,N_8018,N_8002);
or U8202 (N_8202,N_8105,N_8087);
xor U8203 (N_8203,N_8120,N_8047);
or U8204 (N_8204,N_8126,N_8148);
nor U8205 (N_8205,N_8099,N_8095);
nor U8206 (N_8206,N_8056,N_8080);
xnor U8207 (N_8207,N_8098,N_8055);
and U8208 (N_8208,N_8128,N_8076);
nor U8209 (N_8209,N_8005,N_8114);
or U8210 (N_8210,N_8112,N_8151);
or U8211 (N_8211,N_8141,N_8030);
nand U8212 (N_8212,N_8035,N_8094);
or U8213 (N_8213,N_8097,N_8006);
and U8214 (N_8214,N_8084,N_8129);
nand U8215 (N_8215,N_8024,N_8113);
and U8216 (N_8216,N_8081,N_8117);
and U8217 (N_8217,N_8092,N_8091);
xnor U8218 (N_8218,N_8065,N_8054);
and U8219 (N_8219,N_8152,N_8072);
nor U8220 (N_8220,N_8063,N_8096);
and U8221 (N_8221,N_8158,N_8023);
nor U8222 (N_8222,N_8036,N_8147);
nor U8223 (N_8223,N_8115,N_8000);
or U8224 (N_8224,N_8004,N_8060);
nor U8225 (N_8225,N_8142,N_8157);
and U8226 (N_8226,N_8040,N_8139);
nand U8227 (N_8227,N_8022,N_8111);
xnor U8228 (N_8228,N_8089,N_8046);
nor U8229 (N_8229,N_8119,N_8009);
nor U8230 (N_8230,N_8061,N_8020);
and U8231 (N_8231,N_8014,N_8016);
and U8232 (N_8232,N_8108,N_8008);
or U8233 (N_8233,N_8121,N_8133);
nor U8234 (N_8234,N_8122,N_8074);
xor U8235 (N_8235,N_8042,N_8140);
nand U8236 (N_8236,N_8069,N_8071);
and U8237 (N_8237,N_8137,N_8093);
nand U8238 (N_8238,N_8064,N_8104);
nand U8239 (N_8239,N_8082,N_8027);
or U8240 (N_8240,N_8028,N_8069);
or U8241 (N_8241,N_8053,N_8026);
xor U8242 (N_8242,N_8082,N_8150);
or U8243 (N_8243,N_8137,N_8130);
xor U8244 (N_8244,N_8087,N_8049);
xnor U8245 (N_8245,N_8035,N_8121);
nand U8246 (N_8246,N_8116,N_8118);
nand U8247 (N_8247,N_8151,N_8044);
or U8248 (N_8248,N_8058,N_8077);
and U8249 (N_8249,N_8093,N_8139);
nand U8250 (N_8250,N_8071,N_8060);
or U8251 (N_8251,N_8144,N_8114);
nand U8252 (N_8252,N_8083,N_8106);
and U8253 (N_8253,N_8057,N_8125);
and U8254 (N_8254,N_8024,N_8111);
nor U8255 (N_8255,N_8158,N_8065);
nor U8256 (N_8256,N_8027,N_8017);
nand U8257 (N_8257,N_8087,N_8064);
nand U8258 (N_8258,N_8106,N_8113);
nor U8259 (N_8259,N_8105,N_8019);
or U8260 (N_8260,N_8076,N_8005);
xnor U8261 (N_8261,N_8028,N_8049);
nor U8262 (N_8262,N_8100,N_8094);
xor U8263 (N_8263,N_8057,N_8004);
or U8264 (N_8264,N_8107,N_8029);
and U8265 (N_8265,N_8102,N_8156);
xnor U8266 (N_8266,N_8159,N_8081);
and U8267 (N_8267,N_8041,N_8049);
nor U8268 (N_8268,N_8157,N_8087);
and U8269 (N_8269,N_8062,N_8035);
or U8270 (N_8270,N_8070,N_8096);
nor U8271 (N_8271,N_8047,N_8145);
or U8272 (N_8272,N_8064,N_8021);
nor U8273 (N_8273,N_8094,N_8108);
and U8274 (N_8274,N_8037,N_8004);
or U8275 (N_8275,N_8001,N_8099);
nand U8276 (N_8276,N_8098,N_8137);
or U8277 (N_8277,N_8114,N_8038);
and U8278 (N_8278,N_8084,N_8114);
xor U8279 (N_8279,N_8112,N_8137);
xor U8280 (N_8280,N_8019,N_8070);
or U8281 (N_8281,N_8052,N_8087);
nand U8282 (N_8282,N_8127,N_8015);
nor U8283 (N_8283,N_8043,N_8075);
nor U8284 (N_8284,N_8020,N_8003);
or U8285 (N_8285,N_8145,N_8116);
nor U8286 (N_8286,N_8071,N_8153);
and U8287 (N_8287,N_8151,N_8087);
nand U8288 (N_8288,N_8139,N_8016);
xnor U8289 (N_8289,N_8153,N_8141);
and U8290 (N_8290,N_8123,N_8060);
or U8291 (N_8291,N_8119,N_8060);
and U8292 (N_8292,N_8048,N_8089);
or U8293 (N_8293,N_8042,N_8128);
xnor U8294 (N_8294,N_8067,N_8018);
xnor U8295 (N_8295,N_8124,N_8131);
xor U8296 (N_8296,N_8026,N_8106);
and U8297 (N_8297,N_8009,N_8152);
nor U8298 (N_8298,N_8066,N_8128);
xor U8299 (N_8299,N_8005,N_8042);
or U8300 (N_8300,N_8119,N_8158);
nor U8301 (N_8301,N_8107,N_8036);
and U8302 (N_8302,N_8150,N_8112);
and U8303 (N_8303,N_8042,N_8025);
nor U8304 (N_8304,N_8156,N_8023);
and U8305 (N_8305,N_8080,N_8129);
nand U8306 (N_8306,N_8005,N_8109);
nor U8307 (N_8307,N_8118,N_8035);
or U8308 (N_8308,N_8027,N_8153);
or U8309 (N_8309,N_8086,N_8091);
nor U8310 (N_8310,N_8079,N_8066);
and U8311 (N_8311,N_8139,N_8081);
xor U8312 (N_8312,N_8154,N_8013);
xor U8313 (N_8313,N_8074,N_8103);
nand U8314 (N_8314,N_8126,N_8129);
nand U8315 (N_8315,N_8081,N_8151);
or U8316 (N_8316,N_8038,N_8095);
and U8317 (N_8317,N_8061,N_8014);
or U8318 (N_8318,N_8025,N_8137);
and U8319 (N_8319,N_8057,N_8113);
and U8320 (N_8320,N_8246,N_8204);
xnor U8321 (N_8321,N_8219,N_8281);
nor U8322 (N_8322,N_8305,N_8270);
nand U8323 (N_8323,N_8272,N_8189);
nor U8324 (N_8324,N_8293,N_8205);
and U8325 (N_8325,N_8223,N_8256);
or U8326 (N_8326,N_8169,N_8233);
nor U8327 (N_8327,N_8266,N_8307);
nand U8328 (N_8328,N_8261,N_8163);
and U8329 (N_8329,N_8286,N_8250);
nand U8330 (N_8330,N_8226,N_8248);
nand U8331 (N_8331,N_8206,N_8214);
and U8332 (N_8332,N_8242,N_8202);
xor U8333 (N_8333,N_8318,N_8217);
nand U8334 (N_8334,N_8302,N_8284);
or U8335 (N_8335,N_8198,N_8173);
nand U8336 (N_8336,N_8277,N_8231);
xnor U8337 (N_8337,N_8176,N_8292);
nor U8338 (N_8338,N_8186,N_8174);
and U8339 (N_8339,N_8276,N_8168);
or U8340 (N_8340,N_8275,N_8194);
nand U8341 (N_8341,N_8232,N_8222);
nor U8342 (N_8342,N_8264,N_8179);
nand U8343 (N_8343,N_8237,N_8203);
nand U8344 (N_8344,N_8216,N_8192);
nor U8345 (N_8345,N_8290,N_8285);
nor U8346 (N_8346,N_8170,N_8213);
and U8347 (N_8347,N_8265,N_8197);
and U8348 (N_8348,N_8239,N_8236);
xnor U8349 (N_8349,N_8311,N_8271);
nand U8350 (N_8350,N_8225,N_8316);
or U8351 (N_8351,N_8258,N_8251);
or U8352 (N_8352,N_8308,N_8296);
nand U8353 (N_8353,N_8274,N_8228);
nor U8354 (N_8354,N_8294,N_8235);
nand U8355 (N_8355,N_8313,N_8287);
nor U8356 (N_8356,N_8208,N_8200);
and U8357 (N_8357,N_8280,N_8295);
and U8358 (N_8358,N_8196,N_8253);
or U8359 (N_8359,N_8312,N_8221);
and U8360 (N_8360,N_8243,N_8301);
nand U8361 (N_8361,N_8282,N_8193);
xor U8362 (N_8362,N_8184,N_8255);
and U8363 (N_8363,N_8297,N_8240);
nor U8364 (N_8364,N_8288,N_8199);
nand U8365 (N_8365,N_8314,N_8273);
or U8366 (N_8366,N_8269,N_8211);
and U8367 (N_8367,N_8291,N_8289);
xnor U8368 (N_8368,N_8283,N_8183);
nand U8369 (N_8369,N_8165,N_8300);
nor U8370 (N_8370,N_8188,N_8215);
or U8371 (N_8371,N_8209,N_8260);
and U8372 (N_8372,N_8247,N_8254);
and U8373 (N_8373,N_8279,N_8303);
nor U8374 (N_8374,N_8162,N_8160);
xnor U8375 (N_8375,N_8187,N_8185);
nand U8376 (N_8376,N_8201,N_8171);
nor U8377 (N_8377,N_8218,N_8212);
nand U8378 (N_8378,N_8210,N_8241);
nand U8379 (N_8379,N_8268,N_8166);
nand U8380 (N_8380,N_8262,N_8317);
xor U8381 (N_8381,N_8234,N_8229);
and U8382 (N_8382,N_8195,N_8164);
or U8383 (N_8383,N_8224,N_8315);
or U8384 (N_8384,N_8249,N_8263);
nor U8385 (N_8385,N_8180,N_8182);
or U8386 (N_8386,N_8161,N_8309);
and U8387 (N_8387,N_8175,N_8252);
xnor U8388 (N_8388,N_8244,N_8190);
xor U8389 (N_8389,N_8310,N_8177);
or U8390 (N_8390,N_8278,N_8259);
nand U8391 (N_8391,N_8304,N_8267);
xnor U8392 (N_8392,N_8207,N_8220);
or U8393 (N_8393,N_8319,N_8191);
nand U8394 (N_8394,N_8167,N_8172);
and U8395 (N_8395,N_8298,N_8238);
nand U8396 (N_8396,N_8230,N_8306);
and U8397 (N_8397,N_8181,N_8257);
nand U8398 (N_8398,N_8178,N_8299);
nor U8399 (N_8399,N_8245,N_8227);
or U8400 (N_8400,N_8224,N_8209);
nand U8401 (N_8401,N_8204,N_8230);
xor U8402 (N_8402,N_8250,N_8302);
xnor U8403 (N_8403,N_8235,N_8239);
nor U8404 (N_8404,N_8308,N_8278);
nor U8405 (N_8405,N_8170,N_8314);
or U8406 (N_8406,N_8204,N_8195);
nand U8407 (N_8407,N_8197,N_8187);
xnor U8408 (N_8408,N_8234,N_8202);
nor U8409 (N_8409,N_8181,N_8303);
nand U8410 (N_8410,N_8309,N_8187);
nor U8411 (N_8411,N_8189,N_8248);
and U8412 (N_8412,N_8173,N_8304);
nand U8413 (N_8413,N_8296,N_8234);
xor U8414 (N_8414,N_8235,N_8181);
and U8415 (N_8415,N_8214,N_8227);
nand U8416 (N_8416,N_8196,N_8269);
or U8417 (N_8417,N_8192,N_8178);
xnor U8418 (N_8418,N_8253,N_8227);
and U8419 (N_8419,N_8277,N_8305);
xnor U8420 (N_8420,N_8243,N_8250);
nand U8421 (N_8421,N_8183,N_8314);
and U8422 (N_8422,N_8222,N_8253);
or U8423 (N_8423,N_8221,N_8298);
xor U8424 (N_8424,N_8285,N_8200);
nor U8425 (N_8425,N_8303,N_8175);
xor U8426 (N_8426,N_8189,N_8198);
and U8427 (N_8427,N_8288,N_8236);
and U8428 (N_8428,N_8307,N_8196);
xnor U8429 (N_8429,N_8199,N_8296);
xor U8430 (N_8430,N_8285,N_8202);
and U8431 (N_8431,N_8261,N_8164);
nor U8432 (N_8432,N_8272,N_8180);
xnor U8433 (N_8433,N_8196,N_8280);
xnor U8434 (N_8434,N_8177,N_8203);
or U8435 (N_8435,N_8240,N_8258);
or U8436 (N_8436,N_8246,N_8193);
and U8437 (N_8437,N_8175,N_8214);
nand U8438 (N_8438,N_8251,N_8215);
xnor U8439 (N_8439,N_8304,N_8182);
and U8440 (N_8440,N_8254,N_8161);
and U8441 (N_8441,N_8254,N_8294);
and U8442 (N_8442,N_8258,N_8250);
or U8443 (N_8443,N_8310,N_8278);
nor U8444 (N_8444,N_8197,N_8279);
or U8445 (N_8445,N_8239,N_8302);
xor U8446 (N_8446,N_8274,N_8278);
nor U8447 (N_8447,N_8306,N_8259);
and U8448 (N_8448,N_8286,N_8189);
or U8449 (N_8449,N_8177,N_8304);
nand U8450 (N_8450,N_8181,N_8195);
xor U8451 (N_8451,N_8289,N_8198);
and U8452 (N_8452,N_8297,N_8226);
nor U8453 (N_8453,N_8253,N_8186);
xor U8454 (N_8454,N_8246,N_8314);
and U8455 (N_8455,N_8166,N_8265);
or U8456 (N_8456,N_8290,N_8245);
nor U8457 (N_8457,N_8318,N_8280);
or U8458 (N_8458,N_8192,N_8279);
and U8459 (N_8459,N_8193,N_8175);
and U8460 (N_8460,N_8197,N_8285);
and U8461 (N_8461,N_8206,N_8217);
nor U8462 (N_8462,N_8247,N_8310);
or U8463 (N_8463,N_8263,N_8197);
nand U8464 (N_8464,N_8277,N_8163);
or U8465 (N_8465,N_8253,N_8203);
nor U8466 (N_8466,N_8248,N_8181);
xor U8467 (N_8467,N_8165,N_8310);
and U8468 (N_8468,N_8222,N_8264);
nor U8469 (N_8469,N_8276,N_8185);
nand U8470 (N_8470,N_8201,N_8262);
and U8471 (N_8471,N_8317,N_8173);
and U8472 (N_8472,N_8218,N_8169);
xor U8473 (N_8473,N_8290,N_8259);
nor U8474 (N_8474,N_8308,N_8284);
or U8475 (N_8475,N_8208,N_8175);
or U8476 (N_8476,N_8287,N_8167);
nor U8477 (N_8477,N_8201,N_8242);
and U8478 (N_8478,N_8269,N_8276);
and U8479 (N_8479,N_8270,N_8263);
xor U8480 (N_8480,N_8374,N_8339);
nand U8481 (N_8481,N_8383,N_8461);
xnor U8482 (N_8482,N_8365,N_8345);
nor U8483 (N_8483,N_8358,N_8459);
xor U8484 (N_8484,N_8428,N_8440);
and U8485 (N_8485,N_8340,N_8395);
xnor U8486 (N_8486,N_8433,N_8409);
xor U8487 (N_8487,N_8332,N_8380);
nor U8488 (N_8488,N_8449,N_8391);
or U8489 (N_8489,N_8435,N_8337);
xor U8490 (N_8490,N_8458,N_8410);
nor U8491 (N_8491,N_8400,N_8397);
nand U8492 (N_8492,N_8331,N_8325);
nor U8493 (N_8493,N_8333,N_8450);
and U8494 (N_8494,N_8361,N_8457);
or U8495 (N_8495,N_8447,N_8357);
nand U8496 (N_8496,N_8454,N_8381);
and U8497 (N_8497,N_8322,N_8323);
and U8498 (N_8498,N_8403,N_8349);
or U8499 (N_8499,N_8479,N_8446);
or U8500 (N_8500,N_8402,N_8353);
nor U8501 (N_8501,N_8320,N_8444);
and U8502 (N_8502,N_8388,N_8335);
or U8503 (N_8503,N_8474,N_8470);
or U8504 (N_8504,N_8465,N_8441);
nand U8505 (N_8505,N_8443,N_8367);
xor U8506 (N_8506,N_8419,N_8379);
and U8507 (N_8507,N_8442,N_8412);
and U8508 (N_8508,N_8344,N_8414);
xor U8509 (N_8509,N_8467,N_8434);
nor U8510 (N_8510,N_8392,N_8420);
nor U8511 (N_8511,N_8376,N_8451);
xnor U8512 (N_8512,N_8324,N_8366);
nand U8513 (N_8513,N_8430,N_8452);
xor U8514 (N_8514,N_8437,N_8472);
and U8515 (N_8515,N_8343,N_8477);
nand U8516 (N_8516,N_8359,N_8423);
xnor U8517 (N_8517,N_8355,N_8405);
or U8518 (N_8518,N_8364,N_8464);
xor U8519 (N_8519,N_8363,N_8415);
xor U8520 (N_8520,N_8327,N_8329);
xnor U8521 (N_8521,N_8466,N_8427);
nor U8522 (N_8522,N_8429,N_8378);
nor U8523 (N_8523,N_8417,N_8384);
and U8524 (N_8524,N_8393,N_8445);
nand U8525 (N_8525,N_8387,N_8471);
and U8526 (N_8526,N_8389,N_8407);
nor U8527 (N_8527,N_8326,N_8413);
xor U8528 (N_8528,N_8369,N_8360);
nand U8529 (N_8529,N_8404,N_8373);
and U8530 (N_8530,N_8422,N_8385);
nor U8531 (N_8531,N_8408,N_8438);
nor U8532 (N_8532,N_8426,N_8390);
nor U8533 (N_8533,N_8362,N_8463);
nand U8534 (N_8534,N_8371,N_8411);
nand U8535 (N_8535,N_8336,N_8342);
and U8536 (N_8536,N_8436,N_8416);
and U8537 (N_8537,N_8468,N_8356);
or U8538 (N_8538,N_8341,N_8418);
nor U8539 (N_8539,N_8473,N_8432);
nand U8540 (N_8540,N_8421,N_8460);
xor U8541 (N_8541,N_8456,N_8394);
xnor U8542 (N_8542,N_8334,N_8330);
nor U8543 (N_8543,N_8352,N_8475);
nand U8544 (N_8544,N_8347,N_8396);
or U8545 (N_8545,N_8431,N_8453);
or U8546 (N_8546,N_8351,N_8401);
nand U8547 (N_8547,N_8476,N_8368);
or U8548 (N_8548,N_8439,N_8377);
xnor U8549 (N_8549,N_8399,N_8424);
and U8550 (N_8550,N_8425,N_8350);
and U8551 (N_8551,N_8469,N_8448);
nand U8552 (N_8552,N_8328,N_8338);
xor U8553 (N_8553,N_8398,N_8372);
xnor U8554 (N_8554,N_8382,N_8354);
and U8555 (N_8555,N_8462,N_8478);
and U8556 (N_8556,N_8375,N_8321);
or U8557 (N_8557,N_8348,N_8455);
and U8558 (N_8558,N_8406,N_8346);
and U8559 (N_8559,N_8386,N_8370);
xnor U8560 (N_8560,N_8434,N_8453);
nand U8561 (N_8561,N_8368,N_8365);
xnor U8562 (N_8562,N_8342,N_8355);
xor U8563 (N_8563,N_8347,N_8340);
nand U8564 (N_8564,N_8386,N_8444);
or U8565 (N_8565,N_8360,N_8461);
nor U8566 (N_8566,N_8461,N_8382);
or U8567 (N_8567,N_8454,N_8359);
or U8568 (N_8568,N_8382,N_8375);
nand U8569 (N_8569,N_8465,N_8414);
and U8570 (N_8570,N_8410,N_8456);
and U8571 (N_8571,N_8337,N_8340);
nor U8572 (N_8572,N_8361,N_8320);
xnor U8573 (N_8573,N_8474,N_8343);
and U8574 (N_8574,N_8388,N_8409);
nor U8575 (N_8575,N_8375,N_8423);
nand U8576 (N_8576,N_8386,N_8461);
or U8577 (N_8577,N_8387,N_8417);
nand U8578 (N_8578,N_8461,N_8436);
nand U8579 (N_8579,N_8445,N_8370);
nor U8580 (N_8580,N_8335,N_8346);
nor U8581 (N_8581,N_8411,N_8396);
or U8582 (N_8582,N_8407,N_8357);
xnor U8583 (N_8583,N_8435,N_8348);
xnor U8584 (N_8584,N_8447,N_8475);
or U8585 (N_8585,N_8413,N_8353);
nand U8586 (N_8586,N_8347,N_8432);
and U8587 (N_8587,N_8460,N_8366);
nand U8588 (N_8588,N_8458,N_8391);
xnor U8589 (N_8589,N_8345,N_8329);
or U8590 (N_8590,N_8373,N_8440);
and U8591 (N_8591,N_8425,N_8411);
or U8592 (N_8592,N_8408,N_8462);
nor U8593 (N_8593,N_8389,N_8469);
or U8594 (N_8594,N_8335,N_8466);
nand U8595 (N_8595,N_8448,N_8436);
or U8596 (N_8596,N_8403,N_8369);
nand U8597 (N_8597,N_8406,N_8387);
xor U8598 (N_8598,N_8426,N_8326);
nor U8599 (N_8599,N_8429,N_8433);
and U8600 (N_8600,N_8392,N_8447);
nor U8601 (N_8601,N_8343,N_8341);
nor U8602 (N_8602,N_8381,N_8377);
xor U8603 (N_8603,N_8463,N_8326);
and U8604 (N_8604,N_8418,N_8468);
xnor U8605 (N_8605,N_8466,N_8348);
nand U8606 (N_8606,N_8364,N_8383);
nand U8607 (N_8607,N_8459,N_8338);
nor U8608 (N_8608,N_8380,N_8320);
nor U8609 (N_8609,N_8446,N_8436);
nor U8610 (N_8610,N_8419,N_8444);
or U8611 (N_8611,N_8337,N_8342);
nor U8612 (N_8612,N_8422,N_8378);
nor U8613 (N_8613,N_8374,N_8447);
nand U8614 (N_8614,N_8320,N_8373);
or U8615 (N_8615,N_8414,N_8376);
or U8616 (N_8616,N_8351,N_8468);
or U8617 (N_8617,N_8458,N_8372);
or U8618 (N_8618,N_8438,N_8364);
nand U8619 (N_8619,N_8321,N_8374);
or U8620 (N_8620,N_8418,N_8350);
nand U8621 (N_8621,N_8479,N_8348);
nand U8622 (N_8622,N_8370,N_8422);
xor U8623 (N_8623,N_8398,N_8365);
nand U8624 (N_8624,N_8425,N_8396);
or U8625 (N_8625,N_8368,N_8377);
nand U8626 (N_8626,N_8336,N_8343);
nand U8627 (N_8627,N_8444,N_8414);
and U8628 (N_8628,N_8419,N_8475);
nor U8629 (N_8629,N_8389,N_8346);
nand U8630 (N_8630,N_8371,N_8468);
or U8631 (N_8631,N_8335,N_8367);
nand U8632 (N_8632,N_8398,N_8385);
nor U8633 (N_8633,N_8430,N_8385);
nor U8634 (N_8634,N_8444,N_8375);
and U8635 (N_8635,N_8321,N_8441);
xor U8636 (N_8636,N_8348,N_8426);
or U8637 (N_8637,N_8434,N_8427);
or U8638 (N_8638,N_8357,N_8321);
xnor U8639 (N_8639,N_8365,N_8367);
nor U8640 (N_8640,N_8638,N_8599);
and U8641 (N_8641,N_8534,N_8614);
nand U8642 (N_8642,N_8486,N_8619);
or U8643 (N_8643,N_8547,N_8630);
nor U8644 (N_8644,N_8603,N_8637);
or U8645 (N_8645,N_8594,N_8512);
nand U8646 (N_8646,N_8507,N_8564);
nand U8647 (N_8647,N_8542,N_8553);
or U8648 (N_8648,N_8502,N_8550);
and U8649 (N_8649,N_8569,N_8549);
and U8650 (N_8650,N_8587,N_8496);
nand U8651 (N_8651,N_8598,N_8610);
and U8652 (N_8652,N_8627,N_8636);
nor U8653 (N_8653,N_8501,N_8525);
nand U8654 (N_8654,N_8523,N_8521);
or U8655 (N_8655,N_8607,N_8580);
nand U8656 (N_8656,N_8499,N_8584);
xnor U8657 (N_8657,N_8586,N_8524);
nor U8658 (N_8658,N_8515,N_8608);
xnor U8659 (N_8659,N_8620,N_8557);
nor U8660 (N_8660,N_8517,N_8555);
or U8661 (N_8661,N_8546,N_8572);
or U8662 (N_8662,N_8565,N_8621);
and U8663 (N_8663,N_8560,N_8493);
nor U8664 (N_8664,N_8633,N_8506);
and U8665 (N_8665,N_8576,N_8578);
xnor U8666 (N_8666,N_8497,N_8552);
and U8667 (N_8667,N_8518,N_8537);
nor U8668 (N_8668,N_8551,N_8519);
xnor U8669 (N_8669,N_8577,N_8622);
xnor U8670 (N_8670,N_8590,N_8606);
xnor U8671 (N_8671,N_8612,N_8604);
and U8672 (N_8672,N_8568,N_8487);
nor U8673 (N_8673,N_8535,N_8631);
xnor U8674 (N_8674,N_8532,N_8494);
nor U8675 (N_8675,N_8573,N_8632);
xor U8676 (N_8676,N_8617,N_8513);
and U8677 (N_8677,N_8579,N_8566);
nor U8678 (N_8678,N_8581,N_8480);
xor U8679 (N_8679,N_8591,N_8639);
xor U8680 (N_8680,N_8556,N_8482);
or U8681 (N_8681,N_8489,N_8628);
nand U8682 (N_8682,N_8514,N_8585);
nor U8683 (N_8683,N_8583,N_8540);
nor U8684 (N_8684,N_8624,N_8634);
nor U8685 (N_8685,N_8558,N_8618);
nand U8686 (N_8686,N_8545,N_8561);
xnor U8687 (N_8687,N_8522,N_8548);
xor U8688 (N_8688,N_8543,N_8492);
or U8689 (N_8689,N_8483,N_8623);
nor U8690 (N_8690,N_8505,N_8570);
nor U8691 (N_8691,N_8611,N_8615);
or U8692 (N_8692,N_8495,N_8625);
nand U8693 (N_8693,N_8626,N_8485);
or U8694 (N_8694,N_8530,N_8488);
or U8695 (N_8695,N_8616,N_8559);
and U8696 (N_8696,N_8593,N_8567);
nand U8697 (N_8697,N_8504,N_8605);
xnor U8698 (N_8698,N_8528,N_8529);
or U8699 (N_8699,N_8589,N_8554);
xnor U8700 (N_8700,N_8511,N_8531);
or U8701 (N_8701,N_8490,N_8484);
nor U8702 (N_8702,N_8613,N_8596);
and U8703 (N_8703,N_8562,N_8527);
nand U8704 (N_8704,N_8602,N_8539);
or U8705 (N_8705,N_8541,N_8571);
nand U8706 (N_8706,N_8516,N_8481);
nor U8707 (N_8707,N_8491,N_8597);
or U8708 (N_8708,N_8582,N_8609);
nor U8709 (N_8709,N_8498,N_8509);
or U8710 (N_8710,N_8520,N_8563);
nand U8711 (N_8711,N_8503,N_8600);
nor U8712 (N_8712,N_8526,N_8508);
nand U8713 (N_8713,N_8536,N_8510);
nor U8714 (N_8714,N_8601,N_8595);
nor U8715 (N_8715,N_8629,N_8500);
or U8716 (N_8716,N_8533,N_8538);
and U8717 (N_8717,N_8635,N_8588);
nand U8718 (N_8718,N_8575,N_8574);
and U8719 (N_8719,N_8544,N_8592);
xor U8720 (N_8720,N_8544,N_8527);
nor U8721 (N_8721,N_8622,N_8500);
xor U8722 (N_8722,N_8634,N_8499);
nand U8723 (N_8723,N_8516,N_8496);
or U8724 (N_8724,N_8604,N_8499);
nor U8725 (N_8725,N_8558,N_8624);
or U8726 (N_8726,N_8618,N_8546);
nor U8727 (N_8727,N_8583,N_8608);
nor U8728 (N_8728,N_8573,N_8591);
nor U8729 (N_8729,N_8486,N_8501);
nand U8730 (N_8730,N_8582,N_8590);
xnor U8731 (N_8731,N_8526,N_8494);
nand U8732 (N_8732,N_8584,N_8501);
nor U8733 (N_8733,N_8601,N_8483);
nor U8734 (N_8734,N_8625,N_8634);
and U8735 (N_8735,N_8499,N_8519);
nor U8736 (N_8736,N_8484,N_8612);
and U8737 (N_8737,N_8556,N_8542);
nand U8738 (N_8738,N_8622,N_8492);
or U8739 (N_8739,N_8614,N_8557);
xor U8740 (N_8740,N_8571,N_8597);
nor U8741 (N_8741,N_8552,N_8519);
and U8742 (N_8742,N_8513,N_8481);
nor U8743 (N_8743,N_8587,N_8607);
and U8744 (N_8744,N_8610,N_8631);
nor U8745 (N_8745,N_8578,N_8487);
or U8746 (N_8746,N_8638,N_8585);
and U8747 (N_8747,N_8569,N_8513);
nor U8748 (N_8748,N_8555,N_8582);
nand U8749 (N_8749,N_8561,N_8557);
and U8750 (N_8750,N_8556,N_8624);
xnor U8751 (N_8751,N_8588,N_8578);
xnor U8752 (N_8752,N_8510,N_8591);
or U8753 (N_8753,N_8490,N_8499);
or U8754 (N_8754,N_8484,N_8547);
xnor U8755 (N_8755,N_8600,N_8590);
and U8756 (N_8756,N_8490,N_8619);
or U8757 (N_8757,N_8528,N_8535);
or U8758 (N_8758,N_8485,N_8548);
and U8759 (N_8759,N_8547,N_8530);
or U8760 (N_8760,N_8579,N_8577);
and U8761 (N_8761,N_8602,N_8622);
and U8762 (N_8762,N_8609,N_8602);
and U8763 (N_8763,N_8560,N_8620);
nor U8764 (N_8764,N_8577,N_8482);
and U8765 (N_8765,N_8588,N_8586);
or U8766 (N_8766,N_8596,N_8512);
nor U8767 (N_8767,N_8565,N_8531);
and U8768 (N_8768,N_8616,N_8558);
xnor U8769 (N_8769,N_8560,N_8535);
nor U8770 (N_8770,N_8493,N_8494);
or U8771 (N_8771,N_8540,N_8558);
nor U8772 (N_8772,N_8569,N_8494);
and U8773 (N_8773,N_8490,N_8520);
nor U8774 (N_8774,N_8560,N_8570);
xor U8775 (N_8775,N_8540,N_8632);
xor U8776 (N_8776,N_8557,N_8500);
or U8777 (N_8777,N_8621,N_8584);
nand U8778 (N_8778,N_8577,N_8520);
xor U8779 (N_8779,N_8527,N_8535);
and U8780 (N_8780,N_8625,N_8537);
nand U8781 (N_8781,N_8592,N_8586);
xnor U8782 (N_8782,N_8557,N_8533);
and U8783 (N_8783,N_8523,N_8502);
and U8784 (N_8784,N_8498,N_8502);
or U8785 (N_8785,N_8627,N_8520);
nand U8786 (N_8786,N_8611,N_8626);
nand U8787 (N_8787,N_8611,N_8624);
or U8788 (N_8788,N_8584,N_8481);
and U8789 (N_8789,N_8613,N_8546);
or U8790 (N_8790,N_8568,N_8505);
nand U8791 (N_8791,N_8600,N_8582);
xnor U8792 (N_8792,N_8583,N_8577);
or U8793 (N_8793,N_8566,N_8572);
or U8794 (N_8794,N_8503,N_8483);
nand U8795 (N_8795,N_8608,N_8621);
or U8796 (N_8796,N_8553,N_8552);
nor U8797 (N_8797,N_8547,N_8629);
nor U8798 (N_8798,N_8569,N_8525);
or U8799 (N_8799,N_8522,N_8483);
and U8800 (N_8800,N_8705,N_8645);
or U8801 (N_8801,N_8743,N_8649);
nor U8802 (N_8802,N_8784,N_8775);
or U8803 (N_8803,N_8647,N_8756);
xor U8804 (N_8804,N_8770,N_8776);
xnor U8805 (N_8805,N_8713,N_8772);
nand U8806 (N_8806,N_8642,N_8664);
nor U8807 (N_8807,N_8672,N_8692);
nor U8808 (N_8808,N_8768,N_8774);
and U8809 (N_8809,N_8791,N_8673);
nand U8810 (N_8810,N_8687,N_8667);
xnor U8811 (N_8811,N_8684,N_8754);
xor U8812 (N_8812,N_8735,N_8727);
or U8813 (N_8813,N_8792,N_8704);
or U8814 (N_8814,N_8709,N_8668);
nor U8815 (N_8815,N_8734,N_8749);
nand U8816 (N_8816,N_8737,N_8780);
or U8817 (N_8817,N_8679,N_8662);
xnor U8818 (N_8818,N_8777,N_8757);
xnor U8819 (N_8819,N_8680,N_8766);
or U8820 (N_8820,N_8771,N_8708);
or U8821 (N_8821,N_8648,N_8702);
xor U8822 (N_8822,N_8755,N_8646);
xor U8823 (N_8823,N_8730,N_8694);
nand U8824 (N_8824,N_8751,N_8736);
or U8825 (N_8825,N_8663,N_8782);
nor U8826 (N_8826,N_8701,N_8711);
or U8827 (N_8827,N_8699,N_8718);
nor U8828 (N_8828,N_8674,N_8677);
nor U8829 (N_8829,N_8748,N_8695);
xor U8830 (N_8830,N_8716,N_8712);
or U8831 (N_8831,N_8657,N_8767);
or U8832 (N_8832,N_8783,N_8731);
xnor U8833 (N_8833,N_8707,N_8761);
nor U8834 (N_8834,N_8658,N_8720);
or U8835 (N_8835,N_8799,N_8759);
or U8836 (N_8836,N_8740,N_8671);
nand U8837 (N_8837,N_8725,N_8659);
xnor U8838 (N_8838,N_8765,N_8741);
xor U8839 (N_8839,N_8643,N_8793);
xnor U8840 (N_8840,N_8682,N_8798);
nand U8841 (N_8841,N_8758,N_8656);
nor U8842 (N_8842,N_8760,N_8655);
or U8843 (N_8843,N_8779,N_8742);
and U8844 (N_8844,N_8654,N_8732);
and U8845 (N_8845,N_8660,N_8796);
or U8846 (N_8846,N_8785,N_8681);
xnor U8847 (N_8847,N_8688,N_8726);
or U8848 (N_8848,N_8721,N_8652);
or U8849 (N_8849,N_8722,N_8670);
or U8850 (N_8850,N_8669,N_8703);
nand U8851 (N_8851,N_8745,N_8752);
nand U8852 (N_8852,N_8661,N_8724);
nor U8853 (N_8853,N_8706,N_8697);
nand U8854 (N_8854,N_8653,N_8744);
or U8855 (N_8855,N_8733,N_8650);
or U8856 (N_8856,N_8676,N_8781);
xnor U8857 (N_8857,N_8773,N_8651);
and U8858 (N_8858,N_8675,N_8683);
nand U8859 (N_8859,N_8786,N_8723);
and U8860 (N_8860,N_8690,N_8763);
xnor U8861 (N_8861,N_8729,N_8795);
or U8862 (N_8862,N_8714,N_8700);
nor U8863 (N_8863,N_8693,N_8762);
xor U8864 (N_8864,N_8640,N_8689);
or U8865 (N_8865,N_8794,N_8753);
and U8866 (N_8866,N_8715,N_8686);
and U8867 (N_8867,N_8710,N_8696);
and U8868 (N_8868,N_8797,N_8789);
nand U8869 (N_8869,N_8750,N_8769);
nand U8870 (N_8870,N_8764,N_8685);
nor U8871 (N_8871,N_8787,N_8698);
nand U8872 (N_8872,N_8739,N_8719);
and U8873 (N_8873,N_8790,N_8717);
nor U8874 (N_8874,N_8747,N_8788);
nor U8875 (N_8875,N_8738,N_8728);
or U8876 (N_8876,N_8644,N_8665);
nor U8877 (N_8877,N_8678,N_8666);
nor U8878 (N_8878,N_8691,N_8746);
xnor U8879 (N_8879,N_8778,N_8641);
xnor U8880 (N_8880,N_8788,N_8728);
nor U8881 (N_8881,N_8793,N_8694);
nand U8882 (N_8882,N_8778,N_8773);
or U8883 (N_8883,N_8701,N_8657);
xnor U8884 (N_8884,N_8661,N_8792);
nand U8885 (N_8885,N_8762,N_8768);
nor U8886 (N_8886,N_8720,N_8646);
xor U8887 (N_8887,N_8673,N_8741);
or U8888 (N_8888,N_8724,N_8643);
and U8889 (N_8889,N_8789,N_8671);
nor U8890 (N_8890,N_8724,N_8726);
and U8891 (N_8891,N_8689,N_8688);
nand U8892 (N_8892,N_8727,N_8717);
xor U8893 (N_8893,N_8723,N_8679);
nor U8894 (N_8894,N_8752,N_8793);
or U8895 (N_8895,N_8774,N_8733);
xor U8896 (N_8896,N_8743,N_8762);
xor U8897 (N_8897,N_8744,N_8725);
or U8898 (N_8898,N_8707,N_8708);
xor U8899 (N_8899,N_8744,N_8726);
xor U8900 (N_8900,N_8775,N_8785);
xnor U8901 (N_8901,N_8701,N_8731);
xor U8902 (N_8902,N_8745,N_8715);
and U8903 (N_8903,N_8642,N_8647);
or U8904 (N_8904,N_8797,N_8695);
and U8905 (N_8905,N_8690,N_8770);
xnor U8906 (N_8906,N_8680,N_8742);
xor U8907 (N_8907,N_8685,N_8768);
nor U8908 (N_8908,N_8749,N_8747);
nor U8909 (N_8909,N_8734,N_8735);
or U8910 (N_8910,N_8671,N_8776);
nor U8911 (N_8911,N_8740,N_8715);
nor U8912 (N_8912,N_8752,N_8700);
and U8913 (N_8913,N_8669,N_8645);
and U8914 (N_8914,N_8779,N_8755);
nand U8915 (N_8915,N_8746,N_8732);
nand U8916 (N_8916,N_8794,N_8646);
nor U8917 (N_8917,N_8752,N_8659);
nor U8918 (N_8918,N_8678,N_8694);
xor U8919 (N_8919,N_8753,N_8723);
nor U8920 (N_8920,N_8720,N_8782);
or U8921 (N_8921,N_8781,N_8743);
or U8922 (N_8922,N_8750,N_8749);
or U8923 (N_8923,N_8744,N_8712);
nor U8924 (N_8924,N_8779,N_8724);
xor U8925 (N_8925,N_8656,N_8788);
or U8926 (N_8926,N_8662,N_8785);
or U8927 (N_8927,N_8773,N_8749);
nor U8928 (N_8928,N_8795,N_8745);
and U8929 (N_8929,N_8641,N_8751);
nand U8930 (N_8930,N_8759,N_8763);
and U8931 (N_8931,N_8785,N_8764);
nor U8932 (N_8932,N_8746,N_8774);
and U8933 (N_8933,N_8751,N_8658);
and U8934 (N_8934,N_8758,N_8707);
xnor U8935 (N_8935,N_8655,N_8652);
nand U8936 (N_8936,N_8734,N_8705);
nand U8937 (N_8937,N_8656,N_8678);
nand U8938 (N_8938,N_8776,N_8682);
xor U8939 (N_8939,N_8649,N_8790);
and U8940 (N_8940,N_8727,N_8781);
nand U8941 (N_8941,N_8682,N_8754);
nand U8942 (N_8942,N_8749,N_8706);
xnor U8943 (N_8943,N_8691,N_8792);
xnor U8944 (N_8944,N_8670,N_8681);
nor U8945 (N_8945,N_8755,N_8661);
and U8946 (N_8946,N_8723,N_8781);
xor U8947 (N_8947,N_8731,N_8730);
or U8948 (N_8948,N_8645,N_8764);
xor U8949 (N_8949,N_8715,N_8774);
nor U8950 (N_8950,N_8729,N_8657);
xnor U8951 (N_8951,N_8739,N_8771);
or U8952 (N_8952,N_8658,N_8679);
xnor U8953 (N_8953,N_8787,N_8757);
nor U8954 (N_8954,N_8778,N_8681);
or U8955 (N_8955,N_8742,N_8777);
xor U8956 (N_8956,N_8651,N_8688);
or U8957 (N_8957,N_8759,N_8760);
xor U8958 (N_8958,N_8704,N_8757);
or U8959 (N_8959,N_8788,N_8688);
xnor U8960 (N_8960,N_8812,N_8824);
and U8961 (N_8961,N_8911,N_8802);
nand U8962 (N_8962,N_8846,N_8872);
or U8963 (N_8963,N_8834,N_8871);
or U8964 (N_8964,N_8899,N_8934);
nand U8965 (N_8965,N_8931,N_8827);
or U8966 (N_8966,N_8891,N_8893);
xor U8967 (N_8967,N_8821,N_8877);
nand U8968 (N_8968,N_8907,N_8807);
and U8969 (N_8969,N_8845,N_8947);
and U8970 (N_8970,N_8867,N_8865);
and U8971 (N_8971,N_8830,N_8811);
nand U8972 (N_8972,N_8926,N_8878);
or U8973 (N_8973,N_8916,N_8952);
nor U8974 (N_8974,N_8806,N_8896);
nand U8975 (N_8975,N_8900,N_8924);
xnor U8976 (N_8976,N_8957,N_8912);
nor U8977 (N_8977,N_8919,N_8855);
and U8978 (N_8978,N_8935,N_8895);
and U8979 (N_8979,N_8928,N_8941);
or U8980 (N_8980,N_8879,N_8813);
and U8981 (N_8981,N_8858,N_8853);
nor U8982 (N_8982,N_8923,N_8943);
nand U8983 (N_8983,N_8839,N_8909);
xnor U8984 (N_8984,N_8906,N_8917);
xnor U8985 (N_8985,N_8831,N_8862);
nand U8986 (N_8986,N_8885,N_8949);
xnor U8987 (N_8987,N_8889,N_8860);
nor U8988 (N_8988,N_8874,N_8828);
nand U8989 (N_8989,N_8873,N_8817);
and U8990 (N_8990,N_8914,N_8945);
and U8991 (N_8991,N_8848,N_8892);
and U8992 (N_8992,N_8925,N_8803);
xnor U8993 (N_8993,N_8849,N_8832);
nand U8994 (N_8994,N_8886,N_8842);
or U8995 (N_8995,N_8959,N_8863);
xor U8996 (N_8996,N_8836,N_8838);
nand U8997 (N_8997,N_8823,N_8864);
or U8998 (N_8998,N_8884,N_8944);
xnor U8999 (N_8999,N_8936,N_8956);
and U9000 (N_9000,N_8822,N_8958);
nand U9001 (N_9001,N_8852,N_8829);
nand U9002 (N_9002,N_8804,N_8866);
xnor U9003 (N_9003,N_8887,N_8929);
and U9004 (N_9004,N_8938,N_8951);
nor U9005 (N_9005,N_8946,N_8883);
nand U9006 (N_9006,N_8841,N_8908);
xor U9007 (N_9007,N_8869,N_8901);
and U9008 (N_9008,N_8856,N_8939);
xor U9009 (N_9009,N_8857,N_8875);
xnor U9010 (N_9010,N_8880,N_8882);
xor U9011 (N_9011,N_8921,N_8955);
nand U9012 (N_9012,N_8937,N_8953);
nand U9013 (N_9013,N_8844,N_8833);
xor U9014 (N_9014,N_8905,N_8902);
and U9015 (N_9015,N_8810,N_8835);
nor U9016 (N_9016,N_8801,N_8826);
or U9017 (N_9017,N_8876,N_8805);
nand U9018 (N_9018,N_8897,N_8920);
or U9019 (N_9019,N_8819,N_8913);
xor U9020 (N_9020,N_8870,N_8854);
or U9021 (N_9021,N_8825,N_8904);
nor U9022 (N_9022,N_8888,N_8840);
nor U9023 (N_9023,N_8814,N_8898);
nand U9024 (N_9024,N_8915,N_8903);
nor U9025 (N_9025,N_8932,N_8850);
or U9026 (N_9026,N_8818,N_8950);
or U9027 (N_9027,N_8922,N_8954);
and U9028 (N_9028,N_8942,N_8868);
or U9029 (N_9029,N_8933,N_8910);
nor U9030 (N_9030,N_8809,N_8927);
nand U9031 (N_9031,N_8837,N_8816);
nand U9032 (N_9032,N_8918,N_8894);
nor U9033 (N_9033,N_8940,N_8859);
and U9034 (N_9034,N_8815,N_8861);
and U9035 (N_9035,N_8800,N_8890);
nand U9036 (N_9036,N_8948,N_8820);
nor U9037 (N_9037,N_8843,N_8847);
nand U9038 (N_9038,N_8881,N_8808);
xor U9039 (N_9039,N_8851,N_8930);
xor U9040 (N_9040,N_8901,N_8954);
or U9041 (N_9041,N_8850,N_8894);
or U9042 (N_9042,N_8842,N_8844);
and U9043 (N_9043,N_8934,N_8883);
and U9044 (N_9044,N_8867,N_8880);
nor U9045 (N_9045,N_8909,N_8848);
nor U9046 (N_9046,N_8834,N_8807);
and U9047 (N_9047,N_8813,N_8814);
nand U9048 (N_9048,N_8810,N_8893);
xnor U9049 (N_9049,N_8831,N_8898);
xor U9050 (N_9050,N_8835,N_8958);
nand U9051 (N_9051,N_8883,N_8938);
nor U9052 (N_9052,N_8830,N_8920);
and U9053 (N_9053,N_8813,N_8831);
xnor U9054 (N_9054,N_8812,N_8924);
and U9055 (N_9055,N_8922,N_8849);
nand U9056 (N_9056,N_8852,N_8901);
or U9057 (N_9057,N_8946,N_8800);
nor U9058 (N_9058,N_8855,N_8931);
or U9059 (N_9059,N_8890,N_8954);
nor U9060 (N_9060,N_8910,N_8841);
nand U9061 (N_9061,N_8809,N_8951);
and U9062 (N_9062,N_8958,N_8887);
nor U9063 (N_9063,N_8914,N_8826);
nor U9064 (N_9064,N_8802,N_8934);
and U9065 (N_9065,N_8868,N_8959);
xnor U9066 (N_9066,N_8879,N_8837);
and U9067 (N_9067,N_8880,N_8901);
or U9068 (N_9068,N_8922,N_8875);
and U9069 (N_9069,N_8922,N_8912);
or U9070 (N_9070,N_8847,N_8855);
and U9071 (N_9071,N_8843,N_8868);
xor U9072 (N_9072,N_8834,N_8853);
or U9073 (N_9073,N_8851,N_8891);
or U9074 (N_9074,N_8951,N_8866);
nand U9075 (N_9075,N_8930,N_8862);
or U9076 (N_9076,N_8897,N_8809);
xnor U9077 (N_9077,N_8923,N_8881);
nor U9078 (N_9078,N_8958,N_8878);
or U9079 (N_9079,N_8915,N_8909);
and U9080 (N_9080,N_8908,N_8927);
nand U9081 (N_9081,N_8825,N_8832);
or U9082 (N_9082,N_8950,N_8842);
and U9083 (N_9083,N_8885,N_8889);
nor U9084 (N_9084,N_8889,N_8876);
and U9085 (N_9085,N_8863,N_8853);
xor U9086 (N_9086,N_8911,N_8868);
nand U9087 (N_9087,N_8812,N_8816);
nand U9088 (N_9088,N_8958,N_8915);
nor U9089 (N_9089,N_8903,N_8815);
nand U9090 (N_9090,N_8884,N_8842);
and U9091 (N_9091,N_8911,N_8803);
or U9092 (N_9092,N_8858,N_8881);
or U9093 (N_9093,N_8850,N_8813);
or U9094 (N_9094,N_8834,N_8936);
nor U9095 (N_9095,N_8814,N_8948);
and U9096 (N_9096,N_8924,N_8939);
xnor U9097 (N_9097,N_8800,N_8843);
nand U9098 (N_9098,N_8827,N_8843);
and U9099 (N_9099,N_8864,N_8837);
or U9100 (N_9100,N_8816,N_8852);
xnor U9101 (N_9101,N_8833,N_8898);
or U9102 (N_9102,N_8901,N_8884);
nand U9103 (N_9103,N_8956,N_8927);
xnor U9104 (N_9104,N_8953,N_8933);
xnor U9105 (N_9105,N_8957,N_8809);
and U9106 (N_9106,N_8893,N_8801);
nor U9107 (N_9107,N_8862,N_8909);
nand U9108 (N_9108,N_8914,N_8855);
and U9109 (N_9109,N_8859,N_8895);
and U9110 (N_9110,N_8883,N_8933);
and U9111 (N_9111,N_8891,N_8896);
xnor U9112 (N_9112,N_8928,N_8913);
or U9113 (N_9113,N_8955,N_8891);
and U9114 (N_9114,N_8849,N_8809);
xnor U9115 (N_9115,N_8957,N_8953);
and U9116 (N_9116,N_8959,N_8923);
nand U9117 (N_9117,N_8838,N_8809);
nor U9118 (N_9118,N_8927,N_8814);
and U9119 (N_9119,N_8885,N_8942);
nand U9120 (N_9120,N_9093,N_9033);
or U9121 (N_9121,N_8976,N_9096);
nand U9122 (N_9122,N_9031,N_9043);
xnor U9123 (N_9123,N_9014,N_9022);
nand U9124 (N_9124,N_8975,N_8964);
nor U9125 (N_9125,N_8984,N_9061);
nand U9126 (N_9126,N_9013,N_9002);
xnor U9127 (N_9127,N_9011,N_9001);
nand U9128 (N_9128,N_9098,N_9101);
xnor U9129 (N_9129,N_9051,N_9016);
nor U9130 (N_9130,N_9113,N_9027);
nor U9131 (N_9131,N_9107,N_9094);
xor U9132 (N_9132,N_8987,N_9081);
and U9133 (N_9133,N_9116,N_9077);
and U9134 (N_9134,N_9105,N_9088);
xor U9135 (N_9135,N_9082,N_8982);
xor U9136 (N_9136,N_9036,N_9039);
xor U9137 (N_9137,N_9069,N_8973);
nor U9138 (N_9138,N_8990,N_9059);
nand U9139 (N_9139,N_9026,N_9042);
or U9140 (N_9140,N_8970,N_9119);
or U9141 (N_9141,N_9103,N_9117);
and U9142 (N_9142,N_9006,N_9057);
and U9143 (N_9143,N_9053,N_9060);
nor U9144 (N_9144,N_9032,N_8962);
xor U9145 (N_9145,N_9034,N_8977);
nor U9146 (N_9146,N_8988,N_9092);
nand U9147 (N_9147,N_9019,N_8965);
nor U9148 (N_9148,N_9063,N_9025);
or U9149 (N_9149,N_9003,N_8966);
and U9150 (N_9150,N_9058,N_8969);
xor U9151 (N_9151,N_9055,N_9065);
or U9152 (N_9152,N_9049,N_9047);
nor U9153 (N_9153,N_8993,N_9078);
and U9154 (N_9154,N_9111,N_9109);
nor U9155 (N_9155,N_9010,N_9075);
or U9156 (N_9156,N_9009,N_9108);
nand U9157 (N_9157,N_9045,N_9021);
nor U9158 (N_9158,N_9052,N_8972);
xnor U9159 (N_9159,N_9112,N_9074);
or U9160 (N_9160,N_9087,N_9104);
or U9161 (N_9161,N_9040,N_9017);
or U9162 (N_9162,N_9007,N_9090);
nor U9163 (N_9163,N_9035,N_9038);
xor U9164 (N_9164,N_9068,N_9037);
nand U9165 (N_9165,N_9028,N_9023);
xor U9166 (N_9166,N_8991,N_9102);
xor U9167 (N_9167,N_9067,N_8995);
nand U9168 (N_9168,N_9041,N_8978);
or U9169 (N_9169,N_8971,N_9083);
nor U9170 (N_9170,N_9054,N_9004);
or U9171 (N_9171,N_8981,N_9079);
or U9172 (N_9172,N_9085,N_9114);
and U9173 (N_9173,N_8986,N_9072);
nand U9174 (N_9174,N_9070,N_9066);
nor U9175 (N_9175,N_9008,N_8996);
nand U9176 (N_9176,N_8968,N_8998);
and U9177 (N_9177,N_9050,N_9076);
xnor U9178 (N_9178,N_9030,N_8967);
xnor U9179 (N_9179,N_9029,N_9000);
nand U9180 (N_9180,N_8997,N_9118);
nor U9181 (N_9181,N_8999,N_8963);
nor U9182 (N_9182,N_9091,N_9084);
xnor U9183 (N_9183,N_8989,N_9062);
and U9184 (N_9184,N_8979,N_9099);
nor U9185 (N_9185,N_9095,N_9115);
xor U9186 (N_9186,N_8974,N_9089);
nand U9187 (N_9187,N_9048,N_9110);
and U9188 (N_9188,N_9044,N_9080);
nand U9189 (N_9189,N_9015,N_9012);
nand U9190 (N_9190,N_9071,N_9086);
or U9191 (N_9191,N_9097,N_9020);
or U9192 (N_9192,N_9064,N_9005);
or U9193 (N_9193,N_8992,N_9073);
or U9194 (N_9194,N_9046,N_8961);
xor U9195 (N_9195,N_8983,N_8980);
xor U9196 (N_9196,N_8985,N_9100);
nand U9197 (N_9197,N_9024,N_8994);
nand U9198 (N_9198,N_9106,N_8960);
nor U9199 (N_9199,N_9018,N_9056);
or U9200 (N_9200,N_9072,N_9075);
or U9201 (N_9201,N_9017,N_8992);
nand U9202 (N_9202,N_8970,N_8994);
or U9203 (N_9203,N_9016,N_9101);
xor U9204 (N_9204,N_9073,N_9050);
xnor U9205 (N_9205,N_8982,N_9116);
xor U9206 (N_9206,N_9035,N_9080);
or U9207 (N_9207,N_9113,N_9003);
xor U9208 (N_9208,N_8983,N_8986);
nand U9209 (N_9209,N_8983,N_9082);
and U9210 (N_9210,N_9108,N_9065);
and U9211 (N_9211,N_8963,N_9024);
or U9212 (N_9212,N_9025,N_9024);
xor U9213 (N_9213,N_9006,N_9054);
xnor U9214 (N_9214,N_9079,N_8987);
and U9215 (N_9215,N_9093,N_9113);
and U9216 (N_9216,N_9028,N_9073);
and U9217 (N_9217,N_8968,N_9062);
nand U9218 (N_9218,N_9086,N_9066);
nor U9219 (N_9219,N_9087,N_9023);
nand U9220 (N_9220,N_9021,N_8983);
and U9221 (N_9221,N_9117,N_9116);
nor U9222 (N_9222,N_9051,N_8994);
nand U9223 (N_9223,N_9029,N_9034);
or U9224 (N_9224,N_9023,N_9035);
and U9225 (N_9225,N_9096,N_9047);
nor U9226 (N_9226,N_9101,N_8966);
or U9227 (N_9227,N_8975,N_9119);
and U9228 (N_9228,N_9058,N_9045);
and U9229 (N_9229,N_9022,N_8977);
xnor U9230 (N_9230,N_9040,N_9014);
nand U9231 (N_9231,N_8968,N_9047);
nand U9232 (N_9232,N_9059,N_9002);
xnor U9233 (N_9233,N_9117,N_9036);
xor U9234 (N_9234,N_9042,N_9096);
and U9235 (N_9235,N_9105,N_9048);
nor U9236 (N_9236,N_9040,N_9094);
or U9237 (N_9237,N_9074,N_9104);
or U9238 (N_9238,N_9020,N_8961);
nor U9239 (N_9239,N_9018,N_9043);
nor U9240 (N_9240,N_9100,N_9057);
nor U9241 (N_9241,N_8975,N_9006);
nand U9242 (N_9242,N_9091,N_8965);
xnor U9243 (N_9243,N_9011,N_9106);
xnor U9244 (N_9244,N_9067,N_9075);
xor U9245 (N_9245,N_9083,N_9036);
nor U9246 (N_9246,N_8964,N_9114);
nand U9247 (N_9247,N_9028,N_9060);
xnor U9248 (N_9248,N_9090,N_9057);
nand U9249 (N_9249,N_9074,N_9028);
and U9250 (N_9250,N_9044,N_8968);
or U9251 (N_9251,N_8977,N_8989);
xor U9252 (N_9252,N_9113,N_9021);
or U9253 (N_9253,N_9087,N_9093);
and U9254 (N_9254,N_9112,N_9055);
xor U9255 (N_9255,N_9048,N_9041);
xor U9256 (N_9256,N_9078,N_9091);
or U9257 (N_9257,N_9007,N_8973);
xor U9258 (N_9258,N_9009,N_8984);
xor U9259 (N_9259,N_9109,N_8985);
or U9260 (N_9260,N_9009,N_9036);
xnor U9261 (N_9261,N_9045,N_9038);
nand U9262 (N_9262,N_9034,N_8985);
and U9263 (N_9263,N_9093,N_8993);
nor U9264 (N_9264,N_9084,N_8967);
and U9265 (N_9265,N_9098,N_9067);
and U9266 (N_9266,N_8983,N_8974);
or U9267 (N_9267,N_9005,N_9108);
nor U9268 (N_9268,N_9025,N_9103);
nand U9269 (N_9269,N_9077,N_8970);
nand U9270 (N_9270,N_8972,N_9034);
xor U9271 (N_9271,N_8988,N_9045);
nor U9272 (N_9272,N_9103,N_8980);
nor U9273 (N_9273,N_8993,N_9063);
or U9274 (N_9274,N_9070,N_9000);
and U9275 (N_9275,N_8963,N_9012);
and U9276 (N_9276,N_9035,N_9085);
and U9277 (N_9277,N_9002,N_9020);
nand U9278 (N_9278,N_9005,N_9058);
and U9279 (N_9279,N_9060,N_9063);
or U9280 (N_9280,N_9137,N_9196);
and U9281 (N_9281,N_9175,N_9144);
xnor U9282 (N_9282,N_9190,N_9243);
or U9283 (N_9283,N_9200,N_9134);
or U9284 (N_9284,N_9277,N_9252);
or U9285 (N_9285,N_9145,N_9128);
xnor U9286 (N_9286,N_9260,N_9172);
nor U9287 (N_9287,N_9225,N_9279);
and U9288 (N_9288,N_9141,N_9124);
nor U9289 (N_9289,N_9138,N_9136);
or U9290 (N_9290,N_9207,N_9239);
and U9291 (N_9291,N_9266,N_9253);
and U9292 (N_9292,N_9214,N_9149);
nand U9293 (N_9293,N_9259,N_9199);
nor U9294 (N_9294,N_9127,N_9140);
nand U9295 (N_9295,N_9156,N_9157);
nor U9296 (N_9296,N_9262,N_9256);
nand U9297 (N_9297,N_9209,N_9133);
nor U9298 (N_9298,N_9230,N_9125);
or U9299 (N_9299,N_9274,N_9150);
or U9300 (N_9300,N_9130,N_9168);
or U9301 (N_9301,N_9276,N_9258);
xor U9302 (N_9302,N_9120,N_9203);
nand U9303 (N_9303,N_9263,N_9244);
nor U9304 (N_9304,N_9278,N_9220);
nor U9305 (N_9305,N_9142,N_9192);
nand U9306 (N_9306,N_9170,N_9273);
nand U9307 (N_9307,N_9269,N_9186);
xnor U9308 (N_9308,N_9143,N_9227);
nor U9309 (N_9309,N_9183,N_9268);
xnor U9310 (N_9310,N_9224,N_9267);
nand U9311 (N_9311,N_9148,N_9122);
and U9312 (N_9312,N_9213,N_9221);
xnor U9313 (N_9313,N_9189,N_9195);
nor U9314 (N_9314,N_9235,N_9217);
or U9315 (N_9315,N_9158,N_9210);
and U9316 (N_9316,N_9126,N_9238);
or U9317 (N_9317,N_9167,N_9231);
nand U9318 (N_9318,N_9264,N_9160);
or U9319 (N_9319,N_9237,N_9188);
and U9320 (N_9320,N_9194,N_9201);
nand U9321 (N_9321,N_9132,N_9236);
and U9322 (N_9322,N_9161,N_9204);
nor U9323 (N_9323,N_9152,N_9174);
or U9324 (N_9324,N_9228,N_9162);
nor U9325 (N_9325,N_9271,N_9191);
nor U9326 (N_9326,N_9178,N_9255);
xnor U9327 (N_9327,N_9153,N_9173);
xor U9328 (N_9328,N_9206,N_9121);
nand U9329 (N_9329,N_9123,N_9223);
and U9330 (N_9330,N_9275,N_9242);
or U9331 (N_9331,N_9226,N_9169);
or U9332 (N_9332,N_9185,N_9197);
or U9333 (N_9333,N_9184,N_9250);
or U9334 (N_9334,N_9171,N_9205);
or U9335 (N_9335,N_9215,N_9182);
nand U9336 (N_9336,N_9222,N_9146);
nor U9337 (N_9337,N_9257,N_9247);
and U9338 (N_9338,N_9163,N_9216);
and U9339 (N_9339,N_9234,N_9233);
nand U9340 (N_9340,N_9180,N_9166);
or U9341 (N_9341,N_9193,N_9135);
or U9342 (N_9342,N_9202,N_9151);
nand U9343 (N_9343,N_9229,N_9165);
nor U9344 (N_9344,N_9155,N_9147);
or U9345 (N_9345,N_9232,N_9248);
or U9346 (N_9346,N_9176,N_9249);
nand U9347 (N_9347,N_9159,N_9198);
nand U9348 (N_9348,N_9218,N_9154);
xor U9349 (N_9349,N_9187,N_9246);
and U9350 (N_9350,N_9245,N_9219);
or U9351 (N_9351,N_9131,N_9251);
nor U9352 (N_9352,N_9265,N_9272);
or U9353 (N_9353,N_9211,N_9240);
and U9354 (N_9354,N_9139,N_9177);
nand U9355 (N_9355,N_9179,N_9241);
nor U9356 (N_9356,N_9181,N_9254);
or U9357 (N_9357,N_9164,N_9208);
nand U9358 (N_9358,N_9212,N_9129);
nand U9359 (N_9359,N_9261,N_9270);
xnor U9360 (N_9360,N_9246,N_9214);
and U9361 (N_9361,N_9245,N_9153);
nand U9362 (N_9362,N_9169,N_9238);
nor U9363 (N_9363,N_9215,N_9150);
or U9364 (N_9364,N_9182,N_9217);
or U9365 (N_9365,N_9176,N_9129);
nor U9366 (N_9366,N_9186,N_9182);
and U9367 (N_9367,N_9248,N_9270);
and U9368 (N_9368,N_9235,N_9177);
nor U9369 (N_9369,N_9272,N_9279);
and U9370 (N_9370,N_9259,N_9163);
or U9371 (N_9371,N_9202,N_9253);
and U9372 (N_9372,N_9256,N_9275);
nor U9373 (N_9373,N_9134,N_9249);
and U9374 (N_9374,N_9141,N_9176);
nor U9375 (N_9375,N_9174,N_9201);
nor U9376 (N_9376,N_9248,N_9161);
xor U9377 (N_9377,N_9210,N_9278);
nor U9378 (N_9378,N_9172,N_9123);
xnor U9379 (N_9379,N_9210,N_9192);
xnor U9380 (N_9380,N_9173,N_9222);
or U9381 (N_9381,N_9242,N_9124);
or U9382 (N_9382,N_9197,N_9150);
nor U9383 (N_9383,N_9263,N_9276);
xor U9384 (N_9384,N_9220,N_9196);
and U9385 (N_9385,N_9124,N_9266);
xnor U9386 (N_9386,N_9225,N_9217);
nand U9387 (N_9387,N_9191,N_9205);
and U9388 (N_9388,N_9163,N_9239);
and U9389 (N_9389,N_9276,N_9140);
nor U9390 (N_9390,N_9171,N_9187);
and U9391 (N_9391,N_9214,N_9183);
nor U9392 (N_9392,N_9194,N_9176);
nor U9393 (N_9393,N_9228,N_9157);
and U9394 (N_9394,N_9172,N_9157);
nand U9395 (N_9395,N_9221,N_9143);
and U9396 (N_9396,N_9140,N_9246);
nand U9397 (N_9397,N_9166,N_9131);
xnor U9398 (N_9398,N_9229,N_9137);
xor U9399 (N_9399,N_9160,N_9193);
nor U9400 (N_9400,N_9243,N_9193);
or U9401 (N_9401,N_9179,N_9130);
xor U9402 (N_9402,N_9186,N_9175);
nor U9403 (N_9403,N_9255,N_9121);
nor U9404 (N_9404,N_9149,N_9239);
or U9405 (N_9405,N_9213,N_9130);
or U9406 (N_9406,N_9173,N_9148);
xor U9407 (N_9407,N_9219,N_9171);
or U9408 (N_9408,N_9146,N_9258);
nor U9409 (N_9409,N_9123,N_9213);
or U9410 (N_9410,N_9218,N_9178);
xnor U9411 (N_9411,N_9215,N_9220);
or U9412 (N_9412,N_9263,N_9169);
nor U9413 (N_9413,N_9213,N_9250);
xnor U9414 (N_9414,N_9163,N_9192);
nor U9415 (N_9415,N_9226,N_9124);
or U9416 (N_9416,N_9195,N_9218);
and U9417 (N_9417,N_9255,N_9182);
and U9418 (N_9418,N_9217,N_9150);
or U9419 (N_9419,N_9230,N_9190);
nand U9420 (N_9420,N_9168,N_9277);
nand U9421 (N_9421,N_9204,N_9240);
or U9422 (N_9422,N_9254,N_9163);
or U9423 (N_9423,N_9187,N_9154);
or U9424 (N_9424,N_9170,N_9155);
and U9425 (N_9425,N_9230,N_9134);
xor U9426 (N_9426,N_9219,N_9195);
and U9427 (N_9427,N_9204,N_9170);
and U9428 (N_9428,N_9219,N_9158);
nor U9429 (N_9429,N_9168,N_9278);
xnor U9430 (N_9430,N_9279,N_9172);
and U9431 (N_9431,N_9154,N_9129);
xor U9432 (N_9432,N_9183,N_9252);
xor U9433 (N_9433,N_9256,N_9162);
xnor U9434 (N_9434,N_9247,N_9176);
nor U9435 (N_9435,N_9173,N_9223);
or U9436 (N_9436,N_9232,N_9221);
nand U9437 (N_9437,N_9234,N_9251);
xnor U9438 (N_9438,N_9152,N_9143);
and U9439 (N_9439,N_9144,N_9257);
or U9440 (N_9440,N_9405,N_9385);
nand U9441 (N_9441,N_9436,N_9383);
xor U9442 (N_9442,N_9280,N_9423);
and U9443 (N_9443,N_9340,N_9332);
nor U9444 (N_9444,N_9323,N_9381);
nor U9445 (N_9445,N_9422,N_9439);
or U9446 (N_9446,N_9283,N_9403);
nand U9447 (N_9447,N_9408,N_9398);
nor U9448 (N_9448,N_9367,N_9404);
xnor U9449 (N_9449,N_9418,N_9378);
or U9450 (N_9450,N_9309,N_9434);
nand U9451 (N_9451,N_9391,N_9437);
or U9452 (N_9452,N_9435,N_9400);
and U9453 (N_9453,N_9379,N_9413);
or U9454 (N_9454,N_9319,N_9352);
or U9455 (N_9455,N_9371,N_9397);
or U9456 (N_9456,N_9313,N_9329);
and U9457 (N_9457,N_9353,N_9426);
xor U9458 (N_9458,N_9412,N_9382);
or U9459 (N_9459,N_9419,N_9365);
or U9460 (N_9460,N_9330,N_9284);
and U9461 (N_9461,N_9317,N_9303);
xor U9462 (N_9462,N_9374,N_9314);
and U9463 (N_9463,N_9392,N_9356);
xor U9464 (N_9464,N_9306,N_9399);
or U9465 (N_9465,N_9344,N_9429);
and U9466 (N_9466,N_9351,N_9411);
and U9467 (N_9467,N_9302,N_9376);
or U9468 (N_9468,N_9363,N_9281);
nand U9469 (N_9469,N_9320,N_9359);
and U9470 (N_9470,N_9354,N_9285);
nand U9471 (N_9471,N_9324,N_9312);
xor U9472 (N_9472,N_9318,N_9343);
and U9473 (N_9473,N_9388,N_9282);
nand U9474 (N_9474,N_9311,N_9427);
and U9475 (N_9475,N_9395,N_9360);
nor U9476 (N_9476,N_9377,N_9364);
xor U9477 (N_9477,N_9289,N_9362);
nor U9478 (N_9478,N_9420,N_9372);
nor U9479 (N_9479,N_9328,N_9428);
or U9480 (N_9480,N_9294,N_9401);
or U9481 (N_9481,N_9348,N_9361);
nand U9482 (N_9482,N_9389,N_9342);
or U9483 (N_9483,N_9407,N_9296);
nand U9484 (N_9484,N_9335,N_9357);
nor U9485 (N_9485,N_9415,N_9402);
xnor U9486 (N_9486,N_9396,N_9310);
nand U9487 (N_9487,N_9373,N_9307);
and U9488 (N_9488,N_9358,N_9390);
or U9489 (N_9489,N_9298,N_9325);
nand U9490 (N_9490,N_9286,N_9414);
and U9491 (N_9491,N_9416,N_9337);
nand U9492 (N_9492,N_9386,N_9369);
or U9493 (N_9493,N_9326,N_9336);
nor U9494 (N_9494,N_9305,N_9433);
nand U9495 (N_9495,N_9299,N_9291);
nor U9496 (N_9496,N_9316,N_9301);
or U9497 (N_9497,N_9295,N_9315);
nand U9498 (N_9498,N_9346,N_9304);
nand U9499 (N_9499,N_9293,N_9350);
or U9500 (N_9500,N_9417,N_9334);
and U9501 (N_9501,N_9421,N_9287);
or U9502 (N_9502,N_9394,N_9322);
and U9503 (N_9503,N_9333,N_9424);
nor U9504 (N_9504,N_9380,N_9368);
and U9505 (N_9505,N_9366,N_9339);
nand U9506 (N_9506,N_9425,N_9290);
nor U9507 (N_9507,N_9288,N_9327);
xor U9508 (N_9508,N_9292,N_9338);
nand U9509 (N_9509,N_9375,N_9430);
xnor U9510 (N_9510,N_9410,N_9438);
and U9511 (N_9511,N_9431,N_9308);
and U9512 (N_9512,N_9355,N_9300);
nand U9513 (N_9513,N_9432,N_9406);
or U9514 (N_9514,N_9341,N_9384);
nor U9515 (N_9515,N_9331,N_9349);
and U9516 (N_9516,N_9345,N_9321);
xor U9517 (N_9517,N_9393,N_9370);
xnor U9518 (N_9518,N_9409,N_9297);
nor U9519 (N_9519,N_9347,N_9387);
nand U9520 (N_9520,N_9405,N_9292);
nor U9521 (N_9521,N_9326,N_9390);
or U9522 (N_9522,N_9346,N_9353);
nor U9523 (N_9523,N_9427,N_9296);
nor U9524 (N_9524,N_9288,N_9286);
nand U9525 (N_9525,N_9375,N_9432);
xnor U9526 (N_9526,N_9291,N_9344);
or U9527 (N_9527,N_9331,N_9335);
xor U9528 (N_9528,N_9386,N_9290);
xnor U9529 (N_9529,N_9379,N_9292);
nor U9530 (N_9530,N_9347,N_9297);
nor U9531 (N_9531,N_9379,N_9352);
nand U9532 (N_9532,N_9411,N_9368);
nand U9533 (N_9533,N_9420,N_9320);
nand U9534 (N_9534,N_9341,N_9313);
and U9535 (N_9535,N_9329,N_9325);
nor U9536 (N_9536,N_9295,N_9385);
nand U9537 (N_9537,N_9316,N_9421);
nor U9538 (N_9538,N_9332,N_9309);
and U9539 (N_9539,N_9343,N_9351);
nand U9540 (N_9540,N_9422,N_9342);
and U9541 (N_9541,N_9298,N_9385);
xnor U9542 (N_9542,N_9328,N_9340);
or U9543 (N_9543,N_9373,N_9365);
and U9544 (N_9544,N_9344,N_9297);
and U9545 (N_9545,N_9356,N_9401);
and U9546 (N_9546,N_9318,N_9422);
and U9547 (N_9547,N_9344,N_9412);
nand U9548 (N_9548,N_9399,N_9421);
xnor U9549 (N_9549,N_9386,N_9306);
nor U9550 (N_9550,N_9327,N_9386);
xor U9551 (N_9551,N_9389,N_9374);
xnor U9552 (N_9552,N_9376,N_9370);
and U9553 (N_9553,N_9342,N_9297);
nand U9554 (N_9554,N_9348,N_9383);
xor U9555 (N_9555,N_9361,N_9333);
nor U9556 (N_9556,N_9359,N_9376);
nor U9557 (N_9557,N_9368,N_9388);
or U9558 (N_9558,N_9358,N_9383);
xor U9559 (N_9559,N_9357,N_9427);
nand U9560 (N_9560,N_9374,N_9376);
nand U9561 (N_9561,N_9328,N_9392);
and U9562 (N_9562,N_9386,N_9291);
nor U9563 (N_9563,N_9291,N_9372);
nand U9564 (N_9564,N_9289,N_9283);
nand U9565 (N_9565,N_9310,N_9299);
nor U9566 (N_9566,N_9337,N_9315);
xor U9567 (N_9567,N_9329,N_9349);
or U9568 (N_9568,N_9350,N_9307);
xor U9569 (N_9569,N_9286,N_9416);
xor U9570 (N_9570,N_9358,N_9352);
and U9571 (N_9571,N_9415,N_9420);
nand U9572 (N_9572,N_9356,N_9385);
xor U9573 (N_9573,N_9420,N_9345);
and U9574 (N_9574,N_9400,N_9380);
nand U9575 (N_9575,N_9325,N_9337);
xor U9576 (N_9576,N_9293,N_9404);
nor U9577 (N_9577,N_9408,N_9315);
nand U9578 (N_9578,N_9366,N_9415);
nor U9579 (N_9579,N_9431,N_9395);
xor U9580 (N_9580,N_9395,N_9411);
nor U9581 (N_9581,N_9347,N_9287);
and U9582 (N_9582,N_9281,N_9431);
nand U9583 (N_9583,N_9385,N_9317);
and U9584 (N_9584,N_9400,N_9438);
or U9585 (N_9585,N_9327,N_9373);
nor U9586 (N_9586,N_9402,N_9343);
or U9587 (N_9587,N_9369,N_9418);
or U9588 (N_9588,N_9382,N_9347);
nand U9589 (N_9589,N_9407,N_9307);
and U9590 (N_9590,N_9280,N_9375);
nand U9591 (N_9591,N_9345,N_9382);
nand U9592 (N_9592,N_9374,N_9331);
or U9593 (N_9593,N_9351,N_9287);
xor U9594 (N_9594,N_9408,N_9321);
nor U9595 (N_9595,N_9358,N_9366);
nand U9596 (N_9596,N_9296,N_9364);
or U9597 (N_9597,N_9339,N_9391);
nand U9598 (N_9598,N_9356,N_9285);
and U9599 (N_9599,N_9330,N_9424);
xor U9600 (N_9600,N_9500,N_9561);
nand U9601 (N_9601,N_9595,N_9507);
or U9602 (N_9602,N_9453,N_9526);
nand U9603 (N_9603,N_9505,N_9599);
nand U9604 (N_9604,N_9522,N_9537);
nand U9605 (N_9605,N_9482,N_9539);
nor U9606 (N_9606,N_9553,N_9536);
or U9607 (N_9607,N_9502,N_9441);
nor U9608 (N_9608,N_9517,N_9558);
nand U9609 (N_9609,N_9503,N_9549);
or U9610 (N_9610,N_9470,N_9544);
nor U9611 (N_9611,N_9473,N_9515);
and U9612 (N_9612,N_9475,N_9509);
nand U9613 (N_9613,N_9487,N_9566);
and U9614 (N_9614,N_9510,N_9560);
or U9615 (N_9615,N_9591,N_9569);
nand U9616 (N_9616,N_9581,N_9585);
nand U9617 (N_9617,N_9512,N_9520);
or U9618 (N_9618,N_9449,N_9496);
nor U9619 (N_9619,N_9546,N_9547);
xor U9620 (N_9620,N_9493,N_9456);
and U9621 (N_9621,N_9538,N_9523);
or U9622 (N_9622,N_9540,N_9463);
xor U9623 (N_9623,N_9532,N_9511);
xor U9624 (N_9624,N_9490,N_9469);
and U9625 (N_9625,N_9545,N_9530);
nand U9626 (N_9626,N_9527,N_9455);
xnor U9627 (N_9627,N_9444,N_9506);
and U9628 (N_9628,N_9471,N_9548);
xor U9629 (N_9629,N_9529,N_9590);
nand U9630 (N_9630,N_9461,N_9524);
nand U9631 (N_9631,N_9594,N_9464);
or U9632 (N_9632,N_9584,N_9534);
xnor U9633 (N_9633,N_9459,N_9488);
nor U9634 (N_9634,N_9597,N_9516);
nor U9635 (N_9635,N_9443,N_9592);
and U9636 (N_9636,N_9467,N_9484);
nor U9637 (N_9637,N_9447,N_9562);
xnor U9638 (N_9638,N_9448,N_9497);
and U9639 (N_9639,N_9450,N_9579);
or U9640 (N_9640,N_9565,N_9474);
or U9641 (N_9641,N_9481,N_9542);
or U9642 (N_9642,N_9472,N_9468);
or U9643 (N_9643,N_9479,N_9483);
xor U9644 (N_9644,N_9452,N_9501);
xnor U9645 (N_9645,N_9596,N_9589);
nand U9646 (N_9646,N_9478,N_9578);
or U9647 (N_9647,N_9580,N_9531);
xnor U9648 (N_9648,N_9513,N_9462);
and U9649 (N_9649,N_9573,N_9528);
and U9650 (N_9650,N_9586,N_9550);
nor U9651 (N_9651,N_9535,N_9466);
and U9652 (N_9652,N_9567,N_9489);
nor U9653 (N_9653,N_9495,N_9559);
nand U9654 (N_9654,N_9445,N_9525);
nand U9655 (N_9655,N_9518,N_9477);
and U9656 (N_9656,N_9451,N_9494);
nor U9657 (N_9657,N_9446,N_9454);
and U9658 (N_9658,N_9555,N_9588);
or U9659 (N_9659,N_9563,N_9491);
or U9660 (N_9660,N_9485,N_9486);
or U9661 (N_9661,N_9521,N_9577);
and U9662 (N_9662,N_9572,N_9504);
or U9663 (N_9663,N_9498,N_9465);
and U9664 (N_9664,N_9557,N_9568);
xnor U9665 (N_9665,N_9554,N_9582);
or U9666 (N_9666,N_9458,N_9440);
and U9667 (N_9667,N_9514,N_9480);
and U9668 (N_9668,N_9574,N_9499);
nand U9669 (N_9669,N_9575,N_9552);
nor U9670 (N_9670,N_9476,N_9508);
nor U9671 (N_9671,N_9457,N_9593);
or U9672 (N_9672,N_9543,N_9533);
nor U9673 (N_9673,N_9541,N_9570);
nor U9674 (N_9674,N_9583,N_9519);
nor U9675 (N_9675,N_9551,N_9564);
nor U9676 (N_9676,N_9442,N_9587);
or U9677 (N_9677,N_9598,N_9576);
and U9678 (N_9678,N_9460,N_9492);
nand U9679 (N_9679,N_9556,N_9571);
and U9680 (N_9680,N_9528,N_9544);
xor U9681 (N_9681,N_9522,N_9466);
nand U9682 (N_9682,N_9557,N_9493);
or U9683 (N_9683,N_9588,N_9579);
and U9684 (N_9684,N_9444,N_9553);
or U9685 (N_9685,N_9516,N_9588);
xor U9686 (N_9686,N_9562,N_9445);
xnor U9687 (N_9687,N_9515,N_9532);
or U9688 (N_9688,N_9522,N_9586);
nand U9689 (N_9689,N_9581,N_9502);
and U9690 (N_9690,N_9532,N_9553);
or U9691 (N_9691,N_9526,N_9566);
or U9692 (N_9692,N_9520,N_9456);
nor U9693 (N_9693,N_9597,N_9488);
nand U9694 (N_9694,N_9585,N_9595);
nor U9695 (N_9695,N_9594,N_9504);
xnor U9696 (N_9696,N_9483,N_9453);
or U9697 (N_9697,N_9553,N_9521);
xnor U9698 (N_9698,N_9576,N_9559);
xnor U9699 (N_9699,N_9598,N_9509);
nor U9700 (N_9700,N_9446,N_9519);
nor U9701 (N_9701,N_9556,N_9521);
nand U9702 (N_9702,N_9485,N_9463);
nor U9703 (N_9703,N_9552,N_9456);
xnor U9704 (N_9704,N_9463,N_9538);
and U9705 (N_9705,N_9474,N_9564);
nor U9706 (N_9706,N_9499,N_9563);
or U9707 (N_9707,N_9526,N_9493);
xnor U9708 (N_9708,N_9563,N_9477);
nand U9709 (N_9709,N_9458,N_9462);
or U9710 (N_9710,N_9459,N_9485);
and U9711 (N_9711,N_9513,N_9570);
nand U9712 (N_9712,N_9503,N_9449);
nand U9713 (N_9713,N_9441,N_9524);
and U9714 (N_9714,N_9444,N_9598);
or U9715 (N_9715,N_9486,N_9594);
or U9716 (N_9716,N_9443,N_9577);
xor U9717 (N_9717,N_9538,N_9593);
nor U9718 (N_9718,N_9442,N_9511);
xor U9719 (N_9719,N_9578,N_9459);
xor U9720 (N_9720,N_9576,N_9528);
and U9721 (N_9721,N_9501,N_9497);
nand U9722 (N_9722,N_9480,N_9528);
xnor U9723 (N_9723,N_9448,N_9596);
and U9724 (N_9724,N_9492,N_9579);
nor U9725 (N_9725,N_9494,N_9517);
and U9726 (N_9726,N_9581,N_9501);
or U9727 (N_9727,N_9486,N_9598);
nand U9728 (N_9728,N_9480,N_9532);
xor U9729 (N_9729,N_9510,N_9580);
nor U9730 (N_9730,N_9445,N_9469);
nand U9731 (N_9731,N_9588,N_9477);
nor U9732 (N_9732,N_9553,N_9506);
and U9733 (N_9733,N_9570,N_9523);
and U9734 (N_9734,N_9550,N_9564);
nor U9735 (N_9735,N_9494,N_9575);
and U9736 (N_9736,N_9545,N_9495);
and U9737 (N_9737,N_9564,N_9498);
and U9738 (N_9738,N_9445,N_9450);
nand U9739 (N_9739,N_9544,N_9514);
and U9740 (N_9740,N_9450,N_9520);
or U9741 (N_9741,N_9443,N_9586);
and U9742 (N_9742,N_9531,N_9476);
nand U9743 (N_9743,N_9454,N_9554);
and U9744 (N_9744,N_9587,N_9507);
xor U9745 (N_9745,N_9503,N_9523);
nor U9746 (N_9746,N_9529,N_9540);
xor U9747 (N_9747,N_9453,N_9566);
or U9748 (N_9748,N_9582,N_9596);
or U9749 (N_9749,N_9544,N_9462);
nor U9750 (N_9750,N_9566,N_9493);
and U9751 (N_9751,N_9490,N_9499);
nor U9752 (N_9752,N_9592,N_9473);
or U9753 (N_9753,N_9519,N_9549);
nand U9754 (N_9754,N_9551,N_9467);
or U9755 (N_9755,N_9486,N_9483);
nor U9756 (N_9756,N_9445,N_9566);
and U9757 (N_9757,N_9472,N_9544);
or U9758 (N_9758,N_9571,N_9504);
or U9759 (N_9759,N_9505,N_9503);
xor U9760 (N_9760,N_9712,N_9609);
xor U9761 (N_9761,N_9752,N_9616);
and U9762 (N_9762,N_9690,N_9678);
nand U9763 (N_9763,N_9756,N_9733);
xor U9764 (N_9764,N_9699,N_9742);
nand U9765 (N_9765,N_9611,N_9704);
xor U9766 (N_9766,N_9727,N_9757);
and U9767 (N_9767,N_9643,N_9716);
and U9768 (N_9768,N_9746,N_9607);
or U9769 (N_9769,N_9653,N_9606);
or U9770 (N_9770,N_9696,N_9626);
xnor U9771 (N_9771,N_9750,N_9655);
nor U9772 (N_9772,N_9738,N_9623);
xnor U9773 (N_9773,N_9720,N_9633);
or U9774 (N_9774,N_9627,N_9753);
or U9775 (N_9775,N_9719,N_9714);
nor U9776 (N_9776,N_9689,N_9702);
or U9777 (N_9777,N_9637,N_9730);
nor U9778 (N_9778,N_9735,N_9620);
nor U9779 (N_9779,N_9644,N_9603);
nor U9780 (N_9780,N_9686,N_9651);
and U9781 (N_9781,N_9741,N_9658);
or U9782 (N_9782,N_9662,N_9649);
or U9783 (N_9783,N_9729,N_9688);
nand U9784 (N_9784,N_9635,N_9639);
nand U9785 (N_9785,N_9724,N_9731);
or U9786 (N_9786,N_9612,N_9671);
xnor U9787 (N_9787,N_9692,N_9661);
and U9788 (N_9788,N_9695,N_9728);
nor U9789 (N_9789,N_9749,N_9706);
and U9790 (N_9790,N_9732,N_9715);
nand U9791 (N_9791,N_9657,N_9717);
and U9792 (N_9792,N_9605,N_9600);
and U9793 (N_9793,N_9648,N_9755);
nor U9794 (N_9794,N_9659,N_9745);
and U9795 (N_9795,N_9647,N_9718);
or U9796 (N_9796,N_9632,N_9666);
xor U9797 (N_9797,N_9621,N_9602);
nor U9798 (N_9798,N_9721,N_9613);
and U9799 (N_9799,N_9663,N_9664);
and U9800 (N_9800,N_9673,N_9675);
xor U9801 (N_9801,N_9610,N_9665);
xnor U9802 (N_9802,N_9744,N_9711);
nand U9803 (N_9803,N_9725,N_9748);
nand U9804 (N_9804,N_9685,N_9737);
nand U9805 (N_9805,N_9629,N_9743);
and U9806 (N_9806,N_9604,N_9669);
nand U9807 (N_9807,N_9670,N_9646);
and U9808 (N_9808,N_9687,N_9624);
or U9809 (N_9809,N_9722,N_9740);
xor U9810 (N_9810,N_9608,N_9638);
nor U9811 (N_9811,N_9619,N_9680);
nand U9812 (N_9812,N_9751,N_9694);
and U9813 (N_9813,N_9734,N_9754);
and U9814 (N_9814,N_9640,N_9622);
and U9815 (N_9815,N_9708,N_9630);
xor U9816 (N_9816,N_9652,N_9726);
nand U9817 (N_9817,N_9723,N_9677);
nor U9818 (N_9818,N_9709,N_9713);
nor U9819 (N_9819,N_9682,N_9736);
xor U9820 (N_9820,N_9618,N_9698);
xnor U9821 (N_9821,N_9703,N_9674);
xnor U9822 (N_9822,N_9628,N_9693);
nor U9823 (N_9823,N_9668,N_9683);
xnor U9824 (N_9824,N_9697,N_9701);
nor U9825 (N_9825,N_9700,N_9667);
and U9826 (N_9826,N_9691,N_9617);
xnor U9827 (N_9827,N_9615,N_9747);
and U9828 (N_9828,N_9631,N_9705);
or U9829 (N_9829,N_9641,N_9707);
nand U9830 (N_9830,N_9660,N_9614);
nor U9831 (N_9831,N_9601,N_9676);
xor U9832 (N_9832,N_9759,N_9758);
xnor U9833 (N_9833,N_9654,N_9710);
nand U9834 (N_9834,N_9625,N_9642);
nor U9835 (N_9835,N_9634,N_9636);
and U9836 (N_9836,N_9739,N_9684);
and U9837 (N_9837,N_9650,N_9681);
nor U9838 (N_9838,N_9656,N_9672);
nand U9839 (N_9839,N_9679,N_9645);
nand U9840 (N_9840,N_9671,N_9730);
and U9841 (N_9841,N_9605,N_9643);
nand U9842 (N_9842,N_9745,N_9728);
or U9843 (N_9843,N_9755,N_9669);
nor U9844 (N_9844,N_9642,N_9732);
nand U9845 (N_9845,N_9727,N_9627);
or U9846 (N_9846,N_9615,N_9730);
nor U9847 (N_9847,N_9606,N_9737);
nor U9848 (N_9848,N_9699,N_9700);
and U9849 (N_9849,N_9758,N_9639);
or U9850 (N_9850,N_9679,N_9750);
nor U9851 (N_9851,N_9611,N_9681);
xnor U9852 (N_9852,N_9748,N_9678);
xor U9853 (N_9853,N_9722,N_9752);
xor U9854 (N_9854,N_9688,N_9702);
xor U9855 (N_9855,N_9733,N_9727);
nand U9856 (N_9856,N_9706,N_9710);
nand U9857 (N_9857,N_9663,N_9701);
nor U9858 (N_9858,N_9730,N_9706);
nor U9859 (N_9859,N_9676,N_9658);
or U9860 (N_9860,N_9606,N_9673);
nand U9861 (N_9861,N_9668,N_9728);
or U9862 (N_9862,N_9719,N_9726);
xnor U9863 (N_9863,N_9753,N_9714);
xor U9864 (N_9864,N_9671,N_9684);
nor U9865 (N_9865,N_9688,N_9673);
nor U9866 (N_9866,N_9741,N_9655);
and U9867 (N_9867,N_9698,N_9600);
and U9868 (N_9868,N_9617,N_9727);
or U9869 (N_9869,N_9604,N_9654);
or U9870 (N_9870,N_9747,N_9731);
nand U9871 (N_9871,N_9745,N_9620);
and U9872 (N_9872,N_9655,N_9686);
or U9873 (N_9873,N_9725,N_9632);
nand U9874 (N_9874,N_9619,N_9648);
nor U9875 (N_9875,N_9634,N_9742);
nor U9876 (N_9876,N_9698,N_9728);
xnor U9877 (N_9877,N_9692,N_9618);
xnor U9878 (N_9878,N_9646,N_9655);
nor U9879 (N_9879,N_9696,N_9712);
and U9880 (N_9880,N_9719,N_9693);
or U9881 (N_9881,N_9754,N_9658);
and U9882 (N_9882,N_9750,N_9721);
nor U9883 (N_9883,N_9659,N_9649);
nand U9884 (N_9884,N_9629,N_9607);
and U9885 (N_9885,N_9650,N_9754);
and U9886 (N_9886,N_9716,N_9740);
and U9887 (N_9887,N_9600,N_9625);
or U9888 (N_9888,N_9676,N_9725);
xor U9889 (N_9889,N_9714,N_9755);
or U9890 (N_9890,N_9615,N_9708);
nor U9891 (N_9891,N_9742,N_9692);
and U9892 (N_9892,N_9619,N_9690);
xnor U9893 (N_9893,N_9758,N_9755);
and U9894 (N_9894,N_9634,N_9746);
nand U9895 (N_9895,N_9666,N_9636);
xor U9896 (N_9896,N_9622,N_9712);
nand U9897 (N_9897,N_9667,N_9651);
xnor U9898 (N_9898,N_9683,N_9648);
xor U9899 (N_9899,N_9679,N_9662);
nor U9900 (N_9900,N_9646,N_9618);
or U9901 (N_9901,N_9721,N_9693);
and U9902 (N_9902,N_9731,N_9686);
and U9903 (N_9903,N_9632,N_9613);
and U9904 (N_9904,N_9609,N_9692);
xnor U9905 (N_9905,N_9618,N_9664);
nor U9906 (N_9906,N_9737,N_9727);
nor U9907 (N_9907,N_9716,N_9750);
nor U9908 (N_9908,N_9621,N_9630);
nor U9909 (N_9909,N_9732,N_9694);
or U9910 (N_9910,N_9740,N_9689);
or U9911 (N_9911,N_9617,N_9625);
xor U9912 (N_9912,N_9719,N_9603);
or U9913 (N_9913,N_9642,N_9682);
or U9914 (N_9914,N_9631,N_9662);
and U9915 (N_9915,N_9748,N_9611);
nand U9916 (N_9916,N_9700,N_9690);
nand U9917 (N_9917,N_9723,N_9737);
or U9918 (N_9918,N_9660,N_9701);
nand U9919 (N_9919,N_9640,N_9632);
nand U9920 (N_9920,N_9775,N_9889);
nor U9921 (N_9921,N_9895,N_9865);
or U9922 (N_9922,N_9811,N_9887);
nor U9923 (N_9923,N_9906,N_9762);
or U9924 (N_9924,N_9820,N_9819);
nand U9925 (N_9925,N_9872,N_9910);
nand U9926 (N_9926,N_9907,N_9912);
nand U9927 (N_9927,N_9822,N_9783);
nor U9928 (N_9928,N_9792,N_9899);
xnor U9929 (N_9929,N_9799,N_9826);
and U9930 (N_9930,N_9830,N_9864);
or U9931 (N_9931,N_9852,N_9903);
or U9932 (N_9932,N_9857,N_9861);
or U9933 (N_9933,N_9888,N_9883);
nand U9934 (N_9934,N_9781,N_9904);
and U9935 (N_9935,N_9840,N_9770);
nor U9936 (N_9936,N_9841,N_9782);
nor U9937 (N_9937,N_9764,N_9765);
xnor U9938 (N_9938,N_9803,N_9870);
xor U9939 (N_9939,N_9867,N_9854);
or U9940 (N_9940,N_9890,N_9869);
and U9941 (N_9941,N_9821,N_9886);
nor U9942 (N_9942,N_9800,N_9901);
nor U9943 (N_9943,N_9892,N_9860);
nand U9944 (N_9944,N_9918,N_9900);
xor U9945 (N_9945,N_9894,N_9838);
xnor U9946 (N_9946,N_9911,N_9847);
xor U9947 (N_9947,N_9810,N_9813);
xor U9948 (N_9948,N_9913,N_9815);
and U9949 (N_9949,N_9881,N_9795);
xnor U9950 (N_9950,N_9808,N_9804);
nand U9951 (N_9951,N_9885,N_9824);
nand U9952 (N_9952,N_9849,N_9837);
and U9953 (N_9953,N_9862,N_9761);
xnor U9954 (N_9954,N_9863,N_9916);
nor U9955 (N_9955,N_9853,N_9835);
and U9956 (N_9956,N_9891,N_9798);
nor U9957 (N_9957,N_9796,N_9794);
or U9958 (N_9958,N_9790,N_9914);
nand U9959 (N_9959,N_9766,N_9768);
or U9960 (N_9960,N_9919,N_9845);
and U9961 (N_9961,N_9801,N_9915);
nand U9962 (N_9962,N_9877,N_9848);
and U9963 (N_9963,N_9873,N_9784);
xor U9964 (N_9964,N_9880,N_9823);
and U9965 (N_9965,N_9855,N_9909);
xnor U9966 (N_9966,N_9763,N_9844);
or U9967 (N_9967,N_9831,N_9769);
and U9968 (N_9968,N_9917,N_9875);
xnor U9969 (N_9969,N_9817,N_9874);
nor U9970 (N_9970,N_9818,N_9876);
xnor U9971 (N_9971,N_9898,N_9825);
nor U9972 (N_9972,N_9882,N_9905);
and U9973 (N_9973,N_9805,N_9828);
or U9974 (N_9974,N_9786,N_9858);
and U9975 (N_9975,N_9832,N_9773);
nand U9976 (N_9976,N_9776,N_9787);
xnor U9977 (N_9977,N_9908,N_9779);
or U9978 (N_9978,N_9829,N_9791);
nor U9979 (N_9979,N_9816,N_9851);
nand U9980 (N_9980,N_9850,N_9859);
xnor U9981 (N_9981,N_9897,N_9893);
and U9982 (N_9982,N_9902,N_9789);
or U9983 (N_9983,N_9785,N_9767);
nor U9984 (N_9984,N_9884,N_9793);
xor U9985 (N_9985,N_9760,N_9802);
nand U9986 (N_9986,N_9797,N_9809);
nand U9987 (N_9987,N_9812,N_9780);
xnor U9988 (N_9988,N_9788,N_9806);
xor U9989 (N_9989,N_9807,N_9839);
nand U9990 (N_9990,N_9833,N_9771);
xnor U9991 (N_9991,N_9778,N_9846);
or U9992 (N_9992,N_9834,N_9777);
xor U9993 (N_9993,N_9856,N_9871);
and U9994 (N_9994,N_9827,N_9836);
nand U9995 (N_9995,N_9842,N_9772);
and U9996 (N_9996,N_9879,N_9896);
and U9997 (N_9997,N_9843,N_9814);
and U9998 (N_9998,N_9866,N_9868);
nor U9999 (N_9999,N_9774,N_9878);
or U10000 (N_10000,N_9897,N_9760);
xnor U10001 (N_10001,N_9871,N_9845);
and U10002 (N_10002,N_9812,N_9883);
and U10003 (N_10003,N_9877,N_9897);
or U10004 (N_10004,N_9775,N_9814);
or U10005 (N_10005,N_9797,N_9815);
xor U10006 (N_10006,N_9827,N_9829);
nor U10007 (N_10007,N_9845,N_9908);
xnor U10008 (N_10008,N_9820,N_9903);
nand U10009 (N_10009,N_9909,N_9901);
xor U10010 (N_10010,N_9853,N_9833);
and U10011 (N_10011,N_9846,N_9762);
nor U10012 (N_10012,N_9824,N_9877);
and U10013 (N_10013,N_9817,N_9788);
nor U10014 (N_10014,N_9784,N_9789);
xnor U10015 (N_10015,N_9908,N_9887);
or U10016 (N_10016,N_9801,N_9895);
and U10017 (N_10017,N_9874,N_9821);
nor U10018 (N_10018,N_9774,N_9795);
or U10019 (N_10019,N_9807,N_9789);
or U10020 (N_10020,N_9805,N_9774);
nand U10021 (N_10021,N_9914,N_9792);
or U10022 (N_10022,N_9894,N_9780);
nand U10023 (N_10023,N_9766,N_9908);
nor U10024 (N_10024,N_9908,N_9904);
nor U10025 (N_10025,N_9814,N_9836);
xnor U10026 (N_10026,N_9822,N_9873);
and U10027 (N_10027,N_9760,N_9819);
and U10028 (N_10028,N_9890,N_9918);
nand U10029 (N_10029,N_9767,N_9789);
and U10030 (N_10030,N_9850,N_9917);
or U10031 (N_10031,N_9866,N_9863);
and U10032 (N_10032,N_9859,N_9833);
nor U10033 (N_10033,N_9826,N_9825);
xnor U10034 (N_10034,N_9895,N_9849);
and U10035 (N_10035,N_9882,N_9885);
and U10036 (N_10036,N_9862,N_9908);
nand U10037 (N_10037,N_9803,N_9891);
and U10038 (N_10038,N_9817,N_9882);
nor U10039 (N_10039,N_9883,N_9902);
nor U10040 (N_10040,N_9858,N_9917);
or U10041 (N_10041,N_9811,N_9782);
nor U10042 (N_10042,N_9911,N_9870);
nand U10043 (N_10043,N_9874,N_9781);
nand U10044 (N_10044,N_9778,N_9771);
or U10045 (N_10045,N_9877,N_9833);
nand U10046 (N_10046,N_9855,N_9875);
and U10047 (N_10047,N_9823,N_9830);
nor U10048 (N_10048,N_9769,N_9802);
nor U10049 (N_10049,N_9776,N_9883);
nor U10050 (N_10050,N_9782,N_9873);
and U10051 (N_10051,N_9798,N_9818);
or U10052 (N_10052,N_9766,N_9835);
xnor U10053 (N_10053,N_9779,N_9899);
and U10054 (N_10054,N_9836,N_9847);
or U10055 (N_10055,N_9883,N_9804);
nor U10056 (N_10056,N_9799,N_9821);
nand U10057 (N_10057,N_9862,N_9856);
nand U10058 (N_10058,N_9816,N_9768);
and U10059 (N_10059,N_9796,N_9869);
nand U10060 (N_10060,N_9880,N_9814);
or U10061 (N_10061,N_9880,N_9800);
nand U10062 (N_10062,N_9897,N_9866);
nand U10063 (N_10063,N_9839,N_9850);
and U10064 (N_10064,N_9885,N_9823);
nor U10065 (N_10065,N_9873,N_9806);
nand U10066 (N_10066,N_9824,N_9831);
nor U10067 (N_10067,N_9882,N_9875);
or U10068 (N_10068,N_9913,N_9892);
xor U10069 (N_10069,N_9823,N_9902);
nor U10070 (N_10070,N_9875,N_9818);
nor U10071 (N_10071,N_9916,N_9770);
nand U10072 (N_10072,N_9768,N_9845);
and U10073 (N_10073,N_9886,N_9895);
nand U10074 (N_10074,N_9863,N_9829);
or U10075 (N_10075,N_9894,N_9816);
nor U10076 (N_10076,N_9883,N_9898);
nor U10077 (N_10077,N_9872,N_9824);
nand U10078 (N_10078,N_9809,N_9887);
or U10079 (N_10079,N_9768,N_9774);
or U10080 (N_10080,N_9927,N_10001);
xor U10081 (N_10081,N_9920,N_10048);
and U10082 (N_10082,N_10028,N_10072);
nor U10083 (N_10083,N_9990,N_9979);
xor U10084 (N_10084,N_10035,N_9921);
nand U10085 (N_10085,N_9975,N_10004);
nand U10086 (N_10086,N_9950,N_9951);
nand U10087 (N_10087,N_10046,N_9931);
or U10088 (N_10088,N_9993,N_9992);
or U10089 (N_10089,N_10036,N_9966);
xor U10090 (N_10090,N_10038,N_10008);
xor U10091 (N_10091,N_9922,N_9971);
xor U10092 (N_10092,N_10064,N_10029);
xor U10093 (N_10093,N_9954,N_9976);
and U10094 (N_10094,N_9928,N_9985);
nor U10095 (N_10095,N_9970,N_9941);
nand U10096 (N_10096,N_10059,N_10023);
nand U10097 (N_10097,N_9969,N_10055);
nand U10098 (N_10098,N_10002,N_10044);
and U10099 (N_10099,N_10034,N_10015);
and U10100 (N_10100,N_9960,N_10077);
and U10101 (N_10101,N_10027,N_10071);
or U10102 (N_10102,N_9999,N_9972);
or U10103 (N_10103,N_9989,N_10049);
and U10104 (N_10104,N_10051,N_9946);
and U10105 (N_10105,N_9964,N_9959);
xnor U10106 (N_10106,N_9998,N_10057);
nor U10107 (N_10107,N_9978,N_9952);
and U10108 (N_10108,N_9924,N_9962);
nand U10109 (N_10109,N_9935,N_9937);
and U10110 (N_10110,N_9925,N_9987);
nand U10111 (N_10111,N_10007,N_9949);
nand U10112 (N_10112,N_10032,N_9997);
or U10113 (N_10113,N_9967,N_10022);
or U10114 (N_10114,N_9994,N_9961);
and U10115 (N_10115,N_10079,N_10040);
xor U10116 (N_10116,N_10005,N_10019);
nand U10117 (N_10117,N_10061,N_9932);
and U10118 (N_10118,N_10068,N_10024);
xor U10119 (N_10119,N_9986,N_10073);
xnor U10120 (N_10120,N_9939,N_9926);
or U10121 (N_10121,N_10076,N_9968);
xor U10122 (N_10122,N_10065,N_10050);
nand U10123 (N_10123,N_10006,N_9923);
and U10124 (N_10124,N_9963,N_10012);
xor U10125 (N_10125,N_9995,N_9945);
nor U10126 (N_10126,N_10031,N_10025);
nand U10127 (N_10127,N_10060,N_9956);
and U10128 (N_10128,N_9940,N_9958);
xnor U10129 (N_10129,N_9980,N_9944);
or U10130 (N_10130,N_9977,N_10010);
xnor U10131 (N_10131,N_10003,N_9948);
xor U10132 (N_10132,N_10039,N_10030);
nand U10133 (N_10133,N_10013,N_9988);
xnor U10134 (N_10134,N_10056,N_10000);
nand U10135 (N_10135,N_9953,N_10041);
or U10136 (N_10136,N_9929,N_10014);
and U10137 (N_10137,N_10067,N_10058);
nor U10138 (N_10138,N_10016,N_10033);
or U10139 (N_10139,N_10042,N_9938);
and U10140 (N_10140,N_10037,N_10045);
or U10141 (N_10141,N_9973,N_10021);
or U10142 (N_10142,N_10063,N_9955);
nor U10143 (N_10143,N_10070,N_9996);
and U10144 (N_10144,N_10052,N_10009);
nor U10145 (N_10145,N_10069,N_10053);
or U10146 (N_10146,N_9974,N_10054);
nor U10147 (N_10147,N_9982,N_9934);
or U10148 (N_10148,N_10011,N_10074);
and U10149 (N_10149,N_10075,N_9942);
and U10150 (N_10150,N_9933,N_9936);
and U10151 (N_10151,N_9943,N_10043);
or U10152 (N_10152,N_9947,N_9983);
nor U10153 (N_10153,N_10078,N_9991);
or U10154 (N_10154,N_10026,N_10020);
nand U10155 (N_10155,N_9957,N_9930);
or U10156 (N_10156,N_9981,N_10062);
nor U10157 (N_10157,N_9984,N_10018);
or U10158 (N_10158,N_10017,N_10066);
nor U10159 (N_10159,N_10047,N_9965);
or U10160 (N_10160,N_10021,N_10044);
and U10161 (N_10161,N_10007,N_10070);
xnor U10162 (N_10162,N_9949,N_9997);
xnor U10163 (N_10163,N_10024,N_10032);
xor U10164 (N_10164,N_9972,N_10001);
nand U10165 (N_10165,N_9948,N_9982);
xnor U10166 (N_10166,N_9964,N_10031);
or U10167 (N_10167,N_10054,N_10019);
nand U10168 (N_10168,N_9962,N_10028);
nor U10169 (N_10169,N_10010,N_10065);
nor U10170 (N_10170,N_10027,N_10078);
nor U10171 (N_10171,N_10071,N_10070);
xor U10172 (N_10172,N_10056,N_10015);
or U10173 (N_10173,N_9987,N_9988);
xor U10174 (N_10174,N_10013,N_10044);
nor U10175 (N_10175,N_10049,N_10036);
nand U10176 (N_10176,N_10029,N_9981);
nand U10177 (N_10177,N_10004,N_9970);
or U10178 (N_10178,N_9975,N_9995);
xnor U10179 (N_10179,N_9964,N_9954);
xnor U10180 (N_10180,N_10063,N_10037);
or U10181 (N_10181,N_10077,N_10020);
and U10182 (N_10182,N_9948,N_9994);
or U10183 (N_10183,N_9959,N_10077);
nand U10184 (N_10184,N_10065,N_9976);
xor U10185 (N_10185,N_10069,N_10047);
nand U10186 (N_10186,N_9930,N_10013);
nor U10187 (N_10187,N_9963,N_9986);
nand U10188 (N_10188,N_10069,N_10059);
and U10189 (N_10189,N_10047,N_10024);
xnor U10190 (N_10190,N_10030,N_9978);
xor U10191 (N_10191,N_10027,N_10020);
or U10192 (N_10192,N_10009,N_10066);
nor U10193 (N_10193,N_10078,N_9946);
nand U10194 (N_10194,N_9952,N_9926);
nand U10195 (N_10195,N_10078,N_10044);
xor U10196 (N_10196,N_10001,N_10013);
nand U10197 (N_10197,N_10069,N_10040);
xor U10198 (N_10198,N_9986,N_9926);
and U10199 (N_10199,N_9951,N_9944);
and U10200 (N_10200,N_9967,N_10037);
xnor U10201 (N_10201,N_10028,N_10036);
nor U10202 (N_10202,N_9933,N_9971);
and U10203 (N_10203,N_9922,N_10077);
xor U10204 (N_10204,N_9996,N_9923);
nor U10205 (N_10205,N_10075,N_9925);
nor U10206 (N_10206,N_9932,N_10071);
and U10207 (N_10207,N_10079,N_10025);
or U10208 (N_10208,N_10075,N_10062);
xor U10209 (N_10209,N_10052,N_9956);
xnor U10210 (N_10210,N_9933,N_9980);
or U10211 (N_10211,N_10078,N_10036);
and U10212 (N_10212,N_10035,N_10031);
and U10213 (N_10213,N_10036,N_10040);
or U10214 (N_10214,N_9929,N_9969);
nand U10215 (N_10215,N_10042,N_9983);
nand U10216 (N_10216,N_10040,N_9965);
or U10217 (N_10217,N_9997,N_10034);
nor U10218 (N_10218,N_10061,N_9941);
nand U10219 (N_10219,N_9930,N_9928);
nor U10220 (N_10220,N_10079,N_9979);
or U10221 (N_10221,N_10021,N_10063);
xnor U10222 (N_10222,N_10048,N_9952);
and U10223 (N_10223,N_9993,N_9958);
nor U10224 (N_10224,N_9940,N_10047);
nor U10225 (N_10225,N_9987,N_9972);
and U10226 (N_10226,N_9982,N_9998);
nor U10227 (N_10227,N_9942,N_9953);
nand U10228 (N_10228,N_10073,N_9988);
xor U10229 (N_10229,N_9948,N_10012);
xor U10230 (N_10230,N_10063,N_10028);
nand U10231 (N_10231,N_10028,N_10032);
nand U10232 (N_10232,N_9974,N_10067);
and U10233 (N_10233,N_10026,N_9971);
xor U10234 (N_10234,N_10048,N_9947);
xnor U10235 (N_10235,N_10031,N_10043);
nand U10236 (N_10236,N_9960,N_9946);
and U10237 (N_10237,N_9965,N_9969);
nand U10238 (N_10238,N_9962,N_10054);
nand U10239 (N_10239,N_9956,N_10005);
and U10240 (N_10240,N_10199,N_10089);
nor U10241 (N_10241,N_10119,N_10135);
and U10242 (N_10242,N_10084,N_10188);
nor U10243 (N_10243,N_10136,N_10131);
and U10244 (N_10244,N_10232,N_10215);
and U10245 (N_10245,N_10201,N_10193);
and U10246 (N_10246,N_10151,N_10112);
or U10247 (N_10247,N_10158,N_10192);
nand U10248 (N_10248,N_10127,N_10085);
or U10249 (N_10249,N_10137,N_10210);
or U10250 (N_10250,N_10183,N_10176);
and U10251 (N_10251,N_10107,N_10145);
nor U10252 (N_10252,N_10214,N_10115);
and U10253 (N_10253,N_10080,N_10098);
xor U10254 (N_10254,N_10090,N_10169);
and U10255 (N_10255,N_10223,N_10106);
and U10256 (N_10256,N_10194,N_10110);
and U10257 (N_10257,N_10190,N_10155);
nand U10258 (N_10258,N_10118,N_10224);
and U10259 (N_10259,N_10165,N_10149);
nand U10260 (N_10260,N_10160,N_10126);
xnor U10261 (N_10261,N_10229,N_10086);
nor U10262 (N_10262,N_10175,N_10164);
or U10263 (N_10263,N_10082,N_10206);
nand U10264 (N_10264,N_10227,N_10228);
or U10265 (N_10265,N_10230,N_10200);
xor U10266 (N_10266,N_10134,N_10088);
and U10267 (N_10267,N_10221,N_10182);
xnor U10268 (N_10268,N_10217,N_10195);
and U10269 (N_10269,N_10141,N_10130);
nor U10270 (N_10270,N_10102,N_10148);
nand U10271 (N_10271,N_10108,N_10197);
and U10272 (N_10272,N_10180,N_10226);
or U10273 (N_10273,N_10125,N_10124);
and U10274 (N_10274,N_10101,N_10144);
xor U10275 (N_10275,N_10219,N_10128);
or U10276 (N_10276,N_10189,N_10212);
and U10277 (N_10277,N_10139,N_10205);
nand U10278 (N_10278,N_10095,N_10233);
nor U10279 (N_10279,N_10161,N_10093);
nor U10280 (N_10280,N_10147,N_10167);
xnor U10281 (N_10281,N_10116,N_10109);
or U10282 (N_10282,N_10187,N_10092);
nand U10283 (N_10283,N_10186,N_10097);
xor U10284 (N_10284,N_10216,N_10174);
nand U10285 (N_10285,N_10154,N_10171);
and U10286 (N_10286,N_10168,N_10191);
nand U10287 (N_10287,N_10142,N_10178);
nor U10288 (N_10288,N_10091,N_10150);
xnor U10289 (N_10289,N_10202,N_10099);
nand U10290 (N_10290,N_10105,N_10133);
and U10291 (N_10291,N_10179,N_10143);
nand U10292 (N_10292,N_10113,N_10218);
nor U10293 (N_10293,N_10083,N_10157);
xnor U10294 (N_10294,N_10121,N_10170);
nor U10295 (N_10295,N_10159,N_10172);
nand U10296 (N_10296,N_10184,N_10103);
and U10297 (N_10297,N_10122,N_10185);
nand U10298 (N_10298,N_10239,N_10203);
and U10299 (N_10299,N_10163,N_10213);
and U10300 (N_10300,N_10177,N_10204);
xor U10301 (N_10301,N_10104,N_10081);
or U10302 (N_10302,N_10123,N_10231);
xnor U10303 (N_10303,N_10153,N_10140);
nand U10304 (N_10304,N_10209,N_10132);
and U10305 (N_10305,N_10096,N_10225);
xor U10306 (N_10306,N_10235,N_10129);
xor U10307 (N_10307,N_10207,N_10146);
nor U10308 (N_10308,N_10211,N_10111);
xor U10309 (N_10309,N_10196,N_10120);
nor U10310 (N_10310,N_10156,N_10138);
nor U10311 (N_10311,N_10220,N_10087);
xnor U10312 (N_10312,N_10238,N_10222);
or U10313 (N_10313,N_10198,N_10236);
or U10314 (N_10314,N_10152,N_10117);
nand U10315 (N_10315,N_10181,N_10208);
nand U10316 (N_10316,N_10094,N_10166);
nor U10317 (N_10317,N_10162,N_10100);
xor U10318 (N_10318,N_10114,N_10237);
nor U10319 (N_10319,N_10173,N_10234);
and U10320 (N_10320,N_10203,N_10237);
or U10321 (N_10321,N_10239,N_10101);
nor U10322 (N_10322,N_10106,N_10220);
and U10323 (N_10323,N_10134,N_10218);
nand U10324 (N_10324,N_10131,N_10155);
nand U10325 (N_10325,N_10146,N_10192);
nor U10326 (N_10326,N_10133,N_10214);
xnor U10327 (N_10327,N_10200,N_10138);
nand U10328 (N_10328,N_10192,N_10137);
nand U10329 (N_10329,N_10194,N_10208);
and U10330 (N_10330,N_10109,N_10230);
xnor U10331 (N_10331,N_10104,N_10189);
xor U10332 (N_10332,N_10159,N_10160);
or U10333 (N_10333,N_10225,N_10159);
or U10334 (N_10334,N_10169,N_10173);
or U10335 (N_10335,N_10186,N_10182);
xnor U10336 (N_10336,N_10231,N_10132);
xnor U10337 (N_10337,N_10203,N_10094);
or U10338 (N_10338,N_10219,N_10110);
xor U10339 (N_10339,N_10133,N_10210);
nor U10340 (N_10340,N_10199,N_10194);
and U10341 (N_10341,N_10137,N_10207);
nor U10342 (N_10342,N_10229,N_10218);
nor U10343 (N_10343,N_10096,N_10150);
nor U10344 (N_10344,N_10224,N_10128);
nand U10345 (N_10345,N_10217,N_10228);
nand U10346 (N_10346,N_10200,N_10214);
or U10347 (N_10347,N_10191,N_10233);
or U10348 (N_10348,N_10185,N_10179);
or U10349 (N_10349,N_10196,N_10139);
xnor U10350 (N_10350,N_10147,N_10196);
or U10351 (N_10351,N_10192,N_10186);
and U10352 (N_10352,N_10096,N_10083);
nand U10353 (N_10353,N_10133,N_10230);
xnor U10354 (N_10354,N_10176,N_10231);
or U10355 (N_10355,N_10180,N_10135);
or U10356 (N_10356,N_10191,N_10105);
xnor U10357 (N_10357,N_10162,N_10093);
and U10358 (N_10358,N_10166,N_10181);
xnor U10359 (N_10359,N_10128,N_10153);
nor U10360 (N_10360,N_10122,N_10192);
nand U10361 (N_10361,N_10131,N_10220);
and U10362 (N_10362,N_10086,N_10181);
nor U10363 (N_10363,N_10190,N_10159);
or U10364 (N_10364,N_10217,N_10202);
nor U10365 (N_10365,N_10201,N_10121);
or U10366 (N_10366,N_10148,N_10229);
nand U10367 (N_10367,N_10212,N_10166);
or U10368 (N_10368,N_10094,N_10119);
nand U10369 (N_10369,N_10209,N_10197);
xor U10370 (N_10370,N_10091,N_10126);
and U10371 (N_10371,N_10129,N_10171);
or U10372 (N_10372,N_10136,N_10162);
nor U10373 (N_10373,N_10196,N_10159);
xor U10374 (N_10374,N_10176,N_10147);
nand U10375 (N_10375,N_10095,N_10156);
xor U10376 (N_10376,N_10187,N_10206);
nand U10377 (N_10377,N_10226,N_10124);
and U10378 (N_10378,N_10136,N_10174);
nor U10379 (N_10379,N_10087,N_10123);
or U10380 (N_10380,N_10098,N_10142);
or U10381 (N_10381,N_10181,N_10129);
or U10382 (N_10382,N_10218,N_10199);
and U10383 (N_10383,N_10144,N_10103);
or U10384 (N_10384,N_10098,N_10235);
nand U10385 (N_10385,N_10111,N_10164);
or U10386 (N_10386,N_10112,N_10087);
nor U10387 (N_10387,N_10142,N_10118);
nand U10388 (N_10388,N_10155,N_10219);
xnor U10389 (N_10389,N_10205,N_10089);
nor U10390 (N_10390,N_10201,N_10188);
xnor U10391 (N_10391,N_10111,N_10081);
xor U10392 (N_10392,N_10154,N_10116);
nand U10393 (N_10393,N_10187,N_10083);
nor U10394 (N_10394,N_10192,N_10147);
nand U10395 (N_10395,N_10231,N_10236);
nand U10396 (N_10396,N_10176,N_10154);
nand U10397 (N_10397,N_10091,N_10177);
or U10398 (N_10398,N_10139,N_10127);
nand U10399 (N_10399,N_10189,N_10207);
or U10400 (N_10400,N_10332,N_10308);
nand U10401 (N_10401,N_10300,N_10281);
nand U10402 (N_10402,N_10262,N_10317);
nor U10403 (N_10403,N_10241,N_10278);
xnor U10404 (N_10404,N_10390,N_10258);
xor U10405 (N_10405,N_10394,N_10369);
nand U10406 (N_10406,N_10357,N_10259);
or U10407 (N_10407,N_10368,N_10244);
and U10408 (N_10408,N_10253,N_10383);
nor U10409 (N_10409,N_10337,N_10265);
or U10410 (N_10410,N_10256,N_10292);
nand U10411 (N_10411,N_10354,N_10306);
xor U10412 (N_10412,N_10377,N_10257);
nor U10413 (N_10413,N_10371,N_10260);
and U10414 (N_10414,N_10284,N_10378);
and U10415 (N_10415,N_10330,N_10269);
and U10416 (N_10416,N_10388,N_10318);
nor U10417 (N_10417,N_10326,N_10352);
and U10418 (N_10418,N_10261,N_10341);
nand U10419 (N_10419,N_10267,N_10327);
nor U10420 (N_10420,N_10315,N_10302);
or U10421 (N_10421,N_10283,N_10333);
or U10422 (N_10422,N_10339,N_10307);
nor U10423 (N_10423,N_10243,N_10392);
or U10424 (N_10424,N_10366,N_10347);
nand U10425 (N_10425,N_10344,N_10310);
nand U10426 (N_10426,N_10381,N_10293);
nor U10427 (N_10427,N_10255,N_10364);
or U10428 (N_10428,N_10282,N_10309);
nor U10429 (N_10429,N_10277,N_10248);
nand U10430 (N_10430,N_10303,N_10320);
xnor U10431 (N_10431,N_10270,N_10304);
nand U10432 (N_10432,N_10274,N_10275);
or U10433 (N_10433,N_10245,N_10386);
nor U10434 (N_10434,N_10335,N_10319);
nor U10435 (N_10435,N_10398,N_10296);
and U10436 (N_10436,N_10328,N_10289);
or U10437 (N_10437,N_10374,N_10387);
nor U10438 (N_10438,N_10365,N_10246);
nor U10439 (N_10439,N_10349,N_10373);
xor U10440 (N_10440,N_10251,N_10323);
or U10441 (N_10441,N_10351,N_10345);
or U10442 (N_10442,N_10362,N_10252);
or U10443 (N_10443,N_10359,N_10297);
xnor U10444 (N_10444,N_10372,N_10264);
nor U10445 (N_10445,N_10240,N_10271);
nand U10446 (N_10446,N_10272,N_10280);
and U10447 (N_10447,N_10290,N_10375);
nand U10448 (N_10448,N_10384,N_10342);
and U10449 (N_10449,N_10355,N_10343);
or U10450 (N_10450,N_10393,N_10363);
xnor U10451 (N_10451,N_10370,N_10353);
and U10452 (N_10452,N_10321,N_10395);
nand U10453 (N_10453,N_10360,N_10379);
nor U10454 (N_10454,N_10322,N_10348);
xor U10455 (N_10455,N_10350,N_10356);
xnor U10456 (N_10456,N_10334,N_10268);
and U10457 (N_10457,N_10346,N_10399);
xnor U10458 (N_10458,N_10305,N_10263);
nand U10459 (N_10459,N_10358,N_10336);
nor U10460 (N_10460,N_10329,N_10331);
xor U10461 (N_10461,N_10279,N_10382);
nand U10462 (N_10462,N_10295,N_10276);
nor U10463 (N_10463,N_10249,N_10298);
xor U10464 (N_10464,N_10250,N_10242);
or U10465 (N_10465,N_10294,N_10247);
and U10466 (N_10466,N_10312,N_10285);
nor U10467 (N_10467,N_10288,N_10391);
or U10468 (N_10468,N_10273,N_10299);
and U10469 (N_10469,N_10311,N_10316);
nand U10470 (N_10470,N_10286,N_10314);
or U10471 (N_10471,N_10396,N_10266);
nand U10472 (N_10472,N_10376,N_10301);
or U10473 (N_10473,N_10380,N_10313);
and U10474 (N_10474,N_10367,N_10287);
nand U10475 (N_10475,N_10389,N_10291);
xnor U10476 (N_10476,N_10361,N_10324);
nand U10477 (N_10477,N_10385,N_10338);
and U10478 (N_10478,N_10340,N_10397);
nor U10479 (N_10479,N_10325,N_10254);
xor U10480 (N_10480,N_10321,N_10293);
or U10481 (N_10481,N_10258,N_10364);
nand U10482 (N_10482,N_10368,N_10385);
nand U10483 (N_10483,N_10333,N_10397);
xnor U10484 (N_10484,N_10268,N_10274);
xor U10485 (N_10485,N_10376,N_10261);
or U10486 (N_10486,N_10375,N_10258);
nand U10487 (N_10487,N_10327,N_10274);
xnor U10488 (N_10488,N_10268,N_10254);
or U10489 (N_10489,N_10387,N_10271);
xnor U10490 (N_10490,N_10296,N_10312);
or U10491 (N_10491,N_10248,N_10361);
and U10492 (N_10492,N_10344,N_10307);
or U10493 (N_10493,N_10326,N_10284);
or U10494 (N_10494,N_10355,N_10258);
nor U10495 (N_10495,N_10379,N_10292);
xor U10496 (N_10496,N_10353,N_10287);
or U10497 (N_10497,N_10391,N_10267);
nand U10498 (N_10498,N_10256,N_10272);
and U10499 (N_10499,N_10251,N_10304);
and U10500 (N_10500,N_10354,N_10298);
nor U10501 (N_10501,N_10348,N_10331);
or U10502 (N_10502,N_10356,N_10255);
or U10503 (N_10503,N_10268,N_10342);
nor U10504 (N_10504,N_10286,N_10254);
or U10505 (N_10505,N_10261,N_10295);
nor U10506 (N_10506,N_10346,N_10283);
nor U10507 (N_10507,N_10312,N_10326);
nor U10508 (N_10508,N_10253,N_10275);
and U10509 (N_10509,N_10274,N_10336);
nand U10510 (N_10510,N_10242,N_10359);
xor U10511 (N_10511,N_10279,N_10352);
or U10512 (N_10512,N_10300,N_10380);
nand U10513 (N_10513,N_10266,N_10309);
xor U10514 (N_10514,N_10335,N_10343);
nor U10515 (N_10515,N_10330,N_10293);
nand U10516 (N_10516,N_10285,N_10324);
xor U10517 (N_10517,N_10247,N_10252);
nand U10518 (N_10518,N_10321,N_10386);
or U10519 (N_10519,N_10273,N_10377);
nor U10520 (N_10520,N_10351,N_10385);
xnor U10521 (N_10521,N_10289,N_10357);
or U10522 (N_10522,N_10381,N_10243);
xnor U10523 (N_10523,N_10386,N_10360);
or U10524 (N_10524,N_10375,N_10275);
xnor U10525 (N_10525,N_10246,N_10278);
and U10526 (N_10526,N_10341,N_10355);
and U10527 (N_10527,N_10290,N_10356);
or U10528 (N_10528,N_10348,N_10376);
nand U10529 (N_10529,N_10326,N_10397);
and U10530 (N_10530,N_10315,N_10372);
xor U10531 (N_10531,N_10291,N_10318);
nor U10532 (N_10532,N_10245,N_10350);
xnor U10533 (N_10533,N_10378,N_10254);
nand U10534 (N_10534,N_10370,N_10331);
and U10535 (N_10535,N_10328,N_10302);
and U10536 (N_10536,N_10341,N_10350);
or U10537 (N_10537,N_10260,N_10339);
and U10538 (N_10538,N_10268,N_10348);
nand U10539 (N_10539,N_10319,N_10379);
xnor U10540 (N_10540,N_10300,N_10394);
nor U10541 (N_10541,N_10294,N_10252);
and U10542 (N_10542,N_10330,N_10345);
nand U10543 (N_10543,N_10369,N_10345);
nor U10544 (N_10544,N_10317,N_10335);
and U10545 (N_10545,N_10286,N_10338);
xnor U10546 (N_10546,N_10283,N_10396);
nand U10547 (N_10547,N_10284,N_10398);
or U10548 (N_10548,N_10259,N_10278);
nor U10549 (N_10549,N_10346,N_10280);
nand U10550 (N_10550,N_10315,N_10333);
nand U10551 (N_10551,N_10292,N_10357);
nor U10552 (N_10552,N_10336,N_10327);
nand U10553 (N_10553,N_10280,N_10375);
and U10554 (N_10554,N_10341,N_10366);
nor U10555 (N_10555,N_10306,N_10258);
or U10556 (N_10556,N_10379,N_10397);
nor U10557 (N_10557,N_10331,N_10336);
or U10558 (N_10558,N_10287,N_10288);
nand U10559 (N_10559,N_10262,N_10250);
and U10560 (N_10560,N_10498,N_10454);
or U10561 (N_10561,N_10502,N_10419);
and U10562 (N_10562,N_10558,N_10485);
and U10563 (N_10563,N_10553,N_10457);
and U10564 (N_10564,N_10471,N_10480);
xnor U10565 (N_10565,N_10543,N_10533);
nand U10566 (N_10566,N_10479,N_10446);
nor U10567 (N_10567,N_10510,N_10519);
nor U10568 (N_10568,N_10492,N_10433);
nand U10569 (N_10569,N_10469,N_10504);
xnor U10570 (N_10570,N_10464,N_10437);
nand U10571 (N_10571,N_10451,N_10501);
nand U10572 (N_10572,N_10465,N_10414);
nor U10573 (N_10573,N_10466,N_10551);
or U10574 (N_10574,N_10412,N_10431);
xor U10575 (N_10575,N_10539,N_10439);
xnor U10576 (N_10576,N_10441,N_10531);
nand U10577 (N_10577,N_10449,N_10517);
or U10578 (N_10578,N_10518,N_10421);
and U10579 (N_10579,N_10483,N_10452);
and U10580 (N_10580,N_10536,N_10408);
or U10581 (N_10581,N_10534,N_10470);
xnor U10582 (N_10582,N_10538,N_10512);
nand U10583 (N_10583,N_10448,N_10508);
and U10584 (N_10584,N_10425,N_10490);
nand U10585 (N_10585,N_10499,N_10511);
nand U10586 (N_10586,N_10491,N_10557);
xor U10587 (N_10587,N_10467,N_10436);
xnor U10588 (N_10588,N_10528,N_10420);
or U10589 (N_10589,N_10521,N_10404);
xor U10590 (N_10590,N_10423,N_10405);
nand U10591 (N_10591,N_10406,N_10427);
xor U10592 (N_10592,N_10442,N_10520);
xnor U10593 (N_10593,N_10489,N_10545);
nand U10594 (N_10594,N_10507,N_10494);
nand U10595 (N_10595,N_10424,N_10463);
or U10596 (N_10596,N_10552,N_10440);
nand U10597 (N_10597,N_10546,N_10447);
nor U10598 (N_10598,N_10453,N_10478);
xor U10599 (N_10599,N_10411,N_10555);
or U10600 (N_10600,N_10473,N_10559);
or U10601 (N_10601,N_10401,N_10455);
nor U10602 (N_10602,N_10526,N_10450);
nand U10603 (N_10603,N_10477,N_10487);
xor U10604 (N_10604,N_10549,N_10472);
xor U10605 (N_10605,N_10410,N_10488);
nand U10606 (N_10606,N_10429,N_10444);
nor U10607 (N_10607,N_10428,N_10461);
or U10608 (N_10608,N_10475,N_10443);
nor U10609 (N_10609,N_10497,N_10418);
and U10610 (N_10610,N_10547,N_10407);
xnor U10611 (N_10611,N_10481,N_10415);
and U10612 (N_10612,N_10459,N_10482);
nor U10613 (N_10613,N_10493,N_10513);
xnor U10614 (N_10614,N_10525,N_10400);
nor U10615 (N_10615,N_10435,N_10484);
and U10616 (N_10616,N_10514,N_10474);
or U10617 (N_10617,N_10542,N_10527);
or U10618 (N_10618,N_10432,N_10403);
and U10619 (N_10619,N_10548,N_10458);
xnor U10620 (N_10620,N_10416,N_10495);
nor U10621 (N_10621,N_10529,N_10506);
and U10622 (N_10622,N_10530,N_10522);
nand U10623 (N_10623,N_10426,N_10541);
nand U10624 (N_10624,N_10413,N_10500);
nand U10625 (N_10625,N_10544,N_10476);
nand U10626 (N_10626,N_10554,N_10417);
nand U10627 (N_10627,N_10422,N_10516);
nor U10628 (N_10628,N_10468,N_10535);
xnor U10629 (N_10629,N_10456,N_10438);
nor U10630 (N_10630,N_10409,N_10402);
xnor U10631 (N_10631,N_10540,N_10503);
or U10632 (N_10632,N_10515,N_10460);
nor U10633 (N_10633,N_10523,N_10486);
or U10634 (N_10634,N_10430,N_10524);
nand U10635 (N_10635,N_10509,N_10550);
nand U10636 (N_10636,N_10496,N_10537);
xnor U10637 (N_10637,N_10556,N_10445);
xnor U10638 (N_10638,N_10434,N_10505);
nor U10639 (N_10639,N_10532,N_10462);
xor U10640 (N_10640,N_10420,N_10478);
nor U10641 (N_10641,N_10463,N_10499);
and U10642 (N_10642,N_10440,N_10476);
or U10643 (N_10643,N_10412,N_10451);
nor U10644 (N_10644,N_10486,N_10485);
nand U10645 (N_10645,N_10471,N_10521);
or U10646 (N_10646,N_10548,N_10525);
nor U10647 (N_10647,N_10441,N_10548);
or U10648 (N_10648,N_10431,N_10409);
nor U10649 (N_10649,N_10482,N_10464);
nor U10650 (N_10650,N_10522,N_10424);
and U10651 (N_10651,N_10411,N_10515);
or U10652 (N_10652,N_10521,N_10530);
or U10653 (N_10653,N_10484,N_10478);
xnor U10654 (N_10654,N_10517,N_10444);
xor U10655 (N_10655,N_10543,N_10536);
or U10656 (N_10656,N_10500,N_10513);
or U10657 (N_10657,N_10406,N_10522);
nor U10658 (N_10658,N_10457,N_10410);
nand U10659 (N_10659,N_10451,N_10510);
nand U10660 (N_10660,N_10505,N_10547);
or U10661 (N_10661,N_10547,N_10538);
or U10662 (N_10662,N_10553,N_10423);
or U10663 (N_10663,N_10500,N_10471);
or U10664 (N_10664,N_10523,N_10476);
xnor U10665 (N_10665,N_10487,N_10514);
and U10666 (N_10666,N_10520,N_10448);
nor U10667 (N_10667,N_10454,N_10472);
and U10668 (N_10668,N_10497,N_10489);
nor U10669 (N_10669,N_10547,N_10457);
nor U10670 (N_10670,N_10507,N_10496);
xnor U10671 (N_10671,N_10502,N_10518);
nand U10672 (N_10672,N_10412,N_10407);
and U10673 (N_10673,N_10480,N_10427);
or U10674 (N_10674,N_10429,N_10465);
nand U10675 (N_10675,N_10556,N_10524);
or U10676 (N_10676,N_10488,N_10490);
nor U10677 (N_10677,N_10442,N_10559);
and U10678 (N_10678,N_10446,N_10499);
nor U10679 (N_10679,N_10405,N_10510);
nor U10680 (N_10680,N_10499,N_10410);
or U10681 (N_10681,N_10479,N_10478);
nand U10682 (N_10682,N_10546,N_10423);
nand U10683 (N_10683,N_10525,N_10552);
and U10684 (N_10684,N_10423,N_10489);
xnor U10685 (N_10685,N_10546,N_10485);
nand U10686 (N_10686,N_10472,N_10428);
xnor U10687 (N_10687,N_10558,N_10513);
xnor U10688 (N_10688,N_10500,N_10426);
and U10689 (N_10689,N_10483,N_10523);
and U10690 (N_10690,N_10511,N_10506);
nor U10691 (N_10691,N_10502,N_10472);
nor U10692 (N_10692,N_10550,N_10546);
or U10693 (N_10693,N_10509,N_10516);
nor U10694 (N_10694,N_10545,N_10516);
nor U10695 (N_10695,N_10556,N_10474);
and U10696 (N_10696,N_10447,N_10404);
nand U10697 (N_10697,N_10477,N_10506);
nor U10698 (N_10698,N_10521,N_10483);
and U10699 (N_10699,N_10403,N_10525);
nor U10700 (N_10700,N_10437,N_10541);
and U10701 (N_10701,N_10514,N_10466);
nor U10702 (N_10702,N_10489,N_10407);
xnor U10703 (N_10703,N_10445,N_10470);
and U10704 (N_10704,N_10538,N_10557);
and U10705 (N_10705,N_10471,N_10498);
or U10706 (N_10706,N_10452,N_10444);
xor U10707 (N_10707,N_10463,N_10404);
nand U10708 (N_10708,N_10549,N_10558);
and U10709 (N_10709,N_10522,N_10450);
nand U10710 (N_10710,N_10541,N_10506);
and U10711 (N_10711,N_10516,N_10470);
or U10712 (N_10712,N_10497,N_10425);
nand U10713 (N_10713,N_10559,N_10467);
xnor U10714 (N_10714,N_10488,N_10528);
nand U10715 (N_10715,N_10400,N_10402);
xor U10716 (N_10716,N_10521,N_10458);
and U10717 (N_10717,N_10508,N_10421);
nor U10718 (N_10718,N_10433,N_10556);
xnor U10719 (N_10719,N_10556,N_10483);
nand U10720 (N_10720,N_10709,N_10583);
or U10721 (N_10721,N_10665,N_10572);
nand U10722 (N_10722,N_10632,N_10687);
xor U10723 (N_10723,N_10619,N_10618);
xor U10724 (N_10724,N_10664,N_10561);
or U10725 (N_10725,N_10634,N_10574);
nand U10726 (N_10726,N_10564,N_10568);
xnor U10727 (N_10727,N_10717,N_10601);
xor U10728 (N_10728,N_10600,N_10567);
and U10729 (N_10729,N_10651,N_10595);
or U10730 (N_10730,N_10616,N_10690);
nor U10731 (N_10731,N_10688,N_10625);
nor U10732 (N_10732,N_10683,N_10656);
nand U10733 (N_10733,N_10654,N_10629);
and U10734 (N_10734,N_10640,N_10686);
nand U10735 (N_10735,N_10606,N_10694);
and U10736 (N_10736,N_10679,N_10695);
and U10737 (N_10737,N_10716,N_10628);
nor U10738 (N_10738,N_10672,N_10660);
or U10739 (N_10739,N_10612,N_10699);
nand U10740 (N_10740,N_10597,N_10698);
nand U10741 (N_10741,N_10650,N_10702);
and U10742 (N_10742,N_10594,N_10569);
xor U10743 (N_10743,N_10577,N_10638);
xor U10744 (N_10744,N_10701,N_10696);
or U10745 (N_10745,N_10667,N_10676);
nand U10746 (N_10746,N_10666,N_10570);
or U10747 (N_10747,N_10635,N_10605);
nor U10748 (N_10748,N_10566,N_10621);
nand U10749 (N_10749,N_10693,N_10593);
and U10750 (N_10750,N_10704,N_10707);
xnor U10751 (N_10751,N_10607,N_10675);
and U10752 (N_10752,N_10586,N_10692);
nand U10753 (N_10753,N_10718,N_10579);
xnor U10754 (N_10754,N_10587,N_10663);
xnor U10755 (N_10755,N_10604,N_10715);
nor U10756 (N_10756,N_10691,N_10642);
nor U10757 (N_10757,N_10598,N_10649);
nand U10758 (N_10758,N_10706,N_10661);
or U10759 (N_10759,N_10578,N_10596);
nand U10760 (N_10760,N_10637,N_10653);
xnor U10761 (N_10761,N_10573,N_10631);
nand U10762 (N_10762,N_10622,N_10617);
nor U10763 (N_10763,N_10677,N_10668);
nand U10764 (N_10764,N_10627,N_10655);
and U10765 (N_10765,N_10719,N_10610);
nor U10766 (N_10766,N_10592,N_10647);
nor U10767 (N_10767,N_10571,N_10697);
or U10768 (N_10768,N_10575,N_10611);
nand U10769 (N_10769,N_10590,N_10711);
xnor U10770 (N_10770,N_10685,N_10560);
nand U10771 (N_10771,N_10581,N_10636);
nor U10772 (N_10772,N_10585,N_10576);
nand U10773 (N_10773,N_10714,N_10609);
nand U10774 (N_10774,N_10680,N_10710);
xor U10775 (N_10775,N_10670,N_10620);
and U10776 (N_10776,N_10602,N_10563);
and U10777 (N_10777,N_10580,N_10626);
nor U10778 (N_10778,N_10682,N_10582);
or U10779 (N_10779,N_10633,N_10659);
or U10780 (N_10780,N_10703,N_10684);
or U10781 (N_10781,N_10652,N_10623);
and U10782 (N_10782,N_10562,N_10678);
nor U10783 (N_10783,N_10671,N_10641);
xnor U10784 (N_10784,N_10657,N_10624);
or U10785 (N_10785,N_10681,N_10643);
nand U10786 (N_10786,N_10591,N_10708);
or U10787 (N_10787,N_10630,N_10648);
or U10788 (N_10788,N_10674,N_10658);
and U10789 (N_10789,N_10603,N_10700);
or U10790 (N_10790,N_10589,N_10662);
or U10791 (N_10791,N_10689,N_10645);
nand U10792 (N_10792,N_10614,N_10588);
nand U10793 (N_10793,N_10613,N_10705);
nor U10794 (N_10794,N_10713,N_10646);
nor U10795 (N_10795,N_10615,N_10584);
xor U10796 (N_10796,N_10639,N_10712);
or U10797 (N_10797,N_10608,N_10599);
xor U10798 (N_10798,N_10669,N_10565);
nor U10799 (N_10799,N_10644,N_10673);
xnor U10800 (N_10800,N_10702,N_10634);
or U10801 (N_10801,N_10679,N_10590);
or U10802 (N_10802,N_10656,N_10568);
xor U10803 (N_10803,N_10680,N_10622);
nor U10804 (N_10804,N_10610,N_10693);
xor U10805 (N_10805,N_10669,N_10716);
nand U10806 (N_10806,N_10641,N_10669);
nor U10807 (N_10807,N_10599,N_10659);
or U10808 (N_10808,N_10682,N_10684);
nand U10809 (N_10809,N_10613,N_10586);
xor U10810 (N_10810,N_10664,N_10629);
or U10811 (N_10811,N_10693,N_10704);
nor U10812 (N_10812,N_10679,N_10606);
xor U10813 (N_10813,N_10650,N_10566);
nor U10814 (N_10814,N_10625,N_10684);
nand U10815 (N_10815,N_10708,N_10581);
nor U10816 (N_10816,N_10564,N_10687);
or U10817 (N_10817,N_10698,N_10626);
and U10818 (N_10818,N_10699,N_10653);
xor U10819 (N_10819,N_10579,N_10569);
or U10820 (N_10820,N_10583,N_10579);
or U10821 (N_10821,N_10570,N_10636);
nand U10822 (N_10822,N_10569,N_10641);
or U10823 (N_10823,N_10610,N_10714);
and U10824 (N_10824,N_10581,N_10619);
or U10825 (N_10825,N_10617,N_10653);
or U10826 (N_10826,N_10586,N_10622);
and U10827 (N_10827,N_10593,N_10607);
or U10828 (N_10828,N_10613,N_10711);
and U10829 (N_10829,N_10600,N_10597);
nand U10830 (N_10830,N_10600,N_10662);
or U10831 (N_10831,N_10694,N_10684);
or U10832 (N_10832,N_10603,N_10605);
nand U10833 (N_10833,N_10638,N_10640);
nand U10834 (N_10834,N_10699,N_10661);
nand U10835 (N_10835,N_10710,N_10592);
and U10836 (N_10836,N_10588,N_10580);
nand U10837 (N_10837,N_10623,N_10583);
nand U10838 (N_10838,N_10696,N_10643);
nand U10839 (N_10839,N_10675,N_10630);
nand U10840 (N_10840,N_10642,N_10659);
xnor U10841 (N_10841,N_10601,N_10645);
xor U10842 (N_10842,N_10618,N_10654);
or U10843 (N_10843,N_10625,N_10676);
nor U10844 (N_10844,N_10671,N_10638);
xor U10845 (N_10845,N_10713,N_10593);
nand U10846 (N_10846,N_10615,N_10636);
nand U10847 (N_10847,N_10694,N_10633);
nor U10848 (N_10848,N_10600,N_10685);
nor U10849 (N_10849,N_10574,N_10593);
nor U10850 (N_10850,N_10655,N_10577);
nand U10851 (N_10851,N_10655,N_10601);
or U10852 (N_10852,N_10664,N_10693);
nand U10853 (N_10853,N_10697,N_10708);
xor U10854 (N_10854,N_10672,N_10575);
or U10855 (N_10855,N_10610,N_10709);
and U10856 (N_10856,N_10686,N_10716);
nor U10857 (N_10857,N_10661,N_10605);
or U10858 (N_10858,N_10616,N_10699);
nand U10859 (N_10859,N_10646,N_10650);
xor U10860 (N_10860,N_10574,N_10592);
nor U10861 (N_10861,N_10635,N_10626);
or U10862 (N_10862,N_10659,N_10574);
nand U10863 (N_10863,N_10700,N_10630);
or U10864 (N_10864,N_10629,N_10607);
xnor U10865 (N_10865,N_10665,N_10692);
nand U10866 (N_10866,N_10713,N_10589);
xor U10867 (N_10867,N_10685,N_10579);
xor U10868 (N_10868,N_10635,N_10687);
xor U10869 (N_10869,N_10576,N_10579);
or U10870 (N_10870,N_10719,N_10659);
nor U10871 (N_10871,N_10645,N_10594);
or U10872 (N_10872,N_10719,N_10714);
xor U10873 (N_10873,N_10624,N_10584);
or U10874 (N_10874,N_10582,N_10627);
and U10875 (N_10875,N_10610,N_10618);
xnor U10876 (N_10876,N_10583,N_10666);
or U10877 (N_10877,N_10563,N_10645);
nor U10878 (N_10878,N_10622,N_10640);
or U10879 (N_10879,N_10625,N_10600);
nand U10880 (N_10880,N_10861,N_10759);
and U10881 (N_10881,N_10870,N_10821);
nor U10882 (N_10882,N_10858,N_10752);
or U10883 (N_10883,N_10864,N_10806);
xor U10884 (N_10884,N_10804,N_10868);
nand U10885 (N_10885,N_10787,N_10818);
xnor U10886 (N_10886,N_10731,N_10740);
and U10887 (N_10887,N_10746,N_10734);
nand U10888 (N_10888,N_10828,N_10801);
or U10889 (N_10889,N_10748,N_10741);
xnor U10890 (N_10890,N_10812,N_10807);
and U10891 (N_10891,N_10797,N_10765);
xor U10892 (N_10892,N_10859,N_10729);
and U10893 (N_10893,N_10875,N_10863);
and U10894 (N_10894,N_10814,N_10779);
or U10895 (N_10895,N_10776,N_10832);
or U10896 (N_10896,N_10736,N_10774);
nor U10897 (N_10897,N_10869,N_10795);
xnor U10898 (N_10898,N_10728,N_10830);
or U10899 (N_10899,N_10811,N_10761);
xnor U10900 (N_10900,N_10844,N_10788);
nor U10901 (N_10901,N_10846,N_10874);
nand U10902 (N_10902,N_10809,N_10792);
nand U10903 (N_10903,N_10857,N_10835);
nand U10904 (N_10904,N_10841,N_10791);
nand U10905 (N_10905,N_10839,N_10726);
xnor U10906 (N_10906,N_10725,N_10815);
and U10907 (N_10907,N_10860,N_10800);
nand U10908 (N_10908,N_10782,N_10866);
xnor U10909 (N_10909,N_10789,N_10850);
nor U10910 (N_10910,N_10724,N_10876);
xnor U10911 (N_10911,N_10786,N_10849);
and U10912 (N_10912,N_10780,N_10784);
or U10913 (N_10913,N_10769,N_10754);
and U10914 (N_10914,N_10878,N_10827);
or U10915 (N_10915,N_10744,N_10767);
and U10916 (N_10916,N_10723,N_10772);
xor U10917 (N_10917,N_10735,N_10873);
xnor U10918 (N_10918,N_10764,N_10785);
xnor U10919 (N_10919,N_10848,N_10824);
nand U10920 (N_10920,N_10766,N_10753);
and U10921 (N_10921,N_10773,N_10837);
and U10922 (N_10922,N_10853,N_10798);
nor U10923 (N_10923,N_10838,N_10799);
and U10924 (N_10924,N_10803,N_10879);
nor U10925 (N_10925,N_10721,N_10756);
xor U10926 (N_10926,N_10867,N_10822);
and U10927 (N_10927,N_10790,N_10840);
or U10928 (N_10928,N_10727,N_10856);
xor U10929 (N_10929,N_10777,N_10862);
and U10930 (N_10930,N_10749,N_10820);
xor U10931 (N_10931,N_10750,N_10722);
nor U10932 (N_10932,N_10833,N_10851);
nor U10933 (N_10933,N_10732,N_10738);
and U10934 (N_10934,N_10743,N_10778);
nor U10935 (N_10935,N_10737,N_10826);
xor U10936 (N_10936,N_10808,N_10842);
and U10937 (N_10937,N_10745,N_10810);
and U10938 (N_10938,N_10834,N_10775);
nor U10939 (N_10939,N_10771,N_10854);
nor U10940 (N_10940,N_10758,N_10831);
nand U10941 (N_10941,N_10872,N_10847);
xnor U10942 (N_10942,N_10730,N_10813);
xor U10943 (N_10943,N_10836,N_10768);
xor U10944 (N_10944,N_10855,N_10783);
and U10945 (N_10945,N_10877,N_10762);
or U10946 (N_10946,N_10793,N_10825);
xnor U10947 (N_10947,N_10733,N_10760);
nand U10948 (N_10948,N_10829,N_10802);
and U10949 (N_10949,N_10751,N_10757);
nor U10950 (N_10950,N_10805,N_10742);
or U10951 (N_10951,N_10770,N_10843);
and U10952 (N_10952,N_10794,N_10819);
nand U10953 (N_10953,N_10845,N_10739);
nor U10954 (N_10954,N_10720,N_10816);
xor U10955 (N_10955,N_10865,N_10817);
nor U10956 (N_10956,N_10871,N_10781);
or U10957 (N_10957,N_10823,N_10796);
xnor U10958 (N_10958,N_10747,N_10852);
xor U10959 (N_10959,N_10763,N_10755);
and U10960 (N_10960,N_10855,N_10849);
and U10961 (N_10961,N_10736,N_10758);
nand U10962 (N_10962,N_10770,N_10820);
and U10963 (N_10963,N_10808,N_10765);
xnor U10964 (N_10964,N_10745,N_10760);
or U10965 (N_10965,N_10744,N_10799);
or U10966 (N_10966,N_10778,N_10789);
nor U10967 (N_10967,N_10734,N_10813);
or U10968 (N_10968,N_10840,N_10789);
nor U10969 (N_10969,N_10793,N_10875);
nand U10970 (N_10970,N_10810,N_10876);
xor U10971 (N_10971,N_10778,N_10874);
nand U10972 (N_10972,N_10738,N_10807);
and U10973 (N_10973,N_10724,N_10866);
nand U10974 (N_10974,N_10868,N_10781);
and U10975 (N_10975,N_10816,N_10803);
and U10976 (N_10976,N_10877,N_10825);
nand U10977 (N_10977,N_10787,N_10831);
nor U10978 (N_10978,N_10824,N_10758);
nand U10979 (N_10979,N_10831,N_10729);
or U10980 (N_10980,N_10878,N_10835);
nor U10981 (N_10981,N_10831,N_10870);
xnor U10982 (N_10982,N_10786,N_10864);
nor U10983 (N_10983,N_10753,N_10845);
nor U10984 (N_10984,N_10858,N_10782);
nor U10985 (N_10985,N_10824,N_10825);
nand U10986 (N_10986,N_10858,N_10831);
nor U10987 (N_10987,N_10781,N_10813);
nand U10988 (N_10988,N_10720,N_10837);
nor U10989 (N_10989,N_10744,N_10772);
or U10990 (N_10990,N_10730,N_10725);
nor U10991 (N_10991,N_10774,N_10799);
nand U10992 (N_10992,N_10781,N_10768);
or U10993 (N_10993,N_10737,N_10755);
xor U10994 (N_10994,N_10827,N_10782);
nand U10995 (N_10995,N_10777,N_10783);
nor U10996 (N_10996,N_10792,N_10745);
and U10997 (N_10997,N_10810,N_10723);
xnor U10998 (N_10998,N_10765,N_10824);
xor U10999 (N_10999,N_10867,N_10786);
nand U11000 (N_11000,N_10843,N_10778);
nand U11001 (N_11001,N_10872,N_10734);
or U11002 (N_11002,N_10819,N_10856);
nand U11003 (N_11003,N_10859,N_10746);
nand U11004 (N_11004,N_10768,N_10766);
nor U11005 (N_11005,N_10830,N_10774);
xnor U11006 (N_11006,N_10854,N_10753);
or U11007 (N_11007,N_10806,N_10740);
nand U11008 (N_11008,N_10736,N_10727);
nand U11009 (N_11009,N_10819,N_10833);
xor U11010 (N_11010,N_10848,N_10750);
nand U11011 (N_11011,N_10822,N_10799);
nor U11012 (N_11012,N_10807,N_10834);
nor U11013 (N_11013,N_10837,N_10795);
or U11014 (N_11014,N_10751,N_10794);
nor U11015 (N_11015,N_10804,N_10835);
or U11016 (N_11016,N_10796,N_10721);
nor U11017 (N_11017,N_10800,N_10806);
xor U11018 (N_11018,N_10734,N_10845);
xnor U11019 (N_11019,N_10720,N_10725);
nand U11020 (N_11020,N_10730,N_10829);
nor U11021 (N_11021,N_10773,N_10830);
xnor U11022 (N_11022,N_10798,N_10828);
xor U11023 (N_11023,N_10735,N_10752);
xnor U11024 (N_11024,N_10749,N_10804);
nor U11025 (N_11025,N_10785,N_10731);
nor U11026 (N_11026,N_10757,N_10772);
xor U11027 (N_11027,N_10790,N_10820);
xnor U11028 (N_11028,N_10867,N_10737);
and U11029 (N_11029,N_10772,N_10785);
xnor U11030 (N_11030,N_10749,N_10791);
and U11031 (N_11031,N_10772,N_10848);
and U11032 (N_11032,N_10764,N_10829);
and U11033 (N_11033,N_10800,N_10861);
nor U11034 (N_11034,N_10860,N_10798);
nor U11035 (N_11035,N_10837,N_10870);
nand U11036 (N_11036,N_10874,N_10776);
nor U11037 (N_11037,N_10870,N_10784);
xnor U11038 (N_11038,N_10775,N_10769);
nand U11039 (N_11039,N_10810,N_10835);
nand U11040 (N_11040,N_10892,N_10902);
nor U11041 (N_11041,N_10924,N_10980);
and U11042 (N_11042,N_11022,N_10944);
and U11043 (N_11043,N_10885,N_10925);
xor U11044 (N_11044,N_11006,N_10936);
or U11045 (N_11045,N_10880,N_10927);
and U11046 (N_11046,N_10958,N_10966);
xnor U11047 (N_11047,N_10981,N_10881);
nand U11048 (N_11048,N_10913,N_10912);
or U11049 (N_11049,N_11035,N_10928);
nor U11050 (N_11050,N_10973,N_10900);
or U11051 (N_11051,N_10992,N_10897);
xor U11052 (N_11052,N_10931,N_10988);
nand U11053 (N_11053,N_11020,N_10914);
or U11054 (N_11054,N_10984,N_10976);
or U11055 (N_11055,N_10887,N_10956);
nor U11056 (N_11056,N_10895,N_10933);
and U11057 (N_11057,N_10985,N_10957);
nor U11058 (N_11058,N_11023,N_10923);
or U11059 (N_11059,N_10882,N_10899);
and U11060 (N_11060,N_10905,N_10962);
nand U11061 (N_11061,N_10948,N_10911);
and U11062 (N_11062,N_10888,N_10995);
or U11063 (N_11063,N_10954,N_11026);
nand U11064 (N_11064,N_10916,N_10907);
nor U11065 (N_11065,N_10996,N_10896);
or U11066 (N_11066,N_11007,N_10953);
nor U11067 (N_11067,N_10974,N_11025);
xor U11068 (N_11068,N_10978,N_10909);
xnor U11069 (N_11069,N_11030,N_10910);
xnor U11070 (N_11070,N_10891,N_10965);
xor U11071 (N_11071,N_11010,N_11034);
nand U11072 (N_11072,N_10938,N_11019);
and U11073 (N_11073,N_10918,N_10898);
nand U11074 (N_11074,N_10975,N_10951);
xor U11075 (N_11075,N_10935,N_10982);
nor U11076 (N_11076,N_10937,N_10952);
nor U11077 (N_11077,N_10964,N_10960);
and U11078 (N_11078,N_11039,N_10959);
nor U11079 (N_11079,N_11011,N_10943);
nor U11080 (N_11080,N_10886,N_10919);
or U11081 (N_11081,N_11033,N_11027);
nor U11082 (N_11082,N_10929,N_11018);
or U11083 (N_11083,N_10920,N_11029);
nand U11084 (N_11084,N_10986,N_10945);
nor U11085 (N_11085,N_10983,N_10998);
and U11086 (N_11086,N_10915,N_11032);
xor U11087 (N_11087,N_11000,N_11016);
nor U11088 (N_11088,N_10989,N_10921);
nor U11089 (N_11089,N_10967,N_10926);
xnor U11090 (N_11090,N_10949,N_10941);
or U11091 (N_11091,N_11031,N_11012);
and U11092 (N_11092,N_11015,N_11028);
nor U11093 (N_11093,N_11036,N_10971);
nand U11094 (N_11094,N_10979,N_11024);
nor U11095 (N_11095,N_11037,N_11004);
nand U11096 (N_11096,N_10997,N_10968);
and U11097 (N_11097,N_10884,N_10894);
or U11098 (N_11098,N_10950,N_10890);
or U11099 (N_11099,N_10939,N_11017);
or U11100 (N_11100,N_10901,N_10947);
and U11101 (N_11101,N_11014,N_11002);
and U11102 (N_11102,N_10977,N_10930);
or U11103 (N_11103,N_10889,N_11003);
nand U11104 (N_11104,N_10970,N_10946);
or U11105 (N_11105,N_10903,N_11005);
nor U11106 (N_11106,N_11001,N_10955);
and U11107 (N_11107,N_10972,N_10994);
or U11108 (N_11108,N_10963,N_10990);
xnor U11109 (N_11109,N_10987,N_10917);
xnor U11110 (N_11110,N_10906,N_11008);
nor U11111 (N_11111,N_10893,N_10883);
or U11112 (N_11112,N_11013,N_10904);
and U11113 (N_11113,N_10908,N_10999);
and U11114 (N_11114,N_10940,N_11038);
nor U11115 (N_11115,N_10991,N_10932);
or U11116 (N_11116,N_10934,N_11021);
and U11117 (N_11117,N_11009,N_10969);
nor U11118 (N_11118,N_10961,N_10993);
xnor U11119 (N_11119,N_10942,N_10922);
xor U11120 (N_11120,N_10942,N_10972);
xor U11121 (N_11121,N_10979,N_10922);
nand U11122 (N_11122,N_10922,N_10971);
nand U11123 (N_11123,N_10896,N_10906);
or U11124 (N_11124,N_10984,N_10969);
nor U11125 (N_11125,N_10899,N_11013);
nor U11126 (N_11126,N_10897,N_10937);
or U11127 (N_11127,N_10998,N_10951);
xnor U11128 (N_11128,N_10993,N_10990);
nand U11129 (N_11129,N_10993,N_11024);
and U11130 (N_11130,N_10930,N_10922);
nor U11131 (N_11131,N_10989,N_10984);
or U11132 (N_11132,N_10887,N_10892);
nor U11133 (N_11133,N_10964,N_10934);
and U11134 (N_11134,N_10882,N_11031);
or U11135 (N_11135,N_10995,N_11016);
nor U11136 (N_11136,N_10980,N_10977);
nand U11137 (N_11137,N_10996,N_10899);
and U11138 (N_11138,N_11030,N_11038);
nor U11139 (N_11139,N_10950,N_11005);
or U11140 (N_11140,N_10934,N_10986);
nand U11141 (N_11141,N_10936,N_10882);
or U11142 (N_11142,N_11034,N_10891);
nor U11143 (N_11143,N_11019,N_10894);
xor U11144 (N_11144,N_11027,N_10954);
nand U11145 (N_11145,N_11015,N_10948);
xnor U11146 (N_11146,N_10950,N_10960);
xnor U11147 (N_11147,N_10938,N_10955);
nand U11148 (N_11148,N_10945,N_10965);
or U11149 (N_11149,N_11037,N_10882);
and U11150 (N_11150,N_10972,N_11016);
and U11151 (N_11151,N_11020,N_10917);
or U11152 (N_11152,N_10943,N_10940);
nor U11153 (N_11153,N_10926,N_10933);
or U11154 (N_11154,N_10942,N_10903);
nand U11155 (N_11155,N_11033,N_10904);
or U11156 (N_11156,N_11008,N_10888);
nand U11157 (N_11157,N_10985,N_10981);
or U11158 (N_11158,N_10908,N_10934);
or U11159 (N_11159,N_10932,N_10947);
nor U11160 (N_11160,N_10940,N_10984);
nand U11161 (N_11161,N_10897,N_10941);
and U11162 (N_11162,N_10926,N_10912);
and U11163 (N_11163,N_11007,N_11016);
xor U11164 (N_11164,N_10985,N_10894);
nor U11165 (N_11165,N_10891,N_11030);
and U11166 (N_11166,N_11019,N_10969);
nor U11167 (N_11167,N_10947,N_10883);
xor U11168 (N_11168,N_10887,N_11005);
nand U11169 (N_11169,N_10963,N_10916);
and U11170 (N_11170,N_11018,N_10991);
and U11171 (N_11171,N_10903,N_10990);
xnor U11172 (N_11172,N_11026,N_10989);
xor U11173 (N_11173,N_10930,N_10957);
and U11174 (N_11174,N_11008,N_10908);
or U11175 (N_11175,N_11005,N_10991);
or U11176 (N_11176,N_10942,N_10909);
nand U11177 (N_11177,N_10979,N_10889);
nand U11178 (N_11178,N_10958,N_10911);
nor U11179 (N_11179,N_10906,N_10933);
or U11180 (N_11180,N_10896,N_10998);
nor U11181 (N_11181,N_11013,N_10908);
or U11182 (N_11182,N_10927,N_11005);
xnor U11183 (N_11183,N_10906,N_10991);
nor U11184 (N_11184,N_10989,N_10917);
nand U11185 (N_11185,N_10986,N_10963);
and U11186 (N_11186,N_10925,N_10931);
xnor U11187 (N_11187,N_11015,N_10900);
nand U11188 (N_11188,N_10949,N_10990);
xnor U11189 (N_11189,N_10920,N_10955);
nand U11190 (N_11190,N_10974,N_10959);
nand U11191 (N_11191,N_10884,N_10973);
and U11192 (N_11192,N_11023,N_10903);
nand U11193 (N_11193,N_10981,N_10927);
nand U11194 (N_11194,N_10933,N_11031);
xor U11195 (N_11195,N_10947,N_10894);
nand U11196 (N_11196,N_11012,N_10927);
and U11197 (N_11197,N_11002,N_10926);
xnor U11198 (N_11198,N_10942,N_11004);
and U11199 (N_11199,N_11010,N_10898);
or U11200 (N_11200,N_11086,N_11083);
xor U11201 (N_11201,N_11127,N_11118);
nand U11202 (N_11202,N_11191,N_11189);
or U11203 (N_11203,N_11080,N_11162);
nand U11204 (N_11204,N_11051,N_11053);
and U11205 (N_11205,N_11062,N_11193);
and U11206 (N_11206,N_11199,N_11185);
xnor U11207 (N_11207,N_11197,N_11181);
xor U11208 (N_11208,N_11098,N_11131);
xor U11209 (N_11209,N_11078,N_11151);
and U11210 (N_11210,N_11190,N_11161);
or U11211 (N_11211,N_11154,N_11071);
nor U11212 (N_11212,N_11043,N_11050);
nor U11213 (N_11213,N_11066,N_11110);
and U11214 (N_11214,N_11124,N_11088);
nor U11215 (N_11215,N_11113,N_11158);
nor U11216 (N_11216,N_11040,N_11076);
nor U11217 (N_11217,N_11145,N_11064);
xor U11218 (N_11218,N_11093,N_11128);
nor U11219 (N_11219,N_11049,N_11107);
and U11220 (N_11220,N_11070,N_11090);
and U11221 (N_11221,N_11123,N_11069);
and U11222 (N_11222,N_11100,N_11108);
and U11223 (N_11223,N_11099,N_11058);
and U11224 (N_11224,N_11101,N_11041);
and U11225 (N_11225,N_11106,N_11065);
nor U11226 (N_11226,N_11104,N_11075);
or U11227 (N_11227,N_11055,N_11175);
and U11228 (N_11228,N_11091,N_11116);
nand U11229 (N_11229,N_11094,N_11188);
nor U11230 (N_11230,N_11112,N_11081);
or U11231 (N_11231,N_11172,N_11173);
nor U11232 (N_11232,N_11138,N_11186);
nand U11233 (N_11233,N_11120,N_11117);
nor U11234 (N_11234,N_11177,N_11044);
and U11235 (N_11235,N_11157,N_11178);
and U11236 (N_11236,N_11130,N_11109);
xnor U11237 (N_11237,N_11060,N_11160);
nor U11238 (N_11238,N_11056,N_11115);
nand U11239 (N_11239,N_11103,N_11059);
nand U11240 (N_11240,N_11129,N_11140);
nand U11241 (N_11241,N_11159,N_11144);
and U11242 (N_11242,N_11196,N_11139);
xor U11243 (N_11243,N_11169,N_11136);
xnor U11244 (N_11244,N_11152,N_11195);
nor U11245 (N_11245,N_11052,N_11167);
and U11246 (N_11246,N_11174,N_11184);
xnor U11247 (N_11247,N_11163,N_11135);
or U11248 (N_11248,N_11121,N_11133);
xnor U11249 (N_11249,N_11054,N_11150);
xor U11250 (N_11250,N_11179,N_11048);
xnor U11251 (N_11251,N_11180,N_11143);
nor U11252 (N_11252,N_11182,N_11105);
nor U11253 (N_11253,N_11155,N_11156);
nand U11254 (N_11254,N_11102,N_11097);
and U11255 (N_11255,N_11089,N_11063);
and U11256 (N_11256,N_11057,N_11082);
nand U11257 (N_11257,N_11148,N_11192);
or U11258 (N_11258,N_11068,N_11149);
and U11259 (N_11259,N_11176,N_11198);
nor U11260 (N_11260,N_11072,N_11164);
xnor U11261 (N_11261,N_11045,N_11153);
xnor U11262 (N_11262,N_11077,N_11141);
or U11263 (N_11263,N_11170,N_11165);
nand U11264 (N_11264,N_11046,N_11084);
and U11265 (N_11265,N_11111,N_11079);
nand U11266 (N_11266,N_11142,N_11134);
nand U11267 (N_11267,N_11114,N_11073);
nor U11268 (N_11268,N_11171,N_11122);
nor U11269 (N_11269,N_11047,N_11126);
or U11270 (N_11270,N_11146,N_11125);
nand U11271 (N_11271,N_11067,N_11166);
and U11272 (N_11272,N_11137,N_11187);
nor U11273 (N_11273,N_11147,N_11132);
nor U11274 (N_11274,N_11095,N_11119);
nand U11275 (N_11275,N_11061,N_11096);
xor U11276 (N_11276,N_11074,N_11042);
nand U11277 (N_11277,N_11087,N_11092);
nand U11278 (N_11278,N_11194,N_11168);
or U11279 (N_11279,N_11085,N_11183);
nand U11280 (N_11280,N_11179,N_11150);
and U11281 (N_11281,N_11113,N_11071);
nor U11282 (N_11282,N_11123,N_11175);
nand U11283 (N_11283,N_11066,N_11067);
nand U11284 (N_11284,N_11128,N_11144);
and U11285 (N_11285,N_11051,N_11087);
or U11286 (N_11286,N_11182,N_11144);
xnor U11287 (N_11287,N_11149,N_11120);
or U11288 (N_11288,N_11143,N_11109);
xnor U11289 (N_11289,N_11074,N_11087);
and U11290 (N_11290,N_11091,N_11177);
nand U11291 (N_11291,N_11106,N_11133);
xor U11292 (N_11292,N_11103,N_11137);
nand U11293 (N_11293,N_11072,N_11165);
nor U11294 (N_11294,N_11053,N_11106);
and U11295 (N_11295,N_11081,N_11051);
nor U11296 (N_11296,N_11089,N_11076);
xnor U11297 (N_11297,N_11114,N_11143);
or U11298 (N_11298,N_11130,N_11185);
xor U11299 (N_11299,N_11072,N_11127);
and U11300 (N_11300,N_11145,N_11123);
nor U11301 (N_11301,N_11060,N_11180);
or U11302 (N_11302,N_11153,N_11105);
xnor U11303 (N_11303,N_11199,N_11165);
xnor U11304 (N_11304,N_11141,N_11061);
or U11305 (N_11305,N_11089,N_11120);
and U11306 (N_11306,N_11075,N_11114);
nor U11307 (N_11307,N_11042,N_11063);
nand U11308 (N_11308,N_11061,N_11189);
xor U11309 (N_11309,N_11093,N_11136);
nor U11310 (N_11310,N_11092,N_11140);
and U11311 (N_11311,N_11144,N_11122);
xnor U11312 (N_11312,N_11190,N_11165);
and U11313 (N_11313,N_11045,N_11084);
nor U11314 (N_11314,N_11166,N_11121);
or U11315 (N_11315,N_11149,N_11115);
or U11316 (N_11316,N_11064,N_11166);
or U11317 (N_11317,N_11113,N_11085);
xor U11318 (N_11318,N_11082,N_11149);
or U11319 (N_11319,N_11083,N_11167);
or U11320 (N_11320,N_11132,N_11181);
nor U11321 (N_11321,N_11107,N_11081);
or U11322 (N_11322,N_11093,N_11147);
or U11323 (N_11323,N_11139,N_11081);
xnor U11324 (N_11324,N_11124,N_11051);
or U11325 (N_11325,N_11192,N_11126);
nand U11326 (N_11326,N_11055,N_11192);
nand U11327 (N_11327,N_11063,N_11165);
and U11328 (N_11328,N_11194,N_11086);
and U11329 (N_11329,N_11049,N_11134);
nand U11330 (N_11330,N_11164,N_11154);
xor U11331 (N_11331,N_11190,N_11172);
and U11332 (N_11332,N_11104,N_11161);
and U11333 (N_11333,N_11109,N_11060);
xor U11334 (N_11334,N_11171,N_11198);
or U11335 (N_11335,N_11110,N_11165);
or U11336 (N_11336,N_11057,N_11153);
and U11337 (N_11337,N_11167,N_11117);
and U11338 (N_11338,N_11052,N_11113);
or U11339 (N_11339,N_11108,N_11154);
xnor U11340 (N_11340,N_11105,N_11163);
nand U11341 (N_11341,N_11081,N_11083);
xnor U11342 (N_11342,N_11134,N_11136);
and U11343 (N_11343,N_11196,N_11130);
or U11344 (N_11344,N_11083,N_11043);
and U11345 (N_11345,N_11094,N_11127);
nand U11346 (N_11346,N_11073,N_11076);
nand U11347 (N_11347,N_11192,N_11165);
and U11348 (N_11348,N_11100,N_11110);
nor U11349 (N_11349,N_11084,N_11079);
and U11350 (N_11350,N_11055,N_11188);
xnor U11351 (N_11351,N_11066,N_11157);
nand U11352 (N_11352,N_11168,N_11164);
and U11353 (N_11353,N_11166,N_11072);
nor U11354 (N_11354,N_11046,N_11165);
xnor U11355 (N_11355,N_11103,N_11104);
xor U11356 (N_11356,N_11136,N_11167);
and U11357 (N_11357,N_11080,N_11041);
xor U11358 (N_11358,N_11187,N_11147);
nand U11359 (N_11359,N_11162,N_11133);
nand U11360 (N_11360,N_11354,N_11314);
nor U11361 (N_11361,N_11277,N_11344);
xnor U11362 (N_11362,N_11234,N_11300);
or U11363 (N_11363,N_11356,N_11342);
nand U11364 (N_11364,N_11238,N_11301);
xor U11365 (N_11365,N_11228,N_11321);
and U11366 (N_11366,N_11340,N_11259);
nand U11367 (N_11367,N_11288,N_11231);
nor U11368 (N_11368,N_11313,N_11303);
nand U11369 (N_11369,N_11355,N_11248);
and U11370 (N_11370,N_11233,N_11309);
nand U11371 (N_11371,N_11275,N_11346);
nor U11372 (N_11372,N_11345,N_11208);
nor U11373 (N_11373,N_11261,N_11251);
and U11374 (N_11374,N_11333,N_11212);
and U11375 (N_11375,N_11265,N_11331);
or U11376 (N_11376,N_11278,N_11337);
or U11377 (N_11377,N_11257,N_11310);
xnor U11378 (N_11378,N_11217,N_11292);
nand U11379 (N_11379,N_11247,N_11357);
nand U11380 (N_11380,N_11267,N_11326);
xnor U11381 (N_11381,N_11211,N_11243);
nand U11382 (N_11382,N_11287,N_11341);
nor U11383 (N_11383,N_11282,N_11245);
xor U11384 (N_11384,N_11317,N_11249);
nand U11385 (N_11385,N_11335,N_11242);
nor U11386 (N_11386,N_11237,N_11350);
nor U11387 (N_11387,N_11329,N_11306);
and U11388 (N_11388,N_11283,N_11284);
nor U11389 (N_11389,N_11347,N_11236);
and U11390 (N_11390,N_11320,N_11264);
or U11391 (N_11391,N_11200,N_11268);
nand U11392 (N_11392,N_11305,N_11297);
or U11393 (N_11393,N_11271,N_11304);
or U11394 (N_11394,N_11227,N_11244);
nor U11395 (N_11395,N_11316,N_11307);
xnor U11396 (N_11396,N_11235,N_11299);
xnor U11397 (N_11397,N_11328,N_11296);
nor U11398 (N_11398,N_11215,N_11323);
nor U11399 (N_11399,N_11325,N_11281);
nand U11400 (N_11400,N_11239,N_11339);
nor U11401 (N_11401,N_11302,N_11260);
nand U11402 (N_11402,N_11241,N_11222);
xor U11403 (N_11403,N_11358,N_11338);
nor U11404 (N_11404,N_11359,N_11308);
or U11405 (N_11405,N_11312,N_11322);
and U11406 (N_11406,N_11298,N_11226);
nand U11407 (N_11407,N_11221,N_11294);
and U11408 (N_11408,N_11258,N_11279);
xor U11409 (N_11409,N_11295,N_11280);
xnor U11410 (N_11410,N_11210,N_11262);
nand U11411 (N_11411,N_11327,N_11270);
nand U11412 (N_11412,N_11351,N_11254);
nor U11413 (N_11413,N_11223,N_11240);
nand U11414 (N_11414,N_11213,N_11311);
nand U11415 (N_11415,N_11207,N_11209);
nor U11416 (N_11416,N_11202,N_11269);
and U11417 (N_11417,N_11224,N_11343);
or U11418 (N_11418,N_11205,N_11290);
nand U11419 (N_11419,N_11289,N_11246);
nand U11420 (N_11420,N_11218,N_11255);
and U11421 (N_11421,N_11336,N_11225);
nand U11422 (N_11422,N_11285,N_11286);
nor U11423 (N_11423,N_11324,N_11276);
or U11424 (N_11424,N_11272,N_11266);
nor U11425 (N_11425,N_11230,N_11253);
or U11426 (N_11426,N_11204,N_11332);
xor U11427 (N_11427,N_11252,N_11352);
and U11428 (N_11428,N_11273,N_11220);
nand U11429 (N_11429,N_11353,N_11330);
nand U11430 (N_11430,N_11206,N_11315);
or U11431 (N_11431,N_11203,N_11319);
nand U11432 (N_11432,N_11263,N_11232);
xnor U11433 (N_11433,N_11348,N_11250);
and U11434 (N_11434,N_11291,N_11214);
xor U11435 (N_11435,N_11256,N_11334);
nand U11436 (N_11436,N_11219,N_11229);
and U11437 (N_11437,N_11274,N_11216);
xnor U11438 (N_11438,N_11349,N_11318);
xnor U11439 (N_11439,N_11201,N_11293);
nand U11440 (N_11440,N_11312,N_11260);
xor U11441 (N_11441,N_11305,N_11238);
and U11442 (N_11442,N_11288,N_11273);
and U11443 (N_11443,N_11264,N_11330);
nor U11444 (N_11444,N_11248,N_11305);
nor U11445 (N_11445,N_11210,N_11205);
nor U11446 (N_11446,N_11243,N_11205);
xor U11447 (N_11447,N_11333,N_11310);
xnor U11448 (N_11448,N_11231,N_11339);
nand U11449 (N_11449,N_11327,N_11273);
nor U11450 (N_11450,N_11275,N_11358);
and U11451 (N_11451,N_11208,N_11219);
and U11452 (N_11452,N_11246,N_11334);
nor U11453 (N_11453,N_11243,N_11270);
and U11454 (N_11454,N_11270,N_11252);
and U11455 (N_11455,N_11251,N_11266);
or U11456 (N_11456,N_11353,N_11218);
nand U11457 (N_11457,N_11293,N_11314);
nor U11458 (N_11458,N_11241,N_11244);
or U11459 (N_11459,N_11263,N_11255);
xor U11460 (N_11460,N_11278,N_11261);
or U11461 (N_11461,N_11308,N_11246);
and U11462 (N_11462,N_11249,N_11267);
or U11463 (N_11463,N_11229,N_11322);
nand U11464 (N_11464,N_11282,N_11302);
xnor U11465 (N_11465,N_11354,N_11313);
or U11466 (N_11466,N_11305,N_11262);
nor U11467 (N_11467,N_11311,N_11223);
or U11468 (N_11468,N_11345,N_11218);
and U11469 (N_11469,N_11206,N_11299);
or U11470 (N_11470,N_11242,N_11222);
or U11471 (N_11471,N_11221,N_11280);
or U11472 (N_11472,N_11215,N_11318);
and U11473 (N_11473,N_11236,N_11278);
or U11474 (N_11474,N_11303,N_11295);
nor U11475 (N_11475,N_11232,N_11358);
xnor U11476 (N_11476,N_11245,N_11323);
nand U11477 (N_11477,N_11319,N_11311);
xor U11478 (N_11478,N_11244,N_11315);
nand U11479 (N_11479,N_11261,N_11339);
nor U11480 (N_11480,N_11233,N_11319);
nand U11481 (N_11481,N_11301,N_11302);
xor U11482 (N_11482,N_11268,N_11348);
xnor U11483 (N_11483,N_11214,N_11205);
or U11484 (N_11484,N_11346,N_11287);
and U11485 (N_11485,N_11327,N_11240);
or U11486 (N_11486,N_11307,N_11302);
xnor U11487 (N_11487,N_11229,N_11232);
xnor U11488 (N_11488,N_11322,N_11219);
nand U11489 (N_11489,N_11251,N_11326);
and U11490 (N_11490,N_11334,N_11265);
and U11491 (N_11491,N_11229,N_11349);
and U11492 (N_11492,N_11275,N_11318);
nor U11493 (N_11493,N_11258,N_11237);
or U11494 (N_11494,N_11347,N_11301);
nand U11495 (N_11495,N_11296,N_11279);
nor U11496 (N_11496,N_11307,N_11251);
nor U11497 (N_11497,N_11283,N_11290);
nor U11498 (N_11498,N_11238,N_11303);
or U11499 (N_11499,N_11275,N_11329);
and U11500 (N_11500,N_11234,N_11338);
nand U11501 (N_11501,N_11205,N_11342);
nand U11502 (N_11502,N_11289,N_11341);
nor U11503 (N_11503,N_11201,N_11342);
nand U11504 (N_11504,N_11299,N_11214);
nand U11505 (N_11505,N_11206,N_11223);
xnor U11506 (N_11506,N_11273,N_11330);
xnor U11507 (N_11507,N_11231,N_11253);
or U11508 (N_11508,N_11212,N_11295);
or U11509 (N_11509,N_11253,N_11333);
xnor U11510 (N_11510,N_11281,N_11280);
nor U11511 (N_11511,N_11277,N_11305);
nor U11512 (N_11512,N_11353,N_11271);
xor U11513 (N_11513,N_11352,N_11356);
or U11514 (N_11514,N_11359,N_11283);
or U11515 (N_11515,N_11222,N_11221);
nand U11516 (N_11516,N_11278,N_11275);
nor U11517 (N_11517,N_11261,N_11227);
nand U11518 (N_11518,N_11249,N_11315);
xor U11519 (N_11519,N_11242,N_11354);
xor U11520 (N_11520,N_11502,N_11368);
xor U11521 (N_11521,N_11397,N_11395);
and U11522 (N_11522,N_11492,N_11470);
and U11523 (N_11523,N_11366,N_11391);
and U11524 (N_11524,N_11414,N_11386);
or U11525 (N_11525,N_11394,N_11387);
nor U11526 (N_11526,N_11493,N_11474);
or U11527 (N_11527,N_11392,N_11458);
and U11528 (N_11528,N_11477,N_11385);
or U11529 (N_11529,N_11503,N_11370);
nand U11530 (N_11530,N_11425,N_11419);
nand U11531 (N_11531,N_11409,N_11390);
or U11532 (N_11532,N_11465,N_11420);
or U11533 (N_11533,N_11508,N_11518);
and U11534 (N_11534,N_11369,N_11371);
or U11535 (N_11535,N_11475,N_11367);
nor U11536 (N_11536,N_11444,N_11380);
or U11537 (N_11537,N_11483,N_11360);
nor U11538 (N_11538,N_11401,N_11450);
and U11539 (N_11539,N_11512,N_11399);
xor U11540 (N_11540,N_11376,N_11519);
nor U11541 (N_11541,N_11382,N_11457);
or U11542 (N_11542,N_11490,N_11421);
nor U11543 (N_11543,N_11495,N_11476);
or U11544 (N_11544,N_11473,N_11393);
nand U11545 (N_11545,N_11375,N_11484);
xnor U11546 (N_11546,N_11515,N_11383);
nor U11547 (N_11547,N_11441,N_11374);
xor U11548 (N_11548,N_11491,N_11511);
xor U11549 (N_11549,N_11428,N_11389);
nand U11550 (N_11550,N_11417,N_11378);
nor U11551 (N_11551,N_11373,N_11415);
nand U11552 (N_11552,N_11468,N_11498);
and U11553 (N_11553,N_11361,N_11388);
or U11554 (N_11554,N_11488,N_11422);
xnor U11555 (N_11555,N_11497,N_11471);
xnor U11556 (N_11556,N_11424,N_11451);
or U11557 (N_11557,N_11403,N_11440);
or U11558 (N_11558,N_11442,N_11411);
nand U11559 (N_11559,N_11501,N_11400);
xnor U11560 (N_11560,N_11460,N_11446);
or U11561 (N_11561,N_11453,N_11410);
or U11562 (N_11562,N_11384,N_11506);
and U11563 (N_11563,N_11485,N_11472);
and U11564 (N_11564,N_11447,N_11456);
nor U11565 (N_11565,N_11407,N_11429);
and U11566 (N_11566,N_11412,N_11402);
nor U11567 (N_11567,N_11364,N_11396);
nand U11568 (N_11568,N_11459,N_11433);
or U11569 (N_11569,N_11455,N_11449);
nor U11570 (N_11570,N_11513,N_11418);
nor U11571 (N_11571,N_11365,N_11504);
nor U11572 (N_11572,N_11436,N_11517);
xor U11573 (N_11573,N_11462,N_11416);
xnor U11574 (N_11574,N_11467,N_11486);
nand U11575 (N_11575,N_11408,N_11480);
xnor U11576 (N_11576,N_11505,N_11398);
xnor U11577 (N_11577,N_11466,N_11464);
xnor U11578 (N_11578,N_11481,N_11372);
nor U11579 (N_11579,N_11431,N_11496);
nor U11580 (N_11580,N_11439,N_11463);
nor U11581 (N_11581,N_11432,N_11379);
nand U11582 (N_11582,N_11426,N_11404);
and U11583 (N_11583,N_11507,N_11509);
or U11584 (N_11584,N_11514,N_11377);
or U11585 (N_11585,N_11434,N_11438);
nand U11586 (N_11586,N_11499,N_11500);
nor U11587 (N_11587,N_11448,N_11405);
nand U11588 (N_11588,N_11381,N_11363);
xnor U11589 (N_11589,N_11362,N_11406);
xor U11590 (N_11590,N_11452,N_11443);
nand U11591 (N_11591,N_11437,N_11494);
nor U11592 (N_11592,N_11435,N_11454);
xnor U11593 (N_11593,N_11423,N_11516);
xor U11594 (N_11594,N_11489,N_11430);
nand U11595 (N_11595,N_11479,N_11487);
or U11596 (N_11596,N_11461,N_11482);
xnor U11597 (N_11597,N_11469,N_11427);
nand U11598 (N_11598,N_11445,N_11413);
xnor U11599 (N_11599,N_11478,N_11510);
xnor U11600 (N_11600,N_11445,N_11451);
and U11601 (N_11601,N_11395,N_11474);
and U11602 (N_11602,N_11389,N_11366);
nand U11603 (N_11603,N_11421,N_11417);
xor U11604 (N_11604,N_11470,N_11373);
and U11605 (N_11605,N_11508,N_11465);
nand U11606 (N_11606,N_11404,N_11382);
xor U11607 (N_11607,N_11412,N_11469);
nor U11608 (N_11608,N_11429,N_11367);
nand U11609 (N_11609,N_11423,N_11395);
xnor U11610 (N_11610,N_11438,N_11396);
nor U11611 (N_11611,N_11405,N_11386);
and U11612 (N_11612,N_11368,N_11507);
nand U11613 (N_11613,N_11408,N_11510);
or U11614 (N_11614,N_11504,N_11412);
nor U11615 (N_11615,N_11440,N_11452);
nor U11616 (N_11616,N_11399,N_11489);
and U11617 (N_11617,N_11399,N_11360);
or U11618 (N_11618,N_11464,N_11507);
or U11619 (N_11619,N_11504,N_11390);
and U11620 (N_11620,N_11430,N_11376);
nor U11621 (N_11621,N_11517,N_11380);
xor U11622 (N_11622,N_11508,N_11517);
nor U11623 (N_11623,N_11430,N_11456);
or U11624 (N_11624,N_11368,N_11403);
xnor U11625 (N_11625,N_11435,N_11455);
nor U11626 (N_11626,N_11504,N_11498);
nor U11627 (N_11627,N_11486,N_11420);
xnor U11628 (N_11628,N_11426,N_11399);
xor U11629 (N_11629,N_11370,N_11485);
nor U11630 (N_11630,N_11515,N_11384);
or U11631 (N_11631,N_11373,N_11393);
xnor U11632 (N_11632,N_11371,N_11416);
xor U11633 (N_11633,N_11487,N_11476);
xnor U11634 (N_11634,N_11436,N_11433);
and U11635 (N_11635,N_11445,N_11487);
or U11636 (N_11636,N_11434,N_11424);
nor U11637 (N_11637,N_11415,N_11504);
nor U11638 (N_11638,N_11455,N_11416);
nor U11639 (N_11639,N_11499,N_11385);
nand U11640 (N_11640,N_11400,N_11418);
and U11641 (N_11641,N_11473,N_11419);
xnor U11642 (N_11642,N_11481,N_11432);
nand U11643 (N_11643,N_11449,N_11385);
or U11644 (N_11644,N_11486,N_11387);
nand U11645 (N_11645,N_11465,N_11505);
or U11646 (N_11646,N_11462,N_11483);
and U11647 (N_11647,N_11466,N_11424);
nor U11648 (N_11648,N_11466,N_11384);
nand U11649 (N_11649,N_11419,N_11469);
or U11650 (N_11650,N_11412,N_11360);
xor U11651 (N_11651,N_11402,N_11475);
or U11652 (N_11652,N_11507,N_11385);
nand U11653 (N_11653,N_11409,N_11451);
nor U11654 (N_11654,N_11469,N_11479);
xnor U11655 (N_11655,N_11374,N_11442);
xor U11656 (N_11656,N_11431,N_11429);
and U11657 (N_11657,N_11412,N_11450);
nand U11658 (N_11658,N_11453,N_11462);
nand U11659 (N_11659,N_11497,N_11509);
nor U11660 (N_11660,N_11387,N_11370);
and U11661 (N_11661,N_11385,N_11489);
or U11662 (N_11662,N_11470,N_11430);
nor U11663 (N_11663,N_11392,N_11491);
or U11664 (N_11664,N_11439,N_11436);
nor U11665 (N_11665,N_11512,N_11443);
and U11666 (N_11666,N_11478,N_11409);
or U11667 (N_11667,N_11474,N_11451);
and U11668 (N_11668,N_11497,N_11398);
or U11669 (N_11669,N_11508,N_11434);
xnor U11670 (N_11670,N_11494,N_11393);
xor U11671 (N_11671,N_11493,N_11449);
nor U11672 (N_11672,N_11460,N_11371);
xor U11673 (N_11673,N_11386,N_11427);
nor U11674 (N_11674,N_11479,N_11435);
or U11675 (N_11675,N_11478,N_11434);
xnor U11676 (N_11676,N_11391,N_11454);
and U11677 (N_11677,N_11378,N_11385);
nor U11678 (N_11678,N_11362,N_11430);
nor U11679 (N_11679,N_11410,N_11371);
xor U11680 (N_11680,N_11579,N_11564);
and U11681 (N_11681,N_11605,N_11656);
nor U11682 (N_11682,N_11647,N_11536);
or U11683 (N_11683,N_11526,N_11664);
xnor U11684 (N_11684,N_11589,N_11658);
and U11685 (N_11685,N_11562,N_11584);
and U11686 (N_11686,N_11637,N_11549);
nor U11687 (N_11687,N_11672,N_11677);
nor U11688 (N_11688,N_11555,N_11648);
xnor U11689 (N_11689,N_11546,N_11551);
xnor U11690 (N_11690,N_11643,N_11569);
and U11691 (N_11691,N_11548,N_11652);
nand U11692 (N_11692,N_11626,N_11570);
and U11693 (N_11693,N_11642,N_11523);
xnor U11694 (N_11694,N_11678,N_11629);
nand U11695 (N_11695,N_11611,N_11668);
and U11696 (N_11696,N_11657,N_11665);
nor U11697 (N_11697,N_11630,N_11571);
and U11698 (N_11698,N_11527,N_11674);
nor U11699 (N_11699,N_11604,N_11640);
or U11700 (N_11700,N_11635,N_11596);
xnor U11701 (N_11701,N_11618,N_11659);
nand U11702 (N_11702,N_11653,N_11651);
nor U11703 (N_11703,N_11554,N_11610);
xor U11704 (N_11704,N_11671,N_11561);
nor U11705 (N_11705,N_11619,N_11560);
nand U11706 (N_11706,N_11661,N_11603);
xnor U11707 (N_11707,N_11633,N_11645);
or U11708 (N_11708,N_11631,N_11616);
or U11709 (N_11709,N_11607,N_11593);
nand U11710 (N_11710,N_11534,N_11552);
xnor U11711 (N_11711,N_11634,N_11575);
xor U11712 (N_11712,N_11553,N_11639);
nor U11713 (N_11713,N_11537,N_11543);
xnor U11714 (N_11714,N_11675,N_11595);
and U11715 (N_11715,N_11614,N_11565);
nor U11716 (N_11716,N_11583,N_11559);
nand U11717 (N_11717,N_11567,N_11649);
nor U11718 (N_11718,N_11623,N_11542);
nor U11719 (N_11719,N_11606,N_11663);
nor U11720 (N_11720,N_11679,N_11524);
xnor U11721 (N_11721,N_11625,N_11620);
xor U11722 (N_11722,N_11590,N_11621);
or U11723 (N_11723,N_11545,N_11597);
nand U11724 (N_11724,N_11550,N_11577);
xor U11725 (N_11725,N_11608,N_11572);
nor U11726 (N_11726,N_11521,N_11573);
xnor U11727 (N_11727,N_11588,N_11609);
and U11728 (N_11728,N_11615,N_11528);
nor U11729 (N_11729,N_11641,N_11632);
or U11730 (N_11730,N_11628,N_11585);
and U11731 (N_11731,N_11594,N_11592);
nor U11732 (N_11732,N_11578,N_11676);
nor U11733 (N_11733,N_11587,N_11522);
nand U11734 (N_11734,N_11581,N_11644);
or U11735 (N_11735,N_11580,N_11636);
nand U11736 (N_11736,N_11612,N_11539);
nand U11737 (N_11737,N_11638,N_11624);
nor U11738 (N_11738,N_11673,N_11667);
xor U11739 (N_11739,N_11654,N_11655);
and U11740 (N_11740,N_11582,N_11541);
xnor U11741 (N_11741,N_11576,N_11669);
and U11742 (N_11742,N_11556,N_11650);
xor U11743 (N_11743,N_11627,N_11613);
or U11744 (N_11744,N_11602,N_11533);
and U11745 (N_11745,N_11600,N_11520);
and U11746 (N_11746,N_11563,N_11662);
nand U11747 (N_11747,N_11586,N_11617);
xor U11748 (N_11748,N_11574,N_11660);
or U11749 (N_11749,N_11538,N_11532);
or U11750 (N_11750,N_11622,N_11568);
xor U11751 (N_11751,N_11531,N_11535);
xor U11752 (N_11752,N_11599,N_11547);
or U11753 (N_11753,N_11529,N_11566);
and U11754 (N_11754,N_11557,N_11530);
and U11755 (N_11755,N_11601,N_11670);
nand U11756 (N_11756,N_11525,N_11646);
and U11757 (N_11757,N_11598,N_11558);
or U11758 (N_11758,N_11666,N_11544);
nor U11759 (N_11759,N_11591,N_11540);
xor U11760 (N_11760,N_11578,N_11616);
nor U11761 (N_11761,N_11570,N_11627);
and U11762 (N_11762,N_11620,N_11594);
and U11763 (N_11763,N_11552,N_11632);
and U11764 (N_11764,N_11604,N_11607);
xor U11765 (N_11765,N_11641,N_11642);
nor U11766 (N_11766,N_11546,N_11527);
nor U11767 (N_11767,N_11541,N_11569);
or U11768 (N_11768,N_11588,N_11603);
and U11769 (N_11769,N_11644,N_11627);
nand U11770 (N_11770,N_11619,N_11646);
nand U11771 (N_11771,N_11663,N_11602);
or U11772 (N_11772,N_11562,N_11528);
nor U11773 (N_11773,N_11581,N_11605);
and U11774 (N_11774,N_11643,N_11545);
or U11775 (N_11775,N_11595,N_11622);
nor U11776 (N_11776,N_11602,N_11646);
nor U11777 (N_11777,N_11526,N_11559);
nor U11778 (N_11778,N_11585,N_11654);
nand U11779 (N_11779,N_11520,N_11545);
and U11780 (N_11780,N_11593,N_11553);
nand U11781 (N_11781,N_11677,N_11598);
xnor U11782 (N_11782,N_11630,N_11651);
or U11783 (N_11783,N_11574,N_11532);
nor U11784 (N_11784,N_11544,N_11577);
nand U11785 (N_11785,N_11555,N_11549);
and U11786 (N_11786,N_11556,N_11581);
or U11787 (N_11787,N_11584,N_11574);
or U11788 (N_11788,N_11642,N_11598);
and U11789 (N_11789,N_11558,N_11589);
and U11790 (N_11790,N_11662,N_11638);
xor U11791 (N_11791,N_11539,N_11566);
nand U11792 (N_11792,N_11660,N_11617);
xor U11793 (N_11793,N_11661,N_11551);
xnor U11794 (N_11794,N_11622,N_11545);
and U11795 (N_11795,N_11530,N_11659);
nand U11796 (N_11796,N_11662,N_11668);
or U11797 (N_11797,N_11597,N_11539);
nand U11798 (N_11798,N_11668,N_11570);
or U11799 (N_11799,N_11573,N_11556);
xor U11800 (N_11800,N_11555,N_11561);
xnor U11801 (N_11801,N_11675,N_11573);
nand U11802 (N_11802,N_11627,N_11548);
nand U11803 (N_11803,N_11526,N_11637);
and U11804 (N_11804,N_11571,N_11659);
nor U11805 (N_11805,N_11588,N_11524);
nand U11806 (N_11806,N_11546,N_11584);
xnor U11807 (N_11807,N_11649,N_11553);
or U11808 (N_11808,N_11564,N_11576);
or U11809 (N_11809,N_11578,N_11634);
nand U11810 (N_11810,N_11535,N_11592);
and U11811 (N_11811,N_11670,N_11529);
and U11812 (N_11812,N_11541,N_11678);
nand U11813 (N_11813,N_11619,N_11550);
nor U11814 (N_11814,N_11614,N_11645);
nand U11815 (N_11815,N_11631,N_11537);
nand U11816 (N_11816,N_11601,N_11662);
and U11817 (N_11817,N_11626,N_11606);
and U11818 (N_11818,N_11619,N_11623);
xor U11819 (N_11819,N_11568,N_11585);
nand U11820 (N_11820,N_11649,N_11620);
or U11821 (N_11821,N_11574,N_11669);
xor U11822 (N_11822,N_11539,N_11649);
xnor U11823 (N_11823,N_11667,N_11610);
nand U11824 (N_11824,N_11564,N_11596);
or U11825 (N_11825,N_11581,N_11627);
and U11826 (N_11826,N_11606,N_11547);
and U11827 (N_11827,N_11549,N_11677);
nor U11828 (N_11828,N_11592,N_11639);
xor U11829 (N_11829,N_11676,N_11543);
nor U11830 (N_11830,N_11572,N_11581);
nand U11831 (N_11831,N_11583,N_11551);
nor U11832 (N_11832,N_11623,N_11538);
nor U11833 (N_11833,N_11590,N_11667);
nand U11834 (N_11834,N_11619,N_11570);
xnor U11835 (N_11835,N_11607,N_11531);
or U11836 (N_11836,N_11585,N_11552);
and U11837 (N_11837,N_11563,N_11553);
or U11838 (N_11838,N_11586,N_11606);
xor U11839 (N_11839,N_11523,N_11568);
nor U11840 (N_11840,N_11690,N_11683);
or U11841 (N_11841,N_11703,N_11775);
and U11842 (N_11842,N_11780,N_11720);
or U11843 (N_11843,N_11810,N_11697);
and U11844 (N_11844,N_11808,N_11693);
and U11845 (N_11845,N_11816,N_11832);
xnor U11846 (N_11846,N_11730,N_11751);
or U11847 (N_11847,N_11798,N_11826);
or U11848 (N_11848,N_11709,N_11834);
and U11849 (N_11849,N_11820,N_11839);
nand U11850 (N_11850,N_11721,N_11795);
or U11851 (N_11851,N_11803,N_11745);
nand U11852 (N_11852,N_11755,N_11728);
xor U11853 (N_11853,N_11778,N_11747);
xnor U11854 (N_11854,N_11764,N_11696);
xor U11855 (N_11855,N_11726,N_11699);
nand U11856 (N_11856,N_11741,N_11701);
nand U11857 (N_11857,N_11742,N_11811);
nor U11858 (N_11858,N_11744,N_11794);
or U11859 (N_11859,N_11765,N_11743);
nand U11860 (N_11860,N_11753,N_11799);
or U11861 (N_11861,N_11768,N_11823);
nand U11862 (N_11862,N_11783,N_11700);
nand U11863 (N_11863,N_11817,N_11707);
and U11864 (N_11864,N_11788,N_11824);
nor U11865 (N_11865,N_11702,N_11757);
nor U11866 (N_11866,N_11695,N_11711);
or U11867 (N_11867,N_11722,N_11784);
and U11868 (N_11868,N_11772,N_11828);
and U11869 (N_11869,N_11705,N_11756);
and U11870 (N_11870,N_11719,N_11710);
nor U11871 (N_11871,N_11750,N_11681);
or U11872 (N_11872,N_11797,N_11807);
xor U11873 (N_11873,N_11727,N_11774);
xor U11874 (N_11874,N_11689,N_11831);
nand U11875 (N_11875,N_11773,N_11746);
and U11876 (N_11876,N_11793,N_11818);
xor U11877 (N_11877,N_11754,N_11680);
or U11878 (N_11878,N_11776,N_11740);
nor U11879 (N_11879,N_11724,N_11806);
and U11880 (N_11880,N_11713,N_11825);
and U11881 (N_11881,N_11805,N_11704);
and U11882 (N_11882,N_11830,N_11682);
xnor U11883 (N_11883,N_11769,N_11827);
and U11884 (N_11884,N_11833,N_11706);
or U11885 (N_11885,N_11761,N_11759);
nand U11886 (N_11886,N_11800,N_11725);
nor U11887 (N_11887,N_11716,N_11789);
or U11888 (N_11888,N_11785,N_11767);
nor U11889 (N_11889,N_11692,N_11779);
xor U11890 (N_11890,N_11766,N_11782);
nand U11891 (N_11891,N_11698,N_11685);
and U11892 (N_11892,N_11763,N_11762);
nor U11893 (N_11893,N_11714,N_11758);
nor U11894 (N_11894,N_11687,N_11815);
nor U11895 (N_11895,N_11787,N_11717);
or U11896 (N_11896,N_11708,N_11760);
nand U11897 (N_11897,N_11802,N_11691);
nand U11898 (N_11898,N_11771,N_11790);
or U11899 (N_11899,N_11801,N_11737);
xor U11900 (N_11900,N_11712,N_11781);
nor U11901 (N_11901,N_11770,N_11804);
xor U11902 (N_11902,N_11812,N_11729);
or U11903 (N_11903,N_11735,N_11752);
and U11904 (N_11904,N_11684,N_11686);
nand U11905 (N_11905,N_11777,N_11814);
xnor U11906 (N_11906,N_11723,N_11813);
nor U11907 (N_11907,N_11809,N_11738);
and U11908 (N_11908,N_11715,N_11796);
xor U11909 (N_11909,N_11821,N_11694);
or U11910 (N_11910,N_11748,N_11838);
nor U11911 (N_11911,N_11835,N_11819);
nand U11912 (N_11912,N_11688,N_11731);
and U11913 (N_11913,N_11734,N_11836);
or U11914 (N_11914,N_11739,N_11792);
xor U11915 (N_11915,N_11837,N_11786);
or U11916 (N_11916,N_11822,N_11791);
nand U11917 (N_11917,N_11733,N_11829);
or U11918 (N_11918,N_11749,N_11732);
nand U11919 (N_11919,N_11718,N_11736);
nor U11920 (N_11920,N_11819,N_11696);
or U11921 (N_11921,N_11799,N_11767);
xnor U11922 (N_11922,N_11736,N_11687);
and U11923 (N_11923,N_11783,N_11800);
or U11924 (N_11924,N_11779,N_11687);
nand U11925 (N_11925,N_11826,N_11761);
or U11926 (N_11926,N_11695,N_11738);
and U11927 (N_11927,N_11733,N_11822);
nor U11928 (N_11928,N_11700,N_11769);
or U11929 (N_11929,N_11772,N_11750);
xor U11930 (N_11930,N_11775,N_11835);
or U11931 (N_11931,N_11718,N_11738);
xnor U11932 (N_11932,N_11801,N_11791);
nor U11933 (N_11933,N_11682,N_11804);
nand U11934 (N_11934,N_11767,N_11694);
and U11935 (N_11935,N_11799,N_11805);
or U11936 (N_11936,N_11694,N_11725);
or U11937 (N_11937,N_11717,N_11786);
and U11938 (N_11938,N_11741,N_11772);
or U11939 (N_11939,N_11682,N_11706);
or U11940 (N_11940,N_11803,N_11705);
nand U11941 (N_11941,N_11680,N_11763);
nand U11942 (N_11942,N_11814,N_11708);
or U11943 (N_11943,N_11838,N_11739);
xor U11944 (N_11944,N_11789,N_11717);
nor U11945 (N_11945,N_11744,N_11779);
xnor U11946 (N_11946,N_11736,N_11815);
nand U11947 (N_11947,N_11811,N_11821);
nor U11948 (N_11948,N_11720,N_11738);
nor U11949 (N_11949,N_11705,N_11680);
or U11950 (N_11950,N_11749,N_11711);
nor U11951 (N_11951,N_11791,N_11826);
xor U11952 (N_11952,N_11737,N_11778);
and U11953 (N_11953,N_11710,N_11750);
or U11954 (N_11954,N_11773,N_11686);
or U11955 (N_11955,N_11742,N_11766);
or U11956 (N_11956,N_11790,N_11780);
or U11957 (N_11957,N_11828,N_11728);
or U11958 (N_11958,N_11833,N_11815);
xor U11959 (N_11959,N_11702,N_11696);
xor U11960 (N_11960,N_11687,N_11698);
nand U11961 (N_11961,N_11737,N_11699);
nand U11962 (N_11962,N_11736,N_11822);
nor U11963 (N_11963,N_11788,N_11772);
nand U11964 (N_11964,N_11795,N_11800);
or U11965 (N_11965,N_11703,N_11755);
and U11966 (N_11966,N_11779,N_11699);
nor U11967 (N_11967,N_11777,N_11701);
xnor U11968 (N_11968,N_11728,N_11775);
nand U11969 (N_11969,N_11802,N_11804);
nand U11970 (N_11970,N_11707,N_11691);
nor U11971 (N_11971,N_11795,N_11824);
nor U11972 (N_11972,N_11784,N_11787);
and U11973 (N_11973,N_11818,N_11729);
xor U11974 (N_11974,N_11711,N_11687);
nand U11975 (N_11975,N_11774,N_11733);
nand U11976 (N_11976,N_11709,N_11787);
or U11977 (N_11977,N_11779,N_11756);
nand U11978 (N_11978,N_11708,N_11721);
nand U11979 (N_11979,N_11720,N_11800);
nor U11980 (N_11980,N_11741,N_11767);
xor U11981 (N_11981,N_11730,N_11688);
nor U11982 (N_11982,N_11722,N_11751);
and U11983 (N_11983,N_11771,N_11698);
or U11984 (N_11984,N_11747,N_11774);
nor U11985 (N_11985,N_11776,N_11833);
and U11986 (N_11986,N_11802,N_11723);
nor U11987 (N_11987,N_11809,N_11761);
nand U11988 (N_11988,N_11838,N_11707);
or U11989 (N_11989,N_11829,N_11832);
xor U11990 (N_11990,N_11770,N_11795);
xor U11991 (N_11991,N_11813,N_11719);
or U11992 (N_11992,N_11688,N_11838);
nand U11993 (N_11993,N_11684,N_11773);
and U11994 (N_11994,N_11746,N_11698);
or U11995 (N_11995,N_11805,N_11695);
nand U11996 (N_11996,N_11768,N_11745);
nand U11997 (N_11997,N_11810,N_11698);
nor U11998 (N_11998,N_11683,N_11756);
nor U11999 (N_11999,N_11715,N_11754);
xnor U12000 (N_12000,N_11919,N_11881);
nand U12001 (N_12001,N_11963,N_11943);
and U12002 (N_12002,N_11849,N_11939);
or U12003 (N_12003,N_11884,N_11955);
or U12004 (N_12004,N_11970,N_11999);
xor U12005 (N_12005,N_11897,N_11941);
nor U12006 (N_12006,N_11893,N_11902);
nand U12007 (N_12007,N_11974,N_11858);
nor U12008 (N_12008,N_11954,N_11910);
nor U12009 (N_12009,N_11985,N_11869);
nand U12010 (N_12010,N_11924,N_11950);
xor U12011 (N_12011,N_11940,N_11867);
and U12012 (N_12012,N_11885,N_11935);
or U12013 (N_12013,N_11853,N_11908);
nor U12014 (N_12014,N_11918,N_11856);
nor U12015 (N_12015,N_11993,N_11952);
nor U12016 (N_12016,N_11972,N_11976);
nand U12017 (N_12017,N_11872,N_11945);
nand U12018 (N_12018,N_11882,N_11862);
nand U12019 (N_12019,N_11937,N_11930);
nand U12020 (N_12020,N_11973,N_11883);
nor U12021 (N_12021,N_11887,N_11863);
nor U12022 (N_12022,N_11942,N_11980);
and U12023 (N_12023,N_11975,N_11953);
or U12024 (N_12024,N_11889,N_11984);
nand U12025 (N_12025,N_11957,N_11964);
xnor U12026 (N_12026,N_11966,N_11944);
nand U12027 (N_12027,N_11923,N_11900);
and U12028 (N_12028,N_11947,N_11852);
nand U12029 (N_12029,N_11979,N_11914);
nand U12030 (N_12030,N_11875,N_11899);
and U12031 (N_12031,N_11895,N_11892);
and U12032 (N_12032,N_11912,N_11840);
nand U12033 (N_12033,N_11842,N_11932);
and U12034 (N_12034,N_11991,N_11846);
nor U12035 (N_12035,N_11988,N_11864);
nor U12036 (N_12036,N_11938,N_11967);
nor U12037 (N_12037,N_11845,N_11956);
nor U12038 (N_12038,N_11989,N_11987);
nand U12039 (N_12039,N_11907,N_11866);
xor U12040 (N_12040,N_11896,N_11934);
or U12041 (N_12041,N_11874,N_11949);
and U12042 (N_12042,N_11871,N_11903);
nand U12043 (N_12043,N_11982,N_11904);
nand U12044 (N_12044,N_11898,N_11848);
and U12045 (N_12045,N_11913,N_11909);
nor U12046 (N_12046,N_11905,N_11946);
xnor U12047 (N_12047,N_11890,N_11994);
or U12048 (N_12048,N_11844,N_11958);
nand U12049 (N_12049,N_11880,N_11977);
xor U12050 (N_12050,N_11917,N_11951);
or U12051 (N_12051,N_11877,N_11873);
nor U12052 (N_12052,N_11841,N_11929);
nand U12053 (N_12053,N_11981,N_11927);
or U12054 (N_12054,N_11901,N_11983);
and U12055 (N_12055,N_11990,N_11855);
and U12056 (N_12056,N_11916,N_11965);
nand U12057 (N_12057,N_11879,N_11948);
nor U12058 (N_12058,N_11978,N_11933);
xnor U12059 (N_12059,N_11996,N_11891);
and U12060 (N_12060,N_11854,N_11921);
nor U12061 (N_12061,N_11878,N_11931);
or U12062 (N_12062,N_11998,N_11857);
xnor U12063 (N_12063,N_11961,N_11886);
nor U12064 (N_12064,N_11959,N_11920);
nand U12065 (N_12065,N_11925,N_11870);
nor U12066 (N_12066,N_11995,N_11865);
nand U12067 (N_12067,N_11915,N_11971);
or U12068 (N_12068,N_11992,N_11859);
xnor U12069 (N_12069,N_11847,N_11936);
or U12070 (N_12070,N_11860,N_11868);
or U12071 (N_12071,N_11906,N_11843);
and U12072 (N_12072,N_11876,N_11926);
nand U12073 (N_12073,N_11861,N_11962);
or U12074 (N_12074,N_11997,N_11986);
xor U12075 (N_12075,N_11969,N_11888);
xnor U12076 (N_12076,N_11960,N_11850);
or U12077 (N_12077,N_11911,N_11851);
nor U12078 (N_12078,N_11922,N_11894);
nor U12079 (N_12079,N_11928,N_11968);
and U12080 (N_12080,N_11927,N_11854);
xnor U12081 (N_12081,N_11952,N_11840);
nor U12082 (N_12082,N_11951,N_11963);
xnor U12083 (N_12083,N_11879,N_11870);
or U12084 (N_12084,N_11970,N_11885);
or U12085 (N_12085,N_11866,N_11992);
nor U12086 (N_12086,N_11847,N_11921);
nand U12087 (N_12087,N_11951,N_11855);
and U12088 (N_12088,N_11932,N_11996);
xor U12089 (N_12089,N_11841,N_11899);
nand U12090 (N_12090,N_11864,N_11948);
or U12091 (N_12091,N_11942,N_11953);
xor U12092 (N_12092,N_11966,N_11876);
nor U12093 (N_12093,N_11974,N_11949);
nor U12094 (N_12094,N_11998,N_11957);
and U12095 (N_12095,N_11932,N_11870);
nor U12096 (N_12096,N_11962,N_11914);
or U12097 (N_12097,N_11875,N_11923);
nand U12098 (N_12098,N_11945,N_11847);
nor U12099 (N_12099,N_11988,N_11977);
xnor U12100 (N_12100,N_11840,N_11996);
nand U12101 (N_12101,N_11934,N_11984);
nand U12102 (N_12102,N_11937,N_11910);
or U12103 (N_12103,N_11889,N_11979);
nand U12104 (N_12104,N_11871,N_11887);
or U12105 (N_12105,N_11859,N_11977);
nor U12106 (N_12106,N_11945,N_11853);
xor U12107 (N_12107,N_11926,N_11872);
nor U12108 (N_12108,N_11898,N_11861);
or U12109 (N_12109,N_11870,N_11991);
xor U12110 (N_12110,N_11876,N_11950);
nor U12111 (N_12111,N_11950,N_11992);
nand U12112 (N_12112,N_11920,N_11994);
nor U12113 (N_12113,N_11868,N_11967);
or U12114 (N_12114,N_11957,N_11853);
and U12115 (N_12115,N_11934,N_11892);
xnor U12116 (N_12116,N_11926,N_11857);
or U12117 (N_12117,N_11958,N_11873);
or U12118 (N_12118,N_11889,N_11897);
and U12119 (N_12119,N_11896,N_11939);
nand U12120 (N_12120,N_11885,N_11983);
and U12121 (N_12121,N_11996,N_11895);
xor U12122 (N_12122,N_11994,N_11906);
and U12123 (N_12123,N_11944,N_11919);
xnor U12124 (N_12124,N_11952,N_11851);
and U12125 (N_12125,N_11873,N_11966);
xnor U12126 (N_12126,N_11943,N_11955);
xnor U12127 (N_12127,N_11933,N_11937);
nand U12128 (N_12128,N_11876,N_11928);
nor U12129 (N_12129,N_11890,N_11850);
and U12130 (N_12130,N_11848,N_11880);
nand U12131 (N_12131,N_11937,N_11868);
or U12132 (N_12132,N_11845,N_11967);
and U12133 (N_12133,N_11876,N_11854);
nor U12134 (N_12134,N_11931,N_11894);
nor U12135 (N_12135,N_11843,N_11983);
nor U12136 (N_12136,N_11991,N_11961);
nand U12137 (N_12137,N_11868,N_11904);
xnor U12138 (N_12138,N_11954,N_11898);
xor U12139 (N_12139,N_11902,N_11860);
xnor U12140 (N_12140,N_11870,N_11923);
or U12141 (N_12141,N_11845,N_11957);
nand U12142 (N_12142,N_11943,N_11884);
or U12143 (N_12143,N_11909,N_11903);
xor U12144 (N_12144,N_11902,N_11945);
and U12145 (N_12145,N_11952,N_11871);
nand U12146 (N_12146,N_11943,N_11996);
nand U12147 (N_12147,N_11861,N_11878);
nor U12148 (N_12148,N_11842,N_11883);
nor U12149 (N_12149,N_11979,N_11988);
xor U12150 (N_12150,N_11930,N_11841);
xor U12151 (N_12151,N_11971,N_11983);
and U12152 (N_12152,N_11954,N_11887);
nand U12153 (N_12153,N_11904,N_11963);
nand U12154 (N_12154,N_11864,N_11961);
and U12155 (N_12155,N_11985,N_11912);
or U12156 (N_12156,N_11903,N_11950);
or U12157 (N_12157,N_11986,N_11951);
nand U12158 (N_12158,N_11873,N_11895);
nor U12159 (N_12159,N_11843,N_11854);
nor U12160 (N_12160,N_12086,N_12035);
nand U12161 (N_12161,N_12047,N_12131);
and U12162 (N_12162,N_12049,N_12121);
xor U12163 (N_12163,N_12120,N_12130);
or U12164 (N_12164,N_12038,N_12122);
and U12165 (N_12165,N_12031,N_12013);
xor U12166 (N_12166,N_12139,N_12071);
xnor U12167 (N_12167,N_12029,N_12081);
or U12168 (N_12168,N_12052,N_12114);
or U12169 (N_12169,N_12152,N_12073);
nor U12170 (N_12170,N_12011,N_12060);
or U12171 (N_12171,N_12144,N_12094);
xnor U12172 (N_12172,N_12063,N_12002);
and U12173 (N_12173,N_12022,N_12075);
nor U12174 (N_12174,N_12111,N_12159);
xor U12175 (N_12175,N_12003,N_12030);
or U12176 (N_12176,N_12040,N_12100);
nor U12177 (N_12177,N_12053,N_12048);
and U12178 (N_12178,N_12024,N_12057);
and U12179 (N_12179,N_12091,N_12090);
and U12180 (N_12180,N_12147,N_12112);
nor U12181 (N_12181,N_12136,N_12001);
and U12182 (N_12182,N_12129,N_12046);
xnor U12183 (N_12183,N_12007,N_12043);
xnor U12184 (N_12184,N_12110,N_12140);
xnor U12185 (N_12185,N_12123,N_12061);
xnor U12186 (N_12186,N_12142,N_12115);
nor U12187 (N_12187,N_12125,N_12074);
nor U12188 (N_12188,N_12021,N_12055);
xnor U12189 (N_12189,N_12085,N_12020);
nor U12190 (N_12190,N_12019,N_12133);
and U12191 (N_12191,N_12016,N_12044);
nand U12192 (N_12192,N_12067,N_12155);
nand U12193 (N_12193,N_12103,N_12072);
nand U12194 (N_12194,N_12156,N_12037);
and U12195 (N_12195,N_12098,N_12143);
nand U12196 (N_12196,N_12033,N_12006);
nor U12197 (N_12197,N_12080,N_12153);
nand U12198 (N_12198,N_12065,N_12045);
nand U12199 (N_12199,N_12004,N_12087);
nor U12200 (N_12200,N_12096,N_12146);
xnor U12201 (N_12201,N_12127,N_12008);
and U12202 (N_12202,N_12124,N_12088);
nand U12203 (N_12203,N_12119,N_12041);
and U12204 (N_12204,N_12066,N_12076);
xor U12205 (N_12205,N_12069,N_12106);
and U12206 (N_12206,N_12104,N_12054);
xor U12207 (N_12207,N_12015,N_12117);
and U12208 (N_12208,N_12032,N_12138);
nor U12209 (N_12209,N_12056,N_12134);
nand U12210 (N_12210,N_12026,N_12089);
xor U12211 (N_12211,N_12034,N_12078);
nor U12212 (N_12212,N_12150,N_12099);
nor U12213 (N_12213,N_12018,N_12107);
xnor U12214 (N_12214,N_12126,N_12102);
nand U12215 (N_12215,N_12009,N_12010);
xor U12216 (N_12216,N_12093,N_12014);
nor U12217 (N_12217,N_12042,N_12051);
or U12218 (N_12218,N_12083,N_12157);
or U12219 (N_12219,N_12023,N_12084);
nor U12220 (N_12220,N_12109,N_12027);
xnor U12221 (N_12221,N_12036,N_12068);
xnor U12222 (N_12222,N_12148,N_12154);
or U12223 (N_12223,N_12132,N_12141);
or U12224 (N_12224,N_12118,N_12058);
or U12225 (N_12225,N_12105,N_12097);
or U12226 (N_12226,N_12050,N_12077);
nor U12227 (N_12227,N_12070,N_12079);
xnor U12228 (N_12228,N_12017,N_12064);
nand U12229 (N_12229,N_12059,N_12082);
nor U12230 (N_12230,N_12113,N_12028);
nand U12231 (N_12231,N_12025,N_12151);
nor U12232 (N_12232,N_12005,N_12128);
nand U12233 (N_12233,N_12158,N_12092);
or U12234 (N_12234,N_12145,N_12135);
xor U12235 (N_12235,N_12000,N_12095);
or U12236 (N_12236,N_12062,N_12116);
xnor U12237 (N_12237,N_12137,N_12012);
nor U12238 (N_12238,N_12108,N_12101);
nor U12239 (N_12239,N_12149,N_12039);
and U12240 (N_12240,N_12070,N_12101);
and U12241 (N_12241,N_12076,N_12111);
and U12242 (N_12242,N_12060,N_12009);
nor U12243 (N_12243,N_12106,N_12016);
nor U12244 (N_12244,N_12114,N_12073);
or U12245 (N_12245,N_12015,N_12112);
and U12246 (N_12246,N_12062,N_12127);
or U12247 (N_12247,N_12089,N_12110);
nand U12248 (N_12248,N_12096,N_12011);
nor U12249 (N_12249,N_12126,N_12131);
xor U12250 (N_12250,N_12103,N_12014);
and U12251 (N_12251,N_12050,N_12107);
xnor U12252 (N_12252,N_12010,N_12007);
xnor U12253 (N_12253,N_12138,N_12103);
and U12254 (N_12254,N_12060,N_12117);
or U12255 (N_12255,N_12128,N_12040);
and U12256 (N_12256,N_12154,N_12106);
nor U12257 (N_12257,N_12097,N_12081);
and U12258 (N_12258,N_12075,N_12027);
xor U12259 (N_12259,N_12033,N_12036);
and U12260 (N_12260,N_12052,N_12039);
and U12261 (N_12261,N_12070,N_12131);
nand U12262 (N_12262,N_12010,N_12069);
or U12263 (N_12263,N_12012,N_12068);
nand U12264 (N_12264,N_12072,N_12086);
xnor U12265 (N_12265,N_12003,N_12066);
or U12266 (N_12266,N_12118,N_12088);
or U12267 (N_12267,N_12025,N_12131);
or U12268 (N_12268,N_12121,N_12037);
nand U12269 (N_12269,N_12158,N_12105);
nor U12270 (N_12270,N_12115,N_12042);
or U12271 (N_12271,N_12088,N_12109);
xor U12272 (N_12272,N_12021,N_12156);
and U12273 (N_12273,N_12117,N_12039);
nor U12274 (N_12274,N_12158,N_12069);
or U12275 (N_12275,N_12046,N_12081);
nand U12276 (N_12276,N_12148,N_12080);
or U12277 (N_12277,N_12087,N_12056);
xor U12278 (N_12278,N_12042,N_12126);
nor U12279 (N_12279,N_12148,N_12036);
xnor U12280 (N_12280,N_12130,N_12037);
xor U12281 (N_12281,N_12093,N_12003);
or U12282 (N_12282,N_12092,N_12021);
nor U12283 (N_12283,N_12036,N_12046);
or U12284 (N_12284,N_12101,N_12038);
nor U12285 (N_12285,N_12081,N_12035);
nor U12286 (N_12286,N_12153,N_12044);
and U12287 (N_12287,N_12060,N_12129);
xor U12288 (N_12288,N_12077,N_12114);
nor U12289 (N_12289,N_12009,N_12058);
xor U12290 (N_12290,N_12138,N_12159);
or U12291 (N_12291,N_12135,N_12120);
nand U12292 (N_12292,N_12150,N_12055);
xnor U12293 (N_12293,N_12037,N_12066);
nor U12294 (N_12294,N_12159,N_12093);
nand U12295 (N_12295,N_12071,N_12049);
nor U12296 (N_12296,N_12048,N_12129);
nand U12297 (N_12297,N_12122,N_12063);
or U12298 (N_12298,N_12126,N_12019);
nand U12299 (N_12299,N_12084,N_12082);
xnor U12300 (N_12300,N_12117,N_12051);
or U12301 (N_12301,N_12152,N_12037);
nor U12302 (N_12302,N_12109,N_12159);
nor U12303 (N_12303,N_12091,N_12139);
and U12304 (N_12304,N_12101,N_12017);
nor U12305 (N_12305,N_12029,N_12136);
nand U12306 (N_12306,N_12141,N_12000);
or U12307 (N_12307,N_12010,N_12076);
xor U12308 (N_12308,N_12113,N_12002);
or U12309 (N_12309,N_12120,N_12145);
nor U12310 (N_12310,N_12156,N_12082);
xnor U12311 (N_12311,N_12051,N_12070);
and U12312 (N_12312,N_12117,N_12076);
and U12313 (N_12313,N_12010,N_12060);
nor U12314 (N_12314,N_12042,N_12095);
nor U12315 (N_12315,N_12099,N_12067);
and U12316 (N_12316,N_12111,N_12149);
and U12317 (N_12317,N_12060,N_12105);
or U12318 (N_12318,N_12068,N_12096);
nand U12319 (N_12319,N_12032,N_12102);
nor U12320 (N_12320,N_12231,N_12305);
and U12321 (N_12321,N_12246,N_12255);
or U12322 (N_12322,N_12276,N_12248);
nor U12323 (N_12323,N_12295,N_12259);
nor U12324 (N_12324,N_12256,N_12173);
nor U12325 (N_12325,N_12217,N_12170);
xnor U12326 (N_12326,N_12313,N_12279);
nor U12327 (N_12327,N_12281,N_12241);
xor U12328 (N_12328,N_12280,N_12219);
xnor U12329 (N_12329,N_12273,N_12227);
or U12330 (N_12330,N_12267,N_12202);
or U12331 (N_12331,N_12270,N_12167);
and U12332 (N_12332,N_12300,N_12196);
xor U12333 (N_12333,N_12315,N_12229);
and U12334 (N_12334,N_12260,N_12211);
xor U12335 (N_12335,N_12275,N_12171);
nand U12336 (N_12336,N_12177,N_12232);
nor U12337 (N_12337,N_12191,N_12181);
xor U12338 (N_12338,N_12206,N_12296);
xor U12339 (N_12339,N_12309,N_12292);
and U12340 (N_12340,N_12164,N_12258);
xnor U12341 (N_12341,N_12249,N_12168);
xnor U12342 (N_12342,N_12200,N_12286);
nor U12343 (N_12343,N_12180,N_12314);
nand U12344 (N_12344,N_12183,N_12230);
xnor U12345 (N_12345,N_12182,N_12185);
and U12346 (N_12346,N_12222,N_12287);
nand U12347 (N_12347,N_12175,N_12221);
xor U12348 (N_12348,N_12186,N_12274);
xnor U12349 (N_12349,N_12162,N_12224);
and U12350 (N_12350,N_12238,N_12318);
or U12351 (N_12351,N_12311,N_12242);
and U12352 (N_12352,N_12178,N_12223);
and U12353 (N_12353,N_12236,N_12294);
or U12354 (N_12354,N_12262,N_12207);
xor U12355 (N_12355,N_12301,N_12165);
xnor U12356 (N_12356,N_12205,N_12298);
xnor U12357 (N_12357,N_12306,N_12233);
or U12358 (N_12358,N_12188,N_12302);
or U12359 (N_12359,N_12297,N_12316);
xor U12360 (N_12360,N_12247,N_12197);
nand U12361 (N_12361,N_12278,N_12269);
or U12362 (N_12362,N_12289,N_12216);
xnor U12363 (N_12363,N_12271,N_12198);
xnor U12364 (N_12364,N_12199,N_12214);
and U12365 (N_12365,N_12293,N_12254);
nor U12366 (N_12366,N_12209,N_12245);
and U12367 (N_12367,N_12250,N_12203);
and U12368 (N_12368,N_12303,N_12237);
or U12369 (N_12369,N_12174,N_12253);
and U12370 (N_12370,N_12261,N_12252);
nand U12371 (N_12371,N_12218,N_12304);
nand U12372 (N_12372,N_12290,N_12194);
or U12373 (N_12373,N_12277,N_12235);
and U12374 (N_12374,N_12251,N_12166);
nor U12375 (N_12375,N_12208,N_12244);
or U12376 (N_12376,N_12213,N_12282);
or U12377 (N_12377,N_12257,N_12263);
nor U12378 (N_12378,N_12226,N_12299);
or U12379 (N_12379,N_12319,N_12310);
nand U12380 (N_12380,N_12169,N_12243);
nor U12381 (N_12381,N_12239,N_12193);
or U12382 (N_12382,N_12283,N_12220);
or U12383 (N_12383,N_12161,N_12266);
nor U12384 (N_12384,N_12176,N_12272);
nand U12385 (N_12385,N_12264,N_12184);
nor U12386 (N_12386,N_12288,N_12228);
or U12387 (N_12387,N_12210,N_12172);
nand U12388 (N_12388,N_12225,N_12179);
nand U12389 (N_12389,N_12268,N_12312);
and U12390 (N_12390,N_12201,N_12160);
and U12391 (N_12391,N_12212,N_12215);
and U12392 (N_12392,N_12189,N_12308);
nand U12393 (N_12393,N_12265,N_12234);
xor U12394 (N_12394,N_12291,N_12240);
and U12395 (N_12395,N_12187,N_12317);
nand U12396 (N_12396,N_12285,N_12190);
or U12397 (N_12397,N_12195,N_12204);
nor U12398 (N_12398,N_12192,N_12307);
or U12399 (N_12399,N_12163,N_12284);
nor U12400 (N_12400,N_12274,N_12196);
nand U12401 (N_12401,N_12261,N_12193);
or U12402 (N_12402,N_12279,N_12160);
nor U12403 (N_12403,N_12268,N_12187);
and U12404 (N_12404,N_12250,N_12223);
or U12405 (N_12405,N_12213,N_12290);
xnor U12406 (N_12406,N_12217,N_12239);
or U12407 (N_12407,N_12167,N_12282);
and U12408 (N_12408,N_12212,N_12181);
nor U12409 (N_12409,N_12271,N_12204);
or U12410 (N_12410,N_12244,N_12188);
nor U12411 (N_12411,N_12234,N_12270);
or U12412 (N_12412,N_12276,N_12318);
nand U12413 (N_12413,N_12253,N_12173);
or U12414 (N_12414,N_12175,N_12213);
or U12415 (N_12415,N_12221,N_12176);
or U12416 (N_12416,N_12214,N_12262);
or U12417 (N_12417,N_12220,N_12178);
nand U12418 (N_12418,N_12288,N_12285);
or U12419 (N_12419,N_12302,N_12213);
nor U12420 (N_12420,N_12189,N_12213);
or U12421 (N_12421,N_12211,N_12247);
xor U12422 (N_12422,N_12245,N_12234);
xnor U12423 (N_12423,N_12318,N_12312);
and U12424 (N_12424,N_12193,N_12191);
or U12425 (N_12425,N_12280,N_12314);
nor U12426 (N_12426,N_12282,N_12231);
or U12427 (N_12427,N_12215,N_12226);
nor U12428 (N_12428,N_12278,N_12232);
and U12429 (N_12429,N_12218,N_12290);
and U12430 (N_12430,N_12281,N_12269);
and U12431 (N_12431,N_12202,N_12255);
or U12432 (N_12432,N_12295,N_12190);
nand U12433 (N_12433,N_12306,N_12240);
xor U12434 (N_12434,N_12216,N_12199);
nor U12435 (N_12435,N_12271,N_12257);
xor U12436 (N_12436,N_12290,N_12293);
or U12437 (N_12437,N_12285,N_12304);
and U12438 (N_12438,N_12284,N_12233);
xor U12439 (N_12439,N_12191,N_12245);
nand U12440 (N_12440,N_12194,N_12256);
nor U12441 (N_12441,N_12267,N_12188);
xor U12442 (N_12442,N_12225,N_12274);
nor U12443 (N_12443,N_12255,N_12180);
nand U12444 (N_12444,N_12212,N_12200);
and U12445 (N_12445,N_12309,N_12207);
nand U12446 (N_12446,N_12216,N_12273);
and U12447 (N_12447,N_12305,N_12220);
nor U12448 (N_12448,N_12285,N_12161);
and U12449 (N_12449,N_12265,N_12252);
or U12450 (N_12450,N_12187,N_12209);
xnor U12451 (N_12451,N_12206,N_12233);
nand U12452 (N_12452,N_12286,N_12166);
nor U12453 (N_12453,N_12259,N_12270);
xnor U12454 (N_12454,N_12217,N_12318);
nand U12455 (N_12455,N_12169,N_12285);
xor U12456 (N_12456,N_12177,N_12240);
xnor U12457 (N_12457,N_12255,N_12162);
nand U12458 (N_12458,N_12193,N_12287);
or U12459 (N_12459,N_12215,N_12218);
or U12460 (N_12460,N_12312,N_12195);
and U12461 (N_12461,N_12166,N_12202);
nand U12462 (N_12462,N_12231,N_12190);
nand U12463 (N_12463,N_12208,N_12313);
or U12464 (N_12464,N_12212,N_12174);
and U12465 (N_12465,N_12293,N_12267);
or U12466 (N_12466,N_12270,N_12276);
and U12467 (N_12467,N_12294,N_12263);
or U12468 (N_12468,N_12300,N_12166);
and U12469 (N_12469,N_12281,N_12294);
and U12470 (N_12470,N_12217,N_12242);
xnor U12471 (N_12471,N_12229,N_12269);
nor U12472 (N_12472,N_12197,N_12227);
nor U12473 (N_12473,N_12319,N_12259);
or U12474 (N_12474,N_12278,N_12170);
nor U12475 (N_12475,N_12229,N_12205);
or U12476 (N_12476,N_12319,N_12266);
nor U12477 (N_12477,N_12230,N_12270);
and U12478 (N_12478,N_12290,N_12284);
and U12479 (N_12479,N_12279,N_12268);
xor U12480 (N_12480,N_12456,N_12358);
xnor U12481 (N_12481,N_12376,N_12425);
or U12482 (N_12482,N_12459,N_12477);
nand U12483 (N_12483,N_12475,N_12443);
nor U12484 (N_12484,N_12328,N_12372);
nand U12485 (N_12485,N_12397,N_12402);
or U12486 (N_12486,N_12360,N_12453);
nor U12487 (N_12487,N_12466,N_12342);
nand U12488 (N_12488,N_12463,N_12321);
nand U12489 (N_12489,N_12324,N_12359);
nand U12490 (N_12490,N_12391,N_12355);
or U12491 (N_12491,N_12384,N_12447);
or U12492 (N_12492,N_12353,N_12411);
nor U12493 (N_12493,N_12435,N_12418);
nor U12494 (N_12494,N_12464,N_12472);
xnor U12495 (N_12495,N_12406,N_12415);
xnor U12496 (N_12496,N_12437,N_12461);
nand U12497 (N_12497,N_12420,N_12403);
and U12498 (N_12498,N_12362,N_12326);
and U12499 (N_12499,N_12433,N_12338);
nand U12500 (N_12500,N_12454,N_12450);
nor U12501 (N_12501,N_12408,N_12457);
nand U12502 (N_12502,N_12331,N_12323);
and U12503 (N_12503,N_12439,N_12381);
xnor U12504 (N_12504,N_12400,N_12401);
nand U12505 (N_12505,N_12465,N_12413);
and U12506 (N_12506,N_12394,N_12399);
and U12507 (N_12507,N_12366,N_12458);
nand U12508 (N_12508,N_12478,N_12462);
xor U12509 (N_12509,N_12417,N_12377);
xor U12510 (N_12510,N_12373,N_12452);
or U12511 (N_12511,N_12378,N_12455);
or U12512 (N_12512,N_12379,N_12442);
nand U12513 (N_12513,N_12410,N_12333);
nand U12514 (N_12514,N_12392,N_12339);
or U12515 (N_12515,N_12441,N_12448);
or U12516 (N_12516,N_12395,N_12354);
nor U12517 (N_12517,N_12389,N_12347);
or U12518 (N_12518,N_12430,N_12361);
xnor U12519 (N_12519,N_12421,N_12468);
and U12520 (N_12520,N_12369,N_12367);
or U12521 (N_12521,N_12404,N_12346);
nor U12522 (N_12522,N_12387,N_12329);
or U12523 (N_12523,N_12340,N_12446);
xor U12524 (N_12524,N_12336,N_12335);
nor U12525 (N_12525,N_12344,N_12393);
xnor U12526 (N_12526,N_12390,N_12436);
nand U12527 (N_12527,N_12434,N_12325);
nor U12528 (N_12528,N_12451,N_12382);
or U12529 (N_12529,N_12467,N_12423);
nand U12530 (N_12530,N_12380,N_12405);
or U12531 (N_12531,N_12473,N_12334);
xor U12532 (N_12532,N_12352,N_12445);
and U12533 (N_12533,N_12368,N_12460);
xor U12534 (N_12534,N_12357,N_12426);
nand U12535 (N_12535,N_12419,N_12471);
nor U12536 (N_12536,N_12412,N_12383);
nor U12537 (N_12537,N_12337,N_12327);
nand U12538 (N_12538,N_12385,N_12374);
xor U12539 (N_12539,N_12427,N_12440);
xor U12540 (N_12540,N_12375,N_12438);
and U12541 (N_12541,N_12414,N_12388);
or U12542 (N_12542,N_12429,N_12469);
or U12543 (N_12543,N_12363,N_12474);
nor U12544 (N_12544,N_12332,N_12386);
xnor U12545 (N_12545,N_12476,N_12345);
or U12546 (N_12546,N_12351,N_12349);
and U12547 (N_12547,N_12364,N_12444);
or U12548 (N_12548,N_12479,N_12416);
xnor U12549 (N_12549,N_12449,N_12356);
and U12550 (N_12550,N_12432,N_12396);
xnor U12551 (N_12551,N_12370,N_12428);
and U12552 (N_12552,N_12350,N_12424);
nand U12553 (N_12553,N_12470,N_12348);
nor U12554 (N_12554,N_12398,N_12320);
nor U12555 (N_12555,N_12330,N_12409);
and U12556 (N_12556,N_12407,N_12365);
xnor U12557 (N_12557,N_12371,N_12343);
xnor U12558 (N_12558,N_12341,N_12431);
and U12559 (N_12559,N_12322,N_12422);
nand U12560 (N_12560,N_12470,N_12415);
nand U12561 (N_12561,N_12366,N_12378);
or U12562 (N_12562,N_12388,N_12403);
or U12563 (N_12563,N_12411,N_12324);
nand U12564 (N_12564,N_12428,N_12453);
or U12565 (N_12565,N_12383,N_12422);
xor U12566 (N_12566,N_12373,N_12400);
and U12567 (N_12567,N_12453,N_12367);
or U12568 (N_12568,N_12443,N_12423);
nand U12569 (N_12569,N_12328,N_12392);
nand U12570 (N_12570,N_12357,N_12331);
xor U12571 (N_12571,N_12414,N_12439);
or U12572 (N_12572,N_12378,N_12371);
nand U12573 (N_12573,N_12369,N_12476);
nand U12574 (N_12574,N_12439,N_12462);
nor U12575 (N_12575,N_12348,N_12329);
and U12576 (N_12576,N_12442,N_12413);
nor U12577 (N_12577,N_12338,N_12340);
nor U12578 (N_12578,N_12384,N_12429);
and U12579 (N_12579,N_12421,N_12426);
or U12580 (N_12580,N_12334,N_12394);
and U12581 (N_12581,N_12378,N_12343);
nor U12582 (N_12582,N_12393,N_12389);
nor U12583 (N_12583,N_12414,N_12456);
nand U12584 (N_12584,N_12359,N_12450);
or U12585 (N_12585,N_12434,N_12431);
nand U12586 (N_12586,N_12408,N_12353);
xor U12587 (N_12587,N_12397,N_12394);
xnor U12588 (N_12588,N_12414,N_12360);
or U12589 (N_12589,N_12396,N_12328);
xnor U12590 (N_12590,N_12459,N_12424);
or U12591 (N_12591,N_12343,N_12413);
and U12592 (N_12592,N_12440,N_12394);
and U12593 (N_12593,N_12342,N_12429);
or U12594 (N_12594,N_12419,N_12475);
or U12595 (N_12595,N_12370,N_12408);
nor U12596 (N_12596,N_12408,N_12410);
nor U12597 (N_12597,N_12339,N_12473);
xor U12598 (N_12598,N_12334,N_12401);
nor U12599 (N_12599,N_12429,N_12435);
or U12600 (N_12600,N_12426,N_12373);
nor U12601 (N_12601,N_12456,N_12357);
nand U12602 (N_12602,N_12325,N_12457);
and U12603 (N_12603,N_12350,N_12469);
or U12604 (N_12604,N_12425,N_12336);
and U12605 (N_12605,N_12440,N_12449);
nor U12606 (N_12606,N_12343,N_12324);
or U12607 (N_12607,N_12339,N_12406);
or U12608 (N_12608,N_12441,N_12427);
or U12609 (N_12609,N_12406,N_12380);
nand U12610 (N_12610,N_12402,N_12351);
nand U12611 (N_12611,N_12443,N_12322);
or U12612 (N_12612,N_12397,N_12449);
nand U12613 (N_12613,N_12344,N_12322);
or U12614 (N_12614,N_12449,N_12399);
or U12615 (N_12615,N_12414,N_12356);
nor U12616 (N_12616,N_12432,N_12463);
or U12617 (N_12617,N_12459,N_12343);
or U12618 (N_12618,N_12462,N_12389);
and U12619 (N_12619,N_12436,N_12355);
nand U12620 (N_12620,N_12334,N_12398);
nand U12621 (N_12621,N_12477,N_12385);
nand U12622 (N_12622,N_12402,N_12360);
xor U12623 (N_12623,N_12332,N_12459);
xor U12624 (N_12624,N_12383,N_12370);
nor U12625 (N_12625,N_12367,N_12476);
and U12626 (N_12626,N_12446,N_12457);
nand U12627 (N_12627,N_12398,N_12339);
nand U12628 (N_12628,N_12328,N_12420);
nor U12629 (N_12629,N_12376,N_12397);
and U12630 (N_12630,N_12449,N_12320);
nor U12631 (N_12631,N_12400,N_12464);
xnor U12632 (N_12632,N_12356,N_12334);
nor U12633 (N_12633,N_12463,N_12361);
and U12634 (N_12634,N_12348,N_12345);
xnor U12635 (N_12635,N_12330,N_12465);
or U12636 (N_12636,N_12477,N_12327);
and U12637 (N_12637,N_12454,N_12455);
nor U12638 (N_12638,N_12360,N_12340);
nand U12639 (N_12639,N_12427,N_12324);
nor U12640 (N_12640,N_12503,N_12580);
and U12641 (N_12641,N_12540,N_12552);
nor U12642 (N_12642,N_12636,N_12592);
nand U12643 (N_12643,N_12551,N_12511);
and U12644 (N_12644,N_12595,N_12598);
and U12645 (N_12645,N_12597,N_12624);
and U12646 (N_12646,N_12618,N_12589);
and U12647 (N_12647,N_12559,N_12521);
or U12648 (N_12648,N_12531,N_12532);
nor U12649 (N_12649,N_12523,N_12575);
nor U12650 (N_12650,N_12518,N_12558);
and U12651 (N_12651,N_12554,N_12534);
nand U12652 (N_12652,N_12601,N_12520);
and U12653 (N_12653,N_12494,N_12612);
xor U12654 (N_12654,N_12508,N_12538);
and U12655 (N_12655,N_12505,N_12553);
nor U12656 (N_12656,N_12504,N_12615);
xnor U12657 (N_12657,N_12513,N_12610);
xnor U12658 (N_12658,N_12555,N_12510);
xor U12659 (N_12659,N_12500,N_12544);
and U12660 (N_12660,N_12560,N_12635);
xnor U12661 (N_12661,N_12509,N_12539);
xnor U12662 (N_12662,N_12585,N_12578);
and U12663 (N_12663,N_12491,N_12495);
xnor U12664 (N_12664,N_12625,N_12634);
xor U12665 (N_12665,N_12614,N_12501);
nand U12666 (N_12666,N_12527,N_12608);
nand U12667 (N_12667,N_12631,N_12633);
xor U12668 (N_12668,N_12543,N_12564);
or U12669 (N_12669,N_12599,N_12571);
or U12670 (N_12670,N_12567,N_12570);
and U12671 (N_12671,N_12481,N_12547);
nor U12672 (N_12672,N_12581,N_12621);
nor U12673 (N_12673,N_12561,N_12506);
nor U12674 (N_12674,N_12619,N_12632);
xnor U12675 (N_12675,N_12548,N_12576);
or U12676 (N_12676,N_12622,N_12535);
nand U12677 (N_12677,N_12620,N_12623);
nand U12678 (N_12678,N_12573,N_12587);
nor U12679 (N_12679,N_12613,N_12603);
xnor U12680 (N_12680,N_12566,N_12512);
xor U12681 (N_12681,N_12606,N_12563);
or U12682 (N_12682,N_12528,N_12591);
nor U12683 (N_12683,N_12630,N_12515);
or U12684 (N_12684,N_12607,N_12556);
xnor U12685 (N_12685,N_12482,N_12583);
nand U12686 (N_12686,N_12568,N_12577);
nor U12687 (N_12687,N_12499,N_12529);
or U12688 (N_12688,N_12516,N_12498);
or U12689 (N_12689,N_12617,N_12545);
nand U12690 (N_12690,N_12569,N_12492);
and U12691 (N_12691,N_12483,N_12557);
xor U12692 (N_12692,N_12605,N_12480);
nor U12693 (N_12693,N_12550,N_12594);
nor U12694 (N_12694,N_12637,N_12488);
nor U12695 (N_12695,N_12486,N_12507);
or U12696 (N_12696,N_12562,N_12639);
nand U12697 (N_12697,N_12530,N_12522);
nor U12698 (N_12698,N_12541,N_12593);
xnor U12699 (N_12699,N_12590,N_12524);
nand U12700 (N_12700,N_12616,N_12604);
nand U12701 (N_12701,N_12537,N_12497);
and U12702 (N_12702,N_12586,N_12493);
and U12703 (N_12703,N_12542,N_12517);
nand U12704 (N_12704,N_12602,N_12629);
and U12705 (N_12705,N_12549,N_12609);
xor U12706 (N_12706,N_12490,N_12514);
nand U12707 (N_12707,N_12536,N_12489);
nand U12708 (N_12708,N_12638,N_12582);
or U12709 (N_12709,N_12626,N_12584);
nor U12710 (N_12710,N_12579,N_12519);
nor U12711 (N_12711,N_12496,N_12546);
and U12712 (N_12712,N_12565,N_12627);
or U12713 (N_12713,N_12600,N_12611);
nor U12714 (N_12714,N_12526,N_12628);
nor U12715 (N_12715,N_12588,N_12533);
nand U12716 (N_12716,N_12572,N_12485);
nand U12717 (N_12717,N_12525,N_12484);
nand U12718 (N_12718,N_12596,N_12487);
or U12719 (N_12719,N_12574,N_12502);
nand U12720 (N_12720,N_12551,N_12593);
xor U12721 (N_12721,N_12570,N_12512);
or U12722 (N_12722,N_12600,N_12556);
and U12723 (N_12723,N_12497,N_12571);
nor U12724 (N_12724,N_12507,N_12581);
nor U12725 (N_12725,N_12480,N_12520);
nor U12726 (N_12726,N_12573,N_12623);
and U12727 (N_12727,N_12560,N_12581);
xor U12728 (N_12728,N_12488,N_12591);
xor U12729 (N_12729,N_12530,N_12541);
or U12730 (N_12730,N_12553,N_12531);
or U12731 (N_12731,N_12608,N_12627);
nor U12732 (N_12732,N_12617,N_12563);
nand U12733 (N_12733,N_12622,N_12513);
nor U12734 (N_12734,N_12554,N_12498);
and U12735 (N_12735,N_12629,N_12609);
nor U12736 (N_12736,N_12591,N_12623);
and U12737 (N_12737,N_12631,N_12484);
xnor U12738 (N_12738,N_12503,N_12515);
nor U12739 (N_12739,N_12510,N_12546);
and U12740 (N_12740,N_12498,N_12639);
nand U12741 (N_12741,N_12505,N_12619);
xor U12742 (N_12742,N_12541,N_12504);
nor U12743 (N_12743,N_12576,N_12563);
nor U12744 (N_12744,N_12533,N_12524);
or U12745 (N_12745,N_12492,N_12596);
and U12746 (N_12746,N_12585,N_12609);
or U12747 (N_12747,N_12545,N_12587);
and U12748 (N_12748,N_12518,N_12539);
xnor U12749 (N_12749,N_12567,N_12508);
nand U12750 (N_12750,N_12583,N_12587);
xnor U12751 (N_12751,N_12590,N_12512);
nor U12752 (N_12752,N_12545,N_12608);
and U12753 (N_12753,N_12617,N_12505);
nand U12754 (N_12754,N_12506,N_12504);
xnor U12755 (N_12755,N_12491,N_12626);
xor U12756 (N_12756,N_12494,N_12625);
nor U12757 (N_12757,N_12562,N_12532);
or U12758 (N_12758,N_12614,N_12636);
nand U12759 (N_12759,N_12613,N_12585);
nor U12760 (N_12760,N_12485,N_12579);
nand U12761 (N_12761,N_12638,N_12605);
and U12762 (N_12762,N_12590,N_12499);
xnor U12763 (N_12763,N_12633,N_12543);
and U12764 (N_12764,N_12638,N_12557);
nand U12765 (N_12765,N_12618,N_12606);
xor U12766 (N_12766,N_12561,N_12573);
nand U12767 (N_12767,N_12575,N_12542);
and U12768 (N_12768,N_12572,N_12533);
nor U12769 (N_12769,N_12530,N_12593);
nor U12770 (N_12770,N_12612,N_12528);
nor U12771 (N_12771,N_12605,N_12639);
or U12772 (N_12772,N_12480,N_12536);
nand U12773 (N_12773,N_12539,N_12514);
and U12774 (N_12774,N_12491,N_12529);
xor U12775 (N_12775,N_12542,N_12530);
or U12776 (N_12776,N_12523,N_12603);
and U12777 (N_12777,N_12576,N_12616);
xor U12778 (N_12778,N_12549,N_12506);
and U12779 (N_12779,N_12594,N_12576);
xor U12780 (N_12780,N_12541,N_12629);
nor U12781 (N_12781,N_12618,N_12492);
or U12782 (N_12782,N_12546,N_12551);
xnor U12783 (N_12783,N_12510,N_12526);
or U12784 (N_12784,N_12507,N_12606);
nor U12785 (N_12785,N_12553,N_12481);
or U12786 (N_12786,N_12485,N_12539);
or U12787 (N_12787,N_12565,N_12602);
nor U12788 (N_12788,N_12540,N_12618);
and U12789 (N_12789,N_12601,N_12515);
or U12790 (N_12790,N_12610,N_12499);
nand U12791 (N_12791,N_12563,N_12539);
xnor U12792 (N_12792,N_12573,N_12577);
nand U12793 (N_12793,N_12487,N_12517);
xor U12794 (N_12794,N_12606,N_12593);
nand U12795 (N_12795,N_12618,N_12620);
or U12796 (N_12796,N_12564,N_12506);
nor U12797 (N_12797,N_12551,N_12491);
and U12798 (N_12798,N_12558,N_12533);
and U12799 (N_12799,N_12547,N_12586);
xnor U12800 (N_12800,N_12764,N_12696);
nor U12801 (N_12801,N_12646,N_12718);
xor U12802 (N_12802,N_12794,N_12702);
xor U12803 (N_12803,N_12651,N_12752);
nor U12804 (N_12804,N_12647,N_12674);
nor U12805 (N_12805,N_12797,N_12687);
or U12806 (N_12806,N_12678,N_12686);
nand U12807 (N_12807,N_12644,N_12776);
nor U12808 (N_12808,N_12737,N_12736);
xor U12809 (N_12809,N_12682,N_12768);
or U12810 (N_12810,N_12705,N_12789);
xor U12811 (N_12811,N_12675,N_12712);
and U12812 (N_12812,N_12679,N_12784);
nand U12813 (N_12813,N_12798,N_12688);
xnor U12814 (N_12814,N_12668,N_12761);
or U12815 (N_12815,N_12643,N_12719);
nor U12816 (N_12816,N_12763,N_12795);
nor U12817 (N_12817,N_12706,N_12750);
nor U12818 (N_12818,N_12779,N_12726);
or U12819 (N_12819,N_12656,N_12670);
xor U12820 (N_12820,N_12648,N_12690);
nand U12821 (N_12821,N_12707,N_12650);
and U12822 (N_12822,N_12765,N_12665);
xnor U12823 (N_12823,N_12741,N_12756);
or U12824 (N_12824,N_12772,N_12669);
and U12825 (N_12825,N_12703,N_12673);
xor U12826 (N_12826,N_12698,N_12672);
nor U12827 (N_12827,N_12728,N_12739);
or U12828 (N_12828,N_12774,N_12695);
or U12829 (N_12829,N_12641,N_12713);
or U12830 (N_12830,N_12676,N_12775);
and U12831 (N_12831,N_12783,N_12704);
nor U12832 (N_12832,N_12693,N_12773);
xnor U12833 (N_12833,N_12716,N_12645);
nor U12834 (N_12834,N_12727,N_12720);
nand U12835 (N_12835,N_12640,N_12666);
and U12836 (N_12836,N_12732,N_12697);
xor U12837 (N_12837,N_12721,N_12725);
xor U12838 (N_12838,N_12754,N_12746);
nor U12839 (N_12839,N_12724,N_12662);
and U12840 (N_12840,N_12663,N_12778);
nand U12841 (N_12841,N_12755,N_12711);
nor U12842 (N_12842,N_12661,N_12745);
xor U12843 (N_12843,N_12683,N_12791);
xor U12844 (N_12844,N_12664,N_12654);
xnor U12845 (N_12845,N_12762,N_12731);
nand U12846 (N_12846,N_12792,N_12652);
nand U12847 (N_12847,N_12692,N_12677);
or U12848 (N_12848,N_12691,N_12760);
xnor U12849 (N_12849,N_12799,N_12748);
nand U12850 (N_12850,N_12708,N_12767);
and U12851 (N_12851,N_12786,N_12742);
nand U12852 (N_12852,N_12722,N_12684);
nor U12853 (N_12853,N_12667,N_12642);
nand U12854 (N_12854,N_12733,N_12714);
and U12855 (N_12855,N_12771,N_12759);
or U12856 (N_12856,N_12758,N_12782);
nand U12857 (N_12857,N_12790,N_12735);
or U12858 (N_12858,N_12657,N_12671);
xor U12859 (N_12859,N_12658,N_12738);
nor U12860 (N_12860,N_12694,N_12749);
nor U12861 (N_12861,N_12715,N_12788);
xnor U12862 (N_12862,N_12780,N_12777);
xnor U12863 (N_12863,N_12717,N_12660);
and U12864 (N_12864,N_12649,N_12734);
or U12865 (N_12865,N_12699,N_12653);
xnor U12866 (N_12866,N_12729,N_12769);
nor U12867 (N_12867,N_12744,N_12730);
nand U12868 (N_12868,N_12781,N_12710);
nand U12869 (N_12869,N_12743,N_12685);
and U12870 (N_12870,N_12753,N_12785);
and U12871 (N_12871,N_12723,N_12793);
nand U12872 (N_12872,N_12740,N_12680);
nor U12873 (N_12873,N_12655,N_12751);
xor U12874 (N_12874,N_12796,N_12747);
and U12875 (N_12875,N_12700,N_12689);
xnor U12876 (N_12876,N_12757,N_12766);
xor U12877 (N_12877,N_12770,N_12681);
nand U12878 (N_12878,N_12787,N_12659);
nor U12879 (N_12879,N_12701,N_12709);
and U12880 (N_12880,N_12766,N_12730);
and U12881 (N_12881,N_12676,N_12741);
xnor U12882 (N_12882,N_12640,N_12717);
xnor U12883 (N_12883,N_12779,N_12646);
nand U12884 (N_12884,N_12665,N_12701);
xnor U12885 (N_12885,N_12745,N_12697);
and U12886 (N_12886,N_12712,N_12775);
nor U12887 (N_12887,N_12772,N_12650);
or U12888 (N_12888,N_12714,N_12666);
and U12889 (N_12889,N_12700,N_12741);
or U12890 (N_12890,N_12644,N_12799);
or U12891 (N_12891,N_12736,N_12676);
xnor U12892 (N_12892,N_12703,N_12649);
xor U12893 (N_12893,N_12666,N_12693);
or U12894 (N_12894,N_12652,N_12693);
nor U12895 (N_12895,N_12722,N_12726);
or U12896 (N_12896,N_12704,N_12792);
xnor U12897 (N_12897,N_12685,N_12740);
or U12898 (N_12898,N_12649,N_12777);
and U12899 (N_12899,N_12674,N_12676);
nor U12900 (N_12900,N_12786,N_12739);
or U12901 (N_12901,N_12663,N_12738);
and U12902 (N_12902,N_12793,N_12715);
xnor U12903 (N_12903,N_12655,N_12757);
nand U12904 (N_12904,N_12739,N_12656);
or U12905 (N_12905,N_12754,N_12730);
or U12906 (N_12906,N_12765,N_12762);
nand U12907 (N_12907,N_12738,N_12766);
and U12908 (N_12908,N_12667,N_12761);
and U12909 (N_12909,N_12695,N_12674);
nor U12910 (N_12910,N_12792,N_12715);
or U12911 (N_12911,N_12749,N_12729);
xor U12912 (N_12912,N_12656,N_12759);
and U12913 (N_12913,N_12784,N_12753);
and U12914 (N_12914,N_12688,N_12785);
or U12915 (N_12915,N_12776,N_12730);
xnor U12916 (N_12916,N_12705,N_12648);
or U12917 (N_12917,N_12770,N_12760);
nand U12918 (N_12918,N_12744,N_12662);
or U12919 (N_12919,N_12662,N_12794);
or U12920 (N_12920,N_12703,N_12668);
and U12921 (N_12921,N_12674,N_12659);
nand U12922 (N_12922,N_12738,N_12685);
or U12923 (N_12923,N_12708,N_12706);
nor U12924 (N_12924,N_12786,N_12796);
and U12925 (N_12925,N_12715,N_12719);
nor U12926 (N_12926,N_12750,N_12768);
nand U12927 (N_12927,N_12719,N_12786);
and U12928 (N_12928,N_12791,N_12751);
xor U12929 (N_12929,N_12653,N_12680);
nor U12930 (N_12930,N_12759,N_12712);
or U12931 (N_12931,N_12666,N_12770);
nor U12932 (N_12932,N_12684,N_12799);
nor U12933 (N_12933,N_12745,N_12743);
nor U12934 (N_12934,N_12654,N_12726);
nor U12935 (N_12935,N_12762,N_12691);
xnor U12936 (N_12936,N_12734,N_12672);
and U12937 (N_12937,N_12700,N_12746);
xnor U12938 (N_12938,N_12689,N_12674);
nor U12939 (N_12939,N_12674,N_12697);
and U12940 (N_12940,N_12762,N_12661);
or U12941 (N_12941,N_12642,N_12652);
nor U12942 (N_12942,N_12780,N_12722);
or U12943 (N_12943,N_12720,N_12685);
nor U12944 (N_12944,N_12699,N_12672);
and U12945 (N_12945,N_12712,N_12782);
and U12946 (N_12946,N_12717,N_12767);
nand U12947 (N_12947,N_12698,N_12708);
nand U12948 (N_12948,N_12667,N_12640);
nor U12949 (N_12949,N_12664,N_12643);
and U12950 (N_12950,N_12715,N_12783);
or U12951 (N_12951,N_12757,N_12761);
xor U12952 (N_12952,N_12659,N_12666);
and U12953 (N_12953,N_12654,N_12728);
nor U12954 (N_12954,N_12731,N_12729);
and U12955 (N_12955,N_12733,N_12682);
and U12956 (N_12956,N_12735,N_12761);
and U12957 (N_12957,N_12678,N_12644);
and U12958 (N_12958,N_12781,N_12770);
nand U12959 (N_12959,N_12674,N_12759);
or U12960 (N_12960,N_12842,N_12932);
or U12961 (N_12961,N_12954,N_12851);
nor U12962 (N_12962,N_12836,N_12877);
nor U12963 (N_12963,N_12894,N_12807);
xnor U12964 (N_12964,N_12918,N_12818);
nand U12965 (N_12965,N_12853,N_12866);
nand U12966 (N_12966,N_12862,N_12899);
nor U12967 (N_12967,N_12887,N_12924);
nand U12968 (N_12968,N_12831,N_12893);
nand U12969 (N_12969,N_12897,N_12857);
nand U12970 (N_12970,N_12947,N_12868);
nor U12971 (N_12971,N_12870,N_12910);
or U12972 (N_12972,N_12871,N_12959);
or U12973 (N_12973,N_12815,N_12811);
and U12974 (N_12974,N_12940,N_12948);
and U12975 (N_12975,N_12944,N_12881);
xor U12976 (N_12976,N_12907,N_12895);
or U12977 (N_12977,N_12905,N_12854);
nand U12978 (N_12978,N_12847,N_12911);
xor U12979 (N_12979,N_12922,N_12845);
xor U12980 (N_12980,N_12900,N_12852);
nand U12981 (N_12981,N_12810,N_12951);
nor U12982 (N_12982,N_12873,N_12902);
or U12983 (N_12983,N_12813,N_12823);
xnor U12984 (N_12984,N_12912,N_12952);
and U12985 (N_12985,N_12927,N_12826);
and U12986 (N_12986,N_12943,N_12957);
nand U12987 (N_12987,N_12822,N_12803);
xnor U12988 (N_12988,N_12861,N_12830);
or U12989 (N_12989,N_12889,N_12812);
nor U12990 (N_12990,N_12921,N_12950);
xnor U12991 (N_12991,N_12901,N_12869);
or U12992 (N_12992,N_12829,N_12945);
or U12993 (N_12993,N_12834,N_12896);
or U12994 (N_12994,N_12875,N_12955);
xor U12995 (N_12995,N_12883,N_12953);
xor U12996 (N_12996,N_12814,N_12878);
xnor U12997 (N_12997,N_12928,N_12913);
xor U12998 (N_12998,N_12956,N_12809);
or U12999 (N_12999,N_12939,N_12936);
or U13000 (N_13000,N_12864,N_12856);
or U13001 (N_13001,N_12890,N_12863);
and U13002 (N_13002,N_12879,N_12867);
xor U13003 (N_13003,N_12929,N_12839);
or U13004 (N_13004,N_12806,N_12872);
nand U13005 (N_13005,N_12888,N_12828);
nand U13006 (N_13006,N_12804,N_12808);
and U13007 (N_13007,N_12833,N_12906);
nand U13008 (N_13008,N_12919,N_12848);
and U13009 (N_13009,N_12805,N_12909);
nand U13010 (N_13010,N_12832,N_12920);
nand U13011 (N_13011,N_12802,N_12882);
nand U13012 (N_13012,N_12855,N_12930);
and U13013 (N_13013,N_12819,N_12937);
nand U13014 (N_13014,N_12898,N_12840);
or U13015 (N_13015,N_12800,N_12865);
or U13016 (N_13016,N_12820,N_12935);
nor U13017 (N_13017,N_12859,N_12850);
and U13018 (N_13018,N_12821,N_12903);
nand U13019 (N_13019,N_12843,N_12884);
or U13020 (N_13020,N_12860,N_12874);
nand U13021 (N_13021,N_12931,N_12914);
xor U13022 (N_13022,N_12958,N_12925);
nor U13023 (N_13023,N_12825,N_12824);
nand U13024 (N_13024,N_12838,N_12827);
nand U13025 (N_13025,N_12801,N_12917);
or U13026 (N_13026,N_12841,N_12938);
nand U13027 (N_13027,N_12885,N_12946);
xnor U13028 (N_13028,N_12942,N_12849);
nor U13029 (N_13029,N_12949,N_12816);
xor U13030 (N_13030,N_12908,N_12876);
nand U13031 (N_13031,N_12934,N_12844);
xnor U13032 (N_13032,N_12837,N_12933);
nand U13033 (N_13033,N_12904,N_12880);
nor U13034 (N_13034,N_12892,N_12923);
or U13035 (N_13035,N_12817,N_12858);
and U13036 (N_13036,N_12915,N_12846);
or U13037 (N_13037,N_12886,N_12926);
and U13038 (N_13038,N_12835,N_12916);
and U13039 (N_13039,N_12941,N_12891);
nand U13040 (N_13040,N_12833,N_12859);
nand U13041 (N_13041,N_12939,N_12856);
xor U13042 (N_13042,N_12924,N_12921);
xnor U13043 (N_13043,N_12926,N_12839);
or U13044 (N_13044,N_12881,N_12855);
and U13045 (N_13045,N_12902,N_12925);
nand U13046 (N_13046,N_12873,N_12812);
nand U13047 (N_13047,N_12924,N_12927);
nor U13048 (N_13048,N_12823,N_12857);
nor U13049 (N_13049,N_12865,N_12911);
or U13050 (N_13050,N_12905,N_12871);
and U13051 (N_13051,N_12894,N_12883);
nand U13052 (N_13052,N_12827,N_12941);
xor U13053 (N_13053,N_12910,N_12894);
nor U13054 (N_13054,N_12930,N_12854);
nand U13055 (N_13055,N_12940,N_12878);
nor U13056 (N_13056,N_12863,N_12806);
nor U13057 (N_13057,N_12865,N_12818);
xor U13058 (N_13058,N_12913,N_12846);
nand U13059 (N_13059,N_12829,N_12802);
xnor U13060 (N_13060,N_12848,N_12840);
nor U13061 (N_13061,N_12830,N_12914);
and U13062 (N_13062,N_12875,N_12865);
or U13063 (N_13063,N_12868,N_12943);
and U13064 (N_13064,N_12814,N_12927);
nor U13065 (N_13065,N_12949,N_12850);
nand U13066 (N_13066,N_12870,N_12807);
nand U13067 (N_13067,N_12808,N_12949);
nor U13068 (N_13068,N_12879,N_12938);
xnor U13069 (N_13069,N_12915,N_12889);
and U13070 (N_13070,N_12887,N_12953);
nand U13071 (N_13071,N_12823,N_12878);
nand U13072 (N_13072,N_12847,N_12822);
xor U13073 (N_13073,N_12804,N_12827);
or U13074 (N_13074,N_12878,N_12875);
nand U13075 (N_13075,N_12848,N_12957);
nand U13076 (N_13076,N_12872,N_12847);
xnor U13077 (N_13077,N_12840,N_12833);
or U13078 (N_13078,N_12909,N_12947);
nor U13079 (N_13079,N_12953,N_12956);
xnor U13080 (N_13080,N_12803,N_12865);
and U13081 (N_13081,N_12870,N_12876);
nand U13082 (N_13082,N_12841,N_12832);
nor U13083 (N_13083,N_12856,N_12806);
xor U13084 (N_13084,N_12894,N_12842);
nor U13085 (N_13085,N_12874,N_12842);
and U13086 (N_13086,N_12909,N_12861);
or U13087 (N_13087,N_12832,N_12925);
nand U13088 (N_13088,N_12823,N_12915);
nand U13089 (N_13089,N_12895,N_12874);
or U13090 (N_13090,N_12866,N_12806);
nand U13091 (N_13091,N_12941,N_12955);
and U13092 (N_13092,N_12801,N_12848);
nand U13093 (N_13093,N_12802,N_12933);
xnor U13094 (N_13094,N_12917,N_12939);
nand U13095 (N_13095,N_12886,N_12821);
nand U13096 (N_13096,N_12954,N_12843);
and U13097 (N_13097,N_12857,N_12866);
nand U13098 (N_13098,N_12897,N_12819);
and U13099 (N_13099,N_12809,N_12807);
nand U13100 (N_13100,N_12844,N_12891);
nor U13101 (N_13101,N_12833,N_12890);
xnor U13102 (N_13102,N_12938,N_12821);
xnor U13103 (N_13103,N_12842,N_12837);
or U13104 (N_13104,N_12850,N_12829);
xor U13105 (N_13105,N_12882,N_12871);
xnor U13106 (N_13106,N_12832,N_12857);
nand U13107 (N_13107,N_12947,N_12805);
and U13108 (N_13108,N_12954,N_12923);
xor U13109 (N_13109,N_12893,N_12926);
nand U13110 (N_13110,N_12885,N_12958);
or U13111 (N_13111,N_12950,N_12954);
xor U13112 (N_13112,N_12854,N_12805);
and U13113 (N_13113,N_12835,N_12935);
xnor U13114 (N_13114,N_12904,N_12955);
and U13115 (N_13115,N_12907,N_12825);
and U13116 (N_13116,N_12869,N_12849);
and U13117 (N_13117,N_12861,N_12931);
nor U13118 (N_13118,N_12800,N_12806);
or U13119 (N_13119,N_12821,N_12862);
or U13120 (N_13120,N_13097,N_13099);
xor U13121 (N_13121,N_12971,N_12963);
xor U13122 (N_13122,N_13050,N_13066);
nand U13123 (N_13123,N_12989,N_13009);
or U13124 (N_13124,N_13044,N_12962);
and U13125 (N_13125,N_13023,N_13000);
nor U13126 (N_13126,N_13033,N_12976);
nor U13127 (N_13127,N_13042,N_13024);
nor U13128 (N_13128,N_13016,N_12975);
and U13129 (N_13129,N_12991,N_13080);
nand U13130 (N_13130,N_13071,N_13012);
xnor U13131 (N_13131,N_13086,N_12995);
xor U13132 (N_13132,N_12998,N_13063);
xnor U13133 (N_13133,N_13106,N_12994);
nor U13134 (N_13134,N_13112,N_13020);
and U13135 (N_13135,N_13007,N_13003);
nor U13136 (N_13136,N_12979,N_12967);
nand U13137 (N_13137,N_13072,N_13059);
and U13138 (N_13138,N_12993,N_13095);
xor U13139 (N_13139,N_13002,N_13111);
and U13140 (N_13140,N_13008,N_13021);
nor U13141 (N_13141,N_13026,N_13055);
xor U13142 (N_13142,N_12972,N_13038);
or U13143 (N_13143,N_13025,N_13093);
nand U13144 (N_13144,N_12977,N_13067);
nand U13145 (N_13145,N_13028,N_12983);
and U13146 (N_13146,N_13001,N_12992);
and U13147 (N_13147,N_13117,N_13114);
and U13148 (N_13148,N_12999,N_13079);
nand U13149 (N_13149,N_13041,N_13010);
xnor U13150 (N_13150,N_13083,N_13015);
and U13151 (N_13151,N_13094,N_12985);
and U13152 (N_13152,N_13075,N_13078);
xnor U13153 (N_13153,N_13036,N_13104);
and U13154 (N_13154,N_13013,N_13074);
or U13155 (N_13155,N_13107,N_13032);
nand U13156 (N_13156,N_13060,N_12984);
or U13157 (N_13157,N_13088,N_13054);
and U13158 (N_13158,N_12964,N_12970);
nand U13159 (N_13159,N_13037,N_12982);
xor U13160 (N_13160,N_13053,N_13014);
or U13161 (N_13161,N_13089,N_13061);
and U13162 (N_13162,N_12974,N_13085);
nand U13163 (N_13163,N_13049,N_13052);
or U13164 (N_13164,N_12965,N_13057);
xor U13165 (N_13165,N_12981,N_13034);
nand U13166 (N_13166,N_13030,N_13087);
and U13167 (N_13167,N_13076,N_12961);
nand U13168 (N_13168,N_13103,N_13022);
nand U13169 (N_13169,N_13043,N_13109);
xor U13170 (N_13170,N_13098,N_13019);
xor U13171 (N_13171,N_12978,N_13064);
and U13172 (N_13172,N_13119,N_12990);
xor U13173 (N_13173,N_13058,N_12986);
nor U13174 (N_13174,N_13069,N_13116);
xor U13175 (N_13175,N_13084,N_13082);
and U13176 (N_13176,N_12980,N_13105);
nand U13177 (N_13177,N_13005,N_13100);
xor U13178 (N_13178,N_13110,N_13115);
nor U13179 (N_13179,N_13068,N_13118);
nor U13180 (N_13180,N_13081,N_12969);
nand U13181 (N_13181,N_13045,N_13073);
or U13182 (N_13182,N_13113,N_12973);
xor U13183 (N_13183,N_13006,N_13027);
nand U13184 (N_13184,N_12996,N_13048);
or U13185 (N_13185,N_12960,N_12988);
and U13186 (N_13186,N_13011,N_13065);
and U13187 (N_13187,N_13108,N_13101);
and U13188 (N_13188,N_13102,N_12987);
nor U13189 (N_13189,N_13004,N_13092);
nor U13190 (N_13190,N_13077,N_12966);
and U13191 (N_13191,N_13017,N_13090);
or U13192 (N_13192,N_13062,N_13035);
xor U13193 (N_13193,N_13056,N_13091);
or U13194 (N_13194,N_13031,N_13029);
nand U13195 (N_13195,N_13047,N_13096);
or U13196 (N_13196,N_13070,N_13039);
or U13197 (N_13197,N_12968,N_13051);
xnor U13198 (N_13198,N_13046,N_12997);
or U13199 (N_13199,N_13018,N_13040);
xnor U13200 (N_13200,N_13107,N_13091);
or U13201 (N_13201,N_13090,N_13030);
nor U13202 (N_13202,N_12999,N_13077);
or U13203 (N_13203,N_13005,N_13118);
or U13204 (N_13204,N_13052,N_13033);
and U13205 (N_13205,N_13102,N_13016);
and U13206 (N_13206,N_13114,N_13019);
xor U13207 (N_13207,N_13099,N_12979);
nor U13208 (N_13208,N_12972,N_13047);
and U13209 (N_13209,N_13019,N_12981);
or U13210 (N_13210,N_12983,N_13039);
xnor U13211 (N_13211,N_13009,N_12992);
or U13212 (N_13212,N_13035,N_13043);
or U13213 (N_13213,N_12999,N_13094);
nor U13214 (N_13214,N_13059,N_13001);
or U13215 (N_13215,N_13071,N_12962);
xnor U13216 (N_13216,N_13044,N_13115);
nor U13217 (N_13217,N_13080,N_12968);
or U13218 (N_13218,N_13052,N_13004);
or U13219 (N_13219,N_13057,N_12990);
nand U13220 (N_13220,N_12982,N_12963);
nand U13221 (N_13221,N_13027,N_13077);
nand U13222 (N_13222,N_13089,N_12998);
nor U13223 (N_13223,N_13063,N_13095);
xor U13224 (N_13224,N_13025,N_13109);
and U13225 (N_13225,N_13035,N_13016);
nand U13226 (N_13226,N_13013,N_13061);
xnor U13227 (N_13227,N_13072,N_13095);
and U13228 (N_13228,N_13013,N_13079);
nor U13229 (N_13229,N_13055,N_13039);
or U13230 (N_13230,N_13113,N_13033);
xor U13231 (N_13231,N_13092,N_12986);
and U13232 (N_13232,N_13104,N_13043);
nand U13233 (N_13233,N_13013,N_13004);
xnor U13234 (N_13234,N_13039,N_13083);
nor U13235 (N_13235,N_12998,N_13076);
nor U13236 (N_13236,N_12985,N_12975);
nor U13237 (N_13237,N_12961,N_13077);
and U13238 (N_13238,N_12984,N_13079);
xnor U13239 (N_13239,N_13000,N_13032);
or U13240 (N_13240,N_13084,N_12991);
and U13241 (N_13241,N_13029,N_13088);
xor U13242 (N_13242,N_12991,N_13098);
xor U13243 (N_13243,N_13096,N_13075);
or U13244 (N_13244,N_13070,N_13049);
or U13245 (N_13245,N_13102,N_13035);
nand U13246 (N_13246,N_13023,N_12998);
or U13247 (N_13247,N_12995,N_13008);
nand U13248 (N_13248,N_12987,N_13098);
xor U13249 (N_13249,N_13039,N_13044);
and U13250 (N_13250,N_13116,N_13071);
or U13251 (N_13251,N_13073,N_13113);
nor U13252 (N_13252,N_13071,N_13088);
nor U13253 (N_13253,N_12974,N_12963);
nor U13254 (N_13254,N_12975,N_13064);
nand U13255 (N_13255,N_12981,N_13101);
xor U13256 (N_13256,N_13105,N_13036);
xnor U13257 (N_13257,N_12967,N_12989);
xnor U13258 (N_13258,N_12997,N_13001);
nand U13259 (N_13259,N_13074,N_13113);
or U13260 (N_13260,N_12996,N_12985);
nor U13261 (N_13261,N_13055,N_12960);
xor U13262 (N_13262,N_13084,N_13107);
or U13263 (N_13263,N_13116,N_12991);
xor U13264 (N_13264,N_13089,N_13099);
nand U13265 (N_13265,N_13009,N_13103);
nor U13266 (N_13266,N_12988,N_13023);
and U13267 (N_13267,N_13025,N_13074);
and U13268 (N_13268,N_13099,N_13005);
and U13269 (N_13269,N_13079,N_13035);
nor U13270 (N_13270,N_13032,N_13003);
nand U13271 (N_13271,N_13015,N_13011);
and U13272 (N_13272,N_13117,N_12977);
nor U13273 (N_13273,N_13061,N_13104);
and U13274 (N_13274,N_13063,N_12978);
xnor U13275 (N_13275,N_13056,N_12986);
and U13276 (N_13276,N_13029,N_12996);
nor U13277 (N_13277,N_13074,N_13104);
and U13278 (N_13278,N_13061,N_13016);
and U13279 (N_13279,N_13104,N_13101);
or U13280 (N_13280,N_13142,N_13221);
and U13281 (N_13281,N_13202,N_13257);
or U13282 (N_13282,N_13239,N_13178);
or U13283 (N_13283,N_13185,N_13217);
nor U13284 (N_13284,N_13154,N_13131);
nor U13285 (N_13285,N_13124,N_13259);
nand U13286 (N_13286,N_13220,N_13245);
or U13287 (N_13287,N_13275,N_13197);
xor U13288 (N_13288,N_13238,N_13193);
nand U13289 (N_13289,N_13180,N_13125);
xor U13290 (N_13290,N_13147,N_13153);
xnor U13291 (N_13291,N_13137,N_13122);
or U13292 (N_13292,N_13121,N_13167);
nand U13293 (N_13293,N_13132,N_13272);
and U13294 (N_13294,N_13252,N_13133);
nand U13295 (N_13295,N_13258,N_13278);
and U13296 (N_13296,N_13173,N_13236);
and U13297 (N_13297,N_13253,N_13208);
xor U13298 (N_13298,N_13191,N_13189);
or U13299 (N_13299,N_13279,N_13267);
or U13300 (N_13300,N_13145,N_13234);
nand U13301 (N_13301,N_13261,N_13138);
or U13302 (N_13302,N_13175,N_13251);
xor U13303 (N_13303,N_13210,N_13225);
and U13304 (N_13304,N_13213,N_13172);
and U13305 (N_13305,N_13196,N_13266);
or U13306 (N_13306,N_13222,N_13195);
nor U13307 (N_13307,N_13166,N_13155);
nor U13308 (N_13308,N_13143,N_13174);
xor U13309 (N_13309,N_13148,N_13273);
nor U13310 (N_13310,N_13128,N_13216);
nand U13311 (N_13311,N_13201,N_13264);
nand U13312 (N_13312,N_13235,N_13246);
nand U13313 (N_13313,N_13186,N_13149);
or U13314 (N_13314,N_13150,N_13228);
or U13315 (N_13315,N_13194,N_13255);
or U13316 (N_13316,N_13209,N_13232);
nor U13317 (N_13317,N_13270,N_13223);
xnor U13318 (N_13318,N_13237,N_13199);
and U13319 (N_13319,N_13152,N_13157);
xnor U13320 (N_13320,N_13229,N_13248);
or U13321 (N_13321,N_13120,N_13215);
nand U13322 (N_13322,N_13187,N_13226);
xnor U13323 (N_13323,N_13161,N_13244);
nand U13324 (N_13324,N_13269,N_13190);
xor U13325 (N_13325,N_13224,N_13200);
or U13326 (N_13326,N_13126,N_13205);
nand U13327 (N_13327,N_13140,N_13231);
or U13328 (N_13328,N_13129,N_13182);
and U13329 (N_13329,N_13162,N_13268);
nand U13330 (N_13330,N_13158,N_13274);
nand U13331 (N_13331,N_13168,N_13276);
nor U13332 (N_13332,N_13170,N_13179);
xor U13333 (N_13333,N_13159,N_13139);
and U13334 (N_13334,N_13206,N_13135);
xnor U13335 (N_13335,N_13260,N_13256);
xor U13336 (N_13336,N_13227,N_13151);
xnor U13337 (N_13337,N_13136,N_13241);
and U13338 (N_13338,N_13123,N_13203);
xor U13339 (N_13339,N_13204,N_13130);
or U13340 (N_13340,N_13277,N_13127);
nand U13341 (N_13341,N_13249,N_13156);
nor U13342 (N_13342,N_13247,N_13164);
or U13343 (N_13343,N_13230,N_13233);
and U13344 (N_13344,N_13198,N_13192);
nand U13345 (N_13345,N_13271,N_13141);
nor U13346 (N_13346,N_13165,N_13212);
xor U13347 (N_13347,N_13254,N_13265);
and U13348 (N_13348,N_13218,N_13242);
or U13349 (N_13349,N_13214,N_13171);
or U13350 (N_13350,N_13134,N_13184);
xnor U13351 (N_13351,N_13163,N_13262);
nand U13352 (N_13352,N_13183,N_13181);
or U13353 (N_13353,N_13240,N_13250);
and U13354 (N_13354,N_13176,N_13177);
or U13355 (N_13355,N_13144,N_13263);
xnor U13356 (N_13356,N_13219,N_13169);
nor U13357 (N_13357,N_13207,N_13160);
nand U13358 (N_13358,N_13188,N_13146);
xnor U13359 (N_13359,N_13211,N_13243);
and U13360 (N_13360,N_13222,N_13237);
nor U13361 (N_13361,N_13153,N_13248);
and U13362 (N_13362,N_13129,N_13214);
nor U13363 (N_13363,N_13207,N_13265);
or U13364 (N_13364,N_13240,N_13210);
or U13365 (N_13365,N_13270,N_13164);
nor U13366 (N_13366,N_13269,N_13135);
xnor U13367 (N_13367,N_13182,N_13279);
or U13368 (N_13368,N_13166,N_13124);
nor U13369 (N_13369,N_13273,N_13275);
and U13370 (N_13370,N_13129,N_13248);
and U13371 (N_13371,N_13153,N_13250);
or U13372 (N_13372,N_13131,N_13153);
xor U13373 (N_13373,N_13143,N_13167);
or U13374 (N_13374,N_13261,N_13130);
nand U13375 (N_13375,N_13172,N_13237);
xor U13376 (N_13376,N_13125,N_13148);
nor U13377 (N_13377,N_13198,N_13165);
and U13378 (N_13378,N_13255,N_13248);
and U13379 (N_13379,N_13276,N_13187);
xor U13380 (N_13380,N_13246,N_13199);
and U13381 (N_13381,N_13152,N_13179);
xor U13382 (N_13382,N_13196,N_13175);
and U13383 (N_13383,N_13176,N_13271);
and U13384 (N_13384,N_13179,N_13211);
and U13385 (N_13385,N_13218,N_13257);
and U13386 (N_13386,N_13200,N_13262);
or U13387 (N_13387,N_13121,N_13177);
xnor U13388 (N_13388,N_13210,N_13211);
or U13389 (N_13389,N_13206,N_13165);
or U13390 (N_13390,N_13158,N_13237);
and U13391 (N_13391,N_13196,N_13246);
nor U13392 (N_13392,N_13131,N_13138);
and U13393 (N_13393,N_13249,N_13168);
or U13394 (N_13394,N_13123,N_13215);
and U13395 (N_13395,N_13211,N_13256);
and U13396 (N_13396,N_13240,N_13181);
nand U13397 (N_13397,N_13224,N_13147);
and U13398 (N_13398,N_13166,N_13167);
nor U13399 (N_13399,N_13265,N_13235);
nor U13400 (N_13400,N_13259,N_13180);
nor U13401 (N_13401,N_13186,N_13225);
nor U13402 (N_13402,N_13278,N_13165);
nor U13403 (N_13403,N_13278,N_13157);
xor U13404 (N_13404,N_13154,N_13158);
or U13405 (N_13405,N_13253,N_13169);
nor U13406 (N_13406,N_13120,N_13150);
xor U13407 (N_13407,N_13225,N_13216);
or U13408 (N_13408,N_13186,N_13220);
or U13409 (N_13409,N_13273,N_13260);
nand U13410 (N_13410,N_13150,N_13236);
and U13411 (N_13411,N_13219,N_13159);
nand U13412 (N_13412,N_13277,N_13196);
xnor U13413 (N_13413,N_13161,N_13167);
nand U13414 (N_13414,N_13274,N_13178);
nand U13415 (N_13415,N_13141,N_13221);
nor U13416 (N_13416,N_13247,N_13218);
xnor U13417 (N_13417,N_13259,N_13240);
nand U13418 (N_13418,N_13223,N_13177);
or U13419 (N_13419,N_13180,N_13208);
nand U13420 (N_13420,N_13276,N_13229);
or U13421 (N_13421,N_13214,N_13254);
and U13422 (N_13422,N_13209,N_13241);
nand U13423 (N_13423,N_13174,N_13211);
and U13424 (N_13424,N_13204,N_13243);
nand U13425 (N_13425,N_13138,N_13180);
xor U13426 (N_13426,N_13238,N_13262);
nor U13427 (N_13427,N_13120,N_13205);
and U13428 (N_13428,N_13173,N_13273);
or U13429 (N_13429,N_13235,N_13189);
xor U13430 (N_13430,N_13219,N_13136);
nand U13431 (N_13431,N_13143,N_13279);
nor U13432 (N_13432,N_13183,N_13161);
nand U13433 (N_13433,N_13145,N_13120);
and U13434 (N_13434,N_13176,N_13220);
nor U13435 (N_13435,N_13209,N_13222);
nor U13436 (N_13436,N_13186,N_13156);
or U13437 (N_13437,N_13254,N_13276);
and U13438 (N_13438,N_13276,N_13158);
and U13439 (N_13439,N_13268,N_13144);
and U13440 (N_13440,N_13328,N_13300);
nor U13441 (N_13441,N_13305,N_13437);
nor U13442 (N_13442,N_13391,N_13409);
and U13443 (N_13443,N_13315,N_13417);
or U13444 (N_13444,N_13311,N_13334);
nand U13445 (N_13445,N_13291,N_13384);
or U13446 (N_13446,N_13349,N_13286);
and U13447 (N_13447,N_13280,N_13321);
and U13448 (N_13448,N_13307,N_13297);
and U13449 (N_13449,N_13374,N_13287);
nor U13450 (N_13450,N_13314,N_13325);
nor U13451 (N_13451,N_13419,N_13304);
xor U13452 (N_13452,N_13352,N_13302);
or U13453 (N_13453,N_13290,N_13296);
or U13454 (N_13454,N_13295,N_13401);
or U13455 (N_13455,N_13331,N_13299);
or U13456 (N_13456,N_13337,N_13430);
xnor U13457 (N_13457,N_13285,N_13399);
and U13458 (N_13458,N_13412,N_13421);
xor U13459 (N_13459,N_13336,N_13416);
or U13460 (N_13460,N_13365,N_13429);
or U13461 (N_13461,N_13432,N_13434);
nand U13462 (N_13462,N_13306,N_13415);
nor U13463 (N_13463,N_13406,N_13340);
nor U13464 (N_13464,N_13301,N_13342);
or U13465 (N_13465,N_13338,N_13375);
xor U13466 (N_13466,N_13383,N_13358);
or U13467 (N_13467,N_13322,N_13390);
nand U13468 (N_13468,N_13402,N_13392);
xnor U13469 (N_13469,N_13425,N_13389);
or U13470 (N_13470,N_13403,N_13319);
nand U13471 (N_13471,N_13424,N_13317);
nand U13472 (N_13472,N_13363,N_13353);
or U13473 (N_13473,N_13376,N_13318);
nor U13474 (N_13474,N_13366,N_13386);
or U13475 (N_13475,N_13354,N_13393);
nor U13476 (N_13476,N_13382,N_13379);
and U13477 (N_13477,N_13388,N_13438);
nand U13478 (N_13478,N_13281,N_13293);
nor U13479 (N_13479,N_13436,N_13378);
and U13480 (N_13480,N_13369,N_13368);
and U13481 (N_13481,N_13335,N_13345);
and U13482 (N_13482,N_13360,N_13398);
or U13483 (N_13483,N_13431,N_13404);
or U13484 (N_13484,N_13405,N_13394);
xnor U13485 (N_13485,N_13326,N_13284);
nor U13486 (N_13486,N_13371,N_13288);
or U13487 (N_13487,N_13292,N_13426);
nand U13488 (N_13488,N_13364,N_13303);
xnor U13489 (N_13489,N_13413,N_13414);
nand U13490 (N_13490,N_13370,N_13312);
nand U13491 (N_13491,N_13408,N_13330);
nor U13492 (N_13492,N_13410,N_13346);
nor U13493 (N_13493,N_13324,N_13313);
nor U13494 (N_13494,N_13373,N_13418);
and U13495 (N_13495,N_13367,N_13423);
and U13496 (N_13496,N_13294,N_13381);
or U13497 (N_13497,N_13355,N_13348);
nor U13498 (N_13498,N_13396,N_13411);
xnor U13499 (N_13499,N_13377,N_13356);
nor U13500 (N_13500,N_13309,N_13359);
and U13501 (N_13501,N_13316,N_13283);
nand U13502 (N_13502,N_13435,N_13372);
nand U13503 (N_13503,N_13339,N_13343);
or U13504 (N_13504,N_13433,N_13310);
and U13505 (N_13505,N_13427,N_13351);
xnor U13506 (N_13506,N_13407,N_13387);
nor U13507 (N_13507,N_13439,N_13400);
nand U13508 (N_13508,N_13327,N_13344);
nand U13509 (N_13509,N_13347,N_13385);
and U13510 (N_13510,N_13329,N_13282);
nand U13511 (N_13511,N_13298,N_13397);
xnor U13512 (N_13512,N_13332,N_13357);
nand U13513 (N_13513,N_13362,N_13289);
nor U13514 (N_13514,N_13350,N_13395);
xnor U13515 (N_13515,N_13380,N_13323);
nor U13516 (N_13516,N_13320,N_13341);
nand U13517 (N_13517,N_13422,N_13308);
nand U13518 (N_13518,N_13361,N_13428);
nor U13519 (N_13519,N_13420,N_13333);
and U13520 (N_13520,N_13426,N_13357);
or U13521 (N_13521,N_13331,N_13427);
nand U13522 (N_13522,N_13418,N_13430);
nand U13523 (N_13523,N_13337,N_13325);
xnor U13524 (N_13524,N_13345,N_13369);
nand U13525 (N_13525,N_13374,N_13320);
nor U13526 (N_13526,N_13336,N_13378);
and U13527 (N_13527,N_13414,N_13399);
and U13528 (N_13528,N_13308,N_13385);
and U13529 (N_13529,N_13378,N_13348);
or U13530 (N_13530,N_13314,N_13394);
nor U13531 (N_13531,N_13307,N_13347);
or U13532 (N_13532,N_13286,N_13376);
or U13533 (N_13533,N_13400,N_13402);
or U13534 (N_13534,N_13414,N_13321);
or U13535 (N_13535,N_13419,N_13432);
nand U13536 (N_13536,N_13412,N_13330);
xor U13537 (N_13537,N_13367,N_13311);
xnor U13538 (N_13538,N_13420,N_13319);
or U13539 (N_13539,N_13358,N_13370);
xor U13540 (N_13540,N_13364,N_13343);
nor U13541 (N_13541,N_13409,N_13312);
and U13542 (N_13542,N_13354,N_13283);
nor U13543 (N_13543,N_13357,N_13363);
xor U13544 (N_13544,N_13280,N_13320);
nor U13545 (N_13545,N_13283,N_13330);
nor U13546 (N_13546,N_13389,N_13431);
and U13547 (N_13547,N_13281,N_13321);
and U13548 (N_13548,N_13302,N_13299);
xor U13549 (N_13549,N_13301,N_13365);
nor U13550 (N_13550,N_13399,N_13352);
xor U13551 (N_13551,N_13337,N_13312);
nor U13552 (N_13552,N_13405,N_13363);
nor U13553 (N_13553,N_13318,N_13384);
xnor U13554 (N_13554,N_13437,N_13316);
nand U13555 (N_13555,N_13390,N_13357);
nor U13556 (N_13556,N_13385,N_13359);
or U13557 (N_13557,N_13345,N_13370);
and U13558 (N_13558,N_13360,N_13401);
xnor U13559 (N_13559,N_13389,N_13418);
nand U13560 (N_13560,N_13436,N_13377);
or U13561 (N_13561,N_13361,N_13312);
or U13562 (N_13562,N_13368,N_13291);
nor U13563 (N_13563,N_13394,N_13385);
nand U13564 (N_13564,N_13340,N_13313);
nor U13565 (N_13565,N_13332,N_13388);
and U13566 (N_13566,N_13326,N_13354);
nor U13567 (N_13567,N_13298,N_13422);
xor U13568 (N_13568,N_13364,N_13350);
and U13569 (N_13569,N_13414,N_13433);
nand U13570 (N_13570,N_13343,N_13354);
and U13571 (N_13571,N_13281,N_13370);
nor U13572 (N_13572,N_13399,N_13395);
nor U13573 (N_13573,N_13377,N_13402);
nand U13574 (N_13574,N_13438,N_13390);
nand U13575 (N_13575,N_13377,N_13354);
nand U13576 (N_13576,N_13424,N_13414);
or U13577 (N_13577,N_13337,N_13367);
nand U13578 (N_13578,N_13379,N_13289);
or U13579 (N_13579,N_13366,N_13334);
or U13580 (N_13580,N_13392,N_13399);
or U13581 (N_13581,N_13281,N_13418);
nor U13582 (N_13582,N_13418,N_13412);
xor U13583 (N_13583,N_13327,N_13320);
or U13584 (N_13584,N_13433,N_13287);
xor U13585 (N_13585,N_13359,N_13374);
and U13586 (N_13586,N_13324,N_13387);
nor U13587 (N_13587,N_13293,N_13332);
xnor U13588 (N_13588,N_13347,N_13351);
and U13589 (N_13589,N_13377,N_13293);
xnor U13590 (N_13590,N_13304,N_13407);
nor U13591 (N_13591,N_13340,N_13314);
xnor U13592 (N_13592,N_13308,N_13292);
nand U13593 (N_13593,N_13344,N_13345);
and U13594 (N_13594,N_13420,N_13309);
nand U13595 (N_13595,N_13366,N_13412);
nor U13596 (N_13596,N_13402,N_13435);
and U13597 (N_13597,N_13343,N_13375);
and U13598 (N_13598,N_13285,N_13408);
nor U13599 (N_13599,N_13345,N_13375);
xor U13600 (N_13600,N_13472,N_13458);
nand U13601 (N_13601,N_13561,N_13521);
nor U13602 (N_13602,N_13571,N_13443);
nor U13603 (N_13603,N_13459,N_13471);
nand U13604 (N_13604,N_13509,N_13485);
xnor U13605 (N_13605,N_13511,N_13499);
nor U13606 (N_13606,N_13558,N_13582);
or U13607 (N_13607,N_13560,N_13502);
or U13608 (N_13608,N_13504,N_13514);
and U13609 (N_13609,N_13552,N_13475);
xnor U13610 (N_13610,N_13454,N_13526);
nand U13611 (N_13611,N_13455,N_13587);
and U13612 (N_13612,N_13528,N_13501);
xor U13613 (N_13613,N_13577,N_13545);
xnor U13614 (N_13614,N_13462,N_13556);
xnor U13615 (N_13615,N_13522,N_13595);
nand U13616 (N_13616,N_13481,N_13478);
nand U13617 (N_13617,N_13566,N_13555);
and U13618 (N_13618,N_13540,N_13541);
and U13619 (N_13619,N_13529,N_13483);
xnor U13620 (N_13620,N_13453,N_13533);
and U13621 (N_13621,N_13574,N_13447);
and U13622 (N_13622,N_13470,N_13508);
and U13623 (N_13623,N_13538,N_13477);
or U13624 (N_13624,N_13591,N_13512);
xor U13625 (N_13625,N_13482,N_13518);
nor U13626 (N_13626,N_13583,N_13452);
nand U13627 (N_13627,N_13489,N_13564);
nand U13628 (N_13628,N_13527,N_13559);
nand U13629 (N_13629,N_13542,N_13519);
or U13630 (N_13630,N_13570,N_13565);
or U13631 (N_13631,N_13479,N_13568);
nor U13632 (N_13632,N_13513,N_13491);
nor U13633 (N_13633,N_13449,N_13503);
nand U13634 (N_13634,N_13493,N_13547);
and U13635 (N_13635,N_13579,N_13534);
or U13636 (N_13636,N_13554,N_13525);
nand U13637 (N_13637,N_13578,N_13457);
nand U13638 (N_13638,N_13563,N_13498);
or U13639 (N_13639,N_13451,N_13446);
xnor U13640 (N_13640,N_13496,N_13590);
xor U13641 (N_13641,N_13494,N_13569);
xnor U13642 (N_13642,N_13549,N_13450);
or U13643 (N_13643,N_13575,N_13573);
nor U13644 (N_13644,N_13473,N_13581);
or U13645 (N_13645,N_13536,N_13572);
and U13646 (N_13646,N_13497,N_13585);
and U13647 (N_13647,N_13445,N_13539);
xor U13648 (N_13648,N_13535,N_13480);
and U13649 (N_13649,N_13500,N_13466);
or U13650 (N_13650,N_13476,N_13507);
nor U13651 (N_13651,N_13546,N_13505);
and U13652 (N_13652,N_13488,N_13557);
xor U13653 (N_13653,N_13510,N_13593);
and U13654 (N_13654,N_13598,N_13567);
nand U13655 (N_13655,N_13440,N_13463);
and U13656 (N_13656,N_13495,N_13467);
xor U13657 (N_13657,N_13456,N_13490);
nor U13658 (N_13658,N_13531,N_13594);
and U13659 (N_13659,N_13589,N_13441);
or U13660 (N_13660,N_13544,N_13515);
or U13661 (N_13661,N_13516,N_13469);
or U13662 (N_13662,N_13592,N_13576);
nand U13663 (N_13663,N_13537,N_13586);
or U13664 (N_13664,N_13448,N_13465);
xor U13665 (N_13665,N_13468,N_13461);
xnor U13666 (N_13666,N_13597,N_13486);
and U13667 (N_13667,N_13484,N_13460);
xor U13668 (N_13668,N_13442,N_13548);
and U13669 (N_13669,N_13524,N_13523);
xor U13670 (N_13670,N_13492,N_13474);
xnor U13671 (N_13671,N_13553,N_13599);
xor U13672 (N_13672,N_13530,N_13532);
xor U13673 (N_13673,N_13506,N_13584);
or U13674 (N_13674,N_13551,N_13580);
or U13675 (N_13675,N_13596,N_13464);
or U13676 (N_13676,N_13517,N_13543);
nor U13677 (N_13677,N_13520,N_13550);
nor U13678 (N_13678,N_13444,N_13562);
or U13679 (N_13679,N_13487,N_13588);
or U13680 (N_13680,N_13512,N_13563);
or U13681 (N_13681,N_13457,N_13555);
and U13682 (N_13682,N_13530,N_13462);
xor U13683 (N_13683,N_13523,N_13553);
nor U13684 (N_13684,N_13561,N_13562);
or U13685 (N_13685,N_13569,N_13555);
nor U13686 (N_13686,N_13584,N_13540);
or U13687 (N_13687,N_13578,N_13524);
xor U13688 (N_13688,N_13462,N_13584);
nand U13689 (N_13689,N_13501,N_13492);
nor U13690 (N_13690,N_13479,N_13455);
xnor U13691 (N_13691,N_13453,N_13526);
xor U13692 (N_13692,N_13514,N_13443);
or U13693 (N_13693,N_13463,N_13495);
and U13694 (N_13694,N_13566,N_13480);
and U13695 (N_13695,N_13529,N_13501);
nor U13696 (N_13696,N_13458,N_13589);
nor U13697 (N_13697,N_13516,N_13495);
nor U13698 (N_13698,N_13478,N_13492);
or U13699 (N_13699,N_13491,N_13522);
nor U13700 (N_13700,N_13540,N_13460);
or U13701 (N_13701,N_13525,N_13595);
nand U13702 (N_13702,N_13533,N_13512);
xor U13703 (N_13703,N_13444,N_13574);
and U13704 (N_13704,N_13535,N_13550);
or U13705 (N_13705,N_13494,N_13581);
xor U13706 (N_13706,N_13530,N_13498);
and U13707 (N_13707,N_13584,N_13454);
and U13708 (N_13708,N_13497,N_13508);
nor U13709 (N_13709,N_13459,N_13511);
or U13710 (N_13710,N_13586,N_13511);
nor U13711 (N_13711,N_13519,N_13581);
xor U13712 (N_13712,N_13456,N_13580);
xnor U13713 (N_13713,N_13510,N_13562);
and U13714 (N_13714,N_13544,N_13472);
and U13715 (N_13715,N_13521,N_13590);
and U13716 (N_13716,N_13543,N_13522);
and U13717 (N_13717,N_13506,N_13564);
or U13718 (N_13718,N_13440,N_13501);
nand U13719 (N_13719,N_13485,N_13529);
nand U13720 (N_13720,N_13492,N_13594);
xnor U13721 (N_13721,N_13454,N_13504);
or U13722 (N_13722,N_13532,N_13487);
nor U13723 (N_13723,N_13501,N_13445);
xor U13724 (N_13724,N_13492,N_13510);
and U13725 (N_13725,N_13466,N_13596);
and U13726 (N_13726,N_13508,N_13555);
xnor U13727 (N_13727,N_13524,N_13571);
nand U13728 (N_13728,N_13462,N_13489);
xnor U13729 (N_13729,N_13564,N_13534);
and U13730 (N_13730,N_13578,N_13550);
and U13731 (N_13731,N_13589,N_13509);
nor U13732 (N_13732,N_13587,N_13480);
and U13733 (N_13733,N_13569,N_13497);
xor U13734 (N_13734,N_13483,N_13507);
or U13735 (N_13735,N_13499,N_13488);
and U13736 (N_13736,N_13543,N_13491);
nand U13737 (N_13737,N_13520,N_13464);
or U13738 (N_13738,N_13526,N_13529);
nor U13739 (N_13739,N_13527,N_13473);
and U13740 (N_13740,N_13481,N_13544);
nor U13741 (N_13741,N_13567,N_13501);
xnor U13742 (N_13742,N_13544,N_13546);
xor U13743 (N_13743,N_13461,N_13563);
or U13744 (N_13744,N_13466,N_13526);
or U13745 (N_13745,N_13524,N_13444);
nor U13746 (N_13746,N_13481,N_13503);
and U13747 (N_13747,N_13447,N_13527);
nor U13748 (N_13748,N_13446,N_13497);
xnor U13749 (N_13749,N_13570,N_13443);
nand U13750 (N_13750,N_13465,N_13504);
nor U13751 (N_13751,N_13455,N_13450);
and U13752 (N_13752,N_13521,N_13480);
xnor U13753 (N_13753,N_13547,N_13472);
nand U13754 (N_13754,N_13478,N_13450);
nand U13755 (N_13755,N_13550,N_13494);
xor U13756 (N_13756,N_13595,N_13550);
nand U13757 (N_13757,N_13453,N_13447);
nand U13758 (N_13758,N_13452,N_13562);
or U13759 (N_13759,N_13594,N_13578);
or U13760 (N_13760,N_13679,N_13606);
or U13761 (N_13761,N_13618,N_13654);
xnor U13762 (N_13762,N_13633,N_13600);
nand U13763 (N_13763,N_13673,N_13615);
and U13764 (N_13764,N_13689,N_13655);
nand U13765 (N_13765,N_13639,N_13665);
or U13766 (N_13766,N_13701,N_13660);
xnor U13767 (N_13767,N_13629,N_13626);
or U13768 (N_13768,N_13616,N_13674);
and U13769 (N_13769,N_13641,N_13631);
or U13770 (N_13770,N_13707,N_13727);
xnor U13771 (N_13771,N_13695,N_13601);
and U13772 (N_13772,N_13603,N_13692);
xor U13773 (N_13773,N_13733,N_13656);
or U13774 (N_13774,N_13681,N_13716);
and U13775 (N_13775,N_13737,N_13619);
nand U13776 (N_13776,N_13649,N_13685);
nor U13777 (N_13777,N_13643,N_13604);
and U13778 (N_13778,N_13676,N_13613);
nand U13779 (N_13779,N_13635,N_13640);
nor U13780 (N_13780,N_13696,N_13688);
nor U13781 (N_13781,N_13697,N_13678);
nand U13782 (N_13782,N_13743,N_13651);
or U13783 (N_13783,N_13636,N_13672);
nor U13784 (N_13784,N_13622,N_13637);
and U13785 (N_13785,N_13617,N_13721);
or U13786 (N_13786,N_13624,N_13730);
or U13787 (N_13787,N_13757,N_13632);
nand U13788 (N_13788,N_13722,N_13715);
xor U13789 (N_13789,N_13608,N_13659);
nand U13790 (N_13790,N_13759,N_13713);
and U13791 (N_13791,N_13718,N_13740);
xor U13792 (N_13792,N_13677,N_13675);
xor U13793 (N_13793,N_13751,N_13682);
xnor U13794 (N_13794,N_13704,N_13712);
and U13795 (N_13795,N_13736,N_13700);
nand U13796 (N_13796,N_13642,N_13714);
and U13797 (N_13797,N_13705,N_13666);
or U13798 (N_13798,N_13630,N_13691);
xor U13799 (N_13799,N_13670,N_13747);
nand U13800 (N_13800,N_13621,N_13738);
or U13801 (N_13801,N_13711,N_13647);
xnor U13802 (N_13802,N_13687,N_13758);
nor U13803 (N_13803,N_13607,N_13653);
nand U13804 (N_13804,N_13690,N_13752);
or U13805 (N_13805,N_13708,N_13650);
nand U13806 (N_13806,N_13703,N_13749);
nand U13807 (N_13807,N_13748,N_13699);
nor U13808 (N_13808,N_13669,N_13694);
or U13809 (N_13809,N_13735,N_13750);
nor U13810 (N_13810,N_13661,N_13657);
nor U13811 (N_13811,N_13734,N_13627);
or U13812 (N_13812,N_13709,N_13753);
and U13813 (N_13813,N_13628,N_13684);
or U13814 (N_13814,N_13664,N_13724);
nor U13815 (N_13815,N_13741,N_13754);
or U13816 (N_13816,N_13732,N_13645);
xor U13817 (N_13817,N_13731,N_13698);
xnor U13818 (N_13818,N_13693,N_13742);
xnor U13819 (N_13819,N_13725,N_13623);
or U13820 (N_13820,N_13620,N_13683);
or U13821 (N_13821,N_13611,N_13671);
or U13822 (N_13822,N_13625,N_13638);
xnor U13823 (N_13823,N_13663,N_13720);
or U13824 (N_13824,N_13667,N_13602);
nor U13825 (N_13825,N_13755,N_13723);
and U13826 (N_13826,N_13680,N_13729);
nand U13827 (N_13827,N_13745,N_13686);
or U13828 (N_13828,N_13614,N_13739);
xor U13829 (N_13829,N_13746,N_13652);
and U13830 (N_13830,N_13612,N_13756);
or U13831 (N_13831,N_13610,N_13605);
nor U13832 (N_13832,N_13662,N_13744);
xor U13833 (N_13833,N_13710,N_13726);
xor U13834 (N_13834,N_13609,N_13702);
nand U13835 (N_13835,N_13706,N_13658);
and U13836 (N_13836,N_13728,N_13648);
or U13837 (N_13837,N_13646,N_13634);
or U13838 (N_13838,N_13668,N_13644);
nor U13839 (N_13839,N_13717,N_13719);
xor U13840 (N_13840,N_13749,N_13651);
nand U13841 (N_13841,N_13669,N_13662);
nand U13842 (N_13842,N_13657,N_13724);
nand U13843 (N_13843,N_13759,N_13749);
xnor U13844 (N_13844,N_13692,N_13606);
or U13845 (N_13845,N_13676,N_13681);
and U13846 (N_13846,N_13662,N_13613);
or U13847 (N_13847,N_13757,N_13750);
xnor U13848 (N_13848,N_13703,N_13641);
or U13849 (N_13849,N_13744,N_13678);
or U13850 (N_13850,N_13646,N_13630);
or U13851 (N_13851,N_13724,N_13645);
or U13852 (N_13852,N_13709,N_13633);
or U13853 (N_13853,N_13748,N_13661);
xnor U13854 (N_13854,N_13602,N_13710);
and U13855 (N_13855,N_13686,N_13611);
nand U13856 (N_13856,N_13696,N_13610);
nand U13857 (N_13857,N_13629,N_13752);
nor U13858 (N_13858,N_13726,N_13648);
nand U13859 (N_13859,N_13643,N_13743);
xnor U13860 (N_13860,N_13691,N_13654);
xor U13861 (N_13861,N_13735,N_13699);
nor U13862 (N_13862,N_13664,N_13620);
and U13863 (N_13863,N_13722,N_13671);
nand U13864 (N_13864,N_13744,N_13693);
or U13865 (N_13865,N_13686,N_13730);
nor U13866 (N_13866,N_13736,N_13749);
nor U13867 (N_13867,N_13651,N_13691);
nor U13868 (N_13868,N_13667,N_13651);
or U13869 (N_13869,N_13661,N_13751);
and U13870 (N_13870,N_13693,N_13749);
nor U13871 (N_13871,N_13661,N_13667);
xnor U13872 (N_13872,N_13753,N_13644);
nand U13873 (N_13873,N_13605,N_13718);
xor U13874 (N_13874,N_13658,N_13613);
and U13875 (N_13875,N_13714,N_13653);
and U13876 (N_13876,N_13744,N_13754);
nand U13877 (N_13877,N_13618,N_13682);
xor U13878 (N_13878,N_13621,N_13706);
nand U13879 (N_13879,N_13706,N_13678);
nand U13880 (N_13880,N_13636,N_13735);
or U13881 (N_13881,N_13654,N_13625);
and U13882 (N_13882,N_13637,N_13745);
or U13883 (N_13883,N_13644,N_13695);
nand U13884 (N_13884,N_13756,N_13749);
nand U13885 (N_13885,N_13709,N_13675);
nor U13886 (N_13886,N_13668,N_13624);
and U13887 (N_13887,N_13694,N_13610);
nor U13888 (N_13888,N_13742,N_13757);
xor U13889 (N_13889,N_13688,N_13739);
xnor U13890 (N_13890,N_13682,N_13741);
nor U13891 (N_13891,N_13717,N_13731);
nand U13892 (N_13892,N_13603,N_13681);
or U13893 (N_13893,N_13706,N_13616);
and U13894 (N_13894,N_13722,N_13673);
or U13895 (N_13895,N_13604,N_13681);
xnor U13896 (N_13896,N_13699,N_13647);
nand U13897 (N_13897,N_13625,N_13741);
or U13898 (N_13898,N_13608,N_13750);
xor U13899 (N_13899,N_13717,N_13716);
and U13900 (N_13900,N_13709,N_13638);
or U13901 (N_13901,N_13625,N_13663);
xor U13902 (N_13902,N_13644,N_13721);
or U13903 (N_13903,N_13627,N_13713);
nor U13904 (N_13904,N_13753,N_13694);
or U13905 (N_13905,N_13693,N_13732);
and U13906 (N_13906,N_13725,N_13753);
and U13907 (N_13907,N_13621,N_13689);
and U13908 (N_13908,N_13741,N_13746);
nor U13909 (N_13909,N_13670,N_13676);
xor U13910 (N_13910,N_13709,N_13738);
xor U13911 (N_13911,N_13729,N_13685);
nand U13912 (N_13912,N_13610,N_13751);
nor U13913 (N_13913,N_13680,N_13713);
xor U13914 (N_13914,N_13636,N_13678);
and U13915 (N_13915,N_13664,N_13618);
or U13916 (N_13916,N_13727,N_13750);
nand U13917 (N_13917,N_13640,N_13649);
xnor U13918 (N_13918,N_13674,N_13602);
and U13919 (N_13919,N_13640,N_13687);
and U13920 (N_13920,N_13838,N_13814);
nor U13921 (N_13921,N_13798,N_13876);
and U13922 (N_13922,N_13856,N_13914);
nand U13923 (N_13923,N_13913,N_13895);
xnor U13924 (N_13924,N_13848,N_13863);
nor U13925 (N_13925,N_13894,N_13802);
and U13926 (N_13926,N_13785,N_13845);
or U13927 (N_13927,N_13760,N_13796);
nand U13928 (N_13928,N_13779,N_13772);
or U13929 (N_13929,N_13824,N_13882);
and U13930 (N_13930,N_13763,N_13832);
or U13931 (N_13931,N_13765,N_13872);
nand U13932 (N_13932,N_13778,N_13771);
or U13933 (N_13933,N_13819,N_13790);
xnor U13934 (N_13934,N_13868,N_13853);
and U13935 (N_13935,N_13918,N_13858);
and U13936 (N_13936,N_13817,N_13829);
nor U13937 (N_13937,N_13855,N_13880);
and U13938 (N_13938,N_13906,N_13916);
nor U13939 (N_13939,N_13823,N_13812);
and U13940 (N_13940,N_13818,N_13892);
or U13941 (N_13941,N_13775,N_13762);
xnor U13942 (N_13942,N_13810,N_13777);
and U13943 (N_13943,N_13839,N_13786);
xnor U13944 (N_13944,N_13893,N_13837);
or U13945 (N_13945,N_13830,N_13862);
or U13946 (N_13946,N_13891,N_13794);
xor U13947 (N_13947,N_13865,N_13854);
and U13948 (N_13948,N_13773,N_13846);
and U13949 (N_13949,N_13903,N_13805);
and U13950 (N_13950,N_13799,N_13890);
nand U13951 (N_13951,N_13813,N_13870);
nor U13952 (N_13952,N_13770,N_13831);
xnor U13953 (N_13953,N_13902,N_13769);
nor U13954 (N_13954,N_13800,N_13761);
or U13955 (N_13955,N_13889,N_13843);
xnor U13956 (N_13956,N_13833,N_13788);
nand U13957 (N_13957,N_13907,N_13910);
or U13958 (N_13958,N_13820,N_13791);
xnor U13959 (N_13959,N_13766,N_13919);
and U13960 (N_13960,N_13896,N_13825);
and U13961 (N_13961,N_13912,N_13797);
nor U13962 (N_13962,N_13901,N_13908);
xnor U13963 (N_13963,N_13809,N_13764);
or U13964 (N_13964,N_13873,N_13789);
and U13965 (N_13965,N_13849,N_13821);
nand U13966 (N_13966,N_13808,N_13864);
nor U13967 (N_13967,N_13780,N_13888);
or U13968 (N_13968,N_13816,N_13822);
and U13969 (N_13969,N_13878,N_13861);
xor U13970 (N_13970,N_13904,N_13776);
or U13971 (N_13971,N_13915,N_13857);
and U13972 (N_13972,N_13840,N_13806);
and U13973 (N_13973,N_13875,N_13917);
nand U13974 (N_13974,N_13782,N_13911);
or U13975 (N_13975,N_13866,N_13909);
nand U13976 (N_13976,N_13774,N_13815);
nand U13977 (N_13977,N_13851,N_13844);
or U13978 (N_13978,N_13898,N_13807);
nor U13979 (N_13979,N_13850,N_13859);
or U13980 (N_13980,N_13869,N_13836);
nor U13981 (N_13981,N_13884,N_13781);
nor U13982 (N_13982,N_13900,N_13828);
and U13983 (N_13983,N_13834,N_13887);
nand U13984 (N_13984,N_13811,N_13767);
nand U13985 (N_13985,N_13877,N_13827);
nand U13986 (N_13986,N_13871,N_13842);
nand U13987 (N_13987,N_13803,N_13768);
nand U13988 (N_13988,N_13835,N_13801);
nand U13989 (N_13989,N_13784,N_13795);
or U13990 (N_13990,N_13787,N_13852);
xor U13991 (N_13991,N_13783,N_13897);
and U13992 (N_13992,N_13826,N_13867);
xor U13993 (N_13993,N_13886,N_13899);
xnor U13994 (N_13994,N_13804,N_13847);
xor U13995 (N_13995,N_13793,N_13905);
and U13996 (N_13996,N_13881,N_13883);
nand U13997 (N_13997,N_13860,N_13874);
and U13998 (N_13998,N_13885,N_13879);
and U13999 (N_13999,N_13841,N_13792);
and U14000 (N_14000,N_13858,N_13821);
or U14001 (N_14001,N_13868,N_13850);
xnor U14002 (N_14002,N_13841,N_13849);
or U14003 (N_14003,N_13830,N_13854);
nor U14004 (N_14004,N_13856,N_13904);
nand U14005 (N_14005,N_13874,N_13866);
xor U14006 (N_14006,N_13782,N_13820);
or U14007 (N_14007,N_13828,N_13795);
xor U14008 (N_14008,N_13908,N_13774);
nand U14009 (N_14009,N_13906,N_13794);
xnor U14010 (N_14010,N_13879,N_13912);
and U14011 (N_14011,N_13896,N_13878);
or U14012 (N_14012,N_13793,N_13868);
and U14013 (N_14013,N_13887,N_13910);
and U14014 (N_14014,N_13911,N_13903);
or U14015 (N_14015,N_13814,N_13773);
nor U14016 (N_14016,N_13850,N_13761);
or U14017 (N_14017,N_13871,N_13905);
nor U14018 (N_14018,N_13893,N_13827);
or U14019 (N_14019,N_13852,N_13912);
or U14020 (N_14020,N_13883,N_13900);
nor U14021 (N_14021,N_13891,N_13767);
and U14022 (N_14022,N_13785,N_13899);
xor U14023 (N_14023,N_13807,N_13881);
or U14024 (N_14024,N_13800,N_13840);
or U14025 (N_14025,N_13888,N_13869);
and U14026 (N_14026,N_13773,N_13836);
nor U14027 (N_14027,N_13840,N_13803);
and U14028 (N_14028,N_13760,N_13870);
and U14029 (N_14029,N_13793,N_13775);
xor U14030 (N_14030,N_13781,N_13806);
nand U14031 (N_14031,N_13801,N_13843);
and U14032 (N_14032,N_13810,N_13869);
and U14033 (N_14033,N_13799,N_13878);
nor U14034 (N_14034,N_13829,N_13851);
nand U14035 (N_14035,N_13760,N_13858);
or U14036 (N_14036,N_13859,N_13897);
or U14037 (N_14037,N_13892,N_13845);
and U14038 (N_14038,N_13768,N_13884);
or U14039 (N_14039,N_13854,N_13847);
nand U14040 (N_14040,N_13898,N_13860);
nor U14041 (N_14041,N_13815,N_13837);
or U14042 (N_14042,N_13868,N_13894);
and U14043 (N_14043,N_13809,N_13858);
nor U14044 (N_14044,N_13858,N_13903);
nand U14045 (N_14045,N_13778,N_13761);
xnor U14046 (N_14046,N_13885,N_13815);
or U14047 (N_14047,N_13911,N_13905);
nor U14048 (N_14048,N_13777,N_13772);
xnor U14049 (N_14049,N_13805,N_13787);
nor U14050 (N_14050,N_13916,N_13808);
nor U14051 (N_14051,N_13857,N_13867);
xnor U14052 (N_14052,N_13778,N_13770);
or U14053 (N_14053,N_13892,N_13899);
nand U14054 (N_14054,N_13904,N_13779);
and U14055 (N_14055,N_13880,N_13801);
nor U14056 (N_14056,N_13808,N_13863);
and U14057 (N_14057,N_13819,N_13914);
or U14058 (N_14058,N_13762,N_13799);
or U14059 (N_14059,N_13816,N_13786);
or U14060 (N_14060,N_13788,N_13870);
xnor U14061 (N_14061,N_13803,N_13865);
xnor U14062 (N_14062,N_13887,N_13821);
nand U14063 (N_14063,N_13886,N_13868);
and U14064 (N_14064,N_13876,N_13763);
nand U14065 (N_14065,N_13887,N_13827);
or U14066 (N_14066,N_13860,N_13895);
xnor U14067 (N_14067,N_13886,N_13880);
and U14068 (N_14068,N_13852,N_13854);
nor U14069 (N_14069,N_13865,N_13796);
and U14070 (N_14070,N_13804,N_13892);
nand U14071 (N_14071,N_13793,N_13897);
nand U14072 (N_14072,N_13861,N_13779);
or U14073 (N_14073,N_13912,N_13771);
xnor U14074 (N_14074,N_13828,N_13792);
xnor U14075 (N_14075,N_13876,N_13850);
and U14076 (N_14076,N_13806,N_13771);
and U14077 (N_14077,N_13804,N_13772);
or U14078 (N_14078,N_13812,N_13810);
nand U14079 (N_14079,N_13792,N_13887);
or U14080 (N_14080,N_14067,N_13927);
nand U14081 (N_14081,N_14000,N_13994);
nand U14082 (N_14082,N_13965,N_13940);
nor U14083 (N_14083,N_14031,N_13976);
nor U14084 (N_14084,N_14052,N_14035);
nor U14085 (N_14085,N_13921,N_13939);
nand U14086 (N_14086,N_14071,N_14012);
nand U14087 (N_14087,N_14019,N_14045);
nor U14088 (N_14088,N_14048,N_14064);
or U14089 (N_14089,N_13999,N_13993);
xor U14090 (N_14090,N_14002,N_13925);
and U14091 (N_14091,N_13978,N_13952);
xor U14092 (N_14092,N_14046,N_13975);
nand U14093 (N_14093,N_14021,N_13946);
nor U14094 (N_14094,N_13937,N_13989);
nor U14095 (N_14095,N_13980,N_13922);
or U14096 (N_14096,N_14077,N_13968);
xor U14097 (N_14097,N_13967,N_13941);
nand U14098 (N_14098,N_14005,N_14009);
or U14099 (N_14099,N_13935,N_14018);
nand U14100 (N_14100,N_13987,N_14032);
nor U14101 (N_14101,N_13972,N_13926);
nand U14102 (N_14102,N_13961,N_14008);
or U14103 (N_14103,N_13981,N_14059);
nor U14104 (N_14104,N_13950,N_14078);
xnor U14105 (N_14105,N_14073,N_13996);
or U14106 (N_14106,N_13948,N_14042);
and U14107 (N_14107,N_14044,N_13990);
or U14108 (N_14108,N_14007,N_13962);
nor U14109 (N_14109,N_14070,N_14039);
nand U14110 (N_14110,N_14013,N_13997);
or U14111 (N_14111,N_14010,N_13988);
or U14112 (N_14112,N_13932,N_13957);
or U14113 (N_14113,N_13938,N_14043);
nand U14114 (N_14114,N_14036,N_14079);
nor U14115 (N_14115,N_13963,N_13929);
and U14116 (N_14116,N_13974,N_13959);
or U14117 (N_14117,N_13953,N_13979);
xor U14118 (N_14118,N_14072,N_13956);
and U14119 (N_14119,N_14037,N_13995);
or U14120 (N_14120,N_14056,N_13966);
and U14121 (N_14121,N_14029,N_13943);
nand U14122 (N_14122,N_14028,N_14017);
nor U14123 (N_14123,N_14057,N_14047);
or U14124 (N_14124,N_14076,N_14055);
nand U14125 (N_14125,N_14023,N_13977);
nor U14126 (N_14126,N_13924,N_13984);
nand U14127 (N_14127,N_13960,N_14058);
nand U14128 (N_14128,N_13973,N_14040);
or U14129 (N_14129,N_14015,N_14068);
and U14130 (N_14130,N_13991,N_14034);
and U14131 (N_14131,N_13969,N_13934);
nand U14132 (N_14132,N_14030,N_14027);
xnor U14133 (N_14133,N_14016,N_14014);
nand U14134 (N_14134,N_14011,N_13923);
and U14135 (N_14135,N_14075,N_13928);
and U14136 (N_14136,N_13986,N_13982);
nand U14137 (N_14137,N_14069,N_14022);
nand U14138 (N_14138,N_14001,N_14025);
xnor U14139 (N_14139,N_13944,N_14038);
xor U14140 (N_14140,N_14003,N_13958);
or U14141 (N_14141,N_14065,N_14024);
and U14142 (N_14142,N_13992,N_13971);
xnor U14143 (N_14143,N_13955,N_14051);
or U14144 (N_14144,N_13998,N_14061);
nor U14145 (N_14145,N_14041,N_13964);
or U14146 (N_14146,N_13920,N_14033);
nand U14147 (N_14147,N_14054,N_14074);
xnor U14148 (N_14148,N_14062,N_13949);
xnor U14149 (N_14149,N_14053,N_13942);
xnor U14150 (N_14150,N_14020,N_13945);
or U14151 (N_14151,N_13931,N_13985);
nor U14152 (N_14152,N_13930,N_13983);
or U14153 (N_14153,N_13951,N_14049);
xor U14154 (N_14154,N_14060,N_14004);
nand U14155 (N_14155,N_13936,N_13970);
and U14156 (N_14156,N_13954,N_14026);
xnor U14157 (N_14157,N_13933,N_14006);
nand U14158 (N_14158,N_13947,N_14066);
nand U14159 (N_14159,N_14063,N_14050);
nor U14160 (N_14160,N_13986,N_14004);
or U14161 (N_14161,N_14061,N_14064);
and U14162 (N_14162,N_14024,N_13982);
nand U14163 (N_14163,N_13994,N_14072);
nand U14164 (N_14164,N_14016,N_13943);
xnor U14165 (N_14165,N_14010,N_13952);
xnor U14166 (N_14166,N_13989,N_13994);
nor U14167 (N_14167,N_14037,N_14051);
nor U14168 (N_14168,N_14061,N_14052);
xor U14169 (N_14169,N_14030,N_13944);
or U14170 (N_14170,N_13948,N_13995);
nor U14171 (N_14171,N_14013,N_13946);
nand U14172 (N_14172,N_14023,N_14059);
and U14173 (N_14173,N_14072,N_14059);
nor U14174 (N_14174,N_13948,N_14065);
nor U14175 (N_14175,N_14015,N_13934);
or U14176 (N_14176,N_14031,N_14011);
xnor U14177 (N_14177,N_13999,N_14038);
nand U14178 (N_14178,N_14037,N_13968);
and U14179 (N_14179,N_14012,N_14028);
nor U14180 (N_14180,N_14051,N_14062);
nand U14181 (N_14181,N_13984,N_13957);
nor U14182 (N_14182,N_13995,N_13984);
nor U14183 (N_14183,N_14010,N_13962);
or U14184 (N_14184,N_13983,N_13998);
and U14185 (N_14185,N_13987,N_14015);
nor U14186 (N_14186,N_14034,N_14041);
or U14187 (N_14187,N_13991,N_13946);
nand U14188 (N_14188,N_13929,N_14064);
or U14189 (N_14189,N_14049,N_13938);
xor U14190 (N_14190,N_13935,N_13968);
nor U14191 (N_14191,N_13976,N_14023);
and U14192 (N_14192,N_13988,N_13999);
nand U14193 (N_14193,N_14026,N_13948);
nand U14194 (N_14194,N_13972,N_13960);
or U14195 (N_14195,N_14041,N_13984);
nor U14196 (N_14196,N_13963,N_14031);
nand U14197 (N_14197,N_13954,N_14048);
and U14198 (N_14198,N_14012,N_13930);
xor U14199 (N_14199,N_13943,N_13941);
xnor U14200 (N_14200,N_14014,N_14022);
nor U14201 (N_14201,N_14052,N_14079);
nor U14202 (N_14202,N_14000,N_14013);
xor U14203 (N_14203,N_13933,N_13927);
xnor U14204 (N_14204,N_13930,N_14068);
xnor U14205 (N_14205,N_14079,N_14046);
and U14206 (N_14206,N_14061,N_13993);
nand U14207 (N_14207,N_14037,N_14042);
nor U14208 (N_14208,N_13968,N_13952);
nand U14209 (N_14209,N_14060,N_13929);
xnor U14210 (N_14210,N_14004,N_13987);
or U14211 (N_14211,N_13996,N_13962);
nand U14212 (N_14212,N_14071,N_14049);
nand U14213 (N_14213,N_13986,N_13965);
xor U14214 (N_14214,N_14010,N_14074);
and U14215 (N_14215,N_14023,N_14039);
xor U14216 (N_14216,N_13945,N_13977);
and U14217 (N_14217,N_13992,N_13952);
and U14218 (N_14218,N_13951,N_14053);
nor U14219 (N_14219,N_13955,N_14031);
xnor U14220 (N_14220,N_13987,N_13957);
or U14221 (N_14221,N_14063,N_13954);
or U14222 (N_14222,N_14037,N_13966);
xor U14223 (N_14223,N_13926,N_14054);
nand U14224 (N_14224,N_13991,N_14052);
nand U14225 (N_14225,N_13929,N_14065);
nor U14226 (N_14226,N_13975,N_13977);
and U14227 (N_14227,N_14004,N_14018);
nand U14228 (N_14228,N_13972,N_14050);
nand U14229 (N_14229,N_14075,N_14037);
and U14230 (N_14230,N_13928,N_14010);
and U14231 (N_14231,N_13970,N_14041);
xnor U14232 (N_14232,N_14076,N_13949);
nand U14233 (N_14233,N_13957,N_14025);
or U14234 (N_14234,N_14003,N_13934);
nor U14235 (N_14235,N_13975,N_13970);
or U14236 (N_14236,N_14050,N_13961);
or U14237 (N_14237,N_14027,N_13973);
nor U14238 (N_14238,N_13942,N_14013);
xor U14239 (N_14239,N_14071,N_14013);
and U14240 (N_14240,N_14202,N_14205);
nand U14241 (N_14241,N_14192,N_14132);
nand U14242 (N_14242,N_14081,N_14218);
and U14243 (N_14243,N_14152,N_14164);
nand U14244 (N_14244,N_14217,N_14210);
or U14245 (N_14245,N_14147,N_14177);
xnor U14246 (N_14246,N_14095,N_14123);
xor U14247 (N_14247,N_14106,N_14102);
nand U14248 (N_14248,N_14206,N_14116);
xnor U14249 (N_14249,N_14150,N_14110);
nor U14250 (N_14250,N_14109,N_14093);
nor U14251 (N_14251,N_14124,N_14238);
nor U14252 (N_14252,N_14134,N_14101);
and U14253 (N_14253,N_14234,N_14149);
and U14254 (N_14254,N_14175,N_14163);
xor U14255 (N_14255,N_14105,N_14138);
xnor U14256 (N_14256,N_14153,N_14199);
nand U14257 (N_14257,N_14173,N_14085);
nand U14258 (N_14258,N_14161,N_14215);
nor U14259 (N_14259,N_14211,N_14219);
or U14260 (N_14260,N_14151,N_14193);
and U14261 (N_14261,N_14100,N_14168);
xor U14262 (N_14262,N_14127,N_14137);
and U14263 (N_14263,N_14170,N_14144);
nor U14264 (N_14264,N_14082,N_14089);
nand U14265 (N_14265,N_14112,N_14117);
nor U14266 (N_14266,N_14115,N_14207);
xor U14267 (N_14267,N_14203,N_14120);
xnor U14268 (N_14268,N_14197,N_14086);
and U14269 (N_14269,N_14183,N_14119);
xor U14270 (N_14270,N_14209,N_14200);
xnor U14271 (N_14271,N_14181,N_14179);
and U14272 (N_14272,N_14180,N_14114);
nand U14273 (N_14273,N_14186,N_14204);
and U14274 (N_14274,N_14226,N_14122);
and U14275 (N_14275,N_14195,N_14229);
xnor U14276 (N_14276,N_14140,N_14104);
xor U14277 (N_14277,N_14220,N_14098);
xor U14278 (N_14278,N_14131,N_14190);
xor U14279 (N_14279,N_14133,N_14191);
and U14280 (N_14280,N_14188,N_14142);
nor U14281 (N_14281,N_14158,N_14182);
nand U14282 (N_14282,N_14231,N_14230);
or U14283 (N_14283,N_14233,N_14194);
nor U14284 (N_14284,N_14185,N_14216);
or U14285 (N_14285,N_14108,N_14171);
nor U14286 (N_14286,N_14232,N_14237);
nand U14287 (N_14287,N_14222,N_14162);
nor U14288 (N_14288,N_14166,N_14097);
nor U14289 (N_14289,N_14224,N_14136);
nor U14290 (N_14290,N_14198,N_14084);
or U14291 (N_14291,N_14223,N_14139);
and U14292 (N_14292,N_14225,N_14184);
or U14293 (N_14293,N_14094,N_14169);
xnor U14294 (N_14294,N_14091,N_14239);
and U14295 (N_14295,N_14107,N_14178);
nor U14296 (N_14296,N_14128,N_14145);
xnor U14297 (N_14297,N_14141,N_14148);
or U14298 (N_14298,N_14214,N_14213);
or U14299 (N_14299,N_14189,N_14146);
or U14300 (N_14300,N_14208,N_14159);
and U14301 (N_14301,N_14099,N_14167);
or U14302 (N_14302,N_14235,N_14157);
xor U14303 (N_14303,N_14111,N_14135);
nand U14304 (N_14304,N_14090,N_14092);
nand U14305 (N_14305,N_14236,N_14129);
xor U14306 (N_14306,N_14156,N_14196);
xor U14307 (N_14307,N_14103,N_14155);
nor U14308 (N_14308,N_14228,N_14174);
and U14309 (N_14309,N_14121,N_14212);
and U14310 (N_14310,N_14083,N_14088);
xnor U14311 (N_14311,N_14165,N_14126);
nand U14312 (N_14312,N_14087,N_14154);
and U14313 (N_14313,N_14201,N_14080);
nand U14314 (N_14314,N_14125,N_14113);
nor U14315 (N_14315,N_14187,N_14176);
or U14316 (N_14316,N_14160,N_14227);
nand U14317 (N_14317,N_14221,N_14172);
xnor U14318 (N_14318,N_14118,N_14096);
nand U14319 (N_14319,N_14143,N_14130);
nand U14320 (N_14320,N_14174,N_14156);
xor U14321 (N_14321,N_14153,N_14090);
nand U14322 (N_14322,N_14113,N_14215);
nand U14323 (N_14323,N_14159,N_14168);
xnor U14324 (N_14324,N_14120,N_14098);
nand U14325 (N_14325,N_14096,N_14167);
nand U14326 (N_14326,N_14094,N_14173);
or U14327 (N_14327,N_14095,N_14156);
and U14328 (N_14328,N_14135,N_14167);
nand U14329 (N_14329,N_14087,N_14094);
and U14330 (N_14330,N_14155,N_14113);
and U14331 (N_14331,N_14119,N_14130);
nor U14332 (N_14332,N_14155,N_14089);
nand U14333 (N_14333,N_14091,N_14211);
nand U14334 (N_14334,N_14128,N_14209);
xor U14335 (N_14335,N_14130,N_14239);
xnor U14336 (N_14336,N_14088,N_14174);
nor U14337 (N_14337,N_14197,N_14192);
and U14338 (N_14338,N_14209,N_14140);
nand U14339 (N_14339,N_14191,N_14110);
xor U14340 (N_14340,N_14089,N_14112);
xor U14341 (N_14341,N_14128,N_14213);
nand U14342 (N_14342,N_14158,N_14220);
nor U14343 (N_14343,N_14104,N_14086);
or U14344 (N_14344,N_14206,N_14161);
xnor U14345 (N_14345,N_14149,N_14238);
and U14346 (N_14346,N_14198,N_14129);
nand U14347 (N_14347,N_14230,N_14193);
nor U14348 (N_14348,N_14167,N_14129);
nand U14349 (N_14349,N_14176,N_14169);
nor U14350 (N_14350,N_14182,N_14157);
and U14351 (N_14351,N_14170,N_14205);
and U14352 (N_14352,N_14170,N_14115);
and U14353 (N_14353,N_14189,N_14117);
or U14354 (N_14354,N_14189,N_14226);
nor U14355 (N_14355,N_14236,N_14103);
xor U14356 (N_14356,N_14177,N_14135);
nor U14357 (N_14357,N_14202,N_14114);
or U14358 (N_14358,N_14170,N_14176);
or U14359 (N_14359,N_14230,N_14133);
and U14360 (N_14360,N_14084,N_14144);
nor U14361 (N_14361,N_14080,N_14169);
xnor U14362 (N_14362,N_14093,N_14172);
nor U14363 (N_14363,N_14122,N_14085);
nand U14364 (N_14364,N_14146,N_14201);
or U14365 (N_14365,N_14199,N_14141);
nand U14366 (N_14366,N_14179,N_14235);
nand U14367 (N_14367,N_14115,N_14191);
nor U14368 (N_14368,N_14124,N_14151);
and U14369 (N_14369,N_14233,N_14084);
nand U14370 (N_14370,N_14193,N_14185);
xnor U14371 (N_14371,N_14124,N_14148);
or U14372 (N_14372,N_14119,N_14164);
xnor U14373 (N_14373,N_14088,N_14100);
and U14374 (N_14374,N_14197,N_14115);
xor U14375 (N_14375,N_14113,N_14114);
or U14376 (N_14376,N_14111,N_14210);
or U14377 (N_14377,N_14170,N_14193);
or U14378 (N_14378,N_14182,N_14231);
and U14379 (N_14379,N_14226,N_14237);
or U14380 (N_14380,N_14176,N_14147);
nand U14381 (N_14381,N_14197,N_14228);
nand U14382 (N_14382,N_14172,N_14234);
nand U14383 (N_14383,N_14130,N_14082);
or U14384 (N_14384,N_14097,N_14228);
or U14385 (N_14385,N_14227,N_14198);
or U14386 (N_14386,N_14092,N_14234);
nand U14387 (N_14387,N_14154,N_14203);
xor U14388 (N_14388,N_14093,N_14192);
or U14389 (N_14389,N_14232,N_14137);
or U14390 (N_14390,N_14126,N_14080);
xor U14391 (N_14391,N_14209,N_14113);
nand U14392 (N_14392,N_14220,N_14087);
xor U14393 (N_14393,N_14082,N_14191);
or U14394 (N_14394,N_14097,N_14164);
xor U14395 (N_14395,N_14095,N_14207);
xnor U14396 (N_14396,N_14218,N_14228);
nand U14397 (N_14397,N_14080,N_14152);
nand U14398 (N_14398,N_14158,N_14123);
or U14399 (N_14399,N_14122,N_14109);
nor U14400 (N_14400,N_14384,N_14355);
or U14401 (N_14401,N_14307,N_14255);
or U14402 (N_14402,N_14338,N_14347);
and U14403 (N_14403,N_14346,N_14391);
or U14404 (N_14404,N_14248,N_14301);
nand U14405 (N_14405,N_14393,N_14372);
or U14406 (N_14406,N_14265,N_14325);
or U14407 (N_14407,N_14277,N_14274);
nand U14408 (N_14408,N_14380,N_14327);
or U14409 (N_14409,N_14365,N_14382);
and U14410 (N_14410,N_14392,N_14354);
xor U14411 (N_14411,N_14398,N_14271);
and U14412 (N_14412,N_14242,N_14319);
nor U14413 (N_14413,N_14333,N_14348);
xor U14414 (N_14414,N_14304,N_14314);
xor U14415 (N_14415,N_14269,N_14373);
nor U14416 (N_14416,N_14290,N_14294);
nand U14417 (N_14417,N_14243,N_14310);
xnor U14418 (N_14418,N_14258,N_14303);
nand U14419 (N_14419,N_14262,N_14363);
or U14420 (N_14420,N_14247,N_14374);
nand U14421 (N_14421,N_14276,N_14289);
nand U14422 (N_14422,N_14273,N_14298);
or U14423 (N_14423,N_14279,N_14246);
or U14424 (N_14424,N_14287,N_14302);
or U14425 (N_14425,N_14379,N_14288);
xor U14426 (N_14426,N_14263,N_14281);
nand U14427 (N_14427,N_14335,N_14352);
and U14428 (N_14428,N_14337,N_14254);
or U14429 (N_14429,N_14369,N_14370);
and U14430 (N_14430,N_14377,N_14383);
nand U14431 (N_14431,N_14351,N_14359);
nand U14432 (N_14432,N_14245,N_14326);
and U14433 (N_14433,N_14394,N_14340);
nor U14434 (N_14434,N_14309,N_14322);
or U14435 (N_14435,N_14388,N_14341);
xnor U14436 (N_14436,N_14381,N_14299);
nand U14437 (N_14437,N_14390,N_14357);
nor U14438 (N_14438,N_14389,N_14280);
nand U14439 (N_14439,N_14285,N_14368);
nor U14440 (N_14440,N_14251,N_14378);
xnor U14441 (N_14441,N_14328,N_14249);
nand U14442 (N_14442,N_14244,N_14259);
nor U14443 (N_14443,N_14257,N_14356);
or U14444 (N_14444,N_14315,N_14344);
xnor U14445 (N_14445,N_14376,N_14358);
and U14446 (N_14446,N_14291,N_14343);
nand U14447 (N_14447,N_14366,N_14240);
nand U14448 (N_14448,N_14396,N_14308);
or U14449 (N_14449,N_14330,N_14399);
and U14450 (N_14450,N_14332,N_14349);
xor U14451 (N_14451,N_14286,N_14334);
or U14452 (N_14452,N_14283,N_14397);
xnor U14453 (N_14453,N_14305,N_14266);
nand U14454 (N_14454,N_14367,N_14360);
nor U14455 (N_14455,N_14264,N_14353);
xor U14456 (N_14456,N_14253,N_14272);
or U14457 (N_14457,N_14342,N_14267);
and U14458 (N_14458,N_14316,N_14278);
nand U14459 (N_14459,N_14261,N_14268);
nand U14460 (N_14460,N_14292,N_14284);
or U14461 (N_14461,N_14241,N_14295);
and U14462 (N_14462,N_14297,N_14345);
xor U14463 (N_14463,N_14260,N_14282);
nand U14464 (N_14464,N_14293,N_14323);
or U14465 (N_14465,N_14320,N_14321);
nor U14466 (N_14466,N_14312,N_14339);
and U14467 (N_14467,N_14306,N_14375);
and U14468 (N_14468,N_14386,N_14364);
xnor U14469 (N_14469,N_14256,N_14275);
xor U14470 (N_14470,N_14270,N_14252);
nor U14471 (N_14471,N_14324,N_14336);
nand U14472 (N_14472,N_14362,N_14296);
xnor U14473 (N_14473,N_14385,N_14371);
xor U14474 (N_14474,N_14311,N_14350);
nand U14475 (N_14475,N_14313,N_14317);
or U14476 (N_14476,N_14331,N_14361);
or U14477 (N_14477,N_14329,N_14395);
xor U14478 (N_14478,N_14300,N_14250);
and U14479 (N_14479,N_14318,N_14387);
nor U14480 (N_14480,N_14280,N_14352);
xnor U14481 (N_14481,N_14303,N_14364);
xor U14482 (N_14482,N_14354,N_14351);
nor U14483 (N_14483,N_14260,N_14241);
xnor U14484 (N_14484,N_14368,N_14394);
nand U14485 (N_14485,N_14370,N_14271);
nor U14486 (N_14486,N_14275,N_14365);
xnor U14487 (N_14487,N_14293,N_14398);
xnor U14488 (N_14488,N_14265,N_14350);
xnor U14489 (N_14489,N_14281,N_14369);
xor U14490 (N_14490,N_14249,N_14274);
and U14491 (N_14491,N_14359,N_14278);
nor U14492 (N_14492,N_14343,N_14295);
nor U14493 (N_14493,N_14351,N_14362);
and U14494 (N_14494,N_14266,N_14257);
or U14495 (N_14495,N_14257,N_14290);
nand U14496 (N_14496,N_14244,N_14398);
xor U14497 (N_14497,N_14280,N_14326);
nand U14498 (N_14498,N_14244,N_14282);
and U14499 (N_14499,N_14358,N_14364);
xor U14500 (N_14500,N_14287,N_14367);
or U14501 (N_14501,N_14346,N_14286);
nand U14502 (N_14502,N_14392,N_14358);
xor U14503 (N_14503,N_14349,N_14354);
or U14504 (N_14504,N_14376,N_14240);
or U14505 (N_14505,N_14332,N_14346);
and U14506 (N_14506,N_14324,N_14316);
nand U14507 (N_14507,N_14308,N_14394);
or U14508 (N_14508,N_14261,N_14281);
or U14509 (N_14509,N_14304,N_14358);
or U14510 (N_14510,N_14263,N_14350);
nand U14511 (N_14511,N_14340,N_14274);
xor U14512 (N_14512,N_14257,N_14352);
xnor U14513 (N_14513,N_14324,N_14303);
or U14514 (N_14514,N_14388,N_14328);
or U14515 (N_14515,N_14251,N_14246);
or U14516 (N_14516,N_14246,N_14366);
and U14517 (N_14517,N_14286,N_14385);
and U14518 (N_14518,N_14359,N_14258);
and U14519 (N_14519,N_14304,N_14320);
nor U14520 (N_14520,N_14386,N_14316);
and U14521 (N_14521,N_14364,N_14277);
xnor U14522 (N_14522,N_14360,N_14286);
nand U14523 (N_14523,N_14266,N_14383);
nor U14524 (N_14524,N_14304,N_14368);
nor U14525 (N_14525,N_14270,N_14353);
or U14526 (N_14526,N_14350,N_14330);
xnor U14527 (N_14527,N_14305,N_14372);
or U14528 (N_14528,N_14366,N_14245);
nor U14529 (N_14529,N_14361,N_14285);
nand U14530 (N_14530,N_14367,N_14378);
xnor U14531 (N_14531,N_14354,N_14346);
and U14532 (N_14532,N_14391,N_14352);
or U14533 (N_14533,N_14353,N_14245);
or U14534 (N_14534,N_14294,N_14347);
and U14535 (N_14535,N_14342,N_14319);
nand U14536 (N_14536,N_14277,N_14332);
nor U14537 (N_14537,N_14284,N_14326);
xnor U14538 (N_14538,N_14394,N_14301);
nand U14539 (N_14539,N_14255,N_14277);
and U14540 (N_14540,N_14346,N_14380);
and U14541 (N_14541,N_14327,N_14356);
or U14542 (N_14542,N_14398,N_14264);
nand U14543 (N_14543,N_14240,N_14377);
xor U14544 (N_14544,N_14240,N_14305);
nand U14545 (N_14545,N_14349,N_14367);
nor U14546 (N_14546,N_14321,N_14376);
xor U14547 (N_14547,N_14320,N_14353);
nor U14548 (N_14548,N_14257,N_14255);
and U14549 (N_14549,N_14318,N_14319);
nor U14550 (N_14550,N_14255,N_14299);
xnor U14551 (N_14551,N_14240,N_14242);
nand U14552 (N_14552,N_14247,N_14255);
nand U14553 (N_14553,N_14329,N_14260);
xor U14554 (N_14554,N_14294,N_14390);
xor U14555 (N_14555,N_14253,N_14375);
nand U14556 (N_14556,N_14360,N_14358);
nor U14557 (N_14557,N_14334,N_14345);
nand U14558 (N_14558,N_14379,N_14254);
xor U14559 (N_14559,N_14282,N_14249);
nand U14560 (N_14560,N_14439,N_14527);
nor U14561 (N_14561,N_14473,N_14438);
or U14562 (N_14562,N_14501,N_14521);
xnor U14563 (N_14563,N_14482,N_14461);
nand U14564 (N_14564,N_14445,N_14433);
or U14565 (N_14565,N_14477,N_14431);
or U14566 (N_14566,N_14426,N_14499);
xor U14567 (N_14567,N_14420,N_14494);
xnor U14568 (N_14568,N_14422,N_14467);
and U14569 (N_14569,N_14469,N_14486);
or U14570 (N_14570,N_14551,N_14429);
xnor U14571 (N_14571,N_14506,N_14530);
and U14572 (N_14572,N_14400,N_14522);
and U14573 (N_14573,N_14479,N_14538);
nor U14574 (N_14574,N_14503,N_14497);
nor U14575 (N_14575,N_14464,N_14512);
nor U14576 (N_14576,N_14437,N_14505);
and U14577 (N_14577,N_14465,N_14476);
xor U14578 (N_14578,N_14423,N_14490);
and U14579 (N_14579,N_14456,N_14504);
nand U14580 (N_14580,N_14519,N_14457);
xor U14581 (N_14581,N_14525,N_14471);
or U14582 (N_14582,N_14509,N_14536);
and U14583 (N_14583,N_14449,N_14411);
and U14584 (N_14584,N_14533,N_14478);
nor U14585 (N_14585,N_14444,N_14502);
nand U14586 (N_14586,N_14414,N_14558);
xnor U14587 (N_14587,N_14495,N_14516);
and U14588 (N_14588,N_14496,N_14401);
and U14589 (N_14589,N_14537,N_14441);
xor U14590 (N_14590,N_14443,N_14498);
and U14591 (N_14591,N_14554,N_14507);
or U14592 (N_14592,N_14466,N_14523);
nor U14593 (N_14593,N_14488,N_14539);
xnor U14594 (N_14594,N_14547,N_14405);
xor U14595 (N_14595,N_14552,N_14404);
or U14596 (N_14596,N_14517,N_14410);
and U14597 (N_14597,N_14485,N_14534);
and U14598 (N_14598,N_14546,N_14542);
and U14599 (N_14599,N_14416,N_14555);
or U14600 (N_14600,N_14408,N_14455);
nor U14601 (N_14601,N_14472,N_14463);
nand U14602 (N_14602,N_14428,N_14425);
nor U14603 (N_14603,N_14417,N_14480);
xnor U14604 (N_14604,N_14511,N_14514);
xor U14605 (N_14605,N_14491,N_14447);
or U14606 (N_14606,N_14556,N_14520);
and U14607 (N_14607,N_14446,N_14435);
or U14608 (N_14608,N_14424,N_14508);
xor U14609 (N_14609,N_14548,N_14470);
xor U14610 (N_14610,N_14500,N_14442);
and U14611 (N_14611,N_14430,N_14483);
and U14612 (N_14612,N_14535,N_14412);
and U14613 (N_14613,N_14557,N_14515);
or U14614 (N_14614,N_14492,N_14559);
xor U14615 (N_14615,N_14526,N_14451);
nor U14616 (N_14616,N_14513,N_14434);
or U14617 (N_14617,N_14532,N_14541);
nand U14618 (N_14618,N_14529,N_14531);
xor U14619 (N_14619,N_14524,N_14450);
xnor U14620 (N_14620,N_14543,N_14402);
nor U14621 (N_14621,N_14481,N_14484);
or U14622 (N_14622,N_14436,N_14493);
or U14623 (N_14623,N_14540,N_14407);
or U14624 (N_14624,N_14487,N_14454);
or U14625 (N_14625,N_14448,N_14510);
nand U14626 (N_14626,N_14549,N_14544);
nor U14627 (N_14627,N_14403,N_14440);
and U14628 (N_14628,N_14489,N_14460);
and U14629 (N_14629,N_14409,N_14406);
nand U14630 (N_14630,N_14474,N_14468);
nand U14631 (N_14631,N_14413,N_14553);
xnor U14632 (N_14632,N_14432,N_14459);
nand U14633 (N_14633,N_14452,N_14415);
nor U14634 (N_14634,N_14518,N_14421);
and U14635 (N_14635,N_14458,N_14418);
nand U14636 (N_14636,N_14475,N_14550);
nand U14637 (N_14637,N_14427,N_14462);
nand U14638 (N_14638,N_14545,N_14419);
nor U14639 (N_14639,N_14453,N_14528);
xor U14640 (N_14640,N_14420,N_14542);
or U14641 (N_14641,N_14460,N_14457);
xor U14642 (N_14642,N_14457,N_14475);
xor U14643 (N_14643,N_14506,N_14519);
xor U14644 (N_14644,N_14451,N_14467);
nor U14645 (N_14645,N_14468,N_14496);
nor U14646 (N_14646,N_14517,N_14491);
and U14647 (N_14647,N_14476,N_14477);
nor U14648 (N_14648,N_14412,N_14500);
or U14649 (N_14649,N_14516,N_14449);
xor U14650 (N_14650,N_14409,N_14503);
nor U14651 (N_14651,N_14495,N_14549);
nor U14652 (N_14652,N_14555,N_14553);
and U14653 (N_14653,N_14515,N_14491);
and U14654 (N_14654,N_14482,N_14498);
nor U14655 (N_14655,N_14442,N_14457);
xnor U14656 (N_14656,N_14498,N_14500);
and U14657 (N_14657,N_14472,N_14515);
and U14658 (N_14658,N_14500,N_14552);
nor U14659 (N_14659,N_14447,N_14462);
and U14660 (N_14660,N_14555,N_14547);
nand U14661 (N_14661,N_14506,N_14489);
xnor U14662 (N_14662,N_14469,N_14400);
nand U14663 (N_14663,N_14432,N_14552);
xor U14664 (N_14664,N_14413,N_14482);
xnor U14665 (N_14665,N_14507,N_14414);
and U14666 (N_14666,N_14477,N_14482);
and U14667 (N_14667,N_14447,N_14514);
or U14668 (N_14668,N_14402,N_14506);
nor U14669 (N_14669,N_14497,N_14449);
or U14670 (N_14670,N_14497,N_14532);
and U14671 (N_14671,N_14470,N_14437);
nand U14672 (N_14672,N_14403,N_14537);
xor U14673 (N_14673,N_14553,N_14478);
xnor U14674 (N_14674,N_14510,N_14556);
or U14675 (N_14675,N_14446,N_14443);
xnor U14676 (N_14676,N_14463,N_14534);
and U14677 (N_14677,N_14539,N_14557);
nor U14678 (N_14678,N_14559,N_14540);
nand U14679 (N_14679,N_14409,N_14518);
or U14680 (N_14680,N_14409,N_14559);
and U14681 (N_14681,N_14484,N_14507);
nand U14682 (N_14682,N_14438,N_14483);
nand U14683 (N_14683,N_14456,N_14542);
nor U14684 (N_14684,N_14413,N_14406);
and U14685 (N_14685,N_14435,N_14449);
nand U14686 (N_14686,N_14445,N_14437);
and U14687 (N_14687,N_14491,N_14429);
xnor U14688 (N_14688,N_14494,N_14547);
nand U14689 (N_14689,N_14412,N_14434);
and U14690 (N_14690,N_14430,N_14429);
xnor U14691 (N_14691,N_14506,N_14490);
and U14692 (N_14692,N_14406,N_14439);
and U14693 (N_14693,N_14450,N_14537);
and U14694 (N_14694,N_14522,N_14464);
or U14695 (N_14695,N_14418,N_14497);
xnor U14696 (N_14696,N_14474,N_14517);
nand U14697 (N_14697,N_14486,N_14434);
nand U14698 (N_14698,N_14484,N_14458);
or U14699 (N_14699,N_14463,N_14435);
and U14700 (N_14700,N_14516,N_14471);
nor U14701 (N_14701,N_14498,N_14466);
and U14702 (N_14702,N_14454,N_14491);
xnor U14703 (N_14703,N_14513,N_14552);
and U14704 (N_14704,N_14487,N_14409);
or U14705 (N_14705,N_14546,N_14455);
nor U14706 (N_14706,N_14539,N_14430);
nand U14707 (N_14707,N_14557,N_14403);
or U14708 (N_14708,N_14499,N_14541);
nor U14709 (N_14709,N_14489,N_14548);
or U14710 (N_14710,N_14495,N_14494);
nand U14711 (N_14711,N_14434,N_14441);
or U14712 (N_14712,N_14545,N_14476);
nor U14713 (N_14713,N_14406,N_14520);
xnor U14714 (N_14714,N_14440,N_14510);
or U14715 (N_14715,N_14499,N_14455);
nand U14716 (N_14716,N_14488,N_14506);
or U14717 (N_14717,N_14557,N_14475);
and U14718 (N_14718,N_14416,N_14550);
xor U14719 (N_14719,N_14517,N_14554);
and U14720 (N_14720,N_14603,N_14662);
nand U14721 (N_14721,N_14669,N_14580);
or U14722 (N_14722,N_14701,N_14710);
nand U14723 (N_14723,N_14686,N_14652);
nor U14724 (N_14724,N_14604,N_14594);
or U14725 (N_14725,N_14632,N_14614);
or U14726 (N_14726,N_14587,N_14621);
and U14727 (N_14727,N_14688,N_14615);
and U14728 (N_14728,N_14576,N_14613);
and U14729 (N_14729,N_14649,N_14646);
and U14730 (N_14730,N_14638,N_14661);
xnor U14731 (N_14731,N_14696,N_14656);
xnor U14732 (N_14732,N_14679,N_14663);
and U14733 (N_14733,N_14709,N_14672);
or U14734 (N_14734,N_14566,N_14597);
nor U14735 (N_14735,N_14637,N_14634);
and U14736 (N_14736,N_14627,N_14591);
xnor U14737 (N_14737,N_14700,N_14602);
xor U14738 (N_14738,N_14673,N_14691);
nor U14739 (N_14739,N_14648,N_14645);
xor U14740 (N_14740,N_14577,N_14714);
xnor U14741 (N_14741,N_14703,N_14573);
xnor U14742 (N_14742,N_14625,N_14647);
xor U14743 (N_14743,N_14631,N_14562);
nor U14744 (N_14744,N_14600,N_14711);
nor U14745 (N_14745,N_14674,N_14639);
nor U14746 (N_14746,N_14707,N_14706);
xor U14747 (N_14747,N_14644,N_14590);
or U14748 (N_14748,N_14579,N_14687);
nand U14749 (N_14749,N_14693,N_14596);
xnor U14750 (N_14750,N_14702,N_14628);
nor U14751 (N_14751,N_14593,N_14713);
or U14752 (N_14752,N_14574,N_14609);
nor U14753 (N_14753,N_14650,N_14623);
and U14754 (N_14754,N_14581,N_14651);
and U14755 (N_14755,N_14681,N_14712);
nand U14756 (N_14756,N_14560,N_14680);
xor U14757 (N_14757,N_14716,N_14629);
xor U14758 (N_14758,N_14698,N_14624);
xnor U14759 (N_14759,N_14689,N_14578);
or U14760 (N_14760,N_14564,N_14563);
nand U14761 (N_14761,N_14616,N_14584);
and U14762 (N_14762,N_14565,N_14641);
and U14763 (N_14763,N_14690,N_14658);
and U14764 (N_14764,N_14588,N_14575);
or U14765 (N_14765,N_14717,N_14595);
or U14766 (N_14766,N_14607,N_14571);
and U14767 (N_14767,N_14660,N_14675);
or U14768 (N_14768,N_14583,N_14642);
nand U14769 (N_14769,N_14635,N_14569);
xor U14770 (N_14770,N_14608,N_14589);
xnor U14771 (N_14771,N_14657,N_14683);
and U14772 (N_14772,N_14668,N_14630);
nand U14773 (N_14773,N_14708,N_14682);
and U14774 (N_14774,N_14685,N_14611);
xnor U14775 (N_14775,N_14666,N_14677);
nor U14776 (N_14776,N_14606,N_14715);
nor U14777 (N_14777,N_14664,N_14655);
xor U14778 (N_14778,N_14699,N_14695);
nor U14779 (N_14779,N_14653,N_14705);
or U14780 (N_14780,N_14620,N_14619);
and U14781 (N_14781,N_14697,N_14636);
nor U14782 (N_14782,N_14570,N_14601);
xor U14783 (N_14783,N_14605,N_14622);
nand U14784 (N_14784,N_14610,N_14665);
or U14785 (N_14785,N_14678,N_14667);
nor U14786 (N_14786,N_14567,N_14612);
xnor U14787 (N_14787,N_14568,N_14704);
nand U14788 (N_14788,N_14692,N_14670);
and U14789 (N_14789,N_14598,N_14684);
or U14790 (N_14790,N_14592,N_14640);
and U14791 (N_14791,N_14694,N_14586);
nand U14792 (N_14792,N_14719,N_14618);
or U14793 (N_14793,N_14633,N_14572);
xor U14794 (N_14794,N_14585,N_14561);
and U14795 (N_14795,N_14617,N_14718);
or U14796 (N_14796,N_14626,N_14659);
and U14797 (N_14797,N_14676,N_14671);
and U14798 (N_14798,N_14643,N_14582);
xnor U14799 (N_14799,N_14654,N_14599);
xor U14800 (N_14800,N_14658,N_14570);
nand U14801 (N_14801,N_14648,N_14571);
nor U14802 (N_14802,N_14575,N_14656);
and U14803 (N_14803,N_14681,N_14641);
nand U14804 (N_14804,N_14695,N_14630);
and U14805 (N_14805,N_14568,N_14574);
nor U14806 (N_14806,N_14574,N_14561);
nor U14807 (N_14807,N_14560,N_14658);
nor U14808 (N_14808,N_14636,N_14604);
and U14809 (N_14809,N_14688,N_14599);
xnor U14810 (N_14810,N_14635,N_14612);
nand U14811 (N_14811,N_14561,N_14717);
nand U14812 (N_14812,N_14694,N_14563);
or U14813 (N_14813,N_14597,N_14677);
and U14814 (N_14814,N_14631,N_14603);
or U14815 (N_14815,N_14718,N_14599);
nand U14816 (N_14816,N_14708,N_14614);
and U14817 (N_14817,N_14705,N_14660);
xor U14818 (N_14818,N_14701,N_14591);
and U14819 (N_14819,N_14571,N_14718);
nor U14820 (N_14820,N_14633,N_14626);
nand U14821 (N_14821,N_14646,N_14581);
nor U14822 (N_14822,N_14707,N_14689);
xor U14823 (N_14823,N_14667,N_14714);
nor U14824 (N_14824,N_14713,N_14643);
or U14825 (N_14825,N_14632,N_14600);
xnor U14826 (N_14826,N_14674,N_14677);
nor U14827 (N_14827,N_14574,N_14707);
nor U14828 (N_14828,N_14669,N_14629);
or U14829 (N_14829,N_14682,N_14701);
xor U14830 (N_14830,N_14704,N_14705);
or U14831 (N_14831,N_14657,N_14709);
nand U14832 (N_14832,N_14574,N_14690);
or U14833 (N_14833,N_14573,N_14709);
or U14834 (N_14834,N_14697,N_14604);
nor U14835 (N_14835,N_14642,N_14654);
and U14836 (N_14836,N_14700,N_14711);
or U14837 (N_14837,N_14562,N_14580);
nand U14838 (N_14838,N_14595,N_14687);
and U14839 (N_14839,N_14596,N_14673);
nor U14840 (N_14840,N_14617,N_14652);
nor U14841 (N_14841,N_14716,N_14701);
nor U14842 (N_14842,N_14578,N_14678);
or U14843 (N_14843,N_14586,N_14560);
and U14844 (N_14844,N_14576,N_14675);
and U14845 (N_14845,N_14677,N_14692);
nor U14846 (N_14846,N_14696,N_14596);
and U14847 (N_14847,N_14600,N_14635);
or U14848 (N_14848,N_14713,N_14708);
or U14849 (N_14849,N_14698,N_14664);
and U14850 (N_14850,N_14594,N_14702);
or U14851 (N_14851,N_14719,N_14658);
and U14852 (N_14852,N_14704,N_14667);
xnor U14853 (N_14853,N_14690,N_14646);
xor U14854 (N_14854,N_14561,N_14579);
or U14855 (N_14855,N_14580,N_14589);
xor U14856 (N_14856,N_14645,N_14689);
nor U14857 (N_14857,N_14623,N_14691);
and U14858 (N_14858,N_14600,N_14630);
nand U14859 (N_14859,N_14583,N_14631);
and U14860 (N_14860,N_14693,N_14627);
or U14861 (N_14861,N_14694,N_14579);
nand U14862 (N_14862,N_14699,N_14581);
nand U14863 (N_14863,N_14719,N_14609);
or U14864 (N_14864,N_14672,N_14578);
nor U14865 (N_14865,N_14643,N_14667);
nor U14866 (N_14866,N_14611,N_14580);
xnor U14867 (N_14867,N_14614,N_14568);
and U14868 (N_14868,N_14717,N_14712);
nand U14869 (N_14869,N_14585,N_14579);
and U14870 (N_14870,N_14649,N_14562);
and U14871 (N_14871,N_14631,N_14699);
nor U14872 (N_14872,N_14562,N_14694);
nand U14873 (N_14873,N_14700,N_14673);
and U14874 (N_14874,N_14668,N_14697);
nand U14875 (N_14875,N_14698,N_14634);
xor U14876 (N_14876,N_14660,N_14599);
xor U14877 (N_14877,N_14634,N_14636);
and U14878 (N_14878,N_14692,N_14618);
nand U14879 (N_14879,N_14678,N_14682);
xor U14880 (N_14880,N_14829,N_14855);
or U14881 (N_14881,N_14872,N_14796);
nand U14882 (N_14882,N_14877,N_14878);
nor U14883 (N_14883,N_14833,N_14739);
and U14884 (N_14884,N_14873,N_14874);
or U14885 (N_14885,N_14861,N_14795);
or U14886 (N_14886,N_14757,N_14814);
and U14887 (N_14887,N_14842,N_14737);
nor U14888 (N_14888,N_14857,N_14759);
and U14889 (N_14889,N_14723,N_14782);
nand U14890 (N_14890,N_14865,N_14845);
nand U14891 (N_14891,N_14791,N_14822);
and U14892 (N_14892,N_14863,N_14787);
and U14893 (N_14893,N_14843,N_14836);
or U14894 (N_14894,N_14762,N_14773);
xor U14895 (N_14895,N_14847,N_14775);
or U14896 (N_14896,N_14850,N_14806);
or U14897 (N_14897,N_14870,N_14741);
or U14898 (N_14898,N_14736,N_14776);
or U14899 (N_14899,N_14751,N_14835);
nor U14900 (N_14900,N_14720,N_14876);
xnor U14901 (N_14901,N_14753,N_14778);
nand U14902 (N_14902,N_14788,N_14760);
nor U14903 (N_14903,N_14837,N_14821);
nor U14904 (N_14904,N_14802,N_14729);
and U14905 (N_14905,N_14823,N_14860);
or U14906 (N_14906,N_14830,N_14746);
nor U14907 (N_14907,N_14811,N_14804);
xor U14908 (N_14908,N_14727,N_14844);
and U14909 (N_14909,N_14783,N_14755);
nand U14910 (N_14910,N_14854,N_14747);
and U14911 (N_14911,N_14828,N_14766);
nand U14912 (N_14912,N_14820,N_14864);
nor U14913 (N_14913,N_14813,N_14725);
or U14914 (N_14914,N_14771,N_14832);
nor U14915 (N_14915,N_14786,N_14834);
or U14916 (N_14916,N_14765,N_14868);
nor U14917 (N_14917,N_14824,N_14790);
nor U14918 (N_14918,N_14721,N_14826);
nand U14919 (N_14919,N_14767,N_14779);
or U14920 (N_14920,N_14867,N_14797);
nor U14921 (N_14921,N_14774,N_14841);
or U14922 (N_14922,N_14740,N_14754);
or U14923 (N_14923,N_14726,N_14858);
or U14924 (N_14924,N_14808,N_14758);
or U14925 (N_14925,N_14848,N_14819);
nor U14926 (N_14926,N_14849,N_14815);
nor U14927 (N_14927,N_14732,N_14856);
and U14928 (N_14928,N_14810,N_14827);
nor U14929 (N_14929,N_14839,N_14871);
or U14930 (N_14930,N_14785,N_14825);
nand U14931 (N_14931,N_14772,N_14724);
xnor U14932 (N_14932,N_14731,N_14735);
nor U14933 (N_14933,N_14807,N_14764);
xor U14934 (N_14934,N_14734,N_14862);
and U14935 (N_14935,N_14879,N_14798);
and U14936 (N_14936,N_14803,N_14780);
and U14937 (N_14937,N_14792,N_14852);
xnor U14938 (N_14938,N_14777,N_14859);
or U14939 (N_14939,N_14745,N_14728);
and U14940 (N_14940,N_14730,N_14816);
and U14941 (N_14941,N_14809,N_14750);
nor U14942 (N_14942,N_14763,N_14784);
and U14943 (N_14943,N_14851,N_14733);
xor U14944 (N_14944,N_14866,N_14875);
nor U14945 (N_14945,N_14800,N_14749);
nand U14946 (N_14946,N_14853,N_14789);
nand U14947 (N_14947,N_14793,N_14769);
nor U14948 (N_14948,N_14743,N_14799);
xor U14949 (N_14949,N_14801,N_14812);
nor U14950 (N_14950,N_14840,N_14761);
nor U14951 (N_14951,N_14748,N_14722);
and U14952 (N_14952,N_14794,N_14817);
and U14953 (N_14953,N_14756,N_14738);
nand U14954 (N_14954,N_14846,N_14752);
nand U14955 (N_14955,N_14869,N_14838);
nand U14956 (N_14956,N_14818,N_14805);
nand U14957 (N_14957,N_14744,N_14768);
nor U14958 (N_14958,N_14781,N_14742);
nand U14959 (N_14959,N_14770,N_14831);
or U14960 (N_14960,N_14842,N_14784);
nand U14961 (N_14961,N_14810,N_14828);
or U14962 (N_14962,N_14814,N_14875);
xor U14963 (N_14963,N_14731,N_14752);
or U14964 (N_14964,N_14876,N_14765);
and U14965 (N_14965,N_14833,N_14859);
nand U14966 (N_14966,N_14878,N_14794);
or U14967 (N_14967,N_14836,N_14753);
or U14968 (N_14968,N_14826,N_14765);
or U14969 (N_14969,N_14814,N_14762);
nand U14970 (N_14970,N_14863,N_14874);
nor U14971 (N_14971,N_14755,N_14746);
xor U14972 (N_14972,N_14854,N_14822);
or U14973 (N_14973,N_14815,N_14768);
and U14974 (N_14974,N_14807,N_14842);
nand U14975 (N_14975,N_14802,N_14747);
and U14976 (N_14976,N_14751,N_14845);
or U14977 (N_14977,N_14845,N_14791);
or U14978 (N_14978,N_14811,N_14722);
and U14979 (N_14979,N_14757,N_14846);
nor U14980 (N_14980,N_14798,N_14795);
xnor U14981 (N_14981,N_14779,N_14784);
and U14982 (N_14982,N_14853,N_14793);
and U14983 (N_14983,N_14848,N_14847);
nand U14984 (N_14984,N_14763,N_14870);
nand U14985 (N_14985,N_14730,N_14825);
nand U14986 (N_14986,N_14753,N_14765);
or U14987 (N_14987,N_14854,N_14865);
or U14988 (N_14988,N_14762,N_14829);
and U14989 (N_14989,N_14770,N_14783);
nand U14990 (N_14990,N_14827,N_14727);
xor U14991 (N_14991,N_14818,N_14728);
nor U14992 (N_14992,N_14734,N_14834);
xnor U14993 (N_14993,N_14731,N_14757);
nand U14994 (N_14994,N_14822,N_14724);
and U14995 (N_14995,N_14781,N_14787);
nor U14996 (N_14996,N_14826,N_14801);
nand U14997 (N_14997,N_14741,N_14774);
nor U14998 (N_14998,N_14813,N_14869);
and U14999 (N_14999,N_14801,N_14845);
nand U15000 (N_15000,N_14734,N_14801);
and U15001 (N_15001,N_14730,N_14836);
xnor U15002 (N_15002,N_14743,N_14727);
xnor U15003 (N_15003,N_14747,N_14845);
and U15004 (N_15004,N_14777,N_14844);
xnor U15005 (N_15005,N_14763,N_14750);
and U15006 (N_15006,N_14845,N_14834);
nand U15007 (N_15007,N_14752,N_14765);
and U15008 (N_15008,N_14740,N_14772);
or U15009 (N_15009,N_14826,N_14850);
xnor U15010 (N_15010,N_14821,N_14878);
nor U15011 (N_15011,N_14765,N_14819);
nor U15012 (N_15012,N_14829,N_14741);
nor U15013 (N_15013,N_14731,N_14771);
xor U15014 (N_15014,N_14722,N_14791);
xor U15015 (N_15015,N_14838,N_14731);
and U15016 (N_15016,N_14746,N_14751);
nand U15017 (N_15017,N_14834,N_14791);
or U15018 (N_15018,N_14724,N_14860);
xor U15019 (N_15019,N_14768,N_14754);
nand U15020 (N_15020,N_14864,N_14730);
and U15021 (N_15021,N_14767,N_14875);
xor U15022 (N_15022,N_14747,N_14831);
xor U15023 (N_15023,N_14807,N_14810);
and U15024 (N_15024,N_14765,N_14823);
nand U15025 (N_15025,N_14825,N_14743);
or U15026 (N_15026,N_14743,N_14765);
and U15027 (N_15027,N_14806,N_14827);
xor U15028 (N_15028,N_14873,N_14879);
nand U15029 (N_15029,N_14866,N_14854);
nor U15030 (N_15030,N_14826,N_14744);
or U15031 (N_15031,N_14744,N_14778);
and U15032 (N_15032,N_14849,N_14833);
and U15033 (N_15033,N_14791,N_14838);
xnor U15034 (N_15034,N_14821,N_14733);
xor U15035 (N_15035,N_14856,N_14799);
nand U15036 (N_15036,N_14825,N_14800);
nand U15037 (N_15037,N_14826,N_14864);
nand U15038 (N_15038,N_14729,N_14789);
and U15039 (N_15039,N_14873,N_14749);
xor U15040 (N_15040,N_14897,N_14953);
and U15041 (N_15041,N_14932,N_14934);
nor U15042 (N_15042,N_14935,N_14965);
nor U15043 (N_15043,N_14975,N_14928);
nand U15044 (N_15044,N_14908,N_14954);
xnor U15045 (N_15045,N_14956,N_14994);
or U15046 (N_15046,N_15014,N_15019);
nand U15047 (N_15047,N_14930,N_14959);
nand U15048 (N_15048,N_15020,N_14986);
or U15049 (N_15049,N_15007,N_14906);
and U15050 (N_15050,N_14915,N_14991);
and U15051 (N_15051,N_14937,N_14923);
nor U15052 (N_15052,N_14983,N_14992);
nand U15053 (N_15053,N_14913,N_14939);
or U15054 (N_15054,N_14885,N_15009);
and U15055 (N_15055,N_14996,N_14922);
or U15056 (N_15056,N_14957,N_14989);
nand U15057 (N_15057,N_14900,N_14898);
and U15058 (N_15058,N_14899,N_15035);
nand U15059 (N_15059,N_14974,N_14893);
and U15060 (N_15060,N_15024,N_14999);
nand U15061 (N_15061,N_14907,N_14942);
or U15062 (N_15062,N_14955,N_14951);
or U15063 (N_15063,N_14921,N_14990);
and U15064 (N_15064,N_15017,N_14909);
nand U15065 (N_15065,N_14917,N_14949);
nor U15066 (N_15066,N_14998,N_15039);
or U15067 (N_15067,N_15004,N_15008);
nand U15068 (N_15068,N_14927,N_14941);
and U15069 (N_15069,N_14887,N_14895);
nor U15070 (N_15070,N_14976,N_14919);
and U15071 (N_15071,N_14972,N_15006);
or U15072 (N_15072,N_14968,N_14982);
nand U15073 (N_15073,N_15028,N_14993);
xnor U15074 (N_15074,N_14914,N_14980);
or U15075 (N_15075,N_14946,N_15001);
and U15076 (N_15076,N_15010,N_15038);
nand U15077 (N_15077,N_14890,N_14910);
nand U15078 (N_15078,N_14926,N_14967);
nand U15079 (N_15079,N_14902,N_14943);
nand U15080 (N_15080,N_14905,N_14966);
and U15081 (N_15081,N_15037,N_14938);
or U15082 (N_15082,N_14901,N_14916);
or U15083 (N_15083,N_15013,N_15025);
and U15084 (N_15084,N_14880,N_14945);
xor U15085 (N_15085,N_14904,N_15002);
xor U15086 (N_15086,N_14948,N_14911);
or U15087 (N_15087,N_15012,N_14984);
and U15088 (N_15088,N_15027,N_14925);
or U15089 (N_15089,N_14912,N_15011);
nor U15090 (N_15090,N_14981,N_14891);
xor U15091 (N_15091,N_15036,N_15034);
or U15092 (N_15092,N_14920,N_15015);
nor U15093 (N_15093,N_14977,N_14987);
nand U15094 (N_15094,N_14963,N_15018);
and U15095 (N_15095,N_14940,N_14952);
xor U15096 (N_15096,N_14979,N_15005);
and U15097 (N_15097,N_14881,N_14936);
or U15098 (N_15098,N_14950,N_15031);
or U15099 (N_15099,N_14918,N_14969);
and U15100 (N_15100,N_14944,N_14933);
nand U15101 (N_15101,N_14964,N_14892);
nor U15102 (N_15102,N_15021,N_14888);
and U15103 (N_15103,N_15016,N_14886);
nor U15104 (N_15104,N_15029,N_15022);
nor U15105 (N_15105,N_15000,N_14988);
xnor U15106 (N_15106,N_14970,N_14997);
nand U15107 (N_15107,N_14894,N_15030);
nor U15108 (N_15108,N_14971,N_14947);
xor U15109 (N_15109,N_15032,N_14973);
or U15110 (N_15110,N_15033,N_15023);
or U15111 (N_15111,N_15026,N_14884);
nand U15112 (N_15112,N_14960,N_14961);
xnor U15113 (N_15113,N_14924,N_15003);
nand U15114 (N_15114,N_14889,N_14958);
nor U15115 (N_15115,N_14985,N_14929);
xor U15116 (N_15116,N_14962,N_14978);
xnor U15117 (N_15117,N_14882,N_14931);
or U15118 (N_15118,N_14883,N_14995);
nand U15119 (N_15119,N_14896,N_14903);
xor U15120 (N_15120,N_14920,N_14938);
xnor U15121 (N_15121,N_14966,N_14911);
nand U15122 (N_15122,N_14896,N_14952);
or U15123 (N_15123,N_14898,N_14902);
nor U15124 (N_15124,N_14924,N_14961);
nand U15125 (N_15125,N_14908,N_14917);
and U15126 (N_15126,N_15003,N_15027);
xnor U15127 (N_15127,N_15003,N_14971);
or U15128 (N_15128,N_14937,N_14911);
and U15129 (N_15129,N_14995,N_14951);
xnor U15130 (N_15130,N_14920,N_14915);
or U15131 (N_15131,N_14895,N_14926);
xor U15132 (N_15132,N_14942,N_14955);
nand U15133 (N_15133,N_15000,N_15032);
or U15134 (N_15134,N_15016,N_14978);
nor U15135 (N_15135,N_15014,N_14899);
nor U15136 (N_15136,N_15002,N_14930);
or U15137 (N_15137,N_14927,N_14900);
nand U15138 (N_15138,N_14971,N_14930);
and U15139 (N_15139,N_15036,N_15011);
xnor U15140 (N_15140,N_14886,N_15023);
and U15141 (N_15141,N_14957,N_14909);
or U15142 (N_15142,N_14952,N_15036);
xnor U15143 (N_15143,N_14909,N_14947);
xor U15144 (N_15144,N_14900,N_14915);
nor U15145 (N_15145,N_15008,N_15006);
nor U15146 (N_15146,N_14983,N_14957);
xnor U15147 (N_15147,N_14939,N_14900);
or U15148 (N_15148,N_14953,N_14913);
nor U15149 (N_15149,N_14917,N_15029);
nor U15150 (N_15150,N_14903,N_14980);
or U15151 (N_15151,N_14919,N_14916);
nor U15152 (N_15152,N_14937,N_14989);
nand U15153 (N_15153,N_14924,N_14910);
nor U15154 (N_15154,N_14913,N_14925);
nand U15155 (N_15155,N_14921,N_14994);
nand U15156 (N_15156,N_14941,N_14961);
xor U15157 (N_15157,N_15023,N_14954);
xor U15158 (N_15158,N_14975,N_15022);
nor U15159 (N_15159,N_15034,N_14986);
nor U15160 (N_15160,N_14983,N_15034);
and U15161 (N_15161,N_14907,N_14957);
or U15162 (N_15162,N_14907,N_14881);
or U15163 (N_15163,N_14999,N_14948);
xor U15164 (N_15164,N_15024,N_14987);
xnor U15165 (N_15165,N_14934,N_15018);
xor U15166 (N_15166,N_15036,N_15014);
xor U15167 (N_15167,N_14957,N_15015);
xnor U15168 (N_15168,N_15032,N_14945);
and U15169 (N_15169,N_15014,N_14976);
or U15170 (N_15170,N_15034,N_14990);
xnor U15171 (N_15171,N_14902,N_15005);
and U15172 (N_15172,N_14975,N_14885);
or U15173 (N_15173,N_14963,N_14994);
nand U15174 (N_15174,N_14897,N_14969);
nor U15175 (N_15175,N_14941,N_14995);
xor U15176 (N_15176,N_14961,N_15021);
xnor U15177 (N_15177,N_14887,N_14993);
nor U15178 (N_15178,N_14963,N_14883);
nand U15179 (N_15179,N_15011,N_14924);
nor U15180 (N_15180,N_15022,N_14964);
xnor U15181 (N_15181,N_15036,N_14956);
or U15182 (N_15182,N_15034,N_15032);
and U15183 (N_15183,N_14885,N_14928);
nor U15184 (N_15184,N_15027,N_14928);
and U15185 (N_15185,N_14999,N_14912);
nor U15186 (N_15186,N_14974,N_14922);
or U15187 (N_15187,N_14910,N_14903);
nor U15188 (N_15188,N_15012,N_15035);
and U15189 (N_15189,N_14991,N_14893);
xor U15190 (N_15190,N_15002,N_14967);
and U15191 (N_15191,N_14980,N_14950);
and U15192 (N_15192,N_14931,N_14881);
nand U15193 (N_15193,N_14920,N_14956);
nand U15194 (N_15194,N_14946,N_14963);
or U15195 (N_15195,N_15018,N_14948);
or U15196 (N_15196,N_14887,N_15025);
or U15197 (N_15197,N_14989,N_14962);
nand U15198 (N_15198,N_14915,N_14904);
or U15199 (N_15199,N_14989,N_14946);
xor U15200 (N_15200,N_15173,N_15128);
nor U15201 (N_15201,N_15146,N_15192);
and U15202 (N_15202,N_15119,N_15102);
nand U15203 (N_15203,N_15111,N_15155);
xnor U15204 (N_15204,N_15114,N_15181);
nor U15205 (N_15205,N_15162,N_15093);
xor U15206 (N_15206,N_15041,N_15169);
nor U15207 (N_15207,N_15077,N_15105);
nand U15208 (N_15208,N_15071,N_15110);
or U15209 (N_15209,N_15183,N_15067);
nor U15210 (N_15210,N_15157,N_15051);
nand U15211 (N_15211,N_15138,N_15060);
nor U15212 (N_15212,N_15124,N_15196);
nand U15213 (N_15213,N_15094,N_15085);
nor U15214 (N_15214,N_15160,N_15062);
and U15215 (N_15215,N_15167,N_15099);
or U15216 (N_15216,N_15141,N_15191);
nor U15217 (N_15217,N_15042,N_15069);
or U15218 (N_15218,N_15190,N_15199);
and U15219 (N_15219,N_15156,N_15040);
nor U15220 (N_15220,N_15166,N_15090);
nand U15221 (N_15221,N_15152,N_15074);
nor U15222 (N_15222,N_15121,N_15115);
and U15223 (N_15223,N_15170,N_15125);
xor U15224 (N_15224,N_15047,N_15043);
nand U15225 (N_15225,N_15061,N_15165);
nor U15226 (N_15226,N_15188,N_15063);
or U15227 (N_15227,N_15055,N_15100);
nor U15228 (N_15228,N_15149,N_15147);
nand U15229 (N_15229,N_15133,N_15186);
and U15230 (N_15230,N_15076,N_15129);
nand U15231 (N_15231,N_15123,N_15044);
xor U15232 (N_15232,N_15104,N_15171);
nand U15233 (N_15233,N_15189,N_15184);
nor U15234 (N_15234,N_15070,N_15134);
and U15235 (N_15235,N_15112,N_15096);
and U15236 (N_15236,N_15127,N_15180);
nor U15237 (N_15237,N_15049,N_15116);
nand U15238 (N_15238,N_15117,N_15084);
and U15239 (N_15239,N_15059,N_15136);
xor U15240 (N_15240,N_15075,N_15187);
nand U15241 (N_15241,N_15176,N_15088);
xnor U15242 (N_15242,N_15080,N_15172);
xor U15243 (N_15243,N_15078,N_15135);
and U15244 (N_15244,N_15109,N_15106);
xor U15245 (N_15245,N_15193,N_15178);
nand U15246 (N_15246,N_15058,N_15198);
and U15247 (N_15247,N_15056,N_15145);
nor U15248 (N_15248,N_15103,N_15097);
nand U15249 (N_15249,N_15045,N_15050);
nand U15250 (N_15250,N_15081,N_15143);
and U15251 (N_15251,N_15066,N_15154);
nor U15252 (N_15252,N_15158,N_15054);
nand U15253 (N_15253,N_15083,N_15086);
xnor U15254 (N_15254,N_15072,N_15150);
xnor U15255 (N_15255,N_15132,N_15140);
nor U15256 (N_15256,N_15091,N_15068);
xor U15257 (N_15257,N_15098,N_15101);
and U15258 (N_15258,N_15175,N_15148);
nand U15259 (N_15259,N_15130,N_15151);
or U15260 (N_15260,N_15064,N_15163);
nand U15261 (N_15261,N_15079,N_15065);
xnor U15262 (N_15262,N_15118,N_15168);
xor U15263 (N_15263,N_15179,N_15185);
nor U15264 (N_15264,N_15120,N_15092);
and U15265 (N_15265,N_15144,N_15137);
xor U15266 (N_15266,N_15122,N_15089);
nand U15267 (N_15267,N_15177,N_15194);
and U15268 (N_15268,N_15108,N_15073);
xnor U15269 (N_15269,N_15052,N_15139);
nand U15270 (N_15270,N_15182,N_15164);
and U15271 (N_15271,N_15057,N_15113);
and U15272 (N_15272,N_15159,N_15095);
nor U15273 (N_15273,N_15174,N_15107);
or U15274 (N_15274,N_15153,N_15142);
and U15275 (N_15275,N_15082,N_15195);
nor U15276 (N_15276,N_15131,N_15046);
nor U15277 (N_15277,N_15197,N_15048);
nand U15278 (N_15278,N_15053,N_15126);
nand U15279 (N_15279,N_15087,N_15161);
xnor U15280 (N_15280,N_15098,N_15068);
or U15281 (N_15281,N_15164,N_15076);
or U15282 (N_15282,N_15165,N_15096);
nand U15283 (N_15283,N_15050,N_15170);
or U15284 (N_15284,N_15186,N_15196);
nand U15285 (N_15285,N_15130,N_15046);
and U15286 (N_15286,N_15085,N_15163);
and U15287 (N_15287,N_15154,N_15137);
nor U15288 (N_15288,N_15159,N_15087);
or U15289 (N_15289,N_15148,N_15165);
and U15290 (N_15290,N_15080,N_15078);
and U15291 (N_15291,N_15071,N_15153);
nand U15292 (N_15292,N_15159,N_15045);
xor U15293 (N_15293,N_15056,N_15187);
nand U15294 (N_15294,N_15067,N_15187);
nand U15295 (N_15295,N_15079,N_15149);
or U15296 (N_15296,N_15059,N_15071);
and U15297 (N_15297,N_15097,N_15148);
nand U15298 (N_15298,N_15184,N_15125);
or U15299 (N_15299,N_15064,N_15199);
nor U15300 (N_15300,N_15070,N_15095);
and U15301 (N_15301,N_15169,N_15128);
or U15302 (N_15302,N_15116,N_15181);
xnor U15303 (N_15303,N_15128,N_15040);
or U15304 (N_15304,N_15145,N_15110);
nand U15305 (N_15305,N_15041,N_15121);
or U15306 (N_15306,N_15052,N_15195);
xor U15307 (N_15307,N_15198,N_15162);
xor U15308 (N_15308,N_15143,N_15160);
xor U15309 (N_15309,N_15086,N_15123);
and U15310 (N_15310,N_15123,N_15060);
nor U15311 (N_15311,N_15043,N_15143);
xor U15312 (N_15312,N_15194,N_15084);
nor U15313 (N_15313,N_15100,N_15052);
xnor U15314 (N_15314,N_15112,N_15126);
xnor U15315 (N_15315,N_15182,N_15112);
or U15316 (N_15316,N_15191,N_15086);
or U15317 (N_15317,N_15115,N_15094);
nor U15318 (N_15318,N_15136,N_15082);
nand U15319 (N_15319,N_15069,N_15047);
nor U15320 (N_15320,N_15091,N_15164);
or U15321 (N_15321,N_15162,N_15091);
nand U15322 (N_15322,N_15133,N_15153);
and U15323 (N_15323,N_15082,N_15192);
nand U15324 (N_15324,N_15154,N_15092);
nor U15325 (N_15325,N_15185,N_15109);
or U15326 (N_15326,N_15164,N_15197);
and U15327 (N_15327,N_15139,N_15103);
and U15328 (N_15328,N_15081,N_15095);
nand U15329 (N_15329,N_15131,N_15109);
nor U15330 (N_15330,N_15063,N_15198);
nor U15331 (N_15331,N_15136,N_15040);
or U15332 (N_15332,N_15184,N_15132);
xnor U15333 (N_15333,N_15108,N_15186);
xor U15334 (N_15334,N_15088,N_15189);
and U15335 (N_15335,N_15189,N_15164);
xnor U15336 (N_15336,N_15148,N_15077);
nand U15337 (N_15337,N_15141,N_15041);
nor U15338 (N_15338,N_15156,N_15118);
xor U15339 (N_15339,N_15098,N_15102);
nor U15340 (N_15340,N_15189,N_15177);
and U15341 (N_15341,N_15090,N_15115);
and U15342 (N_15342,N_15063,N_15058);
nand U15343 (N_15343,N_15076,N_15111);
xnor U15344 (N_15344,N_15182,N_15171);
nor U15345 (N_15345,N_15051,N_15081);
or U15346 (N_15346,N_15148,N_15160);
nor U15347 (N_15347,N_15156,N_15100);
nor U15348 (N_15348,N_15142,N_15126);
and U15349 (N_15349,N_15178,N_15191);
nor U15350 (N_15350,N_15075,N_15190);
or U15351 (N_15351,N_15177,N_15088);
nor U15352 (N_15352,N_15060,N_15161);
and U15353 (N_15353,N_15158,N_15090);
or U15354 (N_15354,N_15079,N_15084);
nand U15355 (N_15355,N_15077,N_15102);
nor U15356 (N_15356,N_15193,N_15192);
xnor U15357 (N_15357,N_15199,N_15173);
nand U15358 (N_15358,N_15054,N_15100);
or U15359 (N_15359,N_15113,N_15110);
nand U15360 (N_15360,N_15291,N_15315);
nand U15361 (N_15361,N_15323,N_15327);
xor U15362 (N_15362,N_15268,N_15350);
nor U15363 (N_15363,N_15285,N_15279);
xor U15364 (N_15364,N_15329,N_15302);
nand U15365 (N_15365,N_15270,N_15335);
xnor U15366 (N_15366,N_15269,N_15313);
nand U15367 (N_15367,N_15214,N_15330);
nor U15368 (N_15368,N_15341,N_15278);
xor U15369 (N_15369,N_15203,N_15276);
nand U15370 (N_15370,N_15227,N_15211);
and U15371 (N_15371,N_15239,N_15282);
xor U15372 (N_15372,N_15243,N_15308);
xnor U15373 (N_15373,N_15314,N_15273);
nor U15374 (N_15374,N_15244,N_15353);
nor U15375 (N_15375,N_15298,N_15263);
nor U15376 (N_15376,N_15326,N_15252);
and U15377 (N_15377,N_15344,N_15320);
or U15378 (N_15378,N_15334,N_15296);
xor U15379 (N_15379,N_15222,N_15259);
and U15380 (N_15380,N_15242,N_15357);
or U15381 (N_15381,N_15289,N_15297);
and U15382 (N_15382,N_15339,N_15256);
nor U15383 (N_15383,N_15359,N_15245);
and U15384 (N_15384,N_15200,N_15286);
nor U15385 (N_15385,N_15241,N_15325);
or U15386 (N_15386,N_15295,N_15292);
or U15387 (N_15387,N_15262,N_15342);
xnor U15388 (N_15388,N_15304,N_15224);
nor U15389 (N_15389,N_15305,N_15293);
nor U15390 (N_15390,N_15358,N_15299);
or U15391 (N_15391,N_15218,N_15319);
nand U15392 (N_15392,N_15281,N_15260);
or U15393 (N_15393,N_15340,N_15231);
nand U15394 (N_15394,N_15254,N_15247);
nor U15395 (N_15395,N_15322,N_15250);
nand U15396 (N_15396,N_15205,N_15215);
nand U15397 (N_15397,N_15294,N_15354);
and U15398 (N_15398,N_15201,N_15347);
or U15399 (N_15399,N_15253,N_15246);
xor U15400 (N_15400,N_15232,N_15223);
xnor U15401 (N_15401,N_15272,N_15346);
nor U15402 (N_15402,N_15275,N_15213);
nand U15403 (N_15403,N_15237,N_15216);
xnor U15404 (N_15404,N_15331,N_15311);
and U15405 (N_15405,N_15235,N_15306);
nand U15406 (N_15406,N_15351,N_15321);
and U15407 (N_15407,N_15349,N_15348);
xnor U15408 (N_15408,N_15290,N_15318);
nand U15409 (N_15409,N_15217,N_15345);
nor U15410 (N_15410,N_15343,N_15312);
or U15411 (N_15411,N_15287,N_15352);
nor U15412 (N_15412,N_15219,N_15257);
xor U15413 (N_15413,N_15206,N_15202);
xor U15414 (N_15414,N_15283,N_15310);
or U15415 (N_15415,N_15249,N_15271);
and U15416 (N_15416,N_15333,N_15355);
nor U15417 (N_15417,N_15274,N_15207);
xor U15418 (N_15418,N_15248,N_15210);
nand U15419 (N_15419,N_15277,N_15225);
nand U15420 (N_15420,N_15303,N_15228);
and U15421 (N_15421,N_15324,N_15328);
or U15422 (N_15422,N_15337,N_15265);
and U15423 (N_15423,N_15212,N_15356);
xor U15424 (N_15424,N_15264,N_15280);
nand U15425 (N_15425,N_15258,N_15208);
or U15426 (N_15426,N_15251,N_15255);
nand U15427 (N_15427,N_15300,N_15236);
or U15428 (N_15428,N_15226,N_15307);
and U15429 (N_15429,N_15234,N_15220);
or U15430 (N_15430,N_15238,N_15229);
and U15431 (N_15431,N_15301,N_15309);
and U15432 (N_15432,N_15266,N_15240);
and U15433 (N_15433,N_15288,N_15221);
and U15434 (N_15434,N_15284,N_15261);
and U15435 (N_15435,N_15338,N_15267);
or U15436 (N_15436,N_15204,N_15317);
and U15437 (N_15437,N_15332,N_15233);
and U15438 (N_15438,N_15336,N_15230);
xnor U15439 (N_15439,N_15316,N_15209);
or U15440 (N_15440,N_15327,N_15356);
or U15441 (N_15441,N_15238,N_15276);
nor U15442 (N_15442,N_15299,N_15219);
and U15443 (N_15443,N_15265,N_15317);
xnor U15444 (N_15444,N_15266,N_15316);
or U15445 (N_15445,N_15302,N_15245);
xnor U15446 (N_15446,N_15204,N_15287);
or U15447 (N_15447,N_15341,N_15253);
nor U15448 (N_15448,N_15343,N_15212);
or U15449 (N_15449,N_15318,N_15343);
and U15450 (N_15450,N_15357,N_15312);
nand U15451 (N_15451,N_15223,N_15324);
or U15452 (N_15452,N_15231,N_15342);
nand U15453 (N_15453,N_15230,N_15238);
nor U15454 (N_15454,N_15227,N_15300);
nor U15455 (N_15455,N_15276,N_15303);
xor U15456 (N_15456,N_15279,N_15288);
and U15457 (N_15457,N_15275,N_15342);
nand U15458 (N_15458,N_15216,N_15277);
xor U15459 (N_15459,N_15307,N_15221);
or U15460 (N_15460,N_15270,N_15309);
nor U15461 (N_15461,N_15286,N_15210);
or U15462 (N_15462,N_15203,N_15235);
nor U15463 (N_15463,N_15206,N_15353);
nor U15464 (N_15464,N_15314,N_15276);
xnor U15465 (N_15465,N_15303,N_15219);
and U15466 (N_15466,N_15355,N_15349);
nor U15467 (N_15467,N_15259,N_15350);
xor U15468 (N_15468,N_15233,N_15334);
nor U15469 (N_15469,N_15270,N_15285);
nand U15470 (N_15470,N_15236,N_15215);
or U15471 (N_15471,N_15241,N_15269);
and U15472 (N_15472,N_15330,N_15339);
or U15473 (N_15473,N_15342,N_15304);
nor U15474 (N_15474,N_15281,N_15227);
nor U15475 (N_15475,N_15213,N_15239);
nor U15476 (N_15476,N_15297,N_15284);
and U15477 (N_15477,N_15330,N_15309);
nor U15478 (N_15478,N_15294,N_15256);
or U15479 (N_15479,N_15260,N_15213);
nand U15480 (N_15480,N_15291,N_15289);
xor U15481 (N_15481,N_15301,N_15353);
or U15482 (N_15482,N_15271,N_15291);
nor U15483 (N_15483,N_15343,N_15230);
or U15484 (N_15484,N_15327,N_15217);
xnor U15485 (N_15485,N_15218,N_15249);
xnor U15486 (N_15486,N_15325,N_15259);
nand U15487 (N_15487,N_15254,N_15325);
and U15488 (N_15488,N_15267,N_15358);
and U15489 (N_15489,N_15209,N_15287);
xnor U15490 (N_15490,N_15288,N_15254);
or U15491 (N_15491,N_15305,N_15312);
or U15492 (N_15492,N_15284,N_15359);
and U15493 (N_15493,N_15354,N_15358);
and U15494 (N_15494,N_15347,N_15250);
nor U15495 (N_15495,N_15356,N_15328);
xnor U15496 (N_15496,N_15234,N_15224);
xnor U15497 (N_15497,N_15216,N_15318);
and U15498 (N_15498,N_15226,N_15317);
and U15499 (N_15499,N_15327,N_15295);
nand U15500 (N_15500,N_15315,N_15234);
xnor U15501 (N_15501,N_15230,N_15286);
and U15502 (N_15502,N_15227,N_15233);
nand U15503 (N_15503,N_15276,N_15322);
nand U15504 (N_15504,N_15231,N_15275);
xnor U15505 (N_15505,N_15227,N_15266);
nand U15506 (N_15506,N_15289,N_15305);
nand U15507 (N_15507,N_15217,N_15344);
nor U15508 (N_15508,N_15290,N_15211);
nand U15509 (N_15509,N_15250,N_15206);
nor U15510 (N_15510,N_15242,N_15236);
xor U15511 (N_15511,N_15279,N_15201);
nor U15512 (N_15512,N_15296,N_15204);
nand U15513 (N_15513,N_15347,N_15338);
xnor U15514 (N_15514,N_15299,N_15311);
nor U15515 (N_15515,N_15338,N_15310);
xor U15516 (N_15516,N_15238,N_15355);
or U15517 (N_15517,N_15203,N_15233);
and U15518 (N_15518,N_15345,N_15257);
xnor U15519 (N_15519,N_15266,N_15202);
and U15520 (N_15520,N_15487,N_15448);
nor U15521 (N_15521,N_15406,N_15443);
nor U15522 (N_15522,N_15436,N_15412);
xor U15523 (N_15523,N_15505,N_15409);
and U15524 (N_15524,N_15365,N_15441);
nor U15525 (N_15525,N_15473,N_15500);
or U15526 (N_15526,N_15425,N_15472);
nor U15527 (N_15527,N_15493,N_15435);
nand U15528 (N_15528,N_15476,N_15457);
or U15529 (N_15529,N_15369,N_15394);
nand U15530 (N_15530,N_15367,N_15494);
or U15531 (N_15531,N_15417,N_15468);
xnor U15532 (N_15532,N_15454,N_15398);
xnor U15533 (N_15533,N_15517,N_15391);
xor U15534 (N_15534,N_15501,N_15383);
nand U15535 (N_15535,N_15467,N_15363);
xor U15536 (N_15536,N_15506,N_15396);
xor U15537 (N_15537,N_15432,N_15447);
nand U15538 (N_15538,N_15478,N_15489);
nand U15539 (N_15539,N_15403,N_15361);
nand U15540 (N_15540,N_15456,N_15382);
and U15541 (N_15541,N_15381,N_15469);
xnor U15542 (N_15542,N_15449,N_15488);
nand U15543 (N_15543,N_15481,N_15480);
nor U15544 (N_15544,N_15392,N_15389);
nor U15545 (N_15545,N_15385,N_15490);
or U15546 (N_15546,N_15410,N_15519);
xnor U15547 (N_15547,N_15399,N_15428);
or U15548 (N_15548,N_15508,N_15462);
xnor U15549 (N_15549,N_15405,N_15495);
nand U15550 (N_15550,N_15444,N_15433);
or U15551 (N_15551,N_15402,N_15373);
and U15552 (N_15552,N_15516,N_15388);
or U15553 (N_15553,N_15368,N_15453);
and U15554 (N_15554,N_15491,N_15463);
and U15555 (N_15555,N_15458,N_15451);
and U15556 (N_15556,N_15423,N_15416);
nand U15557 (N_15557,N_15380,N_15475);
nand U15558 (N_15558,N_15460,N_15459);
nand U15559 (N_15559,N_15397,N_15413);
nor U15560 (N_15560,N_15440,N_15378);
xor U15561 (N_15561,N_15429,N_15513);
nand U15562 (N_15562,N_15366,N_15422);
xnor U15563 (N_15563,N_15420,N_15414);
xor U15564 (N_15564,N_15426,N_15471);
nand U15565 (N_15565,N_15502,N_15384);
or U15566 (N_15566,N_15374,N_15470);
nor U15567 (N_15567,N_15507,N_15503);
and U15568 (N_15568,N_15498,N_15484);
nand U15569 (N_15569,N_15419,N_15427);
nand U15570 (N_15570,N_15492,N_15379);
or U15571 (N_15571,N_15497,N_15465);
nand U15572 (N_15572,N_15464,N_15479);
xnor U15573 (N_15573,N_15496,N_15376);
nand U15574 (N_15574,N_15421,N_15450);
xor U15575 (N_15575,N_15375,N_15370);
nor U15576 (N_15576,N_15390,N_15499);
or U15577 (N_15577,N_15386,N_15482);
and U15578 (N_15578,N_15407,N_15438);
and U15579 (N_15579,N_15400,N_15518);
xnor U15580 (N_15580,N_15442,N_15362);
or U15581 (N_15581,N_15411,N_15418);
xor U15582 (N_15582,N_15377,N_15510);
nor U15583 (N_15583,N_15424,N_15509);
nand U15584 (N_15584,N_15485,N_15515);
and U15585 (N_15585,N_15372,N_15393);
nand U15586 (N_15586,N_15483,N_15408);
nor U15587 (N_15587,N_15461,N_15446);
nand U15588 (N_15588,N_15404,N_15511);
xnor U15589 (N_15589,N_15504,N_15486);
nor U15590 (N_15590,N_15430,N_15401);
and U15591 (N_15591,N_15437,N_15395);
and U15592 (N_15592,N_15474,N_15452);
xor U15593 (N_15593,N_15514,N_15364);
or U15594 (N_15594,N_15387,N_15512);
and U15595 (N_15595,N_15466,N_15445);
nor U15596 (N_15596,N_15360,N_15439);
xnor U15597 (N_15597,N_15477,N_15434);
and U15598 (N_15598,N_15371,N_15415);
xor U15599 (N_15599,N_15455,N_15431);
or U15600 (N_15600,N_15490,N_15510);
nor U15601 (N_15601,N_15519,N_15369);
xnor U15602 (N_15602,N_15510,N_15411);
nor U15603 (N_15603,N_15433,N_15408);
and U15604 (N_15604,N_15413,N_15478);
and U15605 (N_15605,N_15367,N_15498);
and U15606 (N_15606,N_15498,N_15362);
nor U15607 (N_15607,N_15423,N_15381);
and U15608 (N_15608,N_15411,N_15471);
nand U15609 (N_15609,N_15497,N_15385);
or U15610 (N_15610,N_15456,N_15388);
nand U15611 (N_15611,N_15508,N_15504);
or U15612 (N_15612,N_15364,N_15368);
nand U15613 (N_15613,N_15492,N_15484);
nand U15614 (N_15614,N_15375,N_15469);
xnor U15615 (N_15615,N_15477,N_15463);
or U15616 (N_15616,N_15465,N_15372);
or U15617 (N_15617,N_15515,N_15518);
nor U15618 (N_15618,N_15373,N_15385);
and U15619 (N_15619,N_15408,N_15475);
nand U15620 (N_15620,N_15434,N_15453);
xor U15621 (N_15621,N_15424,N_15416);
nand U15622 (N_15622,N_15456,N_15397);
nor U15623 (N_15623,N_15432,N_15398);
and U15624 (N_15624,N_15384,N_15482);
and U15625 (N_15625,N_15416,N_15413);
nor U15626 (N_15626,N_15426,N_15377);
nor U15627 (N_15627,N_15475,N_15407);
or U15628 (N_15628,N_15373,N_15414);
nand U15629 (N_15629,N_15473,N_15465);
xor U15630 (N_15630,N_15426,N_15438);
and U15631 (N_15631,N_15488,N_15512);
nor U15632 (N_15632,N_15455,N_15421);
and U15633 (N_15633,N_15424,N_15502);
nand U15634 (N_15634,N_15448,N_15389);
and U15635 (N_15635,N_15437,N_15402);
nor U15636 (N_15636,N_15459,N_15450);
xor U15637 (N_15637,N_15364,N_15460);
xor U15638 (N_15638,N_15463,N_15391);
and U15639 (N_15639,N_15461,N_15431);
or U15640 (N_15640,N_15441,N_15451);
nand U15641 (N_15641,N_15465,N_15444);
nor U15642 (N_15642,N_15397,N_15377);
nor U15643 (N_15643,N_15383,N_15484);
or U15644 (N_15644,N_15418,N_15472);
xor U15645 (N_15645,N_15458,N_15516);
nand U15646 (N_15646,N_15414,N_15419);
xnor U15647 (N_15647,N_15480,N_15443);
xor U15648 (N_15648,N_15364,N_15360);
nor U15649 (N_15649,N_15445,N_15438);
nor U15650 (N_15650,N_15375,N_15502);
xnor U15651 (N_15651,N_15428,N_15397);
and U15652 (N_15652,N_15511,N_15472);
nor U15653 (N_15653,N_15394,N_15474);
nor U15654 (N_15654,N_15479,N_15482);
and U15655 (N_15655,N_15467,N_15470);
or U15656 (N_15656,N_15478,N_15456);
xor U15657 (N_15657,N_15419,N_15445);
xnor U15658 (N_15658,N_15496,N_15508);
or U15659 (N_15659,N_15466,N_15495);
xor U15660 (N_15660,N_15403,N_15395);
xor U15661 (N_15661,N_15457,N_15516);
and U15662 (N_15662,N_15437,N_15445);
and U15663 (N_15663,N_15496,N_15397);
xor U15664 (N_15664,N_15388,N_15483);
nand U15665 (N_15665,N_15432,N_15468);
or U15666 (N_15666,N_15369,N_15413);
xnor U15667 (N_15667,N_15443,N_15362);
or U15668 (N_15668,N_15415,N_15384);
nor U15669 (N_15669,N_15507,N_15492);
nand U15670 (N_15670,N_15439,N_15487);
and U15671 (N_15671,N_15465,N_15396);
nand U15672 (N_15672,N_15463,N_15379);
and U15673 (N_15673,N_15468,N_15423);
xor U15674 (N_15674,N_15369,N_15431);
xor U15675 (N_15675,N_15374,N_15508);
or U15676 (N_15676,N_15477,N_15432);
nand U15677 (N_15677,N_15501,N_15479);
nor U15678 (N_15678,N_15400,N_15472);
or U15679 (N_15679,N_15468,N_15418);
nand U15680 (N_15680,N_15609,N_15629);
and U15681 (N_15681,N_15530,N_15624);
xor U15682 (N_15682,N_15595,N_15584);
nor U15683 (N_15683,N_15636,N_15621);
or U15684 (N_15684,N_15635,N_15578);
or U15685 (N_15685,N_15658,N_15520);
or U15686 (N_15686,N_15572,N_15529);
or U15687 (N_15687,N_15582,N_15558);
or U15688 (N_15688,N_15649,N_15587);
or U15689 (N_15689,N_15583,N_15652);
nor U15690 (N_15690,N_15677,N_15574);
nand U15691 (N_15691,N_15620,N_15640);
nor U15692 (N_15692,N_15653,N_15638);
or U15693 (N_15693,N_15596,N_15622);
nor U15694 (N_15694,N_15548,N_15580);
or U15695 (N_15695,N_15538,N_15553);
nor U15696 (N_15696,N_15675,N_15614);
nand U15697 (N_15697,N_15656,N_15570);
or U15698 (N_15698,N_15546,N_15642);
and U15699 (N_15699,N_15554,N_15589);
or U15700 (N_15700,N_15634,N_15523);
or U15701 (N_15701,N_15567,N_15559);
or U15702 (N_15702,N_15571,N_15605);
nand U15703 (N_15703,N_15674,N_15602);
and U15704 (N_15704,N_15611,N_15631);
nor U15705 (N_15705,N_15664,N_15542);
or U15706 (N_15706,N_15632,N_15657);
or U15707 (N_15707,N_15627,N_15628);
nand U15708 (N_15708,N_15637,N_15557);
nor U15709 (N_15709,N_15678,N_15537);
xnor U15710 (N_15710,N_15599,N_15643);
nand U15711 (N_15711,N_15598,N_15618);
and U15712 (N_15712,N_15579,N_15650);
nand U15713 (N_15713,N_15594,N_15575);
and U15714 (N_15714,N_15528,N_15607);
nand U15715 (N_15715,N_15564,N_15532);
nor U15716 (N_15716,N_15612,N_15556);
and U15717 (N_15717,N_15534,N_15562);
and U15718 (N_15718,N_15531,N_15619);
and U15719 (N_15719,N_15646,N_15647);
xnor U15720 (N_15720,N_15566,N_15610);
and U15721 (N_15721,N_15616,N_15669);
nor U15722 (N_15722,N_15617,N_15521);
nor U15723 (N_15723,N_15591,N_15670);
nor U15724 (N_15724,N_15539,N_15568);
and U15725 (N_15725,N_15590,N_15565);
and U15726 (N_15726,N_15525,N_15645);
and U15727 (N_15727,N_15577,N_15588);
nor U15728 (N_15728,N_15641,N_15644);
or U15729 (N_15729,N_15555,N_15608);
or U15730 (N_15730,N_15552,N_15673);
nand U15731 (N_15731,N_15547,N_15604);
or U15732 (N_15732,N_15626,N_15600);
nand U15733 (N_15733,N_15625,N_15551);
xor U15734 (N_15734,N_15550,N_15639);
nor U15735 (N_15735,N_15623,N_15662);
nand U15736 (N_15736,N_15661,N_15601);
nor U15737 (N_15737,N_15593,N_15654);
xnor U15738 (N_15738,N_15633,N_15671);
xnor U15739 (N_15739,N_15543,N_15592);
xor U15740 (N_15740,N_15597,N_15659);
or U15741 (N_15741,N_15660,N_15545);
nor U15742 (N_15742,N_15561,N_15667);
nand U15743 (N_15743,N_15651,N_15524);
or U15744 (N_15744,N_15603,N_15576);
nor U15745 (N_15745,N_15549,N_15668);
xor U15746 (N_15746,N_15581,N_15615);
nor U15747 (N_15747,N_15679,N_15655);
or U15748 (N_15748,N_15540,N_15665);
xnor U15749 (N_15749,N_15544,N_15573);
or U15750 (N_15750,N_15522,N_15663);
and U15751 (N_15751,N_15630,N_15613);
or U15752 (N_15752,N_15536,N_15533);
nor U15753 (N_15753,N_15541,N_15569);
xor U15754 (N_15754,N_15586,N_15606);
nor U15755 (N_15755,N_15648,N_15526);
nand U15756 (N_15756,N_15666,N_15527);
nor U15757 (N_15757,N_15676,N_15563);
nand U15758 (N_15758,N_15535,N_15585);
or U15759 (N_15759,N_15560,N_15672);
nor U15760 (N_15760,N_15673,N_15644);
nor U15761 (N_15761,N_15544,N_15638);
nand U15762 (N_15762,N_15648,N_15520);
nor U15763 (N_15763,N_15661,N_15617);
and U15764 (N_15764,N_15665,N_15625);
and U15765 (N_15765,N_15565,N_15615);
or U15766 (N_15766,N_15671,N_15580);
nor U15767 (N_15767,N_15552,N_15630);
and U15768 (N_15768,N_15628,N_15647);
nand U15769 (N_15769,N_15601,N_15643);
and U15770 (N_15770,N_15581,N_15587);
nor U15771 (N_15771,N_15622,N_15630);
xor U15772 (N_15772,N_15618,N_15611);
nand U15773 (N_15773,N_15644,N_15616);
nor U15774 (N_15774,N_15596,N_15605);
or U15775 (N_15775,N_15563,N_15624);
or U15776 (N_15776,N_15553,N_15587);
xor U15777 (N_15777,N_15575,N_15560);
nand U15778 (N_15778,N_15601,N_15679);
nor U15779 (N_15779,N_15573,N_15539);
nand U15780 (N_15780,N_15564,N_15548);
nand U15781 (N_15781,N_15596,N_15612);
xnor U15782 (N_15782,N_15563,N_15626);
nand U15783 (N_15783,N_15520,N_15544);
xnor U15784 (N_15784,N_15605,N_15663);
or U15785 (N_15785,N_15654,N_15565);
and U15786 (N_15786,N_15677,N_15606);
nand U15787 (N_15787,N_15679,N_15599);
nor U15788 (N_15788,N_15581,N_15558);
nor U15789 (N_15789,N_15545,N_15653);
and U15790 (N_15790,N_15578,N_15588);
or U15791 (N_15791,N_15623,N_15650);
or U15792 (N_15792,N_15532,N_15563);
and U15793 (N_15793,N_15661,N_15637);
xor U15794 (N_15794,N_15612,N_15520);
xor U15795 (N_15795,N_15527,N_15553);
or U15796 (N_15796,N_15564,N_15627);
nand U15797 (N_15797,N_15632,N_15641);
nand U15798 (N_15798,N_15667,N_15574);
and U15799 (N_15799,N_15592,N_15544);
nor U15800 (N_15800,N_15654,N_15656);
xor U15801 (N_15801,N_15638,N_15547);
and U15802 (N_15802,N_15624,N_15639);
nor U15803 (N_15803,N_15555,N_15535);
nor U15804 (N_15804,N_15589,N_15625);
and U15805 (N_15805,N_15545,N_15603);
nor U15806 (N_15806,N_15592,N_15550);
nor U15807 (N_15807,N_15544,N_15570);
or U15808 (N_15808,N_15521,N_15649);
nand U15809 (N_15809,N_15602,N_15589);
or U15810 (N_15810,N_15605,N_15528);
or U15811 (N_15811,N_15529,N_15585);
and U15812 (N_15812,N_15543,N_15532);
nor U15813 (N_15813,N_15551,N_15636);
nor U15814 (N_15814,N_15612,N_15609);
and U15815 (N_15815,N_15647,N_15659);
nor U15816 (N_15816,N_15648,N_15596);
nand U15817 (N_15817,N_15660,N_15533);
and U15818 (N_15818,N_15671,N_15531);
or U15819 (N_15819,N_15642,N_15533);
or U15820 (N_15820,N_15557,N_15520);
nor U15821 (N_15821,N_15539,N_15530);
nand U15822 (N_15822,N_15625,N_15664);
xnor U15823 (N_15823,N_15619,N_15641);
and U15824 (N_15824,N_15674,N_15569);
or U15825 (N_15825,N_15624,N_15568);
and U15826 (N_15826,N_15668,N_15645);
and U15827 (N_15827,N_15678,N_15668);
nand U15828 (N_15828,N_15603,N_15556);
nand U15829 (N_15829,N_15520,N_15575);
and U15830 (N_15830,N_15557,N_15620);
and U15831 (N_15831,N_15582,N_15608);
and U15832 (N_15832,N_15567,N_15637);
xnor U15833 (N_15833,N_15532,N_15617);
nor U15834 (N_15834,N_15608,N_15547);
and U15835 (N_15835,N_15529,N_15592);
xnor U15836 (N_15836,N_15574,N_15594);
nor U15837 (N_15837,N_15615,N_15528);
nor U15838 (N_15838,N_15610,N_15633);
xor U15839 (N_15839,N_15620,N_15583);
nor U15840 (N_15840,N_15788,N_15722);
xnor U15841 (N_15841,N_15829,N_15725);
nor U15842 (N_15842,N_15783,N_15692);
nor U15843 (N_15843,N_15735,N_15814);
nand U15844 (N_15844,N_15716,N_15750);
or U15845 (N_15845,N_15701,N_15693);
nor U15846 (N_15846,N_15766,N_15773);
nor U15847 (N_15847,N_15708,N_15782);
xor U15848 (N_15848,N_15820,N_15821);
nor U15849 (N_15849,N_15792,N_15784);
or U15850 (N_15850,N_15752,N_15724);
nand U15851 (N_15851,N_15819,N_15823);
nor U15852 (N_15852,N_15780,N_15777);
or U15853 (N_15853,N_15713,N_15700);
and U15854 (N_15854,N_15739,N_15738);
xor U15855 (N_15855,N_15786,N_15745);
or U15856 (N_15856,N_15791,N_15753);
or U15857 (N_15857,N_15680,N_15808);
nand U15858 (N_15858,N_15754,N_15732);
or U15859 (N_15859,N_15683,N_15800);
xor U15860 (N_15860,N_15838,N_15710);
xnor U15861 (N_15861,N_15768,N_15833);
nor U15862 (N_15862,N_15759,N_15822);
or U15863 (N_15863,N_15825,N_15801);
xor U15864 (N_15864,N_15761,N_15682);
or U15865 (N_15865,N_15815,N_15699);
nand U15866 (N_15866,N_15771,N_15781);
or U15867 (N_15867,N_15685,N_15799);
and U15868 (N_15868,N_15764,N_15830);
and U15869 (N_15869,N_15807,N_15796);
nand U15870 (N_15870,N_15778,N_15810);
nor U15871 (N_15871,N_15737,N_15828);
nand U15872 (N_15872,N_15795,N_15748);
xor U15873 (N_15873,N_15703,N_15787);
and U15874 (N_15874,N_15695,N_15718);
nand U15875 (N_15875,N_15818,N_15751);
or U15876 (N_15876,N_15803,N_15834);
nand U15877 (N_15877,N_15756,N_15690);
nand U15878 (N_15878,N_15811,N_15704);
nor U15879 (N_15879,N_15826,N_15714);
or U15880 (N_15880,N_15733,N_15736);
nand U15881 (N_15881,N_15698,N_15762);
nand U15882 (N_15882,N_15793,N_15746);
xnor U15883 (N_15883,N_15809,N_15835);
nand U15884 (N_15884,N_15757,N_15749);
xnor U15885 (N_15885,N_15707,N_15711);
and U15886 (N_15886,N_15785,N_15839);
or U15887 (N_15887,N_15794,N_15741);
and U15888 (N_15888,N_15790,N_15717);
or U15889 (N_15889,N_15687,N_15758);
xnor U15890 (N_15890,N_15691,N_15805);
nor U15891 (N_15891,N_15775,N_15686);
or U15892 (N_15892,N_15681,N_15767);
or U15893 (N_15893,N_15817,N_15696);
xnor U15894 (N_15894,N_15776,N_15744);
nand U15895 (N_15895,N_15726,N_15727);
or U15896 (N_15896,N_15772,N_15813);
nand U15897 (N_15897,N_15719,N_15702);
and U15898 (N_15898,N_15730,N_15789);
and U15899 (N_15899,N_15731,N_15774);
xnor U15900 (N_15900,N_15721,N_15779);
nor U15901 (N_15901,N_15769,N_15715);
or U15902 (N_15902,N_15802,N_15684);
nor U15903 (N_15903,N_15709,N_15740);
nor U15904 (N_15904,N_15755,N_15806);
nor U15905 (N_15905,N_15712,N_15697);
nor U15906 (N_15906,N_15694,N_15760);
nand U15907 (N_15907,N_15836,N_15705);
nand U15908 (N_15908,N_15770,N_15723);
and U15909 (N_15909,N_15812,N_15765);
nand U15910 (N_15910,N_15720,N_15763);
xnor U15911 (N_15911,N_15729,N_15734);
and U15912 (N_15912,N_15816,N_15831);
nor U15913 (N_15913,N_15824,N_15747);
and U15914 (N_15914,N_15688,N_15804);
xor U15915 (N_15915,N_15728,N_15706);
or U15916 (N_15916,N_15827,N_15742);
xnor U15917 (N_15917,N_15832,N_15743);
nand U15918 (N_15918,N_15689,N_15797);
or U15919 (N_15919,N_15837,N_15798);
nand U15920 (N_15920,N_15806,N_15694);
nor U15921 (N_15921,N_15718,N_15749);
and U15922 (N_15922,N_15810,N_15772);
and U15923 (N_15923,N_15767,N_15742);
xor U15924 (N_15924,N_15702,N_15772);
and U15925 (N_15925,N_15697,N_15747);
xor U15926 (N_15926,N_15808,N_15771);
xnor U15927 (N_15927,N_15744,N_15689);
xor U15928 (N_15928,N_15689,N_15688);
nand U15929 (N_15929,N_15717,N_15839);
nor U15930 (N_15930,N_15816,N_15778);
xor U15931 (N_15931,N_15803,N_15712);
xor U15932 (N_15932,N_15818,N_15715);
and U15933 (N_15933,N_15735,N_15804);
nand U15934 (N_15934,N_15784,N_15780);
or U15935 (N_15935,N_15762,N_15757);
xnor U15936 (N_15936,N_15810,N_15795);
xor U15937 (N_15937,N_15696,N_15768);
xor U15938 (N_15938,N_15775,N_15744);
and U15939 (N_15939,N_15701,N_15719);
or U15940 (N_15940,N_15831,N_15766);
or U15941 (N_15941,N_15801,N_15717);
and U15942 (N_15942,N_15834,N_15785);
xor U15943 (N_15943,N_15755,N_15692);
nor U15944 (N_15944,N_15767,N_15693);
or U15945 (N_15945,N_15807,N_15701);
nand U15946 (N_15946,N_15733,N_15763);
or U15947 (N_15947,N_15827,N_15733);
or U15948 (N_15948,N_15719,N_15748);
nor U15949 (N_15949,N_15749,N_15786);
nor U15950 (N_15950,N_15720,N_15751);
nor U15951 (N_15951,N_15730,N_15690);
nor U15952 (N_15952,N_15820,N_15707);
xnor U15953 (N_15953,N_15821,N_15708);
xor U15954 (N_15954,N_15804,N_15704);
nor U15955 (N_15955,N_15693,N_15804);
and U15956 (N_15956,N_15696,N_15686);
xnor U15957 (N_15957,N_15728,N_15822);
nand U15958 (N_15958,N_15747,N_15688);
or U15959 (N_15959,N_15819,N_15826);
nor U15960 (N_15960,N_15681,N_15834);
or U15961 (N_15961,N_15831,N_15807);
and U15962 (N_15962,N_15835,N_15810);
nor U15963 (N_15963,N_15693,N_15745);
and U15964 (N_15964,N_15833,N_15775);
and U15965 (N_15965,N_15761,N_15803);
and U15966 (N_15966,N_15708,N_15742);
or U15967 (N_15967,N_15749,N_15799);
nand U15968 (N_15968,N_15798,N_15776);
nand U15969 (N_15969,N_15838,N_15744);
and U15970 (N_15970,N_15748,N_15760);
and U15971 (N_15971,N_15757,N_15784);
nand U15972 (N_15972,N_15790,N_15686);
and U15973 (N_15973,N_15789,N_15739);
nand U15974 (N_15974,N_15753,N_15816);
xor U15975 (N_15975,N_15766,N_15741);
xor U15976 (N_15976,N_15837,N_15755);
nand U15977 (N_15977,N_15781,N_15791);
and U15978 (N_15978,N_15783,N_15751);
xnor U15979 (N_15979,N_15835,N_15749);
xor U15980 (N_15980,N_15704,N_15751);
or U15981 (N_15981,N_15700,N_15694);
nor U15982 (N_15982,N_15694,N_15809);
or U15983 (N_15983,N_15792,N_15731);
nor U15984 (N_15984,N_15836,N_15769);
or U15985 (N_15985,N_15766,N_15769);
or U15986 (N_15986,N_15795,N_15744);
and U15987 (N_15987,N_15685,N_15711);
nand U15988 (N_15988,N_15839,N_15746);
nor U15989 (N_15989,N_15829,N_15790);
or U15990 (N_15990,N_15764,N_15790);
nand U15991 (N_15991,N_15772,N_15734);
and U15992 (N_15992,N_15720,N_15738);
or U15993 (N_15993,N_15818,N_15810);
or U15994 (N_15994,N_15774,N_15788);
nand U15995 (N_15995,N_15707,N_15792);
and U15996 (N_15996,N_15768,N_15692);
nand U15997 (N_15997,N_15836,N_15802);
or U15998 (N_15998,N_15735,N_15728);
nor U15999 (N_15999,N_15680,N_15836);
nor U16000 (N_16000,N_15907,N_15853);
nor U16001 (N_16001,N_15955,N_15997);
nor U16002 (N_16002,N_15916,N_15963);
or U16003 (N_16003,N_15967,N_15867);
nor U16004 (N_16004,N_15979,N_15868);
or U16005 (N_16005,N_15993,N_15861);
and U16006 (N_16006,N_15879,N_15975);
or U16007 (N_16007,N_15902,N_15931);
or U16008 (N_16008,N_15924,N_15982);
or U16009 (N_16009,N_15923,N_15855);
nor U16010 (N_16010,N_15893,N_15912);
or U16011 (N_16011,N_15968,N_15960);
or U16012 (N_16012,N_15922,N_15872);
nor U16013 (N_16013,N_15978,N_15899);
nand U16014 (N_16014,N_15998,N_15952);
nor U16015 (N_16015,N_15886,N_15911);
or U16016 (N_16016,N_15987,N_15949);
xnor U16017 (N_16017,N_15841,N_15986);
xnor U16018 (N_16018,N_15896,N_15973);
nand U16019 (N_16019,N_15983,N_15969);
nand U16020 (N_16020,N_15870,N_15958);
nand U16021 (N_16021,N_15898,N_15883);
nand U16022 (N_16022,N_15876,N_15992);
or U16023 (N_16023,N_15903,N_15890);
nand U16024 (N_16024,N_15974,N_15858);
nor U16025 (N_16025,N_15873,N_15909);
and U16026 (N_16026,N_15932,N_15844);
nand U16027 (N_16027,N_15878,N_15892);
and U16028 (N_16028,N_15865,N_15927);
or U16029 (N_16029,N_15863,N_15919);
and U16030 (N_16030,N_15864,N_15926);
xnor U16031 (N_16031,N_15985,N_15970);
nand U16032 (N_16032,N_15869,N_15906);
and U16033 (N_16033,N_15947,N_15951);
nor U16034 (N_16034,N_15887,N_15846);
xor U16035 (N_16035,N_15891,N_15905);
nor U16036 (N_16036,N_15980,N_15943);
nand U16037 (N_16037,N_15850,N_15874);
and U16038 (N_16038,N_15920,N_15981);
or U16039 (N_16039,N_15957,N_15964);
nor U16040 (N_16040,N_15971,N_15877);
xnor U16041 (N_16041,N_15989,N_15999);
and U16042 (N_16042,N_15965,N_15945);
xnor U16043 (N_16043,N_15953,N_15908);
nor U16044 (N_16044,N_15847,N_15935);
and U16045 (N_16045,N_15882,N_15984);
nor U16046 (N_16046,N_15894,N_15950);
nand U16047 (N_16047,N_15954,N_15994);
xor U16048 (N_16048,N_15862,N_15852);
or U16049 (N_16049,N_15866,N_15854);
or U16050 (N_16050,N_15845,N_15930);
nand U16051 (N_16051,N_15996,N_15995);
or U16052 (N_16052,N_15842,N_15940);
nor U16053 (N_16053,N_15959,N_15962);
xor U16054 (N_16054,N_15961,N_15881);
and U16055 (N_16055,N_15988,N_15897);
and U16056 (N_16056,N_15910,N_15918);
or U16057 (N_16057,N_15929,N_15904);
or U16058 (N_16058,N_15936,N_15848);
or U16059 (N_16059,N_15956,N_15888);
and U16060 (N_16060,N_15991,N_15946);
nor U16061 (N_16061,N_15843,N_15915);
xor U16062 (N_16062,N_15859,N_15851);
nor U16063 (N_16063,N_15928,N_15857);
nor U16064 (N_16064,N_15933,N_15917);
and U16065 (N_16065,N_15934,N_15913);
and U16066 (N_16066,N_15939,N_15885);
xnor U16067 (N_16067,N_15942,N_15990);
and U16068 (N_16068,N_15880,N_15944);
xnor U16069 (N_16069,N_15871,N_15977);
and U16070 (N_16070,N_15938,N_15925);
or U16071 (N_16071,N_15856,N_15976);
nand U16072 (N_16072,N_15840,N_15921);
and U16073 (N_16073,N_15914,N_15937);
nor U16074 (N_16074,N_15889,N_15849);
and U16075 (N_16075,N_15948,N_15895);
and U16076 (N_16076,N_15941,N_15901);
nand U16077 (N_16077,N_15900,N_15875);
and U16078 (N_16078,N_15966,N_15972);
or U16079 (N_16079,N_15884,N_15860);
nor U16080 (N_16080,N_15888,N_15915);
or U16081 (N_16081,N_15953,N_15866);
or U16082 (N_16082,N_15973,N_15920);
xor U16083 (N_16083,N_15878,N_15930);
xnor U16084 (N_16084,N_15897,N_15874);
and U16085 (N_16085,N_15993,N_15855);
nand U16086 (N_16086,N_15887,N_15955);
nand U16087 (N_16087,N_15886,N_15884);
nor U16088 (N_16088,N_15896,N_15917);
and U16089 (N_16089,N_15866,N_15990);
nor U16090 (N_16090,N_15959,N_15886);
nor U16091 (N_16091,N_15886,N_15906);
nor U16092 (N_16092,N_15973,N_15881);
and U16093 (N_16093,N_15977,N_15864);
or U16094 (N_16094,N_15972,N_15883);
nor U16095 (N_16095,N_15889,N_15925);
and U16096 (N_16096,N_15977,N_15992);
xor U16097 (N_16097,N_15999,N_15988);
and U16098 (N_16098,N_15874,N_15918);
xnor U16099 (N_16099,N_15924,N_15894);
nor U16100 (N_16100,N_15941,N_15911);
and U16101 (N_16101,N_15864,N_15840);
nand U16102 (N_16102,N_15972,N_15886);
nor U16103 (N_16103,N_15856,N_15956);
nand U16104 (N_16104,N_15920,N_15963);
and U16105 (N_16105,N_15914,N_15969);
xor U16106 (N_16106,N_15917,N_15874);
nor U16107 (N_16107,N_15868,N_15910);
xnor U16108 (N_16108,N_15930,N_15847);
and U16109 (N_16109,N_15840,N_15936);
xor U16110 (N_16110,N_15861,N_15957);
nor U16111 (N_16111,N_15842,N_15854);
and U16112 (N_16112,N_15916,N_15976);
and U16113 (N_16113,N_15979,N_15962);
nor U16114 (N_16114,N_15865,N_15850);
nand U16115 (N_16115,N_15903,N_15907);
and U16116 (N_16116,N_15905,N_15850);
or U16117 (N_16117,N_15892,N_15885);
nand U16118 (N_16118,N_15961,N_15906);
and U16119 (N_16119,N_15910,N_15992);
and U16120 (N_16120,N_15999,N_15943);
nand U16121 (N_16121,N_15992,N_15903);
or U16122 (N_16122,N_15964,N_15908);
xnor U16123 (N_16123,N_15873,N_15978);
xor U16124 (N_16124,N_15918,N_15986);
or U16125 (N_16125,N_15845,N_15995);
nor U16126 (N_16126,N_15981,N_15945);
nor U16127 (N_16127,N_15982,N_15931);
xnor U16128 (N_16128,N_15967,N_15952);
nand U16129 (N_16129,N_15967,N_15908);
xor U16130 (N_16130,N_15876,N_15893);
or U16131 (N_16131,N_15958,N_15995);
nor U16132 (N_16132,N_15890,N_15854);
xnor U16133 (N_16133,N_15887,N_15938);
and U16134 (N_16134,N_15955,N_15854);
or U16135 (N_16135,N_15951,N_15940);
and U16136 (N_16136,N_15917,N_15885);
xnor U16137 (N_16137,N_15982,N_15962);
xor U16138 (N_16138,N_15866,N_15940);
or U16139 (N_16139,N_15846,N_15974);
and U16140 (N_16140,N_15986,N_15882);
and U16141 (N_16141,N_15910,N_15955);
nor U16142 (N_16142,N_15920,N_15900);
nor U16143 (N_16143,N_15906,N_15841);
nor U16144 (N_16144,N_15959,N_15873);
or U16145 (N_16145,N_15978,N_15853);
nand U16146 (N_16146,N_15905,N_15841);
nand U16147 (N_16147,N_15985,N_15913);
and U16148 (N_16148,N_15896,N_15853);
and U16149 (N_16149,N_15942,N_15860);
or U16150 (N_16150,N_15858,N_15939);
or U16151 (N_16151,N_15933,N_15910);
xnor U16152 (N_16152,N_15949,N_15875);
xnor U16153 (N_16153,N_15988,N_15962);
or U16154 (N_16154,N_15978,N_15842);
nand U16155 (N_16155,N_15995,N_15993);
nand U16156 (N_16156,N_15921,N_15974);
nor U16157 (N_16157,N_15939,N_15877);
nor U16158 (N_16158,N_15965,N_15857);
nor U16159 (N_16159,N_15934,N_15858);
xnor U16160 (N_16160,N_16045,N_16134);
xor U16161 (N_16161,N_16046,N_16070);
or U16162 (N_16162,N_16138,N_16128);
or U16163 (N_16163,N_16145,N_16039);
or U16164 (N_16164,N_16006,N_16086);
xor U16165 (N_16165,N_16021,N_16109);
or U16166 (N_16166,N_16088,N_16118);
xor U16167 (N_16167,N_16065,N_16015);
and U16168 (N_16168,N_16028,N_16114);
or U16169 (N_16169,N_16056,N_16147);
nand U16170 (N_16170,N_16076,N_16053);
nand U16171 (N_16171,N_16071,N_16064);
nor U16172 (N_16172,N_16089,N_16063);
or U16173 (N_16173,N_16069,N_16054);
nor U16174 (N_16174,N_16004,N_16016);
nand U16175 (N_16175,N_16115,N_16121);
nand U16176 (N_16176,N_16062,N_16023);
or U16177 (N_16177,N_16058,N_16090);
and U16178 (N_16178,N_16117,N_16130);
or U16179 (N_16179,N_16119,N_16080);
nor U16180 (N_16180,N_16129,N_16029);
xnor U16181 (N_16181,N_16135,N_16074);
nand U16182 (N_16182,N_16024,N_16104);
and U16183 (N_16183,N_16132,N_16124);
nor U16184 (N_16184,N_16051,N_16018);
nand U16185 (N_16185,N_16055,N_16050);
nor U16186 (N_16186,N_16150,N_16013);
nand U16187 (N_16187,N_16011,N_16068);
xor U16188 (N_16188,N_16151,N_16096);
or U16189 (N_16189,N_16008,N_16093);
xor U16190 (N_16190,N_16052,N_16105);
or U16191 (N_16191,N_16042,N_16146);
nand U16192 (N_16192,N_16005,N_16126);
xnor U16193 (N_16193,N_16154,N_16047);
and U16194 (N_16194,N_16014,N_16033);
nor U16195 (N_16195,N_16152,N_16082);
nand U16196 (N_16196,N_16144,N_16048);
nor U16197 (N_16197,N_16035,N_16116);
or U16198 (N_16198,N_16001,N_16155);
nor U16199 (N_16199,N_16103,N_16097);
and U16200 (N_16200,N_16084,N_16111);
and U16201 (N_16201,N_16106,N_16060);
nand U16202 (N_16202,N_16112,N_16007);
or U16203 (N_16203,N_16153,N_16139);
xnor U16204 (N_16204,N_16000,N_16072);
or U16205 (N_16205,N_16022,N_16158);
xor U16206 (N_16206,N_16057,N_16102);
nor U16207 (N_16207,N_16123,N_16079);
nor U16208 (N_16208,N_16131,N_16003);
nand U16209 (N_16209,N_16020,N_16059);
nand U16210 (N_16210,N_16113,N_16012);
nand U16211 (N_16211,N_16085,N_16099);
nand U16212 (N_16212,N_16075,N_16002);
xor U16213 (N_16213,N_16078,N_16087);
and U16214 (N_16214,N_16032,N_16061);
or U16215 (N_16215,N_16136,N_16067);
or U16216 (N_16216,N_16027,N_16140);
xor U16217 (N_16217,N_16141,N_16125);
and U16218 (N_16218,N_16049,N_16100);
nand U16219 (N_16219,N_16083,N_16092);
nand U16220 (N_16220,N_16041,N_16043);
nor U16221 (N_16221,N_16037,N_16077);
xor U16222 (N_16222,N_16010,N_16019);
or U16223 (N_16223,N_16156,N_16122);
or U16224 (N_16224,N_16036,N_16142);
and U16225 (N_16225,N_16009,N_16017);
nor U16226 (N_16226,N_16081,N_16159);
nor U16227 (N_16227,N_16094,N_16133);
or U16228 (N_16228,N_16073,N_16034);
and U16229 (N_16229,N_16025,N_16108);
and U16230 (N_16230,N_16143,N_16157);
nand U16231 (N_16231,N_16127,N_16120);
nor U16232 (N_16232,N_16107,N_16044);
nor U16233 (N_16233,N_16110,N_16101);
nor U16234 (N_16234,N_16040,N_16149);
nor U16235 (N_16235,N_16091,N_16095);
nand U16236 (N_16236,N_16066,N_16098);
or U16237 (N_16237,N_16148,N_16026);
nand U16238 (N_16238,N_16031,N_16038);
nand U16239 (N_16239,N_16030,N_16137);
xor U16240 (N_16240,N_16132,N_16081);
or U16241 (N_16241,N_16056,N_16089);
nor U16242 (N_16242,N_16131,N_16116);
and U16243 (N_16243,N_16019,N_16151);
and U16244 (N_16244,N_16078,N_16128);
nor U16245 (N_16245,N_16065,N_16111);
xor U16246 (N_16246,N_16078,N_16013);
nand U16247 (N_16247,N_16082,N_16150);
xor U16248 (N_16248,N_16068,N_16040);
or U16249 (N_16249,N_16009,N_16132);
or U16250 (N_16250,N_16121,N_16015);
xor U16251 (N_16251,N_16022,N_16130);
and U16252 (N_16252,N_16036,N_16038);
or U16253 (N_16253,N_16060,N_16038);
xnor U16254 (N_16254,N_16054,N_16094);
xnor U16255 (N_16255,N_16060,N_16103);
or U16256 (N_16256,N_16038,N_16012);
or U16257 (N_16257,N_16080,N_16028);
nor U16258 (N_16258,N_16140,N_16098);
nor U16259 (N_16259,N_16153,N_16150);
xnor U16260 (N_16260,N_16031,N_16013);
nand U16261 (N_16261,N_16159,N_16044);
or U16262 (N_16262,N_16094,N_16154);
xnor U16263 (N_16263,N_16075,N_16027);
xor U16264 (N_16264,N_16126,N_16157);
nor U16265 (N_16265,N_16013,N_16118);
or U16266 (N_16266,N_16059,N_16030);
and U16267 (N_16267,N_16078,N_16148);
nand U16268 (N_16268,N_16011,N_16138);
nor U16269 (N_16269,N_16007,N_16080);
nor U16270 (N_16270,N_16146,N_16089);
nor U16271 (N_16271,N_16139,N_16096);
xor U16272 (N_16272,N_16044,N_16105);
nand U16273 (N_16273,N_16025,N_16061);
and U16274 (N_16274,N_16020,N_16083);
nor U16275 (N_16275,N_16151,N_16003);
nor U16276 (N_16276,N_16103,N_16135);
or U16277 (N_16277,N_16157,N_16125);
nand U16278 (N_16278,N_16080,N_16092);
nor U16279 (N_16279,N_16130,N_16052);
or U16280 (N_16280,N_16115,N_16041);
nand U16281 (N_16281,N_16129,N_16156);
or U16282 (N_16282,N_16035,N_16069);
and U16283 (N_16283,N_16159,N_16098);
nand U16284 (N_16284,N_16137,N_16045);
nand U16285 (N_16285,N_16152,N_16052);
xnor U16286 (N_16286,N_16040,N_16070);
nor U16287 (N_16287,N_16127,N_16039);
nor U16288 (N_16288,N_16093,N_16144);
xor U16289 (N_16289,N_16079,N_16129);
and U16290 (N_16290,N_16043,N_16119);
nor U16291 (N_16291,N_16054,N_16144);
or U16292 (N_16292,N_16152,N_16147);
xor U16293 (N_16293,N_16029,N_16069);
or U16294 (N_16294,N_16135,N_16036);
or U16295 (N_16295,N_16019,N_16120);
nand U16296 (N_16296,N_16006,N_16077);
or U16297 (N_16297,N_16116,N_16056);
nand U16298 (N_16298,N_16125,N_16154);
xor U16299 (N_16299,N_16076,N_16086);
xnor U16300 (N_16300,N_16025,N_16111);
nand U16301 (N_16301,N_16140,N_16026);
nand U16302 (N_16302,N_16052,N_16071);
xor U16303 (N_16303,N_16084,N_16020);
or U16304 (N_16304,N_16128,N_16058);
xor U16305 (N_16305,N_16044,N_16095);
and U16306 (N_16306,N_16101,N_16103);
nor U16307 (N_16307,N_16150,N_16110);
and U16308 (N_16308,N_16098,N_16030);
or U16309 (N_16309,N_16122,N_16141);
or U16310 (N_16310,N_16022,N_16083);
nor U16311 (N_16311,N_16090,N_16022);
or U16312 (N_16312,N_16047,N_16139);
xor U16313 (N_16313,N_16085,N_16084);
or U16314 (N_16314,N_16028,N_16099);
and U16315 (N_16315,N_16062,N_16095);
and U16316 (N_16316,N_16103,N_16026);
nand U16317 (N_16317,N_16112,N_16070);
and U16318 (N_16318,N_16024,N_16154);
nand U16319 (N_16319,N_16099,N_16011);
nor U16320 (N_16320,N_16177,N_16243);
nand U16321 (N_16321,N_16253,N_16160);
nand U16322 (N_16322,N_16302,N_16292);
and U16323 (N_16323,N_16260,N_16319);
nor U16324 (N_16324,N_16267,N_16247);
xor U16325 (N_16325,N_16284,N_16301);
and U16326 (N_16326,N_16303,N_16208);
or U16327 (N_16327,N_16236,N_16297);
xnor U16328 (N_16328,N_16308,N_16300);
nand U16329 (N_16329,N_16161,N_16274);
nor U16330 (N_16330,N_16310,N_16254);
xnor U16331 (N_16331,N_16212,N_16235);
or U16332 (N_16332,N_16217,N_16224);
and U16333 (N_16333,N_16198,N_16172);
nor U16334 (N_16334,N_16227,N_16252);
nand U16335 (N_16335,N_16196,N_16268);
and U16336 (N_16336,N_16294,N_16277);
xnor U16337 (N_16337,N_16289,N_16186);
nand U16338 (N_16338,N_16266,N_16238);
nand U16339 (N_16339,N_16271,N_16209);
nand U16340 (N_16340,N_16317,N_16230);
nor U16341 (N_16341,N_16165,N_16241);
or U16342 (N_16342,N_16187,N_16257);
nand U16343 (N_16343,N_16298,N_16288);
xnor U16344 (N_16344,N_16263,N_16190);
or U16345 (N_16345,N_16201,N_16181);
nand U16346 (N_16346,N_16164,N_16229);
nor U16347 (N_16347,N_16245,N_16293);
nor U16348 (N_16348,N_16269,N_16280);
or U16349 (N_16349,N_16232,N_16216);
nand U16350 (N_16350,N_16228,N_16306);
nor U16351 (N_16351,N_16248,N_16168);
xnor U16352 (N_16352,N_16218,N_16221);
nand U16353 (N_16353,N_16174,N_16299);
and U16354 (N_16354,N_16275,N_16225);
and U16355 (N_16355,N_16205,N_16309);
nor U16356 (N_16356,N_16273,N_16182);
nand U16357 (N_16357,N_16226,N_16210);
and U16358 (N_16358,N_16318,N_16163);
or U16359 (N_16359,N_16315,N_16195);
nor U16360 (N_16360,N_16192,N_16312);
nand U16361 (N_16361,N_16237,N_16202);
nor U16362 (N_16362,N_16214,N_16166);
xnor U16363 (N_16363,N_16240,N_16296);
nor U16364 (N_16364,N_16313,N_16213);
nor U16365 (N_16365,N_16256,N_16261);
nor U16366 (N_16366,N_16215,N_16204);
or U16367 (N_16367,N_16176,N_16222);
or U16368 (N_16368,N_16283,N_16246);
nand U16369 (N_16369,N_16231,N_16220);
or U16370 (N_16370,N_16291,N_16233);
or U16371 (N_16371,N_16203,N_16249);
and U16372 (N_16372,N_16276,N_16170);
and U16373 (N_16373,N_16191,N_16173);
nor U16374 (N_16374,N_16316,N_16239);
nor U16375 (N_16375,N_16279,N_16287);
and U16376 (N_16376,N_16169,N_16207);
and U16377 (N_16377,N_16211,N_16244);
or U16378 (N_16378,N_16206,N_16265);
xnor U16379 (N_16379,N_16285,N_16183);
xor U16380 (N_16380,N_16311,N_16178);
nand U16381 (N_16381,N_16304,N_16171);
nor U16382 (N_16382,N_16295,N_16167);
nor U16383 (N_16383,N_16184,N_16234);
xnor U16384 (N_16384,N_16282,N_16259);
and U16385 (N_16385,N_16242,N_16258);
or U16386 (N_16386,N_16179,N_16278);
xor U16387 (N_16387,N_16188,N_16305);
nor U16388 (N_16388,N_16264,N_16194);
xnor U16389 (N_16389,N_16180,N_16281);
or U16390 (N_16390,N_16199,N_16219);
nand U16391 (N_16391,N_16200,N_16290);
nor U16392 (N_16392,N_16193,N_16314);
xnor U16393 (N_16393,N_16185,N_16272);
nor U16394 (N_16394,N_16255,N_16250);
and U16395 (N_16395,N_16286,N_16223);
xor U16396 (N_16396,N_16262,N_16270);
xor U16397 (N_16397,N_16251,N_16307);
and U16398 (N_16398,N_16175,N_16189);
xor U16399 (N_16399,N_16162,N_16197);
and U16400 (N_16400,N_16263,N_16205);
and U16401 (N_16401,N_16292,N_16178);
nor U16402 (N_16402,N_16207,N_16200);
nand U16403 (N_16403,N_16167,N_16283);
or U16404 (N_16404,N_16273,N_16202);
nor U16405 (N_16405,N_16307,N_16184);
xor U16406 (N_16406,N_16210,N_16212);
nor U16407 (N_16407,N_16318,N_16234);
and U16408 (N_16408,N_16187,N_16176);
or U16409 (N_16409,N_16206,N_16307);
nor U16410 (N_16410,N_16162,N_16179);
or U16411 (N_16411,N_16227,N_16280);
and U16412 (N_16412,N_16313,N_16255);
or U16413 (N_16413,N_16292,N_16265);
nand U16414 (N_16414,N_16171,N_16245);
and U16415 (N_16415,N_16253,N_16281);
nand U16416 (N_16416,N_16242,N_16194);
and U16417 (N_16417,N_16273,N_16259);
and U16418 (N_16418,N_16189,N_16271);
and U16419 (N_16419,N_16255,N_16271);
nor U16420 (N_16420,N_16167,N_16231);
or U16421 (N_16421,N_16281,N_16258);
or U16422 (N_16422,N_16314,N_16161);
nor U16423 (N_16423,N_16179,N_16233);
nor U16424 (N_16424,N_16200,N_16263);
nand U16425 (N_16425,N_16261,N_16267);
nor U16426 (N_16426,N_16309,N_16287);
and U16427 (N_16427,N_16243,N_16199);
or U16428 (N_16428,N_16191,N_16246);
and U16429 (N_16429,N_16313,N_16176);
or U16430 (N_16430,N_16210,N_16215);
nor U16431 (N_16431,N_16160,N_16214);
nand U16432 (N_16432,N_16301,N_16177);
xor U16433 (N_16433,N_16199,N_16296);
xor U16434 (N_16434,N_16279,N_16261);
nand U16435 (N_16435,N_16196,N_16298);
or U16436 (N_16436,N_16316,N_16188);
nand U16437 (N_16437,N_16302,N_16311);
or U16438 (N_16438,N_16275,N_16317);
and U16439 (N_16439,N_16276,N_16232);
xor U16440 (N_16440,N_16268,N_16208);
and U16441 (N_16441,N_16184,N_16207);
nand U16442 (N_16442,N_16232,N_16307);
nand U16443 (N_16443,N_16201,N_16221);
xor U16444 (N_16444,N_16249,N_16196);
nor U16445 (N_16445,N_16214,N_16257);
nor U16446 (N_16446,N_16220,N_16223);
nor U16447 (N_16447,N_16186,N_16169);
and U16448 (N_16448,N_16268,N_16244);
or U16449 (N_16449,N_16307,N_16219);
or U16450 (N_16450,N_16166,N_16200);
or U16451 (N_16451,N_16282,N_16223);
nand U16452 (N_16452,N_16173,N_16160);
xnor U16453 (N_16453,N_16273,N_16244);
xor U16454 (N_16454,N_16287,N_16286);
nand U16455 (N_16455,N_16303,N_16162);
nor U16456 (N_16456,N_16188,N_16213);
xor U16457 (N_16457,N_16244,N_16299);
or U16458 (N_16458,N_16196,N_16214);
nor U16459 (N_16459,N_16297,N_16204);
nand U16460 (N_16460,N_16203,N_16255);
or U16461 (N_16461,N_16281,N_16207);
xor U16462 (N_16462,N_16192,N_16197);
nor U16463 (N_16463,N_16252,N_16206);
or U16464 (N_16464,N_16309,N_16211);
xnor U16465 (N_16465,N_16236,N_16284);
nand U16466 (N_16466,N_16272,N_16228);
and U16467 (N_16467,N_16167,N_16204);
nor U16468 (N_16468,N_16187,N_16301);
and U16469 (N_16469,N_16168,N_16203);
and U16470 (N_16470,N_16215,N_16257);
nand U16471 (N_16471,N_16164,N_16299);
xor U16472 (N_16472,N_16164,N_16182);
nor U16473 (N_16473,N_16160,N_16259);
or U16474 (N_16474,N_16288,N_16297);
nor U16475 (N_16475,N_16310,N_16180);
nor U16476 (N_16476,N_16281,N_16166);
xnor U16477 (N_16477,N_16270,N_16209);
xor U16478 (N_16478,N_16274,N_16284);
nor U16479 (N_16479,N_16178,N_16168);
xnor U16480 (N_16480,N_16443,N_16472);
or U16481 (N_16481,N_16459,N_16444);
xnor U16482 (N_16482,N_16479,N_16409);
and U16483 (N_16483,N_16360,N_16380);
xor U16484 (N_16484,N_16420,N_16340);
nand U16485 (N_16485,N_16473,N_16469);
and U16486 (N_16486,N_16377,N_16382);
nand U16487 (N_16487,N_16447,N_16437);
or U16488 (N_16488,N_16398,N_16334);
nand U16489 (N_16489,N_16339,N_16478);
xor U16490 (N_16490,N_16435,N_16400);
nor U16491 (N_16491,N_16425,N_16451);
nor U16492 (N_16492,N_16368,N_16337);
nor U16493 (N_16493,N_16441,N_16323);
nand U16494 (N_16494,N_16358,N_16439);
and U16495 (N_16495,N_16404,N_16357);
xnor U16496 (N_16496,N_16397,N_16324);
and U16497 (N_16497,N_16365,N_16412);
nor U16498 (N_16498,N_16448,N_16336);
nor U16499 (N_16499,N_16422,N_16374);
nor U16500 (N_16500,N_16395,N_16430);
nand U16501 (N_16501,N_16442,N_16359);
nand U16502 (N_16502,N_16390,N_16326);
or U16503 (N_16503,N_16333,N_16343);
nor U16504 (N_16504,N_16393,N_16325);
xor U16505 (N_16505,N_16463,N_16366);
nand U16506 (N_16506,N_16349,N_16468);
or U16507 (N_16507,N_16421,N_16428);
nand U16508 (N_16508,N_16351,N_16401);
nor U16509 (N_16509,N_16372,N_16406);
and U16510 (N_16510,N_16440,N_16364);
and U16511 (N_16511,N_16452,N_16474);
xor U16512 (N_16512,N_16402,N_16331);
nor U16513 (N_16513,N_16431,N_16434);
and U16514 (N_16514,N_16385,N_16354);
xor U16515 (N_16515,N_16369,N_16408);
or U16516 (N_16516,N_16477,N_16455);
xor U16517 (N_16517,N_16456,N_16384);
xor U16518 (N_16518,N_16342,N_16426);
nor U16519 (N_16519,N_16405,N_16438);
nor U16520 (N_16520,N_16328,N_16446);
or U16521 (N_16521,N_16461,N_16367);
nand U16522 (N_16522,N_16457,N_16375);
nand U16523 (N_16523,N_16429,N_16458);
nand U16524 (N_16524,N_16427,N_16373);
nor U16525 (N_16525,N_16330,N_16381);
and U16526 (N_16526,N_16403,N_16332);
xor U16527 (N_16527,N_16411,N_16376);
nand U16528 (N_16528,N_16341,N_16462);
or U16529 (N_16529,N_16361,N_16378);
nand U16530 (N_16530,N_16348,N_16416);
or U16531 (N_16531,N_16424,N_16464);
nor U16532 (N_16532,N_16394,N_16356);
nor U16533 (N_16533,N_16387,N_16350);
nor U16534 (N_16534,N_16386,N_16320);
xor U16535 (N_16535,N_16432,N_16345);
or U16536 (N_16536,N_16449,N_16322);
nand U16537 (N_16537,N_16347,N_16355);
and U16538 (N_16538,N_16414,N_16338);
nand U16539 (N_16539,N_16389,N_16392);
nand U16540 (N_16540,N_16379,N_16418);
and U16541 (N_16541,N_16417,N_16419);
nor U16542 (N_16542,N_16383,N_16470);
or U16543 (N_16543,N_16399,N_16453);
and U16544 (N_16544,N_16450,N_16466);
xnor U16545 (N_16545,N_16454,N_16388);
and U16546 (N_16546,N_16475,N_16465);
or U16547 (N_16547,N_16362,N_16467);
nor U16548 (N_16548,N_16413,N_16391);
xor U16549 (N_16549,N_16415,N_16471);
or U16550 (N_16550,N_16344,N_16329);
and U16551 (N_16551,N_16476,N_16407);
xor U16552 (N_16552,N_16371,N_16423);
nand U16553 (N_16553,N_16363,N_16410);
nor U16554 (N_16554,N_16352,N_16346);
xnor U16555 (N_16555,N_16433,N_16335);
xnor U16556 (N_16556,N_16396,N_16445);
or U16557 (N_16557,N_16321,N_16353);
nor U16558 (N_16558,N_16436,N_16370);
nand U16559 (N_16559,N_16327,N_16460);
xor U16560 (N_16560,N_16435,N_16402);
or U16561 (N_16561,N_16339,N_16439);
nand U16562 (N_16562,N_16459,N_16390);
nor U16563 (N_16563,N_16435,N_16422);
nand U16564 (N_16564,N_16453,N_16413);
and U16565 (N_16565,N_16419,N_16422);
or U16566 (N_16566,N_16401,N_16376);
and U16567 (N_16567,N_16414,N_16467);
nor U16568 (N_16568,N_16323,N_16384);
or U16569 (N_16569,N_16410,N_16453);
nand U16570 (N_16570,N_16390,N_16376);
nand U16571 (N_16571,N_16405,N_16359);
and U16572 (N_16572,N_16355,N_16396);
nand U16573 (N_16573,N_16419,N_16390);
and U16574 (N_16574,N_16377,N_16379);
nand U16575 (N_16575,N_16416,N_16432);
and U16576 (N_16576,N_16462,N_16390);
nand U16577 (N_16577,N_16412,N_16398);
nor U16578 (N_16578,N_16356,N_16370);
nand U16579 (N_16579,N_16360,N_16334);
and U16580 (N_16580,N_16378,N_16377);
nor U16581 (N_16581,N_16320,N_16390);
nand U16582 (N_16582,N_16377,N_16372);
or U16583 (N_16583,N_16388,N_16386);
nand U16584 (N_16584,N_16416,N_16436);
and U16585 (N_16585,N_16425,N_16364);
xnor U16586 (N_16586,N_16323,N_16412);
or U16587 (N_16587,N_16338,N_16396);
and U16588 (N_16588,N_16473,N_16322);
and U16589 (N_16589,N_16359,N_16408);
or U16590 (N_16590,N_16417,N_16431);
and U16591 (N_16591,N_16434,N_16385);
nand U16592 (N_16592,N_16366,N_16379);
nand U16593 (N_16593,N_16327,N_16437);
and U16594 (N_16594,N_16434,N_16337);
nand U16595 (N_16595,N_16363,N_16348);
nor U16596 (N_16596,N_16464,N_16472);
nor U16597 (N_16597,N_16368,N_16353);
or U16598 (N_16598,N_16340,N_16365);
or U16599 (N_16599,N_16389,N_16343);
and U16600 (N_16600,N_16377,N_16407);
xnor U16601 (N_16601,N_16444,N_16424);
or U16602 (N_16602,N_16391,N_16441);
or U16603 (N_16603,N_16362,N_16391);
nor U16604 (N_16604,N_16380,N_16416);
nand U16605 (N_16605,N_16331,N_16364);
nand U16606 (N_16606,N_16372,N_16441);
or U16607 (N_16607,N_16358,N_16421);
and U16608 (N_16608,N_16379,N_16451);
nand U16609 (N_16609,N_16361,N_16385);
xor U16610 (N_16610,N_16396,N_16329);
nor U16611 (N_16611,N_16328,N_16465);
or U16612 (N_16612,N_16415,N_16386);
nand U16613 (N_16613,N_16420,N_16407);
xor U16614 (N_16614,N_16427,N_16375);
or U16615 (N_16615,N_16425,N_16354);
nand U16616 (N_16616,N_16373,N_16439);
and U16617 (N_16617,N_16329,N_16359);
nor U16618 (N_16618,N_16373,N_16391);
xnor U16619 (N_16619,N_16348,N_16423);
or U16620 (N_16620,N_16391,N_16460);
xor U16621 (N_16621,N_16476,N_16345);
nor U16622 (N_16622,N_16441,N_16385);
and U16623 (N_16623,N_16429,N_16460);
and U16624 (N_16624,N_16372,N_16447);
and U16625 (N_16625,N_16387,N_16343);
nand U16626 (N_16626,N_16373,N_16364);
xor U16627 (N_16627,N_16414,N_16371);
nor U16628 (N_16628,N_16322,N_16329);
nor U16629 (N_16629,N_16473,N_16432);
and U16630 (N_16630,N_16464,N_16383);
nand U16631 (N_16631,N_16426,N_16448);
or U16632 (N_16632,N_16464,N_16368);
and U16633 (N_16633,N_16452,N_16428);
or U16634 (N_16634,N_16330,N_16326);
and U16635 (N_16635,N_16410,N_16446);
and U16636 (N_16636,N_16465,N_16385);
nand U16637 (N_16637,N_16352,N_16475);
and U16638 (N_16638,N_16396,N_16326);
or U16639 (N_16639,N_16336,N_16412);
and U16640 (N_16640,N_16527,N_16602);
xnor U16641 (N_16641,N_16600,N_16607);
xnor U16642 (N_16642,N_16503,N_16487);
or U16643 (N_16643,N_16614,N_16629);
nor U16644 (N_16644,N_16604,N_16628);
and U16645 (N_16645,N_16554,N_16575);
or U16646 (N_16646,N_16597,N_16561);
xor U16647 (N_16647,N_16612,N_16516);
or U16648 (N_16648,N_16519,N_16549);
or U16649 (N_16649,N_16528,N_16506);
xor U16650 (N_16650,N_16522,N_16583);
xor U16651 (N_16651,N_16489,N_16539);
or U16652 (N_16652,N_16546,N_16529);
xnor U16653 (N_16653,N_16523,N_16552);
and U16654 (N_16654,N_16496,N_16557);
nor U16655 (N_16655,N_16494,N_16555);
or U16656 (N_16656,N_16637,N_16615);
and U16657 (N_16657,N_16515,N_16536);
xnor U16658 (N_16658,N_16572,N_16638);
nor U16659 (N_16659,N_16488,N_16626);
xor U16660 (N_16660,N_16521,N_16556);
or U16661 (N_16661,N_16576,N_16590);
nor U16662 (N_16662,N_16617,N_16574);
and U16663 (N_16663,N_16564,N_16611);
or U16664 (N_16664,N_16510,N_16573);
or U16665 (N_16665,N_16484,N_16543);
nand U16666 (N_16666,N_16622,N_16482);
xnor U16667 (N_16667,N_16565,N_16524);
xnor U16668 (N_16668,N_16605,N_16623);
nor U16669 (N_16669,N_16501,N_16505);
xor U16670 (N_16670,N_16558,N_16625);
nand U16671 (N_16671,N_16571,N_16548);
xnor U16672 (N_16672,N_16589,N_16497);
nor U16673 (N_16673,N_16577,N_16485);
nor U16674 (N_16674,N_16551,N_16631);
or U16675 (N_16675,N_16586,N_16594);
nor U16676 (N_16676,N_16578,N_16582);
nor U16677 (N_16677,N_16636,N_16535);
or U16678 (N_16678,N_16635,N_16483);
or U16679 (N_16679,N_16639,N_16609);
nand U16680 (N_16680,N_16504,N_16585);
and U16681 (N_16681,N_16533,N_16620);
xor U16682 (N_16682,N_16587,N_16512);
and U16683 (N_16683,N_16567,N_16495);
and U16684 (N_16684,N_16526,N_16619);
xor U16685 (N_16685,N_16584,N_16624);
and U16686 (N_16686,N_16570,N_16520);
xnor U16687 (N_16687,N_16599,N_16540);
xnor U16688 (N_16688,N_16525,N_16490);
xor U16689 (N_16689,N_16492,N_16616);
nand U16690 (N_16690,N_16544,N_16507);
or U16691 (N_16691,N_16591,N_16566);
xor U16692 (N_16692,N_16610,N_16502);
xnor U16693 (N_16693,N_16499,N_16630);
nand U16694 (N_16694,N_16598,N_16480);
xnor U16695 (N_16695,N_16559,N_16518);
and U16696 (N_16696,N_16531,N_16627);
nand U16697 (N_16697,N_16592,N_16634);
nor U16698 (N_16698,N_16509,N_16508);
and U16699 (N_16699,N_16517,N_16606);
xnor U16700 (N_16700,N_16481,N_16545);
nor U16701 (N_16701,N_16538,N_16530);
and U16702 (N_16702,N_16560,N_16493);
and U16703 (N_16703,N_16532,N_16542);
nor U16704 (N_16704,N_16593,N_16581);
nor U16705 (N_16705,N_16621,N_16613);
and U16706 (N_16706,N_16500,N_16541);
and U16707 (N_16707,N_16534,N_16580);
xnor U16708 (N_16708,N_16513,N_16514);
and U16709 (N_16709,N_16511,N_16498);
or U16710 (N_16710,N_16537,N_16562);
nor U16711 (N_16711,N_16569,N_16633);
nor U16712 (N_16712,N_16596,N_16491);
nand U16713 (N_16713,N_16550,N_16603);
xor U16714 (N_16714,N_16486,N_16595);
and U16715 (N_16715,N_16618,N_16588);
nand U16716 (N_16716,N_16632,N_16568);
or U16717 (N_16717,N_16579,N_16563);
and U16718 (N_16718,N_16601,N_16547);
xnor U16719 (N_16719,N_16553,N_16608);
or U16720 (N_16720,N_16560,N_16526);
nor U16721 (N_16721,N_16556,N_16607);
xnor U16722 (N_16722,N_16502,N_16568);
xor U16723 (N_16723,N_16502,N_16607);
or U16724 (N_16724,N_16603,N_16487);
and U16725 (N_16725,N_16609,N_16572);
and U16726 (N_16726,N_16620,N_16584);
nor U16727 (N_16727,N_16484,N_16577);
nand U16728 (N_16728,N_16609,N_16502);
nor U16729 (N_16729,N_16490,N_16624);
and U16730 (N_16730,N_16586,N_16507);
or U16731 (N_16731,N_16586,N_16532);
nand U16732 (N_16732,N_16613,N_16513);
nor U16733 (N_16733,N_16540,N_16556);
or U16734 (N_16734,N_16609,N_16543);
nor U16735 (N_16735,N_16543,N_16589);
or U16736 (N_16736,N_16608,N_16610);
xor U16737 (N_16737,N_16485,N_16582);
and U16738 (N_16738,N_16549,N_16584);
nor U16739 (N_16739,N_16527,N_16564);
nand U16740 (N_16740,N_16487,N_16515);
nor U16741 (N_16741,N_16554,N_16627);
and U16742 (N_16742,N_16532,N_16541);
xnor U16743 (N_16743,N_16538,N_16491);
or U16744 (N_16744,N_16560,N_16481);
nor U16745 (N_16745,N_16593,N_16586);
nor U16746 (N_16746,N_16500,N_16597);
and U16747 (N_16747,N_16495,N_16629);
nor U16748 (N_16748,N_16546,N_16548);
and U16749 (N_16749,N_16600,N_16565);
and U16750 (N_16750,N_16513,N_16633);
and U16751 (N_16751,N_16501,N_16607);
nand U16752 (N_16752,N_16578,N_16619);
nand U16753 (N_16753,N_16508,N_16634);
and U16754 (N_16754,N_16633,N_16508);
nand U16755 (N_16755,N_16632,N_16531);
and U16756 (N_16756,N_16500,N_16617);
nor U16757 (N_16757,N_16606,N_16612);
and U16758 (N_16758,N_16484,N_16609);
nand U16759 (N_16759,N_16585,N_16545);
nor U16760 (N_16760,N_16524,N_16615);
and U16761 (N_16761,N_16626,N_16519);
and U16762 (N_16762,N_16508,N_16601);
xnor U16763 (N_16763,N_16632,N_16544);
nand U16764 (N_16764,N_16490,N_16530);
and U16765 (N_16765,N_16557,N_16598);
xor U16766 (N_16766,N_16491,N_16638);
nand U16767 (N_16767,N_16519,N_16571);
or U16768 (N_16768,N_16543,N_16494);
or U16769 (N_16769,N_16504,N_16505);
nand U16770 (N_16770,N_16594,N_16514);
nor U16771 (N_16771,N_16614,N_16506);
xnor U16772 (N_16772,N_16581,N_16515);
or U16773 (N_16773,N_16556,N_16638);
nor U16774 (N_16774,N_16603,N_16579);
or U16775 (N_16775,N_16519,N_16512);
nor U16776 (N_16776,N_16572,N_16600);
or U16777 (N_16777,N_16559,N_16527);
nand U16778 (N_16778,N_16486,N_16628);
and U16779 (N_16779,N_16531,N_16511);
nand U16780 (N_16780,N_16587,N_16624);
nor U16781 (N_16781,N_16613,N_16629);
nor U16782 (N_16782,N_16557,N_16596);
xor U16783 (N_16783,N_16627,N_16534);
and U16784 (N_16784,N_16483,N_16533);
nand U16785 (N_16785,N_16549,N_16510);
nor U16786 (N_16786,N_16536,N_16617);
nand U16787 (N_16787,N_16522,N_16528);
or U16788 (N_16788,N_16526,N_16487);
or U16789 (N_16789,N_16553,N_16572);
and U16790 (N_16790,N_16484,N_16600);
nor U16791 (N_16791,N_16483,N_16531);
xor U16792 (N_16792,N_16561,N_16538);
and U16793 (N_16793,N_16630,N_16512);
or U16794 (N_16794,N_16562,N_16630);
and U16795 (N_16795,N_16507,N_16496);
or U16796 (N_16796,N_16588,N_16634);
nor U16797 (N_16797,N_16544,N_16545);
xnor U16798 (N_16798,N_16537,N_16543);
nor U16799 (N_16799,N_16594,N_16607);
nor U16800 (N_16800,N_16776,N_16764);
nor U16801 (N_16801,N_16741,N_16758);
xnor U16802 (N_16802,N_16690,N_16733);
xnor U16803 (N_16803,N_16675,N_16688);
and U16804 (N_16804,N_16752,N_16661);
nand U16805 (N_16805,N_16712,N_16766);
and U16806 (N_16806,N_16701,N_16677);
nor U16807 (N_16807,N_16706,N_16761);
or U16808 (N_16808,N_16647,N_16643);
nor U16809 (N_16809,N_16757,N_16660);
or U16810 (N_16810,N_16739,N_16659);
xor U16811 (N_16811,N_16645,N_16650);
nor U16812 (N_16812,N_16704,N_16685);
or U16813 (N_16813,N_16779,N_16744);
xor U16814 (N_16814,N_16674,N_16782);
and U16815 (N_16815,N_16730,N_16737);
nor U16816 (N_16816,N_16783,N_16743);
and U16817 (N_16817,N_16662,N_16792);
and U16818 (N_16818,N_16790,N_16716);
nor U16819 (N_16819,N_16795,N_16679);
or U16820 (N_16820,N_16691,N_16784);
nor U16821 (N_16821,N_16732,N_16667);
xor U16822 (N_16822,N_16793,N_16794);
or U16823 (N_16823,N_16759,N_16749);
xnor U16824 (N_16824,N_16665,N_16699);
nand U16825 (N_16825,N_16702,N_16683);
xnor U16826 (N_16826,N_16756,N_16654);
or U16827 (N_16827,N_16709,N_16686);
and U16828 (N_16828,N_16687,N_16676);
nor U16829 (N_16829,N_16781,N_16641);
nor U16830 (N_16830,N_16652,N_16651);
or U16831 (N_16831,N_16672,N_16720);
or U16832 (N_16832,N_16736,N_16775);
nor U16833 (N_16833,N_16678,N_16788);
nand U16834 (N_16834,N_16696,N_16689);
xor U16835 (N_16835,N_16768,N_16767);
nor U16836 (N_16836,N_16723,N_16668);
or U16837 (N_16837,N_16727,N_16791);
xnor U16838 (N_16838,N_16703,N_16785);
xor U16839 (N_16839,N_16762,N_16642);
nor U16840 (N_16840,N_16695,N_16664);
nand U16841 (N_16841,N_16656,N_16708);
or U16842 (N_16842,N_16657,N_16692);
nor U16843 (N_16843,N_16765,N_16771);
or U16844 (N_16844,N_16681,N_16682);
and U16845 (N_16845,N_16747,N_16799);
nand U16846 (N_16846,N_16669,N_16658);
xnor U16847 (N_16847,N_16787,N_16714);
nor U16848 (N_16848,N_16705,N_16748);
and U16849 (N_16849,N_16746,N_16725);
and U16850 (N_16850,N_16763,N_16713);
nand U16851 (N_16851,N_16755,N_16773);
xnor U16852 (N_16852,N_16640,N_16666);
or U16853 (N_16853,N_16789,N_16649);
nand U16854 (N_16854,N_16726,N_16718);
nor U16855 (N_16855,N_16710,N_16769);
xnor U16856 (N_16856,N_16778,N_16796);
nor U16857 (N_16857,N_16700,N_16694);
xnor U16858 (N_16858,N_16719,N_16697);
nand U16859 (N_16859,N_16728,N_16644);
nor U16860 (N_16860,N_16724,N_16715);
and U16861 (N_16861,N_16731,N_16738);
nand U16862 (N_16862,N_16671,N_16751);
nand U16863 (N_16863,N_16774,N_16680);
xor U16864 (N_16864,N_16707,N_16722);
or U16865 (N_16865,N_16777,N_16760);
and U16866 (N_16866,N_16684,N_16655);
nor U16867 (N_16867,N_16693,N_16721);
nand U16868 (N_16868,N_16698,N_16745);
nand U16869 (N_16869,N_16753,N_16797);
and U16870 (N_16870,N_16754,N_16670);
nand U16871 (N_16871,N_16772,N_16742);
nand U16872 (N_16872,N_16663,N_16750);
xor U16873 (N_16873,N_16770,N_16653);
xnor U16874 (N_16874,N_16711,N_16780);
nand U16875 (N_16875,N_16734,N_16646);
xor U16876 (N_16876,N_16798,N_16735);
or U16877 (N_16877,N_16729,N_16740);
and U16878 (N_16878,N_16648,N_16673);
nand U16879 (N_16879,N_16717,N_16786);
and U16880 (N_16880,N_16687,N_16640);
or U16881 (N_16881,N_16771,N_16704);
nor U16882 (N_16882,N_16780,N_16787);
or U16883 (N_16883,N_16653,N_16677);
nand U16884 (N_16884,N_16693,N_16640);
and U16885 (N_16885,N_16716,N_16733);
nand U16886 (N_16886,N_16767,N_16723);
nor U16887 (N_16887,N_16749,N_16652);
and U16888 (N_16888,N_16646,N_16730);
nand U16889 (N_16889,N_16733,N_16735);
or U16890 (N_16890,N_16641,N_16724);
and U16891 (N_16891,N_16708,N_16660);
or U16892 (N_16892,N_16684,N_16781);
nor U16893 (N_16893,N_16761,N_16783);
xor U16894 (N_16894,N_16783,N_16690);
nor U16895 (N_16895,N_16688,N_16703);
xor U16896 (N_16896,N_16687,N_16644);
nand U16897 (N_16897,N_16670,N_16732);
or U16898 (N_16898,N_16647,N_16644);
or U16899 (N_16899,N_16769,N_16799);
nand U16900 (N_16900,N_16789,N_16670);
or U16901 (N_16901,N_16645,N_16689);
nor U16902 (N_16902,N_16645,N_16794);
or U16903 (N_16903,N_16741,N_16799);
nor U16904 (N_16904,N_16675,N_16658);
nand U16905 (N_16905,N_16656,N_16780);
or U16906 (N_16906,N_16681,N_16747);
nor U16907 (N_16907,N_16786,N_16726);
xnor U16908 (N_16908,N_16757,N_16762);
xnor U16909 (N_16909,N_16750,N_16690);
xor U16910 (N_16910,N_16745,N_16774);
xor U16911 (N_16911,N_16747,N_16648);
nand U16912 (N_16912,N_16770,N_16795);
nor U16913 (N_16913,N_16754,N_16663);
and U16914 (N_16914,N_16717,N_16785);
nor U16915 (N_16915,N_16771,N_16732);
nand U16916 (N_16916,N_16730,N_16685);
or U16917 (N_16917,N_16722,N_16781);
nor U16918 (N_16918,N_16737,N_16777);
or U16919 (N_16919,N_16780,N_16714);
nand U16920 (N_16920,N_16666,N_16661);
nor U16921 (N_16921,N_16796,N_16691);
nand U16922 (N_16922,N_16710,N_16709);
nor U16923 (N_16923,N_16756,N_16741);
or U16924 (N_16924,N_16733,N_16678);
nand U16925 (N_16925,N_16744,N_16795);
nand U16926 (N_16926,N_16742,N_16788);
nand U16927 (N_16927,N_16642,N_16682);
nor U16928 (N_16928,N_16657,N_16736);
nand U16929 (N_16929,N_16763,N_16725);
nor U16930 (N_16930,N_16784,N_16727);
or U16931 (N_16931,N_16686,N_16716);
xnor U16932 (N_16932,N_16680,N_16742);
nor U16933 (N_16933,N_16728,N_16753);
and U16934 (N_16934,N_16773,N_16709);
or U16935 (N_16935,N_16725,N_16673);
and U16936 (N_16936,N_16659,N_16693);
and U16937 (N_16937,N_16711,N_16768);
nor U16938 (N_16938,N_16744,N_16681);
xnor U16939 (N_16939,N_16794,N_16729);
xor U16940 (N_16940,N_16780,N_16778);
xor U16941 (N_16941,N_16725,N_16677);
nand U16942 (N_16942,N_16727,N_16699);
xor U16943 (N_16943,N_16709,N_16790);
nor U16944 (N_16944,N_16790,N_16771);
or U16945 (N_16945,N_16696,N_16737);
xnor U16946 (N_16946,N_16741,N_16748);
and U16947 (N_16947,N_16748,N_16683);
nor U16948 (N_16948,N_16747,N_16783);
nand U16949 (N_16949,N_16662,N_16746);
nand U16950 (N_16950,N_16768,N_16728);
or U16951 (N_16951,N_16706,N_16795);
xnor U16952 (N_16952,N_16663,N_16702);
nand U16953 (N_16953,N_16790,N_16789);
and U16954 (N_16954,N_16689,N_16772);
nand U16955 (N_16955,N_16746,N_16696);
nor U16956 (N_16956,N_16763,N_16792);
xnor U16957 (N_16957,N_16789,N_16669);
nor U16958 (N_16958,N_16737,N_16784);
nand U16959 (N_16959,N_16702,N_16707);
or U16960 (N_16960,N_16952,N_16843);
nand U16961 (N_16961,N_16829,N_16947);
or U16962 (N_16962,N_16845,N_16892);
nand U16963 (N_16963,N_16921,N_16899);
nor U16964 (N_16964,N_16854,N_16871);
or U16965 (N_16965,N_16890,N_16933);
xor U16966 (N_16966,N_16918,N_16864);
nor U16967 (N_16967,N_16954,N_16810);
xnor U16968 (N_16968,N_16886,N_16814);
and U16969 (N_16969,N_16941,N_16876);
nor U16970 (N_16970,N_16832,N_16959);
nand U16971 (N_16971,N_16862,N_16953);
or U16972 (N_16972,N_16855,N_16881);
nand U16973 (N_16973,N_16821,N_16875);
or U16974 (N_16974,N_16866,N_16804);
or U16975 (N_16975,N_16884,N_16882);
xor U16976 (N_16976,N_16906,N_16955);
or U16977 (N_16977,N_16831,N_16874);
xor U16978 (N_16978,N_16951,N_16860);
nand U16979 (N_16979,N_16885,N_16840);
or U16980 (N_16980,N_16809,N_16895);
and U16981 (N_16981,N_16807,N_16908);
nand U16982 (N_16982,N_16861,N_16870);
and U16983 (N_16983,N_16846,N_16856);
nand U16984 (N_16984,N_16904,N_16894);
and U16985 (N_16985,N_16813,N_16911);
or U16986 (N_16986,N_16903,N_16834);
or U16987 (N_16987,N_16868,N_16900);
nand U16988 (N_16988,N_16931,N_16818);
nand U16989 (N_16989,N_16896,N_16839);
nand U16990 (N_16990,N_16841,N_16905);
nor U16991 (N_16991,N_16945,N_16880);
and U16992 (N_16992,N_16938,N_16842);
xnor U16993 (N_16993,N_16825,N_16838);
or U16994 (N_16994,N_16949,N_16927);
or U16995 (N_16995,N_16836,N_16936);
nor U16996 (N_16996,N_16958,N_16847);
xor U16997 (N_16997,N_16805,N_16926);
nand U16998 (N_16998,N_16826,N_16893);
nand U16999 (N_16999,N_16942,N_16922);
nand U17000 (N_17000,N_16910,N_16873);
nand U17001 (N_17001,N_16935,N_16923);
xor U17002 (N_17002,N_16928,N_16956);
xor U17003 (N_17003,N_16808,N_16848);
or U17004 (N_17004,N_16858,N_16909);
or U17005 (N_17005,N_16857,N_16828);
nor U17006 (N_17006,N_16901,N_16929);
and U17007 (N_17007,N_16943,N_16849);
and U17008 (N_17008,N_16816,N_16819);
xor U17009 (N_17009,N_16853,N_16865);
or U17010 (N_17010,N_16907,N_16850);
xor U17011 (N_17011,N_16859,N_16925);
and U17012 (N_17012,N_16917,N_16806);
and U17013 (N_17013,N_16802,N_16869);
nor U17014 (N_17014,N_16878,N_16888);
nand U17015 (N_17015,N_16817,N_16891);
nand U17016 (N_17016,N_16950,N_16932);
or U17017 (N_17017,N_16851,N_16914);
nand U17018 (N_17018,N_16822,N_16930);
nand U17019 (N_17019,N_16827,N_16897);
nand U17020 (N_17020,N_16902,N_16934);
nand U17021 (N_17021,N_16820,N_16872);
nand U17022 (N_17022,N_16913,N_16944);
or U17023 (N_17023,N_16948,N_16957);
xor U17024 (N_17024,N_16812,N_16815);
nor U17025 (N_17025,N_16801,N_16889);
nand U17026 (N_17026,N_16887,N_16883);
nor U17027 (N_17027,N_16837,N_16939);
and U17028 (N_17028,N_16811,N_16916);
and U17029 (N_17029,N_16920,N_16833);
or U17030 (N_17030,N_16919,N_16912);
and U17031 (N_17031,N_16877,N_16937);
nand U17032 (N_17032,N_16924,N_16867);
nor U17033 (N_17033,N_16863,N_16835);
nor U17034 (N_17034,N_16946,N_16915);
or U17035 (N_17035,N_16830,N_16823);
nor U17036 (N_17036,N_16824,N_16879);
or U17037 (N_17037,N_16898,N_16852);
nor U17038 (N_17038,N_16803,N_16844);
or U17039 (N_17039,N_16940,N_16800);
nor U17040 (N_17040,N_16919,N_16946);
and U17041 (N_17041,N_16859,N_16866);
and U17042 (N_17042,N_16847,N_16859);
or U17043 (N_17043,N_16890,N_16905);
or U17044 (N_17044,N_16857,N_16944);
nor U17045 (N_17045,N_16953,N_16898);
xnor U17046 (N_17046,N_16946,N_16825);
nor U17047 (N_17047,N_16938,N_16928);
nor U17048 (N_17048,N_16931,N_16867);
xnor U17049 (N_17049,N_16871,N_16902);
and U17050 (N_17050,N_16827,N_16919);
and U17051 (N_17051,N_16831,N_16929);
or U17052 (N_17052,N_16802,N_16906);
xor U17053 (N_17053,N_16909,N_16916);
nor U17054 (N_17054,N_16910,N_16801);
nand U17055 (N_17055,N_16885,N_16925);
and U17056 (N_17056,N_16953,N_16802);
or U17057 (N_17057,N_16815,N_16890);
and U17058 (N_17058,N_16921,N_16841);
nand U17059 (N_17059,N_16930,N_16917);
nor U17060 (N_17060,N_16933,N_16913);
and U17061 (N_17061,N_16889,N_16880);
and U17062 (N_17062,N_16832,N_16916);
nand U17063 (N_17063,N_16863,N_16802);
and U17064 (N_17064,N_16849,N_16858);
nand U17065 (N_17065,N_16904,N_16877);
nor U17066 (N_17066,N_16866,N_16910);
xnor U17067 (N_17067,N_16800,N_16811);
nand U17068 (N_17068,N_16840,N_16936);
nor U17069 (N_17069,N_16906,N_16858);
and U17070 (N_17070,N_16874,N_16830);
nand U17071 (N_17071,N_16881,N_16874);
nand U17072 (N_17072,N_16809,N_16840);
or U17073 (N_17073,N_16929,N_16824);
nor U17074 (N_17074,N_16957,N_16841);
nand U17075 (N_17075,N_16896,N_16868);
nor U17076 (N_17076,N_16805,N_16942);
and U17077 (N_17077,N_16949,N_16950);
xnor U17078 (N_17078,N_16850,N_16882);
nor U17079 (N_17079,N_16831,N_16881);
xnor U17080 (N_17080,N_16910,N_16807);
nor U17081 (N_17081,N_16844,N_16851);
nor U17082 (N_17082,N_16947,N_16938);
or U17083 (N_17083,N_16832,N_16889);
and U17084 (N_17084,N_16925,N_16872);
and U17085 (N_17085,N_16926,N_16882);
or U17086 (N_17086,N_16833,N_16900);
nand U17087 (N_17087,N_16833,N_16881);
or U17088 (N_17088,N_16934,N_16922);
nor U17089 (N_17089,N_16939,N_16880);
nand U17090 (N_17090,N_16885,N_16893);
nor U17091 (N_17091,N_16888,N_16808);
and U17092 (N_17092,N_16862,N_16849);
and U17093 (N_17093,N_16921,N_16829);
nor U17094 (N_17094,N_16837,N_16833);
and U17095 (N_17095,N_16920,N_16835);
xor U17096 (N_17096,N_16873,N_16835);
xnor U17097 (N_17097,N_16808,N_16861);
and U17098 (N_17098,N_16820,N_16800);
nor U17099 (N_17099,N_16886,N_16898);
and U17100 (N_17100,N_16821,N_16920);
or U17101 (N_17101,N_16956,N_16823);
nand U17102 (N_17102,N_16819,N_16859);
or U17103 (N_17103,N_16914,N_16811);
and U17104 (N_17104,N_16947,N_16845);
or U17105 (N_17105,N_16849,N_16802);
nand U17106 (N_17106,N_16860,N_16837);
nor U17107 (N_17107,N_16932,N_16917);
nand U17108 (N_17108,N_16901,N_16838);
or U17109 (N_17109,N_16896,N_16809);
nand U17110 (N_17110,N_16931,N_16925);
xor U17111 (N_17111,N_16832,N_16933);
nand U17112 (N_17112,N_16854,N_16945);
and U17113 (N_17113,N_16955,N_16956);
and U17114 (N_17114,N_16935,N_16949);
nor U17115 (N_17115,N_16823,N_16808);
xnor U17116 (N_17116,N_16924,N_16862);
nand U17117 (N_17117,N_16923,N_16949);
nor U17118 (N_17118,N_16914,N_16801);
and U17119 (N_17119,N_16818,N_16857);
xnor U17120 (N_17120,N_16968,N_17097);
xnor U17121 (N_17121,N_17094,N_17105);
xor U17122 (N_17122,N_17013,N_17052);
xor U17123 (N_17123,N_17075,N_17107);
nand U17124 (N_17124,N_16961,N_17028);
and U17125 (N_17125,N_17071,N_17036);
and U17126 (N_17126,N_17017,N_17106);
nand U17127 (N_17127,N_17108,N_17043);
xnor U17128 (N_17128,N_17099,N_17021);
xnor U17129 (N_17129,N_17114,N_17096);
nand U17130 (N_17130,N_16964,N_17027);
xnor U17131 (N_17131,N_16993,N_16992);
nand U17132 (N_17132,N_17022,N_17115);
nand U17133 (N_17133,N_17041,N_17024);
nor U17134 (N_17134,N_16988,N_17002);
xor U17135 (N_17135,N_17032,N_17104);
nor U17136 (N_17136,N_16975,N_17009);
or U17137 (N_17137,N_17100,N_17039);
nor U17138 (N_17138,N_16970,N_16978);
and U17139 (N_17139,N_17078,N_17083);
nor U17140 (N_17140,N_17018,N_17045);
nand U17141 (N_17141,N_17056,N_17088);
and U17142 (N_17142,N_17110,N_17058);
nand U17143 (N_17143,N_17068,N_17109);
nand U17144 (N_17144,N_16983,N_17029);
nor U17145 (N_17145,N_16963,N_17080);
nand U17146 (N_17146,N_16982,N_16994);
xnor U17147 (N_17147,N_17062,N_17025);
nand U17148 (N_17148,N_16965,N_17069);
nor U17149 (N_17149,N_17067,N_17098);
or U17150 (N_17150,N_17117,N_17015);
nand U17151 (N_17151,N_17046,N_16973);
or U17152 (N_17152,N_17000,N_17079);
or U17153 (N_17153,N_17003,N_16987);
and U17154 (N_17154,N_17035,N_17042);
xnor U17155 (N_17155,N_16986,N_17070);
xor U17156 (N_17156,N_16984,N_17005);
xnor U17157 (N_17157,N_17060,N_17044);
or U17158 (N_17158,N_17040,N_17061);
nor U17159 (N_17159,N_17037,N_17074);
nand U17160 (N_17160,N_17093,N_16995);
nor U17161 (N_17161,N_17053,N_17087);
or U17162 (N_17162,N_17014,N_17048);
or U17163 (N_17163,N_16962,N_16967);
and U17164 (N_17164,N_17111,N_17103);
and U17165 (N_17165,N_17102,N_16969);
nor U17166 (N_17166,N_17008,N_17020);
xor U17167 (N_17167,N_16991,N_17006);
and U17168 (N_17168,N_16976,N_17030);
and U17169 (N_17169,N_16977,N_17063);
xor U17170 (N_17170,N_17101,N_17084);
and U17171 (N_17171,N_17047,N_17086);
nand U17172 (N_17172,N_17089,N_17116);
or U17173 (N_17173,N_17010,N_16985);
xor U17174 (N_17174,N_17072,N_17112);
and U17175 (N_17175,N_17034,N_17085);
nor U17176 (N_17176,N_17055,N_17031);
nor U17177 (N_17177,N_17065,N_17011);
or U17178 (N_17178,N_17050,N_16960);
or U17179 (N_17179,N_17057,N_17090);
xnor U17180 (N_17180,N_16972,N_16990);
nand U17181 (N_17181,N_17019,N_17081);
or U17182 (N_17182,N_17091,N_17049);
nor U17183 (N_17183,N_16980,N_16998);
or U17184 (N_17184,N_17016,N_16981);
and U17185 (N_17185,N_17095,N_16966);
nor U17186 (N_17186,N_17023,N_16974);
nand U17187 (N_17187,N_17119,N_17004);
nand U17188 (N_17188,N_17076,N_17001);
or U17189 (N_17189,N_17026,N_16999);
and U17190 (N_17190,N_17082,N_17059);
nand U17191 (N_17191,N_17033,N_17064);
and U17192 (N_17192,N_17077,N_17054);
nor U17193 (N_17193,N_16979,N_17113);
nor U17194 (N_17194,N_17007,N_16989);
and U17195 (N_17195,N_17066,N_17038);
nor U17196 (N_17196,N_16997,N_16971);
or U17197 (N_17197,N_17092,N_16996);
xor U17198 (N_17198,N_17073,N_17012);
or U17199 (N_17199,N_17118,N_17051);
or U17200 (N_17200,N_16986,N_17006);
nand U17201 (N_17201,N_17111,N_16995);
xor U17202 (N_17202,N_17097,N_17062);
and U17203 (N_17203,N_17003,N_17078);
and U17204 (N_17204,N_17108,N_17076);
xnor U17205 (N_17205,N_17007,N_17119);
xnor U17206 (N_17206,N_17049,N_16974);
or U17207 (N_17207,N_17037,N_17061);
and U17208 (N_17208,N_17012,N_17026);
nor U17209 (N_17209,N_17009,N_17085);
nand U17210 (N_17210,N_17045,N_17055);
and U17211 (N_17211,N_17087,N_16970);
nor U17212 (N_17212,N_17008,N_17023);
or U17213 (N_17213,N_17047,N_17081);
xnor U17214 (N_17214,N_17049,N_17110);
nor U17215 (N_17215,N_17059,N_16995);
or U17216 (N_17216,N_17116,N_17100);
xor U17217 (N_17217,N_17021,N_17066);
nand U17218 (N_17218,N_17112,N_17073);
xor U17219 (N_17219,N_16993,N_17024);
nand U17220 (N_17220,N_16997,N_16985);
and U17221 (N_17221,N_16985,N_16964);
and U17222 (N_17222,N_16990,N_16974);
nand U17223 (N_17223,N_17039,N_17084);
or U17224 (N_17224,N_17025,N_17049);
nor U17225 (N_17225,N_17013,N_17039);
nand U17226 (N_17226,N_16993,N_17105);
xnor U17227 (N_17227,N_17054,N_16997);
or U17228 (N_17228,N_17029,N_17056);
and U17229 (N_17229,N_17101,N_17018);
xnor U17230 (N_17230,N_17026,N_17081);
nor U17231 (N_17231,N_16973,N_16966);
nand U17232 (N_17232,N_17046,N_17014);
or U17233 (N_17233,N_17091,N_17080);
nor U17234 (N_17234,N_16986,N_16975);
and U17235 (N_17235,N_16960,N_16995);
nand U17236 (N_17236,N_16994,N_17031);
and U17237 (N_17237,N_17049,N_16980);
or U17238 (N_17238,N_17116,N_17092);
or U17239 (N_17239,N_17017,N_17104);
and U17240 (N_17240,N_17030,N_17110);
nor U17241 (N_17241,N_17000,N_16978);
nor U17242 (N_17242,N_17023,N_17016);
nand U17243 (N_17243,N_16993,N_17078);
or U17244 (N_17244,N_17071,N_17027);
and U17245 (N_17245,N_17080,N_17110);
nor U17246 (N_17246,N_16960,N_17032);
or U17247 (N_17247,N_17113,N_17086);
xnor U17248 (N_17248,N_17002,N_17073);
nor U17249 (N_17249,N_16960,N_17036);
nor U17250 (N_17250,N_17092,N_16999);
or U17251 (N_17251,N_17003,N_17007);
xor U17252 (N_17252,N_17113,N_17022);
nor U17253 (N_17253,N_17073,N_17078);
xor U17254 (N_17254,N_17068,N_17115);
nor U17255 (N_17255,N_17005,N_17020);
nor U17256 (N_17256,N_17030,N_17096);
nand U17257 (N_17257,N_17053,N_17056);
and U17258 (N_17258,N_17038,N_17079);
xor U17259 (N_17259,N_17041,N_17087);
and U17260 (N_17260,N_16981,N_17043);
nand U17261 (N_17261,N_17112,N_16963);
and U17262 (N_17262,N_17004,N_16974);
or U17263 (N_17263,N_17048,N_17026);
or U17264 (N_17264,N_16970,N_17101);
or U17265 (N_17265,N_17061,N_17046);
and U17266 (N_17266,N_16972,N_17080);
xnor U17267 (N_17267,N_17030,N_17070);
and U17268 (N_17268,N_17116,N_16971);
and U17269 (N_17269,N_16975,N_17041);
nor U17270 (N_17270,N_17085,N_17001);
xnor U17271 (N_17271,N_17037,N_16970);
nand U17272 (N_17272,N_17074,N_17011);
nand U17273 (N_17273,N_17093,N_17076);
nand U17274 (N_17274,N_17024,N_16972);
nand U17275 (N_17275,N_17105,N_16979);
nand U17276 (N_17276,N_17098,N_16997);
nand U17277 (N_17277,N_17093,N_16992);
nor U17278 (N_17278,N_16986,N_17098);
and U17279 (N_17279,N_17081,N_16982);
or U17280 (N_17280,N_17160,N_17260);
nand U17281 (N_17281,N_17183,N_17156);
nand U17282 (N_17282,N_17210,N_17240);
nor U17283 (N_17283,N_17179,N_17182);
nand U17284 (N_17284,N_17237,N_17174);
xnor U17285 (N_17285,N_17132,N_17241);
nand U17286 (N_17286,N_17184,N_17226);
xnor U17287 (N_17287,N_17259,N_17139);
nand U17288 (N_17288,N_17264,N_17242);
or U17289 (N_17289,N_17131,N_17176);
and U17290 (N_17290,N_17196,N_17246);
or U17291 (N_17291,N_17125,N_17239);
and U17292 (N_17292,N_17233,N_17276);
nand U17293 (N_17293,N_17224,N_17231);
xor U17294 (N_17294,N_17140,N_17249);
nor U17295 (N_17295,N_17218,N_17245);
xnor U17296 (N_17296,N_17123,N_17178);
nand U17297 (N_17297,N_17258,N_17262);
and U17298 (N_17298,N_17159,N_17238);
nand U17299 (N_17299,N_17151,N_17212);
nor U17300 (N_17300,N_17211,N_17275);
xor U17301 (N_17301,N_17200,N_17173);
or U17302 (N_17302,N_17177,N_17213);
and U17303 (N_17303,N_17235,N_17143);
and U17304 (N_17304,N_17251,N_17198);
nand U17305 (N_17305,N_17169,N_17199);
xnor U17306 (N_17306,N_17265,N_17161);
xor U17307 (N_17307,N_17120,N_17175);
xor U17308 (N_17308,N_17229,N_17163);
xor U17309 (N_17309,N_17185,N_17150);
and U17310 (N_17310,N_17227,N_17145);
nor U17311 (N_17311,N_17188,N_17267);
or U17312 (N_17312,N_17124,N_17180);
nor U17313 (N_17313,N_17190,N_17127);
and U17314 (N_17314,N_17186,N_17137);
nand U17315 (N_17315,N_17214,N_17257);
xnor U17316 (N_17316,N_17216,N_17195);
nor U17317 (N_17317,N_17144,N_17243);
and U17318 (N_17318,N_17274,N_17278);
nor U17319 (N_17319,N_17219,N_17189);
and U17320 (N_17320,N_17136,N_17148);
nand U17321 (N_17321,N_17134,N_17209);
and U17322 (N_17322,N_17248,N_17166);
nor U17323 (N_17323,N_17220,N_17225);
nand U17324 (N_17324,N_17254,N_17217);
nand U17325 (N_17325,N_17167,N_17263);
xor U17326 (N_17326,N_17222,N_17203);
nand U17327 (N_17327,N_17141,N_17266);
and U17328 (N_17328,N_17256,N_17158);
xnor U17329 (N_17329,N_17232,N_17168);
nand U17330 (N_17330,N_17187,N_17279);
or U17331 (N_17331,N_17128,N_17165);
xor U17332 (N_17332,N_17269,N_17277);
or U17333 (N_17333,N_17154,N_17129);
nor U17334 (N_17334,N_17147,N_17138);
nor U17335 (N_17335,N_17170,N_17121);
and U17336 (N_17336,N_17122,N_17271);
nor U17337 (N_17337,N_17208,N_17223);
nor U17338 (N_17338,N_17172,N_17152);
and U17339 (N_17339,N_17193,N_17261);
and U17340 (N_17340,N_17153,N_17268);
xor U17341 (N_17341,N_17228,N_17272);
nor U17342 (N_17342,N_17215,N_17194);
or U17343 (N_17343,N_17202,N_17171);
nor U17344 (N_17344,N_17191,N_17207);
xor U17345 (N_17345,N_17205,N_17253);
and U17346 (N_17346,N_17162,N_17146);
or U17347 (N_17347,N_17247,N_17126);
nor U17348 (N_17348,N_17197,N_17135);
xor U17349 (N_17349,N_17149,N_17244);
nor U17350 (N_17350,N_17201,N_17130);
xnor U17351 (N_17351,N_17164,N_17250);
nor U17352 (N_17352,N_17221,N_17270);
nor U17353 (N_17353,N_17157,N_17255);
nand U17354 (N_17354,N_17181,N_17155);
xor U17355 (N_17355,N_17192,N_17230);
xor U17356 (N_17356,N_17236,N_17142);
nor U17357 (N_17357,N_17252,N_17133);
nand U17358 (N_17358,N_17206,N_17204);
or U17359 (N_17359,N_17273,N_17234);
xor U17360 (N_17360,N_17185,N_17215);
nand U17361 (N_17361,N_17187,N_17184);
nor U17362 (N_17362,N_17277,N_17247);
nand U17363 (N_17363,N_17155,N_17197);
nor U17364 (N_17364,N_17147,N_17208);
or U17365 (N_17365,N_17249,N_17229);
or U17366 (N_17366,N_17224,N_17128);
and U17367 (N_17367,N_17268,N_17220);
xnor U17368 (N_17368,N_17158,N_17215);
or U17369 (N_17369,N_17244,N_17200);
nand U17370 (N_17370,N_17176,N_17208);
nor U17371 (N_17371,N_17235,N_17207);
and U17372 (N_17372,N_17151,N_17159);
and U17373 (N_17373,N_17268,N_17264);
xnor U17374 (N_17374,N_17183,N_17186);
nor U17375 (N_17375,N_17165,N_17228);
or U17376 (N_17376,N_17229,N_17123);
xnor U17377 (N_17377,N_17207,N_17276);
nand U17378 (N_17378,N_17277,N_17250);
nor U17379 (N_17379,N_17264,N_17250);
nand U17380 (N_17380,N_17175,N_17233);
nor U17381 (N_17381,N_17130,N_17225);
or U17382 (N_17382,N_17205,N_17250);
xor U17383 (N_17383,N_17198,N_17229);
or U17384 (N_17384,N_17130,N_17127);
and U17385 (N_17385,N_17237,N_17179);
nor U17386 (N_17386,N_17175,N_17143);
nor U17387 (N_17387,N_17216,N_17260);
nand U17388 (N_17388,N_17248,N_17217);
and U17389 (N_17389,N_17147,N_17166);
nor U17390 (N_17390,N_17201,N_17123);
or U17391 (N_17391,N_17272,N_17238);
nor U17392 (N_17392,N_17202,N_17274);
xor U17393 (N_17393,N_17260,N_17257);
nand U17394 (N_17394,N_17251,N_17171);
and U17395 (N_17395,N_17252,N_17179);
and U17396 (N_17396,N_17130,N_17233);
nand U17397 (N_17397,N_17176,N_17194);
nand U17398 (N_17398,N_17141,N_17276);
nor U17399 (N_17399,N_17244,N_17207);
xnor U17400 (N_17400,N_17161,N_17179);
or U17401 (N_17401,N_17161,N_17120);
xnor U17402 (N_17402,N_17267,N_17239);
xor U17403 (N_17403,N_17211,N_17232);
or U17404 (N_17404,N_17271,N_17139);
or U17405 (N_17405,N_17173,N_17249);
nand U17406 (N_17406,N_17254,N_17218);
and U17407 (N_17407,N_17253,N_17167);
xor U17408 (N_17408,N_17275,N_17188);
or U17409 (N_17409,N_17205,N_17263);
and U17410 (N_17410,N_17229,N_17210);
nand U17411 (N_17411,N_17146,N_17231);
xor U17412 (N_17412,N_17236,N_17148);
or U17413 (N_17413,N_17185,N_17209);
nand U17414 (N_17414,N_17143,N_17218);
nor U17415 (N_17415,N_17254,N_17121);
and U17416 (N_17416,N_17128,N_17265);
and U17417 (N_17417,N_17242,N_17226);
nor U17418 (N_17418,N_17208,N_17198);
nor U17419 (N_17419,N_17277,N_17197);
xor U17420 (N_17420,N_17191,N_17171);
xor U17421 (N_17421,N_17232,N_17148);
nor U17422 (N_17422,N_17176,N_17210);
xnor U17423 (N_17423,N_17240,N_17170);
nand U17424 (N_17424,N_17279,N_17140);
xnor U17425 (N_17425,N_17176,N_17166);
nand U17426 (N_17426,N_17165,N_17150);
or U17427 (N_17427,N_17228,N_17241);
or U17428 (N_17428,N_17224,N_17248);
nor U17429 (N_17429,N_17238,N_17196);
nand U17430 (N_17430,N_17250,N_17186);
xnor U17431 (N_17431,N_17205,N_17196);
nor U17432 (N_17432,N_17219,N_17211);
and U17433 (N_17433,N_17138,N_17264);
xnor U17434 (N_17434,N_17153,N_17253);
and U17435 (N_17435,N_17187,N_17203);
xor U17436 (N_17436,N_17173,N_17155);
or U17437 (N_17437,N_17248,N_17174);
nor U17438 (N_17438,N_17217,N_17268);
and U17439 (N_17439,N_17183,N_17139);
and U17440 (N_17440,N_17371,N_17362);
and U17441 (N_17441,N_17380,N_17291);
or U17442 (N_17442,N_17424,N_17342);
nor U17443 (N_17443,N_17347,N_17419);
and U17444 (N_17444,N_17413,N_17361);
or U17445 (N_17445,N_17358,N_17377);
nand U17446 (N_17446,N_17389,N_17406);
or U17447 (N_17447,N_17403,N_17285);
or U17448 (N_17448,N_17308,N_17378);
and U17449 (N_17449,N_17396,N_17420);
or U17450 (N_17450,N_17344,N_17373);
or U17451 (N_17451,N_17417,N_17321);
nor U17452 (N_17452,N_17280,N_17348);
and U17453 (N_17453,N_17346,N_17317);
and U17454 (N_17454,N_17282,N_17414);
nand U17455 (N_17455,N_17426,N_17423);
or U17456 (N_17456,N_17350,N_17387);
xnor U17457 (N_17457,N_17401,N_17310);
nand U17458 (N_17458,N_17372,N_17381);
xnor U17459 (N_17459,N_17370,N_17302);
and U17460 (N_17460,N_17306,N_17296);
nand U17461 (N_17461,N_17399,N_17425);
xnor U17462 (N_17462,N_17297,N_17432);
nor U17463 (N_17463,N_17438,N_17300);
or U17464 (N_17464,N_17304,N_17374);
nor U17465 (N_17465,N_17415,N_17405);
nor U17466 (N_17466,N_17412,N_17299);
xor U17467 (N_17467,N_17295,N_17430);
nor U17468 (N_17468,N_17349,N_17334);
and U17469 (N_17469,N_17286,N_17328);
and U17470 (N_17470,N_17393,N_17305);
and U17471 (N_17471,N_17340,N_17422);
xor U17472 (N_17472,N_17368,N_17345);
or U17473 (N_17473,N_17376,N_17289);
nor U17474 (N_17474,N_17407,N_17307);
xor U17475 (N_17475,N_17433,N_17390);
and U17476 (N_17476,N_17322,N_17319);
nand U17477 (N_17477,N_17324,N_17384);
nor U17478 (N_17478,N_17341,N_17335);
xnor U17479 (N_17479,N_17359,N_17292);
xnor U17480 (N_17480,N_17388,N_17431);
xnor U17481 (N_17481,N_17303,N_17339);
xor U17482 (N_17482,N_17416,N_17287);
and U17483 (N_17483,N_17391,N_17318);
nand U17484 (N_17484,N_17395,N_17379);
nor U17485 (N_17485,N_17313,N_17331);
nor U17486 (N_17486,N_17427,N_17309);
or U17487 (N_17487,N_17367,N_17398);
or U17488 (N_17488,N_17394,N_17337);
or U17489 (N_17489,N_17294,N_17366);
nor U17490 (N_17490,N_17437,N_17386);
and U17491 (N_17491,N_17283,N_17323);
nor U17492 (N_17492,N_17392,N_17336);
xor U17493 (N_17493,N_17353,N_17382);
or U17494 (N_17494,N_17311,N_17428);
nor U17495 (N_17495,N_17333,N_17332);
xor U17496 (N_17496,N_17411,N_17288);
nand U17497 (N_17497,N_17439,N_17397);
and U17498 (N_17498,N_17354,N_17436);
and U17499 (N_17499,N_17365,N_17338);
or U17500 (N_17500,N_17434,N_17363);
and U17501 (N_17501,N_17409,N_17315);
nand U17502 (N_17502,N_17404,N_17355);
nor U17503 (N_17503,N_17429,N_17435);
or U17504 (N_17504,N_17402,N_17325);
nand U17505 (N_17505,N_17330,N_17329);
xnor U17506 (N_17506,N_17298,N_17293);
or U17507 (N_17507,N_17400,N_17326);
nor U17508 (N_17508,N_17352,N_17284);
nand U17509 (N_17509,N_17290,N_17356);
xnor U17510 (N_17510,N_17312,N_17281);
or U17511 (N_17511,N_17410,N_17385);
or U17512 (N_17512,N_17418,N_17421);
and U17513 (N_17513,N_17357,N_17343);
xor U17514 (N_17514,N_17375,N_17316);
nand U17515 (N_17515,N_17351,N_17314);
nand U17516 (N_17516,N_17360,N_17301);
xnor U17517 (N_17517,N_17383,N_17327);
or U17518 (N_17518,N_17369,N_17320);
and U17519 (N_17519,N_17364,N_17408);
nor U17520 (N_17520,N_17401,N_17306);
and U17521 (N_17521,N_17378,N_17345);
or U17522 (N_17522,N_17285,N_17361);
nand U17523 (N_17523,N_17410,N_17396);
and U17524 (N_17524,N_17323,N_17413);
nor U17525 (N_17525,N_17295,N_17418);
or U17526 (N_17526,N_17360,N_17403);
or U17527 (N_17527,N_17296,N_17343);
xor U17528 (N_17528,N_17344,N_17435);
xor U17529 (N_17529,N_17319,N_17405);
and U17530 (N_17530,N_17289,N_17301);
or U17531 (N_17531,N_17288,N_17287);
nor U17532 (N_17532,N_17299,N_17346);
or U17533 (N_17533,N_17436,N_17360);
and U17534 (N_17534,N_17427,N_17347);
nor U17535 (N_17535,N_17351,N_17330);
and U17536 (N_17536,N_17282,N_17307);
or U17537 (N_17537,N_17383,N_17401);
and U17538 (N_17538,N_17337,N_17328);
nand U17539 (N_17539,N_17321,N_17286);
xnor U17540 (N_17540,N_17342,N_17338);
nor U17541 (N_17541,N_17314,N_17371);
nor U17542 (N_17542,N_17408,N_17375);
xnor U17543 (N_17543,N_17298,N_17345);
nand U17544 (N_17544,N_17309,N_17348);
nor U17545 (N_17545,N_17332,N_17301);
nor U17546 (N_17546,N_17421,N_17371);
xnor U17547 (N_17547,N_17439,N_17352);
xnor U17548 (N_17548,N_17294,N_17386);
xnor U17549 (N_17549,N_17289,N_17288);
nand U17550 (N_17550,N_17356,N_17357);
xor U17551 (N_17551,N_17423,N_17330);
and U17552 (N_17552,N_17367,N_17370);
and U17553 (N_17553,N_17410,N_17374);
and U17554 (N_17554,N_17345,N_17379);
nor U17555 (N_17555,N_17298,N_17358);
nand U17556 (N_17556,N_17305,N_17392);
nor U17557 (N_17557,N_17297,N_17382);
nor U17558 (N_17558,N_17392,N_17345);
nand U17559 (N_17559,N_17288,N_17420);
or U17560 (N_17560,N_17434,N_17415);
or U17561 (N_17561,N_17411,N_17305);
xnor U17562 (N_17562,N_17422,N_17403);
nand U17563 (N_17563,N_17354,N_17434);
xnor U17564 (N_17564,N_17356,N_17342);
or U17565 (N_17565,N_17424,N_17353);
nor U17566 (N_17566,N_17393,N_17280);
and U17567 (N_17567,N_17317,N_17331);
and U17568 (N_17568,N_17292,N_17370);
nand U17569 (N_17569,N_17414,N_17310);
nand U17570 (N_17570,N_17330,N_17322);
nor U17571 (N_17571,N_17324,N_17355);
xor U17572 (N_17572,N_17336,N_17434);
nand U17573 (N_17573,N_17346,N_17307);
and U17574 (N_17574,N_17422,N_17320);
nand U17575 (N_17575,N_17349,N_17303);
xnor U17576 (N_17576,N_17360,N_17326);
xnor U17577 (N_17577,N_17394,N_17410);
and U17578 (N_17578,N_17310,N_17376);
and U17579 (N_17579,N_17309,N_17303);
nand U17580 (N_17580,N_17385,N_17387);
xor U17581 (N_17581,N_17390,N_17343);
nor U17582 (N_17582,N_17394,N_17427);
nand U17583 (N_17583,N_17289,N_17341);
or U17584 (N_17584,N_17378,N_17303);
nand U17585 (N_17585,N_17350,N_17366);
or U17586 (N_17586,N_17347,N_17422);
nand U17587 (N_17587,N_17422,N_17336);
nand U17588 (N_17588,N_17300,N_17280);
or U17589 (N_17589,N_17318,N_17355);
xnor U17590 (N_17590,N_17280,N_17431);
and U17591 (N_17591,N_17337,N_17402);
or U17592 (N_17592,N_17374,N_17314);
nor U17593 (N_17593,N_17359,N_17356);
and U17594 (N_17594,N_17310,N_17438);
nor U17595 (N_17595,N_17424,N_17333);
and U17596 (N_17596,N_17315,N_17282);
xor U17597 (N_17597,N_17431,N_17305);
and U17598 (N_17598,N_17438,N_17380);
xnor U17599 (N_17599,N_17419,N_17413);
and U17600 (N_17600,N_17566,N_17562);
nor U17601 (N_17601,N_17521,N_17449);
and U17602 (N_17602,N_17499,N_17508);
nor U17603 (N_17603,N_17597,N_17530);
nor U17604 (N_17604,N_17519,N_17505);
nor U17605 (N_17605,N_17460,N_17573);
and U17606 (N_17606,N_17512,N_17586);
xor U17607 (N_17607,N_17464,N_17487);
nand U17608 (N_17608,N_17448,N_17575);
nor U17609 (N_17609,N_17476,N_17495);
nand U17610 (N_17610,N_17493,N_17561);
and U17611 (N_17611,N_17592,N_17537);
or U17612 (N_17612,N_17558,N_17457);
nor U17613 (N_17613,N_17550,N_17444);
nand U17614 (N_17614,N_17582,N_17552);
or U17615 (N_17615,N_17441,N_17516);
or U17616 (N_17616,N_17470,N_17450);
nand U17617 (N_17617,N_17473,N_17443);
or U17618 (N_17618,N_17480,N_17581);
or U17619 (N_17619,N_17452,N_17477);
or U17620 (N_17620,N_17517,N_17502);
nor U17621 (N_17621,N_17445,N_17446);
or U17622 (N_17622,N_17564,N_17478);
or U17623 (N_17623,N_17568,N_17440);
or U17624 (N_17624,N_17580,N_17447);
nand U17625 (N_17625,N_17551,N_17544);
xnor U17626 (N_17626,N_17567,N_17489);
and U17627 (N_17627,N_17529,N_17509);
and U17628 (N_17628,N_17475,N_17442);
and U17629 (N_17629,N_17599,N_17514);
xor U17630 (N_17630,N_17560,N_17485);
or U17631 (N_17631,N_17462,N_17484);
or U17632 (N_17632,N_17593,N_17583);
nand U17633 (N_17633,N_17526,N_17524);
or U17634 (N_17634,N_17589,N_17574);
and U17635 (N_17635,N_17523,N_17468);
xnor U17636 (N_17636,N_17501,N_17466);
nand U17637 (N_17637,N_17503,N_17534);
nor U17638 (N_17638,N_17556,N_17513);
nand U17639 (N_17639,N_17507,N_17483);
xor U17640 (N_17640,N_17553,N_17458);
and U17641 (N_17641,N_17565,N_17541);
xnor U17642 (N_17642,N_17531,N_17571);
or U17643 (N_17643,N_17522,N_17518);
or U17644 (N_17644,N_17596,N_17510);
and U17645 (N_17645,N_17570,N_17532);
and U17646 (N_17646,N_17472,N_17579);
nand U17647 (N_17647,N_17528,N_17549);
nand U17648 (N_17648,N_17527,N_17525);
xnor U17649 (N_17649,N_17572,N_17465);
or U17650 (N_17650,N_17584,N_17591);
nand U17651 (N_17651,N_17535,N_17590);
xor U17652 (N_17652,N_17533,N_17492);
nand U17653 (N_17653,N_17474,N_17498);
nor U17654 (N_17654,N_17577,N_17481);
or U17655 (N_17655,N_17479,N_17486);
nand U17656 (N_17656,N_17540,N_17578);
nand U17657 (N_17657,N_17482,N_17585);
nor U17658 (N_17658,N_17454,N_17557);
or U17659 (N_17659,N_17471,N_17598);
xor U17660 (N_17660,N_17542,N_17555);
nor U17661 (N_17661,N_17451,N_17543);
xnor U17662 (N_17662,N_17548,N_17459);
xnor U17663 (N_17663,N_17511,N_17461);
nand U17664 (N_17664,N_17504,N_17488);
nor U17665 (N_17665,N_17500,N_17539);
and U17666 (N_17666,N_17559,N_17554);
and U17667 (N_17667,N_17545,N_17569);
xor U17668 (N_17668,N_17520,N_17588);
and U17669 (N_17669,N_17595,N_17576);
nand U17670 (N_17670,N_17469,N_17547);
xor U17671 (N_17671,N_17536,N_17453);
nor U17672 (N_17672,N_17455,N_17515);
nor U17673 (N_17673,N_17494,N_17506);
or U17674 (N_17674,N_17496,N_17594);
xor U17675 (N_17675,N_17546,N_17491);
xnor U17676 (N_17676,N_17463,N_17497);
xnor U17677 (N_17677,N_17456,N_17563);
nor U17678 (N_17678,N_17587,N_17467);
nor U17679 (N_17679,N_17538,N_17490);
and U17680 (N_17680,N_17471,N_17547);
and U17681 (N_17681,N_17579,N_17508);
and U17682 (N_17682,N_17477,N_17506);
xor U17683 (N_17683,N_17444,N_17478);
xnor U17684 (N_17684,N_17541,N_17521);
xnor U17685 (N_17685,N_17501,N_17448);
or U17686 (N_17686,N_17447,N_17543);
nor U17687 (N_17687,N_17594,N_17586);
nand U17688 (N_17688,N_17502,N_17584);
and U17689 (N_17689,N_17452,N_17526);
nand U17690 (N_17690,N_17587,N_17525);
or U17691 (N_17691,N_17447,N_17525);
nand U17692 (N_17692,N_17454,N_17556);
xnor U17693 (N_17693,N_17479,N_17441);
nor U17694 (N_17694,N_17507,N_17441);
nor U17695 (N_17695,N_17555,N_17561);
nor U17696 (N_17696,N_17485,N_17557);
nand U17697 (N_17697,N_17536,N_17596);
xnor U17698 (N_17698,N_17524,N_17532);
xnor U17699 (N_17699,N_17557,N_17575);
xnor U17700 (N_17700,N_17506,N_17521);
nand U17701 (N_17701,N_17475,N_17512);
nor U17702 (N_17702,N_17583,N_17464);
and U17703 (N_17703,N_17572,N_17579);
nor U17704 (N_17704,N_17444,N_17480);
xnor U17705 (N_17705,N_17496,N_17579);
and U17706 (N_17706,N_17479,N_17523);
or U17707 (N_17707,N_17534,N_17526);
and U17708 (N_17708,N_17599,N_17546);
or U17709 (N_17709,N_17534,N_17492);
nand U17710 (N_17710,N_17528,N_17589);
and U17711 (N_17711,N_17460,N_17599);
nand U17712 (N_17712,N_17528,N_17522);
nor U17713 (N_17713,N_17562,N_17516);
nor U17714 (N_17714,N_17560,N_17466);
or U17715 (N_17715,N_17585,N_17596);
nor U17716 (N_17716,N_17548,N_17542);
xor U17717 (N_17717,N_17464,N_17531);
nand U17718 (N_17718,N_17552,N_17452);
and U17719 (N_17719,N_17483,N_17532);
nor U17720 (N_17720,N_17503,N_17510);
nand U17721 (N_17721,N_17563,N_17454);
and U17722 (N_17722,N_17521,N_17465);
nor U17723 (N_17723,N_17456,N_17588);
and U17724 (N_17724,N_17519,N_17590);
xor U17725 (N_17725,N_17471,N_17447);
and U17726 (N_17726,N_17512,N_17472);
or U17727 (N_17727,N_17476,N_17579);
nand U17728 (N_17728,N_17514,N_17493);
xnor U17729 (N_17729,N_17563,N_17559);
and U17730 (N_17730,N_17598,N_17526);
nand U17731 (N_17731,N_17490,N_17568);
or U17732 (N_17732,N_17531,N_17539);
or U17733 (N_17733,N_17504,N_17474);
nand U17734 (N_17734,N_17444,N_17534);
and U17735 (N_17735,N_17578,N_17525);
nand U17736 (N_17736,N_17492,N_17498);
nor U17737 (N_17737,N_17518,N_17457);
and U17738 (N_17738,N_17593,N_17534);
nor U17739 (N_17739,N_17500,N_17570);
xor U17740 (N_17740,N_17599,N_17451);
nand U17741 (N_17741,N_17598,N_17594);
and U17742 (N_17742,N_17579,N_17521);
xnor U17743 (N_17743,N_17463,N_17517);
and U17744 (N_17744,N_17549,N_17578);
or U17745 (N_17745,N_17596,N_17558);
xor U17746 (N_17746,N_17543,N_17495);
or U17747 (N_17747,N_17443,N_17458);
and U17748 (N_17748,N_17453,N_17567);
nor U17749 (N_17749,N_17497,N_17590);
or U17750 (N_17750,N_17452,N_17576);
xor U17751 (N_17751,N_17516,N_17571);
nor U17752 (N_17752,N_17529,N_17581);
nand U17753 (N_17753,N_17509,N_17551);
nor U17754 (N_17754,N_17485,N_17453);
nand U17755 (N_17755,N_17476,N_17479);
xor U17756 (N_17756,N_17592,N_17576);
or U17757 (N_17757,N_17536,N_17551);
nor U17758 (N_17758,N_17598,N_17498);
or U17759 (N_17759,N_17532,N_17563);
and U17760 (N_17760,N_17721,N_17630);
nor U17761 (N_17761,N_17734,N_17751);
or U17762 (N_17762,N_17756,N_17740);
nand U17763 (N_17763,N_17674,N_17714);
nand U17764 (N_17764,N_17754,N_17745);
nor U17765 (N_17765,N_17696,N_17733);
nor U17766 (N_17766,N_17729,N_17632);
xor U17767 (N_17767,N_17614,N_17689);
nand U17768 (N_17768,N_17727,N_17669);
and U17769 (N_17769,N_17616,N_17753);
nor U17770 (N_17770,N_17722,N_17750);
nor U17771 (N_17771,N_17724,N_17601);
nor U17772 (N_17772,N_17672,N_17739);
nand U17773 (N_17773,N_17702,N_17715);
nand U17774 (N_17774,N_17752,N_17723);
nand U17775 (N_17775,N_17652,N_17608);
or U17776 (N_17776,N_17638,N_17675);
nand U17777 (N_17777,N_17660,N_17704);
nand U17778 (N_17778,N_17634,N_17617);
nand U17779 (N_17779,N_17755,N_17639);
nand U17780 (N_17780,N_17695,N_17736);
nor U17781 (N_17781,N_17659,N_17662);
or U17782 (N_17782,N_17631,N_17667);
xor U17783 (N_17783,N_17717,N_17694);
and U17784 (N_17784,N_17624,N_17666);
nor U17785 (N_17785,N_17637,N_17613);
and U17786 (N_17786,N_17627,N_17742);
or U17787 (N_17787,N_17730,N_17629);
or U17788 (N_17788,N_17748,N_17758);
nand U17789 (N_17789,N_17757,N_17670);
nand U17790 (N_17790,N_17744,N_17658);
nand U17791 (N_17791,N_17690,N_17684);
and U17792 (N_17792,N_17641,N_17655);
or U17793 (N_17793,N_17607,N_17643);
nor U17794 (N_17794,N_17633,N_17610);
nor U17795 (N_17795,N_17626,N_17625);
nand U17796 (N_17796,N_17686,N_17743);
nor U17797 (N_17797,N_17720,N_17716);
xor U17798 (N_17798,N_17620,N_17651);
nand U17799 (N_17799,N_17703,N_17621);
xnor U17800 (N_17800,N_17680,N_17635);
and U17801 (N_17801,N_17709,N_17713);
nor U17802 (N_17802,N_17678,N_17640);
or U17803 (N_17803,N_17623,N_17600);
or U17804 (N_17804,N_17712,N_17692);
or U17805 (N_17805,N_17691,N_17603);
or U17806 (N_17806,N_17693,N_17653);
or U17807 (N_17807,N_17645,N_17700);
and U17808 (N_17808,N_17622,N_17650);
nor U17809 (N_17809,N_17759,N_17687);
or U17810 (N_17810,N_17731,N_17708);
nand U17811 (N_17811,N_17609,N_17699);
or U17812 (N_17812,N_17719,N_17701);
nand U17813 (N_17813,N_17648,N_17654);
or U17814 (N_17814,N_17698,N_17611);
xor U17815 (N_17815,N_17682,N_17732);
nor U17816 (N_17816,N_17705,N_17649);
xor U17817 (N_17817,N_17728,N_17642);
and U17818 (N_17818,N_17697,N_17663);
nand U17819 (N_17819,N_17668,N_17661);
nor U17820 (N_17820,N_17688,N_17707);
xor U17821 (N_17821,N_17636,N_17615);
nor U17822 (N_17822,N_17747,N_17606);
xnor U17823 (N_17823,N_17683,N_17646);
or U17824 (N_17824,N_17710,N_17673);
or U17825 (N_17825,N_17749,N_17644);
and U17826 (N_17826,N_17618,N_17738);
nor U17827 (N_17827,N_17725,N_17679);
or U17828 (N_17828,N_17718,N_17746);
or U17829 (N_17829,N_17602,N_17605);
nor U17830 (N_17830,N_17671,N_17619);
xor U17831 (N_17831,N_17665,N_17657);
xnor U17832 (N_17832,N_17681,N_17677);
and U17833 (N_17833,N_17604,N_17711);
or U17834 (N_17834,N_17656,N_17735);
xnor U17835 (N_17835,N_17741,N_17706);
nand U17836 (N_17836,N_17647,N_17737);
and U17837 (N_17837,N_17676,N_17685);
and U17838 (N_17838,N_17726,N_17628);
nand U17839 (N_17839,N_17664,N_17612);
nor U17840 (N_17840,N_17603,N_17648);
and U17841 (N_17841,N_17624,N_17615);
nand U17842 (N_17842,N_17674,N_17752);
nor U17843 (N_17843,N_17658,N_17637);
and U17844 (N_17844,N_17711,N_17674);
xor U17845 (N_17845,N_17709,N_17603);
xnor U17846 (N_17846,N_17707,N_17745);
xnor U17847 (N_17847,N_17640,N_17719);
or U17848 (N_17848,N_17745,N_17631);
xnor U17849 (N_17849,N_17603,N_17726);
and U17850 (N_17850,N_17625,N_17606);
or U17851 (N_17851,N_17671,N_17698);
nand U17852 (N_17852,N_17747,N_17755);
xnor U17853 (N_17853,N_17639,N_17707);
or U17854 (N_17854,N_17706,N_17753);
and U17855 (N_17855,N_17718,N_17627);
nand U17856 (N_17856,N_17745,N_17759);
or U17857 (N_17857,N_17637,N_17698);
nor U17858 (N_17858,N_17636,N_17618);
nor U17859 (N_17859,N_17754,N_17713);
and U17860 (N_17860,N_17661,N_17628);
nand U17861 (N_17861,N_17687,N_17650);
nand U17862 (N_17862,N_17726,N_17691);
and U17863 (N_17863,N_17616,N_17615);
nor U17864 (N_17864,N_17624,N_17692);
and U17865 (N_17865,N_17703,N_17668);
xnor U17866 (N_17866,N_17638,N_17691);
or U17867 (N_17867,N_17714,N_17699);
xnor U17868 (N_17868,N_17637,N_17746);
nand U17869 (N_17869,N_17655,N_17757);
nor U17870 (N_17870,N_17605,N_17673);
or U17871 (N_17871,N_17722,N_17705);
nor U17872 (N_17872,N_17610,N_17694);
xnor U17873 (N_17873,N_17623,N_17696);
nor U17874 (N_17874,N_17700,N_17692);
xor U17875 (N_17875,N_17656,N_17668);
and U17876 (N_17876,N_17756,N_17691);
nand U17877 (N_17877,N_17732,N_17610);
and U17878 (N_17878,N_17662,N_17708);
and U17879 (N_17879,N_17629,N_17745);
xor U17880 (N_17880,N_17752,N_17727);
nor U17881 (N_17881,N_17737,N_17689);
nand U17882 (N_17882,N_17733,N_17680);
nor U17883 (N_17883,N_17707,N_17667);
xnor U17884 (N_17884,N_17755,N_17751);
nor U17885 (N_17885,N_17709,N_17690);
or U17886 (N_17886,N_17725,N_17740);
nor U17887 (N_17887,N_17739,N_17699);
nor U17888 (N_17888,N_17617,N_17735);
xor U17889 (N_17889,N_17670,N_17672);
and U17890 (N_17890,N_17692,N_17758);
and U17891 (N_17891,N_17709,N_17660);
or U17892 (N_17892,N_17646,N_17754);
nand U17893 (N_17893,N_17670,N_17617);
nor U17894 (N_17894,N_17711,N_17665);
nand U17895 (N_17895,N_17717,N_17720);
nand U17896 (N_17896,N_17728,N_17683);
or U17897 (N_17897,N_17685,N_17658);
nor U17898 (N_17898,N_17611,N_17681);
xor U17899 (N_17899,N_17621,N_17607);
nand U17900 (N_17900,N_17631,N_17617);
or U17901 (N_17901,N_17603,N_17659);
nor U17902 (N_17902,N_17605,N_17695);
and U17903 (N_17903,N_17743,N_17675);
xor U17904 (N_17904,N_17709,N_17723);
xnor U17905 (N_17905,N_17628,N_17603);
and U17906 (N_17906,N_17629,N_17708);
or U17907 (N_17907,N_17724,N_17680);
and U17908 (N_17908,N_17661,N_17691);
xnor U17909 (N_17909,N_17652,N_17705);
xor U17910 (N_17910,N_17677,N_17614);
or U17911 (N_17911,N_17658,N_17679);
or U17912 (N_17912,N_17740,N_17643);
or U17913 (N_17913,N_17749,N_17610);
nor U17914 (N_17914,N_17626,N_17735);
or U17915 (N_17915,N_17672,N_17743);
nor U17916 (N_17916,N_17721,N_17608);
xnor U17917 (N_17917,N_17625,N_17670);
and U17918 (N_17918,N_17605,N_17662);
nand U17919 (N_17919,N_17665,N_17729);
and U17920 (N_17920,N_17810,N_17912);
and U17921 (N_17921,N_17808,N_17788);
nand U17922 (N_17922,N_17883,N_17872);
or U17923 (N_17923,N_17828,N_17915);
xor U17924 (N_17924,N_17791,N_17901);
or U17925 (N_17925,N_17896,N_17880);
nand U17926 (N_17926,N_17802,N_17878);
nand U17927 (N_17927,N_17794,N_17893);
and U17928 (N_17928,N_17778,N_17816);
or U17929 (N_17929,N_17917,N_17824);
nand U17930 (N_17930,N_17913,N_17780);
xor U17931 (N_17931,N_17787,N_17905);
nor U17932 (N_17932,N_17823,N_17800);
nand U17933 (N_17933,N_17836,N_17786);
nor U17934 (N_17934,N_17907,N_17798);
nor U17935 (N_17935,N_17840,N_17850);
or U17936 (N_17936,N_17783,N_17813);
nor U17937 (N_17937,N_17879,N_17809);
and U17938 (N_17938,N_17849,N_17826);
nand U17939 (N_17939,N_17887,N_17890);
and U17940 (N_17940,N_17868,N_17910);
nand U17941 (N_17941,N_17863,N_17908);
nand U17942 (N_17942,N_17906,N_17785);
xnor U17943 (N_17943,N_17769,N_17861);
xnor U17944 (N_17944,N_17807,N_17857);
nor U17945 (N_17945,N_17875,N_17873);
nor U17946 (N_17946,N_17762,N_17851);
and U17947 (N_17947,N_17889,N_17886);
and U17948 (N_17948,N_17845,N_17792);
and U17949 (N_17949,N_17773,N_17830);
nor U17950 (N_17950,N_17866,N_17843);
and U17951 (N_17951,N_17871,N_17898);
nand U17952 (N_17952,N_17820,N_17877);
or U17953 (N_17953,N_17835,N_17881);
or U17954 (N_17954,N_17795,N_17774);
nand U17955 (N_17955,N_17844,N_17834);
or U17956 (N_17956,N_17888,N_17862);
nor U17957 (N_17957,N_17856,N_17831);
xor U17958 (N_17958,N_17895,N_17860);
and U17959 (N_17959,N_17892,N_17869);
xnor U17960 (N_17960,N_17819,N_17760);
xor U17961 (N_17961,N_17891,N_17918);
or U17962 (N_17962,N_17885,N_17846);
nand U17963 (N_17963,N_17781,N_17867);
or U17964 (N_17964,N_17799,N_17827);
or U17965 (N_17965,N_17822,N_17833);
xnor U17966 (N_17966,N_17796,N_17900);
xnor U17967 (N_17967,N_17801,N_17865);
xnor U17968 (N_17968,N_17852,N_17870);
xor U17969 (N_17969,N_17847,N_17777);
and U17970 (N_17970,N_17776,N_17817);
nand U17971 (N_17971,N_17804,N_17858);
or U17972 (N_17972,N_17837,N_17770);
or U17973 (N_17973,N_17771,N_17818);
nand U17974 (N_17974,N_17812,N_17789);
nor U17975 (N_17975,N_17897,N_17805);
nand U17976 (N_17976,N_17853,N_17784);
nand U17977 (N_17977,N_17876,N_17761);
nor U17978 (N_17978,N_17821,N_17848);
or U17979 (N_17979,N_17864,N_17764);
and U17980 (N_17980,N_17766,N_17829);
xor U17981 (N_17981,N_17768,N_17779);
and U17982 (N_17982,N_17884,N_17814);
nor U17983 (N_17983,N_17911,N_17811);
or U17984 (N_17984,N_17838,N_17825);
xor U17985 (N_17985,N_17832,N_17797);
xnor U17986 (N_17986,N_17904,N_17767);
nand U17987 (N_17987,N_17874,N_17775);
nand U17988 (N_17988,N_17854,N_17899);
nand U17989 (N_17989,N_17765,N_17815);
nor U17990 (N_17990,N_17782,N_17859);
or U17991 (N_17991,N_17916,N_17806);
or U17992 (N_17992,N_17772,N_17855);
xor U17993 (N_17993,N_17882,N_17839);
nand U17994 (N_17994,N_17841,N_17909);
nor U17995 (N_17995,N_17903,N_17790);
xnor U17996 (N_17996,N_17919,N_17894);
and U17997 (N_17997,N_17914,N_17793);
or U17998 (N_17998,N_17902,N_17842);
nand U17999 (N_17999,N_17803,N_17763);
nor U18000 (N_18000,N_17826,N_17823);
xor U18001 (N_18001,N_17784,N_17793);
nand U18002 (N_18002,N_17850,N_17847);
xor U18003 (N_18003,N_17870,N_17875);
nor U18004 (N_18004,N_17778,N_17856);
xor U18005 (N_18005,N_17872,N_17841);
xor U18006 (N_18006,N_17913,N_17774);
and U18007 (N_18007,N_17788,N_17820);
nand U18008 (N_18008,N_17800,N_17863);
nor U18009 (N_18009,N_17783,N_17871);
or U18010 (N_18010,N_17910,N_17763);
xnor U18011 (N_18011,N_17780,N_17776);
and U18012 (N_18012,N_17826,N_17913);
xor U18013 (N_18013,N_17880,N_17870);
and U18014 (N_18014,N_17789,N_17823);
nand U18015 (N_18015,N_17793,N_17897);
and U18016 (N_18016,N_17771,N_17907);
or U18017 (N_18017,N_17768,N_17814);
nand U18018 (N_18018,N_17780,N_17892);
or U18019 (N_18019,N_17876,N_17898);
nand U18020 (N_18020,N_17877,N_17788);
or U18021 (N_18021,N_17906,N_17909);
nor U18022 (N_18022,N_17817,N_17818);
nor U18023 (N_18023,N_17883,N_17809);
and U18024 (N_18024,N_17802,N_17767);
xnor U18025 (N_18025,N_17901,N_17894);
and U18026 (N_18026,N_17815,N_17766);
or U18027 (N_18027,N_17781,N_17888);
nand U18028 (N_18028,N_17780,N_17888);
and U18029 (N_18029,N_17800,N_17812);
nor U18030 (N_18030,N_17900,N_17786);
or U18031 (N_18031,N_17857,N_17912);
nor U18032 (N_18032,N_17801,N_17773);
xor U18033 (N_18033,N_17818,N_17834);
or U18034 (N_18034,N_17787,N_17851);
and U18035 (N_18035,N_17890,N_17889);
nor U18036 (N_18036,N_17767,N_17914);
xnor U18037 (N_18037,N_17914,N_17892);
xor U18038 (N_18038,N_17807,N_17773);
xnor U18039 (N_18039,N_17851,N_17883);
or U18040 (N_18040,N_17901,N_17902);
and U18041 (N_18041,N_17807,N_17817);
and U18042 (N_18042,N_17777,N_17919);
and U18043 (N_18043,N_17902,N_17772);
or U18044 (N_18044,N_17897,N_17858);
or U18045 (N_18045,N_17797,N_17825);
and U18046 (N_18046,N_17879,N_17878);
and U18047 (N_18047,N_17816,N_17774);
and U18048 (N_18048,N_17813,N_17866);
and U18049 (N_18049,N_17831,N_17797);
and U18050 (N_18050,N_17911,N_17840);
nor U18051 (N_18051,N_17808,N_17900);
nor U18052 (N_18052,N_17879,N_17820);
nor U18053 (N_18053,N_17760,N_17867);
and U18054 (N_18054,N_17864,N_17891);
and U18055 (N_18055,N_17786,N_17826);
xnor U18056 (N_18056,N_17836,N_17892);
nor U18057 (N_18057,N_17805,N_17834);
nand U18058 (N_18058,N_17918,N_17820);
nand U18059 (N_18059,N_17771,N_17816);
and U18060 (N_18060,N_17872,N_17853);
or U18061 (N_18061,N_17856,N_17762);
nand U18062 (N_18062,N_17765,N_17828);
or U18063 (N_18063,N_17775,N_17797);
nand U18064 (N_18064,N_17801,N_17883);
or U18065 (N_18065,N_17845,N_17816);
or U18066 (N_18066,N_17807,N_17889);
nor U18067 (N_18067,N_17871,N_17889);
nand U18068 (N_18068,N_17780,N_17813);
xnor U18069 (N_18069,N_17890,N_17913);
or U18070 (N_18070,N_17824,N_17856);
xnor U18071 (N_18071,N_17803,N_17859);
xnor U18072 (N_18072,N_17859,N_17905);
nor U18073 (N_18073,N_17856,N_17870);
xor U18074 (N_18074,N_17848,N_17862);
xnor U18075 (N_18075,N_17852,N_17909);
or U18076 (N_18076,N_17807,N_17823);
and U18077 (N_18077,N_17900,N_17913);
and U18078 (N_18078,N_17803,N_17892);
or U18079 (N_18079,N_17873,N_17783);
or U18080 (N_18080,N_17966,N_18029);
nor U18081 (N_18081,N_17951,N_17932);
or U18082 (N_18082,N_18008,N_17930);
nand U18083 (N_18083,N_18005,N_18057);
nor U18084 (N_18084,N_17922,N_18063);
nand U18085 (N_18085,N_17943,N_18003);
or U18086 (N_18086,N_17974,N_18041);
xnor U18087 (N_18087,N_17978,N_18023);
or U18088 (N_18088,N_17959,N_17992);
nand U18089 (N_18089,N_18025,N_18055);
nand U18090 (N_18090,N_18067,N_18020);
and U18091 (N_18091,N_17969,N_17928);
or U18092 (N_18092,N_18038,N_18032);
or U18093 (N_18093,N_18033,N_18068);
and U18094 (N_18094,N_18026,N_17970);
and U18095 (N_18095,N_18030,N_17926);
nor U18096 (N_18096,N_18037,N_17947);
and U18097 (N_18097,N_18053,N_17984);
xor U18098 (N_18098,N_17968,N_18028);
or U18099 (N_18099,N_17942,N_17954);
nand U18100 (N_18100,N_17962,N_17950);
or U18101 (N_18101,N_17931,N_18064);
or U18102 (N_18102,N_17973,N_18052);
nand U18103 (N_18103,N_17940,N_17971);
and U18104 (N_18104,N_17993,N_18016);
nor U18105 (N_18105,N_17925,N_18010);
and U18106 (N_18106,N_18062,N_17997);
nor U18107 (N_18107,N_18056,N_18024);
xnor U18108 (N_18108,N_18011,N_18061);
and U18109 (N_18109,N_18077,N_17952);
xnor U18110 (N_18110,N_17923,N_17976);
nand U18111 (N_18111,N_18043,N_18022);
or U18112 (N_18112,N_17980,N_17987);
xor U18113 (N_18113,N_18050,N_17946);
or U18114 (N_18114,N_18031,N_18078);
xnor U18115 (N_18115,N_18047,N_18048);
xor U18116 (N_18116,N_18040,N_17988);
or U18117 (N_18117,N_17965,N_18034);
or U18118 (N_18118,N_17972,N_18035);
or U18119 (N_18119,N_17998,N_17982);
xor U18120 (N_18120,N_18072,N_18051);
or U18121 (N_18121,N_17955,N_17957);
or U18122 (N_18122,N_17991,N_18045);
and U18123 (N_18123,N_17989,N_18074);
nand U18124 (N_18124,N_17956,N_17994);
and U18125 (N_18125,N_17927,N_17939);
xor U18126 (N_18126,N_17920,N_18070);
nor U18127 (N_18127,N_18013,N_17967);
nor U18128 (N_18128,N_17929,N_17981);
nand U18129 (N_18129,N_18076,N_17986);
xnor U18130 (N_18130,N_17958,N_17948);
and U18131 (N_18131,N_17999,N_18065);
nor U18132 (N_18132,N_17953,N_18017);
and U18133 (N_18133,N_18060,N_17941);
and U18134 (N_18134,N_18004,N_18069);
and U18135 (N_18135,N_18000,N_17960);
nor U18136 (N_18136,N_17990,N_17996);
xnor U18137 (N_18137,N_18027,N_17963);
xor U18138 (N_18138,N_18018,N_18015);
nand U18139 (N_18139,N_17934,N_17985);
nand U18140 (N_18140,N_17936,N_18039);
xnor U18141 (N_18141,N_18044,N_17937);
xor U18142 (N_18142,N_18073,N_17979);
nand U18143 (N_18143,N_17995,N_18014);
or U18144 (N_18144,N_17933,N_17921);
and U18145 (N_18145,N_17938,N_17924);
or U18146 (N_18146,N_18006,N_18036);
or U18147 (N_18147,N_18009,N_18002);
nor U18148 (N_18148,N_17949,N_18042);
nand U18149 (N_18149,N_18046,N_18071);
nand U18150 (N_18150,N_18001,N_17944);
and U18151 (N_18151,N_18054,N_18058);
nor U18152 (N_18152,N_18021,N_17977);
or U18153 (N_18153,N_17945,N_17983);
and U18154 (N_18154,N_18079,N_18019);
xnor U18155 (N_18155,N_18007,N_18066);
and U18156 (N_18156,N_18075,N_17964);
or U18157 (N_18157,N_18059,N_18012);
nand U18158 (N_18158,N_17935,N_17961);
and U18159 (N_18159,N_17975,N_18049);
nand U18160 (N_18160,N_18056,N_17947);
or U18161 (N_18161,N_17925,N_17994);
nand U18162 (N_18162,N_18016,N_17955);
or U18163 (N_18163,N_18051,N_18006);
nor U18164 (N_18164,N_17953,N_18048);
or U18165 (N_18165,N_17982,N_17980);
or U18166 (N_18166,N_18014,N_18050);
and U18167 (N_18167,N_17976,N_18013);
nor U18168 (N_18168,N_17962,N_17953);
and U18169 (N_18169,N_18069,N_17963);
xnor U18170 (N_18170,N_17949,N_17953);
nand U18171 (N_18171,N_17956,N_17995);
and U18172 (N_18172,N_18023,N_18046);
nor U18173 (N_18173,N_17994,N_18051);
and U18174 (N_18174,N_17954,N_17941);
nor U18175 (N_18175,N_18025,N_17938);
nor U18176 (N_18176,N_17993,N_17973);
and U18177 (N_18177,N_17974,N_18068);
nand U18178 (N_18178,N_17948,N_18040);
xnor U18179 (N_18179,N_17980,N_18002);
and U18180 (N_18180,N_18050,N_17958);
xor U18181 (N_18181,N_17976,N_18029);
nand U18182 (N_18182,N_18071,N_17944);
nor U18183 (N_18183,N_17928,N_17943);
nand U18184 (N_18184,N_17993,N_18054);
nor U18185 (N_18185,N_18002,N_18055);
xor U18186 (N_18186,N_17932,N_18001);
xnor U18187 (N_18187,N_18015,N_18047);
nor U18188 (N_18188,N_17984,N_18069);
and U18189 (N_18189,N_17967,N_17936);
nor U18190 (N_18190,N_18000,N_18013);
nor U18191 (N_18191,N_17926,N_18074);
xnor U18192 (N_18192,N_17935,N_18009);
or U18193 (N_18193,N_17947,N_18034);
and U18194 (N_18194,N_17978,N_17932);
nor U18195 (N_18195,N_17950,N_17957);
or U18196 (N_18196,N_17950,N_18030);
and U18197 (N_18197,N_17949,N_17952);
nor U18198 (N_18198,N_17965,N_18069);
nor U18199 (N_18199,N_18049,N_18040);
nand U18200 (N_18200,N_18019,N_17942);
xor U18201 (N_18201,N_17953,N_17985);
xnor U18202 (N_18202,N_18072,N_18022);
and U18203 (N_18203,N_17924,N_17955);
or U18204 (N_18204,N_18011,N_17949);
xnor U18205 (N_18205,N_17925,N_17993);
nand U18206 (N_18206,N_17985,N_17976);
and U18207 (N_18207,N_17999,N_18049);
nor U18208 (N_18208,N_17988,N_17961);
xnor U18209 (N_18209,N_17953,N_18021);
xnor U18210 (N_18210,N_17948,N_18068);
xor U18211 (N_18211,N_18059,N_18035);
and U18212 (N_18212,N_18033,N_18050);
xor U18213 (N_18213,N_17969,N_17971);
and U18214 (N_18214,N_17936,N_17983);
nor U18215 (N_18215,N_17972,N_17977);
nor U18216 (N_18216,N_17961,N_17933);
nand U18217 (N_18217,N_18077,N_17998);
nand U18218 (N_18218,N_17925,N_18043);
or U18219 (N_18219,N_18029,N_17934);
nor U18220 (N_18220,N_17951,N_17987);
nor U18221 (N_18221,N_18003,N_18021);
nor U18222 (N_18222,N_18015,N_17939);
nor U18223 (N_18223,N_17948,N_18048);
and U18224 (N_18224,N_17997,N_17935);
and U18225 (N_18225,N_17961,N_18015);
xor U18226 (N_18226,N_18047,N_18049);
or U18227 (N_18227,N_17961,N_17951);
or U18228 (N_18228,N_17920,N_18008);
or U18229 (N_18229,N_17932,N_18060);
or U18230 (N_18230,N_18074,N_18005);
xnor U18231 (N_18231,N_18032,N_17994);
xor U18232 (N_18232,N_18008,N_17927);
xor U18233 (N_18233,N_17998,N_18015);
nor U18234 (N_18234,N_17924,N_17996);
or U18235 (N_18235,N_18076,N_18075);
nor U18236 (N_18236,N_17961,N_18007);
nand U18237 (N_18237,N_17994,N_17937);
or U18238 (N_18238,N_17924,N_17954);
xnor U18239 (N_18239,N_17979,N_17955);
and U18240 (N_18240,N_18117,N_18219);
or U18241 (N_18241,N_18083,N_18105);
xor U18242 (N_18242,N_18140,N_18124);
or U18243 (N_18243,N_18141,N_18188);
nor U18244 (N_18244,N_18118,N_18143);
nand U18245 (N_18245,N_18183,N_18090);
nor U18246 (N_18246,N_18130,N_18147);
nand U18247 (N_18247,N_18096,N_18210);
nand U18248 (N_18248,N_18095,N_18205);
xnor U18249 (N_18249,N_18223,N_18165);
xnor U18250 (N_18250,N_18080,N_18217);
and U18251 (N_18251,N_18166,N_18100);
or U18252 (N_18252,N_18198,N_18093);
nor U18253 (N_18253,N_18151,N_18175);
nand U18254 (N_18254,N_18142,N_18137);
and U18255 (N_18255,N_18185,N_18234);
xnor U18256 (N_18256,N_18162,N_18216);
nor U18257 (N_18257,N_18203,N_18215);
or U18258 (N_18258,N_18220,N_18170);
nand U18259 (N_18259,N_18239,N_18094);
nand U18260 (N_18260,N_18156,N_18120);
nor U18261 (N_18261,N_18098,N_18213);
or U18262 (N_18262,N_18089,N_18115);
and U18263 (N_18263,N_18082,N_18121);
nor U18264 (N_18264,N_18152,N_18233);
nor U18265 (N_18265,N_18101,N_18212);
and U18266 (N_18266,N_18214,N_18133);
nor U18267 (N_18267,N_18107,N_18085);
nand U18268 (N_18268,N_18086,N_18110);
or U18269 (N_18269,N_18148,N_18102);
xnor U18270 (N_18270,N_18172,N_18202);
nand U18271 (N_18271,N_18138,N_18211);
and U18272 (N_18272,N_18197,N_18111);
nand U18273 (N_18273,N_18108,N_18139);
and U18274 (N_18274,N_18128,N_18134);
or U18275 (N_18275,N_18081,N_18237);
or U18276 (N_18276,N_18168,N_18208);
and U18277 (N_18277,N_18158,N_18123);
nor U18278 (N_18278,N_18225,N_18125);
or U18279 (N_18279,N_18174,N_18222);
nor U18280 (N_18280,N_18238,N_18160);
or U18281 (N_18281,N_18195,N_18145);
and U18282 (N_18282,N_18109,N_18099);
nor U18283 (N_18283,N_18149,N_18119);
and U18284 (N_18284,N_18224,N_18169);
and U18285 (N_18285,N_18154,N_18182);
or U18286 (N_18286,N_18229,N_18113);
xnor U18287 (N_18287,N_18088,N_18181);
and U18288 (N_18288,N_18227,N_18173);
xor U18289 (N_18289,N_18193,N_18207);
xnor U18290 (N_18290,N_18112,N_18209);
nor U18291 (N_18291,N_18129,N_18230);
or U18292 (N_18292,N_18201,N_18114);
and U18293 (N_18293,N_18159,N_18155);
xnor U18294 (N_18294,N_18231,N_18127);
nand U18295 (N_18295,N_18189,N_18097);
nor U18296 (N_18296,N_18091,N_18132);
nand U18297 (N_18297,N_18186,N_18200);
or U18298 (N_18298,N_18221,N_18164);
xnor U18299 (N_18299,N_18192,N_18150);
or U18300 (N_18300,N_18204,N_18177);
or U18301 (N_18301,N_18218,N_18180);
xnor U18302 (N_18302,N_18194,N_18126);
nand U18303 (N_18303,N_18092,N_18104);
and U18304 (N_18304,N_18232,N_18236);
nand U18305 (N_18305,N_18146,N_18199);
or U18306 (N_18306,N_18228,N_18161);
xnor U18307 (N_18307,N_18135,N_18131);
xnor U18308 (N_18308,N_18206,N_18178);
xor U18309 (N_18309,N_18122,N_18190);
nor U18310 (N_18310,N_18084,N_18187);
and U18311 (N_18311,N_18167,N_18144);
nand U18312 (N_18312,N_18103,N_18184);
nand U18313 (N_18313,N_18171,N_18176);
nand U18314 (N_18314,N_18226,N_18153);
or U18315 (N_18315,N_18106,N_18235);
nand U18316 (N_18316,N_18087,N_18116);
nand U18317 (N_18317,N_18157,N_18179);
and U18318 (N_18318,N_18136,N_18196);
nor U18319 (N_18319,N_18191,N_18163);
or U18320 (N_18320,N_18158,N_18098);
xor U18321 (N_18321,N_18101,N_18156);
xnor U18322 (N_18322,N_18232,N_18146);
nand U18323 (N_18323,N_18112,N_18224);
xnor U18324 (N_18324,N_18081,N_18238);
and U18325 (N_18325,N_18177,N_18163);
nor U18326 (N_18326,N_18188,N_18203);
nor U18327 (N_18327,N_18138,N_18213);
and U18328 (N_18328,N_18200,N_18139);
nor U18329 (N_18329,N_18182,N_18140);
nor U18330 (N_18330,N_18116,N_18083);
nand U18331 (N_18331,N_18140,N_18221);
or U18332 (N_18332,N_18135,N_18111);
nor U18333 (N_18333,N_18211,N_18216);
nor U18334 (N_18334,N_18115,N_18157);
or U18335 (N_18335,N_18106,N_18217);
and U18336 (N_18336,N_18099,N_18153);
nor U18337 (N_18337,N_18151,N_18198);
or U18338 (N_18338,N_18144,N_18143);
nand U18339 (N_18339,N_18153,N_18118);
and U18340 (N_18340,N_18216,N_18144);
xor U18341 (N_18341,N_18194,N_18191);
xor U18342 (N_18342,N_18220,N_18238);
xor U18343 (N_18343,N_18139,N_18136);
and U18344 (N_18344,N_18157,N_18193);
xnor U18345 (N_18345,N_18123,N_18175);
nand U18346 (N_18346,N_18228,N_18154);
and U18347 (N_18347,N_18174,N_18202);
or U18348 (N_18348,N_18197,N_18086);
and U18349 (N_18349,N_18229,N_18176);
and U18350 (N_18350,N_18082,N_18080);
nand U18351 (N_18351,N_18219,N_18209);
and U18352 (N_18352,N_18193,N_18166);
nor U18353 (N_18353,N_18172,N_18158);
nand U18354 (N_18354,N_18123,N_18236);
nor U18355 (N_18355,N_18082,N_18192);
or U18356 (N_18356,N_18177,N_18194);
or U18357 (N_18357,N_18104,N_18233);
and U18358 (N_18358,N_18205,N_18112);
and U18359 (N_18359,N_18128,N_18165);
or U18360 (N_18360,N_18199,N_18157);
and U18361 (N_18361,N_18168,N_18129);
nand U18362 (N_18362,N_18199,N_18219);
xor U18363 (N_18363,N_18207,N_18110);
or U18364 (N_18364,N_18177,N_18107);
xor U18365 (N_18365,N_18178,N_18224);
and U18366 (N_18366,N_18128,N_18141);
or U18367 (N_18367,N_18222,N_18224);
nand U18368 (N_18368,N_18238,N_18161);
xor U18369 (N_18369,N_18235,N_18175);
xnor U18370 (N_18370,N_18096,N_18191);
and U18371 (N_18371,N_18164,N_18203);
nor U18372 (N_18372,N_18158,N_18203);
and U18373 (N_18373,N_18200,N_18130);
or U18374 (N_18374,N_18201,N_18212);
and U18375 (N_18375,N_18107,N_18082);
or U18376 (N_18376,N_18192,N_18086);
xor U18377 (N_18377,N_18173,N_18116);
or U18378 (N_18378,N_18130,N_18174);
nor U18379 (N_18379,N_18129,N_18229);
nand U18380 (N_18380,N_18212,N_18196);
nor U18381 (N_18381,N_18210,N_18211);
nor U18382 (N_18382,N_18226,N_18182);
nand U18383 (N_18383,N_18207,N_18114);
nand U18384 (N_18384,N_18095,N_18197);
nor U18385 (N_18385,N_18107,N_18181);
xnor U18386 (N_18386,N_18086,N_18093);
xor U18387 (N_18387,N_18224,N_18135);
nand U18388 (N_18388,N_18179,N_18232);
nand U18389 (N_18389,N_18221,N_18092);
nand U18390 (N_18390,N_18139,N_18093);
and U18391 (N_18391,N_18164,N_18235);
nand U18392 (N_18392,N_18085,N_18143);
or U18393 (N_18393,N_18175,N_18202);
or U18394 (N_18394,N_18112,N_18231);
or U18395 (N_18395,N_18235,N_18212);
nand U18396 (N_18396,N_18168,N_18100);
and U18397 (N_18397,N_18120,N_18155);
or U18398 (N_18398,N_18219,N_18100);
nor U18399 (N_18399,N_18222,N_18106);
nand U18400 (N_18400,N_18295,N_18244);
nand U18401 (N_18401,N_18366,N_18376);
or U18402 (N_18402,N_18283,N_18292);
nor U18403 (N_18403,N_18320,N_18242);
and U18404 (N_18404,N_18378,N_18276);
or U18405 (N_18405,N_18312,N_18270);
nor U18406 (N_18406,N_18279,N_18371);
and U18407 (N_18407,N_18265,N_18319);
xnor U18408 (N_18408,N_18256,N_18345);
xnor U18409 (N_18409,N_18374,N_18336);
or U18410 (N_18410,N_18309,N_18253);
nor U18411 (N_18411,N_18348,N_18385);
nand U18412 (N_18412,N_18354,N_18264);
and U18413 (N_18413,N_18271,N_18325);
xor U18414 (N_18414,N_18393,N_18373);
xnor U18415 (N_18415,N_18329,N_18307);
and U18416 (N_18416,N_18269,N_18261);
nand U18417 (N_18417,N_18350,N_18394);
or U18418 (N_18418,N_18395,N_18257);
nand U18419 (N_18419,N_18397,N_18268);
and U18420 (N_18420,N_18260,N_18275);
or U18421 (N_18421,N_18344,N_18252);
or U18422 (N_18422,N_18390,N_18273);
nor U18423 (N_18423,N_18249,N_18304);
nand U18424 (N_18424,N_18347,N_18266);
nand U18425 (N_18425,N_18316,N_18298);
or U18426 (N_18426,N_18372,N_18381);
and U18427 (N_18427,N_18301,N_18321);
xor U18428 (N_18428,N_18246,N_18313);
nand U18429 (N_18429,N_18291,N_18379);
nand U18430 (N_18430,N_18251,N_18326);
and U18431 (N_18431,N_18392,N_18310);
xnor U18432 (N_18432,N_18284,N_18388);
xnor U18433 (N_18433,N_18303,N_18367);
or U18434 (N_18434,N_18353,N_18290);
nand U18435 (N_18435,N_18255,N_18258);
xnor U18436 (N_18436,N_18342,N_18331);
nand U18437 (N_18437,N_18360,N_18280);
nor U18438 (N_18438,N_18262,N_18384);
nand U18439 (N_18439,N_18382,N_18287);
nor U18440 (N_18440,N_18240,N_18351);
nand U18441 (N_18441,N_18338,N_18259);
nor U18442 (N_18442,N_18334,N_18274);
nand U18443 (N_18443,N_18386,N_18375);
and U18444 (N_18444,N_18289,N_18306);
or U18445 (N_18445,N_18327,N_18370);
xor U18446 (N_18446,N_18272,N_18300);
or U18447 (N_18447,N_18317,N_18391);
nor U18448 (N_18448,N_18352,N_18356);
and U18449 (N_18449,N_18357,N_18302);
xnor U18450 (N_18450,N_18314,N_18318);
and U18451 (N_18451,N_18340,N_18363);
xor U18452 (N_18452,N_18254,N_18267);
and U18453 (N_18453,N_18365,N_18343);
nor U18454 (N_18454,N_18278,N_18311);
xnor U18455 (N_18455,N_18297,N_18263);
and U18456 (N_18456,N_18355,N_18296);
xnor U18457 (N_18457,N_18294,N_18364);
nand U18458 (N_18458,N_18349,N_18341);
and U18459 (N_18459,N_18399,N_18247);
or U18460 (N_18460,N_18248,N_18377);
xor U18461 (N_18461,N_18332,N_18362);
nor U18462 (N_18462,N_18305,N_18346);
nor U18463 (N_18463,N_18333,N_18361);
xnor U18464 (N_18464,N_18369,N_18398);
nand U18465 (N_18465,N_18285,N_18339);
xnor U18466 (N_18466,N_18293,N_18299);
nand U18467 (N_18467,N_18323,N_18250);
or U18468 (N_18468,N_18245,N_18380);
nand U18469 (N_18469,N_18330,N_18308);
and U18470 (N_18470,N_18359,N_18322);
nand U18471 (N_18471,N_18396,N_18387);
nand U18472 (N_18472,N_18241,N_18383);
nand U18473 (N_18473,N_18368,N_18243);
or U18474 (N_18474,N_18288,N_18337);
nor U18475 (N_18475,N_18328,N_18277);
or U18476 (N_18476,N_18389,N_18315);
and U18477 (N_18477,N_18281,N_18324);
or U18478 (N_18478,N_18282,N_18286);
and U18479 (N_18479,N_18358,N_18335);
nand U18480 (N_18480,N_18301,N_18268);
nor U18481 (N_18481,N_18324,N_18325);
nor U18482 (N_18482,N_18397,N_18391);
nor U18483 (N_18483,N_18257,N_18300);
nor U18484 (N_18484,N_18280,N_18319);
nand U18485 (N_18485,N_18389,N_18394);
or U18486 (N_18486,N_18261,N_18297);
and U18487 (N_18487,N_18242,N_18267);
nor U18488 (N_18488,N_18289,N_18371);
nor U18489 (N_18489,N_18275,N_18314);
and U18490 (N_18490,N_18345,N_18356);
and U18491 (N_18491,N_18373,N_18305);
nor U18492 (N_18492,N_18283,N_18316);
and U18493 (N_18493,N_18341,N_18284);
xor U18494 (N_18494,N_18399,N_18328);
xnor U18495 (N_18495,N_18328,N_18265);
and U18496 (N_18496,N_18262,N_18315);
and U18497 (N_18497,N_18345,N_18292);
or U18498 (N_18498,N_18374,N_18350);
and U18499 (N_18499,N_18269,N_18358);
or U18500 (N_18500,N_18321,N_18373);
or U18501 (N_18501,N_18263,N_18258);
nor U18502 (N_18502,N_18261,N_18248);
nand U18503 (N_18503,N_18372,N_18320);
nor U18504 (N_18504,N_18327,N_18273);
xor U18505 (N_18505,N_18247,N_18384);
nor U18506 (N_18506,N_18378,N_18242);
xnor U18507 (N_18507,N_18266,N_18264);
nand U18508 (N_18508,N_18345,N_18349);
or U18509 (N_18509,N_18265,N_18367);
nor U18510 (N_18510,N_18337,N_18357);
nor U18511 (N_18511,N_18302,N_18263);
nor U18512 (N_18512,N_18258,N_18292);
nor U18513 (N_18513,N_18383,N_18242);
or U18514 (N_18514,N_18260,N_18368);
xnor U18515 (N_18515,N_18390,N_18256);
or U18516 (N_18516,N_18348,N_18389);
nor U18517 (N_18517,N_18271,N_18277);
or U18518 (N_18518,N_18281,N_18358);
and U18519 (N_18519,N_18260,N_18266);
nor U18520 (N_18520,N_18331,N_18379);
nor U18521 (N_18521,N_18342,N_18337);
and U18522 (N_18522,N_18261,N_18360);
nand U18523 (N_18523,N_18279,N_18342);
nor U18524 (N_18524,N_18384,N_18351);
or U18525 (N_18525,N_18280,N_18333);
xnor U18526 (N_18526,N_18346,N_18271);
and U18527 (N_18527,N_18371,N_18328);
xor U18528 (N_18528,N_18345,N_18340);
and U18529 (N_18529,N_18396,N_18240);
nor U18530 (N_18530,N_18282,N_18270);
or U18531 (N_18531,N_18399,N_18267);
nor U18532 (N_18532,N_18361,N_18248);
nor U18533 (N_18533,N_18359,N_18244);
and U18534 (N_18534,N_18316,N_18274);
or U18535 (N_18535,N_18274,N_18391);
and U18536 (N_18536,N_18383,N_18313);
xnor U18537 (N_18537,N_18391,N_18322);
and U18538 (N_18538,N_18330,N_18358);
and U18539 (N_18539,N_18323,N_18259);
nand U18540 (N_18540,N_18314,N_18399);
xor U18541 (N_18541,N_18257,N_18363);
nor U18542 (N_18542,N_18359,N_18330);
xnor U18543 (N_18543,N_18344,N_18333);
or U18544 (N_18544,N_18242,N_18265);
nand U18545 (N_18545,N_18335,N_18300);
nor U18546 (N_18546,N_18389,N_18365);
xor U18547 (N_18547,N_18343,N_18270);
and U18548 (N_18548,N_18260,N_18320);
or U18549 (N_18549,N_18385,N_18316);
and U18550 (N_18550,N_18377,N_18296);
or U18551 (N_18551,N_18326,N_18282);
or U18552 (N_18552,N_18338,N_18250);
xor U18553 (N_18553,N_18382,N_18251);
nand U18554 (N_18554,N_18249,N_18305);
or U18555 (N_18555,N_18297,N_18340);
and U18556 (N_18556,N_18261,N_18384);
nor U18557 (N_18557,N_18371,N_18312);
xor U18558 (N_18558,N_18325,N_18388);
nor U18559 (N_18559,N_18249,N_18277);
xnor U18560 (N_18560,N_18534,N_18519);
or U18561 (N_18561,N_18533,N_18454);
nand U18562 (N_18562,N_18433,N_18481);
xor U18563 (N_18563,N_18476,N_18434);
nor U18564 (N_18564,N_18490,N_18493);
xor U18565 (N_18565,N_18477,N_18409);
and U18566 (N_18566,N_18511,N_18544);
nor U18567 (N_18567,N_18558,N_18497);
nor U18568 (N_18568,N_18529,N_18412);
or U18569 (N_18569,N_18448,N_18553);
xnor U18570 (N_18570,N_18522,N_18542);
xor U18571 (N_18571,N_18479,N_18410);
nand U18572 (N_18572,N_18458,N_18530);
nor U18573 (N_18573,N_18482,N_18469);
xor U18574 (N_18574,N_18506,N_18431);
or U18575 (N_18575,N_18512,N_18452);
nor U18576 (N_18576,N_18543,N_18464);
and U18577 (N_18577,N_18527,N_18403);
nor U18578 (N_18578,N_18461,N_18402);
nor U18579 (N_18579,N_18516,N_18442);
nor U18580 (N_18580,N_18541,N_18438);
xnor U18581 (N_18581,N_18473,N_18429);
nor U18582 (N_18582,N_18449,N_18524);
or U18583 (N_18583,N_18457,N_18540);
or U18584 (N_18584,N_18548,N_18445);
nand U18585 (N_18585,N_18441,N_18414);
nor U18586 (N_18586,N_18455,N_18514);
and U18587 (N_18587,N_18470,N_18510);
xnor U18588 (N_18588,N_18401,N_18420);
xnor U18589 (N_18589,N_18430,N_18509);
or U18590 (N_18590,N_18502,N_18496);
nand U18591 (N_18591,N_18538,N_18494);
or U18592 (N_18592,N_18507,N_18468);
and U18593 (N_18593,N_18480,N_18537);
or U18594 (N_18594,N_18549,N_18499);
nand U18595 (N_18595,N_18484,N_18536);
nand U18596 (N_18596,N_18466,N_18450);
nor U18597 (N_18597,N_18526,N_18525);
nand U18598 (N_18598,N_18460,N_18491);
and U18599 (N_18599,N_18451,N_18475);
and U18600 (N_18600,N_18486,N_18472);
and U18601 (N_18601,N_18417,N_18547);
nand U18602 (N_18602,N_18415,N_18520);
or U18603 (N_18603,N_18453,N_18418);
nand U18604 (N_18604,N_18423,N_18551);
or U18605 (N_18605,N_18413,N_18446);
and U18606 (N_18606,N_18531,N_18424);
xor U18607 (N_18607,N_18463,N_18556);
xor U18608 (N_18608,N_18515,N_18545);
nor U18609 (N_18609,N_18488,N_18421);
nand U18610 (N_18610,N_18444,N_18419);
xor U18611 (N_18611,N_18428,N_18485);
xnor U18612 (N_18612,N_18439,N_18539);
or U18613 (N_18613,N_18503,N_18426);
and U18614 (N_18614,N_18436,N_18513);
nor U18615 (N_18615,N_18443,N_18555);
nand U18616 (N_18616,N_18416,N_18489);
nor U18617 (N_18617,N_18504,N_18546);
and U18618 (N_18618,N_18404,N_18535);
or U18619 (N_18619,N_18523,N_18427);
nand U18620 (N_18620,N_18501,N_18500);
nor U18621 (N_18621,N_18550,N_18467);
nor U18622 (N_18622,N_18405,N_18462);
and U18623 (N_18623,N_18456,N_18517);
nor U18624 (N_18624,N_18411,N_18406);
nand U18625 (N_18625,N_18554,N_18432);
nor U18626 (N_18626,N_18498,N_18487);
xnor U18627 (N_18627,N_18492,N_18440);
or U18628 (N_18628,N_18478,N_18557);
nand U18629 (N_18629,N_18465,N_18447);
xnor U18630 (N_18630,N_18474,N_18508);
or U18631 (N_18631,N_18532,N_18559);
nand U18632 (N_18632,N_18521,N_18407);
nand U18633 (N_18633,N_18425,N_18408);
nand U18634 (N_18634,N_18459,N_18518);
nand U18635 (N_18635,N_18471,N_18437);
and U18636 (N_18636,N_18435,N_18552);
nor U18637 (N_18637,N_18400,N_18528);
and U18638 (N_18638,N_18422,N_18495);
xnor U18639 (N_18639,N_18483,N_18505);
xor U18640 (N_18640,N_18482,N_18523);
or U18641 (N_18641,N_18497,N_18435);
nor U18642 (N_18642,N_18502,N_18480);
nor U18643 (N_18643,N_18529,N_18557);
xor U18644 (N_18644,N_18484,N_18485);
or U18645 (N_18645,N_18415,N_18483);
nor U18646 (N_18646,N_18478,N_18518);
nand U18647 (N_18647,N_18417,N_18542);
and U18648 (N_18648,N_18512,N_18462);
and U18649 (N_18649,N_18539,N_18465);
xor U18650 (N_18650,N_18400,N_18501);
nand U18651 (N_18651,N_18525,N_18460);
nor U18652 (N_18652,N_18486,N_18469);
xnor U18653 (N_18653,N_18446,N_18500);
nor U18654 (N_18654,N_18433,N_18488);
and U18655 (N_18655,N_18428,N_18503);
xor U18656 (N_18656,N_18469,N_18445);
nand U18657 (N_18657,N_18504,N_18423);
and U18658 (N_18658,N_18465,N_18537);
nor U18659 (N_18659,N_18495,N_18470);
or U18660 (N_18660,N_18517,N_18467);
and U18661 (N_18661,N_18515,N_18414);
xor U18662 (N_18662,N_18545,N_18447);
nor U18663 (N_18663,N_18467,N_18453);
nor U18664 (N_18664,N_18519,N_18452);
or U18665 (N_18665,N_18511,N_18499);
and U18666 (N_18666,N_18405,N_18501);
nand U18667 (N_18667,N_18516,N_18437);
nand U18668 (N_18668,N_18415,N_18406);
xnor U18669 (N_18669,N_18442,N_18513);
nand U18670 (N_18670,N_18497,N_18523);
or U18671 (N_18671,N_18531,N_18555);
and U18672 (N_18672,N_18545,N_18525);
nand U18673 (N_18673,N_18559,N_18464);
or U18674 (N_18674,N_18422,N_18473);
nor U18675 (N_18675,N_18511,N_18559);
and U18676 (N_18676,N_18479,N_18477);
and U18677 (N_18677,N_18426,N_18445);
and U18678 (N_18678,N_18469,N_18414);
or U18679 (N_18679,N_18553,N_18495);
or U18680 (N_18680,N_18483,N_18555);
nor U18681 (N_18681,N_18467,N_18488);
nor U18682 (N_18682,N_18426,N_18423);
nand U18683 (N_18683,N_18540,N_18412);
nand U18684 (N_18684,N_18499,N_18470);
and U18685 (N_18685,N_18503,N_18518);
nand U18686 (N_18686,N_18539,N_18529);
nand U18687 (N_18687,N_18408,N_18481);
nand U18688 (N_18688,N_18419,N_18506);
or U18689 (N_18689,N_18456,N_18451);
and U18690 (N_18690,N_18424,N_18513);
or U18691 (N_18691,N_18430,N_18402);
xnor U18692 (N_18692,N_18502,N_18447);
nor U18693 (N_18693,N_18467,N_18502);
nor U18694 (N_18694,N_18486,N_18405);
or U18695 (N_18695,N_18451,N_18527);
nand U18696 (N_18696,N_18536,N_18485);
or U18697 (N_18697,N_18488,N_18490);
nor U18698 (N_18698,N_18525,N_18466);
and U18699 (N_18699,N_18430,N_18486);
nor U18700 (N_18700,N_18526,N_18522);
nor U18701 (N_18701,N_18437,N_18510);
xor U18702 (N_18702,N_18452,N_18417);
nor U18703 (N_18703,N_18437,N_18411);
and U18704 (N_18704,N_18444,N_18475);
nor U18705 (N_18705,N_18518,N_18472);
nand U18706 (N_18706,N_18488,N_18454);
or U18707 (N_18707,N_18557,N_18516);
and U18708 (N_18708,N_18518,N_18493);
and U18709 (N_18709,N_18547,N_18545);
xnor U18710 (N_18710,N_18401,N_18554);
or U18711 (N_18711,N_18511,N_18517);
xor U18712 (N_18712,N_18426,N_18455);
nor U18713 (N_18713,N_18416,N_18409);
nor U18714 (N_18714,N_18423,N_18464);
nand U18715 (N_18715,N_18527,N_18506);
nand U18716 (N_18716,N_18527,N_18479);
or U18717 (N_18717,N_18537,N_18440);
nor U18718 (N_18718,N_18493,N_18520);
and U18719 (N_18719,N_18402,N_18469);
xnor U18720 (N_18720,N_18567,N_18704);
or U18721 (N_18721,N_18579,N_18695);
xor U18722 (N_18722,N_18698,N_18686);
nand U18723 (N_18723,N_18628,N_18633);
or U18724 (N_18724,N_18574,N_18651);
nor U18725 (N_18725,N_18596,N_18636);
nor U18726 (N_18726,N_18621,N_18625);
xor U18727 (N_18727,N_18587,N_18610);
xor U18728 (N_18728,N_18661,N_18662);
xnor U18729 (N_18729,N_18673,N_18649);
xor U18730 (N_18730,N_18577,N_18672);
and U18731 (N_18731,N_18658,N_18639);
and U18732 (N_18732,N_18588,N_18646);
nand U18733 (N_18733,N_18714,N_18643);
or U18734 (N_18734,N_18705,N_18575);
and U18735 (N_18735,N_18681,N_18602);
or U18736 (N_18736,N_18664,N_18583);
xnor U18737 (N_18737,N_18582,N_18683);
and U18738 (N_18738,N_18570,N_18654);
nor U18739 (N_18739,N_18604,N_18612);
nand U18740 (N_18740,N_18709,N_18632);
xor U18741 (N_18741,N_18663,N_18678);
nand U18742 (N_18742,N_18617,N_18690);
nand U18743 (N_18743,N_18707,N_18680);
and U18744 (N_18744,N_18711,N_18679);
and U18745 (N_18745,N_18716,N_18675);
or U18746 (N_18746,N_18631,N_18691);
and U18747 (N_18747,N_18689,N_18605);
xnor U18748 (N_18748,N_18568,N_18569);
and U18749 (N_18749,N_18710,N_18626);
or U18750 (N_18750,N_18589,N_18597);
nor U18751 (N_18751,N_18644,N_18702);
nand U18752 (N_18752,N_18708,N_18692);
nor U18753 (N_18753,N_18667,N_18627);
xnor U18754 (N_18754,N_18655,N_18635);
or U18755 (N_18755,N_18624,N_18677);
nor U18756 (N_18756,N_18674,N_18593);
and U18757 (N_18757,N_18614,N_18685);
nor U18758 (N_18758,N_18562,N_18600);
and U18759 (N_18759,N_18706,N_18585);
nor U18760 (N_18760,N_18630,N_18634);
or U18761 (N_18761,N_18608,N_18609);
and U18762 (N_18762,N_18696,N_18561);
and U18763 (N_18763,N_18670,N_18712);
nand U18764 (N_18764,N_18599,N_18688);
or U18765 (N_18765,N_18697,N_18703);
or U18766 (N_18766,N_18616,N_18648);
and U18767 (N_18767,N_18607,N_18563);
nand U18768 (N_18768,N_18573,N_18606);
nand U18769 (N_18769,N_18642,N_18715);
and U18770 (N_18770,N_18701,N_18629);
xnor U18771 (N_18771,N_18717,N_18700);
nand U18772 (N_18772,N_18718,N_18598);
and U18773 (N_18773,N_18571,N_18578);
xor U18774 (N_18774,N_18671,N_18659);
xnor U18775 (N_18775,N_18668,N_18693);
and U18776 (N_18776,N_18637,N_18613);
and U18777 (N_18777,N_18581,N_18699);
nor U18778 (N_18778,N_18618,N_18653);
xnor U18779 (N_18779,N_18566,N_18687);
or U18780 (N_18780,N_18565,N_18611);
xnor U18781 (N_18781,N_18592,N_18623);
xnor U18782 (N_18782,N_18719,N_18650);
nor U18783 (N_18783,N_18594,N_18591);
nand U18784 (N_18784,N_18590,N_18665);
or U18785 (N_18785,N_18640,N_18586);
xnor U18786 (N_18786,N_18622,N_18684);
or U18787 (N_18787,N_18682,N_18694);
or U18788 (N_18788,N_18656,N_18669);
xor U18789 (N_18789,N_18564,N_18572);
and U18790 (N_18790,N_18645,N_18615);
xor U18791 (N_18791,N_18601,N_18560);
nor U18792 (N_18792,N_18619,N_18603);
or U18793 (N_18793,N_18584,N_18576);
or U18794 (N_18794,N_18713,N_18666);
xor U18795 (N_18795,N_18652,N_18638);
xnor U18796 (N_18796,N_18660,N_18595);
or U18797 (N_18797,N_18641,N_18676);
nand U18798 (N_18798,N_18657,N_18620);
nor U18799 (N_18799,N_18647,N_18580);
or U18800 (N_18800,N_18632,N_18651);
nand U18801 (N_18801,N_18679,N_18680);
or U18802 (N_18802,N_18685,N_18609);
xnor U18803 (N_18803,N_18679,N_18664);
nand U18804 (N_18804,N_18569,N_18636);
nand U18805 (N_18805,N_18668,N_18565);
or U18806 (N_18806,N_18702,N_18642);
nand U18807 (N_18807,N_18561,N_18569);
or U18808 (N_18808,N_18678,N_18698);
xor U18809 (N_18809,N_18566,N_18673);
or U18810 (N_18810,N_18622,N_18630);
or U18811 (N_18811,N_18670,N_18588);
and U18812 (N_18812,N_18714,N_18706);
nor U18813 (N_18813,N_18609,N_18710);
xnor U18814 (N_18814,N_18654,N_18637);
and U18815 (N_18815,N_18569,N_18678);
and U18816 (N_18816,N_18566,N_18600);
xor U18817 (N_18817,N_18670,N_18637);
or U18818 (N_18818,N_18599,N_18665);
and U18819 (N_18819,N_18711,N_18618);
xnor U18820 (N_18820,N_18620,N_18686);
and U18821 (N_18821,N_18587,N_18663);
nor U18822 (N_18822,N_18567,N_18615);
xnor U18823 (N_18823,N_18698,N_18597);
or U18824 (N_18824,N_18618,N_18669);
xnor U18825 (N_18825,N_18673,N_18565);
and U18826 (N_18826,N_18611,N_18579);
nand U18827 (N_18827,N_18560,N_18700);
nor U18828 (N_18828,N_18679,N_18634);
nand U18829 (N_18829,N_18695,N_18692);
and U18830 (N_18830,N_18585,N_18666);
and U18831 (N_18831,N_18567,N_18699);
and U18832 (N_18832,N_18707,N_18618);
xor U18833 (N_18833,N_18565,N_18699);
or U18834 (N_18834,N_18672,N_18563);
nand U18835 (N_18835,N_18684,N_18588);
and U18836 (N_18836,N_18663,N_18679);
and U18837 (N_18837,N_18674,N_18579);
nand U18838 (N_18838,N_18715,N_18580);
nor U18839 (N_18839,N_18607,N_18613);
nand U18840 (N_18840,N_18657,N_18659);
nor U18841 (N_18841,N_18696,N_18652);
xnor U18842 (N_18842,N_18609,N_18666);
xnor U18843 (N_18843,N_18702,N_18599);
nand U18844 (N_18844,N_18690,N_18585);
nand U18845 (N_18845,N_18654,N_18655);
or U18846 (N_18846,N_18654,N_18618);
nand U18847 (N_18847,N_18617,N_18587);
xor U18848 (N_18848,N_18659,N_18585);
xnor U18849 (N_18849,N_18676,N_18659);
or U18850 (N_18850,N_18588,N_18650);
and U18851 (N_18851,N_18692,N_18680);
xnor U18852 (N_18852,N_18628,N_18641);
xnor U18853 (N_18853,N_18655,N_18639);
nor U18854 (N_18854,N_18684,N_18654);
nor U18855 (N_18855,N_18629,N_18658);
or U18856 (N_18856,N_18631,N_18678);
nand U18857 (N_18857,N_18612,N_18567);
xnor U18858 (N_18858,N_18611,N_18615);
xor U18859 (N_18859,N_18675,N_18584);
xnor U18860 (N_18860,N_18582,N_18634);
xor U18861 (N_18861,N_18571,N_18659);
xor U18862 (N_18862,N_18609,N_18573);
nor U18863 (N_18863,N_18592,N_18654);
or U18864 (N_18864,N_18636,N_18688);
nor U18865 (N_18865,N_18644,N_18658);
and U18866 (N_18866,N_18663,N_18573);
xnor U18867 (N_18867,N_18677,N_18675);
xor U18868 (N_18868,N_18681,N_18578);
xor U18869 (N_18869,N_18565,N_18615);
or U18870 (N_18870,N_18562,N_18676);
and U18871 (N_18871,N_18718,N_18657);
xor U18872 (N_18872,N_18698,N_18671);
nand U18873 (N_18873,N_18673,N_18610);
and U18874 (N_18874,N_18655,N_18651);
or U18875 (N_18875,N_18618,N_18688);
nor U18876 (N_18876,N_18709,N_18678);
or U18877 (N_18877,N_18656,N_18681);
and U18878 (N_18878,N_18580,N_18634);
or U18879 (N_18879,N_18589,N_18588);
or U18880 (N_18880,N_18736,N_18831);
or U18881 (N_18881,N_18759,N_18745);
nor U18882 (N_18882,N_18754,N_18852);
nand U18883 (N_18883,N_18766,N_18721);
xor U18884 (N_18884,N_18750,N_18844);
nor U18885 (N_18885,N_18830,N_18791);
xnor U18886 (N_18886,N_18864,N_18738);
xnor U18887 (N_18887,N_18775,N_18764);
or U18888 (N_18888,N_18787,N_18724);
and U18889 (N_18889,N_18833,N_18863);
and U18890 (N_18890,N_18826,N_18836);
xor U18891 (N_18891,N_18794,N_18825);
nor U18892 (N_18892,N_18835,N_18788);
and U18893 (N_18893,N_18756,N_18869);
nand U18894 (N_18894,N_18870,N_18734);
nor U18895 (N_18895,N_18768,N_18757);
nand U18896 (N_18896,N_18808,N_18868);
xor U18897 (N_18897,N_18815,N_18779);
nand U18898 (N_18898,N_18726,N_18873);
and U18899 (N_18899,N_18824,N_18871);
or U18900 (N_18900,N_18729,N_18748);
xnor U18901 (N_18901,N_18781,N_18780);
and U18902 (N_18902,N_18840,N_18733);
and U18903 (N_18903,N_18798,N_18846);
nand U18904 (N_18904,N_18720,N_18742);
xor U18905 (N_18905,N_18799,N_18834);
and U18906 (N_18906,N_18839,N_18829);
or U18907 (N_18907,N_18802,N_18743);
nand U18908 (N_18908,N_18760,N_18805);
nand U18909 (N_18909,N_18803,N_18744);
and U18910 (N_18910,N_18854,N_18811);
xor U18911 (N_18911,N_18741,N_18731);
or U18912 (N_18912,N_18758,N_18849);
nor U18913 (N_18913,N_18827,N_18763);
xor U18914 (N_18914,N_18772,N_18751);
nor U18915 (N_18915,N_18752,N_18774);
nand U18916 (N_18916,N_18874,N_18821);
and U18917 (N_18917,N_18806,N_18876);
xnor U18918 (N_18918,N_18819,N_18816);
and U18919 (N_18919,N_18861,N_18796);
xor U18920 (N_18920,N_18858,N_18786);
xnor U18921 (N_18921,N_18770,N_18812);
or U18922 (N_18922,N_18732,N_18860);
or U18923 (N_18923,N_18793,N_18822);
xor U18924 (N_18924,N_18730,N_18777);
or U18925 (N_18925,N_18867,N_18761);
and U18926 (N_18926,N_18747,N_18776);
or U18927 (N_18927,N_18801,N_18800);
nand U18928 (N_18928,N_18845,N_18878);
or U18929 (N_18929,N_18784,N_18749);
nor U18930 (N_18930,N_18737,N_18875);
nand U18931 (N_18931,N_18820,N_18856);
nor U18932 (N_18932,N_18848,N_18837);
nand U18933 (N_18933,N_18813,N_18790);
nand U18934 (N_18934,N_18722,N_18843);
and U18935 (N_18935,N_18725,N_18728);
and U18936 (N_18936,N_18767,N_18782);
nand U18937 (N_18937,N_18872,N_18771);
nor U18938 (N_18938,N_18851,N_18789);
and U18939 (N_18939,N_18818,N_18866);
nand U18940 (N_18940,N_18740,N_18865);
or U18941 (N_18941,N_18797,N_18823);
xnor U18942 (N_18942,N_18765,N_18735);
nand U18943 (N_18943,N_18809,N_18769);
nor U18944 (N_18944,N_18828,N_18755);
nand U18945 (N_18945,N_18792,N_18841);
xor U18946 (N_18946,N_18804,N_18859);
nand U18947 (N_18947,N_18773,N_18783);
or U18948 (N_18948,N_18807,N_18877);
xor U18949 (N_18949,N_18810,N_18753);
and U18950 (N_18950,N_18817,N_18853);
and U18951 (N_18951,N_18727,N_18879);
or U18952 (N_18952,N_18832,N_18842);
or U18953 (N_18953,N_18723,N_18795);
or U18954 (N_18954,N_18855,N_18739);
and U18955 (N_18955,N_18838,N_18857);
nor U18956 (N_18956,N_18847,N_18814);
or U18957 (N_18957,N_18778,N_18862);
and U18958 (N_18958,N_18785,N_18762);
nand U18959 (N_18959,N_18746,N_18850);
xor U18960 (N_18960,N_18784,N_18751);
nand U18961 (N_18961,N_18827,N_18849);
xor U18962 (N_18962,N_18754,N_18723);
xnor U18963 (N_18963,N_18768,N_18786);
nand U18964 (N_18964,N_18735,N_18779);
xor U18965 (N_18965,N_18845,N_18818);
or U18966 (N_18966,N_18868,N_18767);
or U18967 (N_18967,N_18760,N_18821);
nor U18968 (N_18968,N_18798,N_18814);
xnor U18969 (N_18969,N_18834,N_18829);
and U18970 (N_18970,N_18793,N_18735);
and U18971 (N_18971,N_18852,N_18729);
nand U18972 (N_18972,N_18772,N_18861);
xor U18973 (N_18973,N_18868,N_18727);
and U18974 (N_18974,N_18793,N_18721);
xnor U18975 (N_18975,N_18819,N_18809);
and U18976 (N_18976,N_18787,N_18865);
or U18977 (N_18977,N_18753,N_18737);
or U18978 (N_18978,N_18851,N_18787);
nor U18979 (N_18979,N_18725,N_18833);
and U18980 (N_18980,N_18802,N_18746);
or U18981 (N_18981,N_18790,N_18755);
and U18982 (N_18982,N_18852,N_18763);
xnor U18983 (N_18983,N_18842,N_18740);
and U18984 (N_18984,N_18849,N_18757);
xnor U18985 (N_18985,N_18839,N_18837);
and U18986 (N_18986,N_18736,N_18804);
nand U18987 (N_18987,N_18727,N_18877);
xnor U18988 (N_18988,N_18754,N_18755);
nand U18989 (N_18989,N_18768,N_18874);
nor U18990 (N_18990,N_18782,N_18739);
xnor U18991 (N_18991,N_18762,N_18832);
and U18992 (N_18992,N_18769,N_18876);
xnor U18993 (N_18993,N_18746,N_18771);
nor U18994 (N_18994,N_18879,N_18731);
and U18995 (N_18995,N_18730,N_18769);
or U18996 (N_18996,N_18823,N_18786);
nand U18997 (N_18997,N_18836,N_18864);
or U18998 (N_18998,N_18824,N_18760);
nand U18999 (N_18999,N_18758,N_18727);
and U19000 (N_19000,N_18798,N_18878);
or U19001 (N_19001,N_18848,N_18823);
nand U19002 (N_19002,N_18772,N_18793);
or U19003 (N_19003,N_18769,N_18767);
or U19004 (N_19004,N_18860,N_18734);
or U19005 (N_19005,N_18755,N_18827);
xnor U19006 (N_19006,N_18836,N_18875);
and U19007 (N_19007,N_18738,N_18838);
nand U19008 (N_19008,N_18852,N_18765);
or U19009 (N_19009,N_18833,N_18737);
xor U19010 (N_19010,N_18733,N_18776);
nand U19011 (N_19011,N_18832,N_18837);
nor U19012 (N_19012,N_18786,N_18868);
or U19013 (N_19013,N_18795,N_18861);
or U19014 (N_19014,N_18803,N_18743);
nor U19015 (N_19015,N_18745,N_18772);
nor U19016 (N_19016,N_18825,N_18737);
or U19017 (N_19017,N_18736,N_18872);
and U19018 (N_19018,N_18729,N_18805);
or U19019 (N_19019,N_18811,N_18864);
xor U19020 (N_19020,N_18828,N_18750);
or U19021 (N_19021,N_18831,N_18857);
nor U19022 (N_19022,N_18770,N_18791);
and U19023 (N_19023,N_18732,N_18788);
xor U19024 (N_19024,N_18838,N_18756);
nand U19025 (N_19025,N_18809,N_18829);
or U19026 (N_19026,N_18775,N_18850);
and U19027 (N_19027,N_18801,N_18867);
nand U19028 (N_19028,N_18841,N_18741);
nand U19029 (N_19029,N_18794,N_18733);
xor U19030 (N_19030,N_18800,N_18855);
or U19031 (N_19031,N_18733,N_18721);
or U19032 (N_19032,N_18739,N_18724);
or U19033 (N_19033,N_18769,N_18847);
xnor U19034 (N_19034,N_18800,N_18856);
nand U19035 (N_19035,N_18864,N_18857);
nand U19036 (N_19036,N_18797,N_18745);
nor U19037 (N_19037,N_18825,N_18855);
and U19038 (N_19038,N_18744,N_18830);
and U19039 (N_19039,N_18789,N_18813);
or U19040 (N_19040,N_18903,N_19028);
nor U19041 (N_19041,N_19012,N_18999);
or U19042 (N_19042,N_18936,N_18950);
or U19043 (N_19043,N_18947,N_18937);
or U19044 (N_19044,N_19017,N_18891);
xor U19045 (N_19045,N_18945,N_19011);
nand U19046 (N_19046,N_18926,N_18888);
or U19047 (N_19047,N_19019,N_18884);
and U19048 (N_19048,N_19031,N_18940);
nor U19049 (N_19049,N_18939,N_19002);
or U19050 (N_19050,N_18922,N_18996);
xor U19051 (N_19051,N_18928,N_19023);
xor U19052 (N_19052,N_18898,N_18918);
nor U19053 (N_19053,N_18907,N_18904);
nor U19054 (N_19054,N_18887,N_18913);
and U19055 (N_19055,N_19029,N_18911);
xor U19056 (N_19056,N_19010,N_19009);
nand U19057 (N_19057,N_18932,N_18896);
and U19058 (N_19058,N_18890,N_18984);
nor U19059 (N_19059,N_18925,N_19007);
xor U19060 (N_19060,N_18997,N_18982);
and U19061 (N_19061,N_18920,N_18986);
nor U19062 (N_19062,N_19021,N_19036);
nand U19063 (N_19063,N_18948,N_18927);
nor U19064 (N_19064,N_18953,N_18916);
nor U19065 (N_19065,N_18961,N_18992);
nor U19066 (N_19066,N_18895,N_19001);
nor U19067 (N_19067,N_18956,N_18991);
or U19068 (N_19068,N_19038,N_18931);
nor U19069 (N_19069,N_19015,N_18995);
and U19070 (N_19070,N_18883,N_18899);
nand U19071 (N_19071,N_18942,N_19016);
nor U19072 (N_19072,N_19014,N_19022);
nor U19073 (N_19073,N_18975,N_18981);
nor U19074 (N_19074,N_18957,N_18966);
nand U19075 (N_19075,N_18944,N_19018);
and U19076 (N_19076,N_18909,N_19020);
and U19077 (N_19077,N_18952,N_18990);
or U19078 (N_19078,N_18974,N_18880);
xor U19079 (N_19079,N_18973,N_19006);
or U19080 (N_19080,N_18954,N_19035);
or U19081 (N_19081,N_18900,N_18933);
and U19082 (N_19082,N_19037,N_18959);
nand U19083 (N_19083,N_18946,N_19026);
xor U19084 (N_19084,N_18980,N_18958);
and U19085 (N_19085,N_18960,N_18912);
or U19086 (N_19086,N_18977,N_18979);
or U19087 (N_19087,N_19013,N_19025);
nor U19088 (N_19088,N_18972,N_18915);
or U19089 (N_19089,N_18923,N_18988);
nand U19090 (N_19090,N_18894,N_19024);
or U19091 (N_19091,N_18941,N_18910);
and U19092 (N_19092,N_19039,N_18985);
and U19093 (N_19093,N_18967,N_18987);
xnor U19094 (N_19094,N_18906,N_18978);
nand U19095 (N_19095,N_18897,N_18921);
and U19096 (N_19096,N_19000,N_18892);
or U19097 (N_19097,N_18914,N_18905);
or U19098 (N_19098,N_18938,N_18919);
nand U19099 (N_19099,N_18970,N_18889);
or U19100 (N_19100,N_18969,N_18963);
nor U19101 (N_19101,N_18908,N_18930);
nor U19102 (N_19102,N_18934,N_18924);
nor U19103 (N_19103,N_18951,N_18943);
or U19104 (N_19104,N_19008,N_18929);
nor U19105 (N_19105,N_19034,N_18971);
or U19106 (N_19106,N_18998,N_18965);
nand U19107 (N_19107,N_18886,N_19027);
or U19108 (N_19108,N_18881,N_19030);
xor U19109 (N_19109,N_18882,N_18955);
xnor U19110 (N_19110,N_18993,N_19005);
nor U19111 (N_19111,N_18983,N_18935);
or U19112 (N_19112,N_18962,N_18917);
and U19113 (N_19113,N_19032,N_19004);
xnor U19114 (N_19114,N_19003,N_18976);
nand U19115 (N_19115,N_18994,N_18968);
and U19116 (N_19116,N_18949,N_18964);
nand U19117 (N_19117,N_18901,N_18885);
nand U19118 (N_19118,N_18893,N_19033);
or U19119 (N_19119,N_18902,N_18989);
nor U19120 (N_19120,N_18895,N_18993);
or U19121 (N_19121,N_18992,N_19010);
nand U19122 (N_19122,N_19039,N_19016);
nor U19123 (N_19123,N_19033,N_19002);
nand U19124 (N_19124,N_19032,N_19035);
nand U19125 (N_19125,N_18884,N_18936);
xnor U19126 (N_19126,N_18962,N_18933);
or U19127 (N_19127,N_19009,N_18934);
xnor U19128 (N_19128,N_18940,N_18907);
nand U19129 (N_19129,N_19015,N_18975);
or U19130 (N_19130,N_19003,N_18895);
xnor U19131 (N_19131,N_18992,N_19038);
and U19132 (N_19132,N_18980,N_18994);
xor U19133 (N_19133,N_18886,N_18959);
and U19134 (N_19134,N_18949,N_18928);
or U19135 (N_19135,N_18932,N_18938);
nand U19136 (N_19136,N_18901,N_18960);
xnor U19137 (N_19137,N_18973,N_18934);
xnor U19138 (N_19138,N_18973,N_18985);
nand U19139 (N_19139,N_18936,N_18932);
or U19140 (N_19140,N_18938,N_18964);
nor U19141 (N_19141,N_18920,N_18951);
xor U19142 (N_19142,N_18926,N_18986);
and U19143 (N_19143,N_19004,N_18941);
nor U19144 (N_19144,N_18975,N_18961);
xor U19145 (N_19145,N_18919,N_18937);
nand U19146 (N_19146,N_19024,N_18918);
and U19147 (N_19147,N_18890,N_19021);
nand U19148 (N_19148,N_18895,N_18967);
nor U19149 (N_19149,N_18989,N_18903);
or U19150 (N_19150,N_18907,N_19024);
and U19151 (N_19151,N_18968,N_18950);
nor U19152 (N_19152,N_19015,N_18991);
nor U19153 (N_19153,N_19023,N_18950);
and U19154 (N_19154,N_18993,N_18964);
xnor U19155 (N_19155,N_18885,N_19034);
nand U19156 (N_19156,N_19015,N_18912);
nor U19157 (N_19157,N_18955,N_19038);
nand U19158 (N_19158,N_18891,N_18881);
xor U19159 (N_19159,N_18953,N_18989);
nor U19160 (N_19160,N_18937,N_18948);
or U19161 (N_19161,N_18955,N_19028);
nor U19162 (N_19162,N_18944,N_19039);
and U19163 (N_19163,N_18940,N_18962);
nand U19164 (N_19164,N_18889,N_18908);
nand U19165 (N_19165,N_19003,N_19013);
nor U19166 (N_19166,N_18905,N_18951);
nor U19167 (N_19167,N_19029,N_18994);
and U19168 (N_19168,N_18911,N_19021);
and U19169 (N_19169,N_18939,N_19019);
xnor U19170 (N_19170,N_19038,N_19037);
nand U19171 (N_19171,N_19009,N_19005);
nor U19172 (N_19172,N_18958,N_19028);
xnor U19173 (N_19173,N_18881,N_18977);
nor U19174 (N_19174,N_18966,N_18975);
or U19175 (N_19175,N_18973,N_18990);
nor U19176 (N_19176,N_18965,N_18918);
xor U19177 (N_19177,N_18924,N_18981);
xor U19178 (N_19178,N_19017,N_18913);
nor U19179 (N_19179,N_18928,N_18995);
and U19180 (N_19180,N_18882,N_18959);
or U19181 (N_19181,N_18946,N_18933);
nand U19182 (N_19182,N_18955,N_18970);
or U19183 (N_19183,N_19019,N_18914);
or U19184 (N_19184,N_18954,N_18991);
and U19185 (N_19185,N_18938,N_19011);
nand U19186 (N_19186,N_18918,N_19029);
or U19187 (N_19187,N_18991,N_19000);
nand U19188 (N_19188,N_18951,N_19004);
and U19189 (N_19189,N_18900,N_18999);
and U19190 (N_19190,N_18982,N_19000);
and U19191 (N_19191,N_19016,N_18986);
or U19192 (N_19192,N_19010,N_19000);
nor U19193 (N_19193,N_18912,N_18918);
or U19194 (N_19194,N_19027,N_18984);
and U19195 (N_19195,N_18996,N_18910);
nand U19196 (N_19196,N_18985,N_18967);
nand U19197 (N_19197,N_19036,N_18961);
xor U19198 (N_19198,N_18958,N_18882);
and U19199 (N_19199,N_19033,N_18902);
and U19200 (N_19200,N_19065,N_19162);
xor U19201 (N_19201,N_19056,N_19125);
nor U19202 (N_19202,N_19053,N_19186);
xor U19203 (N_19203,N_19176,N_19054);
nor U19204 (N_19204,N_19120,N_19190);
xnor U19205 (N_19205,N_19100,N_19115);
xor U19206 (N_19206,N_19075,N_19091);
nand U19207 (N_19207,N_19134,N_19069);
nor U19208 (N_19208,N_19127,N_19129);
xnor U19209 (N_19209,N_19042,N_19068);
xor U19210 (N_19210,N_19083,N_19148);
and U19211 (N_19211,N_19116,N_19102);
xnor U19212 (N_19212,N_19169,N_19079);
nor U19213 (N_19213,N_19078,N_19181);
or U19214 (N_19214,N_19117,N_19135);
nand U19215 (N_19215,N_19050,N_19090);
xor U19216 (N_19216,N_19055,N_19092);
and U19217 (N_19217,N_19097,N_19199);
xor U19218 (N_19218,N_19122,N_19153);
nor U19219 (N_19219,N_19142,N_19177);
nand U19220 (N_19220,N_19141,N_19057);
or U19221 (N_19221,N_19151,N_19157);
nor U19222 (N_19222,N_19094,N_19043);
and U19223 (N_19223,N_19072,N_19046);
and U19224 (N_19224,N_19154,N_19052);
nor U19225 (N_19225,N_19156,N_19145);
or U19226 (N_19226,N_19171,N_19098);
or U19227 (N_19227,N_19185,N_19193);
nand U19228 (N_19228,N_19168,N_19073);
nor U19229 (N_19229,N_19191,N_19150);
nor U19230 (N_19230,N_19066,N_19089);
nor U19231 (N_19231,N_19084,N_19188);
or U19232 (N_19232,N_19062,N_19107);
nand U19233 (N_19233,N_19184,N_19058);
nor U19234 (N_19234,N_19165,N_19070);
xnor U19235 (N_19235,N_19197,N_19194);
and U19236 (N_19236,N_19159,N_19067);
nand U19237 (N_19237,N_19140,N_19076);
xor U19238 (N_19238,N_19133,N_19045);
or U19239 (N_19239,N_19187,N_19174);
nand U19240 (N_19240,N_19110,N_19167);
nor U19241 (N_19241,N_19048,N_19096);
nand U19242 (N_19242,N_19059,N_19155);
and U19243 (N_19243,N_19082,N_19114);
xnor U19244 (N_19244,N_19121,N_19189);
nand U19245 (N_19245,N_19182,N_19086);
nand U19246 (N_19246,N_19195,N_19138);
xor U19247 (N_19247,N_19152,N_19160);
xnor U19248 (N_19248,N_19198,N_19063);
nor U19249 (N_19249,N_19074,N_19161);
nor U19250 (N_19250,N_19183,N_19108);
and U19251 (N_19251,N_19132,N_19049);
xnor U19252 (N_19252,N_19128,N_19080);
nand U19253 (N_19253,N_19131,N_19166);
xor U19254 (N_19254,N_19103,N_19137);
or U19255 (N_19255,N_19163,N_19087);
and U19256 (N_19256,N_19064,N_19158);
nor U19257 (N_19257,N_19040,N_19101);
xor U19258 (N_19258,N_19088,N_19144);
or U19259 (N_19259,N_19060,N_19196);
and U19260 (N_19260,N_19077,N_19170);
xnor U19261 (N_19261,N_19051,N_19093);
nor U19262 (N_19262,N_19081,N_19041);
nor U19263 (N_19263,N_19095,N_19139);
nor U19264 (N_19264,N_19130,N_19146);
or U19265 (N_19265,N_19147,N_19047);
and U19266 (N_19266,N_19179,N_19123);
and U19267 (N_19267,N_19112,N_19180);
nor U19268 (N_19268,N_19105,N_19119);
xnor U19269 (N_19269,N_19085,N_19164);
xor U19270 (N_19270,N_19149,N_19126);
nand U19271 (N_19271,N_19118,N_19106);
or U19272 (N_19272,N_19178,N_19173);
nor U19273 (N_19273,N_19172,N_19044);
and U19274 (N_19274,N_19192,N_19175);
or U19275 (N_19275,N_19124,N_19071);
nand U19276 (N_19276,N_19113,N_19109);
xnor U19277 (N_19277,N_19099,N_19111);
and U19278 (N_19278,N_19104,N_19143);
or U19279 (N_19279,N_19061,N_19136);
nor U19280 (N_19280,N_19171,N_19115);
and U19281 (N_19281,N_19188,N_19040);
nor U19282 (N_19282,N_19173,N_19042);
xnor U19283 (N_19283,N_19077,N_19106);
or U19284 (N_19284,N_19086,N_19045);
and U19285 (N_19285,N_19122,N_19059);
or U19286 (N_19286,N_19169,N_19145);
nand U19287 (N_19287,N_19088,N_19128);
xor U19288 (N_19288,N_19143,N_19073);
or U19289 (N_19289,N_19118,N_19099);
nand U19290 (N_19290,N_19150,N_19119);
nand U19291 (N_19291,N_19160,N_19099);
or U19292 (N_19292,N_19129,N_19101);
nand U19293 (N_19293,N_19086,N_19056);
nand U19294 (N_19294,N_19130,N_19138);
nand U19295 (N_19295,N_19114,N_19141);
nand U19296 (N_19296,N_19068,N_19085);
xor U19297 (N_19297,N_19103,N_19098);
xor U19298 (N_19298,N_19057,N_19101);
xnor U19299 (N_19299,N_19126,N_19063);
nor U19300 (N_19300,N_19041,N_19061);
xnor U19301 (N_19301,N_19180,N_19077);
or U19302 (N_19302,N_19103,N_19191);
and U19303 (N_19303,N_19091,N_19181);
or U19304 (N_19304,N_19082,N_19051);
nor U19305 (N_19305,N_19041,N_19111);
nand U19306 (N_19306,N_19090,N_19140);
nand U19307 (N_19307,N_19181,N_19074);
nand U19308 (N_19308,N_19063,N_19111);
or U19309 (N_19309,N_19144,N_19178);
nor U19310 (N_19310,N_19131,N_19084);
xnor U19311 (N_19311,N_19164,N_19130);
or U19312 (N_19312,N_19113,N_19125);
or U19313 (N_19313,N_19182,N_19130);
nand U19314 (N_19314,N_19058,N_19193);
or U19315 (N_19315,N_19102,N_19155);
and U19316 (N_19316,N_19106,N_19111);
xnor U19317 (N_19317,N_19121,N_19166);
xor U19318 (N_19318,N_19112,N_19052);
or U19319 (N_19319,N_19072,N_19162);
nor U19320 (N_19320,N_19083,N_19197);
nand U19321 (N_19321,N_19118,N_19083);
or U19322 (N_19322,N_19071,N_19079);
nor U19323 (N_19323,N_19113,N_19092);
nand U19324 (N_19324,N_19084,N_19071);
or U19325 (N_19325,N_19190,N_19090);
and U19326 (N_19326,N_19174,N_19100);
xor U19327 (N_19327,N_19182,N_19123);
nor U19328 (N_19328,N_19109,N_19044);
xnor U19329 (N_19329,N_19154,N_19171);
and U19330 (N_19330,N_19092,N_19148);
or U19331 (N_19331,N_19080,N_19168);
and U19332 (N_19332,N_19136,N_19187);
nand U19333 (N_19333,N_19122,N_19041);
and U19334 (N_19334,N_19125,N_19076);
xor U19335 (N_19335,N_19187,N_19181);
nor U19336 (N_19336,N_19158,N_19193);
and U19337 (N_19337,N_19138,N_19186);
nand U19338 (N_19338,N_19080,N_19159);
nor U19339 (N_19339,N_19136,N_19124);
nand U19340 (N_19340,N_19157,N_19111);
nor U19341 (N_19341,N_19142,N_19041);
or U19342 (N_19342,N_19125,N_19116);
xnor U19343 (N_19343,N_19146,N_19089);
xor U19344 (N_19344,N_19191,N_19196);
or U19345 (N_19345,N_19179,N_19055);
and U19346 (N_19346,N_19144,N_19191);
nand U19347 (N_19347,N_19164,N_19077);
nor U19348 (N_19348,N_19100,N_19097);
xnor U19349 (N_19349,N_19053,N_19140);
and U19350 (N_19350,N_19079,N_19181);
xor U19351 (N_19351,N_19046,N_19182);
nor U19352 (N_19352,N_19150,N_19154);
xor U19353 (N_19353,N_19067,N_19041);
nor U19354 (N_19354,N_19196,N_19048);
or U19355 (N_19355,N_19168,N_19127);
nor U19356 (N_19356,N_19113,N_19066);
xnor U19357 (N_19357,N_19182,N_19127);
or U19358 (N_19358,N_19047,N_19157);
and U19359 (N_19359,N_19128,N_19056);
and U19360 (N_19360,N_19291,N_19340);
nor U19361 (N_19361,N_19255,N_19276);
xnor U19362 (N_19362,N_19308,N_19279);
or U19363 (N_19363,N_19320,N_19299);
nand U19364 (N_19364,N_19203,N_19201);
nand U19365 (N_19365,N_19322,N_19286);
nor U19366 (N_19366,N_19212,N_19327);
nand U19367 (N_19367,N_19244,N_19314);
and U19368 (N_19368,N_19355,N_19293);
nor U19369 (N_19369,N_19310,N_19338);
xnor U19370 (N_19370,N_19281,N_19270);
and U19371 (N_19371,N_19218,N_19211);
nor U19372 (N_19372,N_19278,N_19348);
nor U19373 (N_19373,N_19221,N_19311);
xnor U19374 (N_19374,N_19336,N_19215);
and U19375 (N_19375,N_19325,N_19300);
nand U19376 (N_19376,N_19248,N_19251);
and U19377 (N_19377,N_19263,N_19238);
nor U19378 (N_19378,N_19297,N_19344);
nor U19379 (N_19379,N_19219,N_19341);
nand U19380 (N_19380,N_19358,N_19245);
xor U19381 (N_19381,N_19249,N_19240);
xnor U19382 (N_19382,N_19326,N_19312);
xnor U19383 (N_19383,N_19342,N_19275);
and U19384 (N_19384,N_19273,N_19306);
nor U19385 (N_19385,N_19284,N_19224);
nand U19386 (N_19386,N_19239,N_19282);
nand U19387 (N_19387,N_19202,N_19307);
and U19388 (N_19388,N_19304,N_19264);
and U19389 (N_19389,N_19208,N_19288);
nand U19390 (N_19390,N_19330,N_19222);
nand U19391 (N_19391,N_19334,N_19315);
xor U19392 (N_19392,N_19209,N_19345);
nor U19393 (N_19393,N_19349,N_19228);
and U19394 (N_19394,N_19247,N_19277);
nor U19395 (N_19395,N_19357,N_19231);
or U19396 (N_19396,N_19259,N_19335);
xnor U19397 (N_19397,N_19226,N_19285);
nor U19398 (N_19398,N_19242,N_19298);
nand U19399 (N_19399,N_19289,N_19271);
or U19400 (N_19400,N_19260,N_19214);
nand U19401 (N_19401,N_19354,N_19294);
xnor U19402 (N_19402,N_19235,N_19267);
nor U19403 (N_19403,N_19266,N_19351);
xor U19404 (N_19404,N_19257,N_19236);
xor U19405 (N_19405,N_19352,N_19232);
xor U19406 (N_19406,N_19204,N_19230);
or U19407 (N_19407,N_19350,N_19225);
xor U19408 (N_19408,N_19272,N_19343);
or U19409 (N_19409,N_19261,N_19265);
or U19410 (N_19410,N_19254,N_19296);
or U19411 (N_19411,N_19280,N_19233);
and U19412 (N_19412,N_19313,N_19292);
and U19413 (N_19413,N_19353,N_19347);
nor U19414 (N_19414,N_19234,N_19333);
and U19415 (N_19415,N_19256,N_19205);
nand U19416 (N_19416,N_19303,N_19305);
nor U19417 (N_19417,N_19274,N_19268);
nor U19418 (N_19418,N_19316,N_19241);
nand U19419 (N_19419,N_19252,N_19302);
xnor U19420 (N_19420,N_19287,N_19283);
nor U19421 (N_19421,N_19328,N_19210);
or U19422 (N_19422,N_19206,N_19290);
or U19423 (N_19423,N_19217,N_19359);
nand U19424 (N_19424,N_19213,N_19246);
nand U19425 (N_19425,N_19321,N_19346);
nand U19426 (N_19426,N_19258,N_19207);
xnor U19427 (N_19427,N_19323,N_19220);
xor U19428 (N_19428,N_19309,N_19216);
nor U19429 (N_19429,N_19301,N_19262);
nor U19430 (N_19430,N_19269,N_19253);
or U19431 (N_19431,N_19243,N_19356);
nor U19432 (N_19432,N_19237,N_19223);
or U19433 (N_19433,N_19329,N_19324);
and U19434 (N_19434,N_19332,N_19331);
or U19435 (N_19435,N_19295,N_19337);
xor U19436 (N_19436,N_19317,N_19339);
nor U19437 (N_19437,N_19200,N_19318);
and U19438 (N_19438,N_19319,N_19227);
xnor U19439 (N_19439,N_19229,N_19250);
nor U19440 (N_19440,N_19200,N_19277);
xor U19441 (N_19441,N_19343,N_19256);
and U19442 (N_19442,N_19262,N_19208);
or U19443 (N_19443,N_19351,N_19239);
and U19444 (N_19444,N_19309,N_19300);
and U19445 (N_19445,N_19262,N_19291);
nor U19446 (N_19446,N_19346,N_19254);
or U19447 (N_19447,N_19258,N_19222);
nand U19448 (N_19448,N_19342,N_19326);
nand U19449 (N_19449,N_19318,N_19358);
or U19450 (N_19450,N_19257,N_19229);
nand U19451 (N_19451,N_19281,N_19217);
xnor U19452 (N_19452,N_19315,N_19278);
or U19453 (N_19453,N_19211,N_19322);
nand U19454 (N_19454,N_19348,N_19310);
and U19455 (N_19455,N_19310,N_19236);
and U19456 (N_19456,N_19213,N_19317);
nand U19457 (N_19457,N_19247,N_19213);
and U19458 (N_19458,N_19210,N_19305);
nand U19459 (N_19459,N_19353,N_19309);
or U19460 (N_19460,N_19343,N_19216);
nor U19461 (N_19461,N_19328,N_19330);
or U19462 (N_19462,N_19296,N_19288);
and U19463 (N_19463,N_19256,N_19222);
nor U19464 (N_19464,N_19268,N_19249);
xnor U19465 (N_19465,N_19217,N_19307);
or U19466 (N_19466,N_19226,N_19296);
or U19467 (N_19467,N_19283,N_19215);
nor U19468 (N_19468,N_19353,N_19214);
or U19469 (N_19469,N_19333,N_19277);
xor U19470 (N_19470,N_19298,N_19295);
or U19471 (N_19471,N_19326,N_19296);
and U19472 (N_19472,N_19261,N_19254);
and U19473 (N_19473,N_19342,N_19306);
nand U19474 (N_19474,N_19258,N_19241);
xor U19475 (N_19475,N_19243,N_19230);
nand U19476 (N_19476,N_19284,N_19342);
nor U19477 (N_19477,N_19247,N_19348);
and U19478 (N_19478,N_19287,N_19254);
and U19479 (N_19479,N_19307,N_19336);
or U19480 (N_19480,N_19298,N_19286);
or U19481 (N_19481,N_19246,N_19277);
xor U19482 (N_19482,N_19270,N_19222);
nor U19483 (N_19483,N_19266,N_19318);
and U19484 (N_19484,N_19266,N_19206);
nand U19485 (N_19485,N_19331,N_19245);
or U19486 (N_19486,N_19356,N_19229);
or U19487 (N_19487,N_19331,N_19251);
and U19488 (N_19488,N_19273,N_19308);
nor U19489 (N_19489,N_19206,N_19326);
nand U19490 (N_19490,N_19253,N_19219);
or U19491 (N_19491,N_19312,N_19330);
xnor U19492 (N_19492,N_19316,N_19324);
xor U19493 (N_19493,N_19352,N_19226);
or U19494 (N_19494,N_19269,N_19205);
xnor U19495 (N_19495,N_19217,N_19336);
xnor U19496 (N_19496,N_19317,N_19233);
nand U19497 (N_19497,N_19355,N_19269);
or U19498 (N_19498,N_19222,N_19232);
xnor U19499 (N_19499,N_19214,N_19299);
or U19500 (N_19500,N_19225,N_19245);
nor U19501 (N_19501,N_19285,N_19201);
or U19502 (N_19502,N_19328,N_19284);
nand U19503 (N_19503,N_19241,N_19278);
and U19504 (N_19504,N_19276,N_19283);
xnor U19505 (N_19505,N_19247,N_19218);
xor U19506 (N_19506,N_19359,N_19226);
nor U19507 (N_19507,N_19267,N_19250);
nand U19508 (N_19508,N_19273,N_19305);
nand U19509 (N_19509,N_19321,N_19283);
and U19510 (N_19510,N_19213,N_19270);
xnor U19511 (N_19511,N_19254,N_19251);
nand U19512 (N_19512,N_19306,N_19270);
or U19513 (N_19513,N_19312,N_19254);
and U19514 (N_19514,N_19315,N_19289);
xnor U19515 (N_19515,N_19207,N_19253);
nand U19516 (N_19516,N_19242,N_19349);
and U19517 (N_19517,N_19325,N_19270);
or U19518 (N_19518,N_19277,N_19233);
xor U19519 (N_19519,N_19337,N_19304);
nand U19520 (N_19520,N_19412,N_19366);
and U19521 (N_19521,N_19463,N_19411);
nand U19522 (N_19522,N_19444,N_19371);
nor U19523 (N_19523,N_19380,N_19399);
nor U19524 (N_19524,N_19458,N_19374);
nor U19525 (N_19525,N_19367,N_19391);
nand U19526 (N_19526,N_19510,N_19402);
xor U19527 (N_19527,N_19477,N_19373);
or U19528 (N_19528,N_19509,N_19483);
xnor U19529 (N_19529,N_19423,N_19401);
nor U19530 (N_19530,N_19454,N_19487);
xor U19531 (N_19531,N_19514,N_19396);
nand U19532 (N_19532,N_19434,N_19460);
nand U19533 (N_19533,N_19448,N_19453);
and U19534 (N_19534,N_19498,N_19455);
nand U19535 (N_19535,N_19485,N_19465);
nand U19536 (N_19536,N_19497,N_19507);
or U19537 (N_19537,N_19408,N_19431);
and U19538 (N_19538,N_19429,N_19418);
nand U19539 (N_19539,N_19386,N_19388);
or U19540 (N_19540,N_19512,N_19414);
nand U19541 (N_19541,N_19370,N_19364);
nand U19542 (N_19542,N_19390,N_19471);
and U19543 (N_19543,N_19372,N_19449);
xnor U19544 (N_19544,N_19428,N_19383);
nor U19545 (N_19545,N_19504,N_19486);
or U19546 (N_19546,N_19457,N_19519);
or U19547 (N_19547,N_19500,N_19502);
nand U19548 (N_19548,N_19480,N_19369);
nand U19549 (N_19549,N_19459,N_19495);
xnor U19550 (N_19550,N_19432,N_19415);
nand U19551 (N_19551,N_19387,N_19475);
nand U19552 (N_19552,N_19476,N_19389);
nand U19553 (N_19553,N_19397,N_19445);
and U19554 (N_19554,N_19461,N_19464);
xnor U19555 (N_19555,N_19481,N_19403);
xnor U19556 (N_19556,N_19368,N_19472);
or U19557 (N_19557,N_19469,N_19484);
xnor U19558 (N_19558,N_19468,N_19362);
nand U19559 (N_19559,N_19377,N_19407);
nor U19560 (N_19560,N_19451,N_19513);
or U19561 (N_19561,N_19490,N_19443);
nor U19562 (N_19562,N_19473,N_19511);
nor U19563 (N_19563,N_19382,N_19491);
nand U19564 (N_19564,N_19506,N_19442);
and U19565 (N_19565,N_19398,N_19438);
or U19566 (N_19566,N_19406,N_19503);
nand U19567 (N_19567,N_19478,N_19517);
and U19568 (N_19568,N_19375,N_19422);
or U19569 (N_19569,N_19400,N_19409);
and U19570 (N_19570,N_19405,N_19395);
nand U19571 (N_19571,N_19426,N_19518);
xnor U19572 (N_19572,N_19505,N_19479);
or U19573 (N_19573,N_19466,N_19441);
xor U19574 (N_19574,N_19413,N_19493);
xor U19575 (N_19575,N_19456,N_19376);
or U19576 (N_19576,N_19416,N_19420);
nand U19577 (N_19577,N_19430,N_19437);
nand U19578 (N_19578,N_19393,N_19433);
nor U19579 (N_19579,N_19381,N_19379);
and U19580 (N_19580,N_19492,N_19392);
nor U19581 (N_19581,N_19446,N_19361);
nand U19582 (N_19582,N_19516,N_19499);
or U19583 (N_19583,N_19436,N_19450);
or U19584 (N_19584,N_19427,N_19470);
or U19585 (N_19585,N_19496,N_19482);
and U19586 (N_19586,N_19501,N_19421);
and U19587 (N_19587,N_19439,N_19378);
nor U19588 (N_19588,N_19488,N_19365);
xor U19589 (N_19589,N_19410,N_19417);
nor U19590 (N_19590,N_19363,N_19515);
xnor U19591 (N_19591,N_19462,N_19394);
nand U19592 (N_19592,N_19404,N_19384);
nor U19593 (N_19593,N_19474,N_19447);
nand U19594 (N_19594,N_19425,N_19435);
nand U19595 (N_19595,N_19467,N_19508);
nor U19596 (N_19596,N_19419,N_19494);
or U19597 (N_19597,N_19489,N_19452);
and U19598 (N_19598,N_19424,N_19440);
nor U19599 (N_19599,N_19385,N_19360);
nand U19600 (N_19600,N_19472,N_19403);
nand U19601 (N_19601,N_19503,N_19432);
and U19602 (N_19602,N_19497,N_19374);
nand U19603 (N_19603,N_19417,N_19512);
nand U19604 (N_19604,N_19417,N_19518);
nor U19605 (N_19605,N_19380,N_19467);
or U19606 (N_19606,N_19400,N_19441);
nand U19607 (N_19607,N_19377,N_19401);
or U19608 (N_19608,N_19476,N_19364);
nor U19609 (N_19609,N_19506,N_19361);
nor U19610 (N_19610,N_19409,N_19429);
nand U19611 (N_19611,N_19382,N_19383);
and U19612 (N_19612,N_19434,N_19452);
nor U19613 (N_19613,N_19425,N_19518);
or U19614 (N_19614,N_19510,N_19392);
or U19615 (N_19615,N_19457,N_19455);
and U19616 (N_19616,N_19475,N_19360);
or U19617 (N_19617,N_19410,N_19450);
xor U19618 (N_19618,N_19389,N_19478);
and U19619 (N_19619,N_19469,N_19444);
xnor U19620 (N_19620,N_19387,N_19458);
nor U19621 (N_19621,N_19505,N_19466);
nor U19622 (N_19622,N_19461,N_19391);
nand U19623 (N_19623,N_19368,N_19374);
or U19624 (N_19624,N_19485,N_19510);
or U19625 (N_19625,N_19403,N_19383);
and U19626 (N_19626,N_19399,N_19411);
xor U19627 (N_19627,N_19456,N_19439);
or U19628 (N_19628,N_19433,N_19449);
or U19629 (N_19629,N_19384,N_19381);
and U19630 (N_19630,N_19489,N_19450);
and U19631 (N_19631,N_19506,N_19517);
nand U19632 (N_19632,N_19484,N_19414);
nor U19633 (N_19633,N_19489,N_19384);
nor U19634 (N_19634,N_19512,N_19514);
nand U19635 (N_19635,N_19453,N_19443);
and U19636 (N_19636,N_19473,N_19461);
and U19637 (N_19637,N_19432,N_19388);
and U19638 (N_19638,N_19393,N_19465);
nand U19639 (N_19639,N_19387,N_19373);
xnor U19640 (N_19640,N_19488,N_19468);
xnor U19641 (N_19641,N_19418,N_19365);
and U19642 (N_19642,N_19489,N_19480);
nor U19643 (N_19643,N_19422,N_19518);
nand U19644 (N_19644,N_19438,N_19373);
xnor U19645 (N_19645,N_19423,N_19453);
and U19646 (N_19646,N_19379,N_19518);
or U19647 (N_19647,N_19422,N_19453);
or U19648 (N_19648,N_19412,N_19384);
and U19649 (N_19649,N_19471,N_19407);
and U19650 (N_19650,N_19463,N_19364);
xnor U19651 (N_19651,N_19423,N_19511);
or U19652 (N_19652,N_19513,N_19420);
xnor U19653 (N_19653,N_19502,N_19406);
xnor U19654 (N_19654,N_19460,N_19506);
nor U19655 (N_19655,N_19518,N_19519);
nor U19656 (N_19656,N_19498,N_19489);
or U19657 (N_19657,N_19483,N_19513);
nand U19658 (N_19658,N_19455,N_19393);
nand U19659 (N_19659,N_19509,N_19421);
nor U19660 (N_19660,N_19424,N_19438);
and U19661 (N_19661,N_19361,N_19428);
or U19662 (N_19662,N_19377,N_19418);
xor U19663 (N_19663,N_19403,N_19438);
nor U19664 (N_19664,N_19471,N_19473);
nand U19665 (N_19665,N_19455,N_19492);
or U19666 (N_19666,N_19368,N_19422);
or U19667 (N_19667,N_19465,N_19427);
xor U19668 (N_19668,N_19517,N_19510);
xor U19669 (N_19669,N_19510,N_19426);
and U19670 (N_19670,N_19406,N_19374);
or U19671 (N_19671,N_19389,N_19390);
nor U19672 (N_19672,N_19391,N_19502);
nor U19673 (N_19673,N_19488,N_19441);
nand U19674 (N_19674,N_19374,N_19443);
xor U19675 (N_19675,N_19425,N_19460);
nand U19676 (N_19676,N_19380,N_19441);
or U19677 (N_19677,N_19366,N_19495);
xnor U19678 (N_19678,N_19365,N_19448);
or U19679 (N_19679,N_19485,N_19498);
xor U19680 (N_19680,N_19526,N_19621);
nand U19681 (N_19681,N_19639,N_19675);
nand U19682 (N_19682,N_19566,N_19599);
and U19683 (N_19683,N_19570,N_19544);
and U19684 (N_19684,N_19541,N_19539);
and U19685 (N_19685,N_19583,N_19647);
or U19686 (N_19686,N_19576,N_19528);
and U19687 (N_19687,N_19565,N_19658);
and U19688 (N_19688,N_19637,N_19534);
xor U19689 (N_19689,N_19582,N_19630);
nand U19690 (N_19690,N_19578,N_19663);
xor U19691 (N_19691,N_19659,N_19626);
nand U19692 (N_19692,N_19623,N_19657);
and U19693 (N_19693,N_19610,N_19633);
nor U19694 (N_19694,N_19646,N_19627);
and U19695 (N_19695,N_19574,N_19554);
or U19696 (N_19696,N_19533,N_19521);
xnor U19697 (N_19697,N_19653,N_19605);
and U19698 (N_19698,N_19677,N_19664);
or U19699 (N_19699,N_19586,N_19560);
nand U19700 (N_19700,N_19580,N_19606);
xnor U19701 (N_19701,N_19593,N_19674);
or U19702 (N_19702,N_19649,N_19611);
xor U19703 (N_19703,N_19549,N_19558);
nor U19704 (N_19704,N_19613,N_19631);
nor U19705 (N_19705,N_19662,N_19625);
nor U19706 (N_19706,N_19601,N_19531);
xnor U19707 (N_19707,N_19594,N_19572);
xnor U19708 (N_19708,N_19543,N_19622);
nand U19709 (N_19709,N_19575,N_19660);
nor U19710 (N_19710,N_19588,N_19569);
nand U19711 (N_19711,N_19634,N_19648);
nor U19712 (N_19712,N_19562,N_19615);
nand U19713 (N_19713,N_19624,N_19671);
xnor U19714 (N_19714,N_19557,N_19589);
nor U19715 (N_19715,N_19596,N_19581);
nor U19716 (N_19716,N_19673,N_19654);
nand U19717 (N_19717,N_19587,N_19666);
or U19718 (N_19718,N_19670,N_19640);
and U19719 (N_19719,N_19603,N_19571);
nor U19720 (N_19720,N_19559,N_19669);
nand U19721 (N_19721,N_19592,N_19584);
and U19722 (N_19722,N_19656,N_19608);
nor U19723 (N_19723,N_19619,N_19598);
or U19724 (N_19724,N_19527,N_19661);
and U19725 (N_19725,N_19564,N_19609);
and U19726 (N_19726,N_19577,N_19600);
nor U19727 (N_19727,N_19641,N_19665);
or U19728 (N_19728,N_19530,N_19595);
nand U19729 (N_19729,N_19645,N_19536);
nand U19730 (N_19730,N_19524,N_19612);
nand U19731 (N_19731,N_19550,N_19602);
nor U19732 (N_19732,N_19607,N_19614);
and U19733 (N_19733,N_19538,N_19650);
or U19734 (N_19734,N_19546,N_19547);
or U19735 (N_19735,N_19667,N_19597);
or U19736 (N_19736,N_19542,N_19561);
and U19737 (N_19737,N_19563,N_19679);
nand U19738 (N_19738,N_19551,N_19556);
nor U19739 (N_19739,N_19590,N_19552);
nor U19740 (N_19740,N_19523,N_19629);
or U19741 (N_19741,N_19620,N_19652);
nor U19742 (N_19742,N_19616,N_19585);
and U19743 (N_19743,N_19522,N_19678);
and U19744 (N_19744,N_19591,N_19540);
nor U19745 (N_19745,N_19555,N_19579);
and U19746 (N_19746,N_19643,N_19553);
or U19747 (N_19747,N_19537,N_19635);
xnor U19748 (N_19748,N_19618,N_19655);
nor U19749 (N_19749,N_19617,N_19525);
nand U19750 (N_19750,N_19644,N_19628);
or U19751 (N_19751,N_19676,N_19636);
and U19752 (N_19752,N_19545,N_19548);
nand U19753 (N_19753,N_19535,N_19529);
xor U19754 (N_19754,N_19651,N_19638);
nor U19755 (N_19755,N_19632,N_19604);
or U19756 (N_19756,N_19642,N_19568);
and U19757 (N_19757,N_19520,N_19672);
and U19758 (N_19758,N_19532,N_19668);
or U19759 (N_19759,N_19573,N_19567);
nor U19760 (N_19760,N_19564,N_19644);
nor U19761 (N_19761,N_19557,N_19584);
and U19762 (N_19762,N_19595,N_19609);
xor U19763 (N_19763,N_19535,N_19664);
xnor U19764 (N_19764,N_19621,N_19603);
nand U19765 (N_19765,N_19643,N_19613);
nand U19766 (N_19766,N_19624,N_19657);
or U19767 (N_19767,N_19562,N_19539);
and U19768 (N_19768,N_19605,N_19520);
xnor U19769 (N_19769,N_19535,N_19545);
and U19770 (N_19770,N_19649,N_19529);
or U19771 (N_19771,N_19536,N_19668);
xnor U19772 (N_19772,N_19600,N_19634);
or U19773 (N_19773,N_19575,N_19541);
nand U19774 (N_19774,N_19563,N_19655);
nor U19775 (N_19775,N_19536,N_19540);
xnor U19776 (N_19776,N_19624,N_19549);
xnor U19777 (N_19777,N_19659,N_19618);
or U19778 (N_19778,N_19633,N_19555);
or U19779 (N_19779,N_19551,N_19537);
nor U19780 (N_19780,N_19677,N_19539);
nand U19781 (N_19781,N_19678,N_19667);
or U19782 (N_19782,N_19622,N_19613);
nor U19783 (N_19783,N_19627,N_19573);
and U19784 (N_19784,N_19557,N_19669);
nor U19785 (N_19785,N_19663,N_19653);
xnor U19786 (N_19786,N_19677,N_19553);
nand U19787 (N_19787,N_19557,N_19671);
or U19788 (N_19788,N_19544,N_19541);
and U19789 (N_19789,N_19661,N_19537);
or U19790 (N_19790,N_19550,N_19677);
nand U19791 (N_19791,N_19671,N_19617);
or U19792 (N_19792,N_19547,N_19591);
nand U19793 (N_19793,N_19561,N_19630);
nand U19794 (N_19794,N_19622,N_19589);
xor U19795 (N_19795,N_19636,N_19578);
nor U19796 (N_19796,N_19533,N_19662);
nand U19797 (N_19797,N_19583,N_19562);
or U19798 (N_19798,N_19651,N_19614);
nor U19799 (N_19799,N_19566,N_19653);
nand U19800 (N_19800,N_19646,N_19639);
nand U19801 (N_19801,N_19627,N_19578);
nor U19802 (N_19802,N_19602,N_19592);
or U19803 (N_19803,N_19593,N_19586);
nor U19804 (N_19804,N_19566,N_19632);
and U19805 (N_19805,N_19626,N_19663);
nor U19806 (N_19806,N_19527,N_19655);
nor U19807 (N_19807,N_19672,N_19549);
and U19808 (N_19808,N_19618,N_19558);
nand U19809 (N_19809,N_19536,N_19535);
nor U19810 (N_19810,N_19645,N_19642);
xor U19811 (N_19811,N_19605,N_19591);
nor U19812 (N_19812,N_19655,N_19522);
or U19813 (N_19813,N_19553,N_19661);
nor U19814 (N_19814,N_19588,N_19606);
xnor U19815 (N_19815,N_19672,N_19637);
nor U19816 (N_19816,N_19668,N_19647);
and U19817 (N_19817,N_19603,N_19641);
or U19818 (N_19818,N_19598,N_19588);
xor U19819 (N_19819,N_19612,N_19609);
nand U19820 (N_19820,N_19637,N_19589);
xnor U19821 (N_19821,N_19572,N_19604);
xor U19822 (N_19822,N_19582,N_19564);
and U19823 (N_19823,N_19621,N_19555);
or U19824 (N_19824,N_19679,N_19659);
and U19825 (N_19825,N_19585,N_19675);
and U19826 (N_19826,N_19546,N_19576);
or U19827 (N_19827,N_19531,N_19678);
and U19828 (N_19828,N_19577,N_19573);
nand U19829 (N_19829,N_19624,N_19604);
or U19830 (N_19830,N_19672,N_19595);
or U19831 (N_19831,N_19585,N_19562);
xor U19832 (N_19832,N_19615,N_19672);
xnor U19833 (N_19833,N_19654,N_19552);
nand U19834 (N_19834,N_19661,N_19641);
xor U19835 (N_19835,N_19672,N_19554);
xnor U19836 (N_19836,N_19582,N_19654);
and U19837 (N_19837,N_19592,N_19597);
nand U19838 (N_19838,N_19659,N_19646);
and U19839 (N_19839,N_19533,N_19631);
and U19840 (N_19840,N_19741,N_19792);
nor U19841 (N_19841,N_19683,N_19803);
nand U19842 (N_19842,N_19806,N_19812);
xnor U19843 (N_19843,N_19719,N_19698);
or U19844 (N_19844,N_19766,N_19770);
xor U19845 (N_19845,N_19691,N_19816);
xor U19846 (N_19846,N_19723,N_19747);
and U19847 (N_19847,N_19831,N_19810);
xnor U19848 (N_19848,N_19815,N_19687);
nand U19849 (N_19849,N_19715,N_19737);
xnor U19850 (N_19850,N_19830,N_19820);
or U19851 (N_19851,N_19799,N_19707);
nor U19852 (N_19852,N_19778,N_19724);
and U19853 (N_19853,N_19712,N_19813);
or U19854 (N_19854,N_19684,N_19811);
xor U19855 (N_19855,N_19727,N_19834);
nand U19856 (N_19856,N_19703,N_19739);
xor U19857 (N_19857,N_19755,N_19769);
nor U19858 (N_19858,N_19725,N_19756);
xor U19859 (N_19859,N_19818,N_19821);
xor U19860 (N_19860,N_19729,N_19751);
nand U19861 (N_19861,N_19711,N_19759);
xnor U19862 (N_19862,N_19686,N_19791);
or U19863 (N_19863,N_19718,N_19728);
nor U19864 (N_19864,N_19825,N_19768);
nor U19865 (N_19865,N_19828,N_19731);
and U19866 (N_19866,N_19693,N_19772);
nand U19867 (N_19867,N_19786,N_19829);
or U19868 (N_19868,N_19742,N_19823);
and U19869 (N_19869,N_19779,N_19798);
and U19870 (N_19870,N_19706,N_19743);
nor U19871 (N_19871,N_19814,N_19685);
xnor U19872 (N_19872,N_19688,N_19767);
nand U19873 (N_19873,N_19757,N_19682);
or U19874 (N_19874,N_19817,N_19714);
xor U19875 (N_19875,N_19762,N_19807);
and U19876 (N_19876,N_19796,N_19705);
and U19877 (N_19877,N_19783,N_19773);
nor U19878 (N_19878,N_19750,N_19819);
or U19879 (N_19879,N_19754,N_19732);
and U19880 (N_19880,N_19835,N_19735);
or U19881 (N_19881,N_19697,N_19805);
xnor U19882 (N_19882,N_19710,N_19744);
or U19883 (N_19883,N_19717,N_19726);
or U19884 (N_19884,N_19701,N_19826);
nand U19885 (N_19885,N_19716,N_19794);
nor U19886 (N_19886,N_19708,N_19837);
and U19887 (N_19887,N_19709,N_19838);
and U19888 (N_19888,N_19721,N_19681);
xnor U19889 (N_19889,N_19696,N_19782);
nand U19890 (N_19890,N_19801,N_19824);
or U19891 (N_19891,N_19775,N_19802);
or U19892 (N_19892,N_19809,N_19761);
or U19893 (N_19893,N_19694,N_19832);
or U19894 (N_19894,N_19800,N_19781);
nand U19895 (N_19895,N_19746,N_19692);
xor U19896 (N_19896,N_19804,N_19733);
xor U19897 (N_19897,N_19784,N_19839);
xor U19898 (N_19898,N_19787,N_19795);
and U19899 (N_19899,N_19699,N_19780);
nor U19900 (N_19900,N_19764,N_19680);
or U19901 (N_19901,N_19753,N_19827);
or U19902 (N_19902,N_19713,N_19695);
nand U19903 (N_19903,N_19752,N_19790);
xnor U19904 (N_19904,N_19771,N_19734);
xor U19905 (N_19905,N_19776,N_19785);
and U19906 (N_19906,N_19788,N_19748);
xnor U19907 (N_19907,N_19777,N_19690);
or U19908 (N_19908,N_19736,N_19760);
and U19909 (N_19909,N_19758,N_19740);
nand U19910 (N_19910,N_19833,N_19730);
nor U19911 (N_19911,N_19822,N_19774);
nor U19912 (N_19912,N_19749,N_19720);
xor U19913 (N_19913,N_19789,N_19797);
nand U19914 (N_19914,N_19722,N_19765);
nand U19915 (N_19915,N_19702,N_19808);
nand U19916 (N_19916,N_19793,N_19689);
nor U19917 (N_19917,N_19745,N_19738);
nand U19918 (N_19918,N_19836,N_19704);
nand U19919 (N_19919,N_19700,N_19763);
or U19920 (N_19920,N_19759,N_19729);
nand U19921 (N_19921,N_19735,N_19743);
nor U19922 (N_19922,N_19782,N_19797);
xor U19923 (N_19923,N_19823,N_19703);
and U19924 (N_19924,N_19775,N_19779);
nand U19925 (N_19925,N_19746,N_19754);
and U19926 (N_19926,N_19748,N_19824);
and U19927 (N_19927,N_19738,N_19820);
nand U19928 (N_19928,N_19687,N_19761);
nand U19929 (N_19929,N_19764,N_19753);
and U19930 (N_19930,N_19733,N_19750);
or U19931 (N_19931,N_19734,N_19759);
or U19932 (N_19932,N_19742,N_19730);
or U19933 (N_19933,N_19762,N_19823);
xor U19934 (N_19934,N_19697,N_19727);
nor U19935 (N_19935,N_19742,N_19810);
xnor U19936 (N_19936,N_19834,N_19798);
nand U19937 (N_19937,N_19780,N_19813);
nor U19938 (N_19938,N_19791,N_19780);
or U19939 (N_19939,N_19790,N_19721);
nor U19940 (N_19940,N_19683,N_19729);
nor U19941 (N_19941,N_19822,N_19814);
xnor U19942 (N_19942,N_19809,N_19692);
and U19943 (N_19943,N_19682,N_19713);
and U19944 (N_19944,N_19797,N_19773);
or U19945 (N_19945,N_19763,N_19789);
nor U19946 (N_19946,N_19682,N_19695);
and U19947 (N_19947,N_19690,N_19786);
xnor U19948 (N_19948,N_19802,N_19781);
and U19949 (N_19949,N_19732,N_19701);
and U19950 (N_19950,N_19722,N_19735);
nand U19951 (N_19951,N_19752,N_19730);
nor U19952 (N_19952,N_19705,N_19722);
and U19953 (N_19953,N_19696,N_19813);
and U19954 (N_19954,N_19808,N_19777);
xor U19955 (N_19955,N_19741,N_19745);
xor U19956 (N_19956,N_19746,N_19786);
nor U19957 (N_19957,N_19687,N_19713);
xor U19958 (N_19958,N_19774,N_19693);
and U19959 (N_19959,N_19778,N_19695);
nor U19960 (N_19960,N_19789,N_19697);
or U19961 (N_19961,N_19815,N_19732);
xor U19962 (N_19962,N_19787,N_19825);
or U19963 (N_19963,N_19747,N_19780);
and U19964 (N_19964,N_19786,N_19681);
nand U19965 (N_19965,N_19746,N_19691);
or U19966 (N_19966,N_19804,N_19799);
or U19967 (N_19967,N_19771,N_19733);
nor U19968 (N_19968,N_19802,N_19722);
xor U19969 (N_19969,N_19712,N_19724);
nor U19970 (N_19970,N_19790,N_19699);
and U19971 (N_19971,N_19685,N_19764);
nand U19972 (N_19972,N_19800,N_19834);
or U19973 (N_19973,N_19723,N_19736);
or U19974 (N_19974,N_19743,N_19763);
and U19975 (N_19975,N_19745,N_19816);
nor U19976 (N_19976,N_19776,N_19809);
or U19977 (N_19977,N_19766,N_19795);
nand U19978 (N_19978,N_19827,N_19769);
xor U19979 (N_19979,N_19695,N_19701);
and U19980 (N_19980,N_19837,N_19839);
nand U19981 (N_19981,N_19686,N_19733);
xnor U19982 (N_19982,N_19745,N_19815);
nand U19983 (N_19983,N_19822,N_19747);
or U19984 (N_19984,N_19773,N_19827);
nor U19985 (N_19985,N_19742,N_19695);
or U19986 (N_19986,N_19703,N_19818);
and U19987 (N_19987,N_19743,N_19779);
and U19988 (N_19988,N_19800,N_19762);
nand U19989 (N_19989,N_19790,N_19821);
nand U19990 (N_19990,N_19729,N_19680);
nand U19991 (N_19991,N_19816,N_19823);
and U19992 (N_19992,N_19825,N_19771);
xnor U19993 (N_19993,N_19698,N_19809);
or U19994 (N_19994,N_19769,N_19724);
nor U19995 (N_19995,N_19798,N_19769);
nor U19996 (N_19996,N_19804,N_19742);
nand U19997 (N_19997,N_19788,N_19838);
nor U19998 (N_19998,N_19816,N_19709);
nand U19999 (N_19999,N_19822,N_19787);
nand UO_0 (O_0,N_19986,N_19981);
nor UO_1 (O_1,N_19945,N_19957);
or UO_2 (O_2,N_19896,N_19859);
or UO_3 (O_3,N_19966,N_19911);
xor UO_4 (O_4,N_19882,N_19931);
and UO_5 (O_5,N_19942,N_19972);
nor UO_6 (O_6,N_19897,N_19925);
or UO_7 (O_7,N_19869,N_19943);
xnor UO_8 (O_8,N_19965,N_19893);
nor UO_9 (O_9,N_19973,N_19849);
and UO_10 (O_10,N_19894,N_19903);
xnor UO_11 (O_11,N_19941,N_19995);
or UO_12 (O_12,N_19851,N_19938);
nand UO_13 (O_13,N_19952,N_19856);
or UO_14 (O_14,N_19919,N_19861);
and UO_15 (O_15,N_19910,N_19977);
nor UO_16 (O_16,N_19914,N_19866);
nand UO_17 (O_17,N_19949,N_19907);
and UO_18 (O_18,N_19992,N_19970);
or UO_19 (O_19,N_19979,N_19927);
xnor UO_20 (O_20,N_19921,N_19918);
nand UO_21 (O_21,N_19864,N_19976);
nor UO_22 (O_22,N_19886,N_19960);
nor UO_23 (O_23,N_19905,N_19985);
or UO_24 (O_24,N_19948,N_19915);
nor UO_25 (O_25,N_19877,N_19974);
and UO_26 (O_26,N_19964,N_19902);
and UO_27 (O_27,N_19889,N_19954);
xor UO_28 (O_28,N_19924,N_19904);
nand UO_29 (O_29,N_19850,N_19999);
xor UO_30 (O_30,N_19855,N_19936);
nand UO_31 (O_31,N_19884,N_19940);
nand UO_32 (O_32,N_19944,N_19852);
or UO_33 (O_33,N_19934,N_19908);
nor UO_34 (O_34,N_19888,N_19917);
or UO_35 (O_35,N_19841,N_19885);
or UO_36 (O_36,N_19874,N_19916);
xor UO_37 (O_37,N_19989,N_19983);
or UO_38 (O_38,N_19891,N_19858);
or UO_39 (O_39,N_19848,N_19840);
or UO_40 (O_40,N_19937,N_19860);
and UO_41 (O_41,N_19857,N_19959);
and UO_42 (O_42,N_19878,N_19879);
nor UO_43 (O_43,N_19843,N_19939);
and UO_44 (O_44,N_19880,N_19984);
or UO_45 (O_45,N_19968,N_19978);
xnor UO_46 (O_46,N_19876,N_19933);
xor UO_47 (O_47,N_19998,N_19871);
nor UO_48 (O_48,N_19920,N_19953);
or UO_49 (O_49,N_19870,N_19887);
or UO_50 (O_50,N_19987,N_19988);
nand UO_51 (O_51,N_19863,N_19956);
or UO_52 (O_52,N_19969,N_19913);
and UO_53 (O_53,N_19967,N_19898);
nand UO_54 (O_54,N_19872,N_19930);
xnor UO_55 (O_55,N_19961,N_19881);
xor UO_56 (O_56,N_19975,N_19895);
nor UO_57 (O_57,N_19862,N_19906);
nor UO_58 (O_58,N_19946,N_19947);
and UO_59 (O_59,N_19963,N_19846);
nor UO_60 (O_60,N_19991,N_19928);
nor UO_61 (O_61,N_19950,N_19890);
or UO_62 (O_62,N_19971,N_19875);
nor UO_63 (O_63,N_19962,N_19867);
nand UO_64 (O_64,N_19923,N_19926);
nor UO_65 (O_65,N_19892,N_19847);
xnor UO_66 (O_66,N_19990,N_19900);
and UO_67 (O_67,N_19994,N_19955);
and UO_68 (O_68,N_19993,N_19980);
nand UO_69 (O_69,N_19883,N_19932);
and UO_70 (O_70,N_19922,N_19845);
and UO_71 (O_71,N_19873,N_19865);
xnor UO_72 (O_72,N_19853,N_19982);
or UO_73 (O_73,N_19899,N_19909);
nand UO_74 (O_74,N_19929,N_19842);
and UO_75 (O_75,N_19951,N_19854);
xor UO_76 (O_76,N_19868,N_19958);
xnor UO_77 (O_77,N_19997,N_19912);
nor UO_78 (O_78,N_19901,N_19996);
nand UO_79 (O_79,N_19844,N_19935);
and UO_80 (O_80,N_19913,N_19934);
and UO_81 (O_81,N_19947,N_19975);
and UO_82 (O_82,N_19981,N_19873);
and UO_83 (O_83,N_19922,N_19965);
or UO_84 (O_84,N_19879,N_19990);
xor UO_85 (O_85,N_19985,N_19927);
or UO_86 (O_86,N_19996,N_19991);
and UO_87 (O_87,N_19905,N_19962);
xor UO_88 (O_88,N_19888,N_19931);
or UO_89 (O_89,N_19890,N_19918);
nor UO_90 (O_90,N_19890,N_19985);
xnor UO_91 (O_91,N_19932,N_19918);
nor UO_92 (O_92,N_19932,N_19876);
or UO_93 (O_93,N_19936,N_19993);
nand UO_94 (O_94,N_19952,N_19914);
or UO_95 (O_95,N_19866,N_19875);
xnor UO_96 (O_96,N_19986,N_19873);
nand UO_97 (O_97,N_19928,N_19894);
nand UO_98 (O_98,N_19991,N_19888);
nor UO_99 (O_99,N_19870,N_19939);
nor UO_100 (O_100,N_19843,N_19977);
xnor UO_101 (O_101,N_19938,N_19993);
xor UO_102 (O_102,N_19878,N_19987);
nor UO_103 (O_103,N_19999,N_19857);
nor UO_104 (O_104,N_19863,N_19994);
nand UO_105 (O_105,N_19984,N_19909);
and UO_106 (O_106,N_19926,N_19856);
xnor UO_107 (O_107,N_19950,N_19854);
nor UO_108 (O_108,N_19892,N_19928);
nor UO_109 (O_109,N_19903,N_19968);
and UO_110 (O_110,N_19993,N_19853);
nor UO_111 (O_111,N_19907,N_19929);
nand UO_112 (O_112,N_19917,N_19928);
xor UO_113 (O_113,N_19977,N_19984);
nor UO_114 (O_114,N_19849,N_19936);
nand UO_115 (O_115,N_19959,N_19969);
or UO_116 (O_116,N_19988,N_19843);
or UO_117 (O_117,N_19872,N_19885);
and UO_118 (O_118,N_19999,N_19841);
xor UO_119 (O_119,N_19989,N_19904);
nand UO_120 (O_120,N_19986,N_19867);
and UO_121 (O_121,N_19971,N_19979);
or UO_122 (O_122,N_19873,N_19899);
nor UO_123 (O_123,N_19864,N_19982);
and UO_124 (O_124,N_19988,N_19984);
xor UO_125 (O_125,N_19932,N_19908);
nand UO_126 (O_126,N_19855,N_19893);
or UO_127 (O_127,N_19918,N_19971);
nor UO_128 (O_128,N_19949,N_19970);
nand UO_129 (O_129,N_19926,N_19996);
nor UO_130 (O_130,N_19861,N_19950);
nand UO_131 (O_131,N_19931,N_19922);
nor UO_132 (O_132,N_19941,N_19894);
nand UO_133 (O_133,N_19931,N_19886);
nand UO_134 (O_134,N_19895,N_19874);
nand UO_135 (O_135,N_19912,N_19887);
nor UO_136 (O_136,N_19889,N_19951);
nor UO_137 (O_137,N_19961,N_19879);
xor UO_138 (O_138,N_19885,N_19909);
xnor UO_139 (O_139,N_19908,N_19847);
or UO_140 (O_140,N_19860,N_19981);
nor UO_141 (O_141,N_19952,N_19909);
nor UO_142 (O_142,N_19842,N_19923);
nor UO_143 (O_143,N_19882,N_19959);
nand UO_144 (O_144,N_19953,N_19870);
xnor UO_145 (O_145,N_19887,N_19975);
nor UO_146 (O_146,N_19872,N_19881);
or UO_147 (O_147,N_19859,N_19989);
xor UO_148 (O_148,N_19877,N_19950);
xor UO_149 (O_149,N_19902,N_19887);
xor UO_150 (O_150,N_19854,N_19949);
and UO_151 (O_151,N_19892,N_19899);
xor UO_152 (O_152,N_19848,N_19935);
and UO_153 (O_153,N_19912,N_19989);
or UO_154 (O_154,N_19884,N_19972);
or UO_155 (O_155,N_19929,N_19911);
nor UO_156 (O_156,N_19858,N_19936);
and UO_157 (O_157,N_19943,N_19971);
xor UO_158 (O_158,N_19912,N_19944);
and UO_159 (O_159,N_19874,N_19902);
or UO_160 (O_160,N_19989,N_19846);
nor UO_161 (O_161,N_19968,N_19926);
xor UO_162 (O_162,N_19868,N_19919);
or UO_163 (O_163,N_19899,N_19961);
nand UO_164 (O_164,N_19947,N_19974);
xor UO_165 (O_165,N_19852,N_19859);
xnor UO_166 (O_166,N_19879,N_19842);
or UO_167 (O_167,N_19855,N_19881);
or UO_168 (O_168,N_19968,N_19944);
and UO_169 (O_169,N_19863,N_19960);
nor UO_170 (O_170,N_19868,N_19929);
nor UO_171 (O_171,N_19965,N_19996);
nand UO_172 (O_172,N_19990,N_19961);
or UO_173 (O_173,N_19984,N_19983);
nor UO_174 (O_174,N_19860,N_19857);
nor UO_175 (O_175,N_19886,N_19850);
nor UO_176 (O_176,N_19965,N_19917);
or UO_177 (O_177,N_19936,N_19879);
nand UO_178 (O_178,N_19950,N_19975);
and UO_179 (O_179,N_19850,N_19905);
or UO_180 (O_180,N_19909,N_19854);
nor UO_181 (O_181,N_19951,N_19972);
or UO_182 (O_182,N_19965,N_19898);
or UO_183 (O_183,N_19936,N_19876);
nand UO_184 (O_184,N_19863,N_19931);
xnor UO_185 (O_185,N_19985,N_19957);
nor UO_186 (O_186,N_19976,N_19919);
and UO_187 (O_187,N_19968,N_19887);
nor UO_188 (O_188,N_19915,N_19978);
and UO_189 (O_189,N_19864,N_19981);
xnor UO_190 (O_190,N_19884,N_19929);
nor UO_191 (O_191,N_19988,N_19968);
nand UO_192 (O_192,N_19918,N_19991);
nand UO_193 (O_193,N_19977,N_19899);
xnor UO_194 (O_194,N_19859,N_19899);
xor UO_195 (O_195,N_19939,N_19919);
and UO_196 (O_196,N_19896,N_19940);
nor UO_197 (O_197,N_19947,N_19953);
xor UO_198 (O_198,N_19969,N_19877);
xnor UO_199 (O_199,N_19891,N_19934);
nor UO_200 (O_200,N_19961,N_19933);
xnor UO_201 (O_201,N_19932,N_19885);
nor UO_202 (O_202,N_19963,N_19974);
xnor UO_203 (O_203,N_19858,N_19973);
or UO_204 (O_204,N_19962,N_19857);
nor UO_205 (O_205,N_19909,N_19852);
xnor UO_206 (O_206,N_19989,N_19942);
nand UO_207 (O_207,N_19840,N_19959);
or UO_208 (O_208,N_19941,N_19933);
and UO_209 (O_209,N_19946,N_19888);
xnor UO_210 (O_210,N_19900,N_19950);
xor UO_211 (O_211,N_19892,N_19909);
xnor UO_212 (O_212,N_19926,N_19869);
xnor UO_213 (O_213,N_19902,N_19927);
and UO_214 (O_214,N_19868,N_19881);
xnor UO_215 (O_215,N_19976,N_19888);
nand UO_216 (O_216,N_19949,N_19863);
nand UO_217 (O_217,N_19923,N_19893);
or UO_218 (O_218,N_19866,N_19863);
nand UO_219 (O_219,N_19878,N_19882);
xor UO_220 (O_220,N_19851,N_19960);
nand UO_221 (O_221,N_19910,N_19937);
nor UO_222 (O_222,N_19953,N_19881);
and UO_223 (O_223,N_19982,N_19908);
and UO_224 (O_224,N_19963,N_19862);
or UO_225 (O_225,N_19930,N_19918);
and UO_226 (O_226,N_19895,N_19910);
and UO_227 (O_227,N_19894,N_19888);
and UO_228 (O_228,N_19921,N_19994);
nand UO_229 (O_229,N_19880,N_19881);
xnor UO_230 (O_230,N_19967,N_19943);
xnor UO_231 (O_231,N_19939,N_19901);
nor UO_232 (O_232,N_19894,N_19902);
xor UO_233 (O_233,N_19969,N_19923);
or UO_234 (O_234,N_19869,N_19874);
xor UO_235 (O_235,N_19841,N_19933);
xnor UO_236 (O_236,N_19907,N_19939);
nand UO_237 (O_237,N_19860,N_19964);
or UO_238 (O_238,N_19986,N_19902);
nor UO_239 (O_239,N_19944,N_19856);
nor UO_240 (O_240,N_19925,N_19980);
nor UO_241 (O_241,N_19848,N_19999);
nor UO_242 (O_242,N_19930,N_19894);
xor UO_243 (O_243,N_19850,N_19986);
nand UO_244 (O_244,N_19900,N_19901);
or UO_245 (O_245,N_19963,N_19951);
or UO_246 (O_246,N_19925,N_19849);
xor UO_247 (O_247,N_19881,N_19852);
or UO_248 (O_248,N_19850,N_19946);
nor UO_249 (O_249,N_19916,N_19975);
nor UO_250 (O_250,N_19927,N_19952);
xnor UO_251 (O_251,N_19971,N_19887);
and UO_252 (O_252,N_19959,N_19876);
and UO_253 (O_253,N_19904,N_19986);
or UO_254 (O_254,N_19997,N_19962);
xnor UO_255 (O_255,N_19932,N_19923);
xnor UO_256 (O_256,N_19949,N_19968);
nor UO_257 (O_257,N_19901,N_19877);
nor UO_258 (O_258,N_19983,N_19948);
nor UO_259 (O_259,N_19900,N_19947);
or UO_260 (O_260,N_19917,N_19920);
xnor UO_261 (O_261,N_19996,N_19855);
or UO_262 (O_262,N_19897,N_19952);
xnor UO_263 (O_263,N_19993,N_19855);
and UO_264 (O_264,N_19852,N_19970);
and UO_265 (O_265,N_19852,N_19949);
xor UO_266 (O_266,N_19915,N_19987);
xor UO_267 (O_267,N_19991,N_19971);
xor UO_268 (O_268,N_19883,N_19918);
and UO_269 (O_269,N_19967,N_19995);
nand UO_270 (O_270,N_19856,N_19916);
or UO_271 (O_271,N_19890,N_19922);
or UO_272 (O_272,N_19942,N_19951);
or UO_273 (O_273,N_19999,N_19974);
nand UO_274 (O_274,N_19949,N_19874);
nand UO_275 (O_275,N_19877,N_19895);
and UO_276 (O_276,N_19976,N_19979);
nor UO_277 (O_277,N_19924,N_19955);
xor UO_278 (O_278,N_19978,N_19910);
xnor UO_279 (O_279,N_19986,N_19870);
and UO_280 (O_280,N_19869,N_19887);
nand UO_281 (O_281,N_19959,N_19953);
and UO_282 (O_282,N_19849,N_19993);
xnor UO_283 (O_283,N_19885,N_19884);
nor UO_284 (O_284,N_19981,N_19975);
or UO_285 (O_285,N_19975,N_19849);
nand UO_286 (O_286,N_19983,N_19927);
nor UO_287 (O_287,N_19933,N_19919);
xor UO_288 (O_288,N_19868,N_19997);
nand UO_289 (O_289,N_19964,N_19976);
and UO_290 (O_290,N_19966,N_19983);
and UO_291 (O_291,N_19981,N_19857);
or UO_292 (O_292,N_19947,N_19988);
nor UO_293 (O_293,N_19947,N_19869);
and UO_294 (O_294,N_19960,N_19872);
xnor UO_295 (O_295,N_19888,N_19868);
or UO_296 (O_296,N_19921,N_19864);
and UO_297 (O_297,N_19966,N_19954);
xnor UO_298 (O_298,N_19996,N_19883);
nand UO_299 (O_299,N_19971,N_19858);
xnor UO_300 (O_300,N_19916,N_19883);
and UO_301 (O_301,N_19978,N_19897);
nand UO_302 (O_302,N_19984,N_19901);
xnor UO_303 (O_303,N_19926,N_19876);
xor UO_304 (O_304,N_19988,N_19989);
nand UO_305 (O_305,N_19912,N_19877);
xor UO_306 (O_306,N_19889,N_19864);
xnor UO_307 (O_307,N_19925,N_19931);
and UO_308 (O_308,N_19981,N_19885);
nor UO_309 (O_309,N_19870,N_19940);
nand UO_310 (O_310,N_19917,N_19930);
or UO_311 (O_311,N_19965,N_19952);
or UO_312 (O_312,N_19892,N_19940);
nor UO_313 (O_313,N_19940,N_19864);
or UO_314 (O_314,N_19938,N_19914);
xor UO_315 (O_315,N_19849,N_19976);
nor UO_316 (O_316,N_19965,N_19861);
nand UO_317 (O_317,N_19997,N_19922);
nor UO_318 (O_318,N_19923,N_19949);
and UO_319 (O_319,N_19980,N_19904);
xnor UO_320 (O_320,N_19971,N_19844);
or UO_321 (O_321,N_19974,N_19903);
and UO_322 (O_322,N_19844,N_19922);
nand UO_323 (O_323,N_19913,N_19947);
nor UO_324 (O_324,N_19967,N_19887);
xor UO_325 (O_325,N_19998,N_19994);
xnor UO_326 (O_326,N_19931,N_19917);
nor UO_327 (O_327,N_19846,N_19874);
nand UO_328 (O_328,N_19961,N_19885);
nand UO_329 (O_329,N_19848,N_19921);
and UO_330 (O_330,N_19967,N_19987);
and UO_331 (O_331,N_19966,N_19943);
nor UO_332 (O_332,N_19945,N_19881);
or UO_333 (O_333,N_19982,N_19963);
or UO_334 (O_334,N_19894,N_19923);
nand UO_335 (O_335,N_19907,N_19957);
nor UO_336 (O_336,N_19877,N_19843);
nor UO_337 (O_337,N_19897,N_19992);
and UO_338 (O_338,N_19961,N_19958);
nand UO_339 (O_339,N_19854,N_19958);
xnor UO_340 (O_340,N_19969,N_19986);
or UO_341 (O_341,N_19988,N_19994);
nor UO_342 (O_342,N_19991,N_19990);
nor UO_343 (O_343,N_19942,N_19993);
nand UO_344 (O_344,N_19853,N_19936);
nor UO_345 (O_345,N_19951,N_19917);
or UO_346 (O_346,N_19977,N_19989);
nand UO_347 (O_347,N_19885,N_19982);
nand UO_348 (O_348,N_19997,N_19891);
nor UO_349 (O_349,N_19866,N_19916);
or UO_350 (O_350,N_19873,N_19945);
or UO_351 (O_351,N_19867,N_19896);
or UO_352 (O_352,N_19994,N_19924);
and UO_353 (O_353,N_19878,N_19960);
nor UO_354 (O_354,N_19907,N_19873);
nand UO_355 (O_355,N_19926,N_19878);
or UO_356 (O_356,N_19866,N_19957);
and UO_357 (O_357,N_19868,N_19994);
and UO_358 (O_358,N_19854,N_19993);
nand UO_359 (O_359,N_19918,N_19962);
and UO_360 (O_360,N_19973,N_19851);
xor UO_361 (O_361,N_19987,N_19958);
nor UO_362 (O_362,N_19958,N_19966);
or UO_363 (O_363,N_19949,N_19991);
xnor UO_364 (O_364,N_19890,N_19897);
nand UO_365 (O_365,N_19845,N_19850);
nor UO_366 (O_366,N_19934,N_19924);
nand UO_367 (O_367,N_19842,N_19897);
nand UO_368 (O_368,N_19967,N_19844);
and UO_369 (O_369,N_19919,N_19989);
and UO_370 (O_370,N_19994,N_19953);
and UO_371 (O_371,N_19936,N_19884);
nand UO_372 (O_372,N_19953,N_19951);
or UO_373 (O_373,N_19956,N_19975);
nor UO_374 (O_374,N_19870,N_19860);
or UO_375 (O_375,N_19933,N_19854);
or UO_376 (O_376,N_19959,N_19846);
nor UO_377 (O_377,N_19855,N_19979);
nand UO_378 (O_378,N_19993,N_19912);
xor UO_379 (O_379,N_19847,N_19926);
nor UO_380 (O_380,N_19900,N_19868);
or UO_381 (O_381,N_19909,N_19868);
nand UO_382 (O_382,N_19865,N_19991);
xnor UO_383 (O_383,N_19865,N_19987);
xor UO_384 (O_384,N_19890,N_19912);
nor UO_385 (O_385,N_19982,N_19951);
xnor UO_386 (O_386,N_19949,N_19855);
nor UO_387 (O_387,N_19987,N_19999);
nand UO_388 (O_388,N_19895,N_19869);
or UO_389 (O_389,N_19988,N_19851);
xnor UO_390 (O_390,N_19851,N_19927);
xor UO_391 (O_391,N_19914,N_19972);
nor UO_392 (O_392,N_19985,N_19958);
xor UO_393 (O_393,N_19998,N_19996);
and UO_394 (O_394,N_19994,N_19956);
xnor UO_395 (O_395,N_19846,N_19844);
nand UO_396 (O_396,N_19950,N_19944);
nor UO_397 (O_397,N_19895,N_19859);
nand UO_398 (O_398,N_19900,N_19883);
or UO_399 (O_399,N_19872,N_19989);
nand UO_400 (O_400,N_19895,N_19907);
and UO_401 (O_401,N_19884,N_19980);
xnor UO_402 (O_402,N_19962,N_19949);
and UO_403 (O_403,N_19988,N_19906);
or UO_404 (O_404,N_19960,N_19901);
and UO_405 (O_405,N_19910,N_19954);
xnor UO_406 (O_406,N_19950,N_19924);
and UO_407 (O_407,N_19979,N_19857);
xnor UO_408 (O_408,N_19899,N_19905);
xnor UO_409 (O_409,N_19890,N_19858);
and UO_410 (O_410,N_19982,N_19996);
xor UO_411 (O_411,N_19877,N_19887);
and UO_412 (O_412,N_19843,N_19883);
nand UO_413 (O_413,N_19900,N_19875);
and UO_414 (O_414,N_19940,N_19882);
or UO_415 (O_415,N_19925,N_19964);
or UO_416 (O_416,N_19853,N_19961);
and UO_417 (O_417,N_19841,N_19998);
nor UO_418 (O_418,N_19878,N_19953);
or UO_419 (O_419,N_19969,N_19882);
or UO_420 (O_420,N_19916,N_19987);
and UO_421 (O_421,N_19951,N_19901);
or UO_422 (O_422,N_19862,N_19865);
nand UO_423 (O_423,N_19943,N_19994);
and UO_424 (O_424,N_19978,N_19960);
nor UO_425 (O_425,N_19990,N_19923);
or UO_426 (O_426,N_19881,N_19960);
and UO_427 (O_427,N_19918,N_19898);
and UO_428 (O_428,N_19971,N_19890);
or UO_429 (O_429,N_19925,N_19984);
xor UO_430 (O_430,N_19953,N_19913);
nand UO_431 (O_431,N_19943,N_19973);
and UO_432 (O_432,N_19973,N_19896);
nor UO_433 (O_433,N_19964,N_19975);
xor UO_434 (O_434,N_19910,N_19926);
or UO_435 (O_435,N_19969,N_19965);
nor UO_436 (O_436,N_19984,N_19948);
or UO_437 (O_437,N_19879,N_19895);
nor UO_438 (O_438,N_19963,N_19910);
nand UO_439 (O_439,N_19905,N_19876);
nor UO_440 (O_440,N_19982,N_19852);
and UO_441 (O_441,N_19868,N_19864);
nand UO_442 (O_442,N_19966,N_19847);
or UO_443 (O_443,N_19951,N_19878);
nand UO_444 (O_444,N_19938,N_19863);
xor UO_445 (O_445,N_19881,N_19904);
xnor UO_446 (O_446,N_19958,N_19990);
nor UO_447 (O_447,N_19973,N_19897);
xor UO_448 (O_448,N_19897,N_19922);
nor UO_449 (O_449,N_19872,N_19963);
xor UO_450 (O_450,N_19997,N_19880);
or UO_451 (O_451,N_19887,N_19943);
and UO_452 (O_452,N_19978,N_19850);
nor UO_453 (O_453,N_19911,N_19899);
xor UO_454 (O_454,N_19890,N_19970);
and UO_455 (O_455,N_19883,N_19980);
or UO_456 (O_456,N_19957,N_19917);
nor UO_457 (O_457,N_19870,N_19919);
xnor UO_458 (O_458,N_19960,N_19897);
xor UO_459 (O_459,N_19993,N_19890);
xnor UO_460 (O_460,N_19874,N_19984);
nand UO_461 (O_461,N_19990,N_19960);
nor UO_462 (O_462,N_19893,N_19999);
nand UO_463 (O_463,N_19844,N_19902);
or UO_464 (O_464,N_19969,N_19889);
nor UO_465 (O_465,N_19880,N_19991);
nand UO_466 (O_466,N_19957,N_19855);
nor UO_467 (O_467,N_19878,N_19958);
nor UO_468 (O_468,N_19860,N_19947);
xor UO_469 (O_469,N_19862,N_19914);
xor UO_470 (O_470,N_19958,N_19879);
nor UO_471 (O_471,N_19943,N_19974);
nand UO_472 (O_472,N_19969,N_19930);
or UO_473 (O_473,N_19989,N_19916);
and UO_474 (O_474,N_19987,N_19970);
xnor UO_475 (O_475,N_19918,N_19915);
xor UO_476 (O_476,N_19847,N_19842);
nor UO_477 (O_477,N_19887,N_19862);
nand UO_478 (O_478,N_19986,N_19872);
nand UO_479 (O_479,N_19974,N_19875);
or UO_480 (O_480,N_19941,N_19948);
nand UO_481 (O_481,N_19865,N_19859);
xnor UO_482 (O_482,N_19996,N_19967);
xnor UO_483 (O_483,N_19840,N_19907);
and UO_484 (O_484,N_19901,N_19934);
nor UO_485 (O_485,N_19948,N_19996);
xor UO_486 (O_486,N_19944,N_19872);
nand UO_487 (O_487,N_19931,N_19960);
and UO_488 (O_488,N_19861,N_19957);
xnor UO_489 (O_489,N_19853,N_19887);
or UO_490 (O_490,N_19844,N_19872);
nor UO_491 (O_491,N_19936,N_19887);
nand UO_492 (O_492,N_19906,N_19898);
and UO_493 (O_493,N_19944,N_19876);
xnor UO_494 (O_494,N_19979,N_19977);
or UO_495 (O_495,N_19967,N_19855);
xor UO_496 (O_496,N_19854,N_19925);
nand UO_497 (O_497,N_19934,N_19892);
nand UO_498 (O_498,N_19913,N_19995);
and UO_499 (O_499,N_19930,N_19982);
or UO_500 (O_500,N_19959,N_19904);
or UO_501 (O_501,N_19954,N_19919);
xnor UO_502 (O_502,N_19950,N_19945);
nand UO_503 (O_503,N_19922,N_19891);
xor UO_504 (O_504,N_19959,N_19919);
nor UO_505 (O_505,N_19990,N_19846);
nand UO_506 (O_506,N_19869,N_19861);
xnor UO_507 (O_507,N_19902,N_19982);
or UO_508 (O_508,N_19842,N_19855);
or UO_509 (O_509,N_19841,N_19844);
xnor UO_510 (O_510,N_19955,N_19932);
nor UO_511 (O_511,N_19929,N_19933);
nor UO_512 (O_512,N_19874,N_19993);
nand UO_513 (O_513,N_19896,N_19891);
nor UO_514 (O_514,N_19904,N_19888);
xnor UO_515 (O_515,N_19858,N_19874);
xor UO_516 (O_516,N_19906,N_19985);
xnor UO_517 (O_517,N_19877,N_19868);
and UO_518 (O_518,N_19973,N_19852);
and UO_519 (O_519,N_19971,N_19897);
xor UO_520 (O_520,N_19842,N_19958);
xor UO_521 (O_521,N_19856,N_19923);
nor UO_522 (O_522,N_19858,N_19913);
or UO_523 (O_523,N_19893,N_19981);
and UO_524 (O_524,N_19987,N_19975);
or UO_525 (O_525,N_19988,N_19873);
or UO_526 (O_526,N_19934,N_19983);
xor UO_527 (O_527,N_19973,N_19864);
nand UO_528 (O_528,N_19919,N_19903);
and UO_529 (O_529,N_19954,N_19912);
xor UO_530 (O_530,N_19984,N_19921);
nand UO_531 (O_531,N_19970,N_19910);
or UO_532 (O_532,N_19844,N_19910);
nand UO_533 (O_533,N_19882,N_19922);
or UO_534 (O_534,N_19869,N_19886);
xnor UO_535 (O_535,N_19916,N_19997);
and UO_536 (O_536,N_19879,N_19968);
or UO_537 (O_537,N_19947,N_19893);
nand UO_538 (O_538,N_19995,N_19962);
nand UO_539 (O_539,N_19888,N_19983);
nand UO_540 (O_540,N_19958,N_19892);
nor UO_541 (O_541,N_19985,N_19911);
xnor UO_542 (O_542,N_19938,N_19905);
nand UO_543 (O_543,N_19908,N_19953);
nor UO_544 (O_544,N_19893,N_19974);
or UO_545 (O_545,N_19861,N_19988);
or UO_546 (O_546,N_19880,N_19922);
nand UO_547 (O_547,N_19943,N_19955);
xnor UO_548 (O_548,N_19961,N_19896);
nor UO_549 (O_549,N_19863,N_19858);
nor UO_550 (O_550,N_19888,N_19893);
nand UO_551 (O_551,N_19871,N_19924);
and UO_552 (O_552,N_19941,N_19978);
nand UO_553 (O_553,N_19974,N_19844);
nor UO_554 (O_554,N_19958,N_19866);
or UO_555 (O_555,N_19997,N_19996);
nand UO_556 (O_556,N_19884,N_19867);
nor UO_557 (O_557,N_19953,N_19907);
nand UO_558 (O_558,N_19901,N_19859);
or UO_559 (O_559,N_19904,N_19893);
nand UO_560 (O_560,N_19938,N_19983);
or UO_561 (O_561,N_19861,N_19927);
nand UO_562 (O_562,N_19984,N_19861);
nor UO_563 (O_563,N_19870,N_19909);
and UO_564 (O_564,N_19929,N_19908);
nor UO_565 (O_565,N_19923,N_19981);
or UO_566 (O_566,N_19995,N_19881);
nor UO_567 (O_567,N_19859,N_19910);
xor UO_568 (O_568,N_19972,N_19987);
nor UO_569 (O_569,N_19987,N_19937);
and UO_570 (O_570,N_19939,N_19866);
xor UO_571 (O_571,N_19916,N_19990);
nand UO_572 (O_572,N_19929,N_19916);
nor UO_573 (O_573,N_19975,N_19863);
and UO_574 (O_574,N_19869,N_19952);
nand UO_575 (O_575,N_19970,N_19961);
nand UO_576 (O_576,N_19888,N_19956);
xor UO_577 (O_577,N_19902,N_19975);
or UO_578 (O_578,N_19944,N_19987);
nand UO_579 (O_579,N_19915,N_19886);
nor UO_580 (O_580,N_19870,N_19922);
xor UO_581 (O_581,N_19933,N_19928);
nor UO_582 (O_582,N_19993,N_19965);
nor UO_583 (O_583,N_19984,N_19938);
nor UO_584 (O_584,N_19939,N_19865);
and UO_585 (O_585,N_19886,N_19983);
xnor UO_586 (O_586,N_19978,N_19900);
xor UO_587 (O_587,N_19929,N_19960);
nor UO_588 (O_588,N_19863,N_19933);
nand UO_589 (O_589,N_19904,N_19965);
xnor UO_590 (O_590,N_19910,N_19871);
nand UO_591 (O_591,N_19901,N_19856);
xnor UO_592 (O_592,N_19841,N_19923);
xor UO_593 (O_593,N_19881,N_19884);
xor UO_594 (O_594,N_19852,N_19937);
or UO_595 (O_595,N_19923,N_19861);
or UO_596 (O_596,N_19933,N_19963);
and UO_597 (O_597,N_19946,N_19867);
nor UO_598 (O_598,N_19867,N_19846);
and UO_599 (O_599,N_19911,N_19910);
and UO_600 (O_600,N_19864,N_19906);
nand UO_601 (O_601,N_19864,N_19960);
nor UO_602 (O_602,N_19891,N_19908);
and UO_603 (O_603,N_19863,N_19895);
nand UO_604 (O_604,N_19953,N_19973);
nor UO_605 (O_605,N_19896,N_19875);
or UO_606 (O_606,N_19964,N_19910);
or UO_607 (O_607,N_19917,N_19913);
or UO_608 (O_608,N_19950,N_19910);
nand UO_609 (O_609,N_19885,N_19916);
nor UO_610 (O_610,N_19947,N_19960);
and UO_611 (O_611,N_19890,N_19996);
and UO_612 (O_612,N_19870,N_19863);
or UO_613 (O_613,N_19863,N_19844);
and UO_614 (O_614,N_19914,N_19847);
nand UO_615 (O_615,N_19950,N_19969);
nor UO_616 (O_616,N_19893,N_19927);
and UO_617 (O_617,N_19895,N_19953);
nand UO_618 (O_618,N_19844,N_19955);
or UO_619 (O_619,N_19870,N_19895);
or UO_620 (O_620,N_19954,N_19931);
xnor UO_621 (O_621,N_19857,N_19849);
xnor UO_622 (O_622,N_19989,N_19841);
nand UO_623 (O_623,N_19872,N_19955);
and UO_624 (O_624,N_19977,N_19863);
xnor UO_625 (O_625,N_19926,N_19972);
and UO_626 (O_626,N_19885,N_19991);
nand UO_627 (O_627,N_19925,N_19955);
xor UO_628 (O_628,N_19906,N_19934);
and UO_629 (O_629,N_19978,N_19972);
nor UO_630 (O_630,N_19980,N_19995);
or UO_631 (O_631,N_19949,N_19846);
xor UO_632 (O_632,N_19921,N_19976);
nand UO_633 (O_633,N_19980,N_19890);
and UO_634 (O_634,N_19912,N_19913);
and UO_635 (O_635,N_19898,N_19964);
xnor UO_636 (O_636,N_19950,N_19840);
nor UO_637 (O_637,N_19861,N_19901);
nand UO_638 (O_638,N_19962,N_19894);
xor UO_639 (O_639,N_19861,N_19886);
nor UO_640 (O_640,N_19996,N_19857);
xnor UO_641 (O_641,N_19844,N_19889);
and UO_642 (O_642,N_19961,N_19984);
and UO_643 (O_643,N_19858,N_19875);
nand UO_644 (O_644,N_19907,N_19888);
nand UO_645 (O_645,N_19935,N_19992);
and UO_646 (O_646,N_19883,N_19912);
nor UO_647 (O_647,N_19997,N_19898);
xnor UO_648 (O_648,N_19843,N_19906);
or UO_649 (O_649,N_19852,N_19921);
xor UO_650 (O_650,N_19994,N_19849);
nor UO_651 (O_651,N_19932,N_19892);
and UO_652 (O_652,N_19984,N_19949);
xnor UO_653 (O_653,N_19851,N_19953);
xnor UO_654 (O_654,N_19867,N_19951);
and UO_655 (O_655,N_19898,N_19924);
xnor UO_656 (O_656,N_19980,N_19952);
xor UO_657 (O_657,N_19906,N_19935);
nand UO_658 (O_658,N_19981,N_19997);
nor UO_659 (O_659,N_19958,N_19869);
nand UO_660 (O_660,N_19858,N_19882);
and UO_661 (O_661,N_19940,N_19904);
xor UO_662 (O_662,N_19865,N_19996);
or UO_663 (O_663,N_19852,N_19959);
nor UO_664 (O_664,N_19913,N_19915);
nor UO_665 (O_665,N_19939,N_19874);
nor UO_666 (O_666,N_19873,N_19956);
or UO_667 (O_667,N_19894,N_19886);
nand UO_668 (O_668,N_19883,N_19922);
or UO_669 (O_669,N_19982,N_19933);
and UO_670 (O_670,N_19893,N_19887);
xnor UO_671 (O_671,N_19849,N_19927);
and UO_672 (O_672,N_19991,N_19951);
xor UO_673 (O_673,N_19920,N_19895);
or UO_674 (O_674,N_19934,N_19928);
nor UO_675 (O_675,N_19854,N_19895);
nor UO_676 (O_676,N_19850,N_19843);
xnor UO_677 (O_677,N_19885,N_19965);
or UO_678 (O_678,N_19971,N_19906);
nor UO_679 (O_679,N_19958,N_19893);
nor UO_680 (O_680,N_19899,N_19856);
nor UO_681 (O_681,N_19847,N_19890);
and UO_682 (O_682,N_19973,N_19934);
xor UO_683 (O_683,N_19999,N_19872);
nand UO_684 (O_684,N_19881,N_19898);
nor UO_685 (O_685,N_19882,N_19984);
and UO_686 (O_686,N_19945,N_19890);
or UO_687 (O_687,N_19918,N_19992);
xor UO_688 (O_688,N_19968,N_19995);
nand UO_689 (O_689,N_19940,N_19944);
nor UO_690 (O_690,N_19851,N_19844);
xnor UO_691 (O_691,N_19857,N_19885);
and UO_692 (O_692,N_19908,N_19911);
nand UO_693 (O_693,N_19954,N_19935);
nor UO_694 (O_694,N_19975,N_19865);
xor UO_695 (O_695,N_19989,N_19843);
xnor UO_696 (O_696,N_19959,N_19987);
nand UO_697 (O_697,N_19933,N_19851);
nor UO_698 (O_698,N_19871,N_19944);
and UO_699 (O_699,N_19948,N_19848);
or UO_700 (O_700,N_19955,N_19983);
and UO_701 (O_701,N_19855,N_19863);
nor UO_702 (O_702,N_19970,N_19907);
xnor UO_703 (O_703,N_19881,N_19864);
and UO_704 (O_704,N_19856,N_19963);
xor UO_705 (O_705,N_19939,N_19978);
nand UO_706 (O_706,N_19859,N_19964);
nor UO_707 (O_707,N_19843,N_19937);
nand UO_708 (O_708,N_19939,N_19904);
nand UO_709 (O_709,N_19983,N_19998);
and UO_710 (O_710,N_19988,N_19970);
and UO_711 (O_711,N_19879,N_19971);
and UO_712 (O_712,N_19952,N_19919);
xnor UO_713 (O_713,N_19985,N_19881);
nor UO_714 (O_714,N_19896,N_19883);
and UO_715 (O_715,N_19844,N_19893);
nor UO_716 (O_716,N_19927,N_19971);
xnor UO_717 (O_717,N_19927,N_19889);
xnor UO_718 (O_718,N_19869,N_19937);
nand UO_719 (O_719,N_19939,N_19953);
nand UO_720 (O_720,N_19909,N_19867);
nor UO_721 (O_721,N_19996,N_19867);
nand UO_722 (O_722,N_19962,N_19929);
nor UO_723 (O_723,N_19938,N_19861);
and UO_724 (O_724,N_19853,N_19861);
xor UO_725 (O_725,N_19937,N_19859);
nor UO_726 (O_726,N_19905,N_19914);
nor UO_727 (O_727,N_19979,N_19955);
xnor UO_728 (O_728,N_19852,N_19857);
nand UO_729 (O_729,N_19920,N_19994);
and UO_730 (O_730,N_19843,N_19854);
nor UO_731 (O_731,N_19940,N_19986);
nand UO_732 (O_732,N_19928,N_19927);
nor UO_733 (O_733,N_19861,N_19889);
and UO_734 (O_734,N_19995,N_19928);
xnor UO_735 (O_735,N_19975,N_19910);
and UO_736 (O_736,N_19968,N_19955);
nand UO_737 (O_737,N_19957,N_19863);
xnor UO_738 (O_738,N_19854,N_19890);
nor UO_739 (O_739,N_19896,N_19983);
xnor UO_740 (O_740,N_19986,N_19974);
xor UO_741 (O_741,N_19868,N_19987);
and UO_742 (O_742,N_19932,N_19987);
nor UO_743 (O_743,N_19924,N_19968);
nand UO_744 (O_744,N_19891,N_19945);
nand UO_745 (O_745,N_19938,N_19948);
nor UO_746 (O_746,N_19951,N_19938);
and UO_747 (O_747,N_19870,N_19917);
and UO_748 (O_748,N_19937,N_19855);
xor UO_749 (O_749,N_19872,N_19908);
nor UO_750 (O_750,N_19865,N_19915);
xnor UO_751 (O_751,N_19957,N_19970);
nor UO_752 (O_752,N_19914,N_19923);
nand UO_753 (O_753,N_19924,N_19927);
xnor UO_754 (O_754,N_19965,N_19856);
or UO_755 (O_755,N_19917,N_19863);
nand UO_756 (O_756,N_19866,N_19923);
xnor UO_757 (O_757,N_19956,N_19921);
or UO_758 (O_758,N_19854,N_19935);
nand UO_759 (O_759,N_19878,N_19942);
and UO_760 (O_760,N_19840,N_19852);
or UO_761 (O_761,N_19918,N_19994);
xor UO_762 (O_762,N_19941,N_19972);
or UO_763 (O_763,N_19962,N_19915);
xor UO_764 (O_764,N_19840,N_19857);
xnor UO_765 (O_765,N_19981,N_19998);
nand UO_766 (O_766,N_19993,N_19883);
nand UO_767 (O_767,N_19926,N_19905);
xor UO_768 (O_768,N_19965,N_19855);
or UO_769 (O_769,N_19893,N_19872);
nor UO_770 (O_770,N_19871,N_19845);
nor UO_771 (O_771,N_19924,N_19930);
nor UO_772 (O_772,N_19851,N_19919);
xor UO_773 (O_773,N_19903,N_19862);
nand UO_774 (O_774,N_19948,N_19935);
nand UO_775 (O_775,N_19954,N_19922);
nor UO_776 (O_776,N_19964,N_19897);
or UO_777 (O_777,N_19961,N_19866);
and UO_778 (O_778,N_19929,N_19950);
nor UO_779 (O_779,N_19958,N_19920);
or UO_780 (O_780,N_19884,N_19858);
or UO_781 (O_781,N_19872,N_19969);
nor UO_782 (O_782,N_19926,N_19927);
xnor UO_783 (O_783,N_19940,N_19901);
nor UO_784 (O_784,N_19892,N_19986);
nand UO_785 (O_785,N_19856,N_19933);
xor UO_786 (O_786,N_19951,N_19927);
and UO_787 (O_787,N_19946,N_19993);
nand UO_788 (O_788,N_19992,N_19951);
and UO_789 (O_789,N_19941,N_19986);
xor UO_790 (O_790,N_19953,N_19903);
or UO_791 (O_791,N_19899,N_19924);
nor UO_792 (O_792,N_19901,N_19989);
xnor UO_793 (O_793,N_19968,N_19928);
nor UO_794 (O_794,N_19919,N_19899);
or UO_795 (O_795,N_19926,N_19855);
and UO_796 (O_796,N_19953,N_19884);
or UO_797 (O_797,N_19984,N_19962);
nand UO_798 (O_798,N_19959,N_19892);
nand UO_799 (O_799,N_19849,N_19855);
and UO_800 (O_800,N_19981,N_19969);
and UO_801 (O_801,N_19946,N_19895);
xor UO_802 (O_802,N_19964,N_19869);
or UO_803 (O_803,N_19947,N_19865);
nand UO_804 (O_804,N_19950,N_19995);
nand UO_805 (O_805,N_19876,N_19965);
or UO_806 (O_806,N_19935,N_19885);
and UO_807 (O_807,N_19886,N_19910);
xor UO_808 (O_808,N_19911,N_19993);
or UO_809 (O_809,N_19928,N_19903);
and UO_810 (O_810,N_19982,N_19861);
xor UO_811 (O_811,N_19970,N_19903);
nand UO_812 (O_812,N_19859,N_19886);
xnor UO_813 (O_813,N_19945,N_19962);
and UO_814 (O_814,N_19884,N_19882);
and UO_815 (O_815,N_19917,N_19960);
or UO_816 (O_816,N_19892,N_19939);
nor UO_817 (O_817,N_19987,N_19888);
nand UO_818 (O_818,N_19926,N_19973);
xor UO_819 (O_819,N_19962,N_19886);
nor UO_820 (O_820,N_19979,N_19841);
xnor UO_821 (O_821,N_19965,N_19915);
or UO_822 (O_822,N_19962,N_19980);
nor UO_823 (O_823,N_19964,N_19982);
and UO_824 (O_824,N_19906,N_19927);
or UO_825 (O_825,N_19907,N_19964);
and UO_826 (O_826,N_19916,N_19943);
xor UO_827 (O_827,N_19918,N_19877);
nor UO_828 (O_828,N_19894,N_19961);
or UO_829 (O_829,N_19909,N_19864);
or UO_830 (O_830,N_19881,N_19946);
or UO_831 (O_831,N_19916,N_19972);
nand UO_832 (O_832,N_19908,N_19902);
or UO_833 (O_833,N_19987,N_19906);
and UO_834 (O_834,N_19957,N_19920);
or UO_835 (O_835,N_19997,N_19856);
nand UO_836 (O_836,N_19886,N_19852);
xor UO_837 (O_837,N_19954,N_19959);
or UO_838 (O_838,N_19945,N_19859);
nor UO_839 (O_839,N_19955,N_19886);
and UO_840 (O_840,N_19910,N_19962);
xnor UO_841 (O_841,N_19857,N_19926);
or UO_842 (O_842,N_19886,N_19967);
nand UO_843 (O_843,N_19863,N_19885);
xor UO_844 (O_844,N_19980,N_19862);
or UO_845 (O_845,N_19879,N_19917);
xnor UO_846 (O_846,N_19903,N_19891);
and UO_847 (O_847,N_19964,N_19962);
or UO_848 (O_848,N_19901,N_19950);
or UO_849 (O_849,N_19995,N_19938);
nor UO_850 (O_850,N_19991,N_19973);
nand UO_851 (O_851,N_19856,N_19864);
or UO_852 (O_852,N_19845,N_19890);
xnor UO_853 (O_853,N_19906,N_19888);
and UO_854 (O_854,N_19976,N_19911);
nand UO_855 (O_855,N_19869,N_19858);
xor UO_856 (O_856,N_19841,N_19912);
or UO_857 (O_857,N_19950,N_19909);
and UO_858 (O_858,N_19919,N_19900);
nor UO_859 (O_859,N_19877,N_19914);
xor UO_860 (O_860,N_19876,N_19934);
nor UO_861 (O_861,N_19925,N_19960);
nand UO_862 (O_862,N_19882,N_19991);
nor UO_863 (O_863,N_19906,N_19952);
or UO_864 (O_864,N_19844,N_19943);
and UO_865 (O_865,N_19909,N_19873);
xnor UO_866 (O_866,N_19993,N_19992);
and UO_867 (O_867,N_19911,N_19920);
and UO_868 (O_868,N_19880,N_19989);
nand UO_869 (O_869,N_19979,N_19952);
or UO_870 (O_870,N_19922,N_19864);
and UO_871 (O_871,N_19989,N_19878);
or UO_872 (O_872,N_19879,N_19865);
or UO_873 (O_873,N_19928,N_19885);
or UO_874 (O_874,N_19843,N_19974);
xnor UO_875 (O_875,N_19906,N_19855);
and UO_876 (O_876,N_19862,N_19970);
or UO_877 (O_877,N_19915,N_19954);
or UO_878 (O_878,N_19953,N_19888);
and UO_879 (O_879,N_19996,N_19843);
and UO_880 (O_880,N_19938,N_19970);
and UO_881 (O_881,N_19869,N_19916);
xor UO_882 (O_882,N_19918,N_19977);
and UO_883 (O_883,N_19995,N_19994);
nand UO_884 (O_884,N_19912,N_19952);
and UO_885 (O_885,N_19944,N_19891);
or UO_886 (O_886,N_19867,N_19914);
xor UO_887 (O_887,N_19860,N_19861);
or UO_888 (O_888,N_19981,N_19897);
and UO_889 (O_889,N_19890,N_19883);
or UO_890 (O_890,N_19892,N_19917);
nand UO_891 (O_891,N_19952,N_19944);
or UO_892 (O_892,N_19860,N_19842);
nand UO_893 (O_893,N_19985,N_19961);
and UO_894 (O_894,N_19996,N_19972);
nand UO_895 (O_895,N_19957,N_19928);
or UO_896 (O_896,N_19886,N_19985);
nor UO_897 (O_897,N_19973,N_19960);
and UO_898 (O_898,N_19863,N_19936);
nand UO_899 (O_899,N_19895,N_19888);
and UO_900 (O_900,N_19999,N_19915);
and UO_901 (O_901,N_19959,N_19948);
xor UO_902 (O_902,N_19925,N_19958);
xnor UO_903 (O_903,N_19855,N_19955);
and UO_904 (O_904,N_19840,N_19895);
and UO_905 (O_905,N_19845,N_19918);
xor UO_906 (O_906,N_19842,N_19931);
nand UO_907 (O_907,N_19886,N_19937);
xnor UO_908 (O_908,N_19869,N_19994);
or UO_909 (O_909,N_19964,N_19983);
and UO_910 (O_910,N_19899,N_19938);
nand UO_911 (O_911,N_19982,N_19907);
and UO_912 (O_912,N_19892,N_19971);
and UO_913 (O_913,N_19991,N_19847);
nand UO_914 (O_914,N_19954,N_19957);
and UO_915 (O_915,N_19926,N_19939);
nand UO_916 (O_916,N_19885,N_19842);
and UO_917 (O_917,N_19939,N_19895);
xnor UO_918 (O_918,N_19890,N_19977);
nor UO_919 (O_919,N_19924,N_19858);
and UO_920 (O_920,N_19978,N_19901);
xnor UO_921 (O_921,N_19848,N_19873);
and UO_922 (O_922,N_19998,N_19951);
nand UO_923 (O_923,N_19867,N_19955);
nand UO_924 (O_924,N_19983,N_19866);
nand UO_925 (O_925,N_19962,N_19858);
or UO_926 (O_926,N_19939,N_19871);
or UO_927 (O_927,N_19913,N_19900);
xor UO_928 (O_928,N_19950,N_19884);
or UO_929 (O_929,N_19967,N_19958);
nor UO_930 (O_930,N_19987,N_19870);
xor UO_931 (O_931,N_19928,N_19874);
or UO_932 (O_932,N_19993,N_19884);
nand UO_933 (O_933,N_19898,N_19870);
nand UO_934 (O_934,N_19934,N_19853);
or UO_935 (O_935,N_19914,N_19998);
nand UO_936 (O_936,N_19961,N_19897);
xnor UO_937 (O_937,N_19933,N_19873);
or UO_938 (O_938,N_19867,N_19847);
xor UO_939 (O_939,N_19841,N_19863);
nand UO_940 (O_940,N_19867,N_19892);
nand UO_941 (O_941,N_19939,N_19909);
xnor UO_942 (O_942,N_19844,N_19871);
nand UO_943 (O_943,N_19912,N_19931);
nand UO_944 (O_944,N_19976,N_19842);
nor UO_945 (O_945,N_19933,N_19957);
or UO_946 (O_946,N_19922,N_19902);
nand UO_947 (O_947,N_19919,N_19898);
nand UO_948 (O_948,N_19974,N_19846);
xnor UO_949 (O_949,N_19948,N_19985);
xnor UO_950 (O_950,N_19999,N_19979);
and UO_951 (O_951,N_19842,N_19963);
and UO_952 (O_952,N_19982,N_19987);
or UO_953 (O_953,N_19987,N_19949);
nand UO_954 (O_954,N_19974,N_19892);
nor UO_955 (O_955,N_19859,N_19867);
nor UO_956 (O_956,N_19905,N_19907);
nand UO_957 (O_957,N_19997,N_19846);
nor UO_958 (O_958,N_19996,N_19848);
nor UO_959 (O_959,N_19871,N_19963);
nor UO_960 (O_960,N_19989,N_19852);
xor UO_961 (O_961,N_19953,N_19898);
nand UO_962 (O_962,N_19898,N_19851);
nand UO_963 (O_963,N_19882,N_19894);
or UO_964 (O_964,N_19888,N_19945);
nand UO_965 (O_965,N_19917,N_19991);
or UO_966 (O_966,N_19882,N_19924);
xnor UO_967 (O_967,N_19989,N_19973);
nand UO_968 (O_968,N_19957,N_19925);
xnor UO_969 (O_969,N_19944,N_19969);
nand UO_970 (O_970,N_19968,N_19962);
nand UO_971 (O_971,N_19947,N_19970);
xor UO_972 (O_972,N_19848,N_19900);
xnor UO_973 (O_973,N_19933,N_19864);
or UO_974 (O_974,N_19860,N_19885);
nand UO_975 (O_975,N_19950,N_19955);
and UO_976 (O_976,N_19894,N_19970);
and UO_977 (O_977,N_19978,N_19886);
and UO_978 (O_978,N_19981,N_19951);
or UO_979 (O_979,N_19994,N_19986);
or UO_980 (O_980,N_19874,N_19960);
xor UO_981 (O_981,N_19907,N_19843);
nand UO_982 (O_982,N_19993,N_19866);
xor UO_983 (O_983,N_19969,N_19903);
and UO_984 (O_984,N_19994,N_19972);
xor UO_985 (O_985,N_19862,N_19958);
or UO_986 (O_986,N_19920,N_19940);
or UO_987 (O_987,N_19953,N_19943);
or UO_988 (O_988,N_19913,N_19861);
or UO_989 (O_989,N_19843,N_19964);
nand UO_990 (O_990,N_19867,N_19972);
or UO_991 (O_991,N_19859,N_19902);
xnor UO_992 (O_992,N_19878,N_19903);
nor UO_993 (O_993,N_19869,N_19981);
nor UO_994 (O_994,N_19934,N_19914);
nor UO_995 (O_995,N_19894,N_19935);
xor UO_996 (O_996,N_19951,N_19903);
or UO_997 (O_997,N_19980,N_19894);
or UO_998 (O_998,N_19918,N_19842);
nand UO_999 (O_999,N_19963,N_19971);
or UO_1000 (O_1000,N_19971,N_19904);
xor UO_1001 (O_1001,N_19915,N_19956);
or UO_1002 (O_1002,N_19936,N_19930);
nand UO_1003 (O_1003,N_19851,N_19878);
and UO_1004 (O_1004,N_19887,N_19858);
xor UO_1005 (O_1005,N_19897,N_19989);
and UO_1006 (O_1006,N_19935,N_19984);
nand UO_1007 (O_1007,N_19848,N_19932);
nor UO_1008 (O_1008,N_19848,N_19971);
xnor UO_1009 (O_1009,N_19880,N_19933);
nand UO_1010 (O_1010,N_19927,N_19954);
or UO_1011 (O_1011,N_19980,N_19935);
nor UO_1012 (O_1012,N_19972,N_19880);
nand UO_1013 (O_1013,N_19896,N_19902);
and UO_1014 (O_1014,N_19960,N_19944);
nor UO_1015 (O_1015,N_19998,N_19896);
xor UO_1016 (O_1016,N_19907,N_19860);
and UO_1017 (O_1017,N_19922,N_19972);
and UO_1018 (O_1018,N_19918,N_19896);
or UO_1019 (O_1019,N_19854,N_19864);
xor UO_1020 (O_1020,N_19937,N_19875);
xor UO_1021 (O_1021,N_19957,N_19984);
xnor UO_1022 (O_1022,N_19941,N_19905);
nor UO_1023 (O_1023,N_19995,N_19910);
or UO_1024 (O_1024,N_19891,N_19847);
xor UO_1025 (O_1025,N_19893,N_19922);
nand UO_1026 (O_1026,N_19862,N_19926);
nor UO_1027 (O_1027,N_19882,N_19995);
xnor UO_1028 (O_1028,N_19872,N_19992);
xor UO_1029 (O_1029,N_19859,N_19866);
or UO_1030 (O_1030,N_19861,N_19896);
nor UO_1031 (O_1031,N_19920,N_19991);
or UO_1032 (O_1032,N_19876,N_19948);
and UO_1033 (O_1033,N_19988,N_19850);
xor UO_1034 (O_1034,N_19996,N_19960);
or UO_1035 (O_1035,N_19947,N_19866);
xor UO_1036 (O_1036,N_19961,N_19968);
xnor UO_1037 (O_1037,N_19870,N_19851);
nand UO_1038 (O_1038,N_19934,N_19954);
xor UO_1039 (O_1039,N_19854,N_19996);
or UO_1040 (O_1040,N_19953,N_19977);
nor UO_1041 (O_1041,N_19899,N_19849);
xnor UO_1042 (O_1042,N_19946,N_19986);
nor UO_1043 (O_1043,N_19859,N_19856);
nand UO_1044 (O_1044,N_19915,N_19979);
or UO_1045 (O_1045,N_19965,N_19992);
and UO_1046 (O_1046,N_19969,N_19880);
nand UO_1047 (O_1047,N_19965,N_19930);
and UO_1048 (O_1048,N_19868,N_19970);
and UO_1049 (O_1049,N_19895,N_19970);
xor UO_1050 (O_1050,N_19902,N_19863);
xor UO_1051 (O_1051,N_19885,N_19891);
xor UO_1052 (O_1052,N_19849,N_19929);
and UO_1053 (O_1053,N_19973,N_19865);
or UO_1054 (O_1054,N_19954,N_19870);
xnor UO_1055 (O_1055,N_19986,N_19999);
nor UO_1056 (O_1056,N_19853,N_19848);
xor UO_1057 (O_1057,N_19966,N_19860);
or UO_1058 (O_1058,N_19917,N_19982);
or UO_1059 (O_1059,N_19982,N_19986);
or UO_1060 (O_1060,N_19904,N_19991);
or UO_1061 (O_1061,N_19861,N_19962);
xnor UO_1062 (O_1062,N_19943,N_19992);
xor UO_1063 (O_1063,N_19994,N_19971);
or UO_1064 (O_1064,N_19853,N_19930);
or UO_1065 (O_1065,N_19852,N_19865);
nor UO_1066 (O_1066,N_19893,N_19850);
nor UO_1067 (O_1067,N_19953,N_19902);
xor UO_1068 (O_1068,N_19917,N_19992);
nand UO_1069 (O_1069,N_19860,N_19971);
or UO_1070 (O_1070,N_19901,N_19957);
nand UO_1071 (O_1071,N_19932,N_19989);
and UO_1072 (O_1072,N_19918,N_19914);
xor UO_1073 (O_1073,N_19914,N_19870);
or UO_1074 (O_1074,N_19884,N_19905);
nor UO_1075 (O_1075,N_19966,N_19869);
or UO_1076 (O_1076,N_19987,N_19977);
nand UO_1077 (O_1077,N_19853,N_19844);
nand UO_1078 (O_1078,N_19970,N_19984);
xnor UO_1079 (O_1079,N_19939,N_19856);
nand UO_1080 (O_1080,N_19999,N_19929);
nor UO_1081 (O_1081,N_19861,N_19989);
nor UO_1082 (O_1082,N_19989,N_19864);
or UO_1083 (O_1083,N_19884,N_19967);
or UO_1084 (O_1084,N_19853,N_19973);
or UO_1085 (O_1085,N_19977,N_19869);
xnor UO_1086 (O_1086,N_19983,N_19946);
xor UO_1087 (O_1087,N_19926,N_19851);
and UO_1088 (O_1088,N_19973,N_19981);
and UO_1089 (O_1089,N_19873,N_19943);
or UO_1090 (O_1090,N_19843,N_19960);
or UO_1091 (O_1091,N_19994,N_19929);
nor UO_1092 (O_1092,N_19894,N_19974);
nand UO_1093 (O_1093,N_19990,N_19945);
nor UO_1094 (O_1094,N_19914,N_19909);
xor UO_1095 (O_1095,N_19986,N_19952);
xnor UO_1096 (O_1096,N_19906,N_19982);
nand UO_1097 (O_1097,N_19999,N_19993);
xnor UO_1098 (O_1098,N_19952,N_19865);
or UO_1099 (O_1099,N_19898,N_19952);
and UO_1100 (O_1100,N_19904,N_19941);
nor UO_1101 (O_1101,N_19865,N_19895);
and UO_1102 (O_1102,N_19900,N_19869);
nand UO_1103 (O_1103,N_19979,N_19888);
xnor UO_1104 (O_1104,N_19841,N_19919);
nand UO_1105 (O_1105,N_19930,N_19899);
or UO_1106 (O_1106,N_19998,N_19879);
and UO_1107 (O_1107,N_19857,N_19932);
and UO_1108 (O_1108,N_19906,N_19905);
nor UO_1109 (O_1109,N_19911,N_19909);
nand UO_1110 (O_1110,N_19913,N_19970);
or UO_1111 (O_1111,N_19840,N_19971);
or UO_1112 (O_1112,N_19951,N_19925);
and UO_1113 (O_1113,N_19947,N_19904);
and UO_1114 (O_1114,N_19888,N_19870);
or UO_1115 (O_1115,N_19946,N_19982);
and UO_1116 (O_1116,N_19948,N_19971);
nand UO_1117 (O_1117,N_19979,N_19917);
xnor UO_1118 (O_1118,N_19966,N_19848);
nand UO_1119 (O_1119,N_19971,N_19953);
and UO_1120 (O_1120,N_19847,N_19872);
nor UO_1121 (O_1121,N_19977,N_19928);
xor UO_1122 (O_1122,N_19879,N_19956);
or UO_1123 (O_1123,N_19994,N_19858);
and UO_1124 (O_1124,N_19967,N_19978);
nand UO_1125 (O_1125,N_19873,N_19919);
and UO_1126 (O_1126,N_19944,N_19867);
and UO_1127 (O_1127,N_19924,N_19884);
xnor UO_1128 (O_1128,N_19909,N_19906);
nor UO_1129 (O_1129,N_19909,N_19863);
or UO_1130 (O_1130,N_19975,N_19841);
and UO_1131 (O_1131,N_19894,N_19907);
and UO_1132 (O_1132,N_19934,N_19881);
nor UO_1133 (O_1133,N_19980,N_19998);
or UO_1134 (O_1134,N_19910,N_19915);
and UO_1135 (O_1135,N_19933,N_19926);
and UO_1136 (O_1136,N_19932,N_19841);
nor UO_1137 (O_1137,N_19958,N_19971);
and UO_1138 (O_1138,N_19869,N_19984);
xnor UO_1139 (O_1139,N_19981,N_19929);
nand UO_1140 (O_1140,N_19958,N_19954);
nand UO_1141 (O_1141,N_19920,N_19965);
xor UO_1142 (O_1142,N_19982,N_19945);
xor UO_1143 (O_1143,N_19980,N_19939);
nor UO_1144 (O_1144,N_19999,N_19925);
nand UO_1145 (O_1145,N_19994,N_19891);
xor UO_1146 (O_1146,N_19854,N_19872);
and UO_1147 (O_1147,N_19854,N_19928);
and UO_1148 (O_1148,N_19958,N_19901);
or UO_1149 (O_1149,N_19960,N_19896);
or UO_1150 (O_1150,N_19990,N_19954);
or UO_1151 (O_1151,N_19859,N_19908);
or UO_1152 (O_1152,N_19915,N_19940);
and UO_1153 (O_1153,N_19981,N_19889);
nor UO_1154 (O_1154,N_19880,N_19857);
xor UO_1155 (O_1155,N_19999,N_19932);
nand UO_1156 (O_1156,N_19981,N_19847);
nor UO_1157 (O_1157,N_19907,N_19947);
or UO_1158 (O_1158,N_19932,N_19891);
or UO_1159 (O_1159,N_19847,N_19886);
nor UO_1160 (O_1160,N_19843,N_19963);
and UO_1161 (O_1161,N_19899,N_19879);
or UO_1162 (O_1162,N_19884,N_19922);
nand UO_1163 (O_1163,N_19979,N_19870);
and UO_1164 (O_1164,N_19920,N_19874);
and UO_1165 (O_1165,N_19879,N_19850);
nand UO_1166 (O_1166,N_19978,N_19992);
and UO_1167 (O_1167,N_19973,N_19995);
nor UO_1168 (O_1168,N_19896,N_19917);
or UO_1169 (O_1169,N_19864,N_19887);
or UO_1170 (O_1170,N_19946,N_19862);
and UO_1171 (O_1171,N_19927,N_19841);
and UO_1172 (O_1172,N_19914,N_19943);
and UO_1173 (O_1173,N_19960,N_19841);
nor UO_1174 (O_1174,N_19974,N_19919);
nand UO_1175 (O_1175,N_19897,N_19974);
nor UO_1176 (O_1176,N_19958,N_19974);
nand UO_1177 (O_1177,N_19914,N_19895);
nor UO_1178 (O_1178,N_19914,N_19926);
and UO_1179 (O_1179,N_19992,N_19869);
nor UO_1180 (O_1180,N_19896,N_19934);
and UO_1181 (O_1181,N_19870,N_19896);
nor UO_1182 (O_1182,N_19882,N_19896);
xor UO_1183 (O_1183,N_19921,N_19946);
or UO_1184 (O_1184,N_19938,N_19911);
nor UO_1185 (O_1185,N_19949,N_19884);
or UO_1186 (O_1186,N_19859,N_19930);
nor UO_1187 (O_1187,N_19901,N_19924);
and UO_1188 (O_1188,N_19989,N_19892);
nor UO_1189 (O_1189,N_19909,N_19945);
and UO_1190 (O_1190,N_19954,N_19844);
nor UO_1191 (O_1191,N_19878,N_19890);
and UO_1192 (O_1192,N_19939,N_19879);
or UO_1193 (O_1193,N_19876,N_19895);
and UO_1194 (O_1194,N_19967,N_19859);
xnor UO_1195 (O_1195,N_19924,N_19895);
nand UO_1196 (O_1196,N_19927,N_19852);
xnor UO_1197 (O_1197,N_19930,N_19912);
nor UO_1198 (O_1198,N_19966,N_19878);
xor UO_1199 (O_1199,N_19969,N_19949);
xnor UO_1200 (O_1200,N_19992,N_19863);
nor UO_1201 (O_1201,N_19959,N_19961);
and UO_1202 (O_1202,N_19940,N_19848);
or UO_1203 (O_1203,N_19932,N_19935);
nor UO_1204 (O_1204,N_19958,N_19918);
and UO_1205 (O_1205,N_19919,N_19935);
xor UO_1206 (O_1206,N_19942,N_19883);
nor UO_1207 (O_1207,N_19965,N_19914);
and UO_1208 (O_1208,N_19897,N_19927);
and UO_1209 (O_1209,N_19934,N_19948);
or UO_1210 (O_1210,N_19984,N_19973);
or UO_1211 (O_1211,N_19972,N_19944);
nor UO_1212 (O_1212,N_19932,N_19940);
nor UO_1213 (O_1213,N_19903,N_19952);
or UO_1214 (O_1214,N_19937,N_19984);
xnor UO_1215 (O_1215,N_19980,N_19895);
nand UO_1216 (O_1216,N_19986,N_19882);
nor UO_1217 (O_1217,N_19840,N_19889);
or UO_1218 (O_1218,N_19860,N_19873);
and UO_1219 (O_1219,N_19885,N_19851);
nand UO_1220 (O_1220,N_19993,N_19904);
nand UO_1221 (O_1221,N_19919,N_19916);
nor UO_1222 (O_1222,N_19874,N_19919);
xnor UO_1223 (O_1223,N_19997,N_19980);
nand UO_1224 (O_1224,N_19936,N_19944);
or UO_1225 (O_1225,N_19937,N_19963);
and UO_1226 (O_1226,N_19876,N_19853);
nor UO_1227 (O_1227,N_19866,N_19991);
nand UO_1228 (O_1228,N_19912,N_19867);
nand UO_1229 (O_1229,N_19892,N_19973);
xnor UO_1230 (O_1230,N_19901,N_19997);
nor UO_1231 (O_1231,N_19978,N_19862);
xnor UO_1232 (O_1232,N_19990,N_19887);
nand UO_1233 (O_1233,N_19957,N_19989);
nor UO_1234 (O_1234,N_19957,N_19996);
or UO_1235 (O_1235,N_19883,N_19949);
nand UO_1236 (O_1236,N_19966,N_19905);
and UO_1237 (O_1237,N_19902,N_19883);
and UO_1238 (O_1238,N_19842,N_19892);
or UO_1239 (O_1239,N_19924,N_19923);
nand UO_1240 (O_1240,N_19931,N_19868);
nor UO_1241 (O_1241,N_19933,N_19935);
or UO_1242 (O_1242,N_19882,N_19869);
xor UO_1243 (O_1243,N_19843,N_19888);
and UO_1244 (O_1244,N_19996,N_19850);
nand UO_1245 (O_1245,N_19921,N_19996);
and UO_1246 (O_1246,N_19941,N_19864);
nand UO_1247 (O_1247,N_19896,N_19948);
or UO_1248 (O_1248,N_19896,N_19846);
or UO_1249 (O_1249,N_19945,N_19866);
or UO_1250 (O_1250,N_19869,N_19938);
nand UO_1251 (O_1251,N_19960,N_19869);
or UO_1252 (O_1252,N_19965,N_19970);
or UO_1253 (O_1253,N_19901,N_19971);
nor UO_1254 (O_1254,N_19960,N_19902);
nand UO_1255 (O_1255,N_19896,N_19989);
xnor UO_1256 (O_1256,N_19880,N_19963);
and UO_1257 (O_1257,N_19849,N_19856);
nand UO_1258 (O_1258,N_19997,N_19975);
or UO_1259 (O_1259,N_19958,N_19994);
xor UO_1260 (O_1260,N_19853,N_19920);
xnor UO_1261 (O_1261,N_19948,N_19987);
or UO_1262 (O_1262,N_19977,N_19942);
nor UO_1263 (O_1263,N_19852,N_19961);
xnor UO_1264 (O_1264,N_19993,N_19974);
nand UO_1265 (O_1265,N_19914,N_19924);
nor UO_1266 (O_1266,N_19851,N_19990);
or UO_1267 (O_1267,N_19894,N_19841);
or UO_1268 (O_1268,N_19998,N_19859);
nor UO_1269 (O_1269,N_19841,N_19935);
and UO_1270 (O_1270,N_19891,N_19968);
and UO_1271 (O_1271,N_19965,N_19981);
nor UO_1272 (O_1272,N_19867,N_19963);
and UO_1273 (O_1273,N_19949,N_19939);
and UO_1274 (O_1274,N_19885,N_19924);
xor UO_1275 (O_1275,N_19849,N_19944);
nand UO_1276 (O_1276,N_19847,N_19916);
xnor UO_1277 (O_1277,N_19888,N_19896);
xnor UO_1278 (O_1278,N_19935,N_19996);
nand UO_1279 (O_1279,N_19952,N_19920);
or UO_1280 (O_1280,N_19864,N_19951);
or UO_1281 (O_1281,N_19916,N_19917);
and UO_1282 (O_1282,N_19948,N_19901);
nor UO_1283 (O_1283,N_19991,N_19961);
or UO_1284 (O_1284,N_19994,N_19934);
nor UO_1285 (O_1285,N_19935,N_19857);
and UO_1286 (O_1286,N_19942,N_19957);
xnor UO_1287 (O_1287,N_19974,N_19998);
xor UO_1288 (O_1288,N_19912,N_19955);
and UO_1289 (O_1289,N_19956,N_19858);
nand UO_1290 (O_1290,N_19994,N_19874);
xnor UO_1291 (O_1291,N_19857,N_19866);
nand UO_1292 (O_1292,N_19904,N_19891);
nor UO_1293 (O_1293,N_19842,N_19961);
and UO_1294 (O_1294,N_19957,N_19971);
nor UO_1295 (O_1295,N_19893,N_19891);
nand UO_1296 (O_1296,N_19921,N_19878);
nor UO_1297 (O_1297,N_19915,N_19846);
or UO_1298 (O_1298,N_19856,N_19869);
and UO_1299 (O_1299,N_19941,N_19930);
xor UO_1300 (O_1300,N_19866,N_19930);
nand UO_1301 (O_1301,N_19914,N_19859);
or UO_1302 (O_1302,N_19919,N_19917);
xor UO_1303 (O_1303,N_19954,N_19985);
nand UO_1304 (O_1304,N_19976,N_19962);
nand UO_1305 (O_1305,N_19998,N_19910);
or UO_1306 (O_1306,N_19962,N_19928);
nor UO_1307 (O_1307,N_19991,N_19842);
xnor UO_1308 (O_1308,N_19954,N_19989);
nor UO_1309 (O_1309,N_19991,N_19945);
nand UO_1310 (O_1310,N_19958,N_19936);
xor UO_1311 (O_1311,N_19971,N_19928);
nor UO_1312 (O_1312,N_19886,N_19898);
nor UO_1313 (O_1313,N_19987,N_19991);
nor UO_1314 (O_1314,N_19983,N_19936);
or UO_1315 (O_1315,N_19911,N_19918);
nand UO_1316 (O_1316,N_19955,N_19958);
and UO_1317 (O_1317,N_19976,N_19974);
xor UO_1318 (O_1318,N_19966,N_19963);
xor UO_1319 (O_1319,N_19860,N_19997);
or UO_1320 (O_1320,N_19873,N_19929);
xnor UO_1321 (O_1321,N_19859,N_19862);
or UO_1322 (O_1322,N_19912,N_19985);
xnor UO_1323 (O_1323,N_19965,N_19868);
or UO_1324 (O_1324,N_19996,N_19914);
nor UO_1325 (O_1325,N_19847,N_19936);
or UO_1326 (O_1326,N_19912,N_19948);
or UO_1327 (O_1327,N_19909,N_19919);
nand UO_1328 (O_1328,N_19934,N_19951);
nand UO_1329 (O_1329,N_19851,N_19869);
nand UO_1330 (O_1330,N_19901,N_19970);
and UO_1331 (O_1331,N_19855,N_19997);
and UO_1332 (O_1332,N_19981,N_19927);
nor UO_1333 (O_1333,N_19878,N_19992);
and UO_1334 (O_1334,N_19978,N_19935);
xor UO_1335 (O_1335,N_19992,N_19883);
nand UO_1336 (O_1336,N_19924,N_19993);
or UO_1337 (O_1337,N_19994,N_19985);
and UO_1338 (O_1338,N_19958,N_19859);
or UO_1339 (O_1339,N_19995,N_19975);
xor UO_1340 (O_1340,N_19989,N_19930);
and UO_1341 (O_1341,N_19922,N_19895);
nand UO_1342 (O_1342,N_19943,N_19960);
or UO_1343 (O_1343,N_19943,N_19981);
and UO_1344 (O_1344,N_19968,N_19892);
xnor UO_1345 (O_1345,N_19930,N_19856);
nor UO_1346 (O_1346,N_19937,N_19919);
xor UO_1347 (O_1347,N_19968,N_19883);
nand UO_1348 (O_1348,N_19990,N_19919);
nor UO_1349 (O_1349,N_19937,N_19961);
and UO_1350 (O_1350,N_19841,N_19959);
xor UO_1351 (O_1351,N_19852,N_19922);
or UO_1352 (O_1352,N_19977,N_19920);
and UO_1353 (O_1353,N_19962,N_19973);
xnor UO_1354 (O_1354,N_19969,N_19914);
xor UO_1355 (O_1355,N_19987,N_19983);
and UO_1356 (O_1356,N_19866,N_19994);
xnor UO_1357 (O_1357,N_19936,N_19949);
xor UO_1358 (O_1358,N_19917,N_19903);
nand UO_1359 (O_1359,N_19853,N_19898);
nor UO_1360 (O_1360,N_19852,N_19861);
and UO_1361 (O_1361,N_19939,N_19932);
nand UO_1362 (O_1362,N_19901,N_19928);
xnor UO_1363 (O_1363,N_19970,N_19877);
xnor UO_1364 (O_1364,N_19991,N_19899);
xor UO_1365 (O_1365,N_19856,N_19988);
nand UO_1366 (O_1366,N_19872,N_19956);
nor UO_1367 (O_1367,N_19893,N_19980);
and UO_1368 (O_1368,N_19850,N_19983);
or UO_1369 (O_1369,N_19949,N_19992);
or UO_1370 (O_1370,N_19889,N_19919);
nand UO_1371 (O_1371,N_19939,N_19992);
nor UO_1372 (O_1372,N_19962,N_19873);
nor UO_1373 (O_1373,N_19912,N_19964);
xor UO_1374 (O_1374,N_19967,N_19994);
or UO_1375 (O_1375,N_19933,N_19949);
nand UO_1376 (O_1376,N_19950,N_19848);
or UO_1377 (O_1377,N_19936,N_19910);
nand UO_1378 (O_1378,N_19844,N_19923);
xnor UO_1379 (O_1379,N_19954,N_19963);
xnor UO_1380 (O_1380,N_19997,N_19999);
and UO_1381 (O_1381,N_19935,N_19905);
nand UO_1382 (O_1382,N_19881,N_19877);
or UO_1383 (O_1383,N_19841,N_19908);
xor UO_1384 (O_1384,N_19995,N_19885);
nand UO_1385 (O_1385,N_19940,N_19998);
nand UO_1386 (O_1386,N_19938,N_19957);
xor UO_1387 (O_1387,N_19959,N_19955);
nor UO_1388 (O_1388,N_19894,N_19893);
and UO_1389 (O_1389,N_19843,N_19876);
and UO_1390 (O_1390,N_19918,N_19853);
and UO_1391 (O_1391,N_19872,N_19910);
and UO_1392 (O_1392,N_19946,N_19870);
nand UO_1393 (O_1393,N_19977,N_19840);
or UO_1394 (O_1394,N_19892,N_19914);
xor UO_1395 (O_1395,N_19981,N_19902);
nand UO_1396 (O_1396,N_19880,N_19866);
nor UO_1397 (O_1397,N_19949,N_19957);
xnor UO_1398 (O_1398,N_19961,N_19979);
and UO_1399 (O_1399,N_19875,N_19892);
or UO_1400 (O_1400,N_19927,N_19891);
or UO_1401 (O_1401,N_19936,N_19992);
and UO_1402 (O_1402,N_19894,N_19876);
and UO_1403 (O_1403,N_19915,N_19881);
and UO_1404 (O_1404,N_19866,N_19864);
or UO_1405 (O_1405,N_19987,N_19862);
nand UO_1406 (O_1406,N_19901,N_19916);
and UO_1407 (O_1407,N_19986,N_19865);
nor UO_1408 (O_1408,N_19911,N_19996);
nand UO_1409 (O_1409,N_19965,N_19889);
nand UO_1410 (O_1410,N_19925,N_19893);
xor UO_1411 (O_1411,N_19930,N_19887);
and UO_1412 (O_1412,N_19971,N_19883);
and UO_1413 (O_1413,N_19929,N_19866);
or UO_1414 (O_1414,N_19968,N_19983);
and UO_1415 (O_1415,N_19990,N_19860);
or UO_1416 (O_1416,N_19908,N_19949);
xnor UO_1417 (O_1417,N_19994,N_19846);
nand UO_1418 (O_1418,N_19877,N_19945);
or UO_1419 (O_1419,N_19985,N_19888);
and UO_1420 (O_1420,N_19908,N_19942);
and UO_1421 (O_1421,N_19860,N_19863);
and UO_1422 (O_1422,N_19981,N_19972);
or UO_1423 (O_1423,N_19880,N_19957);
xor UO_1424 (O_1424,N_19849,N_19863);
nor UO_1425 (O_1425,N_19872,N_19871);
and UO_1426 (O_1426,N_19949,N_19940);
and UO_1427 (O_1427,N_19990,N_19953);
or UO_1428 (O_1428,N_19863,N_19845);
and UO_1429 (O_1429,N_19931,N_19853);
or UO_1430 (O_1430,N_19987,N_19963);
and UO_1431 (O_1431,N_19916,N_19998);
nor UO_1432 (O_1432,N_19950,N_19842);
nand UO_1433 (O_1433,N_19994,N_19938);
or UO_1434 (O_1434,N_19946,N_19849);
nand UO_1435 (O_1435,N_19964,N_19974);
nor UO_1436 (O_1436,N_19977,N_19916);
nand UO_1437 (O_1437,N_19910,N_19905);
nand UO_1438 (O_1438,N_19931,N_19945);
and UO_1439 (O_1439,N_19914,N_19865);
xnor UO_1440 (O_1440,N_19996,N_19983);
and UO_1441 (O_1441,N_19906,N_19965);
xor UO_1442 (O_1442,N_19924,N_19970);
nand UO_1443 (O_1443,N_19960,N_19885);
and UO_1444 (O_1444,N_19964,N_19956);
xor UO_1445 (O_1445,N_19998,N_19881);
nand UO_1446 (O_1446,N_19949,N_19881);
xnor UO_1447 (O_1447,N_19991,N_19958);
nor UO_1448 (O_1448,N_19954,N_19901);
or UO_1449 (O_1449,N_19899,N_19912);
xnor UO_1450 (O_1450,N_19877,N_19862);
nand UO_1451 (O_1451,N_19949,N_19871);
and UO_1452 (O_1452,N_19843,N_19980);
xnor UO_1453 (O_1453,N_19885,N_19996);
nor UO_1454 (O_1454,N_19853,N_19888);
nor UO_1455 (O_1455,N_19981,N_19894);
nor UO_1456 (O_1456,N_19901,N_19851);
and UO_1457 (O_1457,N_19939,N_19942);
and UO_1458 (O_1458,N_19929,N_19953);
and UO_1459 (O_1459,N_19855,N_19983);
nor UO_1460 (O_1460,N_19949,N_19902);
and UO_1461 (O_1461,N_19977,N_19887);
and UO_1462 (O_1462,N_19990,N_19943);
nor UO_1463 (O_1463,N_19910,N_19942);
nand UO_1464 (O_1464,N_19900,N_19956);
and UO_1465 (O_1465,N_19882,N_19846);
nor UO_1466 (O_1466,N_19861,N_19936);
or UO_1467 (O_1467,N_19995,N_19896);
nand UO_1468 (O_1468,N_19939,N_19999);
xor UO_1469 (O_1469,N_19891,N_19841);
and UO_1470 (O_1470,N_19970,N_19850);
and UO_1471 (O_1471,N_19973,N_19895);
nor UO_1472 (O_1472,N_19908,N_19990);
or UO_1473 (O_1473,N_19899,N_19890);
nor UO_1474 (O_1474,N_19891,N_19905);
xnor UO_1475 (O_1475,N_19873,N_19875);
nand UO_1476 (O_1476,N_19988,N_19925);
xor UO_1477 (O_1477,N_19841,N_19985);
nand UO_1478 (O_1478,N_19978,N_19933);
nor UO_1479 (O_1479,N_19927,N_19846);
nor UO_1480 (O_1480,N_19904,N_19968);
and UO_1481 (O_1481,N_19892,N_19863);
nand UO_1482 (O_1482,N_19930,N_19865);
xnor UO_1483 (O_1483,N_19988,N_19962);
or UO_1484 (O_1484,N_19852,N_19910);
nand UO_1485 (O_1485,N_19993,N_19976);
and UO_1486 (O_1486,N_19933,N_19996);
or UO_1487 (O_1487,N_19892,N_19884);
or UO_1488 (O_1488,N_19936,N_19840);
nor UO_1489 (O_1489,N_19878,N_19884);
xor UO_1490 (O_1490,N_19899,N_19937);
nor UO_1491 (O_1491,N_19859,N_19887);
nand UO_1492 (O_1492,N_19863,N_19854);
nand UO_1493 (O_1493,N_19870,N_19857);
and UO_1494 (O_1494,N_19948,N_19965);
xnor UO_1495 (O_1495,N_19911,N_19947);
and UO_1496 (O_1496,N_19909,N_19991);
or UO_1497 (O_1497,N_19841,N_19922);
nand UO_1498 (O_1498,N_19936,N_19875);
nand UO_1499 (O_1499,N_19887,N_19913);
nor UO_1500 (O_1500,N_19962,N_19881);
nor UO_1501 (O_1501,N_19943,N_19961);
or UO_1502 (O_1502,N_19854,N_19989);
nand UO_1503 (O_1503,N_19926,N_19994);
and UO_1504 (O_1504,N_19973,N_19893);
and UO_1505 (O_1505,N_19930,N_19933);
nor UO_1506 (O_1506,N_19860,N_19890);
nand UO_1507 (O_1507,N_19852,N_19925);
nor UO_1508 (O_1508,N_19873,N_19974);
xnor UO_1509 (O_1509,N_19865,N_19970);
or UO_1510 (O_1510,N_19953,N_19930);
or UO_1511 (O_1511,N_19877,N_19988);
or UO_1512 (O_1512,N_19863,N_19905);
nand UO_1513 (O_1513,N_19901,N_19942);
nor UO_1514 (O_1514,N_19943,N_19978);
and UO_1515 (O_1515,N_19872,N_19866);
or UO_1516 (O_1516,N_19856,N_19907);
or UO_1517 (O_1517,N_19924,N_19940);
or UO_1518 (O_1518,N_19850,N_19914);
or UO_1519 (O_1519,N_19897,N_19912);
xnor UO_1520 (O_1520,N_19894,N_19950);
and UO_1521 (O_1521,N_19868,N_19991);
and UO_1522 (O_1522,N_19870,N_19874);
and UO_1523 (O_1523,N_19850,N_19995);
xnor UO_1524 (O_1524,N_19888,N_19889);
nand UO_1525 (O_1525,N_19849,N_19935);
nor UO_1526 (O_1526,N_19986,N_19992);
xnor UO_1527 (O_1527,N_19883,N_19877);
and UO_1528 (O_1528,N_19986,N_19958);
and UO_1529 (O_1529,N_19954,N_19894);
or UO_1530 (O_1530,N_19849,N_19966);
nor UO_1531 (O_1531,N_19933,N_19939);
xnor UO_1532 (O_1532,N_19924,N_19900);
nor UO_1533 (O_1533,N_19975,N_19879);
nand UO_1534 (O_1534,N_19989,N_19849);
and UO_1535 (O_1535,N_19857,N_19987);
nand UO_1536 (O_1536,N_19893,N_19991);
xor UO_1537 (O_1537,N_19975,N_19958);
or UO_1538 (O_1538,N_19974,N_19901);
nand UO_1539 (O_1539,N_19861,N_19845);
xnor UO_1540 (O_1540,N_19933,N_19990);
nor UO_1541 (O_1541,N_19874,N_19907);
or UO_1542 (O_1542,N_19941,N_19847);
nor UO_1543 (O_1543,N_19968,N_19912);
or UO_1544 (O_1544,N_19946,N_19973);
nand UO_1545 (O_1545,N_19880,N_19879);
or UO_1546 (O_1546,N_19896,N_19851);
nor UO_1547 (O_1547,N_19890,N_19933);
nand UO_1548 (O_1548,N_19894,N_19945);
and UO_1549 (O_1549,N_19982,N_19997);
xnor UO_1550 (O_1550,N_19998,N_19935);
nor UO_1551 (O_1551,N_19867,N_19973);
nand UO_1552 (O_1552,N_19844,N_19900);
nand UO_1553 (O_1553,N_19983,N_19972);
xnor UO_1554 (O_1554,N_19974,N_19987);
nand UO_1555 (O_1555,N_19982,N_19846);
nor UO_1556 (O_1556,N_19976,N_19863);
or UO_1557 (O_1557,N_19928,N_19973);
nor UO_1558 (O_1558,N_19944,N_19859);
xnor UO_1559 (O_1559,N_19958,N_19903);
nand UO_1560 (O_1560,N_19930,N_19875);
or UO_1561 (O_1561,N_19854,N_19851);
xnor UO_1562 (O_1562,N_19881,N_19927);
nand UO_1563 (O_1563,N_19949,N_19954);
nor UO_1564 (O_1564,N_19872,N_19876);
nand UO_1565 (O_1565,N_19842,N_19932);
and UO_1566 (O_1566,N_19845,N_19879);
nor UO_1567 (O_1567,N_19915,N_19897);
nor UO_1568 (O_1568,N_19957,N_19896);
and UO_1569 (O_1569,N_19843,N_19916);
nor UO_1570 (O_1570,N_19887,N_19939);
and UO_1571 (O_1571,N_19870,N_19934);
nor UO_1572 (O_1572,N_19903,N_19927);
and UO_1573 (O_1573,N_19957,N_19994);
nor UO_1574 (O_1574,N_19989,N_19948);
or UO_1575 (O_1575,N_19843,N_19947);
or UO_1576 (O_1576,N_19962,N_19908);
or UO_1577 (O_1577,N_19888,N_19855);
xnor UO_1578 (O_1578,N_19882,N_19862);
nor UO_1579 (O_1579,N_19925,N_19942);
or UO_1580 (O_1580,N_19979,N_19966);
and UO_1581 (O_1581,N_19860,N_19864);
or UO_1582 (O_1582,N_19844,N_19961);
nor UO_1583 (O_1583,N_19964,N_19997);
nor UO_1584 (O_1584,N_19877,N_19886);
nand UO_1585 (O_1585,N_19992,N_19871);
nand UO_1586 (O_1586,N_19996,N_19877);
nor UO_1587 (O_1587,N_19918,N_19859);
and UO_1588 (O_1588,N_19903,N_19980);
nor UO_1589 (O_1589,N_19996,N_19976);
or UO_1590 (O_1590,N_19990,N_19944);
xor UO_1591 (O_1591,N_19912,N_19886);
or UO_1592 (O_1592,N_19870,N_19915);
and UO_1593 (O_1593,N_19851,N_19879);
nand UO_1594 (O_1594,N_19849,N_19938);
and UO_1595 (O_1595,N_19884,N_19840);
and UO_1596 (O_1596,N_19889,N_19996);
nor UO_1597 (O_1597,N_19861,N_19871);
nor UO_1598 (O_1598,N_19975,N_19904);
xnor UO_1599 (O_1599,N_19881,N_19841);
xnor UO_1600 (O_1600,N_19924,N_19992);
xnor UO_1601 (O_1601,N_19977,N_19847);
and UO_1602 (O_1602,N_19843,N_19859);
nand UO_1603 (O_1603,N_19884,N_19925);
nor UO_1604 (O_1604,N_19906,N_19953);
xnor UO_1605 (O_1605,N_19873,N_19851);
or UO_1606 (O_1606,N_19905,N_19851);
or UO_1607 (O_1607,N_19975,N_19968);
or UO_1608 (O_1608,N_19973,N_19841);
or UO_1609 (O_1609,N_19945,N_19902);
nand UO_1610 (O_1610,N_19988,N_19938);
nand UO_1611 (O_1611,N_19969,N_19865);
or UO_1612 (O_1612,N_19937,N_19965);
nor UO_1613 (O_1613,N_19867,N_19947);
nor UO_1614 (O_1614,N_19840,N_19957);
nand UO_1615 (O_1615,N_19929,N_19915);
and UO_1616 (O_1616,N_19933,N_19855);
or UO_1617 (O_1617,N_19940,N_19914);
and UO_1618 (O_1618,N_19846,N_19854);
and UO_1619 (O_1619,N_19890,N_19884);
nor UO_1620 (O_1620,N_19918,N_19964);
and UO_1621 (O_1621,N_19861,N_19972);
or UO_1622 (O_1622,N_19912,N_19892);
nand UO_1623 (O_1623,N_19906,N_19925);
and UO_1624 (O_1624,N_19961,N_19996);
and UO_1625 (O_1625,N_19875,N_19870);
xnor UO_1626 (O_1626,N_19879,N_19887);
nor UO_1627 (O_1627,N_19998,N_19852);
xor UO_1628 (O_1628,N_19971,N_19881);
nand UO_1629 (O_1629,N_19974,N_19967);
xnor UO_1630 (O_1630,N_19850,N_19906);
or UO_1631 (O_1631,N_19908,N_19910);
or UO_1632 (O_1632,N_19874,N_19889);
nor UO_1633 (O_1633,N_19954,N_19971);
or UO_1634 (O_1634,N_19918,N_19973);
and UO_1635 (O_1635,N_19905,N_19890);
xor UO_1636 (O_1636,N_19975,N_19944);
xor UO_1637 (O_1637,N_19842,N_19904);
nand UO_1638 (O_1638,N_19991,N_19911);
nor UO_1639 (O_1639,N_19923,N_19908);
nand UO_1640 (O_1640,N_19854,N_19955);
xor UO_1641 (O_1641,N_19898,N_19864);
xor UO_1642 (O_1642,N_19987,N_19933);
nand UO_1643 (O_1643,N_19957,N_19851);
or UO_1644 (O_1644,N_19991,N_19926);
nand UO_1645 (O_1645,N_19918,N_19940);
and UO_1646 (O_1646,N_19950,N_19942);
xor UO_1647 (O_1647,N_19941,N_19943);
nand UO_1648 (O_1648,N_19948,N_19962);
nor UO_1649 (O_1649,N_19997,N_19854);
xnor UO_1650 (O_1650,N_19868,N_19989);
nand UO_1651 (O_1651,N_19895,N_19851);
nand UO_1652 (O_1652,N_19936,N_19905);
and UO_1653 (O_1653,N_19845,N_19974);
xor UO_1654 (O_1654,N_19883,N_19986);
xor UO_1655 (O_1655,N_19851,N_19974);
nand UO_1656 (O_1656,N_19978,N_19930);
xor UO_1657 (O_1657,N_19902,N_19870);
or UO_1658 (O_1658,N_19983,N_19911);
or UO_1659 (O_1659,N_19972,N_19961);
nor UO_1660 (O_1660,N_19999,N_19911);
nand UO_1661 (O_1661,N_19956,N_19945);
and UO_1662 (O_1662,N_19995,N_19982);
or UO_1663 (O_1663,N_19875,N_19878);
nor UO_1664 (O_1664,N_19858,N_19898);
nand UO_1665 (O_1665,N_19984,N_19897);
nor UO_1666 (O_1666,N_19951,N_19876);
xor UO_1667 (O_1667,N_19952,N_19997);
or UO_1668 (O_1668,N_19875,N_19864);
and UO_1669 (O_1669,N_19929,N_19969);
and UO_1670 (O_1670,N_19882,N_19950);
nor UO_1671 (O_1671,N_19987,N_19956);
and UO_1672 (O_1672,N_19967,N_19893);
or UO_1673 (O_1673,N_19954,N_19897);
xor UO_1674 (O_1674,N_19938,N_19903);
nand UO_1675 (O_1675,N_19993,N_19871);
nand UO_1676 (O_1676,N_19960,N_19918);
nand UO_1677 (O_1677,N_19939,N_19938);
nor UO_1678 (O_1678,N_19917,N_19846);
xor UO_1679 (O_1679,N_19967,N_19879);
or UO_1680 (O_1680,N_19940,N_19854);
nand UO_1681 (O_1681,N_19930,N_19991);
or UO_1682 (O_1682,N_19850,N_19934);
nor UO_1683 (O_1683,N_19894,N_19917);
xor UO_1684 (O_1684,N_19916,N_19933);
or UO_1685 (O_1685,N_19903,N_19868);
nand UO_1686 (O_1686,N_19978,N_19923);
nand UO_1687 (O_1687,N_19876,N_19920);
nor UO_1688 (O_1688,N_19917,N_19964);
and UO_1689 (O_1689,N_19998,N_19903);
or UO_1690 (O_1690,N_19986,N_19962);
and UO_1691 (O_1691,N_19842,N_19843);
nor UO_1692 (O_1692,N_19880,N_19965);
xnor UO_1693 (O_1693,N_19952,N_19850);
nor UO_1694 (O_1694,N_19898,N_19987);
and UO_1695 (O_1695,N_19958,N_19982);
and UO_1696 (O_1696,N_19903,N_19877);
nor UO_1697 (O_1697,N_19981,N_19914);
and UO_1698 (O_1698,N_19908,N_19930);
nor UO_1699 (O_1699,N_19892,N_19855);
xnor UO_1700 (O_1700,N_19875,N_19949);
and UO_1701 (O_1701,N_19868,N_19943);
or UO_1702 (O_1702,N_19978,N_19846);
nand UO_1703 (O_1703,N_19951,N_19857);
or UO_1704 (O_1704,N_19960,N_19848);
nor UO_1705 (O_1705,N_19992,N_19971);
nand UO_1706 (O_1706,N_19970,N_19914);
or UO_1707 (O_1707,N_19869,N_19899);
nand UO_1708 (O_1708,N_19984,N_19952);
nand UO_1709 (O_1709,N_19853,N_19927);
nand UO_1710 (O_1710,N_19872,N_19861);
or UO_1711 (O_1711,N_19979,N_19861);
nor UO_1712 (O_1712,N_19931,N_19928);
and UO_1713 (O_1713,N_19844,N_19856);
or UO_1714 (O_1714,N_19844,N_19912);
nand UO_1715 (O_1715,N_19846,N_19868);
and UO_1716 (O_1716,N_19976,N_19876);
nor UO_1717 (O_1717,N_19971,N_19850);
nand UO_1718 (O_1718,N_19929,N_19922);
nand UO_1719 (O_1719,N_19883,N_19974);
or UO_1720 (O_1720,N_19840,N_19873);
and UO_1721 (O_1721,N_19911,N_19887);
xnor UO_1722 (O_1722,N_19946,N_19997);
and UO_1723 (O_1723,N_19910,N_19843);
or UO_1724 (O_1724,N_19988,N_19885);
xnor UO_1725 (O_1725,N_19847,N_19864);
xnor UO_1726 (O_1726,N_19873,N_19876);
nor UO_1727 (O_1727,N_19911,N_19896);
or UO_1728 (O_1728,N_19842,N_19853);
xnor UO_1729 (O_1729,N_19999,N_19994);
or UO_1730 (O_1730,N_19863,N_19985);
nand UO_1731 (O_1731,N_19997,N_19907);
nor UO_1732 (O_1732,N_19928,N_19853);
xor UO_1733 (O_1733,N_19883,N_19898);
and UO_1734 (O_1734,N_19846,N_19937);
xor UO_1735 (O_1735,N_19931,N_19910);
nor UO_1736 (O_1736,N_19907,N_19841);
nor UO_1737 (O_1737,N_19946,N_19958);
or UO_1738 (O_1738,N_19927,N_19948);
xor UO_1739 (O_1739,N_19913,N_19971);
nand UO_1740 (O_1740,N_19893,N_19964);
nor UO_1741 (O_1741,N_19966,N_19925);
or UO_1742 (O_1742,N_19878,N_19949);
nand UO_1743 (O_1743,N_19899,N_19962);
and UO_1744 (O_1744,N_19931,N_19904);
nor UO_1745 (O_1745,N_19877,N_19975);
and UO_1746 (O_1746,N_19891,N_19881);
nand UO_1747 (O_1747,N_19849,N_19985);
or UO_1748 (O_1748,N_19906,N_19890);
or UO_1749 (O_1749,N_19956,N_19996);
nand UO_1750 (O_1750,N_19953,N_19931);
and UO_1751 (O_1751,N_19910,N_19967);
or UO_1752 (O_1752,N_19986,N_19963);
nor UO_1753 (O_1753,N_19926,N_19946);
xnor UO_1754 (O_1754,N_19915,N_19874);
xor UO_1755 (O_1755,N_19905,N_19953);
or UO_1756 (O_1756,N_19855,N_19958);
xnor UO_1757 (O_1757,N_19852,N_19856);
nor UO_1758 (O_1758,N_19971,N_19846);
or UO_1759 (O_1759,N_19911,N_19926);
or UO_1760 (O_1760,N_19920,N_19982);
nand UO_1761 (O_1761,N_19976,N_19904);
nand UO_1762 (O_1762,N_19943,N_19863);
nor UO_1763 (O_1763,N_19944,N_19909);
or UO_1764 (O_1764,N_19999,N_19968);
nor UO_1765 (O_1765,N_19843,N_19874);
nor UO_1766 (O_1766,N_19953,N_19879);
xnor UO_1767 (O_1767,N_19848,N_19988);
nor UO_1768 (O_1768,N_19975,N_19930);
or UO_1769 (O_1769,N_19988,N_19983);
and UO_1770 (O_1770,N_19966,N_19879);
nor UO_1771 (O_1771,N_19906,N_19872);
nand UO_1772 (O_1772,N_19893,N_19982);
or UO_1773 (O_1773,N_19997,N_19933);
or UO_1774 (O_1774,N_19907,N_19852);
or UO_1775 (O_1775,N_19932,N_19968);
nor UO_1776 (O_1776,N_19974,N_19915);
xor UO_1777 (O_1777,N_19955,N_19891);
nand UO_1778 (O_1778,N_19873,N_19895);
nor UO_1779 (O_1779,N_19900,N_19949);
nor UO_1780 (O_1780,N_19943,N_19900);
or UO_1781 (O_1781,N_19855,N_19920);
or UO_1782 (O_1782,N_19946,N_19952);
nand UO_1783 (O_1783,N_19876,N_19917);
xnor UO_1784 (O_1784,N_19860,N_19987);
or UO_1785 (O_1785,N_19895,N_19933);
xnor UO_1786 (O_1786,N_19928,N_19906);
nand UO_1787 (O_1787,N_19920,N_19893);
and UO_1788 (O_1788,N_19995,N_19943);
and UO_1789 (O_1789,N_19961,N_19850);
nor UO_1790 (O_1790,N_19886,N_19902);
and UO_1791 (O_1791,N_19855,N_19864);
nand UO_1792 (O_1792,N_19890,N_19940);
xnor UO_1793 (O_1793,N_19879,N_19957);
nand UO_1794 (O_1794,N_19876,N_19960);
or UO_1795 (O_1795,N_19843,N_19918);
nand UO_1796 (O_1796,N_19860,N_19953);
and UO_1797 (O_1797,N_19961,N_19856);
xnor UO_1798 (O_1798,N_19856,N_19878);
xnor UO_1799 (O_1799,N_19919,N_19869);
xor UO_1800 (O_1800,N_19986,N_19995);
xnor UO_1801 (O_1801,N_19904,N_19883);
nand UO_1802 (O_1802,N_19909,N_19990);
xnor UO_1803 (O_1803,N_19882,N_19928);
and UO_1804 (O_1804,N_19882,N_19844);
nor UO_1805 (O_1805,N_19986,N_19863);
nand UO_1806 (O_1806,N_19845,N_19881);
xnor UO_1807 (O_1807,N_19913,N_19944);
nand UO_1808 (O_1808,N_19980,N_19902);
nor UO_1809 (O_1809,N_19840,N_19923);
nand UO_1810 (O_1810,N_19977,N_19933);
and UO_1811 (O_1811,N_19844,N_19980);
nor UO_1812 (O_1812,N_19980,N_19886);
and UO_1813 (O_1813,N_19844,N_19864);
nor UO_1814 (O_1814,N_19932,N_19973);
xnor UO_1815 (O_1815,N_19886,N_19903);
nand UO_1816 (O_1816,N_19983,N_19919);
nor UO_1817 (O_1817,N_19957,N_19870);
nand UO_1818 (O_1818,N_19931,N_19883);
and UO_1819 (O_1819,N_19908,N_19914);
xor UO_1820 (O_1820,N_19940,N_19973);
or UO_1821 (O_1821,N_19921,N_19919);
and UO_1822 (O_1822,N_19919,N_19904);
nand UO_1823 (O_1823,N_19955,N_19859);
and UO_1824 (O_1824,N_19849,N_19971);
nand UO_1825 (O_1825,N_19975,N_19857);
or UO_1826 (O_1826,N_19875,N_19924);
nand UO_1827 (O_1827,N_19893,N_19949);
nor UO_1828 (O_1828,N_19940,N_19902);
or UO_1829 (O_1829,N_19956,N_19927);
and UO_1830 (O_1830,N_19978,N_19847);
nor UO_1831 (O_1831,N_19873,N_19977);
and UO_1832 (O_1832,N_19963,N_19983);
nor UO_1833 (O_1833,N_19985,N_19852);
nor UO_1834 (O_1834,N_19998,N_19868);
or UO_1835 (O_1835,N_19956,N_19957);
and UO_1836 (O_1836,N_19860,N_19911);
and UO_1837 (O_1837,N_19850,N_19980);
or UO_1838 (O_1838,N_19944,N_19895);
nor UO_1839 (O_1839,N_19862,N_19983);
nand UO_1840 (O_1840,N_19928,N_19988);
nand UO_1841 (O_1841,N_19867,N_19937);
nor UO_1842 (O_1842,N_19955,N_19861);
nor UO_1843 (O_1843,N_19861,N_19969);
nor UO_1844 (O_1844,N_19887,N_19884);
nor UO_1845 (O_1845,N_19841,N_19899);
nor UO_1846 (O_1846,N_19944,N_19875);
or UO_1847 (O_1847,N_19847,N_19960);
or UO_1848 (O_1848,N_19843,N_19933);
or UO_1849 (O_1849,N_19964,N_19965);
nand UO_1850 (O_1850,N_19963,N_19840);
xor UO_1851 (O_1851,N_19981,N_19881);
and UO_1852 (O_1852,N_19965,N_19974);
and UO_1853 (O_1853,N_19995,N_19916);
nor UO_1854 (O_1854,N_19888,N_19848);
or UO_1855 (O_1855,N_19867,N_19885);
xor UO_1856 (O_1856,N_19919,N_19945);
and UO_1857 (O_1857,N_19991,N_19849);
xnor UO_1858 (O_1858,N_19871,N_19956);
or UO_1859 (O_1859,N_19950,N_19951);
xor UO_1860 (O_1860,N_19947,N_19885);
nor UO_1861 (O_1861,N_19988,N_19950);
nor UO_1862 (O_1862,N_19866,N_19926);
or UO_1863 (O_1863,N_19971,N_19870);
nor UO_1864 (O_1864,N_19894,N_19897);
nand UO_1865 (O_1865,N_19964,N_19953);
xor UO_1866 (O_1866,N_19956,N_19842);
nand UO_1867 (O_1867,N_19975,N_19953);
nand UO_1868 (O_1868,N_19988,N_19901);
nand UO_1869 (O_1869,N_19991,N_19900);
nand UO_1870 (O_1870,N_19848,N_19953);
xor UO_1871 (O_1871,N_19890,N_19990);
xnor UO_1872 (O_1872,N_19951,N_19907);
or UO_1873 (O_1873,N_19941,N_19987);
nand UO_1874 (O_1874,N_19901,N_19936);
nand UO_1875 (O_1875,N_19880,N_19961);
xor UO_1876 (O_1876,N_19849,N_19852);
xnor UO_1877 (O_1877,N_19904,N_19994);
nand UO_1878 (O_1878,N_19888,N_19990);
or UO_1879 (O_1879,N_19842,N_19887);
xor UO_1880 (O_1880,N_19847,N_19987);
xnor UO_1881 (O_1881,N_19952,N_19964);
and UO_1882 (O_1882,N_19884,N_19970);
or UO_1883 (O_1883,N_19870,N_19843);
nand UO_1884 (O_1884,N_19976,N_19949);
or UO_1885 (O_1885,N_19842,N_19959);
and UO_1886 (O_1886,N_19884,N_19854);
nor UO_1887 (O_1887,N_19945,N_19887);
nor UO_1888 (O_1888,N_19982,N_19939);
xnor UO_1889 (O_1889,N_19977,N_19874);
xor UO_1890 (O_1890,N_19987,N_19854);
nor UO_1891 (O_1891,N_19876,N_19844);
nor UO_1892 (O_1892,N_19876,N_19879);
or UO_1893 (O_1893,N_19862,N_19943);
xnor UO_1894 (O_1894,N_19911,N_19872);
and UO_1895 (O_1895,N_19892,N_19941);
or UO_1896 (O_1896,N_19891,N_19879);
nor UO_1897 (O_1897,N_19902,N_19974);
xnor UO_1898 (O_1898,N_19940,N_19841);
nand UO_1899 (O_1899,N_19927,N_19945);
nor UO_1900 (O_1900,N_19903,N_19965);
nand UO_1901 (O_1901,N_19861,N_19953);
xnor UO_1902 (O_1902,N_19999,N_19870);
xnor UO_1903 (O_1903,N_19909,N_19875);
xor UO_1904 (O_1904,N_19849,N_19942);
nor UO_1905 (O_1905,N_19915,N_19923);
xnor UO_1906 (O_1906,N_19980,N_19932);
and UO_1907 (O_1907,N_19852,N_19955);
nor UO_1908 (O_1908,N_19976,N_19994);
xnor UO_1909 (O_1909,N_19961,N_19997);
and UO_1910 (O_1910,N_19891,N_19848);
nor UO_1911 (O_1911,N_19870,N_19872);
nand UO_1912 (O_1912,N_19924,N_19909);
nor UO_1913 (O_1913,N_19926,N_19970);
and UO_1914 (O_1914,N_19905,N_19961);
nor UO_1915 (O_1915,N_19888,N_19924);
nor UO_1916 (O_1916,N_19863,N_19923);
nand UO_1917 (O_1917,N_19979,N_19940);
nor UO_1918 (O_1918,N_19960,N_19906);
or UO_1919 (O_1919,N_19897,N_19860);
or UO_1920 (O_1920,N_19928,N_19990);
nand UO_1921 (O_1921,N_19851,N_19956);
and UO_1922 (O_1922,N_19915,N_19963);
and UO_1923 (O_1923,N_19931,N_19956);
xor UO_1924 (O_1924,N_19887,N_19941);
or UO_1925 (O_1925,N_19897,N_19871);
xnor UO_1926 (O_1926,N_19850,N_19872);
nor UO_1927 (O_1927,N_19992,N_19958);
nor UO_1928 (O_1928,N_19948,N_19964);
or UO_1929 (O_1929,N_19965,N_19958);
or UO_1930 (O_1930,N_19858,N_19883);
nor UO_1931 (O_1931,N_19956,N_19846);
or UO_1932 (O_1932,N_19913,N_19919);
xnor UO_1933 (O_1933,N_19878,N_19974);
or UO_1934 (O_1934,N_19991,N_19972);
or UO_1935 (O_1935,N_19921,N_19860);
nand UO_1936 (O_1936,N_19890,N_19926);
nor UO_1937 (O_1937,N_19867,N_19999);
nand UO_1938 (O_1938,N_19991,N_19840);
xnor UO_1939 (O_1939,N_19954,N_19953);
or UO_1940 (O_1940,N_19860,N_19875);
and UO_1941 (O_1941,N_19992,N_19931);
nand UO_1942 (O_1942,N_19998,N_19866);
nand UO_1943 (O_1943,N_19963,N_19967);
xnor UO_1944 (O_1944,N_19882,N_19895);
and UO_1945 (O_1945,N_19952,N_19981);
and UO_1946 (O_1946,N_19935,N_19969);
and UO_1947 (O_1947,N_19894,N_19863);
or UO_1948 (O_1948,N_19927,N_19904);
xor UO_1949 (O_1949,N_19903,N_19866);
and UO_1950 (O_1950,N_19993,N_19947);
xnor UO_1951 (O_1951,N_19915,N_19964);
nand UO_1952 (O_1952,N_19990,N_19856);
xor UO_1953 (O_1953,N_19905,N_19939);
nand UO_1954 (O_1954,N_19878,N_19976);
xnor UO_1955 (O_1955,N_19926,N_19938);
xnor UO_1956 (O_1956,N_19977,N_19967);
or UO_1957 (O_1957,N_19948,N_19942);
nor UO_1958 (O_1958,N_19964,N_19848);
nand UO_1959 (O_1959,N_19867,N_19988);
nor UO_1960 (O_1960,N_19960,N_19948);
or UO_1961 (O_1961,N_19932,N_19896);
nor UO_1962 (O_1962,N_19974,N_19969);
and UO_1963 (O_1963,N_19870,N_19885);
nor UO_1964 (O_1964,N_19979,N_19978);
nand UO_1965 (O_1965,N_19947,N_19963);
xor UO_1966 (O_1966,N_19982,N_19845);
xnor UO_1967 (O_1967,N_19952,N_19893);
nand UO_1968 (O_1968,N_19840,N_19987);
xnor UO_1969 (O_1969,N_19959,N_19990);
and UO_1970 (O_1970,N_19888,N_19994);
or UO_1971 (O_1971,N_19943,N_19843);
nor UO_1972 (O_1972,N_19979,N_19933);
nor UO_1973 (O_1973,N_19932,N_19859);
and UO_1974 (O_1974,N_19860,N_19998);
and UO_1975 (O_1975,N_19935,N_19957);
nand UO_1976 (O_1976,N_19964,N_19995);
or UO_1977 (O_1977,N_19953,N_19844);
and UO_1978 (O_1978,N_19918,N_19878);
and UO_1979 (O_1979,N_19908,N_19947);
nor UO_1980 (O_1980,N_19869,N_19846);
nor UO_1981 (O_1981,N_19876,N_19945);
or UO_1982 (O_1982,N_19887,N_19929);
or UO_1983 (O_1983,N_19860,N_19891);
nor UO_1984 (O_1984,N_19899,N_19848);
xor UO_1985 (O_1985,N_19893,N_19846);
or UO_1986 (O_1986,N_19850,N_19990);
nand UO_1987 (O_1987,N_19920,N_19886);
nor UO_1988 (O_1988,N_19871,N_19903);
nand UO_1989 (O_1989,N_19896,N_19887);
or UO_1990 (O_1990,N_19844,N_19919);
and UO_1991 (O_1991,N_19845,N_19927);
nor UO_1992 (O_1992,N_19996,N_19993);
or UO_1993 (O_1993,N_19980,N_19991);
nand UO_1994 (O_1994,N_19866,N_19976);
nor UO_1995 (O_1995,N_19996,N_19992);
nand UO_1996 (O_1996,N_19962,N_19868);
nor UO_1997 (O_1997,N_19973,N_19958);
nand UO_1998 (O_1998,N_19864,N_19969);
nand UO_1999 (O_1999,N_19924,N_19851);
and UO_2000 (O_2000,N_19917,N_19956);
and UO_2001 (O_2001,N_19912,N_19846);
xnor UO_2002 (O_2002,N_19931,N_19964);
nand UO_2003 (O_2003,N_19899,N_19895);
xnor UO_2004 (O_2004,N_19983,N_19952);
nor UO_2005 (O_2005,N_19867,N_19976);
or UO_2006 (O_2006,N_19979,N_19994);
nor UO_2007 (O_2007,N_19896,N_19877);
and UO_2008 (O_2008,N_19866,N_19931);
xor UO_2009 (O_2009,N_19941,N_19846);
nor UO_2010 (O_2010,N_19848,N_19992);
nand UO_2011 (O_2011,N_19852,N_19914);
and UO_2012 (O_2012,N_19863,N_19898);
nor UO_2013 (O_2013,N_19981,N_19875);
and UO_2014 (O_2014,N_19853,N_19885);
nor UO_2015 (O_2015,N_19971,N_19878);
xor UO_2016 (O_2016,N_19995,N_19912);
nand UO_2017 (O_2017,N_19922,N_19910);
or UO_2018 (O_2018,N_19970,N_19932);
or UO_2019 (O_2019,N_19931,N_19920);
or UO_2020 (O_2020,N_19875,N_19904);
or UO_2021 (O_2021,N_19885,N_19963);
and UO_2022 (O_2022,N_19987,N_19978);
xor UO_2023 (O_2023,N_19965,N_19873);
nor UO_2024 (O_2024,N_19893,N_19984);
or UO_2025 (O_2025,N_19841,N_19860);
and UO_2026 (O_2026,N_19946,N_19878);
or UO_2027 (O_2027,N_19896,N_19929);
and UO_2028 (O_2028,N_19865,N_19976);
or UO_2029 (O_2029,N_19854,N_19973);
nor UO_2030 (O_2030,N_19866,N_19956);
nand UO_2031 (O_2031,N_19927,N_19855);
nor UO_2032 (O_2032,N_19845,N_19992);
nor UO_2033 (O_2033,N_19958,N_19969);
and UO_2034 (O_2034,N_19924,N_19966);
and UO_2035 (O_2035,N_19996,N_19950);
or UO_2036 (O_2036,N_19903,N_19934);
and UO_2037 (O_2037,N_19848,N_19871);
or UO_2038 (O_2038,N_19841,N_19866);
xnor UO_2039 (O_2039,N_19880,N_19883);
xnor UO_2040 (O_2040,N_19918,N_19920);
and UO_2041 (O_2041,N_19963,N_19876);
or UO_2042 (O_2042,N_19911,N_19916);
or UO_2043 (O_2043,N_19995,N_19863);
and UO_2044 (O_2044,N_19981,N_19870);
and UO_2045 (O_2045,N_19869,N_19864);
xnor UO_2046 (O_2046,N_19989,N_19923);
or UO_2047 (O_2047,N_19865,N_19929);
nand UO_2048 (O_2048,N_19900,N_19962);
nand UO_2049 (O_2049,N_19893,N_19864);
nand UO_2050 (O_2050,N_19950,N_19893);
nor UO_2051 (O_2051,N_19990,N_19974);
or UO_2052 (O_2052,N_19881,N_19993);
or UO_2053 (O_2053,N_19889,N_19868);
nor UO_2054 (O_2054,N_19866,N_19901);
and UO_2055 (O_2055,N_19953,N_19980);
and UO_2056 (O_2056,N_19994,N_19860);
xnor UO_2057 (O_2057,N_19983,N_19950);
or UO_2058 (O_2058,N_19917,N_19887);
nand UO_2059 (O_2059,N_19861,N_19946);
xnor UO_2060 (O_2060,N_19931,N_19984);
nand UO_2061 (O_2061,N_19931,N_19981);
nor UO_2062 (O_2062,N_19960,N_19853);
nor UO_2063 (O_2063,N_19972,N_19949);
xnor UO_2064 (O_2064,N_19855,N_19951);
or UO_2065 (O_2065,N_19941,N_19938);
nor UO_2066 (O_2066,N_19866,N_19966);
nand UO_2067 (O_2067,N_19842,N_19983);
and UO_2068 (O_2068,N_19867,N_19922);
xor UO_2069 (O_2069,N_19877,N_19931);
or UO_2070 (O_2070,N_19999,N_19906);
nand UO_2071 (O_2071,N_19897,N_19868);
xnor UO_2072 (O_2072,N_19937,N_19929);
nor UO_2073 (O_2073,N_19845,N_19975);
nand UO_2074 (O_2074,N_19984,N_19963);
xor UO_2075 (O_2075,N_19997,N_19900);
xnor UO_2076 (O_2076,N_19913,N_19896);
and UO_2077 (O_2077,N_19984,N_19915);
nand UO_2078 (O_2078,N_19974,N_19946);
xnor UO_2079 (O_2079,N_19920,N_19933);
and UO_2080 (O_2080,N_19909,N_19949);
xor UO_2081 (O_2081,N_19922,N_19982);
nand UO_2082 (O_2082,N_19942,N_19914);
and UO_2083 (O_2083,N_19915,N_19925);
or UO_2084 (O_2084,N_19848,N_19989);
or UO_2085 (O_2085,N_19841,N_19992);
or UO_2086 (O_2086,N_19882,N_19971);
or UO_2087 (O_2087,N_19892,N_19894);
nor UO_2088 (O_2088,N_19868,N_19862);
nand UO_2089 (O_2089,N_19955,N_19869);
xor UO_2090 (O_2090,N_19873,N_19921);
and UO_2091 (O_2091,N_19905,N_19995);
and UO_2092 (O_2092,N_19907,N_19932);
or UO_2093 (O_2093,N_19994,N_19885);
xor UO_2094 (O_2094,N_19863,N_19896);
nor UO_2095 (O_2095,N_19884,N_19997);
nand UO_2096 (O_2096,N_19942,N_19932);
or UO_2097 (O_2097,N_19901,N_19998);
nor UO_2098 (O_2098,N_19981,N_19934);
or UO_2099 (O_2099,N_19995,N_19923);
xor UO_2100 (O_2100,N_19921,N_19966);
nand UO_2101 (O_2101,N_19925,N_19950);
or UO_2102 (O_2102,N_19917,N_19905);
xor UO_2103 (O_2103,N_19886,N_19885);
nand UO_2104 (O_2104,N_19965,N_19972);
xnor UO_2105 (O_2105,N_19955,N_19866);
and UO_2106 (O_2106,N_19977,N_19991);
xor UO_2107 (O_2107,N_19890,N_19955);
xor UO_2108 (O_2108,N_19913,N_19924);
or UO_2109 (O_2109,N_19889,N_19903);
nand UO_2110 (O_2110,N_19915,N_19850);
and UO_2111 (O_2111,N_19896,N_19906);
and UO_2112 (O_2112,N_19979,N_19893);
or UO_2113 (O_2113,N_19974,N_19879);
nand UO_2114 (O_2114,N_19959,N_19986);
xor UO_2115 (O_2115,N_19885,N_19917);
xor UO_2116 (O_2116,N_19995,N_19930);
or UO_2117 (O_2117,N_19967,N_19926);
xnor UO_2118 (O_2118,N_19867,N_19936);
and UO_2119 (O_2119,N_19928,N_19981);
or UO_2120 (O_2120,N_19928,N_19941);
and UO_2121 (O_2121,N_19862,N_19939);
nor UO_2122 (O_2122,N_19902,N_19963);
xor UO_2123 (O_2123,N_19845,N_19866);
nand UO_2124 (O_2124,N_19973,N_19992);
nor UO_2125 (O_2125,N_19858,N_19859);
and UO_2126 (O_2126,N_19840,N_19908);
nand UO_2127 (O_2127,N_19901,N_19977);
and UO_2128 (O_2128,N_19901,N_19882);
xor UO_2129 (O_2129,N_19842,N_19851);
or UO_2130 (O_2130,N_19950,N_19880);
nor UO_2131 (O_2131,N_19977,N_19853);
and UO_2132 (O_2132,N_19988,N_19862);
and UO_2133 (O_2133,N_19955,N_19894);
or UO_2134 (O_2134,N_19907,N_19850);
or UO_2135 (O_2135,N_19861,N_19922);
and UO_2136 (O_2136,N_19885,N_19992);
nor UO_2137 (O_2137,N_19955,N_19947);
nor UO_2138 (O_2138,N_19910,N_19840);
or UO_2139 (O_2139,N_19916,N_19931);
nor UO_2140 (O_2140,N_19852,N_19950);
or UO_2141 (O_2141,N_19935,N_19991);
xor UO_2142 (O_2142,N_19850,N_19858);
xor UO_2143 (O_2143,N_19991,N_19985);
nand UO_2144 (O_2144,N_19929,N_19983);
and UO_2145 (O_2145,N_19972,N_19967);
and UO_2146 (O_2146,N_19891,N_19925);
xnor UO_2147 (O_2147,N_19989,N_19862);
nor UO_2148 (O_2148,N_19998,N_19928);
xnor UO_2149 (O_2149,N_19879,N_19866);
and UO_2150 (O_2150,N_19897,N_19980);
nor UO_2151 (O_2151,N_19907,N_19842);
or UO_2152 (O_2152,N_19915,N_19953);
nand UO_2153 (O_2153,N_19861,N_19898);
xnor UO_2154 (O_2154,N_19870,N_19951);
xnor UO_2155 (O_2155,N_19840,N_19952);
nand UO_2156 (O_2156,N_19849,N_19908);
and UO_2157 (O_2157,N_19995,N_19898);
xnor UO_2158 (O_2158,N_19978,N_19840);
nor UO_2159 (O_2159,N_19974,N_19904);
xor UO_2160 (O_2160,N_19940,N_19881);
and UO_2161 (O_2161,N_19890,N_19989);
nand UO_2162 (O_2162,N_19895,N_19881);
nor UO_2163 (O_2163,N_19890,N_19924);
nand UO_2164 (O_2164,N_19956,N_19916);
nand UO_2165 (O_2165,N_19930,N_19911);
or UO_2166 (O_2166,N_19942,N_19979);
xor UO_2167 (O_2167,N_19893,N_19992);
xnor UO_2168 (O_2168,N_19857,N_19963);
and UO_2169 (O_2169,N_19897,N_19863);
nand UO_2170 (O_2170,N_19899,N_19894);
nor UO_2171 (O_2171,N_19843,N_19946);
xnor UO_2172 (O_2172,N_19870,N_19973);
and UO_2173 (O_2173,N_19958,N_19888);
nand UO_2174 (O_2174,N_19930,N_19971);
or UO_2175 (O_2175,N_19937,N_19999);
nor UO_2176 (O_2176,N_19844,N_19958);
xnor UO_2177 (O_2177,N_19914,N_19933);
xor UO_2178 (O_2178,N_19846,N_19910);
and UO_2179 (O_2179,N_19849,N_19890);
xor UO_2180 (O_2180,N_19866,N_19935);
nand UO_2181 (O_2181,N_19842,N_19900);
or UO_2182 (O_2182,N_19928,N_19930);
nor UO_2183 (O_2183,N_19966,N_19973);
nand UO_2184 (O_2184,N_19868,N_19930);
xor UO_2185 (O_2185,N_19952,N_19881);
xnor UO_2186 (O_2186,N_19890,N_19957);
nand UO_2187 (O_2187,N_19863,N_19913);
or UO_2188 (O_2188,N_19926,N_19936);
and UO_2189 (O_2189,N_19979,N_19913);
or UO_2190 (O_2190,N_19893,N_19975);
nand UO_2191 (O_2191,N_19939,N_19900);
nand UO_2192 (O_2192,N_19976,N_19943);
or UO_2193 (O_2193,N_19974,N_19884);
xor UO_2194 (O_2194,N_19882,N_19997);
nand UO_2195 (O_2195,N_19990,N_19915);
nand UO_2196 (O_2196,N_19881,N_19850);
nor UO_2197 (O_2197,N_19929,N_19931);
or UO_2198 (O_2198,N_19845,N_19923);
and UO_2199 (O_2199,N_19969,N_19905);
nand UO_2200 (O_2200,N_19878,N_19945);
xnor UO_2201 (O_2201,N_19974,N_19862);
and UO_2202 (O_2202,N_19935,N_19850);
xor UO_2203 (O_2203,N_19925,N_19982);
and UO_2204 (O_2204,N_19968,N_19940);
and UO_2205 (O_2205,N_19933,N_19944);
or UO_2206 (O_2206,N_19878,N_19915);
or UO_2207 (O_2207,N_19848,N_19903);
and UO_2208 (O_2208,N_19909,N_19903);
nor UO_2209 (O_2209,N_19859,N_19993);
or UO_2210 (O_2210,N_19924,N_19928);
nand UO_2211 (O_2211,N_19986,N_19856);
or UO_2212 (O_2212,N_19997,N_19888);
nor UO_2213 (O_2213,N_19857,N_19978);
nand UO_2214 (O_2214,N_19916,N_19857);
xnor UO_2215 (O_2215,N_19869,N_19929);
nor UO_2216 (O_2216,N_19980,N_19912);
and UO_2217 (O_2217,N_19969,N_19976);
xnor UO_2218 (O_2218,N_19945,N_19939);
nor UO_2219 (O_2219,N_19872,N_19975);
nand UO_2220 (O_2220,N_19907,N_19904);
and UO_2221 (O_2221,N_19994,N_19848);
and UO_2222 (O_2222,N_19960,N_19868);
and UO_2223 (O_2223,N_19852,N_19986);
nor UO_2224 (O_2224,N_19968,N_19888);
nand UO_2225 (O_2225,N_19971,N_19941);
xnor UO_2226 (O_2226,N_19854,N_19881);
and UO_2227 (O_2227,N_19875,N_19908);
xnor UO_2228 (O_2228,N_19868,N_19971);
nor UO_2229 (O_2229,N_19842,N_19866);
nand UO_2230 (O_2230,N_19845,N_19943);
xor UO_2231 (O_2231,N_19943,N_19854);
nor UO_2232 (O_2232,N_19929,N_19913);
or UO_2233 (O_2233,N_19915,N_19985);
xor UO_2234 (O_2234,N_19904,N_19929);
or UO_2235 (O_2235,N_19858,N_19930);
nor UO_2236 (O_2236,N_19933,N_19969);
and UO_2237 (O_2237,N_19954,N_19883);
nor UO_2238 (O_2238,N_19965,N_19910);
xor UO_2239 (O_2239,N_19979,N_19921);
or UO_2240 (O_2240,N_19918,N_19943);
xnor UO_2241 (O_2241,N_19900,N_19992);
nand UO_2242 (O_2242,N_19942,N_19931);
nand UO_2243 (O_2243,N_19847,N_19845);
or UO_2244 (O_2244,N_19912,N_19932);
xnor UO_2245 (O_2245,N_19929,N_19955);
and UO_2246 (O_2246,N_19871,N_19894);
nor UO_2247 (O_2247,N_19891,N_19964);
nor UO_2248 (O_2248,N_19907,N_19871);
nor UO_2249 (O_2249,N_19913,N_19937);
or UO_2250 (O_2250,N_19943,N_19985);
nor UO_2251 (O_2251,N_19928,N_19947);
nor UO_2252 (O_2252,N_19913,N_19925);
nand UO_2253 (O_2253,N_19924,N_19948);
nor UO_2254 (O_2254,N_19865,N_19891);
xnor UO_2255 (O_2255,N_19942,N_19926);
xor UO_2256 (O_2256,N_19939,N_19885);
xor UO_2257 (O_2257,N_19958,N_19910);
or UO_2258 (O_2258,N_19844,N_19996);
nor UO_2259 (O_2259,N_19861,N_19954);
nand UO_2260 (O_2260,N_19981,N_19876);
nor UO_2261 (O_2261,N_19848,N_19863);
or UO_2262 (O_2262,N_19880,N_19907);
and UO_2263 (O_2263,N_19922,N_19944);
and UO_2264 (O_2264,N_19968,N_19921);
and UO_2265 (O_2265,N_19861,N_19998);
and UO_2266 (O_2266,N_19873,N_19882);
or UO_2267 (O_2267,N_19861,N_19942);
and UO_2268 (O_2268,N_19954,N_19898);
xor UO_2269 (O_2269,N_19997,N_19991);
and UO_2270 (O_2270,N_19966,N_19859);
xnor UO_2271 (O_2271,N_19871,N_19914);
nor UO_2272 (O_2272,N_19920,N_19882);
xor UO_2273 (O_2273,N_19979,N_19907);
or UO_2274 (O_2274,N_19883,N_19952);
and UO_2275 (O_2275,N_19981,N_19991);
and UO_2276 (O_2276,N_19912,N_19893);
nor UO_2277 (O_2277,N_19868,N_19946);
nand UO_2278 (O_2278,N_19897,N_19879);
or UO_2279 (O_2279,N_19894,N_19984);
or UO_2280 (O_2280,N_19842,N_19996);
xnor UO_2281 (O_2281,N_19928,N_19912);
nand UO_2282 (O_2282,N_19866,N_19913);
nor UO_2283 (O_2283,N_19874,N_19851);
nor UO_2284 (O_2284,N_19928,N_19873);
xor UO_2285 (O_2285,N_19850,N_19981);
and UO_2286 (O_2286,N_19927,N_19885);
xor UO_2287 (O_2287,N_19996,N_19942);
nand UO_2288 (O_2288,N_19959,N_19932);
nand UO_2289 (O_2289,N_19982,N_19868);
xor UO_2290 (O_2290,N_19906,N_19873);
or UO_2291 (O_2291,N_19852,N_19975);
xnor UO_2292 (O_2292,N_19860,N_19846);
xor UO_2293 (O_2293,N_19985,N_19878);
xor UO_2294 (O_2294,N_19965,N_19842);
nor UO_2295 (O_2295,N_19948,N_19907);
or UO_2296 (O_2296,N_19985,N_19887);
xnor UO_2297 (O_2297,N_19965,N_19966);
and UO_2298 (O_2298,N_19871,N_19961);
and UO_2299 (O_2299,N_19886,N_19874);
nand UO_2300 (O_2300,N_19967,N_19959);
nand UO_2301 (O_2301,N_19887,N_19958);
and UO_2302 (O_2302,N_19850,N_19877);
nand UO_2303 (O_2303,N_19954,N_19995);
and UO_2304 (O_2304,N_19938,N_19885);
or UO_2305 (O_2305,N_19965,N_19895);
nor UO_2306 (O_2306,N_19929,N_19967);
nand UO_2307 (O_2307,N_19886,N_19901);
nand UO_2308 (O_2308,N_19908,N_19944);
nor UO_2309 (O_2309,N_19931,N_19940);
and UO_2310 (O_2310,N_19963,N_19975);
nor UO_2311 (O_2311,N_19840,N_19883);
nand UO_2312 (O_2312,N_19858,N_19958);
and UO_2313 (O_2313,N_19860,N_19973);
xnor UO_2314 (O_2314,N_19947,N_19898);
nor UO_2315 (O_2315,N_19976,N_19860);
nor UO_2316 (O_2316,N_19968,N_19974);
and UO_2317 (O_2317,N_19952,N_19961);
nor UO_2318 (O_2318,N_19849,N_19870);
xor UO_2319 (O_2319,N_19857,N_19954);
nand UO_2320 (O_2320,N_19986,N_19983);
nor UO_2321 (O_2321,N_19998,N_19845);
nor UO_2322 (O_2322,N_19870,N_19969);
nor UO_2323 (O_2323,N_19966,N_19882);
nor UO_2324 (O_2324,N_19906,N_19981);
and UO_2325 (O_2325,N_19932,N_19960);
nand UO_2326 (O_2326,N_19895,N_19847);
or UO_2327 (O_2327,N_19945,N_19855);
and UO_2328 (O_2328,N_19947,N_19968);
nand UO_2329 (O_2329,N_19859,N_19939);
xnor UO_2330 (O_2330,N_19950,N_19845);
or UO_2331 (O_2331,N_19904,N_19935);
nand UO_2332 (O_2332,N_19859,N_19848);
and UO_2333 (O_2333,N_19876,N_19911);
and UO_2334 (O_2334,N_19915,N_19933);
nor UO_2335 (O_2335,N_19888,N_19912);
nand UO_2336 (O_2336,N_19903,N_19966);
and UO_2337 (O_2337,N_19875,N_19852);
or UO_2338 (O_2338,N_19858,N_19878);
nor UO_2339 (O_2339,N_19881,N_19902);
or UO_2340 (O_2340,N_19920,N_19967);
or UO_2341 (O_2341,N_19883,N_19920);
or UO_2342 (O_2342,N_19945,N_19935);
nand UO_2343 (O_2343,N_19893,N_19943);
or UO_2344 (O_2344,N_19947,N_19940);
or UO_2345 (O_2345,N_19910,N_19898);
nand UO_2346 (O_2346,N_19920,N_19884);
nor UO_2347 (O_2347,N_19905,N_19963);
xor UO_2348 (O_2348,N_19871,N_19974);
nand UO_2349 (O_2349,N_19971,N_19867);
nand UO_2350 (O_2350,N_19937,N_19868);
or UO_2351 (O_2351,N_19917,N_19998);
nand UO_2352 (O_2352,N_19973,N_19980);
nand UO_2353 (O_2353,N_19883,N_19976);
and UO_2354 (O_2354,N_19907,N_19911);
nand UO_2355 (O_2355,N_19952,N_19990);
nor UO_2356 (O_2356,N_19888,N_19845);
nor UO_2357 (O_2357,N_19901,N_19994);
nand UO_2358 (O_2358,N_19853,N_19991);
xnor UO_2359 (O_2359,N_19968,N_19934);
xnor UO_2360 (O_2360,N_19918,N_19984);
nand UO_2361 (O_2361,N_19863,N_19954);
or UO_2362 (O_2362,N_19879,N_19914);
and UO_2363 (O_2363,N_19911,N_19974);
nand UO_2364 (O_2364,N_19940,N_19936);
or UO_2365 (O_2365,N_19985,N_19990);
nand UO_2366 (O_2366,N_19885,N_19969);
nor UO_2367 (O_2367,N_19946,N_19980);
or UO_2368 (O_2368,N_19859,N_19919);
and UO_2369 (O_2369,N_19860,N_19931);
or UO_2370 (O_2370,N_19898,N_19999);
nor UO_2371 (O_2371,N_19850,N_19929);
xnor UO_2372 (O_2372,N_19979,N_19905);
nor UO_2373 (O_2373,N_19921,N_19841);
nand UO_2374 (O_2374,N_19897,N_19935);
nand UO_2375 (O_2375,N_19868,N_19949);
nor UO_2376 (O_2376,N_19949,N_19925);
and UO_2377 (O_2377,N_19882,N_19889);
and UO_2378 (O_2378,N_19927,N_19909);
nand UO_2379 (O_2379,N_19949,N_19979);
or UO_2380 (O_2380,N_19995,N_19998);
nor UO_2381 (O_2381,N_19881,N_19959);
nand UO_2382 (O_2382,N_19840,N_19954);
nor UO_2383 (O_2383,N_19965,N_19894);
nor UO_2384 (O_2384,N_19876,N_19888);
and UO_2385 (O_2385,N_19990,N_19854);
and UO_2386 (O_2386,N_19906,N_19931);
and UO_2387 (O_2387,N_19848,N_19877);
and UO_2388 (O_2388,N_19853,N_19919);
nand UO_2389 (O_2389,N_19888,N_19982);
nor UO_2390 (O_2390,N_19968,N_19954);
or UO_2391 (O_2391,N_19982,N_19871);
and UO_2392 (O_2392,N_19927,N_19990);
or UO_2393 (O_2393,N_19850,N_19949);
xor UO_2394 (O_2394,N_19998,N_19967);
nand UO_2395 (O_2395,N_19956,N_19854);
or UO_2396 (O_2396,N_19986,N_19947);
nand UO_2397 (O_2397,N_19873,N_19963);
nand UO_2398 (O_2398,N_19929,N_19986);
or UO_2399 (O_2399,N_19964,N_19927);
or UO_2400 (O_2400,N_19907,N_19988);
nand UO_2401 (O_2401,N_19863,N_19950);
nor UO_2402 (O_2402,N_19914,N_19851);
nor UO_2403 (O_2403,N_19907,N_19952);
xnor UO_2404 (O_2404,N_19897,N_19979);
nor UO_2405 (O_2405,N_19932,N_19952);
nor UO_2406 (O_2406,N_19961,N_19845);
nor UO_2407 (O_2407,N_19944,N_19979);
nor UO_2408 (O_2408,N_19856,N_19913);
nand UO_2409 (O_2409,N_19918,N_19865);
nand UO_2410 (O_2410,N_19934,N_19950);
xor UO_2411 (O_2411,N_19974,N_19889);
nand UO_2412 (O_2412,N_19857,N_19862);
or UO_2413 (O_2413,N_19877,N_19874);
nand UO_2414 (O_2414,N_19916,N_19903);
xnor UO_2415 (O_2415,N_19997,N_19988);
and UO_2416 (O_2416,N_19979,N_19865);
nor UO_2417 (O_2417,N_19935,N_19929);
xor UO_2418 (O_2418,N_19926,N_19928);
nand UO_2419 (O_2419,N_19930,N_19956);
nor UO_2420 (O_2420,N_19922,N_19959);
nand UO_2421 (O_2421,N_19944,N_19855);
nand UO_2422 (O_2422,N_19977,N_19941);
and UO_2423 (O_2423,N_19966,N_19962);
nand UO_2424 (O_2424,N_19884,N_19973);
nand UO_2425 (O_2425,N_19896,N_19987);
xor UO_2426 (O_2426,N_19852,N_19912);
nor UO_2427 (O_2427,N_19991,N_19959);
and UO_2428 (O_2428,N_19963,N_19887);
and UO_2429 (O_2429,N_19962,N_19883);
and UO_2430 (O_2430,N_19883,N_19876);
nor UO_2431 (O_2431,N_19889,N_19928);
and UO_2432 (O_2432,N_19987,N_19902);
and UO_2433 (O_2433,N_19998,N_19864);
xor UO_2434 (O_2434,N_19867,N_19841);
nor UO_2435 (O_2435,N_19996,N_19944);
xor UO_2436 (O_2436,N_19868,N_19975);
xnor UO_2437 (O_2437,N_19883,N_19930);
xnor UO_2438 (O_2438,N_19845,N_19957);
nor UO_2439 (O_2439,N_19858,N_19986);
or UO_2440 (O_2440,N_19990,N_19973);
nor UO_2441 (O_2441,N_19990,N_19941);
xor UO_2442 (O_2442,N_19998,N_19887);
xor UO_2443 (O_2443,N_19965,N_19843);
xnor UO_2444 (O_2444,N_19858,N_19978);
or UO_2445 (O_2445,N_19880,N_19860);
xor UO_2446 (O_2446,N_19855,N_19921);
or UO_2447 (O_2447,N_19849,N_19861);
or UO_2448 (O_2448,N_19903,N_19985);
and UO_2449 (O_2449,N_19871,N_19919);
and UO_2450 (O_2450,N_19941,N_19937);
nand UO_2451 (O_2451,N_19873,N_19997);
or UO_2452 (O_2452,N_19980,N_19860);
and UO_2453 (O_2453,N_19962,N_19991);
and UO_2454 (O_2454,N_19869,N_19932);
and UO_2455 (O_2455,N_19845,N_19843);
and UO_2456 (O_2456,N_19917,N_19847);
nand UO_2457 (O_2457,N_19944,N_19868);
and UO_2458 (O_2458,N_19862,N_19912);
xnor UO_2459 (O_2459,N_19897,N_19940);
xor UO_2460 (O_2460,N_19927,N_19936);
nand UO_2461 (O_2461,N_19977,N_19962);
xor UO_2462 (O_2462,N_19853,N_19901);
and UO_2463 (O_2463,N_19932,N_19971);
or UO_2464 (O_2464,N_19926,N_19959);
or UO_2465 (O_2465,N_19956,N_19998);
nor UO_2466 (O_2466,N_19898,N_19996);
xor UO_2467 (O_2467,N_19928,N_19869);
xor UO_2468 (O_2468,N_19949,N_19964);
and UO_2469 (O_2469,N_19915,N_19848);
nand UO_2470 (O_2470,N_19981,N_19854);
xor UO_2471 (O_2471,N_19901,N_19848);
nor UO_2472 (O_2472,N_19874,N_19945);
nand UO_2473 (O_2473,N_19980,N_19949);
or UO_2474 (O_2474,N_19881,N_19924);
nor UO_2475 (O_2475,N_19934,N_19884);
xnor UO_2476 (O_2476,N_19961,N_19848);
nor UO_2477 (O_2477,N_19869,N_19860);
or UO_2478 (O_2478,N_19918,N_19902);
or UO_2479 (O_2479,N_19914,N_19878);
nand UO_2480 (O_2480,N_19854,N_19944);
nor UO_2481 (O_2481,N_19861,N_19858);
nor UO_2482 (O_2482,N_19891,N_19930);
and UO_2483 (O_2483,N_19964,N_19933);
nand UO_2484 (O_2484,N_19919,N_19906);
and UO_2485 (O_2485,N_19865,N_19946);
and UO_2486 (O_2486,N_19940,N_19853);
and UO_2487 (O_2487,N_19959,N_19909);
nor UO_2488 (O_2488,N_19895,N_19967);
nor UO_2489 (O_2489,N_19974,N_19910);
nand UO_2490 (O_2490,N_19849,N_19865);
or UO_2491 (O_2491,N_19916,N_19932);
xnor UO_2492 (O_2492,N_19955,N_19846);
xnor UO_2493 (O_2493,N_19899,N_19852);
nand UO_2494 (O_2494,N_19918,N_19959);
nor UO_2495 (O_2495,N_19852,N_19908);
or UO_2496 (O_2496,N_19898,N_19961);
nand UO_2497 (O_2497,N_19934,N_19971);
and UO_2498 (O_2498,N_19920,N_19859);
xnor UO_2499 (O_2499,N_19980,N_19922);
endmodule