module basic_3000_30000_3500_15_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
and U0 (N_0,In_285,In_1418);
nor U1 (N_1,In_328,In_1702);
nor U2 (N_2,In_1431,In_463);
or U3 (N_3,In_2967,In_2737);
nand U4 (N_4,In_826,In_180);
nand U5 (N_5,In_791,In_1438);
and U6 (N_6,In_1447,In_1518);
nand U7 (N_7,In_2866,In_528);
nor U8 (N_8,In_1338,In_496);
xor U9 (N_9,In_1063,In_821);
nor U10 (N_10,In_777,In_2912);
or U11 (N_11,In_654,In_2342);
or U12 (N_12,In_1594,In_814);
xor U13 (N_13,In_346,In_558);
nand U14 (N_14,In_2131,In_686);
or U15 (N_15,In_2265,In_1358);
nand U16 (N_16,In_977,In_488);
xnor U17 (N_17,In_1632,In_1376);
or U18 (N_18,In_506,In_150);
and U19 (N_19,In_2464,In_790);
nand U20 (N_20,In_2685,In_416);
nand U21 (N_21,In_1432,In_2176);
or U22 (N_22,In_2144,In_667);
nand U23 (N_23,In_1955,In_2742);
and U24 (N_24,In_697,In_2593);
xnor U25 (N_25,In_2202,In_1283);
nor U26 (N_26,In_849,In_1295);
nand U27 (N_27,In_2903,In_1729);
nor U28 (N_28,In_1716,In_1787);
nor U29 (N_29,In_1224,In_342);
xor U30 (N_30,In_194,In_860);
or U31 (N_31,In_1739,In_234);
or U32 (N_32,In_2816,In_2611);
xor U33 (N_33,In_728,In_803);
xor U34 (N_34,In_522,In_934);
nor U35 (N_35,In_1010,In_2288);
or U36 (N_36,In_2774,In_2802);
nand U37 (N_37,In_2601,In_2378);
nand U38 (N_38,In_754,In_337);
xor U39 (N_39,In_1348,In_2318);
and U40 (N_40,In_794,In_1895);
and U41 (N_41,In_1225,In_1142);
or U42 (N_42,In_913,In_73);
or U43 (N_43,In_2430,In_763);
xor U44 (N_44,In_785,In_2920);
xor U45 (N_45,In_321,In_169);
or U46 (N_46,In_1377,In_8);
nor U47 (N_47,In_89,In_502);
xor U48 (N_48,In_2103,In_1948);
nand U49 (N_49,In_1782,In_835);
nand U50 (N_50,In_2456,In_2840);
or U51 (N_51,In_2827,In_2814);
and U52 (N_52,In_751,In_1152);
nand U53 (N_53,In_157,In_2418);
nor U54 (N_54,In_2348,In_1725);
xnor U55 (N_55,In_2076,In_64);
nor U56 (N_56,In_525,In_1000);
nand U57 (N_57,In_1004,In_901);
or U58 (N_58,In_2600,In_2587);
or U59 (N_59,In_415,In_1665);
nor U60 (N_60,In_569,In_607);
nor U61 (N_61,In_943,In_348);
nand U62 (N_62,In_1459,In_1083);
nor U63 (N_63,In_795,In_1668);
or U64 (N_64,In_891,In_1513);
xor U65 (N_65,In_1841,In_2436);
xor U66 (N_66,In_1700,In_244);
nor U67 (N_67,In_131,In_1324);
nand U68 (N_68,In_762,In_2235);
nor U69 (N_69,In_2934,In_2386);
nor U70 (N_70,In_2706,In_465);
nand U71 (N_71,In_355,In_2838);
or U72 (N_72,In_461,In_1687);
and U73 (N_73,In_2639,In_1412);
or U74 (N_74,In_2129,In_322);
or U75 (N_75,In_1918,In_2579);
nor U76 (N_76,In_1273,In_2673);
nor U77 (N_77,In_2613,In_1652);
nor U78 (N_78,In_2495,In_2505);
nand U79 (N_79,In_1608,In_2511);
and U80 (N_80,In_2240,In_1906);
nor U81 (N_81,In_1504,In_112);
and U82 (N_82,In_2382,In_482);
and U83 (N_83,In_1118,In_166);
nand U84 (N_84,In_2198,In_231);
nand U85 (N_85,In_725,In_1603);
nor U86 (N_86,In_2628,In_805);
or U87 (N_87,In_290,In_393);
and U88 (N_88,In_1969,In_1034);
nand U89 (N_89,In_1831,In_2638);
nor U90 (N_90,In_772,In_2224);
or U91 (N_91,In_1445,In_1434);
or U92 (N_92,In_1585,In_1744);
nand U93 (N_93,In_1396,In_1096);
or U94 (N_94,In_1139,In_1171);
or U95 (N_95,In_969,In_1243);
nor U96 (N_96,In_292,In_864);
or U97 (N_97,In_2729,In_707);
and U98 (N_98,In_1961,In_2010);
nand U99 (N_99,In_1014,In_656);
xnor U100 (N_100,In_1367,In_2151);
nand U101 (N_101,In_2463,In_638);
xnor U102 (N_102,In_1884,In_865);
or U103 (N_103,In_1277,In_2126);
or U104 (N_104,In_1202,In_513);
nand U105 (N_105,In_926,In_1487);
and U106 (N_106,In_1246,In_1127);
nand U107 (N_107,In_2405,In_975);
nand U108 (N_108,In_530,In_1631);
nand U109 (N_109,In_916,In_1439);
nand U110 (N_110,In_678,In_2991);
nor U111 (N_111,In_2584,In_1892);
or U112 (N_112,In_1670,In_2283);
nor U113 (N_113,In_2455,In_1065);
nand U114 (N_114,In_2525,In_2752);
and U115 (N_115,In_626,In_640);
xnor U116 (N_116,In_2330,In_771);
or U117 (N_117,In_491,In_1470);
or U118 (N_118,In_2023,In_1592);
or U119 (N_119,In_474,In_1644);
nand U120 (N_120,In_1714,In_1521);
xnor U121 (N_121,In_2458,In_159);
xnor U122 (N_122,In_2810,In_2796);
xor U123 (N_123,In_382,In_6);
and U124 (N_124,In_1320,In_2401);
nor U125 (N_125,In_120,In_389);
nand U126 (N_126,In_957,In_2243);
xnor U127 (N_127,In_295,In_451);
nand U128 (N_128,In_190,In_999);
or U129 (N_129,In_1076,In_178);
nor U130 (N_130,In_433,In_2732);
nor U131 (N_131,In_1617,In_2947);
nand U132 (N_132,In_22,In_2360);
nor U133 (N_133,In_1797,In_2755);
xnor U134 (N_134,In_1624,In_2085);
and U135 (N_135,In_879,In_475);
nand U136 (N_136,In_1336,In_1270);
xor U137 (N_137,In_1872,In_1828);
nor U138 (N_138,In_1168,In_619);
xor U139 (N_139,In_2294,In_1941);
nor U140 (N_140,In_2583,In_570);
xor U141 (N_141,In_761,In_2434);
nand U142 (N_142,In_1741,In_1692);
and U143 (N_143,In_1073,In_1005);
nor U144 (N_144,In_2645,In_13);
or U145 (N_145,In_2177,In_1241);
xnor U146 (N_146,In_1071,In_2306);
or U147 (N_147,In_1141,In_714);
and U148 (N_148,In_1537,In_1512);
nand U149 (N_149,In_1369,In_1253);
nor U150 (N_150,In_2258,In_2052);
xnor U151 (N_151,In_2334,In_2194);
xor U152 (N_152,In_2139,In_1478);
and U153 (N_153,In_224,In_1162);
and U154 (N_154,In_302,In_1737);
xnor U155 (N_155,In_705,In_2345);
and U156 (N_156,In_2766,In_1813);
nor U157 (N_157,In_137,In_153);
or U158 (N_158,In_1688,In_2409);
or U159 (N_159,In_657,In_775);
nor U160 (N_160,In_2309,In_1134);
and U161 (N_161,In_552,In_1068);
nand U162 (N_162,In_1102,In_2536);
nor U163 (N_163,In_12,In_2313);
nand U164 (N_164,In_2308,In_2417);
or U165 (N_165,In_1238,In_1934);
nor U166 (N_166,In_2806,In_127);
nand U167 (N_167,In_521,In_642);
and U168 (N_168,In_1380,In_418);
nor U169 (N_169,In_1720,In_2678);
nand U170 (N_170,In_870,In_2736);
or U171 (N_171,In_294,In_769);
xor U172 (N_172,In_1764,In_2359);
nor U173 (N_173,In_1183,In_130);
and U174 (N_174,In_1953,In_262);
nand U175 (N_175,In_874,In_779);
nand U176 (N_176,In_2841,In_1777);
nor U177 (N_177,In_1494,In_177);
xnor U178 (N_178,In_1411,In_2038);
nor U179 (N_179,In_1448,In_129);
nor U180 (N_180,In_2159,In_2280);
and U181 (N_181,In_1458,In_398);
nand U182 (N_182,In_2670,In_1266);
and U183 (N_183,In_1981,In_2233);
or U184 (N_184,In_2162,In_350);
nor U185 (N_185,In_1811,In_2260);
nand U186 (N_186,In_1900,In_2963);
or U187 (N_187,In_2797,In_1593);
nand U188 (N_188,In_2461,In_457);
and U189 (N_189,In_1482,In_435);
nor U190 (N_190,In_941,In_2142);
nor U191 (N_191,In_2343,In_2237);
nor U192 (N_192,In_1163,In_571);
nor U193 (N_193,In_812,In_1776);
xnor U194 (N_194,In_397,In_1379);
xor U195 (N_195,In_524,In_223);
or U196 (N_196,In_2270,In_1685);
xnor U197 (N_197,In_179,In_1676);
xnor U198 (N_198,In_1326,In_2);
nand U199 (N_199,In_968,In_2962);
nand U200 (N_200,In_989,In_1755);
xor U201 (N_201,In_2094,In_746);
nor U202 (N_202,In_1200,In_2890);
nor U203 (N_203,In_2484,In_2384);
nand U204 (N_204,In_1347,In_1052);
and U205 (N_205,In_2119,In_43);
or U206 (N_206,In_920,In_1192);
nand U207 (N_207,In_1929,In_2508);
nor U208 (N_208,In_2834,In_2435);
nor U209 (N_209,In_2217,In_2146);
nand U210 (N_210,In_2366,In_661);
nor U211 (N_211,In_2250,In_2900);
xor U212 (N_212,In_1852,In_2077);
and U213 (N_213,In_454,In_2823);
xnor U214 (N_214,In_1097,In_550);
xnor U215 (N_215,In_584,In_1977);
xnor U216 (N_216,In_1115,In_2896);
nand U217 (N_217,In_1552,In_2189);
and U218 (N_218,In_26,In_15);
nor U219 (N_219,In_395,In_630);
nand U220 (N_220,In_2067,In_2652);
and U221 (N_221,In_854,In_2376);
or U222 (N_222,In_2744,In_119);
nor U223 (N_223,In_2560,In_1613);
or U224 (N_224,In_287,In_2468);
nand U225 (N_225,In_1706,In_2878);
and U226 (N_226,In_843,In_1511);
or U227 (N_227,In_408,In_1920);
and U228 (N_228,In_2748,In_1765);
xnor U229 (N_229,In_2995,In_2949);
and U230 (N_230,In_2481,In_2355);
and U231 (N_231,In_2447,In_50);
nand U232 (N_232,In_2311,In_1164);
and U233 (N_233,In_2234,In_1230);
xor U234 (N_234,In_238,In_226);
nand U235 (N_235,In_1580,In_855);
nand U236 (N_236,In_2474,In_1337);
and U237 (N_237,In_2801,In_2315);
xor U238 (N_238,In_2341,In_1566);
nand U239 (N_239,In_1880,In_1467);
nor U240 (N_240,In_272,In_31);
xnor U241 (N_241,In_2494,In_2178);
or U242 (N_242,In_978,In_2501);
and U243 (N_243,In_611,In_2180);
and U244 (N_244,In_487,In_721);
and U245 (N_245,In_1849,In_251);
nor U246 (N_246,In_1736,In_1393);
xnor U247 (N_247,In_1529,In_2502);
and U248 (N_248,In_799,In_1444);
xor U249 (N_249,In_1078,In_1159);
nand U250 (N_250,In_2116,In_690);
nand U251 (N_251,In_1589,In_1007);
xor U252 (N_252,In_930,In_2066);
and U253 (N_253,In_2192,In_1008);
and U254 (N_254,In_756,In_49);
and U255 (N_255,In_2822,In_2205);
nor U256 (N_256,In_28,In_2867);
nand U257 (N_257,In_192,In_1032);
xor U258 (N_258,In_2338,In_420);
or U259 (N_259,In_501,In_2413);
nor U260 (N_260,In_737,In_875);
xor U261 (N_261,In_1098,In_745);
nand U262 (N_262,In_2072,In_1724);
nand U263 (N_263,In_2941,In_1313);
nand U264 (N_264,In_1302,In_206);
or U265 (N_265,In_2493,In_2677);
xnor U266 (N_266,In_1888,In_2124);
or U267 (N_267,In_2546,In_1633);
nor U268 (N_268,In_586,In_1796);
xnor U269 (N_269,In_175,In_2985);
nor U270 (N_270,In_1721,In_441);
nand U271 (N_271,In_2016,In_1505);
nand U272 (N_272,In_2290,In_442);
or U273 (N_273,In_2470,In_743);
xor U274 (N_274,In_1229,In_1244);
xnor U275 (N_275,In_1166,In_554);
xor U276 (N_276,In_815,In_1681);
and U277 (N_277,In_593,In_1500);
and U278 (N_278,In_2438,In_2286);
or U279 (N_279,In_1426,In_649);
or U280 (N_280,In_1562,In_1384);
nor U281 (N_281,In_2263,In_2728);
or U282 (N_282,In_2113,In_720);
nor U283 (N_283,In_2305,In_123);
or U284 (N_284,In_214,In_2354);
nor U285 (N_285,In_2577,In_537);
nor U286 (N_286,In_921,In_724);
xnor U287 (N_287,In_2731,In_476);
or U288 (N_288,In_2325,In_92);
nand U289 (N_289,In_1294,In_1218);
nor U290 (N_290,In_1801,In_2689);
xnor U291 (N_291,In_77,In_1194);
or U292 (N_292,In_1824,In_425);
and U293 (N_293,In_2506,In_967);
nor U294 (N_294,In_198,In_2292);
xnor U295 (N_295,In_1655,In_2363);
nand U296 (N_296,In_1758,In_766);
or U297 (N_297,In_2623,In_1323);
or U298 (N_298,In_1417,In_541);
xnor U299 (N_299,In_2765,In_819);
nor U300 (N_300,In_1084,In_1414);
or U301 (N_301,In_635,In_47);
nand U302 (N_302,In_2693,In_10);
nor U303 (N_303,In_1029,In_1406);
or U304 (N_304,In_1922,In_1258);
xnor U305 (N_305,In_1709,In_4);
or U306 (N_306,In_1648,In_716);
and U307 (N_307,In_1345,In_712);
nand U308 (N_308,In_2929,In_2231);
and U309 (N_309,In_2046,In_117);
xnor U310 (N_310,In_1025,In_1394);
and U311 (N_311,In_1666,In_2968);
or U312 (N_312,In_1835,In_2431);
or U313 (N_313,In_986,In_2884);
xor U314 (N_314,In_1599,In_2655);
nand U315 (N_315,In_274,In_776);
or U316 (N_316,In_2711,In_2937);
nand U317 (N_317,In_2479,In_1059);
xnor U318 (N_318,In_1060,In_1208);
and U319 (N_319,In_796,In_1859);
xnor U320 (N_320,In_1196,In_973);
nor U321 (N_321,In_237,In_2277);
or U322 (N_322,In_2065,In_1310);
and U323 (N_323,In_1278,In_1667);
nor U324 (N_324,In_1672,In_1003);
or U325 (N_325,In_878,In_316);
nand U326 (N_326,In_464,In_2559);
and U327 (N_327,In_412,In_2317);
nand U328 (N_328,In_1460,In_1826);
nor U329 (N_329,In_1983,In_2870);
xnor U330 (N_330,In_1501,In_1484);
or U331 (N_331,In_1368,In_2388);
nor U332 (N_332,In_1420,In_514);
nand U333 (N_333,In_392,In_1174);
nand U334 (N_334,In_1534,In_813);
nand U335 (N_335,In_1863,In_2648);
nor U336 (N_336,In_1307,In_2998);
xnor U337 (N_337,In_1693,In_2002);
nand U338 (N_338,In_2381,In_2471);
or U339 (N_339,In_1120,In_1763);
and U340 (N_340,In_825,In_1561);
and U341 (N_341,In_2279,In_1752);
and U342 (N_342,In_2888,In_252);
nor U343 (N_343,In_1261,In_2799);
nand U344 (N_344,In_623,In_468);
nand U345 (N_345,In_1247,In_146);
xor U346 (N_346,In_2757,In_1937);
nand U347 (N_347,In_2773,In_2905);
nor U348 (N_348,In_1611,In_2996);
nand U349 (N_349,In_257,In_2984);
xnor U350 (N_350,In_145,In_2157);
or U351 (N_351,In_844,In_1352);
or U352 (N_352,In_2893,In_1694);
xnor U353 (N_353,In_1292,In_161);
xor U354 (N_354,In_1287,In_125);
nand U355 (N_355,In_1496,In_232);
or U356 (N_356,In_1738,In_1893);
nor U357 (N_357,In_200,In_2898);
and U358 (N_358,In_734,In_1228);
xor U359 (N_359,In_405,In_2931);
or U360 (N_360,In_1242,In_2775);
nand U361 (N_361,In_2102,In_427);
nand U362 (N_362,In_1495,In_256);
nor U363 (N_363,In_2276,In_1933);
and U364 (N_364,In_2246,In_869);
or U365 (N_365,In_665,In_953);
and U366 (N_366,In_1201,In_1104);
and U367 (N_367,In_2674,In_1108);
and U368 (N_368,In_2475,In_917);
and U369 (N_369,In_1361,In_1923);
or U370 (N_370,In_1992,In_2244);
xnor U371 (N_371,In_1802,In_1213);
nand U372 (N_372,In_1645,In_1371);
nor U373 (N_373,In_1753,In_1121);
or U374 (N_374,In_516,In_1761);
and U375 (N_375,In_80,In_2857);
and U376 (N_376,In_313,In_85);
nor U377 (N_377,In_163,In_2120);
and U378 (N_378,In_2022,In_1601);
or U379 (N_379,In_333,In_2078);
nor U380 (N_380,In_2758,In_2156);
and U381 (N_381,In_426,In_663);
nand U382 (N_382,In_1772,In_1891);
and U383 (N_383,In_1359,In_109);
nor U384 (N_384,In_152,In_559);
and U385 (N_385,In_1587,In_1309);
xor U386 (N_386,In_903,In_1205);
and U387 (N_387,In_2125,In_789);
xnor U388 (N_388,In_651,In_2961);
nor U389 (N_389,In_460,In_2203);
or U390 (N_390,In_2873,In_172);
or U391 (N_391,In_543,In_1231);
and U392 (N_392,In_171,In_2432);
xnor U393 (N_393,In_2295,In_1269);
or U394 (N_394,In_2549,In_1179);
and U395 (N_395,In_738,In_360);
nand U396 (N_396,In_1113,In_2186);
and U397 (N_397,In_332,In_240);
nor U398 (N_398,In_1442,In_2974);
or U399 (N_399,In_715,In_2015);
nor U400 (N_400,In_2252,In_347);
or U401 (N_401,In_858,In_2933);
xnor U402 (N_402,In_2112,In_1492);
xor U403 (N_403,In_1701,In_1869);
nor U404 (N_404,In_3,In_1732);
and U405 (N_405,In_594,In_431);
xor U406 (N_406,In_2589,In_2695);
nand U407 (N_407,In_383,In_1583);
and U408 (N_408,In_792,In_1086);
and U409 (N_409,In_2886,In_2020);
or U410 (N_410,In_480,In_1173);
and U411 (N_411,In_281,In_1223);
or U412 (N_412,In_2459,In_1605);
or U413 (N_413,In_1952,In_1082);
xnor U414 (N_414,In_2513,In_1968);
nand U415 (N_415,In_1209,In_1629);
and U416 (N_416,In_1651,In_208);
nand U417 (N_417,In_1297,In_1827);
and U418 (N_418,In_2939,In_24);
nand U419 (N_419,In_2724,In_2013);
nand U420 (N_420,In_691,In_2364);
or U421 (N_421,In_2740,In_2412);
nand U422 (N_422,In_492,In_1069);
xnor U423 (N_423,In_2383,In_582);
nand U424 (N_424,In_2666,In_915);
nor U425 (N_425,In_76,In_1669);
xor U426 (N_426,In_369,In_2457);
xor U427 (N_427,In_1733,In_181);
nor U428 (N_428,In_1040,In_2635);
nand U429 (N_429,In_669,In_2808);
nand U430 (N_430,In_1085,In_149);
xnor U431 (N_431,In_1885,In_2091);
and U432 (N_432,In_1938,In_2215);
or U433 (N_433,In_1836,In_1189);
nor U434 (N_434,In_371,In_99);
and U435 (N_435,In_413,In_1314);
and U436 (N_436,In_2168,In_2056);
xnor U437 (N_437,In_818,In_2352);
nand U438 (N_438,In_939,In_1680);
nand U439 (N_439,In_2289,In_2910);
and U440 (N_440,In_2811,In_2817);
and U441 (N_441,In_199,In_2956);
or U442 (N_442,In_1554,In_1964);
and U443 (N_443,In_882,In_373);
xnor U444 (N_444,In_1606,In_1107);
nand U445 (N_445,In_2096,In_627);
nor U446 (N_446,In_1346,In_905);
xor U447 (N_447,In_2298,In_2351);
and U448 (N_448,In_404,In_719);
xor U449 (N_449,In_1762,In_259);
nor U450 (N_450,In_1564,In_1172);
or U451 (N_451,In_2642,In_2357);
xor U452 (N_452,In_2406,In_2444);
and U453 (N_453,In_250,In_1112);
nand U454 (N_454,In_2656,In_1017);
nand U455 (N_455,In_1105,In_1507);
nand U456 (N_456,In_83,In_1461);
nor U457 (N_457,In_2946,In_440);
and U458 (N_458,In_331,In_2644);
nor U459 (N_459,In_741,In_2966);
xnor U460 (N_460,In_1945,In_2885);
and U461 (N_461,In_338,In_1009);
nor U462 (N_462,In_729,In_2171);
or U463 (N_463,In_1786,In_2173);
and U464 (N_464,In_1609,In_1577);
or U465 (N_465,In_1404,In_141);
nand U466 (N_466,In_2894,In_1449);
xor U467 (N_467,In_2251,In_1905);
xnor U468 (N_468,In_2271,In_538);
xor U469 (N_469,In_1671,In_2195);
and U470 (N_470,In_2622,In_1541);
xor U471 (N_471,In_2738,In_1234);
nor U472 (N_472,In_1865,In_1902);
or U473 (N_473,In_2682,In_2365);
nand U474 (N_474,In_539,In_1590);
and U475 (N_475,In_1597,In_2483);
or U476 (N_476,In_2230,In_1425);
nor U477 (N_477,In_2665,In_2183);
or U478 (N_478,In_2410,In_1144);
nor U479 (N_479,In_2148,In_2981);
and U480 (N_480,In_1019,In_2404);
nor U481 (N_481,In_2953,In_1128);
nor U482 (N_482,In_1704,In_1457);
and U483 (N_483,In_1153,In_60);
xnor U484 (N_484,In_2372,In_271);
nor U485 (N_485,In_1304,In_2637);
nor U486 (N_486,In_1727,In_2904);
or U487 (N_487,In_2557,In_960);
xnor U488 (N_488,In_1110,In_1129);
xor U489 (N_489,In_555,In_2727);
xor U490 (N_490,In_608,In_1634);
and U491 (N_491,In_1532,In_2837);
nand U492 (N_492,In_1976,In_1756);
nor U493 (N_493,In_113,In_1436);
and U494 (N_494,In_48,In_804);
nand U495 (N_495,In_2371,In_800);
nor U496 (N_496,In_2854,In_1176);
and U497 (N_497,In_2080,In_2043);
nor U498 (N_498,In_185,In_86);
and U499 (N_499,In_2293,In_2597);
or U500 (N_500,In_2641,In_1503);
and U501 (N_501,In_2005,In_1871);
and U502 (N_502,In_134,In_101);
nand U503 (N_503,In_600,In_1641);
xnor U504 (N_504,In_2069,In_363);
or U505 (N_505,In_1781,In_1822);
or U506 (N_506,In_811,In_648);
nand U507 (N_507,In_18,In_523);
nor U508 (N_508,In_708,In_622);
nor U509 (N_509,In_573,In_2442);
or U510 (N_510,In_1186,In_907);
nor U511 (N_511,In_1474,In_1889);
xnor U512 (N_512,In_1881,In_1993);
nand U513 (N_513,In_293,In_2190);
nand U514 (N_514,In_1300,In_2979);
nand U515 (N_515,In_381,In_327);
and U516 (N_516,In_2952,In_1257);
xor U517 (N_517,In_1039,In_1028);
xnor U518 (N_518,In_1049,In_1717);
nand U519 (N_519,In_2092,In_2701);
nor U520 (N_520,In_82,In_2696);
and U521 (N_521,In_115,In_1628);
nand U522 (N_522,In_659,In_2296);
nor U523 (N_523,In_515,In_1169);
or U524 (N_524,In_2741,In_2555);
xnor U525 (N_525,In_836,In_2667);
or U526 (N_526,In_2167,In_16);
or U527 (N_527,In_510,In_2539);
and U528 (N_528,In_2024,In_2692);
nor U529 (N_529,In_2218,In_409);
xnor U530 (N_530,In_138,In_1921);
nor U531 (N_531,In_985,In_155);
and U532 (N_532,In_2828,In_1623);
or U533 (N_533,In_2503,In_2662);
or U534 (N_534,In_1473,In_773);
xnor U535 (N_535,In_1077,In_1464);
xor U536 (N_536,In_2489,In_253);
nor U537 (N_537,In_107,In_2895);
xnor U538 (N_538,In_1227,In_1095);
and U539 (N_539,In_2763,In_1264);
nor U540 (N_540,In_824,In_650);
nor U541 (N_541,In_2007,In_2118);
or U542 (N_542,In_1678,In_703);
and U543 (N_543,In_2344,In_1854);
nor U544 (N_544,In_1,In_2747);
xnor U545 (N_545,In_2193,In_2681);
xor U546 (N_546,In_946,In_2115);
and U547 (N_547,In_2165,In_410);
nor U548 (N_548,In_572,In_1991);
xnor U549 (N_549,In_580,In_2544);
or U550 (N_550,In_505,In_438);
xor U551 (N_551,In_861,In_2594);
and U552 (N_552,In_1240,In_7);
and U553 (N_553,In_616,In_1958);
nor U554 (N_554,In_1821,In_2718);
or U555 (N_555,In_1850,In_197);
nand U556 (N_556,In_2958,In_2543);
and U557 (N_557,In_1747,In_1020);
or U558 (N_558,In_209,In_2831);
and U559 (N_559,In_1401,In_1626);
xnor U560 (N_560,In_997,In_2490);
or U561 (N_561,In_618,In_126);
xnor U562 (N_562,In_2255,In_341);
and U563 (N_563,In_1730,In_2362);
nand U564 (N_564,In_2429,In_2921);
and U565 (N_565,In_2184,In_401);
nand U566 (N_566,In_1960,In_2709);
or U567 (N_567,In_1703,In_2319);
or U568 (N_568,In_2856,In_63);
xnor U569 (N_569,In_2045,In_890);
or U570 (N_570,In_1935,In_2440);
nand U571 (N_571,In_1388,In_1663);
xnor U572 (N_572,In_1012,In_191);
xor U573 (N_573,In_2993,In_2138);
nand U574 (N_574,In_1090,In_2390);
nor U575 (N_575,In_1252,In_2730);
xor U576 (N_576,In_2507,In_2196);
nor U577 (N_577,In_17,In_2303);
nand U578 (N_578,In_2819,In_2328);
and U579 (N_579,In_2573,In_992);
or U580 (N_580,In_2919,In_888);
xor U581 (N_581,In_2331,In_2879);
xnor U582 (N_582,In_2152,In_2267);
nand U583 (N_583,In_2812,In_912);
nor U584 (N_584,In_2547,In_1058);
xnor U585 (N_585,In_1894,In_1614);
xor U586 (N_586,In_1259,In_2954);
and U587 (N_587,In_2710,In_254);
nor U588 (N_588,In_1896,In_852);
nor U589 (N_589,In_2874,In_2326);
and U590 (N_590,In_1595,In_1357);
xor U591 (N_591,In_1804,In_41);
nor U592 (N_592,In_949,In_311);
or U593 (N_593,In_1250,In_300);
nand U594 (N_594,In_1351,In_1114);
xor U595 (N_595,In_2104,In_2708);
xor U596 (N_596,In_1116,In_453);
xor U597 (N_597,In_1639,In_2935);
or U598 (N_598,In_1317,In_2445);
nand U599 (N_599,In_1398,In_1080);
nand U600 (N_600,In_1180,In_391);
xnor U601 (N_601,In_1546,In_1050);
nor U602 (N_602,In_2049,In_2705);
and U603 (N_603,In_2735,In_105);
and U604 (N_604,In_1033,In_1638);
nand U605 (N_605,In_2088,In_1553);
or U606 (N_606,In_1220,In_1908);
or U607 (N_607,In_764,In_329);
nor U608 (N_608,In_2163,In_2524);
xnor U609 (N_609,In_2723,In_439);
nand U610 (N_610,In_1378,In_1572);
or U611 (N_611,In_1087,In_2304);
or U612 (N_612,In_1178,In_589);
nor U613 (N_613,In_54,In_1137);
or U614 (N_614,In_1864,In_2522);
nor U615 (N_615,In_2721,In_1342);
nor U616 (N_616,In_494,In_857);
and U617 (N_617,In_2753,In_664);
or U618 (N_618,In_859,In_910);
and U619 (N_619,In_2554,In_1927);
nand U620 (N_620,In_1282,In_658);
or U621 (N_621,In_456,In_2169);
nor U622 (N_622,In_981,In_1520);
xnor U623 (N_623,In_1101,In_1111);
xor U624 (N_624,In_2809,In_1710);
nor U625 (N_625,In_2535,In_982);
or U626 (N_626,In_336,In_551);
or U627 (N_627,In_2262,In_788);
and U628 (N_628,In_55,In_330);
xnor U629 (N_629,In_2373,In_1555);
nor U630 (N_630,In_2229,In_1215);
and U631 (N_631,In_1967,In_1109);
and U632 (N_632,In_1980,In_151);
nor U633 (N_633,In_2241,In_1596);
xnor U634 (N_634,In_1463,In_590);
nor U635 (N_635,In_671,In_1939);
and U636 (N_636,In_1600,In_735);
nand U637 (N_637,In_2795,In_277);
or U638 (N_638,In_2245,In_2563);
nand U639 (N_639,In_599,In_357);
or U640 (N_640,In_604,In_345);
xor U641 (N_641,In_2017,In_1598);
nor U642 (N_642,In_1757,In_1508);
xnor U643 (N_643,In_2839,In_2687);
or U644 (N_644,In_1175,In_1878);
or U645 (N_645,In_1064,In_991);
and U646 (N_646,In_676,In_598);
nor U647 (N_647,In_1898,In_1079);
nand U648 (N_648,In_1198,In_2025);
and U649 (N_649,In_1416,In_780);
or U650 (N_650,In_216,In_1006);
and U651 (N_651,In_980,In_1847);
nor U652 (N_652,In_2562,In_46);
and U653 (N_653,In_2771,In_1604);
nand U654 (N_654,In_1497,In_317);
and U655 (N_655,In_591,In_196);
nand U656 (N_656,In_527,In_2164);
or U657 (N_657,In_2035,In_2266);
nand U658 (N_658,In_1267,In_1767);
or U659 (N_659,In_1851,In_1306);
nor U660 (N_660,In_2626,In_2054);
nand U661 (N_661,In_1479,In_1862);
nand U662 (N_662,In_566,In_900);
nor U663 (N_663,In_1998,In_770);
nand U664 (N_664,In_2282,In_2278);
xnor U665 (N_665,In_219,In_2784);
or U666 (N_666,In_1410,In_1131);
or U667 (N_667,In_560,In_2448);
xor U668 (N_668,In_1441,In_1321);
nor U669 (N_669,In_1092,In_2599);
xor U670 (N_670,In_1212,In_173);
or U671 (N_671,In_1745,In_2788);
or U672 (N_672,In_2604,In_834);
xnor U673 (N_673,In_1199,In_2647);
nand U674 (N_674,In_1191,In_2654);
nor U675 (N_675,In_692,In_87);
nor U676 (N_676,In_2683,In_2932);
nor U677 (N_677,In_2750,In_1773);
nand U678 (N_678,In_1932,In_1743);
or U679 (N_679,In_851,In_2565);
or U680 (N_680,In_2074,In_1588);
and U681 (N_681,In_2845,In_2123);
or U682 (N_682,In_2592,In_1182);
nand U683 (N_683,In_748,In_477);
nor U684 (N_684,In_318,In_1621);
nand U685 (N_685,In_2361,In_621);
xor U686 (N_686,In_1488,In_970);
and U687 (N_687,In_1316,In_2201);
nand U688 (N_688,In_1940,In_2605);
xor U689 (N_689,In_533,In_2284);
nor U690 (N_690,In_1924,In_1047);
nor U691 (N_691,In_1919,In_2454);
nand U692 (N_692,In_1957,In_2803);
and U693 (N_693,In_394,In_2485);
nor U694 (N_694,In_2712,In_696);
xor U695 (N_695,In_563,In_1392);
xnor U696 (N_696,In_38,In_2335);
nor U697 (N_697,In_1675,In_1103);
nor U698 (N_698,In_837,In_1569);
nand U699 (N_699,In_639,In_124);
nor U700 (N_700,In_1653,In_2117);
or U701 (N_701,In_1349,In_2400);
nor U702 (N_702,In_2369,In_1749);
nor U703 (N_703,In_1286,In_1048);
nor U704 (N_704,In_1547,In_2518);
nor U705 (N_705,In_1557,In_144);
and U706 (N_706,In_2392,In_750);
and U707 (N_707,In_221,In_187);
xor U708 (N_708,In_1185,In_2140);
xnor U709 (N_709,In_1053,In_2324);
or U710 (N_710,In_1062,In_111);
and U711 (N_711,In_1966,In_2358);
nand U712 (N_712,In_35,In_148);
or U713 (N_713,In_59,In_2150);
nor U714 (N_714,In_1853,In_2614);
nor U715 (N_715,In_679,In_2733);
and U716 (N_716,In_2624,In_578);
xor U717 (N_717,In_2346,In_2922);
nand U718 (N_718,In_104,In_2316);
nand U719 (N_719,In_248,In_531);
or U720 (N_720,In_1423,In_1002);
nor U721 (N_721,In_2777,In_176);
nor U722 (N_722,In_1271,In_1689);
nor U723 (N_723,In_675,In_2523);
xnor U724 (N_724,In_432,In_1657);
or U725 (N_725,In_2039,In_1126);
nor U726 (N_726,In_942,In_1462);
or U727 (N_727,In_1809,In_1548);
and U728 (N_728,In_1279,In_1057);
xnor U729 (N_729,In_2424,In_2813);
xor U730 (N_730,In_1235,In_188);
nor U731 (N_731,In_876,In_700);
xor U732 (N_732,In_2291,In_2063);
xnor U733 (N_733,In_2553,In_2210);
nand U734 (N_734,In_1181,In_2403);
nand U735 (N_735,In_2965,In_2496);
and U736 (N_736,In_455,In_2608);
xnor U737 (N_737,In_2122,In_2084);
or U738 (N_738,In_1481,In_1284);
xor U739 (N_739,In_755,In_227);
nand U740 (N_740,In_808,In_867);
or U741 (N_741,In_2862,In_2514);
and U742 (N_742,In_213,In_1823);
and U743 (N_743,In_998,In_632);
nand U744 (N_744,In_1799,In_2702);
nor U745 (N_745,In_565,In_585);
xor U746 (N_746,In_615,In_264);
nand U747 (N_747,In_2899,In_1942);
and U748 (N_748,In_2402,In_672);
xnor U749 (N_749,In_1293,In_2452);
nor U750 (N_750,In_2356,In_2135);
and U751 (N_751,In_2769,In_2994);
or U752 (N_752,In_2030,In_354);
nor U753 (N_753,In_1391,In_1237);
or U754 (N_754,In_1818,In_1697);
nor U755 (N_755,In_961,In_1879);
nor U756 (N_756,In_2659,In_2141);
nand U757 (N_757,In_2887,In_20);
nor U758 (N_758,In_423,In_893);
nand U759 (N_759,In_225,In_2876);
and U760 (N_760,In_417,In_2191);
nor U761 (N_761,In_940,In_2913);
and U762 (N_762,In_1407,In_2545);
nor U763 (N_763,In_445,In_2337);
nor U764 (N_764,In_2242,In_948);
nand U765 (N_765,In_702,In_1856);
xnor U766 (N_766,In_2745,In_2399);
xor U767 (N_767,In_39,In_2582);
nor U768 (N_768,In_2699,In_1088);
and U769 (N_769,In_1331,In_140);
xnor U770 (N_770,In_1842,In_2690);
or U771 (N_771,In_269,In_37);
xor U772 (N_772,In_2302,In_2081);
or U773 (N_773,In_2570,In_2794);
nand U774 (N_774,In_908,In_1015);
xor U775 (N_775,In_617,In_2537);
xnor U776 (N_776,In_862,In_1622);
nand U777 (N_777,In_1021,In_955);
or U778 (N_778,In_1066,In_1045);
xor U779 (N_779,In_1876,In_1263);
or U780 (N_780,In_603,In_614);
and U781 (N_781,In_1456,In_1866);
or U782 (N_782,In_1195,In_1914);
nor U783 (N_783,In_2830,In_2101);
or U784 (N_784,In_1798,In_2086);
xnor U785 (N_785,In_2349,In_1586);
xnor U786 (N_786,In_75,In_1046);
nor U787 (N_787,In_2155,In_2098);
nand U788 (N_788,In_1031,In_2586);
xnor U789 (N_789,In_1719,In_53);
and U790 (N_790,In_765,In_1754);
and U791 (N_791,In_1437,In_1452);
and U792 (N_792,In_823,In_2848);
and U793 (N_793,In_1844,In_212);
or U794 (N_794,In_2108,In_1089);
or U795 (N_795,In_2580,In_652);
and U796 (N_796,In_713,In_1742);
nand U797 (N_797,In_2055,In_1576);
and U798 (N_798,In_2720,In_856);
nand U799 (N_799,In_485,In_1477);
xnor U800 (N_800,In_1299,In_1531);
nor U801 (N_801,In_1814,In_2672);
or U802 (N_802,In_1570,In_2492);
nor U803 (N_803,In_2465,In_1366);
and U804 (N_804,In_1022,In_1543);
nand U805 (N_805,In_935,In_1305);
xor U806 (N_806,In_881,In_2734);
xnor U807 (N_807,In_284,In_2509);
or U808 (N_808,In_2397,In_2487);
xor U809 (N_809,In_2609,In_1197);
nand U810 (N_810,In_740,In_2200);
nand U811 (N_811,In_579,In_1728);
or U812 (N_812,In_1542,In_801);
xnor U813 (N_813,In_2793,In_1551);
nand U814 (N_814,In_1343,In_534);
nor U815 (N_815,In_1216,In_1498);
xnor U816 (N_816,In_45,In_1711);
xor U817 (N_817,In_1158,In_526);
nand U818 (N_818,In_1239,In_634);
or U819 (N_819,In_2427,In_2925);
nor U820 (N_820,In_2411,In_2679);
xnor U821 (N_821,In_1429,In_2000);
xnor U822 (N_822,In_1808,In_2865);
xnor U823 (N_823,In_710,In_2232);
and U824 (N_824,In_67,In_1995);
nor U825 (N_825,In_1156,In_951);
or U826 (N_826,In_1734,In_242);
and U827 (N_827,In_1027,In_1760);
or U828 (N_828,In_1268,In_1794);
xor U829 (N_829,In_1860,In_2987);
nand U830 (N_830,In_1815,In_1123);
nor U831 (N_831,In_2497,In_1759);
nor U832 (N_832,In_2861,In_809);
nand U833 (N_833,In_2787,In_1962);
and U834 (N_834,In_1074,In_270);
nor U835 (N_835,In_42,In_1327);
nand U836 (N_836,In_2892,In_1820);
or U837 (N_837,In_1288,In_633);
and U838 (N_838,In_923,In_1916);
xor U839 (N_839,In_1803,In_1303);
nor U840 (N_840,In_362,In_233);
nand U841 (N_841,In_306,In_2147);
xnor U842 (N_842,In_139,In_613);
xor U843 (N_843,In_947,In_918);
or U844 (N_844,In_767,In_275);
xor U845 (N_845,In_2158,In_1713);
or U846 (N_846,In_2254,In_2488);
or U847 (N_847,In_797,In_631);
xnor U848 (N_848,In_732,In_609);
nor U849 (N_849,In_1790,In_2037);
xnor U850 (N_850,In_512,In_959);
nand U851 (N_851,In_928,In_1707);
or U852 (N_852,In_1399,In_1982);
and U853 (N_853,In_247,In_2707);
xnor U854 (N_854,In_1340,In_1325);
or U855 (N_855,In_2451,In_2408);
and U856 (N_856,In_868,In_2595);
and U857 (N_857,In_351,In_1930);
xor U858 (N_858,In_976,In_1536);
or U859 (N_859,In_1705,In_1677);
nand U860 (N_860,In_904,In_1731);
and U861 (N_861,In_1528,In_2527);
nor U862 (N_862,In_2477,In_2500);
and U863 (N_863,In_301,In_816);
and U864 (N_864,In_1540,In_165);
nand U865 (N_865,In_1016,In_303);
or U866 (N_866,In_984,In_807);
xnor U867 (N_867,In_1559,In_540);
nand U868 (N_868,In_1041,In_2686);
xor U869 (N_869,In_2923,In_2453);
nor U870 (N_870,In_1514,In_473);
xnor U871 (N_871,In_334,In_1026);
or U872 (N_872,In_1963,In_840);
nor U873 (N_873,In_863,In_2805);
or U874 (N_874,In_1450,In_370);
nor U875 (N_875,In_2955,In_1954);
xor U876 (N_876,In_2466,In_1499);
nand U877 (N_877,In_2650,In_2548);
or U878 (N_878,In_1490,In_268);
nand U879 (N_879,In_388,In_938);
xnor U880 (N_880,In_2815,In_2100);
nand U881 (N_881,In_32,In_1838);
nor U882 (N_882,In_2520,In_450);
or U883 (N_883,In_1533,In_2868);
nor U884 (N_884,In_1070,In_1779);
xnor U885 (N_885,In_2743,In_2073);
or U886 (N_886,In_1684,In_211);
nor U887 (N_887,In_116,In_1443);
nor U888 (N_888,In_760,In_1311);
nand U889 (N_889,In_1829,In_1903);
nor U890 (N_890,In_1409,In_1296);
nor U891 (N_891,In_1188,In_759);
and U892 (N_892,In_245,In_1055);
xor U893 (N_893,In_1226,In_265);
nand U894 (N_894,In_2079,In_1354);
xnor U895 (N_895,In_2882,In_508);
and U896 (N_896,In_1972,In_1094);
xor U897 (N_897,In_2498,In_950);
nand U898 (N_898,In_1285,In_706);
nor U899 (N_899,In_2990,In_340);
nor U900 (N_900,In_52,In_641);
and U901 (N_901,In_1578,In_1132);
or U902 (N_902,In_489,In_2846);
or U903 (N_903,In_829,In_1091);
nand U904 (N_904,In_2380,In_701);
and U905 (N_905,In_2907,In_1155);
xnor U906 (N_906,In_1769,In_97);
nand U907 (N_907,In_1466,In_898);
and U908 (N_908,In_2542,In_1329);
xnor U909 (N_909,In_1544,In_96);
or U910 (N_910,In_2620,In_583);
xnor U911 (N_911,In_2852,In_2825);
nand U912 (N_912,In_606,In_2336);
nand U913 (N_913,In_532,In_2790);
xnor U914 (N_914,In_927,In_1506);
or U915 (N_915,In_2964,In_974);
xnor U916 (N_916,In_964,In_2136);
or U917 (N_917,In_2786,In_143);
nand U918 (N_918,In_339,In_2864);
nor U919 (N_919,In_886,In_877);
nor U920 (N_920,In_1571,In_289);
xor U921 (N_921,In_1726,In_2467);
or U922 (N_922,In_1771,In_1373);
nand U923 (N_923,In_2110,In_1875);
nand U924 (N_924,In_2633,In_2719);
and U925 (N_925,In_1602,In_2897);
or U926 (N_926,In_2145,In_402);
xor U927 (N_927,In_2832,In_378);
or U928 (N_928,In_2658,In_2174);
or U929 (N_929,In_2726,In_288);
xnor U930 (N_930,In_2598,In_2578);
nor U931 (N_931,In_1615,In_2394);
nor U932 (N_932,In_1735,In_828);
or U933 (N_933,In_1718,In_757);
or U934 (N_934,In_832,In_2441);
or U935 (N_935,In_2375,In_2778);
nor U936 (N_936,In_2761,In_730);
nand U937 (N_937,In_1913,In_324);
or U938 (N_938,In_241,In_846);
or U939 (N_939,In_2216,In_1530);
nand U940 (N_940,In_486,In_399);
nor U941 (N_941,In_147,In_733);
nor U942 (N_942,In_1219,In_1117);
and U943 (N_943,In_1435,In_2090);
and U944 (N_944,In_1440,In_2206);
nor U945 (N_945,In_154,In_367);
nand U946 (N_946,In_1148,In_1845);
xor U947 (N_947,In_443,In_2591);
nor U948 (N_948,In_1428,In_1054);
nand U949 (N_949,In_2688,In_2651);
nor U950 (N_950,In_694,In_1999);
nand U951 (N_951,In_2491,In_1030);
and U952 (N_952,In_2029,In_467);
xor U953 (N_953,In_932,In_2307);
nor U954 (N_954,In_687,In_1951);
xnor U955 (N_955,In_2596,In_2285);
and U956 (N_956,In_1785,In_1928);
nand U957 (N_957,In_574,In_424);
or U958 (N_958,In_564,In_567);
xnor U959 (N_959,In_2379,In_535);
nor U960 (N_960,In_479,In_2333);
nand U961 (N_961,In_69,In_798);
or U962 (N_962,In_2552,In_2050);
nor U963 (N_963,In_1433,In_1335);
or U964 (N_964,In_1036,In_400);
or U965 (N_965,In_2473,In_1360);
and U966 (N_966,In_1151,In_1140);
nand U967 (N_967,In_2109,In_478);
xnor U968 (N_968,In_1682,In_2842);
and U969 (N_969,In_1793,In_802);
xor U970 (N_970,In_158,In_2847);
and U971 (N_971,In_2051,In_2099);
or U972 (N_972,In_2978,In_2754);
xor U973 (N_973,In_1581,In_2127);
nor U974 (N_974,In_2916,In_128);
and U975 (N_975,In_952,In_1125);
nor U976 (N_976,In_597,In_1451);
nor U977 (N_977,In_2154,In_62);
xnor U978 (N_978,In_2930,In_557);
and U979 (N_979,In_784,In_1698);
nor U980 (N_980,In_2209,In_718);
nor U981 (N_981,In_786,In_1255);
or U982 (N_982,In_2001,In_403);
nand U983 (N_983,In_549,In_1556);
nor U984 (N_984,In_298,In_544);
xnor U985 (N_985,In_499,In_2860);
nand U986 (N_986,In_352,In_193);
nor U987 (N_987,In_276,In_0);
and U988 (N_988,In_2197,In_1381);
nor U989 (N_989,In_1364,In_547);
or U990 (N_990,In_629,In_1538);
nor U991 (N_991,In_1915,In_2149);
nand U992 (N_992,In_344,In_364);
nand U993 (N_993,In_2739,In_1944);
or U994 (N_994,In_1043,In_2792);
nor U995 (N_995,In_693,In_1636);
xor U996 (N_996,In_1233,In_1341);
and U997 (N_997,In_2226,In_2936);
and U998 (N_998,In_2989,In_1912);
xnor U999 (N_999,In_684,In_1959);
nand U1000 (N_1000,In_944,In_1819);
xor U1001 (N_1001,In_2948,In_201);
nor U1002 (N_1002,In_1926,In_1650);
nor U1003 (N_1003,In_366,In_44);
and U1004 (N_1004,In_2031,In_2253);
nand U1005 (N_1005,In_1289,In_1509);
nor U1006 (N_1006,In_2880,In_1280);
nand U1007 (N_1007,In_2247,In_902);
nand U1008 (N_1008,In_2980,In_1843);
or U1009 (N_1009,In_1390,In_1917);
nor U1010 (N_1010,In_887,In_2636);
xnor U1011 (N_1011,In_2472,In_758);
nor U1012 (N_1012,In_308,In_972);
nor U1013 (N_1013,In_839,In_358);
xor U1014 (N_1014,In_282,In_2273);
xor U1015 (N_1015,In_466,In_1874);
and U1016 (N_1016,In_2918,In_106);
nand U1017 (N_1017,In_1832,In_2646);
and U1018 (N_1018,In_1422,In_1517);
or U1019 (N_1019,In_310,In_2625);
nand U1020 (N_1020,In_1298,In_1911);
xor U1021 (N_1021,In_830,In_1899);
nand U1022 (N_1022,In_100,In_2133);
nor U1023 (N_1023,In_1778,In_170);
nor U1024 (N_1024,In_2053,In_419);
and U1025 (N_1025,In_2510,In_529);
xor U1026 (N_1026,In_2576,In_2529);
nor U1027 (N_1027,In_279,In_1658);
and U1028 (N_1028,In_1281,In_2512);
nor U1029 (N_1029,In_2347,In_1910);
and U1030 (N_1030,In_688,In_1430);
xnor U1031 (N_1031,In_1413,In_66);
nand U1032 (N_1032,In_2618,In_1567);
nor U1033 (N_1033,In_711,In_1746);
nor U1034 (N_1034,In_2214,In_365);
or U1035 (N_1035,In_2004,In_2257);
xor U1036 (N_1036,In_897,In_312);
nor U1037 (N_1037,In_2439,In_2901);
xor U1038 (N_1038,In_2664,In_1526);
nor U1039 (N_1039,In_1419,In_2663);
or U1040 (N_1040,In_768,In_2643);
nand U1041 (N_1041,In_500,In_810);
nor U1042 (N_1042,In_1775,In_2630);
and U1043 (N_1043,In_1975,In_1591);
nor U1044 (N_1044,In_296,In_2019);
or U1045 (N_1045,In_81,In_646);
or U1046 (N_1046,In_1245,In_220);
nand U1047 (N_1047,In_2211,In_2983);
or U1048 (N_1048,In_1206,In_469);
nor U1049 (N_1049,In_749,In_1839);
or U1050 (N_1050,In_1984,In_845);
nor U1051 (N_1051,In_132,In_437);
and U1052 (N_1052,In_1037,In_561);
xnor U1053 (N_1053,In_1750,In_343);
xnor U1054 (N_1054,In_2208,In_2572);
or U1055 (N_1055,In_945,In_2420);
xor U1056 (N_1056,In_1136,In_1100);
or U1057 (N_1057,In_1522,In_848);
xor U1058 (N_1058,In_1855,In_853);
nand U1059 (N_1059,In_1861,In_2259);
or U1060 (N_1060,In_2619,In_601);
nand U1061 (N_1061,In_778,In_2261);
nand U1062 (N_1062,In_29,In_2915);
or U1063 (N_1063,In_2426,In_1989);
or U1064 (N_1064,In_2213,In_2028);
nand U1065 (N_1065,In_1318,In_2749);
nand U1066 (N_1066,In_1882,In_1943);
or U1067 (N_1067,In_2323,In_1403);
and U1068 (N_1068,In_1262,In_1332);
nor U1069 (N_1069,In_1674,In_2999);
nand U1070 (N_1070,In_2070,In_806);
nor U1071 (N_1071,In_84,In_1475);
and U1072 (N_1072,In_2389,In_752);
xor U1073 (N_1073,In_2181,In_2785);
xor U1074 (N_1074,In_2281,In_1483);
or U1075 (N_1075,In_2106,In_183);
nand U1076 (N_1076,In_263,In_2219);
nor U1077 (N_1077,In_2849,In_1978);
xor U1078 (N_1078,In_2881,In_717);
nand U1079 (N_1079,In_787,In_838);
nor U1080 (N_1080,In_2684,In_375);
nor U1081 (N_1081,In_1353,In_2634);
or U1082 (N_1082,In_51,In_2450);
nand U1083 (N_1083,In_1051,In_1664);
or U1084 (N_1084,In_2564,In_2717);
nor U1085 (N_1085,In_1365,In_353);
xnor U1086 (N_1086,In_2959,In_205);
or U1087 (N_1087,In_2715,In_260);
nor U1088 (N_1088,In_1035,In_1868);
xnor U1089 (N_1089,In_1099,In_581);
xor U1090 (N_1090,In_2287,In_2970);
and U1091 (N_1091,In_2804,In_1395);
nand U1092 (N_1092,In_2657,In_1217);
nand U1093 (N_1093,In_1154,In_2768);
or U1094 (N_1094,In_1146,In_1374);
and U1095 (N_1095,In_1372,In_2569);
or U1096 (N_1096,In_2264,In_2393);
and U1097 (N_1097,In_1886,In_9);
or U1098 (N_1098,In_114,In_602);
xor U1099 (N_1099,In_2855,In_2835);
and U1100 (N_1100,In_1662,In_680);
xor U1101 (N_1101,In_2008,In_65);
and U1102 (N_1102,In_307,In_595);
nand U1103 (N_1103,In_1751,In_1405);
or U1104 (N_1104,In_2301,In_1130);
nor U1105 (N_1105,In_2274,In_896);
nand U1106 (N_1106,In_517,In_747);
or U1107 (N_1107,In_2700,In_744);
nand U1108 (N_1108,In_1549,In_883);
xor U1109 (N_1109,In_1272,In_1160);
or U1110 (N_1110,In_168,In_1203);
nand U1111 (N_1111,In_452,In_286);
nor U1112 (N_1112,In_406,In_2575);
nand U1113 (N_1113,In_685,In_668);
nor U1114 (N_1114,In_1812,In_27);
nand U1115 (N_1115,In_1625,In_1397);
or U1116 (N_1116,In_2350,In_2504);
nor U1117 (N_1117,In_1149,In_2322);
or U1118 (N_1118,In_1986,In_255);
nand U1119 (N_1119,In_2850,In_1619);
xor U1120 (N_1120,In_1333,In_2924);
nor U1121 (N_1121,In_774,In_1476);
nand U1122 (N_1122,In_386,In_2047);
nor U1123 (N_1123,In_871,In_1620);
nor U1124 (N_1124,In_1312,In_1515);
and U1125 (N_1125,In_2058,In_503);
or U1126 (N_1126,In_1579,In_2694);
nand U1127 (N_1127,In_1690,In_1837);
xnor U1128 (N_1128,In_2175,In_1550);
xnor U1129 (N_1129,In_2538,In_2423);
xnor U1130 (N_1130,In_1907,In_68);
nor U1131 (N_1131,In_1389,In_736);
xnor U1132 (N_1132,In_215,In_588);
nand U1133 (N_1133,In_2482,In_2395);
nor U1134 (N_1134,In_723,In_966);
and U1135 (N_1135,In_1119,In_577);
and U1136 (N_1136,In_2928,In_361);
or U1137 (N_1137,In_545,In_1249);
nor U1138 (N_1138,In_283,In_1683);
or U1139 (N_1139,In_1956,In_507);
and U1140 (N_1140,In_372,In_1383);
and U1141 (N_1141,In_2982,In_195);
xnor U1142 (N_1142,In_1468,In_160);
xnor U1143 (N_1143,In_782,In_444);
nor U1144 (N_1144,In_988,In_447);
nand U1145 (N_1145,In_228,In_2516);
or U1146 (N_1146,In_273,In_1539);
or U1147 (N_1147,In_2612,In_156);
nor U1148 (N_1148,In_167,In_2574);
or U1149 (N_1149,In_2697,In_218);
or U1150 (N_1150,In_246,In_1770);
xnor U1151 (N_1151,In_2526,In_1276);
xnor U1152 (N_1152,In_1480,In_2225);
nor U1153 (N_1153,In_2764,In_873);
and U1154 (N_1154,In_979,In_33);
nand U1155 (N_1155,In_1565,In_2671);
and U1156 (N_1156,In_2188,In_1190);
nand U1157 (N_1157,In_2248,In_2691);
xnor U1158 (N_1158,In_493,In_2942);
nor U1159 (N_1159,In_1890,In_2824);
nor U1160 (N_1160,In_793,In_925);
and U1161 (N_1161,In_620,In_2661);
nor U1162 (N_1162,In_110,In_142);
xor U1163 (N_1163,In_1334,In_2275);
and U1164 (N_1164,In_2172,In_1453);
and U1165 (N_1165,In_2725,In_349);
xor U1166 (N_1166,In_820,In_2556);
xnor U1167 (N_1167,In_2869,In_2528);
and U1168 (N_1168,In_2032,In_1584);
nor U1169 (N_1169,In_1023,In_93);
or U1170 (N_1170,In_304,In_2071);
xnor U1171 (N_1171,In_2872,In_1563);
nand U1172 (N_1172,In_2973,In_2992);
or U1173 (N_1173,In_2875,In_1723);
and U1174 (N_1174,In_326,In_1167);
and U1175 (N_1175,In_1236,In_2877);
nor U1176 (N_1176,In_267,In_624);
nor U1177 (N_1177,In_1985,In_434);
nand U1178 (N_1178,In_1184,In_14);
nor U1179 (N_1179,In_384,In_885);
and U1180 (N_1180,In_2062,In_2669);
xnor U1181 (N_1181,In_872,In_118);
xnor U1182 (N_1182,In_1897,In_2268);
and U1183 (N_1183,In_922,In_2629);
and U1184 (N_1184,In_2798,In_2097);
or U1185 (N_1185,In_2704,In_562);
nor U1186 (N_1186,In_71,In_2977);
and U1187 (N_1187,In_990,In_1800);
or U1188 (N_1188,In_2770,In_2914);
and U1189 (N_1189,In_2212,In_266);
or U1190 (N_1190,In_2111,In_2460);
nor U1191 (N_1191,In_1858,In_1840);
or U1192 (N_1192,In_1901,In_1510);
and U1193 (N_1193,In_1165,In_2425);
and U1194 (N_1194,In_481,In_937);
or U1195 (N_1195,In_2329,In_1660);
xnor U1196 (N_1196,In_1024,In_504);
xor U1197 (N_1197,In_2960,In_2036);
xor U1198 (N_1198,In_243,In_2975);
and U1199 (N_1199,In_1408,In_956);
xnor U1200 (N_1200,In_2249,In_983);
nor U1201 (N_1201,In_2027,In_2478);
or U1202 (N_1202,In_2310,In_1319);
xor U1203 (N_1203,In_1883,In_2075);
and U1204 (N_1204,In_1616,In_2068);
nor U1205 (N_1205,In_2676,In_325);
and U1206 (N_1206,In_449,In_1768);
xnor U1207 (N_1207,In_2568,In_1931);
or U1208 (N_1208,In_727,In_1290);
nand U1209 (N_1209,In_2220,In_2179);
nor U1210 (N_1210,In_2781,In_2668);
and U1211 (N_1211,In_884,In_2532);
xnor U1212 (N_1212,In_1308,In_996);
xnor U1213 (N_1213,In_2476,In_446);
and U1214 (N_1214,In_1649,In_189);
and U1215 (N_1215,In_2610,In_1042);
nor U1216 (N_1216,In_677,In_1362);
xnor U1217 (N_1217,In_315,In_495);
nand U1218 (N_1218,In_470,In_2531);
nor U1219 (N_1219,In_2370,In_2844);
nand U1220 (N_1220,In_2541,In_21);
and U1221 (N_1221,In_1524,In_74);
xnor U1222 (N_1222,In_2780,In_1387);
nand U1223 (N_1223,In_895,In_1996);
nor U1224 (N_1224,In_850,In_831);
nor U1225 (N_1225,In_1427,In_2950);
or U1226 (N_1226,In_2581,In_1640);
nor U1227 (N_1227,In_2746,In_1712);
and U1228 (N_1228,In_1485,In_2926);
nand U1229 (N_1229,In_430,In_57);
nand U1230 (N_1230,In_61,In_1810);
and U1231 (N_1231,In_742,In_56);
or U1232 (N_1232,In_704,In_2199);
or U1233 (N_1233,In_1469,In_2836);
xor U1234 (N_1234,In_2986,In_2089);
nand U1235 (N_1235,In_1001,In_23);
or U1236 (N_1236,In_520,In_2550);
or U1237 (N_1237,In_217,In_2236);
nand U1238 (N_1238,In_2107,In_2377);
nor U1239 (N_1239,In_2312,In_2034);
and U1240 (N_1240,In_235,In_91);
and U1241 (N_1241,In_1056,In_2443);
nand U1242 (N_1242,In_2269,In_2061);
or U1243 (N_1243,In_2480,In_695);
nor U1244 (N_1244,In_1909,In_1356);
xor U1245 (N_1245,In_58,In_497);
nor U1246 (N_1246,In_536,In_546);
nor U1247 (N_1247,In_1740,In_2908);
nand U1248 (N_1248,In_297,In_2951);
and U1249 (N_1249,In_670,In_2044);
xor U1250 (N_1250,In_1170,In_542);
and U1251 (N_1251,In_2714,In_1973);
nor U1252 (N_1252,In_30,In_186);
nor U1253 (N_1253,In_377,In_2649);
and U1254 (N_1254,In_122,In_576);
and U1255 (N_1255,In_2807,In_121);
nand U1256 (N_1256,In_1936,In_40);
nand U1257 (N_1257,In_1627,In_1949);
and U1258 (N_1258,In_2006,In_2716);
xor U1259 (N_1259,In_1877,In_1867);
nor U1260 (N_1260,In_2945,In_2134);
nand U1261 (N_1261,In_472,In_1722);
or U1262 (N_1262,In_647,In_2859);
and U1263 (N_1263,In_1661,In_1994);
nand U1264 (N_1264,In_958,In_2166);
nand U1265 (N_1265,In_1519,In_1806);
nor U1266 (N_1266,In_924,In_1135);
or U1267 (N_1267,In_385,In_79);
nand U1268 (N_1268,In_1491,In_1315);
and U1269 (N_1269,In_1679,In_2756);
and U1270 (N_1270,In_11,In_666);
and U1271 (N_1271,In_548,In_636);
or U1272 (N_1272,In_817,In_202);
or U1273 (N_1273,In_894,In_2751);
or U1274 (N_1274,In_2040,In_2327);
nand U1275 (N_1275,In_518,In_2299);
or U1276 (N_1276,In_1795,In_2571);
nand U1277 (N_1277,In_2534,In_2851);
nor U1278 (N_1278,In_1355,In_2519);
nor U1279 (N_1279,In_1857,In_1177);
nand U1280 (N_1280,In_637,In_1691);
xor U1281 (N_1281,In_1833,In_2153);
or U1282 (N_1282,In_1254,In_892);
nand U1283 (N_1283,In_2653,In_962);
and U1284 (N_1284,In_323,In_605);
and U1285 (N_1285,In_2105,In_681);
nor U1286 (N_1286,In_1904,In_2433);
or U1287 (N_1287,In_2160,In_1375);
and U1288 (N_1288,In_2185,In_568);
nor U1289 (N_1289,In_2833,In_1471);
nand U1290 (N_1290,In_1106,In_1545);
nand U1291 (N_1291,In_1848,In_458);
xor U1292 (N_1292,In_19,In_2843);
or U1293 (N_1293,In_422,In_1887);
nor U1294 (N_1294,In_236,In_1791);
nand U1295 (N_1295,In_1807,In_2566);
and U1296 (N_1296,In_2114,In_899);
xnor U1297 (N_1297,In_374,In_833);
or U1298 (N_1298,In_2826,In_2428);
xnor U1299 (N_1299,In_1328,In_1147);
and U1300 (N_1300,In_1400,In_2927);
and U1301 (N_1301,In_291,In_1516);
nand U1302 (N_1302,In_674,In_1637);
nor U1303 (N_1303,In_722,In_88);
nor U1304 (N_1304,In_2561,In_1421);
or U1305 (N_1305,In_2607,In_94);
and U1306 (N_1306,In_2902,In_753);
and U1307 (N_1307,In_2385,In_414);
or U1308 (N_1308,In_2776,In_1946);
or U1309 (N_1309,In_2437,In_2421);
nand U1310 (N_1310,In_2368,In_1446);
and U1311 (N_1311,In_2703,In_1161);
nand U1312 (N_1312,In_2969,In_229);
xnor U1313 (N_1313,In_1011,In_379);
nand U1314 (N_1314,In_2469,In_2041);
nor U1315 (N_1315,In_2938,In_314);
xnor U1316 (N_1316,In_376,In_1256);
nand U1317 (N_1317,In_1817,In_587);
xor U1318 (N_1318,In_889,In_2396);
or U1319 (N_1319,In_459,In_462);
and U1320 (N_1320,In_2540,In_2391);
nand U1321 (N_1321,In_1971,In_931);
xor U1322 (N_1322,In_1612,In_1834);
or U1323 (N_1323,In_511,In_2137);
nor U1324 (N_1324,In_249,In_2132);
or U1325 (N_1325,In_2387,In_1222);
and U1326 (N_1326,In_174,In_1075);
xor U1327 (N_1327,In_1950,In_1792);
nor U1328 (N_1328,In_553,In_909);
nand U1329 (N_1329,In_1987,In_1607);
and U1330 (N_1330,In_309,In_1038);
and U1331 (N_1331,In_847,In_2012);
nor U1332 (N_1332,In_2407,In_1093);
nor U1333 (N_1333,In_994,In_1221);
or U1334 (N_1334,In_1489,In_2616);
nand U1335 (N_1335,In_1654,In_933);
xor U1336 (N_1336,In_2782,In_906);
nand U1337 (N_1337,In_1232,In_1207);
xnor U1338 (N_1338,In_428,In_655);
or U1339 (N_1339,In_1072,In_2003);
and U1340 (N_1340,In_2588,In_2416);
xor U1341 (N_1341,In_1816,In_2971);
xnor U1342 (N_1342,In_2911,In_1339);
xnor U1343 (N_1343,In_421,In_2615);
xnor U1344 (N_1344,In_2533,In_2783);
nor U1345 (N_1345,In_2060,In_653);
xor U1346 (N_1346,In_1780,In_2093);
nand U1347 (N_1347,In_2419,In_2590);
nor U1348 (N_1348,In_645,In_2187);
xor U1349 (N_1349,In_822,In_2228);
xnor U1350 (N_1350,In_133,In_1502);
nor U1351 (N_1351,In_2272,In_709);
xnor U1352 (N_1352,In_689,In_698);
and U1353 (N_1353,In_356,In_880);
and U1354 (N_1354,In_1846,In_1527);
xor U1355 (N_1355,In_1766,In_5);
or U1356 (N_1356,In_2943,In_1214);
xor U1357 (N_1357,In_783,In_2760);
xnor U1358 (N_1358,In_261,In_1535);
nand U1359 (N_1359,In_2818,In_683);
and U1360 (N_1360,In_628,In_781);
nand U1361 (N_1361,In_2221,In_2517);
nand U1362 (N_1362,In_102,In_2713);
xor U1363 (N_1363,In_1783,In_1322);
and U1364 (N_1364,In_483,In_2829);
and U1365 (N_1365,In_72,In_1472);
and U1366 (N_1366,In_210,In_995);
or U1367 (N_1367,In_2095,In_164);
xor U1368 (N_1368,In_2821,In_2087);
and U1369 (N_1369,In_2223,In_1789);
nand U1370 (N_1370,In_136,In_25);
nor U1371 (N_1371,In_2680,In_993);
and U1372 (N_1372,In_1386,In_2083);
and U1373 (N_1373,In_407,In_726);
nand U1374 (N_1374,In_1157,In_842);
xnor U1375 (N_1375,In_2082,In_1870);
nor U1376 (N_1376,In_390,In_1187);
nand U1377 (N_1377,In_987,In_335);
nand U1378 (N_1378,In_2631,In_1525);
and U1379 (N_1379,In_2449,In_2515);
and U1380 (N_1380,In_556,In_2414);
nor U1381 (N_1381,In_2863,In_1454);
nand U1382 (N_1382,In_1708,In_429);
and U1383 (N_1383,In_519,In_184);
or U1384 (N_1384,In_1748,In_2791);
nor U1385 (N_1385,In_2182,In_204);
nand U1386 (N_1386,In_2779,In_1560);
xor U1387 (N_1387,In_2789,In_319);
xor U1388 (N_1388,In_2853,In_965);
nor U1389 (N_1389,In_2499,In_2239);
nor U1390 (N_1390,In_2759,In_1265);
nor U1391 (N_1391,In_103,In_1990);
nand U1392 (N_1392,In_2161,In_95);
and U1393 (N_1393,In_2944,In_1145);
nor U1394 (N_1394,In_1210,In_1830);
nor U1395 (N_1395,In_1018,In_2660);
nand U1396 (N_1396,In_2256,In_1122);
xnor U1397 (N_1397,In_1784,In_2367);
nand U1398 (N_1398,In_2415,In_2042);
nand U1399 (N_1399,In_1081,In_2558);
nor U1400 (N_1400,In_207,In_78);
nor U1401 (N_1401,In_258,In_162);
xor U1402 (N_1402,In_411,In_2698);
xnor U1403 (N_1403,In_954,In_1275);
and U1404 (N_1404,In_625,In_2606);
xor U1405 (N_1405,In_739,In_2988);
nand U1406 (N_1406,In_2627,In_1044);
or U1407 (N_1407,In_2603,In_1988);
or U1408 (N_1408,In_2121,In_2486);
nand U1409 (N_1409,In_1204,In_2143);
xnor U1410 (N_1410,In_2321,In_1067);
or U1411 (N_1411,In_182,In_1013);
or U1412 (N_1412,In_2976,In_1643);
nand U1413 (N_1413,In_936,In_929);
nor U1414 (N_1414,In_1193,In_1486);
or U1415 (N_1415,In_1455,In_1143);
nor U1416 (N_1416,In_2997,In_2858);
or U1417 (N_1417,In_2340,In_2300);
nand U1418 (N_1418,In_2632,In_1696);
nand U1419 (N_1419,In_643,In_2057);
or U1420 (N_1420,In_2320,In_1291);
and U1421 (N_1421,In_2222,In_1493);
nand U1422 (N_1422,In_2018,In_1774);
xnor U1423 (N_1423,In_359,In_1150);
xor U1424 (N_1424,In_1260,In_2602);
or U1425 (N_1425,In_2940,In_1825);
nor U1426 (N_1426,In_2883,In_2207);
nand U1427 (N_1427,In_919,In_1656);
xor U1428 (N_1428,In_592,In_396);
or U1429 (N_1429,In_2009,In_1568);
nor U1430 (N_1430,In_70,In_2772);
nand U1431 (N_1431,In_2048,In_2917);
and U1432 (N_1432,In_1873,In_1363);
and U1433 (N_1433,In_673,In_2871);
nor U1434 (N_1434,In_1947,In_2767);
and U1435 (N_1435,In_2909,In_90);
or U1436 (N_1436,In_1659,In_644);
xnor U1437 (N_1437,In_2462,In_2972);
nand U1438 (N_1438,In_1061,In_1385);
and U1439 (N_1439,In_2339,In_2204);
and U1440 (N_1440,In_1805,In_963);
nand U1441 (N_1441,In_2446,In_2762);
nand U1442 (N_1442,In_1715,In_2170);
xnor U1443 (N_1443,In_2033,In_1695);
or U1444 (N_1444,In_2374,In_2891);
nor U1445 (N_1445,In_1415,In_490);
xnor U1446 (N_1446,In_2314,In_2422);
xnor U1447 (N_1447,In_1965,In_1582);
or U1448 (N_1448,In_596,In_1251);
and U1449 (N_1449,In_911,In_1575);
or U1450 (N_1450,In_1344,In_368);
or U1451 (N_1451,In_299,In_36);
nor U1452 (N_1452,In_1630,In_1610);
nor U1453 (N_1453,In_699,In_1925);
nand U1454 (N_1454,In_2521,In_1274);
nor U1455 (N_1455,In_1124,In_1370);
nand U1456 (N_1456,In_34,In_305);
or U1457 (N_1457,In_222,In_1330);
nor U1458 (N_1458,In_1301,In_841);
xnor U1459 (N_1459,In_471,In_1673);
nand U1460 (N_1460,In_1248,In_2128);
nor U1461 (N_1461,In_610,In_2551);
and U1462 (N_1462,In_278,In_498);
or U1463 (N_1463,In_436,In_1788);
or U1464 (N_1464,In_387,In_731);
and U1465 (N_1465,In_575,In_2889);
or U1466 (N_1466,In_239,In_108);
nand U1467 (N_1467,In_1558,In_866);
or U1468 (N_1468,In_2617,In_2026);
or U1469 (N_1469,In_380,In_1647);
and U1470 (N_1470,In_1523,In_2722);
or U1471 (N_1471,In_1618,In_1635);
nand U1472 (N_1472,In_682,In_2398);
and U1473 (N_1473,In_2011,In_1211);
nand U1474 (N_1474,In_1574,In_484);
nor U1475 (N_1475,In_1974,In_2021);
nor U1476 (N_1476,In_280,In_1646);
nand U1477 (N_1477,In_2238,In_2585);
and U1478 (N_1478,In_2353,In_2064);
and U1479 (N_1479,In_1424,In_2820);
nand U1480 (N_1480,In_1686,In_662);
or U1481 (N_1481,In_1133,In_1350);
nor U1482 (N_1482,In_2130,In_1970);
xor U1483 (N_1483,In_1699,In_1138);
and U1484 (N_1484,In_98,In_1402);
and U1485 (N_1485,In_135,In_1573);
or U1486 (N_1486,In_1465,In_203);
or U1487 (N_1487,In_448,In_2957);
or U1488 (N_1488,In_2800,In_1979);
xnor U1489 (N_1489,In_1382,In_2227);
and U1490 (N_1490,In_971,In_2059);
nor U1491 (N_1491,In_2332,In_2621);
nand U1492 (N_1492,In_2014,In_1642);
and U1493 (N_1493,In_827,In_914);
or U1494 (N_1494,In_660,In_509);
xor U1495 (N_1495,In_612,In_2297);
xor U1496 (N_1496,In_1997,In_2530);
or U1497 (N_1497,In_320,In_2675);
nor U1498 (N_1498,In_2567,In_2906);
and U1499 (N_1499,In_230,In_2640);
nor U1500 (N_1500,In_2602,In_1666);
xnor U1501 (N_1501,In_467,In_1461);
or U1502 (N_1502,In_1555,In_2039);
xor U1503 (N_1503,In_2354,In_2143);
and U1504 (N_1504,In_1721,In_2372);
nor U1505 (N_1505,In_1778,In_851);
and U1506 (N_1506,In_1841,In_1313);
nor U1507 (N_1507,In_1664,In_325);
nor U1508 (N_1508,In_1911,In_568);
or U1509 (N_1509,In_1332,In_1622);
and U1510 (N_1510,In_2259,In_2880);
nand U1511 (N_1511,In_1872,In_1127);
or U1512 (N_1512,In_1619,In_1734);
and U1513 (N_1513,In_2925,In_158);
nand U1514 (N_1514,In_765,In_581);
xor U1515 (N_1515,In_1104,In_302);
and U1516 (N_1516,In_1249,In_2303);
xnor U1517 (N_1517,In_1075,In_239);
or U1518 (N_1518,In_2723,In_581);
xor U1519 (N_1519,In_2258,In_1026);
or U1520 (N_1520,In_2961,In_2591);
and U1521 (N_1521,In_1700,In_1801);
xor U1522 (N_1522,In_1140,In_2642);
and U1523 (N_1523,In_2189,In_956);
or U1524 (N_1524,In_629,In_1990);
nor U1525 (N_1525,In_429,In_2201);
xor U1526 (N_1526,In_2139,In_1346);
nor U1527 (N_1527,In_103,In_2791);
or U1528 (N_1528,In_1904,In_2196);
nor U1529 (N_1529,In_627,In_268);
and U1530 (N_1530,In_2746,In_2629);
nor U1531 (N_1531,In_886,In_1532);
or U1532 (N_1532,In_771,In_1879);
nor U1533 (N_1533,In_601,In_344);
or U1534 (N_1534,In_1924,In_2614);
and U1535 (N_1535,In_2378,In_2912);
or U1536 (N_1536,In_1371,In_355);
xnor U1537 (N_1537,In_1849,In_2255);
nor U1538 (N_1538,In_252,In_453);
nor U1539 (N_1539,In_1651,In_1451);
and U1540 (N_1540,In_2682,In_2427);
xnor U1541 (N_1541,In_1778,In_749);
or U1542 (N_1542,In_2617,In_1255);
or U1543 (N_1543,In_2564,In_432);
nor U1544 (N_1544,In_2587,In_1404);
and U1545 (N_1545,In_861,In_977);
nor U1546 (N_1546,In_466,In_376);
and U1547 (N_1547,In_1230,In_291);
nor U1548 (N_1548,In_405,In_326);
nor U1549 (N_1549,In_1027,In_2829);
nand U1550 (N_1550,In_2657,In_2487);
or U1551 (N_1551,In_874,In_2486);
nor U1552 (N_1552,In_2285,In_2986);
and U1553 (N_1553,In_1395,In_333);
and U1554 (N_1554,In_1748,In_2330);
and U1555 (N_1555,In_1002,In_1674);
or U1556 (N_1556,In_589,In_1329);
nor U1557 (N_1557,In_2772,In_47);
nor U1558 (N_1558,In_719,In_53);
nand U1559 (N_1559,In_1490,In_1240);
nand U1560 (N_1560,In_604,In_407);
and U1561 (N_1561,In_2523,In_1762);
nand U1562 (N_1562,In_2051,In_2067);
nand U1563 (N_1563,In_797,In_574);
or U1564 (N_1564,In_480,In_1233);
nor U1565 (N_1565,In_171,In_2146);
nand U1566 (N_1566,In_654,In_2819);
nor U1567 (N_1567,In_123,In_507);
and U1568 (N_1568,In_1753,In_2058);
and U1569 (N_1569,In_1902,In_2079);
nand U1570 (N_1570,In_2537,In_1063);
and U1571 (N_1571,In_1382,In_1567);
nand U1572 (N_1572,In_920,In_130);
and U1573 (N_1573,In_2300,In_1246);
nand U1574 (N_1574,In_116,In_2983);
or U1575 (N_1575,In_415,In_2602);
nand U1576 (N_1576,In_1033,In_2052);
nand U1577 (N_1577,In_822,In_1319);
nand U1578 (N_1578,In_2905,In_201);
nand U1579 (N_1579,In_197,In_2201);
or U1580 (N_1580,In_766,In_383);
xor U1581 (N_1581,In_1939,In_1937);
nand U1582 (N_1582,In_1706,In_362);
nand U1583 (N_1583,In_1290,In_57);
nand U1584 (N_1584,In_1255,In_746);
nand U1585 (N_1585,In_1548,In_2519);
and U1586 (N_1586,In_1712,In_1476);
xor U1587 (N_1587,In_383,In_225);
or U1588 (N_1588,In_2191,In_259);
or U1589 (N_1589,In_1275,In_2596);
nor U1590 (N_1590,In_2189,In_119);
xnor U1591 (N_1591,In_2821,In_440);
or U1592 (N_1592,In_2085,In_1989);
nor U1593 (N_1593,In_2396,In_1397);
or U1594 (N_1594,In_486,In_2668);
nor U1595 (N_1595,In_1326,In_2936);
or U1596 (N_1596,In_461,In_868);
and U1597 (N_1597,In_2593,In_1099);
xor U1598 (N_1598,In_2592,In_328);
nand U1599 (N_1599,In_2676,In_1210);
or U1600 (N_1600,In_1519,In_401);
and U1601 (N_1601,In_1603,In_140);
xnor U1602 (N_1602,In_964,In_958);
nor U1603 (N_1603,In_1034,In_436);
or U1604 (N_1604,In_1944,In_860);
nand U1605 (N_1605,In_445,In_5);
xnor U1606 (N_1606,In_6,In_2488);
or U1607 (N_1607,In_669,In_2702);
nor U1608 (N_1608,In_2052,In_2825);
xnor U1609 (N_1609,In_1546,In_1027);
or U1610 (N_1610,In_570,In_2886);
xnor U1611 (N_1611,In_2065,In_1690);
xnor U1612 (N_1612,In_2355,In_22);
nor U1613 (N_1613,In_5,In_2707);
xor U1614 (N_1614,In_30,In_1674);
or U1615 (N_1615,In_1878,In_2234);
nor U1616 (N_1616,In_2388,In_2610);
xnor U1617 (N_1617,In_74,In_1208);
and U1618 (N_1618,In_647,In_1251);
and U1619 (N_1619,In_1315,In_1803);
nor U1620 (N_1620,In_661,In_1256);
xnor U1621 (N_1621,In_2418,In_2558);
nand U1622 (N_1622,In_877,In_1725);
and U1623 (N_1623,In_1924,In_522);
and U1624 (N_1624,In_2575,In_659);
xor U1625 (N_1625,In_1992,In_882);
and U1626 (N_1626,In_2301,In_1408);
or U1627 (N_1627,In_1801,In_2546);
nand U1628 (N_1628,In_420,In_186);
or U1629 (N_1629,In_1275,In_1891);
nand U1630 (N_1630,In_1566,In_1054);
and U1631 (N_1631,In_1535,In_2004);
and U1632 (N_1632,In_1819,In_1067);
or U1633 (N_1633,In_902,In_2171);
nand U1634 (N_1634,In_2574,In_2470);
and U1635 (N_1635,In_2233,In_396);
nor U1636 (N_1636,In_1042,In_1255);
xor U1637 (N_1637,In_1726,In_2897);
nor U1638 (N_1638,In_2993,In_480);
nand U1639 (N_1639,In_1530,In_2712);
nor U1640 (N_1640,In_2126,In_1735);
and U1641 (N_1641,In_2239,In_343);
and U1642 (N_1642,In_2373,In_1287);
and U1643 (N_1643,In_1141,In_2100);
nand U1644 (N_1644,In_2421,In_2831);
xnor U1645 (N_1645,In_2948,In_2239);
xnor U1646 (N_1646,In_608,In_1663);
nor U1647 (N_1647,In_2149,In_1378);
xnor U1648 (N_1648,In_2971,In_410);
nand U1649 (N_1649,In_1669,In_1404);
xor U1650 (N_1650,In_534,In_1180);
nand U1651 (N_1651,In_2328,In_999);
nand U1652 (N_1652,In_1706,In_2702);
nor U1653 (N_1653,In_280,In_511);
or U1654 (N_1654,In_652,In_1057);
nand U1655 (N_1655,In_280,In_2199);
nor U1656 (N_1656,In_1482,In_1650);
or U1657 (N_1657,In_1624,In_224);
or U1658 (N_1658,In_786,In_2432);
and U1659 (N_1659,In_328,In_599);
or U1660 (N_1660,In_568,In_2639);
and U1661 (N_1661,In_1656,In_877);
or U1662 (N_1662,In_2267,In_1046);
xnor U1663 (N_1663,In_125,In_926);
xnor U1664 (N_1664,In_661,In_1902);
or U1665 (N_1665,In_923,In_2516);
or U1666 (N_1666,In_1197,In_170);
and U1667 (N_1667,In_2061,In_317);
nor U1668 (N_1668,In_1637,In_2216);
or U1669 (N_1669,In_128,In_1822);
and U1670 (N_1670,In_1331,In_135);
or U1671 (N_1671,In_1002,In_191);
xnor U1672 (N_1672,In_359,In_978);
nand U1673 (N_1673,In_2447,In_1470);
xor U1674 (N_1674,In_1706,In_1283);
nand U1675 (N_1675,In_2051,In_26);
nand U1676 (N_1676,In_1051,In_1526);
nor U1677 (N_1677,In_1412,In_896);
nand U1678 (N_1678,In_1614,In_116);
nor U1679 (N_1679,In_1448,In_509);
nand U1680 (N_1680,In_347,In_411);
xor U1681 (N_1681,In_2442,In_1044);
or U1682 (N_1682,In_563,In_2416);
xor U1683 (N_1683,In_1451,In_2695);
or U1684 (N_1684,In_998,In_670);
or U1685 (N_1685,In_532,In_2999);
and U1686 (N_1686,In_487,In_2185);
nor U1687 (N_1687,In_2691,In_2104);
or U1688 (N_1688,In_437,In_431);
nor U1689 (N_1689,In_1593,In_2944);
nor U1690 (N_1690,In_1405,In_494);
nand U1691 (N_1691,In_1952,In_1109);
or U1692 (N_1692,In_1964,In_733);
nor U1693 (N_1693,In_2575,In_2462);
or U1694 (N_1694,In_220,In_530);
xnor U1695 (N_1695,In_1269,In_387);
nor U1696 (N_1696,In_1571,In_1192);
nand U1697 (N_1697,In_1368,In_2792);
xor U1698 (N_1698,In_2612,In_61);
nor U1699 (N_1699,In_807,In_1741);
and U1700 (N_1700,In_1286,In_5);
or U1701 (N_1701,In_2556,In_1717);
nor U1702 (N_1702,In_191,In_1914);
xnor U1703 (N_1703,In_623,In_2765);
and U1704 (N_1704,In_2033,In_2411);
or U1705 (N_1705,In_537,In_2581);
and U1706 (N_1706,In_386,In_2657);
nand U1707 (N_1707,In_1291,In_2581);
or U1708 (N_1708,In_1302,In_1381);
nand U1709 (N_1709,In_2048,In_1191);
nand U1710 (N_1710,In_2821,In_390);
or U1711 (N_1711,In_1621,In_1513);
nand U1712 (N_1712,In_2366,In_1605);
xor U1713 (N_1713,In_2070,In_1170);
nor U1714 (N_1714,In_154,In_1258);
or U1715 (N_1715,In_2866,In_27);
xor U1716 (N_1716,In_1550,In_335);
nand U1717 (N_1717,In_2638,In_1533);
nand U1718 (N_1718,In_2459,In_313);
or U1719 (N_1719,In_2317,In_556);
xnor U1720 (N_1720,In_361,In_2759);
nor U1721 (N_1721,In_508,In_367);
nor U1722 (N_1722,In_2764,In_1863);
nand U1723 (N_1723,In_476,In_2530);
nand U1724 (N_1724,In_2418,In_1302);
nor U1725 (N_1725,In_1211,In_608);
nor U1726 (N_1726,In_2365,In_664);
nor U1727 (N_1727,In_2871,In_1071);
xnor U1728 (N_1728,In_1423,In_877);
nand U1729 (N_1729,In_1718,In_1312);
xor U1730 (N_1730,In_219,In_2896);
nand U1731 (N_1731,In_787,In_805);
nand U1732 (N_1732,In_1348,In_2915);
xnor U1733 (N_1733,In_2807,In_1663);
nor U1734 (N_1734,In_2554,In_1445);
xor U1735 (N_1735,In_206,In_570);
nand U1736 (N_1736,In_2075,In_1861);
or U1737 (N_1737,In_779,In_997);
or U1738 (N_1738,In_845,In_2745);
xnor U1739 (N_1739,In_1256,In_457);
xor U1740 (N_1740,In_2608,In_2777);
nor U1741 (N_1741,In_1685,In_131);
xor U1742 (N_1742,In_2449,In_228);
or U1743 (N_1743,In_1347,In_2971);
xor U1744 (N_1744,In_258,In_233);
and U1745 (N_1745,In_2641,In_467);
and U1746 (N_1746,In_451,In_1933);
xnor U1747 (N_1747,In_1929,In_2659);
nor U1748 (N_1748,In_1905,In_2653);
xor U1749 (N_1749,In_1304,In_2049);
nor U1750 (N_1750,In_2902,In_474);
nor U1751 (N_1751,In_2527,In_826);
nor U1752 (N_1752,In_918,In_208);
and U1753 (N_1753,In_1328,In_1790);
or U1754 (N_1754,In_849,In_2981);
nor U1755 (N_1755,In_544,In_2035);
xor U1756 (N_1756,In_803,In_674);
nand U1757 (N_1757,In_543,In_449);
and U1758 (N_1758,In_2252,In_684);
nand U1759 (N_1759,In_2448,In_2837);
or U1760 (N_1760,In_2688,In_2334);
xor U1761 (N_1761,In_2396,In_210);
nor U1762 (N_1762,In_567,In_1228);
xor U1763 (N_1763,In_324,In_2852);
and U1764 (N_1764,In_2450,In_2202);
nor U1765 (N_1765,In_664,In_1950);
xor U1766 (N_1766,In_1187,In_1048);
and U1767 (N_1767,In_306,In_2936);
or U1768 (N_1768,In_1224,In_1585);
nand U1769 (N_1769,In_530,In_1930);
xnor U1770 (N_1770,In_1564,In_1184);
xnor U1771 (N_1771,In_248,In_2003);
and U1772 (N_1772,In_901,In_2000);
nand U1773 (N_1773,In_1808,In_1771);
and U1774 (N_1774,In_820,In_21);
nor U1775 (N_1775,In_1900,In_2213);
or U1776 (N_1776,In_1492,In_2884);
or U1777 (N_1777,In_2362,In_878);
xor U1778 (N_1778,In_2621,In_1911);
xor U1779 (N_1779,In_854,In_2488);
or U1780 (N_1780,In_1333,In_1051);
or U1781 (N_1781,In_2227,In_2323);
nor U1782 (N_1782,In_1800,In_452);
nand U1783 (N_1783,In_29,In_2804);
nand U1784 (N_1784,In_1270,In_229);
nand U1785 (N_1785,In_1007,In_16);
nand U1786 (N_1786,In_2484,In_2390);
and U1787 (N_1787,In_359,In_1641);
nand U1788 (N_1788,In_1374,In_2982);
xor U1789 (N_1789,In_849,In_736);
xor U1790 (N_1790,In_2940,In_1613);
nand U1791 (N_1791,In_246,In_247);
or U1792 (N_1792,In_953,In_2339);
nor U1793 (N_1793,In_1682,In_398);
and U1794 (N_1794,In_2171,In_1917);
or U1795 (N_1795,In_426,In_2893);
and U1796 (N_1796,In_1704,In_698);
nor U1797 (N_1797,In_369,In_1589);
or U1798 (N_1798,In_1466,In_1727);
or U1799 (N_1799,In_521,In_1827);
xor U1800 (N_1800,In_2487,In_2430);
or U1801 (N_1801,In_1960,In_566);
nand U1802 (N_1802,In_1438,In_1382);
xor U1803 (N_1803,In_2217,In_771);
xnor U1804 (N_1804,In_2801,In_433);
nand U1805 (N_1805,In_822,In_1115);
nor U1806 (N_1806,In_777,In_2659);
nor U1807 (N_1807,In_345,In_1714);
nor U1808 (N_1808,In_583,In_1809);
or U1809 (N_1809,In_1611,In_700);
nor U1810 (N_1810,In_95,In_2121);
nor U1811 (N_1811,In_1459,In_2203);
nand U1812 (N_1812,In_993,In_2013);
or U1813 (N_1813,In_823,In_1380);
and U1814 (N_1814,In_1249,In_438);
xor U1815 (N_1815,In_62,In_1799);
xor U1816 (N_1816,In_1965,In_2389);
and U1817 (N_1817,In_611,In_1117);
nor U1818 (N_1818,In_1576,In_1961);
or U1819 (N_1819,In_706,In_261);
and U1820 (N_1820,In_1466,In_487);
nand U1821 (N_1821,In_2126,In_645);
nand U1822 (N_1822,In_117,In_2135);
xor U1823 (N_1823,In_2534,In_1764);
xnor U1824 (N_1824,In_961,In_1970);
or U1825 (N_1825,In_1239,In_1125);
xor U1826 (N_1826,In_1740,In_2150);
or U1827 (N_1827,In_1436,In_2634);
nand U1828 (N_1828,In_1037,In_1032);
xor U1829 (N_1829,In_1694,In_69);
or U1830 (N_1830,In_493,In_689);
and U1831 (N_1831,In_662,In_268);
or U1832 (N_1832,In_63,In_278);
xor U1833 (N_1833,In_1400,In_1753);
xor U1834 (N_1834,In_2060,In_1411);
nor U1835 (N_1835,In_304,In_1293);
nor U1836 (N_1836,In_2366,In_1351);
or U1837 (N_1837,In_557,In_2171);
nor U1838 (N_1838,In_2093,In_1501);
nor U1839 (N_1839,In_2972,In_303);
nand U1840 (N_1840,In_2235,In_1176);
xor U1841 (N_1841,In_1632,In_1477);
xor U1842 (N_1842,In_2928,In_320);
nand U1843 (N_1843,In_1287,In_2757);
or U1844 (N_1844,In_1337,In_36);
nand U1845 (N_1845,In_2823,In_2044);
nor U1846 (N_1846,In_446,In_801);
and U1847 (N_1847,In_2370,In_232);
or U1848 (N_1848,In_750,In_1702);
or U1849 (N_1849,In_182,In_979);
and U1850 (N_1850,In_70,In_227);
and U1851 (N_1851,In_1194,In_341);
xor U1852 (N_1852,In_1435,In_818);
or U1853 (N_1853,In_997,In_395);
and U1854 (N_1854,In_1381,In_2524);
nand U1855 (N_1855,In_2706,In_463);
xor U1856 (N_1856,In_430,In_180);
xnor U1857 (N_1857,In_2808,In_1351);
and U1858 (N_1858,In_2290,In_2785);
nor U1859 (N_1859,In_2688,In_1693);
nor U1860 (N_1860,In_2676,In_2929);
nand U1861 (N_1861,In_1410,In_2191);
xor U1862 (N_1862,In_1215,In_2594);
or U1863 (N_1863,In_2716,In_824);
and U1864 (N_1864,In_1294,In_2870);
and U1865 (N_1865,In_1855,In_1446);
nor U1866 (N_1866,In_2768,In_1210);
or U1867 (N_1867,In_815,In_2654);
nor U1868 (N_1868,In_2581,In_1753);
nor U1869 (N_1869,In_125,In_2259);
and U1870 (N_1870,In_1570,In_2386);
and U1871 (N_1871,In_844,In_1175);
nand U1872 (N_1872,In_315,In_1578);
nor U1873 (N_1873,In_1645,In_1175);
and U1874 (N_1874,In_108,In_2850);
nand U1875 (N_1875,In_1081,In_11);
nor U1876 (N_1876,In_898,In_276);
nand U1877 (N_1877,In_1334,In_1140);
or U1878 (N_1878,In_293,In_2633);
nor U1879 (N_1879,In_1657,In_1060);
xnor U1880 (N_1880,In_622,In_927);
nor U1881 (N_1881,In_1989,In_1204);
xor U1882 (N_1882,In_2136,In_1021);
nor U1883 (N_1883,In_2576,In_2874);
nor U1884 (N_1884,In_664,In_2030);
or U1885 (N_1885,In_2783,In_1451);
nand U1886 (N_1886,In_2342,In_230);
xor U1887 (N_1887,In_708,In_513);
and U1888 (N_1888,In_2278,In_2189);
nand U1889 (N_1889,In_668,In_976);
xor U1890 (N_1890,In_2564,In_1564);
nor U1891 (N_1891,In_1088,In_108);
xor U1892 (N_1892,In_1516,In_1150);
nand U1893 (N_1893,In_1348,In_759);
xor U1894 (N_1894,In_1470,In_2814);
or U1895 (N_1895,In_804,In_1183);
or U1896 (N_1896,In_696,In_2397);
xor U1897 (N_1897,In_1675,In_1912);
and U1898 (N_1898,In_1275,In_2820);
nand U1899 (N_1899,In_1070,In_357);
nor U1900 (N_1900,In_314,In_1749);
or U1901 (N_1901,In_2353,In_2866);
or U1902 (N_1902,In_2049,In_2153);
nor U1903 (N_1903,In_320,In_283);
nand U1904 (N_1904,In_263,In_199);
nor U1905 (N_1905,In_1565,In_303);
and U1906 (N_1906,In_2248,In_2300);
and U1907 (N_1907,In_392,In_49);
xnor U1908 (N_1908,In_1435,In_2055);
and U1909 (N_1909,In_2506,In_534);
nand U1910 (N_1910,In_987,In_2026);
nor U1911 (N_1911,In_714,In_2595);
and U1912 (N_1912,In_1053,In_2256);
nand U1913 (N_1913,In_1676,In_1702);
or U1914 (N_1914,In_1971,In_2497);
nand U1915 (N_1915,In_905,In_761);
nand U1916 (N_1916,In_432,In_977);
and U1917 (N_1917,In_1618,In_95);
or U1918 (N_1918,In_2692,In_522);
or U1919 (N_1919,In_416,In_137);
xnor U1920 (N_1920,In_842,In_1141);
xnor U1921 (N_1921,In_2554,In_1972);
xor U1922 (N_1922,In_624,In_13);
xnor U1923 (N_1923,In_2312,In_1248);
and U1924 (N_1924,In_1024,In_1556);
and U1925 (N_1925,In_2091,In_897);
or U1926 (N_1926,In_792,In_821);
or U1927 (N_1927,In_2781,In_562);
nand U1928 (N_1928,In_2244,In_615);
and U1929 (N_1929,In_833,In_1285);
or U1930 (N_1930,In_1228,In_112);
and U1931 (N_1931,In_1625,In_1748);
and U1932 (N_1932,In_897,In_2251);
or U1933 (N_1933,In_1327,In_65);
nand U1934 (N_1934,In_2987,In_34);
xnor U1935 (N_1935,In_2064,In_114);
and U1936 (N_1936,In_2724,In_506);
nor U1937 (N_1937,In_1886,In_317);
nand U1938 (N_1938,In_1673,In_2074);
and U1939 (N_1939,In_2386,In_1756);
xor U1940 (N_1940,In_2569,In_2716);
or U1941 (N_1941,In_1185,In_1435);
nand U1942 (N_1942,In_2299,In_2779);
or U1943 (N_1943,In_1877,In_1314);
or U1944 (N_1944,In_1427,In_40);
nor U1945 (N_1945,In_508,In_783);
nand U1946 (N_1946,In_191,In_798);
or U1947 (N_1947,In_1693,In_1516);
xor U1948 (N_1948,In_1202,In_265);
xnor U1949 (N_1949,In_2046,In_1465);
or U1950 (N_1950,In_2032,In_2287);
or U1951 (N_1951,In_2508,In_88);
xnor U1952 (N_1952,In_129,In_2259);
nor U1953 (N_1953,In_1152,In_1306);
and U1954 (N_1954,In_1527,In_1480);
xor U1955 (N_1955,In_808,In_562);
xor U1956 (N_1956,In_453,In_623);
or U1957 (N_1957,In_1333,In_710);
or U1958 (N_1958,In_342,In_2291);
nor U1959 (N_1959,In_380,In_2202);
xnor U1960 (N_1960,In_59,In_1254);
nand U1961 (N_1961,In_561,In_850);
or U1962 (N_1962,In_345,In_2638);
nor U1963 (N_1963,In_2393,In_294);
xnor U1964 (N_1964,In_910,In_950);
nor U1965 (N_1965,In_2791,In_34);
xor U1966 (N_1966,In_325,In_1256);
nand U1967 (N_1967,In_577,In_805);
and U1968 (N_1968,In_2835,In_315);
nor U1969 (N_1969,In_2682,In_2481);
nand U1970 (N_1970,In_2992,In_2158);
and U1971 (N_1971,In_1833,In_2261);
nor U1972 (N_1972,In_572,In_1528);
and U1973 (N_1973,In_779,In_2689);
and U1974 (N_1974,In_2340,In_960);
nor U1975 (N_1975,In_2700,In_639);
nand U1976 (N_1976,In_2201,In_446);
or U1977 (N_1977,In_963,In_2623);
xnor U1978 (N_1978,In_665,In_2972);
and U1979 (N_1979,In_796,In_1960);
xor U1980 (N_1980,In_664,In_956);
xnor U1981 (N_1981,In_372,In_2500);
and U1982 (N_1982,In_2619,In_297);
nor U1983 (N_1983,In_1287,In_2531);
and U1984 (N_1984,In_1431,In_1634);
and U1985 (N_1985,In_1713,In_1585);
xor U1986 (N_1986,In_1737,In_1190);
and U1987 (N_1987,In_2700,In_1979);
nand U1988 (N_1988,In_1098,In_1121);
xor U1989 (N_1989,In_2554,In_2721);
or U1990 (N_1990,In_1611,In_1897);
xnor U1991 (N_1991,In_2611,In_316);
xor U1992 (N_1992,In_2822,In_64);
nor U1993 (N_1993,In_1650,In_2399);
nor U1994 (N_1994,In_2462,In_1365);
xnor U1995 (N_1995,In_2876,In_1215);
xor U1996 (N_1996,In_2936,In_540);
and U1997 (N_1997,In_1769,In_1192);
nor U1998 (N_1998,In_662,In_1);
nand U1999 (N_1999,In_1553,In_1352);
or U2000 (N_2000,N_39,N_1675);
or U2001 (N_2001,N_1739,N_1581);
nand U2002 (N_2002,N_58,N_800);
and U2003 (N_2003,N_311,N_1598);
or U2004 (N_2004,N_1859,N_725);
xnor U2005 (N_2005,N_426,N_615);
nor U2006 (N_2006,N_1555,N_1792);
xor U2007 (N_2007,N_959,N_1536);
xor U2008 (N_2008,N_861,N_1038);
or U2009 (N_2009,N_604,N_1127);
nand U2010 (N_2010,N_666,N_1452);
nand U2011 (N_2011,N_823,N_1152);
or U2012 (N_2012,N_1828,N_1800);
and U2013 (N_2013,N_696,N_808);
nor U2014 (N_2014,N_1296,N_339);
nor U2015 (N_2015,N_1063,N_565);
or U2016 (N_2016,N_299,N_191);
or U2017 (N_2017,N_1669,N_1707);
nor U2018 (N_2018,N_173,N_1387);
xnor U2019 (N_2019,N_967,N_957);
nand U2020 (N_2020,N_297,N_480);
nand U2021 (N_2021,N_810,N_1723);
nand U2022 (N_2022,N_607,N_1637);
nor U2023 (N_2023,N_649,N_64);
and U2024 (N_2024,N_1138,N_356);
nand U2025 (N_2025,N_1733,N_1622);
nand U2026 (N_2026,N_1579,N_1280);
nand U2027 (N_2027,N_1758,N_1606);
or U2028 (N_2028,N_1922,N_933);
or U2029 (N_2029,N_1010,N_1345);
nor U2030 (N_2030,N_1766,N_1070);
nor U2031 (N_2031,N_1718,N_1066);
xnor U2032 (N_2032,N_1664,N_161);
and U2033 (N_2033,N_1678,N_1483);
or U2034 (N_2034,N_1183,N_730);
nor U2035 (N_2035,N_281,N_611);
and U2036 (N_2036,N_205,N_1780);
and U2037 (N_2037,N_1001,N_1174);
or U2038 (N_2038,N_33,N_786);
and U2039 (N_2039,N_1545,N_150);
or U2040 (N_2040,N_37,N_446);
nand U2041 (N_2041,N_714,N_335);
or U2042 (N_2042,N_359,N_1013);
and U2043 (N_2043,N_247,N_134);
xnor U2044 (N_2044,N_306,N_1926);
nor U2045 (N_2045,N_818,N_507);
nand U2046 (N_2046,N_345,N_589);
and U2047 (N_2047,N_1119,N_934);
or U2048 (N_2048,N_427,N_1429);
nand U2049 (N_2049,N_1794,N_49);
and U2050 (N_2050,N_682,N_1176);
nand U2051 (N_2051,N_1500,N_1959);
nand U2052 (N_2052,N_357,N_314);
nand U2053 (N_2053,N_1779,N_1473);
nor U2054 (N_2054,N_1956,N_1488);
nor U2055 (N_2055,N_417,N_464);
nand U2056 (N_2056,N_1254,N_962);
nor U2057 (N_2057,N_1065,N_459);
and U2058 (N_2058,N_1680,N_1411);
and U2059 (N_2059,N_1023,N_1930);
xor U2060 (N_2060,N_224,N_32);
xor U2061 (N_2061,N_470,N_1860);
nor U2062 (N_2062,N_1952,N_1671);
nand U2063 (N_2063,N_997,N_453);
and U2064 (N_2064,N_1507,N_119);
xor U2065 (N_2065,N_530,N_1998);
nand U2066 (N_2066,N_966,N_391);
xnor U2067 (N_2067,N_576,N_544);
nor U2068 (N_2068,N_1289,N_1279);
or U2069 (N_2069,N_746,N_1416);
or U2070 (N_2070,N_1297,N_892);
nand U2071 (N_2071,N_1706,N_1619);
xnor U2072 (N_2072,N_239,N_1761);
and U2073 (N_2073,N_1201,N_286);
and U2074 (N_2074,N_1661,N_31);
or U2075 (N_2075,N_697,N_59);
and U2076 (N_2076,N_77,N_1658);
nor U2077 (N_2077,N_938,N_1951);
and U2078 (N_2078,N_274,N_1463);
xnor U2079 (N_2079,N_1133,N_1027);
and U2080 (N_2080,N_881,N_1564);
nand U2081 (N_2081,N_988,N_1260);
nor U2082 (N_2082,N_656,N_659);
nor U2083 (N_2083,N_1479,N_630);
or U2084 (N_2084,N_768,N_1881);
xnor U2085 (N_2085,N_414,N_1018);
nand U2086 (N_2086,N_1143,N_1550);
nand U2087 (N_2087,N_592,N_1660);
xor U2088 (N_2088,N_1314,N_1367);
nand U2089 (N_2089,N_1921,N_727);
nand U2090 (N_2090,N_1547,N_597);
xor U2091 (N_2091,N_1724,N_371);
or U2092 (N_2092,N_1571,N_321);
or U2093 (N_2093,N_703,N_1182);
nor U2094 (N_2094,N_159,N_1643);
nand U2095 (N_2095,N_474,N_509);
xor U2096 (N_2096,N_1745,N_372);
and U2097 (N_2097,N_1316,N_1394);
and U2098 (N_2098,N_375,N_1272);
xnor U2099 (N_2099,N_575,N_1121);
or U2100 (N_2100,N_147,N_148);
nor U2101 (N_2101,N_140,N_863);
or U2102 (N_2102,N_911,N_1135);
nor U2103 (N_2103,N_925,N_1358);
and U2104 (N_2104,N_226,N_1556);
and U2105 (N_2105,N_403,N_1087);
and U2106 (N_2106,N_1770,N_756);
and U2107 (N_2107,N_1667,N_61);
nor U2108 (N_2108,N_1246,N_586);
or U2109 (N_2109,N_1697,N_1050);
xnor U2110 (N_2110,N_203,N_1113);
nor U2111 (N_2111,N_608,N_1361);
xor U2112 (N_2112,N_495,N_1496);
nand U2113 (N_2113,N_418,N_1047);
xor U2114 (N_2114,N_486,N_1195);
nor U2115 (N_2115,N_1436,N_1576);
nand U2116 (N_2116,N_1041,N_385);
and U2117 (N_2117,N_580,N_1891);
xnor U2118 (N_2118,N_1508,N_904);
or U2119 (N_2119,N_621,N_977);
nand U2120 (N_2120,N_1693,N_1491);
nand U2121 (N_2121,N_767,N_1422);
nand U2122 (N_2122,N_1168,N_388);
nand U2123 (N_2123,N_1222,N_132);
nor U2124 (N_2124,N_1906,N_1625);
nor U2125 (N_2125,N_326,N_496);
xnor U2126 (N_2126,N_1273,N_201);
and U2127 (N_2127,N_112,N_1553);
or U2128 (N_2128,N_781,N_1798);
and U2129 (N_2129,N_1386,N_1595);
nor U2130 (N_2130,N_884,N_1437);
and U2131 (N_2131,N_1392,N_1778);
and U2132 (N_2132,N_1155,N_1799);
nand U2133 (N_2133,N_518,N_1459);
and U2134 (N_2134,N_1224,N_185);
xor U2135 (N_2135,N_587,N_436);
nand U2136 (N_2136,N_1223,N_1966);
and U2137 (N_2137,N_1321,N_614);
xnor U2138 (N_2138,N_1626,N_53);
nand U2139 (N_2139,N_318,N_994);
nand U2140 (N_2140,N_1858,N_916);
nor U2141 (N_2141,N_1325,N_844);
or U2142 (N_2142,N_1151,N_429);
nand U2143 (N_2143,N_1080,N_260);
and U2144 (N_2144,N_1274,N_873);
or U2145 (N_2145,N_413,N_1282);
or U2146 (N_2146,N_794,N_1048);
xnor U2147 (N_2147,N_1957,N_1665);
nand U2148 (N_2148,N_1291,N_1343);
xnor U2149 (N_2149,N_1097,N_277);
nand U2150 (N_2150,N_368,N_1942);
nand U2151 (N_2151,N_489,N_1944);
nor U2152 (N_2152,N_1374,N_747);
and U2153 (N_2153,N_513,N_1600);
and U2154 (N_2154,N_1501,N_1456);
xor U2155 (N_2155,N_13,N_954);
and U2156 (N_2156,N_491,N_141);
and U2157 (N_2157,N_1668,N_519);
or U2158 (N_2158,N_200,N_895);
xor U2159 (N_2159,N_1160,N_1318);
and U2160 (N_2160,N_1397,N_36);
nand U2161 (N_2161,N_840,N_120);
nand U2162 (N_2162,N_729,N_1574);
nand U2163 (N_2163,N_1278,N_1524);
xnor U2164 (N_2164,N_7,N_1029);
xor U2165 (N_2165,N_724,N_1652);
nor U2166 (N_2166,N_1692,N_1315);
nor U2167 (N_2167,N_1356,N_1610);
nand U2168 (N_2168,N_126,N_499);
nand U2169 (N_2169,N_1819,N_710);
nand U2170 (N_2170,N_1431,N_228);
nor U2171 (N_2171,N_1695,N_1457);
nor U2172 (N_2172,N_673,N_1025);
nand U2173 (N_2173,N_1214,N_947);
or U2174 (N_2174,N_868,N_1283);
or U2175 (N_2175,N_1403,N_145);
and U2176 (N_2176,N_1982,N_582);
nand U2177 (N_2177,N_744,N_324);
nor U2178 (N_2178,N_1110,N_914);
or U2179 (N_2179,N_633,N_1599);
nand U2180 (N_2180,N_1931,N_348);
xnor U2181 (N_2181,N_483,N_1578);
and U2182 (N_2182,N_1713,N_590);
and U2183 (N_2183,N_1776,N_1084);
or U2184 (N_2184,N_1051,N_287);
nand U2185 (N_2185,N_1002,N_215);
nor U2186 (N_2186,N_1352,N_733);
nor U2187 (N_2187,N_1977,N_1878);
or U2188 (N_2188,N_1910,N_867);
nor U2189 (N_2189,N_643,N_38);
nand U2190 (N_2190,N_680,N_1519);
nand U2191 (N_2191,N_569,N_1360);
or U2192 (N_2192,N_1469,N_1955);
xor U2193 (N_2193,N_1357,N_660);
nand U2194 (N_2194,N_851,N_1915);
nand U2195 (N_2195,N_931,N_1885);
xor U2196 (N_2196,N_1268,N_1607);
and U2197 (N_2197,N_1364,N_1414);
xor U2198 (N_2198,N_1848,N_1383);
and U2199 (N_2199,N_435,N_748);
nor U2200 (N_2200,N_1552,N_1771);
nor U2201 (N_2201,N_117,N_54);
nand U2202 (N_2202,N_1845,N_1935);
xor U2203 (N_2203,N_785,N_628);
and U2204 (N_2204,N_285,N_476);
nor U2205 (N_2205,N_1221,N_1270);
and U2206 (N_2206,N_1727,N_1980);
or U2207 (N_2207,N_504,N_1188);
nand U2208 (N_2208,N_1109,N_813);
xor U2209 (N_2209,N_635,N_296);
nand U2210 (N_2210,N_1918,N_1755);
xor U2211 (N_2211,N_494,N_1218);
xnor U2212 (N_2212,N_273,N_872);
or U2213 (N_2213,N_960,N_1642);
and U2214 (N_2214,N_1130,N_1091);
xnor U2215 (N_2215,N_197,N_1613);
or U2216 (N_2216,N_1332,N_1624);
nand U2217 (N_2217,N_232,N_1638);
nor U2218 (N_2218,N_1014,N_1686);
and U2219 (N_2219,N_1996,N_871);
nor U2220 (N_2220,N_1145,N_1477);
nand U2221 (N_2221,N_801,N_266);
and U2222 (N_2222,N_1995,N_848);
nand U2223 (N_2223,N_1482,N_99);
or U2224 (N_2224,N_1015,N_915);
and U2225 (N_2225,N_858,N_340);
nor U2226 (N_2226,N_1107,N_674);
xor U2227 (N_2227,N_1310,N_1516);
xnor U2228 (N_2228,N_883,N_1169);
and U2229 (N_2229,N_764,N_1540);
nor U2230 (N_2230,N_1728,N_165);
and U2231 (N_2231,N_1445,N_1227);
or U2232 (N_2232,N_1717,N_1543);
nand U2233 (N_2233,N_788,N_1630);
nor U2234 (N_2234,N_1565,N_1238);
nor U2235 (N_2235,N_671,N_650);
xnor U2236 (N_2236,N_815,N_520);
xor U2237 (N_2237,N_998,N_1096);
or U2238 (N_2238,N_254,N_1265);
nand U2239 (N_2239,N_220,N_1991);
or U2240 (N_2240,N_986,N_1299);
nor U2241 (N_2241,N_1016,N_731);
xor U2242 (N_2242,N_1824,N_620);
and U2243 (N_2243,N_1653,N_434);
and U2244 (N_2244,N_1334,N_619);
xnor U2245 (N_2245,N_1163,N_1655);
or U2246 (N_2246,N_1628,N_1967);
nand U2247 (N_2247,N_1061,N_1011);
nor U2248 (N_2248,N_539,N_543);
nor U2249 (N_2249,N_538,N_1461);
or U2250 (N_2250,N_1495,N_1648);
nand U2251 (N_2251,N_1088,N_617);
or U2252 (N_2252,N_949,N_1920);
nand U2253 (N_2253,N_854,N_458);
and U2254 (N_2254,N_1382,N_985);
nand U2255 (N_2255,N_1984,N_151);
nand U2256 (N_2256,N_1243,N_1287);
and U2257 (N_2257,N_1114,N_279);
and U2258 (N_2258,N_353,N_1970);
nand U2259 (N_2259,N_1705,N_121);
nand U2260 (N_2260,N_551,N_1961);
nor U2261 (N_2261,N_9,N_1415);
or U2262 (N_2262,N_689,N_751);
or U2263 (N_2263,N_1651,N_1303);
nor U2264 (N_2264,N_81,N_877);
and U2265 (N_2265,N_1186,N_820);
or U2266 (N_2266,N_1795,N_1498);
nand U2267 (N_2267,N_236,N_199);
or U2268 (N_2268,N_1144,N_1408);
nand U2269 (N_2269,N_51,N_248);
or U2270 (N_2270,N_1492,N_264);
and U2271 (N_2271,N_338,N_94);
or U2272 (N_2272,N_1376,N_1286);
nor U2273 (N_2273,N_641,N_1816);
nor U2274 (N_2274,N_1217,N_1657);
xor U2275 (N_2275,N_1340,N_22);
nor U2276 (N_2276,N_1663,N_1939);
or U2277 (N_2277,N_1378,N_96);
and U2278 (N_2278,N_723,N_987);
xor U2279 (N_2279,N_157,N_761);
and U2280 (N_2280,N_154,N_1808);
nand U2281 (N_2281,N_1810,N_455);
and U2282 (N_2282,N_826,N_108);
and U2283 (N_2283,N_1818,N_1975);
nand U2284 (N_2284,N_1008,N_1596);
nor U2285 (N_2285,N_969,N_1703);
nor U2286 (N_2286,N_1572,N_1781);
and U2287 (N_2287,N_1988,N_1894);
nor U2288 (N_2288,N_890,N_950);
and U2289 (N_2289,N_24,N_879);
xnor U2290 (N_2290,N_278,N_25);
nand U2291 (N_2291,N_655,N_1990);
nand U2292 (N_2292,N_624,N_1216);
xor U2293 (N_2293,N_462,N_903);
and U2294 (N_2294,N_553,N_770);
and U2295 (N_2295,N_263,N_677);
or U2296 (N_2296,N_1583,N_1264);
nor U2297 (N_2297,N_43,N_647);
or U2298 (N_2298,N_1765,N_719);
and U2299 (N_2299,N_1069,N_1700);
nand U2300 (N_2300,N_1000,N_222);
xnor U2301 (N_2301,N_244,N_1647);
nor U2302 (N_2302,N_1177,N_466);
and U2303 (N_2303,N_705,N_713);
nor U2304 (N_2304,N_503,N_920);
or U2305 (N_2305,N_1769,N_924);
nand U2306 (N_2306,N_704,N_574);
or U2307 (N_2307,N_1573,N_1229);
nand U2308 (N_2308,N_10,N_1803);
and U2309 (N_2309,N_1850,N_798);
nand U2310 (N_2310,N_1554,N_1099);
xnor U2311 (N_2311,N_1814,N_1381);
nor U2312 (N_2312,N_1231,N_1896);
and U2313 (N_2313,N_275,N_736);
nor U2314 (N_2314,N_415,N_1040);
or U2315 (N_2315,N_1225,N_1538);
nor U2316 (N_2316,N_1587,N_1094);
and U2317 (N_2317,N_690,N_506);
nand U2318 (N_2318,N_717,N_406);
nor U2319 (N_2319,N_1568,N_93);
and U2320 (N_2320,N_523,N_238);
and U2321 (N_2321,N_164,N_1523);
nand U2322 (N_2322,N_765,N_901);
and U2323 (N_2323,N_533,N_1396);
and U2324 (N_2324,N_1992,N_1417);
nand U2325 (N_2325,N_835,N_802);
nand U2326 (N_2326,N_125,N_156);
or U2327 (N_2327,N_627,N_830);
or U2328 (N_2328,N_1876,N_521);
nor U2329 (N_2329,N_1932,N_760);
or U2330 (N_2330,N_1368,N_57);
and U2331 (N_2331,N_548,N_795);
nand U2332 (N_2332,N_62,N_1673);
or U2333 (N_2333,N_1319,N_443);
xnor U2334 (N_2334,N_47,N_1748);
xor U2335 (N_2335,N_846,N_566);
nand U2336 (N_2336,N_1480,N_831);
xor U2337 (N_2337,N_1406,N_836);
or U2338 (N_2338,N_629,N_1385);
and U2339 (N_2339,N_1275,N_1732);
xor U2340 (N_2340,N_1430,N_1730);
nor U2341 (N_2341,N_1923,N_1276);
and U2342 (N_2342,N_632,N_1913);
nor U2343 (N_2343,N_639,N_1353);
and U2344 (N_2344,N_596,N_1756);
nand U2345 (N_2345,N_1446,N_445);
nand U2346 (N_2346,N_928,N_8);
nor U2347 (N_2347,N_180,N_251);
or U2348 (N_2348,N_482,N_1078);
nand U2349 (N_2349,N_1136,N_1989);
nor U2350 (N_2350,N_30,N_1140);
nor U2351 (N_2351,N_564,N_1393);
nor U2352 (N_2352,N_358,N_1502);
or U2353 (N_2353,N_327,N_1342);
nor U2354 (N_2354,N_1714,N_19);
and U2355 (N_2355,N_1968,N_945);
or U2356 (N_2356,N_1442,N_1106);
xnor U2357 (N_2357,N_1672,N_1277);
nor U2358 (N_2358,N_1559,N_1787);
xnor U2359 (N_2359,N_613,N_243);
and U2360 (N_2360,N_268,N_910);
xnor U2361 (N_2361,N_995,N_369);
or U2362 (N_2362,N_668,N_927);
nand U2363 (N_2363,N_583,N_571);
or U2364 (N_2364,N_379,N_1884);
xnor U2365 (N_2365,N_1699,N_1490);
nor U2366 (N_2366,N_1937,N_308);
nor U2367 (N_2367,N_430,N_1839);
nand U2368 (N_2368,N_1149,N_780);
and U2369 (N_2369,N_1997,N_1561);
nor U2370 (N_2370,N_1060,N_1308);
and U2371 (N_2371,N_282,N_1082);
or U2372 (N_2372,N_1199,N_1339);
or U2373 (N_2373,N_1467,N_130);
and U2374 (N_2374,N_1586,N_252);
and U2375 (N_2375,N_1028,N_618);
xnor U2376 (N_2376,N_160,N_1458);
and U2377 (N_2377,N_1782,N_532);
nor U2378 (N_2378,N_407,N_1077);
or U2379 (N_2379,N_1439,N_397);
xor U2380 (N_2380,N_718,N_420);
xor U2381 (N_2381,N_594,N_1420);
nand U2382 (N_2382,N_1054,N_259);
xnor U2383 (N_2383,N_1954,N_1632);
nand U2384 (N_2384,N_317,N_1418);
and U2385 (N_2385,N_208,N_142);
nand U2386 (N_2386,N_1683,N_1399);
and U2387 (N_2387,N_1030,N_1081);
nor U2388 (N_2388,N_905,N_1233);
or U2389 (N_2389,N_1880,N_694);
xnor U2390 (N_2390,N_1941,N_1752);
nand U2391 (N_2391,N_1244,N_822);
and U2392 (N_2392,N_1962,N_1840);
nand U2393 (N_2393,N_796,N_399);
nor U2394 (N_2394,N_351,N_876);
and U2395 (N_2395,N_400,N_1307);
nand U2396 (N_2396,N_1662,N_1972);
or U2397 (N_2397,N_838,N_442);
xnor U2398 (N_2398,N_75,N_1902);
nor U2399 (N_2399,N_231,N_1022);
nand U2400 (N_2400,N_12,N_390);
and U2401 (N_2401,N_1940,N_1949);
xor U2402 (N_2402,N_1148,N_227);
nor U2403 (N_2403,N_1964,N_1074);
and U2404 (N_2404,N_149,N_1617);
nand U2405 (N_2405,N_177,N_567);
or U2406 (N_2406,N_1533,N_819);
nor U2407 (N_2407,N_948,N_1875);
nor U2408 (N_2408,N_1377,N_515);
nand U2409 (N_2409,N_490,N_750);
or U2410 (N_2410,N_1602,N_207);
nand U2411 (N_2411,N_393,N_1423);
or U2412 (N_2412,N_961,N_45);
nor U2413 (N_2413,N_896,N_1391);
and U2414 (N_2414,N_245,N_769);
nor U2415 (N_2415,N_1236,N_1142);
or U2416 (N_2416,N_706,N_1812);
xor U2417 (N_2417,N_753,N_433);
nor U2418 (N_2418,N_842,N_1293);
nor U2419 (N_2419,N_939,N_958);
nor U2420 (N_2420,N_109,N_1641);
xnor U2421 (N_2421,N_1232,N_849);
and U2422 (N_2422,N_1122,N_1741);
or U2423 (N_2423,N_1679,N_591);
nand U2424 (N_2424,N_1973,N_488);
and U2425 (N_2425,N_1688,N_1908);
nand U2426 (N_2426,N_1373,N_128);
nor U2427 (N_2427,N_395,N_21);
xnor U2428 (N_2428,N_1235,N_667);
or U2429 (N_2429,N_1404,N_1846);
xor U2430 (N_2430,N_562,N_1836);
or U2431 (N_2431,N_811,N_561);
or U2432 (N_2432,N_584,N_79);
nor U2433 (N_2433,N_527,N_1604);
or U2434 (N_2434,N_558,N_1009);
nand U2435 (N_2435,N_1330,N_1306);
nor U2436 (N_2436,N_46,N_1659);
and U2437 (N_2437,N_1936,N_1154);
or U2438 (N_2438,N_1202,N_288);
nand U2439 (N_2439,N_766,N_1476);
xor U2440 (N_2440,N_1702,N_841);
xnor U2441 (N_2441,N_1359,N_1751);
xnor U2442 (N_2442,N_1434,N_797);
nand U2443 (N_2443,N_1100,N_793);
xnor U2444 (N_2444,N_803,N_106);
nor U2445 (N_2445,N_757,N_313);
and U2446 (N_2446,N_531,N_1395);
or U2447 (N_2447,N_941,N_888);
and U2448 (N_2448,N_1212,N_373);
xnor U2449 (N_2449,N_783,N_1012);
and U2450 (N_2450,N_1046,N_241);
nor U2451 (N_2451,N_89,N_1076);
or U2452 (N_2452,N_363,N_1527);
xnor U2453 (N_2453,N_83,N_964);
nand U2454 (N_2454,N_1825,N_331);
or U2455 (N_2455,N_720,N_1883);
xor U2456 (N_2456,N_1337,N_267);
nor U2457 (N_2457,N_170,N_346);
and U2458 (N_2458,N_891,N_300);
nand U2459 (N_2459,N_40,N_1822);
xor U2460 (N_2460,N_864,N_1993);
xor U2461 (N_2461,N_573,N_739);
or U2462 (N_2462,N_606,N_1150);
xnor U2463 (N_2463,N_1654,N_332);
nor U2464 (N_2464,N_726,N_1440);
or U2465 (N_2465,N_944,N_648);
and U2466 (N_2466,N_669,N_143);
nor U2467 (N_2467,N_885,N_741);
or U2468 (N_2468,N_475,N_742);
xor U2469 (N_2469,N_1472,N_1497);
and U2470 (N_2470,N_1187,N_1026);
xnor U2471 (N_2471,N_1245,N_14);
and U2472 (N_2472,N_1089,N_182);
nor U2473 (N_2473,N_1609,N_1558);
or U2474 (N_2474,N_425,N_250);
nand U2475 (N_2475,N_1020,N_889);
nand U2476 (N_2476,N_773,N_805);
nor U2477 (N_2477,N_1656,N_1447);
and U2478 (N_2478,N_1698,N_1783);
or U2479 (N_2479,N_1105,N_1288);
or U2480 (N_2480,N_1892,N_1075);
or U2481 (N_2481,N_138,N_153);
and U2482 (N_2482,N_1948,N_602);
nand U2483 (N_2483,N_1017,N_1083);
or U2484 (N_2484,N_1098,N_1379);
or U2485 (N_2485,N_1336,N_1721);
or U2486 (N_2486,N_1517,N_105);
and U2487 (N_2487,N_942,N_1058);
xor U2488 (N_2488,N_355,N_1102);
nand U2489 (N_2489,N_262,N_1178);
nand U2490 (N_2490,N_1175,N_257);
and U2491 (N_2491,N_1852,N_1033);
and U2492 (N_2492,N_86,N_700);
or U2493 (N_2493,N_70,N_255);
or U2494 (N_2494,N_752,N_1433);
nor U2495 (N_2495,N_1092,N_246);
xor U2496 (N_2496,N_181,N_1294);
and U2497 (N_2497,N_1608,N_1475);
xnor U2498 (N_2498,N_71,N_214);
nand U2499 (N_2499,N_1635,N_325);
xnor U2500 (N_2500,N_1979,N_1466);
nor U2501 (N_2501,N_167,N_1826);
xnor U2502 (N_2502,N_683,N_1534);
nand U2503 (N_2503,N_1398,N_1849);
nand U2504 (N_2504,N_1919,N_758);
and U2505 (N_2505,N_1179,N_15);
or U2506 (N_2506,N_69,N_1184);
nand U2507 (N_2507,N_1676,N_107);
or U2508 (N_2508,N_444,N_508);
or U2509 (N_2509,N_392,N_1313);
nor U2510 (N_2510,N_919,N_172);
nand U2511 (N_2511,N_1485,N_194);
or U2512 (N_2512,N_1575,N_1068);
nor U2513 (N_2513,N_1943,N_777);
nand U2514 (N_2514,N_1854,N_1520);
or U2515 (N_2515,N_1513,N_1384);
or U2516 (N_2516,N_1510,N_695);
and U2517 (N_2517,N_1166,N_1811);
nand U2518 (N_2518,N_209,N_1899);
nor U2519 (N_2519,N_1633,N_1329);
nor U2520 (N_2520,N_487,N_1690);
nand U2521 (N_2521,N_1509,N_500);
nor U2522 (N_2522,N_1710,N_129);
nand U2523 (N_2523,N_1258,N_1219);
and U2524 (N_2524,N_1311,N_1685);
xnor U2525 (N_2525,N_972,N_1909);
nand U2526 (N_2526,N_404,N_1588);
and U2527 (N_2527,N_1252,N_541);
or U2528 (N_2528,N_588,N_1032);
xor U2529 (N_2529,N_1847,N_333);
nor U2530 (N_2530,N_82,N_1317);
nand U2531 (N_2531,N_1347,N_234);
nor U2532 (N_2532,N_1388,N_1059);
and U2533 (N_2533,N_1546,N_505);
or U2534 (N_2534,N_1969,N_1370);
nor U2535 (N_2535,N_412,N_1090);
nand U2536 (N_2536,N_76,N_787);
nor U2537 (N_2537,N_1117,N_1725);
xnor U2538 (N_2538,N_97,N_271);
nor U2539 (N_2539,N_843,N_276);
and U2540 (N_2540,N_1247,N_1890);
nand U2541 (N_2541,N_131,N_1147);
and U2542 (N_2542,N_374,N_1261);
nand U2543 (N_2543,N_196,N_616);
nand U2544 (N_2544,N_1837,N_1521);
or U2545 (N_2545,N_850,N_665);
or U2546 (N_2546,N_1355,N_290);
xnor U2547 (N_2547,N_1185,N_1499);
or U2548 (N_2548,N_1003,N_1341);
or U2549 (N_2549,N_1454,N_991);
nor U2550 (N_2550,N_526,N_1981);
xor U2551 (N_2551,N_307,N_1478);
nand U2552 (N_2552,N_1872,N_1985);
nand U2553 (N_2553,N_100,N_354);
xnor U2554 (N_2554,N_1207,N_862);
nor U2555 (N_2555,N_419,N_78);
xnor U2556 (N_2556,N_1104,N_1131);
nand U2557 (N_2557,N_1530,N_1743);
and U2558 (N_2558,N_599,N_347);
nor U2559 (N_2559,N_1815,N_852);
xor U2560 (N_2560,N_41,N_416);
and U2561 (N_2561,N_1210,N_1162);
nor U2562 (N_2562,N_1400,N_1537);
nand U2563 (N_2563,N_310,N_114);
and U2564 (N_2564,N_1284,N_1731);
nand U2565 (N_2565,N_568,N_195);
or U2566 (N_2566,N_1950,N_1271);
nand U2567 (N_2567,N_1844,N_240);
nor U2568 (N_2568,N_893,N_923);
nand U2569 (N_2569,N_1958,N_1916);
xor U2570 (N_2570,N_124,N_28);
and U2571 (N_2571,N_1670,N_980);
nor U2572 (N_2572,N_1464,N_918);
nor U2573 (N_2573,N_118,N_233);
or U2574 (N_2574,N_1156,N_1594);
and U2575 (N_2575,N_676,N_206);
xnor U2576 (N_2576,N_328,N_1465);
or U2577 (N_2577,N_992,N_743);
or U2578 (N_2578,N_1226,N_341);
nand U2579 (N_2579,N_179,N_1868);
or U2580 (N_2580,N_1871,N_651);
or U2581 (N_2581,N_1865,N_1869);
xnor U2582 (N_2582,N_450,N_524);
nand U2583 (N_2583,N_789,N_383);
nand U2584 (N_2584,N_921,N_91);
nor U2585 (N_2585,N_859,N_1734);
nor U2586 (N_2586,N_983,N_493);
xnor U2587 (N_2587,N_1775,N_225);
xor U2588 (N_2588,N_1443,N_1511);
or U2589 (N_2589,N_479,N_1085);
nor U2590 (N_2590,N_737,N_219);
nand U2591 (N_2591,N_387,N_316);
and U2592 (N_2592,N_935,N_1426);
nand U2593 (N_2593,N_740,N_1928);
xor U2594 (N_2594,N_171,N_216);
or U2595 (N_2595,N_1324,N_1640);
nor U2596 (N_2596,N_360,N_1006);
and U2597 (N_2597,N_817,N_1945);
nand U2598 (N_2598,N_1644,N_1206);
xor U2599 (N_2599,N_952,N_814);
nand U2600 (N_2600,N_1471,N_292);
and U2601 (N_2601,N_204,N_1905);
and U2602 (N_2602,N_1666,N_692);
or U2603 (N_2603,N_1934,N_291);
nor U2604 (N_2604,N_784,N_386);
or U2605 (N_2605,N_1867,N_211);
xor U2606 (N_2606,N_1354,N_42);
or U2607 (N_2607,N_559,N_34);
xnor U2608 (N_2608,N_1257,N_85);
and U2609 (N_2609,N_320,N_492);
nand U2610 (N_2610,N_1912,N_654);
or U2611 (N_2611,N_60,N_1914);
or U2612 (N_2612,N_1532,N_409);
xnor U2613 (N_2613,N_1366,N_217);
nor U2614 (N_2614,N_1203,N_1621);
or U2615 (N_2615,N_1021,N_6);
or U2616 (N_2616,N_304,N_408);
nand U2617 (N_2617,N_283,N_1749);
or U2618 (N_2618,N_1548,N_1164);
and U2619 (N_2619,N_698,N_1525);
nand U2620 (N_2620,N_293,N_1593);
nand U2621 (N_2621,N_790,N_44);
nor U2622 (N_2622,N_1539,N_1253);
nor U2623 (N_2623,N_1994,N_965);
xor U2624 (N_2624,N_1448,N_806);
and U2625 (N_2625,N_887,N_389);
nand U2626 (N_2626,N_1582,N_1763);
xor U2627 (N_2627,N_472,N_1052);
xor U2628 (N_2628,N_661,N_642);
xor U2629 (N_2629,N_1298,N_525);
or U2630 (N_2630,N_563,N_1504);
or U2631 (N_2631,N_498,N_330);
xnor U2632 (N_2632,N_993,N_401);
or U2633 (N_2633,N_1125,N_1777);
or U2634 (N_2634,N_855,N_213);
xor U2635 (N_2635,N_845,N_163);
xnor U2636 (N_2636,N_1736,N_678);
xnor U2637 (N_2637,N_1924,N_869);
or U2638 (N_2638,N_440,N_684);
or U2639 (N_2639,N_1784,N_133);
nor U2640 (N_2640,N_111,N_396);
xnor U2641 (N_2641,N_1614,N_65);
and U2642 (N_2642,N_1841,N_1116);
or U2643 (N_2643,N_912,N_187);
and U2644 (N_2644,N_1889,N_1494);
xor U2645 (N_2645,N_186,N_1925);
nor U2646 (N_2646,N_1412,N_634);
and U2647 (N_2647,N_1338,N_1419);
or U2648 (N_2648,N_1198,N_1677);
and U2649 (N_2649,N_155,N_829);
nor U2650 (N_2650,N_1759,N_1933);
nor U2651 (N_2651,N_1863,N_1432);
xor U2652 (N_2652,N_1806,N_193);
xor U2653 (N_2653,N_996,N_1372);
xnor U2654 (N_2654,N_1864,N_1965);
nor U2655 (N_2655,N_679,N_973);
and U2656 (N_2656,N_432,N_80);
nor U2657 (N_2657,N_16,N_137);
or U2658 (N_2658,N_1470,N_930);
or U2659 (N_2659,N_1629,N_1590);
nand U2660 (N_2660,N_897,N_1866);
or U2661 (N_2661,N_832,N_716);
nor U2662 (N_2662,N_560,N_249);
nor U2663 (N_2663,N_1196,N_688);
nor U2664 (N_2664,N_547,N_577);
nand U2665 (N_2665,N_1740,N_336);
or U2666 (N_2666,N_572,N_636);
and U2667 (N_2667,N_1879,N_497);
xor U2668 (N_2668,N_693,N_1882);
or U2669 (N_2669,N_1256,N_202);
or U2670 (N_2670,N_1351,N_600);
xnor U2671 (N_2671,N_422,N_11);
and U2672 (N_2672,N_1737,N_1322);
nor U2673 (N_2673,N_74,N_183);
or U2674 (N_2674,N_1897,N_272);
xor U2675 (N_2675,N_653,N_349);
nand U2676 (N_2676,N_970,N_1281);
nor U2677 (N_2677,N_672,N_1333);
nand U2678 (N_2678,N_837,N_484);
or U2679 (N_2679,N_535,N_732);
nor U2680 (N_2680,N_101,N_1486);
nor U2681 (N_2681,N_1073,N_1108);
nand U2682 (N_2682,N_122,N_1189);
and U2683 (N_2683,N_1251,N_975);
and U2684 (N_2684,N_1618,N_622);
nor U2685 (N_2685,N_1079,N_1093);
nor U2686 (N_2686,N_102,N_1259);
xor U2687 (N_2687,N_192,N_1760);
nand U2688 (N_2688,N_1165,N_609);
nand U2689 (N_2689,N_1005,N_652);
or U2690 (N_2690,N_1817,N_1407);
nand U2691 (N_2691,N_1712,N_242);
nor U2692 (N_2692,N_1460,N_168);
xor U2693 (N_2693,N_1754,N_1999);
nand U2694 (N_2694,N_886,N_212);
or U2695 (N_2695,N_1362,N_92);
and U2696 (N_2696,N_771,N_473);
and U2697 (N_2697,N_343,N_1560);
nor U2698 (N_2698,N_1190,N_1757);
xor U2699 (N_2699,N_1305,N_540);
or U2700 (N_2700,N_1772,N_378);
and U2701 (N_2701,N_1870,N_1804);
nor U2702 (N_2702,N_315,N_1438);
and U2703 (N_2703,N_309,N_1823);
nor U2704 (N_2704,N_1290,N_946);
nand U2705 (N_2705,N_1312,N_711);
nand U2706 (N_2706,N_605,N_344);
xor U2707 (N_2707,N_1976,N_612);
nand U2708 (N_2708,N_762,N_50);
or U2709 (N_2709,N_1788,N_218);
xor U2710 (N_2710,N_702,N_441);
xnor U2711 (N_2711,N_828,N_1269);
nor U2712 (N_2712,N_1036,N_1067);
nor U2713 (N_2713,N_1375,N_1200);
and U2714 (N_2714,N_1584,N_979);
and U2715 (N_2715,N_1413,N_1515);
nor U2716 (N_2716,N_1627,N_48);
nand U2717 (N_2717,N_1886,N_1983);
nor U2718 (N_2718,N_1620,N_439);
or U2719 (N_2719,N_1790,N_1696);
xor U2720 (N_2720,N_549,N_176);
nand U2721 (N_2721,N_402,N_1128);
and U2722 (N_2722,N_1829,N_1544);
xnor U2723 (N_2723,N_900,N_1946);
or U2724 (N_2724,N_1181,N_687);
nand U2725 (N_2725,N_1141,N_699);
nand U2726 (N_2726,N_1518,N_898);
nand U2727 (N_2727,N_856,N_782);
or U2728 (N_2728,N_169,N_1821);
nor U2729 (N_2729,N_715,N_1220);
or U2730 (N_2730,N_1369,N_1645);
and U2731 (N_2731,N_123,N_305);
nor U2732 (N_2732,N_1450,N_280);
nor U2733 (N_2733,N_734,N_1421);
nand U2734 (N_2734,N_477,N_302);
or U2735 (N_2735,N_1044,N_827);
and U2736 (N_2736,N_1228,N_1842);
or U2737 (N_2737,N_502,N_1623);
or U2738 (N_2738,N_926,N_27);
and U2739 (N_2739,N_1424,N_1684);
nor U2740 (N_2740,N_1024,N_1292);
and U2741 (N_2741,N_1039,N_261);
nand U2742 (N_2742,N_1597,N_645);
or U2743 (N_2743,N_1636,N_1820);
and U2744 (N_2744,N_555,N_749);
and U2745 (N_2745,N_940,N_1159);
or U2746 (N_2746,N_1791,N_68);
or U2747 (N_2747,N_1487,N_162);
nand U2748 (N_2748,N_1953,N_1715);
and U2749 (N_2749,N_550,N_712);
nand U2750 (N_2750,N_755,N_999);
nand U2751 (N_2751,N_1681,N_1529);
or U2752 (N_2752,N_657,N_1158);
xnor U2753 (N_2753,N_235,N_866);
xnor U2754 (N_2754,N_337,N_1729);
nor U2755 (N_2755,N_1716,N_1455);
nor U2756 (N_2756,N_874,N_1650);
and U2757 (N_2757,N_381,N_556);
or U2758 (N_2758,N_67,N_857);
xor U2759 (N_2759,N_557,N_198);
or U2760 (N_2760,N_1043,N_1735);
nand U2761 (N_2761,N_1577,N_1402);
nand U2762 (N_2762,N_809,N_1134);
xnor U2763 (N_2763,N_1132,N_899);
nand U2764 (N_2764,N_1535,N_1255);
or U2765 (N_2765,N_1,N_664);
xor U2766 (N_2766,N_1861,N_1911);
and U2767 (N_2767,N_1045,N_451);
and U2768 (N_2768,N_631,N_1197);
xor U2769 (N_2769,N_485,N_1631);
and U2770 (N_2770,N_1522,N_312);
and U2771 (N_2771,N_1851,N_989);
nand U2772 (N_2772,N_2,N_229);
xor U2773 (N_2773,N_158,N_411);
nand U2774 (N_2774,N_1927,N_1960);
nor U2775 (N_2775,N_511,N_256);
nor U2776 (N_2776,N_1674,N_1250);
nand U2777 (N_2777,N_1767,N_1126);
xnor U2778 (N_2778,N_364,N_460);
and U2779 (N_2779,N_1694,N_906);
and U2780 (N_2780,N_115,N_640);
nor U2781 (N_2781,N_626,N_1528);
nand U2782 (N_2782,N_405,N_90);
nand U2783 (N_2783,N_1230,N_517);
xor U2784 (N_2784,N_1785,N_1615);
or U2785 (N_2785,N_974,N_870);
xnor U2786 (N_2786,N_5,N_956);
xnor U2787 (N_2787,N_1938,N_20);
nor U2788 (N_2788,N_1764,N_289);
nand U2789 (N_2789,N_1649,N_1240);
xor U2790 (N_2790,N_1738,N_1474);
nand U2791 (N_2791,N_510,N_230);
nor U2792 (N_2792,N_1585,N_1365);
xor U2793 (N_2793,N_116,N_481);
and U2794 (N_2794,N_1888,N_1349);
or U2795 (N_2795,N_1512,N_1211);
nor U2796 (N_2796,N_1557,N_779);
nor U2797 (N_2797,N_1320,N_1401);
or U2798 (N_2798,N_1646,N_522);
and U2799 (N_2799,N_127,N_237);
nor U2800 (N_2800,N_1441,N_174);
and U2801 (N_2801,N_303,N_1720);
xnor U2802 (N_2802,N_1428,N_110);
nand U2803 (N_2803,N_447,N_189);
nor U2804 (N_2804,N_1526,N_398);
nor U2805 (N_2805,N_1301,N_839);
nand U2806 (N_2806,N_1542,N_1285);
and U2807 (N_2807,N_1805,N_663);
nor U2808 (N_2808,N_1862,N_1209);
nor U2809 (N_2809,N_791,N_804);
nand U2810 (N_2810,N_735,N_1853);
and U2811 (N_2811,N_922,N_1689);
nand U2812 (N_2812,N_1037,N_361);
nand U2813 (N_2813,N_1747,N_1801);
or U2814 (N_2814,N_570,N_184);
nand U2815 (N_2815,N_469,N_1974);
and U2816 (N_2816,N_152,N_685);
or U2817 (N_2817,N_1350,N_1567);
xnor U2818 (N_2818,N_0,N_1262);
nor U2819 (N_2819,N_1566,N_468);
nor U2820 (N_2820,N_465,N_1887);
and U2821 (N_2821,N_552,N_728);
or U2822 (N_2822,N_270,N_1267);
and U2823 (N_2823,N_1589,N_772);
xor U2824 (N_2824,N_1762,N_467);
or U2825 (N_2825,N_423,N_1753);
or U2826 (N_2826,N_1266,N_410);
or U2827 (N_2827,N_63,N_691);
nand U2828 (N_2828,N_1592,N_833);
nor U2829 (N_2829,N_1917,N_1057);
xor U2830 (N_2830,N_1843,N_638);
xor U2831 (N_2831,N_1170,N_662);
nand U2832 (N_2832,N_1124,N_298);
xor U2833 (N_2833,N_1832,N_269);
and U2834 (N_2834,N_812,N_1193);
nor U2835 (N_2835,N_17,N_721);
or U2836 (N_2836,N_908,N_585);
or U2837 (N_2837,N_1904,N_438);
nand U2838 (N_2838,N_1768,N_1295);
xor U2839 (N_2839,N_1462,N_593);
nand U2840 (N_2840,N_1505,N_35);
and U2841 (N_2841,N_1489,N_431);
xor U2842 (N_2842,N_1612,N_1019);
nor U2843 (N_2843,N_1208,N_978);
xnor U2844 (N_2844,N_1963,N_1056);
xnor U2845 (N_2845,N_1603,N_1389);
nand U2846 (N_2846,N_428,N_644);
and U2847 (N_2847,N_545,N_456);
xnor U2848 (N_2848,N_382,N_937);
nor U2849 (N_2849,N_1205,N_1086);
nand U2850 (N_2850,N_1112,N_1493);
and U2851 (N_2851,N_501,N_1773);
and U2852 (N_2852,N_1072,N_637);
nor U2853 (N_2853,N_603,N_18);
or U2854 (N_2854,N_1813,N_1118);
nor U2855 (N_2855,N_834,N_1153);
nand U2856 (N_2856,N_1947,N_1742);
or U2857 (N_2857,N_210,N_968);
and U2858 (N_2858,N_625,N_1797);
or U2859 (N_2859,N_1549,N_1835);
nand U2860 (N_2860,N_853,N_166);
nor U2861 (N_2861,N_816,N_1172);
nand U2862 (N_2862,N_1405,N_1893);
nand U2863 (N_2863,N_452,N_146);
and U2864 (N_2864,N_1263,N_29);
xor U2865 (N_2865,N_1129,N_87);
or U2866 (N_2866,N_1838,N_1327);
or U2867 (N_2867,N_1503,N_880);
or U2868 (N_2868,N_1346,N_4);
or U2869 (N_2869,N_294,N_377);
nand U2870 (N_2870,N_1173,N_878);
xnor U2871 (N_2871,N_1874,N_56);
and U2872 (N_2872,N_1691,N_362);
or U2873 (N_2873,N_1123,N_1380);
xnor U2874 (N_2874,N_1304,N_1514);
and U2875 (N_2875,N_929,N_534);
xor U2876 (N_2876,N_437,N_774);
nor U2877 (N_2877,N_322,N_514);
and U2878 (N_2878,N_1802,N_754);
and U2879 (N_2879,N_1895,N_1444);
and U2880 (N_2880,N_955,N_825);
nor U2881 (N_2881,N_284,N_1371);
nor U2882 (N_2882,N_66,N_221);
xor U2883 (N_2883,N_424,N_701);
nand U2884 (N_2884,N_1191,N_1827);
or U2885 (N_2885,N_776,N_1481);
and U2886 (N_2886,N_546,N_708);
nor U2887 (N_2887,N_1986,N_1591);
xor U2888 (N_2888,N_3,N_88);
and U2889 (N_2889,N_1071,N_1055);
xnor U2890 (N_2890,N_529,N_1601);
nand U2891 (N_2891,N_722,N_1157);
xnor U2892 (N_2892,N_882,N_981);
nor U2893 (N_2893,N_1453,N_675);
or U2894 (N_2894,N_301,N_1241);
nor U2895 (N_2895,N_1719,N_95);
or U2896 (N_2896,N_976,N_1562);
and U2897 (N_2897,N_73,N_55);
nor U2898 (N_2898,N_917,N_951);
xor U2899 (N_2899,N_847,N_902);
xor U2900 (N_2900,N_707,N_1856);
xor U2901 (N_2901,N_1744,N_365);
xnor U2902 (N_2902,N_136,N_1855);
nand U2903 (N_2903,N_1563,N_265);
nand U2904 (N_2904,N_1309,N_1569);
and U2905 (N_2905,N_1900,N_907);
or U2906 (N_2906,N_1115,N_26);
and U2907 (N_2907,N_144,N_646);
nor U2908 (N_2908,N_963,N_528);
xnor U2909 (N_2909,N_1701,N_982);
nor U2910 (N_2910,N_1898,N_457);
and U2911 (N_2911,N_1331,N_516);
and U2912 (N_2912,N_1363,N_223);
or U2913 (N_2913,N_598,N_860);
xor U2914 (N_2914,N_1161,N_894);
nand U2915 (N_2915,N_1323,N_1335);
xnor U2916 (N_2916,N_578,N_376);
and U2917 (N_2917,N_681,N_1611);
nor U2918 (N_2918,N_1204,N_1809);
nor U2919 (N_2919,N_188,N_253);
xor U2920 (N_2920,N_1167,N_763);
xor U2921 (N_2921,N_1634,N_1035);
xnor U2922 (N_2922,N_1807,N_792);
nor U2923 (N_2923,N_1242,N_1605);
and U2924 (N_2924,N_52,N_1834);
and U2925 (N_2925,N_1796,N_1239);
xnor U2926 (N_2926,N_1427,N_778);
or U2927 (N_2927,N_478,N_821);
nor U2928 (N_2928,N_370,N_1746);
nor U2929 (N_2929,N_1901,N_1053);
xnor U2930 (N_2930,N_1726,N_1570);
and U2931 (N_2931,N_352,N_1484);
or U2932 (N_2932,N_1435,N_1468);
nor U2933 (N_2933,N_1300,N_1390);
and U2934 (N_2934,N_865,N_1137);
nor U2935 (N_2935,N_1095,N_1302);
nand U2936 (N_2936,N_1101,N_463);
nor U2937 (N_2937,N_461,N_1857);
nand U2938 (N_2938,N_799,N_670);
nor U2939 (N_2939,N_1146,N_384);
or U2940 (N_2940,N_1031,N_1616);
and U2941 (N_2941,N_104,N_1833);
nand U2942 (N_2942,N_807,N_1682);
xnor U2943 (N_2943,N_1708,N_971);
or U2944 (N_2944,N_1111,N_295);
xor U2945 (N_2945,N_579,N_1215);
or U2946 (N_2946,N_1903,N_542);
or U2947 (N_2947,N_775,N_319);
and U2948 (N_2948,N_1580,N_1237);
nor U2949 (N_2949,N_1722,N_1180);
xnor U2950 (N_2950,N_366,N_1103);
xor U2951 (N_2951,N_139,N_990);
and U2952 (N_2952,N_1786,N_686);
and U2953 (N_2953,N_623,N_943);
or U2954 (N_2954,N_1249,N_658);
and U2955 (N_2955,N_953,N_909);
nor U2956 (N_2956,N_454,N_1531);
nor U2957 (N_2957,N_1410,N_745);
or U2958 (N_2958,N_1831,N_1213);
and U2959 (N_2959,N_1344,N_1194);
xor U2960 (N_2960,N_1425,N_581);
nor U2961 (N_2961,N_1687,N_448);
or U2962 (N_2962,N_1750,N_1978);
xnor U2963 (N_2963,N_512,N_709);
nor U2964 (N_2964,N_1449,N_1971);
nor U2965 (N_2965,N_98,N_135);
nor U2966 (N_2966,N_1873,N_932);
and U2967 (N_2967,N_875,N_1711);
xnor U2968 (N_2968,N_190,N_1830);
or U2969 (N_2969,N_984,N_329);
xnor U2970 (N_2970,N_554,N_342);
xnor U2971 (N_2971,N_323,N_23);
and U2972 (N_2972,N_1007,N_334);
and U2973 (N_2973,N_1042,N_1004);
nor U2974 (N_2974,N_1171,N_1639);
nand U2975 (N_2975,N_1049,N_1541);
and U2976 (N_2976,N_471,N_258);
nor U2977 (N_2977,N_1774,N_394);
xnor U2978 (N_2978,N_1234,N_84);
nand U2979 (N_2979,N_1326,N_595);
xnor U2980 (N_2980,N_1248,N_1034);
xnor U2981 (N_2981,N_113,N_1328);
or U2982 (N_2982,N_601,N_1348);
nand U2983 (N_2983,N_1709,N_610);
xnor U2984 (N_2984,N_421,N_1793);
nand U2985 (N_2985,N_1062,N_1907);
nor U2986 (N_2986,N_178,N_913);
or U2987 (N_2987,N_536,N_759);
nor U2988 (N_2988,N_103,N_1987);
xnor U2989 (N_2989,N_1139,N_1409);
nand U2990 (N_2990,N_380,N_1120);
nor U2991 (N_2991,N_1789,N_1929);
xnor U2992 (N_2992,N_1877,N_1551);
nor U2993 (N_2993,N_1192,N_936);
nor U2994 (N_2994,N_1451,N_1704);
nor U2995 (N_2995,N_72,N_824);
xnor U2996 (N_2996,N_1064,N_1506);
or U2997 (N_2997,N_537,N_738);
nand U2998 (N_2998,N_175,N_449);
and U2999 (N_2999,N_367,N_350);
or U3000 (N_3000,N_1496,N_1798);
xnor U3001 (N_3001,N_1825,N_196);
nor U3002 (N_3002,N_607,N_1975);
nor U3003 (N_3003,N_907,N_1951);
and U3004 (N_3004,N_341,N_196);
nand U3005 (N_3005,N_732,N_994);
nand U3006 (N_3006,N_158,N_1512);
nor U3007 (N_3007,N_156,N_1174);
or U3008 (N_3008,N_234,N_1876);
nor U3009 (N_3009,N_918,N_205);
and U3010 (N_3010,N_1423,N_720);
and U3011 (N_3011,N_1283,N_932);
nand U3012 (N_3012,N_357,N_64);
or U3013 (N_3013,N_129,N_832);
xor U3014 (N_3014,N_947,N_1802);
nor U3015 (N_3015,N_1069,N_773);
or U3016 (N_3016,N_1806,N_1280);
xor U3017 (N_3017,N_1953,N_1061);
nand U3018 (N_3018,N_638,N_1257);
nand U3019 (N_3019,N_799,N_831);
or U3020 (N_3020,N_1511,N_1398);
or U3021 (N_3021,N_638,N_1692);
nand U3022 (N_3022,N_1286,N_1634);
nor U3023 (N_3023,N_1780,N_1459);
and U3024 (N_3024,N_94,N_1308);
xor U3025 (N_3025,N_889,N_849);
and U3026 (N_3026,N_1897,N_1492);
or U3027 (N_3027,N_651,N_245);
or U3028 (N_3028,N_579,N_657);
nand U3029 (N_3029,N_299,N_1736);
nor U3030 (N_3030,N_576,N_1868);
nor U3031 (N_3031,N_133,N_472);
and U3032 (N_3032,N_595,N_639);
nand U3033 (N_3033,N_1267,N_987);
nor U3034 (N_3034,N_86,N_353);
nand U3035 (N_3035,N_849,N_945);
or U3036 (N_3036,N_1074,N_1058);
xnor U3037 (N_3037,N_1413,N_1826);
nor U3038 (N_3038,N_1066,N_51);
nor U3039 (N_3039,N_847,N_1577);
or U3040 (N_3040,N_176,N_1078);
nand U3041 (N_3041,N_902,N_1779);
nand U3042 (N_3042,N_752,N_817);
or U3043 (N_3043,N_553,N_949);
nand U3044 (N_3044,N_795,N_419);
nor U3045 (N_3045,N_1837,N_1421);
nand U3046 (N_3046,N_303,N_148);
or U3047 (N_3047,N_1022,N_1544);
nand U3048 (N_3048,N_332,N_1923);
nand U3049 (N_3049,N_338,N_197);
nor U3050 (N_3050,N_1301,N_690);
and U3051 (N_3051,N_1452,N_181);
or U3052 (N_3052,N_990,N_1096);
or U3053 (N_3053,N_361,N_1159);
nor U3054 (N_3054,N_17,N_1061);
xor U3055 (N_3055,N_720,N_174);
xor U3056 (N_3056,N_722,N_1634);
nor U3057 (N_3057,N_1506,N_41);
xor U3058 (N_3058,N_1902,N_192);
nor U3059 (N_3059,N_415,N_657);
and U3060 (N_3060,N_268,N_909);
or U3061 (N_3061,N_279,N_1739);
nand U3062 (N_3062,N_788,N_1619);
nor U3063 (N_3063,N_1122,N_1111);
nand U3064 (N_3064,N_71,N_513);
or U3065 (N_3065,N_1783,N_1811);
or U3066 (N_3066,N_1363,N_1162);
and U3067 (N_3067,N_1047,N_947);
nor U3068 (N_3068,N_146,N_550);
and U3069 (N_3069,N_56,N_673);
nor U3070 (N_3070,N_1609,N_343);
nand U3071 (N_3071,N_973,N_544);
xor U3072 (N_3072,N_1945,N_593);
or U3073 (N_3073,N_910,N_441);
xnor U3074 (N_3074,N_886,N_1818);
nor U3075 (N_3075,N_1032,N_485);
nand U3076 (N_3076,N_1174,N_1899);
or U3077 (N_3077,N_1784,N_920);
or U3078 (N_3078,N_591,N_1934);
nand U3079 (N_3079,N_1259,N_812);
or U3080 (N_3080,N_435,N_796);
xnor U3081 (N_3081,N_774,N_449);
and U3082 (N_3082,N_1205,N_487);
nand U3083 (N_3083,N_9,N_6);
and U3084 (N_3084,N_1354,N_1890);
or U3085 (N_3085,N_1717,N_1892);
or U3086 (N_3086,N_1124,N_1278);
nand U3087 (N_3087,N_1394,N_591);
and U3088 (N_3088,N_264,N_486);
nor U3089 (N_3089,N_1846,N_1220);
or U3090 (N_3090,N_1648,N_37);
nor U3091 (N_3091,N_866,N_1397);
or U3092 (N_3092,N_1273,N_456);
nand U3093 (N_3093,N_353,N_1676);
and U3094 (N_3094,N_428,N_164);
nand U3095 (N_3095,N_535,N_1237);
nor U3096 (N_3096,N_129,N_1291);
nand U3097 (N_3097,N_404,N_1067);
or U3098 (N_3098,N_392,N_1699);
nand U3099 (N_3099,N_1533,N_1493);
or U3100 (N_3100,N_579,N_1787);
xor U3101 (N_3101,N_189,N_251);
xnor U3102 (N_3102,N_181,N_732);
nor U3103 (N_3103,N_1128,N_235);
xnor U3104 (N_3104,N_1728,N_979);
nand U3105 (N_3105,N_1192,N_1099);
xnor U3106 (N_3106,N_1504,N_615);
or U3107 (N_3107,N_1836,N_1901);
nand U3108 (N_3108,N_1468,N_1727);
xnor U3109 (N_3109,N_86,N_1083);
nand U3110 (N_3110,N_1937,N_916);
or U3111 (N_3111,N_1197,N_1611);
nor U3112 (N_3112,N_682,N_107);
or U3113 (N_3113,N_840,N_711);
or U3114 (N_3114,N_109,N_549);
or U3115 (N_3115,N_377,N_1367);
and U3116 (N_3116,N_340,N_366);
nand U3117 (N_3117,N_1203,N_1536);
or U3118 (N_3118,N_307,N_647);
nor U3119 (N_3119,N_1200,N_237);
and U3120 (N_3120,N_776,N_1120);
xnor U3121 (N_3121,N_1759,N_1179);
or U3122 (N_3122,N_1611,N_1178);
nor U3123 (N_3123,N_379,N_1025);
nand U3124 (N_3124,N_1921,N_543);
xnor U3125 (N_3125,N_805,N_175);
nor U3126 (N_3126,N_1175,N_1540);
and U3127 (N_3127,N_506,N_1318);
and U3128 (N_3128,N_245,N_1065);
nor U3129 (N_3129,N_1991,N_229);
or U3130 (N_3130,N_1208,N_1974);
and U3131 (N_3131,N_1061,N_1332);
nand U3132 (N_3132,N_77,N_1906);
or U3133 (N_3133,N_1269,N_1379);
xor U3134 (N_3134,N_961,N_1920);
nand U3135 (N_3135,N_710,N_955);
nand U3136 (N_3136,N_1233,N_1953);
nand U3137 (N_3137,N_263,N_20);
nand U3138 (N_3138,N_1811,N_1563);
nand U3139 (N_3139,N_1648,N_68);
or U3140 (N_3140,N_622,N_1652);
xor U3141 (N_3141,N_1369,N_1163);
nor U3142 (N_3142,N_859,N_537);
nand U3143 (N_3143,N_1550,N_1158);
and U3144 (N_3144,N_1892,N_1425);
and U3145 (N_3145,N_1077,N_20);
nand U3146 (N_3146,N_648,N_971);
and U3147 (N_3147,N_1270,N_1278);
nand U3148 (N_3148,N_812,N_854);
and U3149 (N_3149,N_1437,N_1963);
or U3150 (N_3150,N_1431,N_428);
nor U3151 (N_3151,N_869,N_671);
nor U3152 (N_3152,N_628,N_108);
xnor U3153 (N_3153,N_136,N_586);
nand U3154 (N_3154,N_1063,N_779);
xor U3155 (N_3155,N_1068,N_344);
nor U3156 (N_3156,N_1528,N_638);
and U3157 (N_3157,N_810,N_768);
nor U3158 (N_3158,N_555,N_552);
and U3159 (N_3159,N_765,N_1204);
and U3160 (N_3160,N_201,N_1514);
or U3161 (N_3161,N_1853,N_511);
and U3162 (N_3162,N_1714,N_1552);
nor U3163 (N_3163,N_347,N_971);
xor U3164 (N_3164,N_864,N_1759);
or U3165 (N_3165,N_122,N_183);
nand U3166 (N_3166,N_1428,N_1179);
and U3167 (N_3167,N_133,N_730);
nand U3168 (N_3168,N_960,N_1649);
and U3169 (N_3169,N_1770,N_1653);
nor U3170 (N_3170,N_135,N_1563);
and U3171 (N_3171,N_903,N_124);
nor U3172 (N_3172,N_1559,N_1085);
and U3173 (N_3173,N_243,N_1919);
nand U3174 (N_3174,N_554,N_595);
and U3175 (N_3175,N_647,N_130);
nand U3176 (N_3176,N_1807,N_967);
nand U3177 (N_3177,N_734,N_1603);
and U3178 (N_3178,N_1778,N_131);
or U3179 (N_3179,N_79,N_1940);
nor U3180 (N_3180,N_36,N_1904);
and U3181 (N_3181,N_1184,N_1092);
and U3182 (N_3182,N_1749,N_1347);
nand U3183 (N_3183,N_826,N_430);
nor U3184 (N_3184,N_1831,N_1724);
xnor U3185 (N_3185,N_1638,N_1885);
xnor U3186 (N_3186,N_557,N_30);
or U3187 (N_3187,N_405,N_486);
nor U3188 (N_3188,N_1911,N_527);
or U3189 (N_3189,N_472,N_108);
xnor U3190 (N_3190,N_664,N_764);
or U3191 (N_3191,N_1344,N_1908);
xnor U3192 (N_3192,N_1577,N_1618);
or U3193 (N_3193,N_236,N_1285);
and U3194 (N_3194,N_1576,N_539);
xnor U3195 (N_3195,N_1298,N_1307);
nor U3196 (N_3196,N_257,N_684);
xnor U3197 (N_3197,N_159,N_554);
nand U3198 (N_3198,N_1746,N_753);
xnor U3199 (N_3199,N_18,N_677);
xnor U3200 (N_3200,N_1775,N_1702);
xnor U3201 (N_3201,N_1054,N_1107);
or U3202 (N_3202,N_1949,N_1247);
nor U3203 (N_3203,N_85,N_1508);
xor U3204 (N_3204,N_1771,N_539);
nor U3205 (N_3205,N_1722,N_1238);
or U3206 (N_3206,N_1601,N_124);
nor U3207 (N_3207,N_70,N_324);
and U3208 (N_3208,N_1637,N_532);
nand U3209 (N_3209,N_459,N_407);
nand U3210 (N_3210,N_1484,N_1555);
nand U3211 (N_3211,N_1056,N_241);
nor U3212 (N_3212,N_650,N_1715);
nor U3213 (N_3213,N_1718,N_207);
or U3214 (N_3214,N_156,N_1018);
nor U3215 (N_3215,N_124,N_228);
and U3216 (N_3216,N_1129,N_1650);
and U3217 (N_3217,N_1205,N_520);
nand U3218 (N_3218,N_139,N_291);
and U3219 (N_3219,N_1052,N_209);
nor U3220 (N_3220,N_532,N_58);
and U3221 (N_3221,N_1954,N_18);
xor U3222 (N_3222,N_1379,N_732);
nor U3223 (N_3223,N_1367,N_1288);
or U3224 (N_3224,N_1771,N_1431);
nor U3225 (N_3225,N_447,N_1183);
nand U3226 (N_3226,N_1627,N_993);
and U3227 (N_3227,N_116,N_181);
nand U3228 (N_3228,N_68,N_163);
and U3229 (N_3229,N_450,N_599);
nand U3230 (N_3230,N_1112,N_706);
xnor U3231 (N_3231,N_1271,N_1865);
nand U3232 (N_3232,N_288,N_618);
nor U3233 (N_3233,N_1385,N_1640);
nand U3234 (N_3234,N_1322,N_1350);
nor U3235 (N_3235,N_954,N_397);
nand U3236 (N_3236,N_213,N_1672);
nor U3237 (N_3237,N_1561,N_1224);
xor U3238 (N_3238,N_1235,N_220);
nor U3239 (N_3239,N_504,N_303);
nor U3240 (N_3240,N_1942,N_1323);
xor U3241 (N_3241,N_783,N_1135);
nor U3242 (N_3242,N_641,N_203);
nor U3243 (N_3243,N_506,N_1384);
nand U3244 (N_3244,N_764,N_1215);
xnor U3245 (N_3245,N_832,N_580);
and U3246 (N_3246,N_1932,N_169);
nor U3247 (N_3247,N_1069,N_481);
nand U3248 (N_3248,N_1423,N_1472);
or U3249 (N_3249,N_959,N_9);
nor U3250 (N_3250,N_226,N_1222);
or U3251 (N_3251,N_639,N_1316);
and U3252 (N_3252,N_809,N_165);
and U3253 (N_3253,N_1195,N_770);
nor U3254 (N_3254,N_717,N_293);
and U3255 (N_3255,N_501,N_679);
and U3256 (N_3256,N_1746,N_295);
xor U3257 (N_3257,N_1231,N_434);
xnor U3258 (N_3258,N_1622,N_54);
and U3259 (N_3259,N_1685,N_1129);
or U3260 (N_3260,N_208,N_744);
nor U3261 (N_3261,N_275,N_1495);
and U3262 (N_3262,N_1176,N_551);
or U3263 (N_3263,N_1679,N_1655);
nor U3264 (N_3264,N_24,N_1644);
nor U3265 (N_3265,N_700,N_1943);
nor U3266 (N_3266,N_117,N_1759);
and U3267 (N_3267,N_1936,N_1456);
nand U3268 (N_3268,N_1093,N_1688);
xor U3269 (N_3269,N_672,N_716);
or U3270 (N_3270,N_178,N_520);
nor U3271 (N_3271,N_1856,N_1811);
and U3272 (N_3272,N_1577,N_1025);
or U3273 (N_3273,N_1461,N_1203);
xor U3274 (N_3274,N_1508,N_1391);
nand U3275 (N_3275,N_1315,N_773);
nor U3276 (N_3276,N_1204,N_1104);
xnor U3277 (N_3277,N_466,N_1880);
and U3278 (N_3278,N_1986,N_1479);
and U3279 (N_3279,N_1885,N_1955);
or U3280 (N_3280,N_914,N_182);
nor U3281 (N_3281,N_1087,N_106);
or U3282 (N_3282,N_342,N_765);
and U3283 (N_3283,N_1776,N_374);
and U3284 (N_3284,N_509,N_389);
nand U3285 (N_3285,N_524,N_214);
xor U3286 (N_3286,N_51,N_198);
xor U3287 (N_3287,N_1933,N_478);
nand U3288 (N_3288,N_1353,N_1872);
or U3289 (N_3289,N_354,N_769);
nor U3290 (N_3290,N_1560,N_1487);
xor U3291 (N_3291,N_1430,N_839);
or U3292 (N_3292,N_1441,N_313);
xor U3293 (N_3293,N_861,N_1150);
or U3294 (N_3294,N_1252,N_1640);
nor U3295 (N_3295,N_565,N_583);
nor U3296 (N_3296,N_280,N_1240);
and U3297 (N_3297,N_1653,N_248);
or U3298 (N_3298,N_1773,N_419);
or U3299 (N_3299,N_965,N_1401);
xnor U3300 (N_3300,N_1523,N_928);
and U3301 (N_3301,N_682,N_1868);
and U3302 (N_3302,N_260,N_1025);
or U3303 (N_3303,N_952,N_483);
xnor U3304 (N_3304,N_1764,N_967);
nand U3305 (N_3305,N_965,N_1499);
or U3306 (N_3306,N_1130,N_16);
nor U3307 (N_3307,N_1666,N_1973);
or U3308 (N_3308,N_1631,N_1875);
xor U3309 (N_3309,N_294,N_539);
or U3310 (N_3310,N_1558,N_1093);
or U3311 (N_3311,N_1666,N_1141);
or U3312 (N_3312,N_536,N_237);
xor U3313 (N_3313,N_1774,N_1344);
xor U3314 (N_3314,N_218,N_1874);
nand U3315 (N_3315,N_1692,N_167);
and U3316 (N_3316,N_1427,N_1559);
nor U3317 (N_3317,N_82,N_1820);
nor U3318 (N_3318,N_499,N_1755);
or U3319 (N_3319,N_1588,N_1469);
xor U3320 (N_3320,N_515,N_1891);
nand U3321 (N_3321,N_1297,N_1625);
or U3322 (N_3322,N_1536,N_1086);
nor U3323 (N_3323,N_103,N_750);
nor U3324 (N_3324,N_1586,N_815);
nor U3325 (N_3325,N_1502,N_1084);
nor U3326 (N_3326,N_1526,N_450);
or U3327 (N_3327,N_71,N_1467);
nand U3328 (N_3328,N_1080,N_1377);
xnor U3329 (N_3329,N_546,N_1149);
xnor U3330 (N_3330,N_107,N_475);
nand U3331 (N_3331,N_1838,N_995);
nand U3332 (N_3332,N_525,N_1794);
or U3333 (N_3333,N_1460,N_1297);
or U3334 (N_3334,N_465,N_1363);
and U3335 (N_3335,N_291,N_238);
and U3336 (N_3336,N_1693,N_1276);
and U3337 (N_3337,N_912,N_1103);
and U3338 (N_3338,N_1916,N_1887);
or U3339 (N_3339,N_1763,N_507);
nor U3340 (N_3340,N_1680,N_1581);
and U3341 (N_3341,N_1728,N_1741);
xnor U3342 (N_3342,N_760,N_1010);
or U3343 (N_3343,N_687,N_596);
and U3344 (N_3344,N_1975,N_1124);
nand U3345 (N_3345,N_418,N_1087);
xnor U3346 (N_3346,N_1597,N_724);
or U3347 (N_3347,N_371,N_1117);
nor U3348 (N_3348,N_1517,N_838);
xor U3349 (N_3349,N_1987,N_708);
nand U3350 (N_3350,N_444,N_1127);
and U3351 (N_3351,N_1297,N_290);
or U3352 (N_3352,N_606,N_203);
or U3353 (N_3353,N_1185,N_1241);
xor U3354 (N_3354,N_864,N_306);
or U3355 (N_3355,N_582,N_269);
and U3356 (N_3356,N_1914,N_1370);
or U3357 (N_3357,N_917,N_762);
nand U3358 (N_3358,N_1041,N_406);
and U3359 (N_3359,N_1609,N_842);
or U3360 (N_3360,N_1236,N_1593);
nor U3361 (N_3361,N_376,N_1003);
or U3362 (N_3362,N_745,N_1612);
xor U3363 (N_3363,N_1584,N_1618);
or U3364 (N_3364,N_1608,N_1345);
and U3365 (N_3365,N_1710,N_293);
xnor U3366 (N_3366,N_801,N_1753);
and U3367 (N_3367,N_289,N_363);
nor U3368 (N_3368,N_764,N_1850);
or U3369 (N_3369,N_166,N_551);
nand U3370 (N_3370,N_1892,N_1601);
xnor U3371 (N_3371,N_1572,N_841);
nand U3372 (N_3372,N_1443,N_1387);
and U3373 (N_3373,N_1590,N_1888);
nand U3374 (N_3374,N_1322,N_1920);
or U3375 (N_3375,N_239,N_309);
nand U3376 (N_3376,N_1799,N_1920);
nor U3377 (N_3377,N_361,N_1079);
xor U3378 (N_3378,N_9,N_1200);
nor U3379 (N_3379,N_18,N_875);
and U3380 (N_3380,N_1167,N_618);
or U3381 (N_3381,N_1680,N_191);
nor U3382 (N_3382,N_1486,N_1649);
nor U3383 (N_3383,N_1680,N_438);
and U3384 (N_3384,N_1575,N_744);
nand U3385 (N_3385,N_962,N_1697);
and U3386 (N_3386,N_1525,N_1153);
nor U3387 (N_3387,N_681,N_477);
nand U3388 (N_3388,N_1019,N_1091);
nor U3389 (N_3389,N_857,N_1132);
nor U3390 (N_3390,N_1433,N_1767);
and U3391 (N_3391,N_96,N_1099);
nand U3392 (N_3392,N_11,N_176);
nor U3393 (N_3393,N_1914,N_116);
or U3394 (N_3394,N_1676,N_322);
xnor U3395 (N_3395,N_1626,N_1961);
nor U3396 (N_3396,N_1623,N_849);
xnor U3397 (N_3397,N_269,N_1010);
nor U3398 (N_3398,N_1660,N_208);
nand U3399 (N_3399,N_640,N_225);
and U3400 (N_3400,N_1702,N_390);
xnor U3401 (N_3401,N_462,N_38);
or U3402 (N_3402,N_1575,N_1595);
nand U3403 (N_3403,N_1738,N_1131);
xnor U3404 (N_3404,N_1126,N_684);
and U3405 (N_3405,N_1812,N_301);
nand U3406 (N_3406,N_1540,N_414);
or U3407 (N_3407,N_1208,N_677);
nor U3408 (N_3408,N_605,N_940);
and U3409 (N_3409,N_302,N_1572);
nor U3410 (N_3410,N_579,N_1866);
xnor U3411 (N_3411,N_913,N_133);
and U3412 (N_3412,N_531,N_1832);
nor U3413 (N_3413,N_1926,N_864);
nand U3414 (N_3414,N_1447,N_907);
nand U3415 (N_3415,N_702,N_976);
or U3416 (N_3416,N_907,N_1667);
xor U3417 (N_3417,N_226,N_340);
or U3418 (N_3418,N_1004,N_1513);
nand U3419 (N_3419,N_719,N_1911);
or U3420 (N_3420,N_1109,N_772);
and U3421 (N_3421,N_1100,N_882);
nor U3422 (N_3422,N_1522,N_1733);
or U3423 (N_3423,N_602,N_1876);
nand U3424 (N_3424,N_861,N_1815);
or U3425 (N_3425,N_1310,N_496);
nand U3426 (N_3426,N_1322,N_1223);
nand U3427 (N_3427,N_255,N_1288);
nor U3428 (N_3428,N_583,N_1023);
xor U3429 (N_3429,N_607,N_1346);
nand U3430 (N_3430,N_741,N_1544);
or U3431 (N_3431,N_1656,N_1532);
nor U3432 (N_3432,N_918,N_170);
nand U3433 (N_3433,N_772,N_262);
and U3434 (N_3434,N_309,N_1376);
or U3435 (N_3435,N_1584,N_1047);
nor U3436 (N_3436,N_319,N_331);
or U3437 (N_3437,N_971,N_778);
and U3438 (N_3438,N_1519,N_632);
xnor U3439 (N_3439,N_1721,N_1322);
xnor U3440 (N_3440,N_1837,N_549);
or U3441 (N_3441,N_647,N_855);
nand U3442 (N_3442,N_1096,N_542);
nand U3443 (N_3443,N_1468,N_1123);
and U3444 (N_3444,N_1234,N_1352);
and U3445 (N_3445,N_1247,N_717);
or U3446 (N_3446,N_992,N_215);
xor U3447 (N_3447,N_59,N_798);
nand U3448 (N_3448,N_1880,N_998);
nor U3449 (N_3449,N_547,N_387);
and U3450 (N_3450,N_357,N_906);
and U3451 (N_3451,N_341,N_997);
or U3452 (N_3452,N_1467,N_1027);
nor U3453 (N_3453,N_242,N_1632);
xnor U3454 (N_3454,N_758,N_1589);
xor U3455 (N_3455,N_1353,N_548);
nor U3456 (N_3456,N_395,N_441);
nor U3457 (N_3457,N_1241,N_479);
nor U3458 (N_3458,N_969,N_20);
or U3459 (N_3459,N_1829,N_1064);
and U3460 (N_3460,N_507,N_1470);
or U3461 (N_3461,N_360,N_440);
and U3462 (N_3462,N_1559,N_1977);
and U3463 (N_3463,N_777,N_747);
or U3464 (N_3464,N_1299,N_1484);
xnor U3465 (N_3465,N_1994,N_203);
or U3466 (N_3466,N_1342,N_1833);
nand U3467 (N_3467,N_1469,N_616);
xnor U3468 (N_3468,N_1831,N_1673);
nor U3469 (N_3469,N_1778,N_1934);
and U3470 (N_3470,N_1671,N_1172);
and U3471 (N_3471,N_44,N_1912);
and U3472 (N_3472,N_306,N_1205);
or U3473 (N_3473,N_1035,N_1299);
nand U3474 (N_3474,N_540,N_1704);
or U3475 (N_3475,N_1990,N_1561);
nor U3476 (N_3476,N_282,N_1069);
and U3477 (N_3477,N_699,N_674);
xnor U3478 (N_3478,N_1665,N_1094);
or U3479 (N_3479,N_1450,N_1760);
nor U3480 (N_3480,N_1159,N_1210);
nand U3481 (N_3481,N_1493,N_525);
xnor U3482 (N_3482,N_1991,N_1433);
nand U3483 (N_3483,N_1543,N_689);
nand U3484 (N_3484,N_53,N_1467);
xor U3485 (N_3485,N_833,N_576);
nand U3486 (N_3486,N_1051,N_882);
and U3487 (N_3487,N_1477,N_1455);
xor U3488 (N_3488,N_1246,N_1123);
or U3489 (N_3489,N_813,N_727);
and U3490 (N_3490,N_561,N_1261);
nand U3491 (N_3491,N_705,N_1112);
nor U3492 (N_3492,N_1051,N_1662);
nor U3493 (N_3493,N_145,N_207);
xor U3494 (N_3494,N_87,N_1139);
xor U3495 (N_3495,N_1046,N_1957);
or U3496 (N_3496,N_571,N_1234);
xnor U3497 (N_3497,N_83,N_351);
and U3498 (N_3498,N_829,N_214);
or U3499 (N_3499,N_529,N_1320);
and U3500 (N_3500,N_1366,N_168);
nor U3501 (N_3501,N_1116,N_276);
or U3502 (N_3502,N_1904,N_1047);
or U3503 (N_3503,N_1414,N_1723);
xnor U3504 (N_3504,N_391,N_1028);
nand U3505 (N_3505,N_1701,N_546);
and U3506 (N_3506,N_828,N_1685);
or U3507 (N_3507,N_1066,N_1157);
xor U3508 (N_3508,N_1974,N_759);
or U3509 (N_3509,N_1628,N_120);
xnor U3510 (N_3510,N_137,N_638);
nor U3511 (N_3511,N_879,N_591);
nand U3512 (N_3512,N_1889,N_929);
nor U3513 (N_3513,N_335,N_435);
xor U3514 (N_3514,N_1116,N_1130);
or U3515 (N_3515,N_1950,N_394);
xnor U3516 (N_3516,N_462,N_1222);
xor U3517 (N_3517,N_1221,N_1992);
nand U3518 (N_3518,N_1089,N_951);
or U3519 (N_3519,N_1126,N_818);
and U3520 (N_3520,N_1463,N_682);
xor U3521 (N_3521,N_508,N_1418);
and U3522 (N_3522,N_291,N_466);
or U3523 (N_3523,N_1120,N_481);
xnor U3524 (N_3524,N_1124,N_1899);
nand U3525 (N_3525,N_884,N_71);
or U3526 (N_3526,N_1804,N_185);
or U3527 (N_3527,N_1452,N_1501);
and U3528 (N_3528,N_394,N_172);
nor U3529 (N_3529,N_923,N_1963);
xnor U3530 (N_3530,N_1336,N_1541);
nand U3531 (N_3531,N_1909,N_1458);
and U3532 (N_3532,N_233,N_1203);
xor U3533 (N_3533,N_456,N_650);
nand U3534 (N_3534,N_222,N_1163);
or U3535 (N_3535,N_384,N_1652);
nor U3536 (N_3536,N_279,N_118);
nor U3537 (N_3537,N_1332,N_832);
nand U3538 (N_3538,N_917,N_988);
and U3539 (N_3539,N_31,N_627);
and U3540 (N_3540,N_1350,N_1172);
nand U3541 (N_3541,N_1306,N_1093);
nand U3542 (N_3542,N_1081,N_1836);
and U3543 (N_3543,N_1561,N_941);
and U3544 (N_3544,N_1356,N_1488);
nand U3545 (N_3545,N_1809,N_1550);
or U3546 (N_3546,N_221,N_653);
xor U3547 (N_3547,N_1073,N_1145);
xor U3548 (N_3548,N_1809,N_504);
or U3549 (N_3549,N_1518,N_1187);
nor U3550 (N_3550,N_428,N_1498);
xor U3551 (N_3551,N_263,N_650);
and U3552 (N_3552,N_1121,N_1792);
and U3553 (N_3553,N_236,N_940);
nor U3554 (N_3554,N_234,N_985);
and U3555 (N_3555,N_1539,N_159);
nor U3556 (N_3556,N_1408,N_1714);
nor U3557 (N_3557,N_1096,N_1487);
and U3558 (N_3558,N_1296,N_1056);
nand U3559 (N_3559,N_1110,N_177);
xnor U3560 (N_3560,N_835,N_1451);
or U3561 (N_3561,N_120,N_965);
xnor U3562 (N_3562,N_1956,N_1768);
or U3563 (N_3563,N_1318,N_1822);
and U3564 (N_3564,N_179,N_1118);
nor U3565 (N_3565,N_38,N_253);
and U3566 (N_3566,N_311,N_1742);
or U3567 (N_3567,N_1276,N_304);
and U3568 (N_3568,N_1556,N_148);
nand U3569 (N_3569,N_1631,N_5);
and U3570 (N_3570,N_55,N_875);
nand U3571 (N_3571,N_934,N_996);
nand U3572 (N_3572,N_1387,N_223);
nand U3573 (N_3573,N_1332,N_378);
nor U3574 (N_3574,N_74,N_1094);
nand U3575 (N_3575,N_1066,N_1258);
nor U3576 (N_3576,N_248,N_423);
nand U3577 (N_3577,N_1881,N_1172);
or U3578 (N_3578,N_1815,N_1561);
or U3579 (N_3579,N_1908,N_1569);
or U3580 (N_3580,N_1270,N_844);
and U3581 (N_3581,N_1329,N_255);
and U3582 (N_3582,N_1726,N_1220);
nand U3583 (N_3583,N_552,N_102);
and U3584 (N_3584,N_1714,N_76);
and U3585 (N_3585,N_126,N_712);
and U3586 (N_3586,N_741,N_411);
or U3587 (N_3587,N_490,N_830);
and U3588 (N_3588,N_1178,N_77);
xor U3589 (N_3589,N_1701,N_424);
nand U3590 (N_3590,N_1927,N_913);
and U3591 (N_3591,N_601,N_1483);
or U3592 (N_3592,N_1701,N_374);
nor U3593 (N_3593,N_1538,N_1764);
nand U3594 (N_3594,N_1847,N_167);
xor U3595 (N_3595,N_1590,N_748);
and U3596 (N_3596,N_481,N_1390);
or U3597 (N_3597,N_245,N_1020);
nand U3598 (N_3598,N_1200,N_979);
and U3599 (N_3599,N_1129,N_26);
nand U3600 (N_3600,N_1289,N_1942);
nand U3601 (N_3601,N_386,N_1963);
and U3602 (N_3602,N_1429,N_670);
xnor U3603 (N_3603,N_1172,N_1189);
nand U3604 (N_3604,N_1727,N_31);
and U3605 (N_3605,N_1719,N_1671);
or U3606 (N_3606,N_1898,N_675);
nand U3607 (N_3607,N_504,N_1517);
or U3608 (N_3608,N_871,N_210);
and U3609 (N_3609,N_1177,N_1856);
xnor U3610 (N_3610,N_435,N_893);
nor U3611 (N_3611,N_914,N_1614);
nand U3612 (N_3612,N_632,N_190);
and U3613 (N_3613,N_915,N_322);
nand U3614 (N_3614,N_1680,N_597);
xnor U3615 (N_3615,N_1224,N_1763);
and U3616 (N_3616,N_1005,N_839);
xor U3617 (N_3617,N_1320,N_753);
xnor U3618 (N_3618,N_787,N_1106);
xor U3619 (N_3619,N_97,N_827);
nor U3620 (N_3620,N_645,N_878);
and U3621 (N_3621,N_1366,N_1966);
and U3622 (N_3622,N_557,N_1857);
and U3623 (N_3623,N_564,N_948);
nor U3624 (N_3624,N_774,N_1258);
and U3625 (N_3625,N_44,N_528);
nor U3626 (N_3626,N_1994,N_1823);
nand U3627 (N_3627,N_865,N_207);
xnor U3628 (N_3628,N_227,N_1035);
xor U3629 (N_3629,N_1094,N_541);
nand U3630 (N_3630,N_89,N_865);
and U3631 (N_3631,N_1111,N_1259);
and U3632 (N_3632,N_600,N_1498);
or U3633 (N_3633,N_772,N_1716);
nor U3634 (N_3634,N_668,N_1196);
nor U3635 (N_3635,N_1342,N_1446);
and U3636 (N_3636,N_1912,N_716);
nor U3637 (N_3637,N_1006,N_743);
nor U3638 (N_3638,N_361,N_248);
xnor U3639 (N_3639,N_1784,N_1027);
and U3640 (N_3640,N_435,N_1378);
and U3641 (N_3641,N_1486,N_1615);
and U3642 (N_3642,N_167,N_1755);
xor U3643 (N_3643,N_889,N_1634);
or U3644 (N_3644,N_1180,N_808);
nor U3645 (N_3645,N_136,N_420);
and U3646 (N_3646,N_131,N_500);
and U3647 (N_3647,N_1378,N_1725);
and U3648 (N_3648,N_1951,N_1133);
nor U3649 (N_3649,N_79,N_796);
nand U3650 (N_3650,N_555,N_1457);
or U3651 (N_3651,N_751,N_186);
or U3652 (N_3652,N_704,N_1238);
nor U3653 (N_3653,N_556,N_325);
xnor U3654 (N_3654,N_1791,N_661);
or U3655 (N_3655,N_32,N_582);
or U3656 (N_3656,N_1922,N_1036);
xnor U3657 (N_3657,N_1622,N_604);
and U3658 (N_3658,N_986,N_201);
xor U3659 (N_3659,N_1405,N_339);
nor U3660 (N_3660,N_123,N_1972);
xnor U3661 (N_3661,N_787,N_1802);
xor U3662 (N_3662,N_476,N_3);
nor U3663 (N_3663,N_512,N_949);
nand U3664 (N_3664,N_1514,N_681);
nor U3665 (N_3665,N_789,N_1505);
nand U3666 (N_3666,N_1588,N_71);
xor U3667 (N_3667,N_869,N_1430);
nor U3668 (N_3668,N_785,N_1744);
nand U3669 (N_3669,N_961,N_1297);
and U3670 (N_3670,N_656,N_1373);
or U3671 (N_3671,N_1830,N_1293);
nor U3672 (N_3672,N_106,N_105);
nor U3673 (N_3673,N_1958,N_187);
or U3674 (N_3674,N_574,N_1032);
xor U3675 (N_3675,N_1114,N_544);
xnor U3676 (N_3676,N_1785,N_788);
nor U3677 (N_3677,N_1029,N_787);
nor U3678 (N_3678,N_1981,N_1410);
and U3679 (N_3679,N_1630,N_183);
or U3680 (N_3680,N_1099,N_750);
xnor U3681 (N_3681,N_243,N_1580);
nor U3682 (N_3682,N_577,N_1782);
nor U3683 (N_3683,N_1040,N_764);
nor U3684 (N_3684,N_389,N_254);
xor U3685 (N_3685,N_1525,N_1451);
and U3686 (N_3686,N_1629,N_1780);
or U3687 (N_3687,N_86,N_969);
xor U3688 (N_3688,N_58,N_1763);
or U3689 (N_3689,N_131,N_1227);
xnor U3690 (N_3690,N_430,N_1669);
nor U3691 (N_3691,N_1440,N_1694);
nand U3692 (N_3692,N_1926,N_1892);
nand U3693 (N_3693,N_544,N_1789);
xnor U3694 (N_3694,N_949,N_1478);
nor U3695 (N_3695,N_1471,N_1361);
nor U3696 (N_3696,N_926,N_720);
nor U3697 (N_3697,N_1131,N_1446);
nor U3698 (N_3698,N_1654,N_978);
or U3699 (N_3699,N_587,N_966);
or U3700 (N_3700,N_1795,N_939);
nor U3701 (N_3701,N_419,N_1745);
nor U3702 (N_3702,N_1295,N_539);
and U3703 (N_3703,N_813,N_868);
and U3704 (N_3704,N_523,N_179);
nand U3705 (N_3705,N_311,N_1663);
nand U3706 (N_3706,N_1631,N_510);
or U3707 (N_3707,N_623,N_1111);
nand U3708 (N_3708,N_1586,N_155);
xor U3709 (N_3709,N_1421,N_147);
nand U3710 (N_3710,N_931,N_721);
or U3711 (N_3711,N_1617,N_31);
and U3712 (N_3712,N_1741,N_1944);
nand U3713 (N_3713,N_1828,N_1380);
nand U3714 (N_3714,N_1599,N_374);
nor U3715 (N_3715,N_854,N_361);
and U3716 (N_3716,N_533,N_1976);
nand U3717 (N_3717,N_468,N_1502);
nand U3718 (N_3718,N_294,N_1489);
nand U3719 (N_3719,N_1271,N_1200);
and U3720 (N_3720,N_100,N_223);
nand U3721 (N_3721,N_982,N_1339);
and U3722 (N_3722,N_1991,N_1746);
xnor U3723 (N_3723,N_471,N_254);
nor U3724 (N_3724,N_691,N_1998);
nor U3725 (N_3725,N_304,N_1219);
nand U3726 (N_3726,N_357,N_657);
nor U3727 (N_3727,N_76,N_1179);
nand U3728 (N_3728,N_1454,N_1094);
nor U3729 (N_3729,N_401,N_1462);
xnor U3730 (N_3730,N_624,N_359);
nand U3731 (N_3731,N_664,N_1877);
nand U3732 (N_3732,N_171,N_286);
or U3733 (N_3733,N_608,N_1075);
nand U3734 (N_3734,N_1303,N_1027);
nand U3735 (N_3735,N_683,N_763);
xnor U3736 (N_3736,N_1068,N_13);
and U3737 (N_3737,N_471,N_935);
nor U3738 (N_3738,N_1888,N_1865);
nand U3739 (N_3739,N_1262,N_1785);
nor U3740 (N_3740,N_1369,N_14);
nor U3741 (N_3741,N_1614,N_1271);
and U3742 (N_3742,N_304,N_1322);
xor U3743 (N_3743,N_1612,N_1403);
and U3744 (N_3744,N_1639,N_1804);
or U3745 (N_3745,N_174,N_278);
and U3746 (N_3746,N_1001,N_348);
xnor U3747 (N_3747,N_267,N_936);
nand U3748 (N_3748,N_270,N_1282);
or U3749 (N_3749,N_101,N_488);
nor U3750 (N_3750,N_527,N_788);
xor U3751 (N_3751,N_194,N_330);
nand U3752 (N_3752,N_1359,N_1247);
and U3753 (N_3753,N_841,N_1079);
nor U3754 (N_3754,N_857,N_1797);
nand U3755 (N_3755,N_282,N_331);
nor U3756 (N_3756,N_1261,N_491);
nor U3757 (N_3757,N_615,N_261);
nor U3758 (N_3758,N_1619,N_1513);
xor U3759 (N_3759,N_1688,N_1756);
or U3760 (N_3760,N_1159,N_473);
nor U3761 (N_3761,N_774,N_1033);
xnor U3762 (N_3762,N_1721,N_1282);
nand U3763 (N_3763,N_282,N_1204);
or U3764 (N_3764,N_1158,N_351);
and U3765 (N_3765,N_594,N_1687);
nand U3766 (N_3766,N_1386,N_1011);
or U3767 (N_3767,N_478,N_1241);
nand U3768 (N_3768,N_375,N_646);
and U3769 (N_3769,N_397,N_1736);
nand U3770 (N_3770,N_1751,N_226);
xor U3771 (N_3771,N_561,N_822);
and U3772 (N_3772,N_1168,N_1716);
and U3773 (N_3773,N_1075,N_1847);
or U3774 (N_3774,N_266,N_491);
xor U3775 (N_3775,N_1987,N_904);
xnor U3776 (N_3776,N_390,N_312);
nor U3777 (N_3777,N_149,N_1222);
and U3778 (N_3778,N_1989,N_1980);
xor U3779 (N_3779,N_838,N_963);
xor U3780 (N_3780,N_1849,N_1184);
and U3781 (N_3781,N_1109,N_706);
or U3782 (N_3782,N_1266,N_800);
and U3783 (N_3783,N_426,N_1838);
and U3784 (N_3784,N_1248,N_183);
nand U3785 (N_3785,N_877,N_1833);
xnor U3786 (N_3786,N_1687,N_1667);
nor U3787 (N_3787,N_989,N_694);
and U3788 (N_3788,N_312,N_838);
nand U3789 (N_3789,N_1643,N_1306);
or U3790 (N_3790,N_397,N_1304);
xor U3791 (N_3791,N_1837,N_1122);
or U3792 (N_3792,N_640,N_652);
nor U3793 (N_3793,N_354,N_621);
xor U3794 (N_3794,N_287,N_1790);
and U3795 (N_3795,N_540,N_1745);
xor U3796 (N_3796,N_38,N_1919);
xor U3797 (N_3797,N_1351,N_605);
nand U3798 (N_3798,N_1484,N_521);
nor U3799 (N_3799,N_1982,N_1588);
nor U3800 (N_3800,N_223,N_1048);
nor U3801 (N_3801,N_703,N_1384);
nor U3802 (N_3802,N_1701,N_1592);
xnor U3803 (N_3803,N_1197,N_335);
xor U3804 (N_3804,N_938,N_77);
xor U3805 (N_3805,N_1164,N_404);
nor U3806 (N_3806,N_1767,N_1892);
and U3807 (N_3807,N_890,N_1516);
and U3808 (N_3808,N_1873,N_1024);
xor U3809 (N_3809,N_1734,N_413);
xnor U3810 (N_3810,N_949,N_457);
and U3811 (N_3811,N_53,N_1816);
nor U3812 (N_3812,N_1161,N_147);
nor U3813 (N_3813,N_1063,N_436);
xnor U3814 (N_3814,N_609,N_582);
or U3815 (N_3815,N_101,N_1079);
xnor U3816 (N_3816,N_1254,N_1955);
and U3817 (N_3817,N_145,N_1122);
nor U3818 (N_3818,N_758,N_1002);
and U3819 (N_3819,N_1555,N_426);
or U3820 (N_3820,N_293,N_1854);
nor U3821 (N_3821,N_439,N_1546);
and U3822 (N_3822,N_1051,N_1546);
xnor U3823 (N_3823,N_1220,N_1008);
xor U3824 (N_3824,N_1495,N_1772);
nand U3825 (N_3825,N_1534,N_1542);
xnor U3826 (N_3826,N_1021,N_1989);
or U3827 (N_3827,N_174,N_731);
and U3828 (N_3828,N_190,N_1863);
or U3829 (N_3829,N_1998,N_977);
nand U3830 (N_3830,N_1269,N_1795);
or U3831 (N_3831,N_270,N_37);
nand U3832 (N_3832,N_1699,N_1059);
nor U3833 (N_3833,N_117,N_1640);
or U3834 (N_3834,N_1981,N_399);
nand U3835 (N_3835,N_852,N_1878);
xor U3836 (N_3836,N_724,N_1155);
xnor U3837 (N_3837,N_52,N_725);
xor U3838 (N_3838,N_304,N_359);
and U3839 (N_3839,N_1765,N_594);
nor U3840 (N_3840,N_1638,N_1144);
nand U3841 (N_3841,N_71,N_1460);
or U3842 (N_3842,N_1049,N_142);
xnor U3843 (N_3843,N_755,N_242);
xnor U3844 (N_3844,N_1135,N_129);
and U3845 (N_3845,N_1040,N_1556);
nand U3846 (N_3846,N_1708,N_114);
nand U3847 (N_3847,N_185,N_176);
nor U3848 (N_3848,N_1277,N_460);
or U3849 (N_3849,N_1378,N_1823);
and U3850 (N_3850,N_592,N_578);
nand U3851 (N_3851,N_1259,N_1017);
and U3852 (N_3852,N_163,N_1331);
nand U3853 (N_3853,N_455,N_1758);
and U3854 (N_3854,N_1771,N_1641);
nand U3855 (N_3855,N_1199,N_850);
xor U3856 (N_3856,N_1945,N_158);
nor U3857 (N_3857,N_243,N_152);
nand U3858 (N_3858,N_75,N_1124);
nand U3859 (N_3859,N_536,N_451);
xnor U3860 (N_3860,N_1082,N_463);
and U3861 (N_3861,N_131,N_1884);
nand U3862 (N_3862,N_234,N_75);
xnor U3863 (N_3863,N_1008,N_8);
xnor U3864 (N_3864,N_181,N_103);
nand U3865 (N_3865,N_1698,N_1079);
xnor U3866 (N_3866,N_1287,N_535);
and U3867 (N_3867,N_1163,N_1672);
and U3868 (N_3868,N_484,N_1465);
or U3869 (N_3869,N_634,N_932);
and U3870 (N_3870,N_1372,N_1071);
nor U3871 (N_3871,N_626,N_585);
and U3872 (N_3872,N_911,N_1843);
or U3873 (N_3873,N_1406,N_807);
or U3874 (N_3874,N_954,N_1357);
or U3875 (N_3875,N_17,N_92);
nor U3876 (N_3876,N_1496,N_1604);
nand U3877 (N_3877,N_200,N_1897);
xnor U3878 (N_3878,N_1577,N_29);
nor U3879 (N_3879,N_1794,N_793);
nand U3880 (N_3880,N_41,N_1582);
nor U3881 (N_3881,N_1672,N_1288);
and U3882 (N_3882,N_822,N_396);
xnor U3883 (N_3883,N_405,N_1268);
and U3884 (N_3884,N_750,N_218);
nor U3885 (N_3885,N_1486,N_1733);
nor U3886 (N_3886,N_1081,N_809);
nand U3887 (N_3887,N_1493,N_26);
nor U3888 (N_3888,N_1625,N_1224);
xnor U3889 (N_3889,N_1177,N_48);
xnor U3890 (N_3890,N_1176,N_937);
nand U3891 (N_3891,N_1604,N_1790);
nor U3892 (N_3892,N_1634,N_1547);
or U3893 (N_3893,N_1722,N_1430);
and U3894 (N_3894,N_1052,N_1421);
nand U3895 (N_3895,N_1087,N_1105);
or U3896 (N_3896,N_489,N_1940);
nand U3897 (N_3897,N_1985,N_1905);
nor U3898 (N_3898,N_370,N_706);
xor U3899 (N_3899,N_964,N_1748);
xor U3900 (N_3900,N_1924,N_901);
nand U3901 (N_3901,N_1245,N_1262);
nand U3902 (N_3902,N_1619,N_844);
nor U3903 (N_3903,N_1334,N_1273);
nor U3904 (N_3904,N_1118,N_586);
nor U3905 (N_3905,N_140,N_1387);
or U3906 (N_3906,N_305,N_545);
and U3907 (N_3907,N_1616,N_1768);
or U3908 (N_3908,N_1508,N_1735);
xor U3909 (N_3909,N_1093,N_1414);
nor U3910 (N_3910,N_1007,N_1847);
xor U3911 (N_3911,N_759,N_193);
or U3912 (N_3912,N_326,N_1969);
nand U3913 (N_3913,N_741,N_325);
and U3914 (N_3914,N_1794,N_1835);
xor U3915 (N_3915,N_1459,N_1309);
nand U3916 (N_3916,N_1909,N_1912);
nor U3917 (N_3917,N_703,N_1859);
and U3918 (N_3918,N_1491,N_1546);
nor U3919 (N_3919,N_827,N_1079);
nand U3920 (N_3920,N_537,N_17);
xor U3921 (N_3921,N_735,N_1405);
nor U3922 (N_3922,N_1950,N_1518);
or U3923 (N_3923,N_1866,N_1563);
nand U3924 (N_3924,N_1554,N_1659);
and U3925 (N_3925,N_372,N_1408);
nor U3926 (N_3926,N_1609,N_1282);
nand U3927 (N_3927,N_1110,N_449);
nand U3928 (N_3928,N_1796,N_1237);
nand U3929 (N_3929,N_1901,N_4);
xor U3930 (N_3930,N_1750,N_1140);
xor U3931 (N_3931,N_1381,N_631);
nand U3932 (N_3932,N_277,N_1804);
nor U3933 (N_3933,N_1183,N_1070);
nand U3934 (N_3934,N_1326,N_903);
and U3935 (N_3935,N_1164,N_1035);
xor U3936 (N_3936,N_1569,N_13);
nor U3937 (N_3937,N_924,N_23);
xnor U3938 (N_3938,N_30,N_990);
nor U3939 (N_3939,N_1677,N_1992);
and U3940 (N_3940,N_1993,N_1480);
or U3941 (N_3941,N_684,N_1774);
nor U3942 (N_3942,N_1892,N_1598);
nand U3943 (N_3943,N_1005,N_149);
nand U3944 (N_3944,N_1344,N_1193);
nand U3945 (N_3945,N_220,N_1099);
and U3946 (N_3946,N_1882,N_1951);
xor U3947 (N_3947,N_667,N_1522);
nor U3948 (N_3948,N_1635,N_1424);
xnor U3949 (N_3949,N_1484,N_1850);
or U3950 (N_3950,N_1207,N_1554);
nor U3951 (N_3951,N_1516,N_337);
nand U3952 (N_3952,N_1134,N_695);
nor U3953 (N_3953,N_1791,N_1921);
or U3954 (N_3954,N_801,N_1439);
and U3955 (N_3955,N_1144,N_1186);
and U3956 (N_3956,N_974,N_351);
nor U3957 (N_3957,N_976,N_71);
or U3958 (N_3958,N_456,N_186);
nand U3959 (N_3959,N_1909,N_94);
nand U3960 (N_3960,N_1142,N_590);
nand U3961 (N_3961,N_1218,N_549);
nand U3962 (N_3962,N_1117,N_498);
and U3963 (N_3963,N_811,N_729);
nand U3964 (N_3964,N_25,N_662);
nand U3965 (N_3965,N_930,N_79);
nor U3966 (N_3966,N_230,N_1497);
nor U3967 (N_3967,N_293,N_1297);
and U3968 (N_3968,N_863,N_1900);
xor U3969 (N_3969,N_618,N_598);
nand U3970 (N_3970,N_40,N_1918);
and U3971 (N_3971,N_1529,N_943);
xnor U3972 (N_3972,N_870,N_236);
or U3973 (N_3973,N_287,N_1370);
or U3974 (N_3974,N_1180,N_929);
xor U3975 (N_3975,N_883,N_1598);
and U3976 (N_3976,N_527,N_1753);
nor U3977 (N_3977,N_714,N_963);
xor U3978 (N_3978,N_992,N_862);
and U3979 (N_3979,N_1186,N_1319);
and U3980 (N_3980,N_5,N_1166);
xnor U3981 (N_3981,N_23,N_958);
xnor U3982 (N_3982,N_1280,N_1692);
and U3983 (N_3983,N_1181,N_462);
or U3984 (N_3984,N_54,N_1432);
nor U3985 (N_3985,N_1517,N_1452);
nor U3986 (N_3986,N_781,N_1622);
xnor U3987 (N_3987,N_698,N_860);
or U3988 (N_3988,N_698,N_1034);
nand U3989 (N_3989,N_891,N_1222);
nand U3990 (N_3990,N_1118,N_1225);
xor U3991 (N_3991,N_369,N_324);
nor U3992 (N_3992,N_1093,N_1644);
or U3993 (N_3993,N_1845,N_894);
and U3994 (N_3994,N_11,N_1062);
nand U3995 (N_3995,N_1140,N_625);
nor U3996 (N_3996,N_869,N_1220);
xnor U3997 (N_3997,N_1441,N_1343);
nand U3998 (N_3998,N_1123,N_442);
or U3999 (N_3999,N_155,N_784);
nor U4000 (N_4000,N_3724,N_3825);
nor U4001 (N_4001,N_2994,N_3135);
or U4002 (N_4002,N_3469,N_3874);
nand U4003 (N_4003,N_3915,N_2169);
or U4004 (N_4004,N_3523,N_2409);
and U4005 (N_4005,N_2864,N_2332);
xor U4006 (N_4006,N_2513,N_3981);
or U4007 (N_4007,N_2254,N_3948);
nand U4008 (N_4008,N_2711,N_3835);
nand U4009 (N_4009,N_2860,N_3176);
nor U4010 (N_4010,N_3892,N_2760);
xnor U4011 (N_4011,N_3195,N_2003);
and U4012 (N_4012,N_3620,N_3403);
and U4013 (N_4013,N_3569,N_3732);
xnor U4014 (N_4014,N_2488,N_2142);
nor U4015 (N_4015,N_2316,N_3170);
or U4016 (N_4016,N_3952,N_2081);
nand U4017 (N_4017,N_2080,N_3198);
xnor U4018 (N_4018,N_2649,N_2404);
or U4019 (N_4019,N_3386,N_3010);
nor U4020 (N_4020,N_3248,N_2917);
and U4021 (N_4021,N_3986,N_2295);
nor U4022 (N_4022,N_2782,N_2951);
or U4023 (N_4023,N_2174,N_2021);
nand U4024 (N_4024,N_2212,N_3687);
and U4025 (N_4025,N_2996,N_3039);
or U4026 (N_4026,N_3896,N_3490);
xnor U4027 (N_4027,N_2894,N_2798);
xor U4028 (N_4028,N_3739,N_3211);
nor U4029 (N_4029,N_3029,N_3435);
or U4030 (N_4030,N_2286,N_3798);
xnor U4031 (N_4031,N_2669,N_2294);
nor U4032 (N_4032,N_3373,N_3617);
nor U4033 (N_4033,N_2434,N_2065);
xnor U4034 (N_4034,N_2334,N_2412);
xor U4035 (N_4035,N_3224,N_2333);
nand U4036 (N_4036,N_2886,N_2852);
and U4037 (N_4037,N_3820,N_3559);
or U4038 (N_4038,N_2448,N_3396);
nand U4039 (N_4039,N_3872,N_3974);
or U4040 (N_4040,N_3716,N_2125);
xor U4041 (N_4041,N_3991,N_2561);
nand U4042 (N_4042,N_3249,N_2878);
and U4043 (N_4043,N_2024,N_2238);
xor U4044 (N_4044,N_2571,N_2490);
nor U4045 (N_4045,N_3429,N_2050);
and U4046 (N_4046,N_2223,N_2370);
or U4047 (N_4047,N_3661,N_2030);
or U4048 (N_4048,N_2397,N_3286);
xnor U4049 (N_4049,N_2704,N_2202);
nand U4050 (N_4050,N_3810,N_3444);
and U4051 (N_4051,N_2845,N_3426);
nand U4052 (N_4052,N_2098,N_3281);
nand U4053 (N_4053,N_3893,N_3168);
and U4054 (N_4054,N_2369,N_2350);
nand U4055 (N_4055,N_2918,N_2361);
nor U4056 (N_4056,N_2981,N_2577);
nor U4057 (N_4057,N_3078,N_2725);
nor U4058 (N_4058,N_3901,N_2703);
nand U4059 (N_4059,N_3508,N_2411);
nand U4060 (N_4060,N_3236,N_3936);
nor U4061 (N_4061,N_3314,N_2367);
nor U4062 (N_4062,N_3899,N_3301);
and U4063 (N_4063,N_2670,N_2763);
or U4064 (N_4064,N_2802,N_2803);
nand U4065 (N_4065,N_2797,N_3250);
or U4066 (N_4066,N_2259,N_2118);
nand U4067 (N_4067,N_2642,N_2336);
nor U4068 (N_4068,N_2041,N_2237);
and U4069 (N_4069,N_3399,N_2129);
nor U4070 (N_4070,N_2667,N_3088);
and U4071 (N_4071,N_2427,N_2534);
nor U4072 (N_4072,N_3514,N_2780);
nor U4073 (N_4073,N_3621,N_3196);
or U4074 (N_4074,N_2558,N_3934);
or U4075 (N_4075,N_2884,N_2476);
nor U4076 (N_4076,N_2074,N_2487);
xnor U4077 (N_4077,N_2430,N_2728);
xnor U4078 (N_4078,N_2993,N_2665);
nor U4079 (N_4079,N_3594,N_2340);
and U4080 (N_4080,N_3863,N_2343);
or U4081 (N_4081,N_2468,N_3200);
nor U4082 (N_4082,N_3162,N_3031);
or U4083 (N_4083,N_2550,N_3455);
xnor U4084 (N_4084,N_2700,N_3417);
or U4085 (N_4085,N_2281,N_2058);
nand U4086 (N_4086,N_2748,N_2541);
xor U4087 (N_4087,N_2114,N_3876);
or U4088 (N_4088,N_2262,N_3853);
xor U4089 (N_4089,N_3292,N_2222);
or U4090 (N_4090,N_3273,N_2651);
or U4091 (N_4091,N_3451,N_3146);
or U4092 (N_4092,N_2140,N_2526);
nor U4093 (N_4093,N_3040,N_2495);
nand U4094 (N_4094,N_3173,N_2616);
xnor U4095 (N_4095,N_3919,N_3751);
xnor U4096 (N_4096,N_2473,N_3930);
nor U4097 (N_4097,N_3808,N_3885);
xnor U4098 (N_4098,N_3027,N_3870);
and U4099 (N_4099,N_2239,N_3718);
and U4100 (N_4100,N_3118,N_3125);
nand U4101 (N_4101,N_2516,N_3165);
and U4102 (N_4102,N_2750,N_2233);
nand U4103 (N_4103,N_2127,N_3091);
nand U4104 (N_4104,N_3487,N_2761);
nand U4105 (N_4105,N_3231,N_2005);
xor U4106 (N_4106,N_3365,N_3954);
or U4107 (N_4107,N_2596,N_3655);
xnor U4108 (N_4108,N_3374,N_2392);
or U4109 (N_4109,N_2927,N_3436);
nor U4110 (N_4110,N_3616,N_2979);
xnor U4111 (N_4111,N_2063,N_2055);
and U4112 (N_4112,N_2292,N_2889);
and U4113 (N_4113,N_2199,N_2554);
nor U4114 (N_4114,N_2868,N_2958);
nor U4115 (N_4115,N_2315,N_3245);
nand U4116 (N_4116,N_2244,N_3615);
nor U4117 (N_4117,N_2668,N_3159);
or U4118 (N_4118,N_2584,N_3833);
xor U4119 (N_4119,N_2814,N_2829);
or U4120 (N_4120,N_3153,N_3675);
and U4121 (N_4121,N_2610,N_3836);
nand U4122 (N_4122,N_3580,N_3511);
nand U4123 (N_4123,N_2120,N_3440);
nor U4124 (N_4124,N_3058,N_2091);
and U4125 (N_4125,N_2141,N_2349);
nand U4126 (N_4126,N_3680,N_3345);
nand U4127 (N_4127,N_2085,N_3821);
nand U4128 (N_4128,N_3787,N_3096);
xor U4129 (N_4129,N_3119,N_2679);
nor U4130 (N_4130,N_2047,N_2335);
and U4131 (N_4131,N_3271,N_3395);
nor U4132 (N_4132,N_2973,N_3461);
and U4133 (N_4133,N_2096,N_3834);
and U4134 (N_4134,N_2329,N_3762);
xnor U4135 (N_4135,N_2776,N_2337);
nand U4136 (N_4136,N_2092,N_2539);
nor U4137 (N_4137,N_2301,N_2460);
nor U4138 (N_4138,N_3638,N_2304);
nor U4139 (N_4139,N_3938,N_2756);
or U4140 (N_4140,N_2614,N_2822);
nor U4141 (N_4141,N_2842,N_3847);
xor U4142 (N_4142,N_2194,N_2529);
nor U4143 (N_4143,N_2611,N_3969);
xor U4144 (N_4144,N_2263,N_2471);
nor U4145 (N_4145,N_3804,N_2276);
nand U4146 (N_4146,N_3139,N_3849);
and U4147 (N_4147,N_3012,N_2699);
xor U4148 (N_4148,N_3987,N_3026);
nand U4149 (N_4149,N_3341,N_3698);
xor U4150 (N_4150,N_2248,N_3375);
nor U4151 (N_4151,N_2483,N_2546);
and U4152 (N_4152,N_3690,N_3607);
or U4153 (N_4153,N_3629,N_2201);
nand U4154 (N_4154,N_3203,N_2481);
nand U4155 (N_4155,N_2597,N_3439);
and U4156 (N_4156,N_3356,N_3920);
and U4157 (N_4157,N_2772,N_2514);
nand U4158 (N_4158,N_3121,N_3912);
nor U4159 (N_4159,N_3117,N_3667);
nand U4160 (N_4160,N_3316,N_3729);
or U4161 (N_4161,N_2582,N_3209);
nor U4162 (N_4162,N_3644,N_2119);
xnor U4163 (N_4163,N_2873,N_2454);
nand U4164 (N_4164,N_3238,N_3421);
or U4165 (N_4165,N_3926,N_3388);
or U4166 (N_4166,N_3343,N_2870);
nor U4167 (N_4167,N_2923,N_2877);
xnor U4168 (N_4168,N_2757,N_2507);
or U4169 (N_4169,N_3054,N_3895);
xnor U4170 (N_4170,N_2737,N_3784);
xnor U4171 (N_4171,N_3643,N_2986);
and U4172 (N_4172,N_3958,N_2988);
and U4173 (N_4173,N_3537,N_2089);
nand U4174 (N_4174,N_3366,N_3449);
nand U4175 (N_4175,N_3811,N_3144);
and U4176 (N_4176,N_3087,N_3550);
or U4177 (N_4177,N_3637,N_3601);
xnor U4178 (N_4178,N_2817,N_2419);
nand U4179 (N_4179,N_2104,N_2648);
nor U4180 (N_4180,N_2061,N_3014);
nand U4181 (N_4181,N_2265,N_3297);
nor U4182 (N_4182,N_2250,N_3325);
nor U4183 (N_4183,N_2339,N_3190);
xnor U4184 (N_4184,N_3060,N_3664);
and U4185 (N_4185,N_3829,N_3113);
nand U4186 (N_4186,N_3864,N_2779);
and U4187 (N_4187,N_3504,N_3480);
or U4188 (N_4188,N_2804,N_2941);
and U4189 (N_4189,N_3855,N_3393);
or U4190 (N_4190,N_2747,N_3112);
xor U4191 (N_4191,N_3351,N_3788);
and U4192 (N_4192,N_3315,N_2173);
and U4193 (N_4193,N_2245,N_2026);
nand U4194 (N_4194,N_3364,N_2903);
nand U4195 (N_4195,N_2307,N_3790);
xnor U4196 (N_4196,N_3069,N_2338);
or U4197 (N_4197,N_2390,N_3433);
nand U4198 (N_4198,N_3673,N_3080);
xnor U4199 (N_4199,N_2135,N_2207);
nor U4200 (N_4200,N_2844,N_3130);
and U4201 (N_4201,N_3897,N_2847);
nor U4202 (N_4202,N_3319,N_2686);
nand U4203 (N_4203,N_3984,N_3579);
xor U4204 (N_4204,N_2759,N_3323);
nand U4205 (N_4205,N_2948,N_3921);
xnor U4206 (N_4206,N_3856,N_2474);
xnor U4207 (N_4207,N_3081,N_3858);
nor U4208 (N_4208,N_2498,N_2708);
or U4209 (N_4209,N_3558,N_2579);
xnor U4210 (N_4210,N_2676,N_2684);
and U4211 (N_4211,N_2151,N_2874);
and U4212 (N_4212,N_2892,N_3285);
and U4213 (N_4213,N_2690,N_2106);
nor U4214 (N_4214,N_2808,N_3419);
nor U4215 (N_4215,N_2060,N_3941);
and U4216 (N_4216,N_3799,N_3838);
nand U4217 (N_4217,N_2306,N_3484);
nand U4218 (N_4218,N_2843,N_3172);
nand U4219 (N_4219,N_2240,N_3515);
nor U4220 (N_4220,N_3813,N_2028);
or U4221 (N_4221,N_3785,N_3385);
or U4222 (N_4222,N_2858,N_2522);
nor U4223 (N_4223,N_2583,N_3783);
nor U4224 (N_4224,N_2574,N_3613);
xor U4225 (N_4225,N_2570,N_3715);
and U4226 (N_4226,N_3767,N_2038);
and U4227 (N_4227,N_3534,N_3309);
nor U4228 (N_4228,N_2603,N_3128);
nand U4229 (N_4229,N_3400,N_3928);
nor U4230 (N_4230,N_3630,N_3650);
nor U4231 (N_4231,N_3802,N_3931);
xnor U4232 (N_4232,N_3567,N_3358);
nand U4233 (N_4233,N_3660,N_3264);
xor U4234 (N_4234,N_2710,N_3542);
xor U4235 (N_4235,N_2658,N_3244);
and U4236 (N_4236,N_2009,N_3572);
xnor U4237 (N_4237,N_2987,N_3884);
and U4238 (N_4238,N_2485,N_3797);
nand U4239 (N_4239,N_2621,N_3837);
nand U4240 (N_4240,N_2171,N_3126);
xor U4241 (N_4241,N_3635,N_2447);
or U4242 (N_4242,N_2898,N_3988);
nand U4243 (N_4243,N_3432,N_2224);
and U4244 (N_4244,N_3532,N_2653);
xor U4245 (N_4245,N_3553,N_2660);
or U4246 (N_4246,N_3493,N_2615);
and U4247 (N_4247,N_2424,N_3267);
xnor U4248 (N_4248,N_3993,N_3462);
and U4249 (N_4249,N_2497,N_2914);
nor U4250 (N_4250,N_2609,N_3663);
and U4251 (N_4251,N_2938,N_2954);
nand U4252 (N_4252,N_2293,N_3329);
or U4253 (N_4253,N_3679,N_2732);
xnor U4254 (N_4254,N_3181,N_3258);
nor U4255 (N_4255,N_3720,N_2416);
xnor U4256 (N_4256,N_2880,N_2403);
nor U4257 (N_4257,N_3548,N_3473);
or U4258 (N_4258,N_3075,N_3456);
and U4259 (N_4259,N_3642,N_3591);
nor U4260 (N_4260,N_3727,N_3148);
nand U4261 (N_4261,N_2657,N_2272);
nand U4262 (N_4262,N_2879,N_3669);
and U4263 (N_4263,N_2753,N_2791);
nor U4264 (N_4264,N_3295,N_3092);
nand U4265 (N_4265,N_2287,N_3702);
nor U4266 (N_4266,N_2552,N_2749);
nor U4267 (N_4267,N_2432,N_2425);
xor U4268 (N_4268,N_2949,N_2176);
nand U4269 (N_4269,N_3155,N_3229);
xnor U4270 (N_4270,N_3447,N_2565);
or U4271 (N_4271,N_3768,N_3735);
or U4272 (N_4272,N_2206,N_2439);
xor U4273 (N_4273,N_3955,N_3791);
nand U4274 (N_4274,N_2040,N_2643);
nand U4275 (N_4275,N_3158,N_2645);
nor U4276 (N_4276,N_3270,N_2608);
and U4277 (N_4277,N_3083,N_2511);
xnor U4278 (N_4278,N_3015,N_2602);
and U4279 (N_4279,N_3730,N_2891);
and U4280 (N_4280,N_3357,N_2156);
nor U4281 (N_4281,N_3482,N_3488);
nand U4282 (N_4282,N_2590,N_2277);
or U4283 (N_4283,N_2183,N_2991);
nand U4284 (N_4284,N_2509,N_2943);
and U4285 (N_4285,N_2527,N_2214);
xor U4286 (N_4286,N_3061,N_3627);
and U4287 (N_4287,N_2123,N_3757);
or U4288 (N_4288,N_2429,N_2778);
or U4289 (N_4289,N_2956,N_3846);
nor U4290 (N_4290,N_3632,N_2291);
xnor U4291 (N_4291,N_3565,N_3098);
and U4292 (N_4292,N_2867,N_3071);
xnor U4293 (N_4293,N_3976,N_3753);
or U4294 (N_4294,N_3084,N_2130);
or U4295 (N_4295,N_2515,N_2461);
or U4296 (N_4296,N_2396,N_2152);
xor U4297 (N_4297,N_3932,N_3000);
or U4298 (N_4298,N_2832,N_2045);
nor U4299 (N_4299,N_3648,N_3734);
nor U4300 (N_4300,N_2472,N_3547);
nand U4301 (N_4301,N_2652,N_3894);
or U4302 (N_4302,N_2888,N_3873);
nor U4303 (N_4303,N_3105,N_2117);
nand U4304 (N_4304,N_3654,N_2523);
nand U4305 (N_4305,N_3242,N_3459);
or U4306 (N_4306,N_2729,N_3710);
and U4307 (N_4307,N_2840,N_2099);
or U4308 (N_4308,N_3134,N_2209);
xnor U4309 (N_4309,N_2528,N_3577);
nand U4310 (N_4310,N_2157,N_3945);
or U4311 (N_4311,N_3862,N_3247);
nor U4312 (N_4312,N_3854,N_2132);
and U4313 (N_4313,N_3034,N_2268);
or U4314 (N_4314,N_2012,N_3683);
nand U4315 (N_4315,N_2128,N_3398);
and U4316 (N_4316,N_2758,N_3481);
and U4317 (N_4317,N_3259,N_3771);
and U4318 (N_4318,N_2136,N_2296);
nor U4319 (N_4319,N_2654,N_3850);
and U4320 (N_4320,N_3496,N_2475);
nand U4321 (N_4321,N_3342,N_3688);
nand U4322 (N_4322,N_2636,N_3145);
nand U4323 (N_4323,N_3832,N_3222);
xor U4324 (N_4324,N_2557,N_2232);
nor U4325 (N_4325,N_3033,N_2809);
xor U4326 (N_4326,N_2635,N_2064);
or U4327 (N_4327,N_3066,N_2221);
nor U4328 (N_4328,N_2542,N_3218);
or U4329 (N_4329,N_2251,N_2613);
xnor U4330 (N_4330,N_3423,N_2944);
and U4331 (N_4331,N_3234,N_3127);
xnor U4332 (N_4332,N_3230,N_2204);
and U4333 (N_4333,N_3305,N_2231);
and U4334 (N_4334,N_3282,N_3082);
xor U4335 (N_4335,N_3180,N_3561);
nor U4336 (N_4336,N_3549,N_3086);
and U4337 (N_4337,N_2167,N_3521);
or U4338 (N_4338,N_3213,N_3546);
xor U4339 (N_4339,N_2088,N_2155);
xnor U4340 (N_4340,N_3312,N_2764);
or U4341 (N_4341,N_2712,N_3420);
xnor U4342 (N_4342,N_2588,N_2462);
and U4343 (N_4343,N_3882,N_3517);
or U4344 (N_4344,N_3296,N_2482);
xnor U4345 (N_4345,N_2193,N_2995);
nor U4346 (N_4346,N_3210,N_3073);
or U4347 (N_4347,N_2743,N_3494);
and U4348 (N_4348,N_3840,N_2674);
nand U4349 (N_4349,N_3707,N_3516);
and U4350 (N_4350,N_2717,N_3933);
or U4351 (N_4351,N_2444,N_2885);
and U4352 (N_4352,N_3631,N_2755);
and U4353 (N_4353,N_2752,N_2664);
nand U4354 (N_4354,N_3805,N_3843);
xor U4355 (N_4355,N_2671,N_2510);
nand U4356 (N_4356,N_2963,N_2213);
nand U4357 (N_4357,N_2044,N_3918);
nand U4358 (N_4358,N_3951,N_2386);
or U4359 (N_4359,N_2347,N_2626);
xor U4360 (N_4360,N_2524,N_2812);
nand U4361 (N_4361,N_2586,N_2966);
nor U4362 (N_4362,N_3043,N_2869);
nand U4363 (N_4363,N_2039,N_3841);
nand U4364 (N_4364,N_2399,N_3977);
and U4365 (N_4365,N_3205,N_3886);
or U4366 (N_4366,N_3002,N_3431);
nor U4367 (N_4367,N_2433,N_2631);
or U4368 (N_4368,N_3020,N_3774);
nand U4369 (N_4369,N_2856,N_3208);
nor U4370 (N_4370,N_2795,N_3826);
xnor U4371 (N_4371,N_3781,N_3293);
nand U4372 (N_4372,N_3411,N_3370);
nor U4373 (N_4373,N_3275,N_2773);
or U4374 (N_4374,N_2113,N_3506);
or U4375 (N_4375,N_3652,N_3335);
nand U4376 (N_4376,N_3906,N_3848);
or U4377 (N_4377,N_2675,N_3543);
and U4378 (N_4378,N_3404,N_2727);
nor U4379 (N_4379,N_3752,N_2324);
nor U4380 (N_4380,N_2883,N_2477);
nand U4381 (N_4381,N_3064,N_3666);
or U4382 (N_4382,N_3717,N_3041);
and U4383 (N_4383,N_3646,N_2378);
and U4384 (N_4384,N_3037,N_3662);
or U4385 (N_4385,N_3967,N_3177);
nor U4386 (N_4386,N_3240,N_3383);
nor U4387 (N_4387,N_3691,N_2464);
nand U4388 (N_4388,N_3649,N_3007);
and U4389 (N_4389,N_3483,N_2910);
and U4390 (N_4390,N_3289,N_3334);
nor U4391 (N_4391,N_2833,N_2325);
nand U4392 (N_4392,N_3507,N_3830);
and U4393 (N_4393,N_2203,N_3857);
xor U4394 (N_4394,N_2179,N_2693);
nor U4395 (N_4395,N_2016,N_3819);
and U4396 (N_4396,N_2159,N_2500);
and U4397 (N_4397,N_3780,N_3280);
xnor U4398 (N_4398,N_2521,N_2368);
and U4399 (N_4399,N_2813,N_3937);
xor U4400 (N_4400,N_3300,N_2312);
xor U4401 (N_4401,N_2682,N_2721);
nand U4402 (N_4402,N_2154,N_2714);
and U4403 (N_4403,N_3583,N_2980);
and U4404 (N_4404,N_3812,N_3094);
xnor U4405 (N_4405,N_3390,N_3725);
and U4406 (N_4406,N_3239,N_3681);
nand U4407 (N_4407,N_3243,N_2048);
and U4408 (N_4408,N_2855,N_2936);
nor U4409 (N_4409,N_2133,N_2034);
xor U4410 (N_4410,N_2875,N_2924);
nand U4411 (N_4411,N_3363,N_3944);
nand U4412 (N_4412,N_2971,N_2990);
xor U4413 (N_4413,N_2318,N_3274);
nand U4414 (N_4414,N_3413,N_2578);
nor U4415 (N_4415,N_3103,N_2831);
or U4416 (N_4416,N_3497,N_3700);
xor U4417 (N_4417,N_2359,N_3570);
or U4418 (N_4418,N_2544,N_3589);
or U4419 (N_4419,N_3923,N_3437);
nand U4420 (N_4420,N_2930,N_3733);
and U4421 (N_4421,N_3202,N_3776);
and U4422 (N_4422,N_2928,N_2256);
or U4423 (N_4423,N_3880,N_3038);
and U4424 (N_4424,N_2535,N_2501);
nand U4425 (N_4425,N_2862,N_2899);
nand U4426 (N_4426,N_3792,N_2299);
nor U4427 (N_4427,N_3745,N_3478);
nor U4428 (N_4428,N_2865,N_2457);
nand U4429 (N_4429,N_2345,N_3979);
nor U4430 (N_4430,N_2177,N_3332);
and U4431 (N_4431,N_2478,N_3904);
and U4432 (N_4432,N_3582,N_3339);
nand U4433 (N_4433,N_3595,N_2762);
nand U4434 (N_4434,N_3452,N_3994);
and U4435 (N_4435,N_3610,N_3048);
xnor U4436 (N_4436,N_2519,N_2115);
nand U4437 (N_4437,N_2087,N_3871);
and U4438 (N_4438,N_3965,N_2147);
xor U4439 (N_4439,N_3686,N_2093);
or U4440 (N_4440,N_3076,N_3868);
and U4441 (N_4441,N_3949,N_3056);
or U4442 (N_4442,N_3839,N_3817);
nor U4443 (N_4443,N_2919,N_3133);
xnor U4444 (N_4444,N_2228,N_3255);
nor U4445 (N_4445,N_2742,N_3141);
or U4446 (N_4446,N_3174,N_3869);
xor U4447 (N_4447,N_3612,N_3903);
or U4448 (N_4448,N_2111,N_2163);
xnor U4449 (N_4449,N_2056,N_3809);
nor U4450 (N_4450,N_2681,N_3641);
or U4451 (N_4451,N_2164,N_2101);
xnor U4452 (N_4452,N_2342,N_2137);
xnor U4453 (N_4453,N_3376,N_3775);
nor U4454 (N_4454,N_3881,N_3844);
nand U4455 (N_4455,N_3536,N_3586);
xor U4456 (N_4456,N_3711,N_2382);
nor U4457 (N_4457,N_2707,N_2997);
and U4458 (N_4458,N_3657,N_3454);
and U4459 (N_4459,N_3021,N_3226);
nand U4460 (N_4460,N_3694,N_2960);
or U4461 (N_4461,N_3197,N_3605);
nand U4462 (N_4462,N_2967,N_3268);
or U4463 (N_4463,N_3922,N_2053);
nor U4464 (N_4464,N_3909,N_3337);
and U4465 (N_4465,N_3132,N_3438);
nor U4466 (N_4466,N_2575,N_3055);
nand U4467 (N_4467,N_2953,N_3059);
and U4468 (N_4468,N_3120,N_2623);
nor U4469 (N_4469,N_3192,N_3025);
nand U4470 (N_4470,N_2071,N_3171);
and U4471 (N_4471,N_3260,N_2556);
xnor U4472 (N_4472,N_2321,N_2783);
xnor U4473 (N_4473,N_3053,N_3138);
nand U4474 (N_4474,N_2957,N_2008);
or U4475 (N_4475,N_3505,N_2746);
nand U4476 (N_4476,N_2902,N_3878);
and U4477 (N_4477,N_2442,N_3194);
and U4478 (N_4478,N_2310,N_2002);
or U4479 (N_4479,N_3495,N_3044);
nand U4480 (N_4480,N_3685,N_2601);
nand U4481 (N_4481,N_2922,N_2955);
and U4482 (N_4482,N_3371,N_3418);
nor U4483 (N_4483,N_2790,N_3394);
xor U4484 (N_4484,N_3634,N_3578);
and U4485 (N_4485,N_3525,N_3879);
or U4486 (N_4486,N_3384,N_3344);
and U4487 (N_4487,N_3011,N_2850);
xor U4488 (N_4488,N_3806,N_2929);
nand U4489 (N_4489,N_2916,N_3184);
or U4490 (N_4490,N_3831,N_3624);
or U4491 (N_4491,N_2627,N_3818);
and U4492 (N_4492,N_2961,N_3584);
nand U4493 (N_4493,N_3412,N_3430);
nor U4494 (N_4494,N_2269,N_2508);
nand U4495 (N_4495,N_2453,N_3032);
and U4496 (N_4496,N_3109,N_3475);
nand U4497 (N_4497,N_3814,N_3522);
nor U4498 (N_4498,N_3354,N_2323);
or U4499 (N_4499,N_2059,N_3552);
and U4500 (N_4500,N_3304,N_3468);
nor U4501 (N_4501,N_3924,N_3050);
nor U4502 (N_4502,N_2205,N_3816);
and U4503 (N_4503,N_2150,N_2218);
nor U4504 (N_4504,N_3311,N_3307);
xnor U4505 (N_4505,N_2904,N_2054);
or U4506 (N_4506,N_3535,N_3587);
or U4507 (N_4507,N_3860,N_2400);
xor U4508 (N_4508,N_3095,N_2706);
nor U4509 (N_4509,N_2290,N_3758);
and U4510 (N_4510,N_3623,N_3598);
nand U4511 (N_4511,N_3501,N_3703);
and U4512 (N_4512,N_2793,N_2861);
nor U4513 (N_4513,N_3308,N_3362);
nor U4514 (N_4514,N_3235,N_2859);
nand U4515 (N_4515,N_3175,N_3154);
or U4516 (N_4516,N_2109,N_3326);
nor U4517 (N_4517,N_3150,N_2017);
and U4518 (N_4518,N_2458,N_2090);
xor U4519 (N_4519,N_3336,N_2915);
nand U4520 (N_4520,N_3966,N_2502);
xor U4521 (N_4521,N_2572,N_2580);
or U4522 (N_4522,N_2959,N_2624);
nand U4523 (N_4523,N_3187,N_2644);
xor U4524 (N_4524,N_2950,N_2383);
xor U4525 (N_4525,N_3477,N_3246);
or U4526 (N_4526,N_2605,N_3980);
nor U4527 (N_4527,N_3327,N_3990);
and U4528 (N_4528,N_3983,N_3877);
nand U4529 (N_4529,N_2010,N_2385);
nand U4530 (N_4530,N_2823,N_2168);
xor U4531 (N_4531,N_2440,N_2229);
or U4532 (N_4532,N_2407,N_2366);
xnor U4533 (N_4533,N_2965,N_3223);
and U4534 (N_4534,N_3193,N_2815);
or U4535 (N_4535,N_2470,N_3262);
and U4536 (N_4536,N_3405,N_2110);
nor U4537 (N_4537,N_2116,N_3265);
nor U4538 (N_4538,N_2042,N_3701);
and U4539 (N_4539,N_3626,N_2165);
nor U4540 (N_4540,N_2138,N_2718);
xnor U4541 (N_4541,N_2662,N_3407);
and U4542 (N_4542,N_2243,N_3428);
and U4543 (N_4543,N_3953,N_3140);
nor U4544 (N_4544,N_3361,N_3530);
nand U4545 (N_4545,N_2673,N_2545);
and U4546 (N_4546,N_3749,N_2694);
nor U4547 (N_4547,N_3602,N_3353);
nor U4548 (N_4548,N_2633,N_2871);
xnor U4549 (N_4549,N_2210,N_2170);
or U4550 (N_4550,N_3867,N_2100);
or U4551 (N_4551,N_3346,N_2765);
xnor U4552 (N_4552,N_2274,N_2456);
nand U4553 (N_4553,N_2279,N_3217);
xnor U4554 (N_4554,N_2781,N_2225);
nor U4555 (N_4555,N_2446,N_3367);
nand U4556 (N_4556,N_3151,N_2849);
nor U4557 (N_4557,N_3051,N_2387);
nor U4558 (N_4558,N_2536,N_2217);
and U4559 (N_4559,N_3328,N_2405);
nor U4560 (N_4560,N_2406,N_2896);
and U4561 (N_4561,N_2486,N_2247);
xnor U4562 (N_4562,N_3704,N_3588);
or U4563 (N_4563,N_3731,N_2158);
xnor U4564 (N_4564,N_3204,N_2082);
or U4565 (N_4565,N_2661,N_2364);
and U4566 (N_4566,N_3368,N_2692);
nand U4567 (N_4567,N_3699,N_3712);
nand U4568 (N_4568,N_2697,N_2564);
nor U4569 (N_4569,N_3410,N_3269);
or U4570 (N_4570,N_3303,N_3509);
or U4571 (N_4571,N_3476,N_3324);
nand U4572 (N_4572,N_2494,N_2720);
xnor U4573 (N_4573,N_3251,N_2650);
and U4574 (N_4574,N_3065,N_3101);
nand U4575 (N_4575,N_2469,N_2078);
xor U4576 (N_4576,N_2768,N_2374);
xor U4577 (N_4577,N_3443,N_2422);
nor U4578 (N_4578,N_2567,N_3706);
nand U4579 (N_4579,N_2413,N_3902);
and U4580 (N_4580,N_3746,N_3458);
xor U4581 (N_4581,N_2190,N_3564);
nand U4582 (N_4582,N_2198,N_2241);
xor U4583 (N_4583,N_3442,N_3973);
nor U4584 (N_4584,N_2076,N_2261);
nand U4585 (N_4585,N_2197,N_2124);
and U4586 (N_4586,N_3261,N_3914);
or U4587 (N_4587,N_2362,N_3453);
or U4588 (N_4588,N_3645,N_3377);
nor U4589 (N_4589,N_2380,N_2402);
nor U4590 (N_4590,N_3018,N_2022);
nand U4591 (N_4591,N_3737,N_3968);
nor U4592 (N_4592,N_3381,N_3424);
nand U4593 (N_4593,N_2426,N_2573);
nand U4594 (N_4594,N_3489,N_2319);
xor U4595 (N_4595,N_2134,N_2935);
xnor U4596 (N_4596,N_3057,N_2282);
nor U4597 (N_4597,N_2219,N_3290);
or U4598 (N_4598,N_2549,N_2266);
nor U4599 (N_4599,N_3284,N_2437);
and U4600 (N_4600,N_3975,N_3072);
nor U4601 (N_4601,N_2827,N_3227);
nor U4602 (N_4602,N_2070,N_2787);
nand U4603 (N_4603,N_2445,N_2414);
nor U4604 (N_4604,N_2381,N_2267);
and U4605 (N_4605,N_3152,N_3003);
or U4606 (N_4606,N_2418,N_3079);
nand U4607 (N_4607,N_2751,N_2834);
nor U4608 (N_4608,N_2678,N_3513);
and U4609 (N_4609,N_3322,N_3161);
nand U4610 (N_4610,N_3360,N_2784);
nand U4611 (N_4611,N_3013,N_2122);
nand U4612 (N_4612,N_2139,N_2095);
or U4613 (N_4613,N_2043,N_2799);
or U4614 (N_4614,N_2467,N_2503);
or U4615 (N_4615,N_3277,N_2057);
or U4616 (N_4616,N_3518,N_2192);
nand U4617 (N_4617,N_2025,N_2893);
xor U4618 (N_4618,N_2186,N_3590);
nor U4619 (N_4619,N_2970,N_3907);
xor U4620 (N_4620,N_3985,N_2230);
nor U4621 (N_4621,N_3359,N_2484);
xnor U4622 (N_4622,N_2459,N_3708);
nor U4623 (N_4623,N_2612,N_3004);
or U4624 (N_4624,N_3684,N_3131);
or U4625 (N_4625,N_2270,N_2585);
and U4626 (N_4626,N_2866,N_2525);
nand U4627 (N_4627,N_3167,N_3391);
nor U4628 (N_4628,N_2235,N_3340);
nor U4629 (N_4629,N_2680,N_2103);
and U4630 (N_4630,N_3408,N_3622);
and U4631 (N_4631,N_2075,N_3416);
nand U4632 (N_4632,N_2032,N_3471);
xnor U4633 (N_4633,N_3759,N_2789);
nor U4634 (N_4634,N_3531,N_2463);
xor U4635 (N_4635,N_3330,N_3472);
and U4636 (N_4636,N_3036,N_3766);
and U4637 (N_4637,N_3996,N_3755);
nor U4638 (N_4638,N_2906,N_3693);
nor U4639 (N_4639,N_3962,N_3705);
nor U4640 (N_4640,N_2450,N_3122);
and U4641 (N_4641,N_2741,N_2105);
xor U4642 (N_4642,N_2672,N_2146);
xnor U4643 (N_4643,N_2908,N_2466);
or U4644 (N_4644,N_3670,N_2818);
nor U4645 (N_4645,N_2853,N_3115);
nand U4646 (N_4646,N_3035,N_3640);
or U4647 (N_4647,N_3166,N_3942);
or U4648 (N_4648,N_2805,N_3191);
nor U4649 (N_4649,N_2688,N_2972);
nand U4650 (N_4650,N_2227,N_2300);
xor U4651 (N_4651,N_3499,N_3574);
xnor U4652 (N_4652,N_2607,N_2298);
or U4653 (N_4653,N_3911,N_3085);
xnor U4654 (N_4654,N_2144,N_3378);
nand U4655 (N_4655,N_2617,N_3448);
xnor U4656 (N_4656,N_2195,N_3186);
xnor U4657 (N_4657,N_2801,N_2998);
or U4658 (N_4658,N_2532,N_3581);
or U4659 (N_4659,N_2512,N_2492);
nor U4660 (N_4660,N_2530,N_3793);
or U4661 (N_4661,N_3266,N_3957);
and U4662 (N_4662,N_3163,N_2548);
nand U4663 (N_4663,N_3333,N_3692);
nand U4664 (N_4664,N_2901,N_2593);
nor U4665 (N_4665,N_3845,N_2271);
nand U4666 (N_4666,N_3560,N_3777);
nand U4667 (N_4667,N_2848,N_3149);
nor U4668 (N_4668,N_2794,N_3738);
and U4669 (N_4669,N_3414,N_3219);
xor U4670 (N_4670,N_2622,N_3183);
or U4671 (N_4671,N_2730,N_3741);
and U4672 (N_4672,N_2331,N_3422);
and U4673 (N_4673,N_3556,N_2200);
nor U4674 (N_4674,N_2828,N_3677);
nor U4675 (N_4675,N_2052,N_2766);
nand U4676 (N_4676,N_2441,N_2006);
or U4677 (N_4677,N_3568,N_3827);
nand U4678 (N_4678,N_3136,N_3380);
or U4679 (N_4679,N_2777,N_2846);
or U4680 (N_4680,N_3563,N_3750);
xnor U4681 (N_4681,N_2890,N_3714);
xnor U4682 (N_4682,N_2807,N_3279);
nor U4683 (N_4683,N_3769,N_2107);
nor U4684 (N_4684,N_2835,N_3900);
xor U4685 (N_4685,N_3425,N_2563);
or U4686 (N_4686,N_3557,N_2945);
or U4687 (N_4687,N_2920,N_2733);
xor U4688 (N_4688,N_3971,N_3929);
or U4689 (N_4689,N_2632,N_3045);
and U4690 (N_4690,N_3999,N_3479);
xor U4691 (N_4691,N_2377,N_2351);
xnor U4692 (N_4692,N_2280,N_3726);
nor U4693 (N_4693,N_2531,N_3023);
nor U4694 (N_4694,N_3108,N_2452);
or U4695 (N_4695,N_3110,N_2517);
nor U4696 (N_4696,N_3789,N_2771);
nand U4697 (N_4697,N_3465,N_3956);
nand U4698 (N_4698,N_3352,N_3347);
nor U4699 (N_4699,N_2029,N_3935);
nand U4700 (N_4700,N_3474,N_3111);
nand U4701 (N_4701,N_3349,N_2999);
and U4702 (N_4702,N_3551,N_3653);
xor U4703 (N_4703,N_3940,N_3178);
nand U4704 (N_4704,N_3214,N_3485);
or U4705 (N_4705,N_2538,N_3313);
xnor U4706 (N_4706,N_3947,N_2691);
nand U4707 (N_4707,N_3665,N_2249);
nor U4708 (N_4708,N_2320,N_2131);
nor U4709 (N_4709,N_2825,N_3288);
and U4710 (N_4710,N_3022,N_2398);
and U4711 (N_4711,N_2208,N_2677);
nor U4712 (N_4712,N_3992,N_3528);
nor U4713 (N_4713,N_3916,N_2084);
xnor U4714 (N_4714,N_2560,N_3287);
xnor U4715 (N_4715,N_3318,N_2925);
or U4716 (N_4716,N_2162,N_2305);
xor U4717 (N_4717,N_3597,N_2863);
xnor U4718 (N_4718,N_2705,N_2984);
or U4719 (N_4719,N_2148,N_3674);
xor U4720 (N_4720,N_2666,N_3392);
and U4721 (N_4721,N_2327,N_2695);
xor U4722 (N_4722,N_3068,N_3946);
xnor U4723 (N_4723,N_2255,N_2685);
nor U4724 (N_4724,N_3409,N_2978);
nand U4725 (N_4725,N_2365,N_2395);
or U4726 (N_4726,N_3636,N_3672);
nand U4727 (N_4727,N_3042,N_2946);
nor U4728 (N_4728,N_3253,N_3639);
and U4729 (N_4729,N_2143,N_2775);
or U4730 (N_4730,N_3822,N_2068);
or U4731 (N_4731,N_3348,N_3441);
xnor U4732 (N_4732,N_3470,N_3467);
nor U4733 (N_4733,N_2188,N_2638);
nand U4734 (N_4734,N_2505,N_2912);
nand U4735 (N_4735,N_2947,N_2819);
and U4736 (N_4736,N_3321,N_2253);
xnor U4737 (N_4737,N_2792,N_2417);
xnor U4738 (N_4738,N_2628,N_3502);
nand U4739 (N_4739,N_3823,N_2599);
or U4740 (N_4740,N_3046,N_3875);
nor U4741 (N_4741,N_3599,N_2410);
and U4742 (N_4742,N_2435,N_3350);
or U4743 (N_4743,N_2184,N_3866);
and U4744 (N_4744,N_2011,N_2220);
nand U4745 (N_4745,N_2036,N_2926);
and U4746 (N_4746,N_2800,N_3216);
and U4747 (N_4747,N_2185,N_2698);
or U4748 (N_4748,N_2360,N_3647);
and U4749 (N_4749,N_2992,N_3179);
and U4750 (N_4750,N_3124,N_2289);
or U4751 (N_4751,N_3256,N_3052);
nor U4752 (N_4752,N_3207,N_2499);
or U4753 (N_4753,N_3524,N_2576);
nand U4754 (N_4754,N_2121,N_2983);
nor U4755 (N_4755,N_3457,N_2178);
and U4756 (N_4756,N_3910,N_3689);
nor U4757 (N_4757,N_3596,N_2985);
nor U4758 (N_4758,N_3943,N_3861);
xor U4759 (N_4759,N_2389,N_2543);
nand U4760 (N_4760,N_2313,N_2587);
nor U4761 (N_4761,N_3221,N_3355);
and U4762 (N_4762,N_2656,N_3939);
nor U4763 (N_4763,N_2937,N_3659);
xnor U4764 (N_4764,N_3963,N_2285);
and U4765 (N_4765,N_2149,N_3019);
or U4766 (N_4766,N_3142,N_2246);
nor U4767 (N_4767,N_2600,N_3049);
nand U4768 (N_4768,N_3748,N_2932);
nor U4769 (N_4769,N_3157,N_2655);
nand U4770 (N_4770,N_3434,N_3618);
xnor U4771 (N_4771,N_2049,N_2000);
nand U4772 (N_4772,N_3310,N_3756);
or U4773 (N_4773,N_2637,N_3995);
or U4774 (N_4774,N_2145,N_2562);
nand U4775 (N_4775,N_3890,N_2465);
xnor U4776 (N_4776,N_3761,N_3107);
or U4777 (N_4777,N_3678,N_3593);
nor U4778 (N_4778,N_2083,N_2234);
and U4779 (N_4779,N_2479,N_3006);
or U4780 (N_4780,N_2344,N_3106);
nand U4781 (N_4781,N_2001,N_2646);
xor U4782 (N_4782,N_2189,N_2236);
nor U4783 (N_4783,N_3533,N_2566);
and U4784 (N_4784,N_2592,N_3077);
nand U4785 (N_4785,N_3828,N_2931);
xor U4786 (N_4786,N_3220,N_2423);
nand U4787 (N_4787,N_2640,N_2302);
nand U4788 (N_4788,N_3540,N_2606);
nor U4789 (N_4789,N_2735,N_2066);
or U4790 (N_4790,N_3573,N_3656);
or U4791 (N_4791,N_3575,N_2072);
xor U4792 (N_4792,N_3016,N_2537);
nand U4793 (N_4793,N_2372,N_2569);
or U4794 (N_4794,N_2939,N_2489);
xor U4795 (N_4795,N_3241,N_2035);
or U4796 (N_4796,N_3628,N_3772);
xor U4797 (N_4797,N_2264,N_2887);
xor U4798 (N_4798,N_2373,N_2363);
nor U4799 (N_4799,N_2547,N_3100);
xor U4800 (N_4800,N_3427,N_2767);
or U4801 (N_4801,N_2982,N_2352);
and U4802 (N_4802,N_3529,N_2014);
xor U4803 (N_4803,N_3067,N_3611);
nand U4804 (N_4804,N_3070,N_3740);
and U4805 (N_4805,N_2326,N_2211);
nand U4806 (N_4806,N_2810,N_2976);
nor U4807 (N_4807,N_2112,N_2384);
nand U4808 (N_4808,N_2443,N_2258);
nor U4809 (N_4809,N_2242,N_2734);
and U4810 (N_4810,N_2806,N_2689);
nor U4811 (N_4811,N_3466,N_2311);
and U4812 (N_4812,N_2709,N_3778);
nand U4813 (N_4813,N_2436,N_3491);
xor U4814 (N_4814,N_3294,N_2553);
nor U4815 (N_4815,N_2379,N_2739);
nand U4816 (N_4816,N_3539,N_2018);
nand U4817 (N_4817,N_3961,N_3765);
and U4818 (N_4818,N_3089,N_2153);
and U4819 (N_4819,N_3276,N_3545);
and U4820 (N_4820,N_2826,N_2455);
or U4821 (N_4821,N_3614,N_2921);
nor U4822 (N_4822,N_3600,N_2077);
or U4823 (N_4823,N_3782,N_2785);
and U4824 (N_4824,N_3317,N_3188);
nor U4825 (N_4825,N_3492,N_2394);
and U4826 (N_4826,N_3445,N_3074);
nor U4827 (N_4827,N_2196,N_3382);
nor U4828 (N_4828,N_2226,N_2166);
nor U4829 (N_4829,N_3608,N_2252);
or U4830 (N_4830,N_3199,N_3554);
and U4831 (N_4831,N_3415,N_3406);
nor U4832 (N_4832,N_3320,N_2540);
xor U4833 (N_4833,N_2421,N_3695);
or U4834 (N_4834,N_3450,N_2353);
nor U4835 (N_4835,N_3298,N_2401);
nand U4836 (N_4836,N_2770,N_3760);
nor U4837 (N_4837,N_2882,N_2371);
xnor U4838 (N_4838,N_3989,N_3562);
nor U4839 (N_4839,N_3538,N_3090);
nand U4840 (N_4840,N_3544,N_2715);
nor U4841 (N_4841,N_2774,N_3212);
nand U4842 (N_4842,N_2391,N_3576);
xnor U4843 (N_4843,N_3713,N_3801);
nand U4844 (N_4844,N_3585,N_2013);
nand U4845 (N_4845,N_3851,N_2278);
or U4846 (N_4846,N_2905,N_3905);
and U4847 (N_4847,N_2097,N_2897);
nand U4848 (N_4848,N_2620,N_3169);
and U4849 (N_4849,N_3143,N_3779);
nor U4850 (N_4850,N_3728,N_3742);
nand U4851 (N_4851,N_3024,N_2736);
nor U4852 (N_4852,N_2303,N_2907);
nand U4853 (N_4853,N_2094,N_3736);
or U4854 (N_4854,N_3913,N_2595);
nand U4855 (N_4855,N_3254,N_2215);
nand U4856 (N_4856,N_3446,N_2288);
nor U4857 (N_4857,N_3744,N_3097);
and U4858 (N_4858,N_3526,N_3369);
and U4859 (N_4859,N_2881,N_2027);
or U4860 (N_4860,N_2480,N_2160);
xor U4861 (N_4861,N_2346,N_3807);
nand U4862 (N_4862,N_3795,N_3764);
or U4863 (N_4863,N_3763,N_3651);
and U4864 (N_4864,N_2322,N_3658);
nand U4865 (N_4865,N_3603,N_2745);
or U4866 (N_4866,N_3008,N_2952);
and U4867 (N_4867,N_3541,N_3232);
xor U4868 (N_4868,N_3225,N_2428);
nand U4869 (N_4869,N_2589,N_3964);
and U4870 (N_4870,N_2641,N_3093);
nor U4871 (N_4871,N_2824,N_3189);
xnor U4872 (N_4872,N_3682,N_3233);
nand U4873 (N_4873,N_3160,N_3773);
nand U4874 (N_4874,N_3009,N_3001);
nor U4875 (N_4875,N_3865,N_2375);
nand U4876 (N_4876,N_3917,N_2533);
xnor U4877 (N_4877,N_3291,N_3786);
nor U4878 (N_4878,N_2273,N_3719);
xnor U4879 (N_4879,N_2004,N_3201);
xor U4880 (N_4880,N_2431,N_2895);
or U4881 (N_4881,N_2046,N_2297);
nor U4882 (N_4882,N_2598,N_2260);
xor U4883 (N_4883,N_2355,N_2659);
nor U4884 (N_4884,N_2716,N_2308);
nand U4885 (N_4885,N_2837,N_2438);
nand U4886 (N_4886,N_2559,N_3800);
or U4887 (N_4887,N_3722,N_2974);
and U4888 (N_4888,N_2518,N_2647);
xnor U4889 (N_4889,N_3185,N_3512);
xnor U4890 (N_4890,N_2900,N_2722);
and U4891 (N_4891,N_3114,N_3500);
nand U4892 (N_4892,N_2393,N_2968);
nand U4893 (N_4893,N_3102,N_2015);
nand U4894 (N_4894,N_3721,N_2275);
or U4895 (N_4895,N_2738,N_3464);
and U4896 (N_4896,N_3555,N_3676);
and U4897 (N_4897,N_3566,N_2520);
or U4898 (N_4898,N_2619,N_3263);
nor U4899 (N_4899,N_3609,N_2630);
nor U4900 (N_4900,N_2341,N_3272);
and U4901 (N_4901,N_2257,N_2663);
xnor U4902 (N_4902,N_3062,N_3402);
and U4903 (N_4903,N_2839,N_2415);
or U4904 (N_4904,N_2909,N_2872);
nand U4905 (N_4905,N_3123,N_2356);
xor U4906 (N_4906,N_3842,N_2216);
nor U4907 (N_4907,N_2182,N_2449);
nand U4908 (N_4908,N_3604,N_3889);
xnor U4909 (N_4909,N_2740,N_3228);
xor U4910 (N_4910,N_2062,N_2811);
or U4911 (N_4911,N_3387,N_3891);
xnor U4912 (N_4912,N_3815,N_2857);
nor U4913 (N_4913,N_2591,N_3116);
nor U4914 (N_4914,N_3803,N_2713);
xnor U4915 (N_4915,N_2788,N_3005);
or U4916 (N_4916,N_2504,N_2031);
nor U4917 (N_4917,N_3824,N_2551);
or U4918 (N_4918,N_2317,N_2568);
nor U4919 (N_4919,N_2161,N_3397);
nand U4920 (N_4920,N_3147,N_3302);
nand U4921 (N_4921,N_2187,N_2820);
nand U4922 (N_4922,N_2816,N_3696);
xor U4923 (N_4923,N_2019,N_2821);
xnor U4924 (N_4924,N_2020,N_3997);
xor U4925 (N_4925,N_3137,N_2309);
and U4926 (N_4926,N_3063,N_2977);
xnor U4927 (N_4927,N_3498,N_3709);
or U4928 (N_4928,N_3182,N_3883);
and U4929 (N_4929,N_2108,N_2838);
xor U4930 (N_4930,N_3510,N_3927);
nand U4931 (N_4931,N_2073,N_3743);
xor U4932 (N_4932,N_3206,N_3257);
nor U4933 (N_4933,N_2328,N_3633);
xnor U4934 (N_4934,N_2933,N_2942);
xor U4935 (N_4935,N_3982,N_2067);
nor U4936 (N_4936,N_2033,N_2408);
nor U4937 (N_4937,N_3164,N_2069);
or U4938 (N_4938,N_2934,N_2180);
xnor U4939 (N_4939,N_3671,N_3960);
and U4940 (N_4940,N_2358,N_3852);
nor U4941 (N_4941,N_2191,N_2796);
and U4942 (N_4942,N_3970,N_3503);
nand U4943 (N_4943,N_2851,N_2314);
nor U4944 (N_4944,N_3571,N_2007);
xnor U4945 (N_4945,N_2594,N_3104);
and U4946 (N_4946,N_3460,N_2604);
nand U4947 (N_4947,N_3237,N_2975);
and U4948 (N_4948,N_3754,N_3306);
xor U4949 (N_4949,N_2181,N_3747);
or U4950 (N_4950,N_3978,N_2687);
and U4951 (N_4951,N_3338,N_3486);
nor U4952 (N_4952,N_2023,N_2702);
nor U4953 (N_4953,N_2496,N_3794);
or U4954 (N_4954,N_3887,N_2723);
or U4955 (N_4955,N_2696,N_2639);
and U4956 (N_4956,N_2420,N_2940);
nor U4957 (N_4957,N_3030,N_2493);
xnor U4958 (N_4958,N_3527,N_2726);
nand U4959 (N_4959,N_2911,N_2283);
xor U4960 (N_4960,N_2506,N_2854);
and U4961 (N_4961,N_3796,N_3028);
nand U4962 (N_4962,N_2876,N_3723);
xnor U4963 (N_4963,N_2962,N_3859);
nor U4964 (N_4964,N_3379,N_3215);
and U4965 (N_4965,N_3017,N_3463);
nand U4966 (N_4966,N_2830,N_2634);
nand U4967 (N_4967,N_3519,N_2079);
and U4968 (N_4968,N_3372,N_2126);
and U4969 (N_4969,N_2841,N_3156);
xnor U4970 (N_4970,N_2102,N_2989);
xnor U4971 (N_4971,N_2701,N_2330);
xor U4972 (N_4972,N_3770,N_3129);
and U4973 (N_4973,N_2051,N_3925);
or U4974 (N_4974,N_3252,N_2719);
xnor U4975 (N_4975,N_3389,N_3047);
xnor U4976 (N_4976,N_3697,N_2491);
nor U4977 (N_4977,N_3950,N_2581);
nor U4978 (N_4978,N_2683,N_3099);
xnor U4979 (N_4979,N_2388,N_3998);
xnor U4980 (N_4980,N_3625,N_2555);
xor U4981 (N_4981,N_3888,N_2769);
or U4982 (N_4982,N_2451,N_3401);
xor U4983 (N_4983,N_3972,N_3619);
nor U4984 (N_4984,N_2964,N_2786);
nand U4985 (N_4985,N_2754,N_3606);
and U4986 (N_4986,N_2348,N_2175);
or U4987 (N_4987,N_3278,N_3283);
and U4988 (N_4988,N_3668,N_2913);
nand U4989 (N_4989,N_2969,N_3520);
and U4990 (N_4990,N_2086,N_2744);
xor U4991 (N_4991,N_2836,N_3959);
nor U4992 (N_4992,N_3592,N_2357);
xnor U4993 (N_4993,N_2629,N_2731);
or U4994 (N_4994,N_2376,N_2172);
nand U4995 (N_4995,N_2724,N_3331);
nand U4996 (N_4996,N_2618,N_2037);
nand U4997 (N_4997,N_2625,N_3898);
nor U4998 (N_4998,N_3299,N_3908);
xor U4999 (N_4999,N_2284,N_2354);
or U5000 (N_5000,N_3963,N_3596);
or U5001 (N_5001,N_3673,N_2849);
xor U5002 (N_5002,N_3839,N_3864);
xor U5003 (N_5003,N_2186,N_2061);
xnor U5004 (N_5004,N_2528,N_2081);
xor U5005 (N_5005,N_3935,N_3504);
xnor U5006 (N_5006,N_3490,N_2196);
and U5007 (N_5007,N_3470,N_2726);
nand U5008 (N_5008,N_3333,N_3385);
nand U5009 (N_5009,N_2954,N_2720);
nand U5010 (N_5010,N_3774,N_3553);
and U5011 (N_5011,N_2630,N_3526);
xor U5012 (N_5012,N_2808,N_2368);
nor U5013 (N_5013,N_3355,N_2227);
nor U5014 (N_5014,N_3974,N_2907);
and U5015 (N_5015,N_3379,N_2073);
and U5016 (N_5016,N_3385,N_3162);
and U5017 (N_5017,N_2278,N_2925);
nand U5018 (N_5018,N_3820,N_3682);
or U5019 (N_5019,N_3762,N_3171);
or U5020 (N_5020,N_2786,N_3863);
nand U5021 (N_5021,N_3148,N_2633);
nor U5022 (N_5022,N_3326,N_3759);
nor U5023 (N_5023,N_2981,N_2564);
or U5024 (N_5024,N_3891,N_3112);
and U5025 (N_5025,N_3603,N_3823);
nand U5026 (N_5026,N_3808,N_3602);
and U5027 (N_5027,N_2919,N_2061);
xor U5028 (N_5028,N_2136,N_3535);
xnor U5029 (N_5029,N_3296,N_2411);
and U5030 (N_5030,N_3550,N_3433);
nand U5031 (N_5031,N_3386,N_2904);
nor U5032 (N_5032,N_3030,N_3551);
or U5033 (N_5033,N_2771,N_2824);
xor U5034 (N_5034,N_3838,N_3723);
xor U5035 (N_5035,N_3826,N_3028);
nand U5036 (N_5036,N_2295,N_3741);
or U5037 (N_5037,N_3585,N_3150);
and U5038 (N_5038,N_2810,N_2659);
xor U5039 (N_5039,N_3999,N_2159);
nand U5040 (N_5040,N_2760,N_3339);
or U5041 (N_5041,N_3504,N_2728);
and U5042 (N_5042,N_2762,N_3397);
and U5043 (N_5043,N_2286,N_3019);
nand U5044 (N_5044,N_2212,N_2022);
nor U5045 (N_5045,N_2549,N_3424);
and U5046 (N_5046,N_2522,N_2231);
and U5047 (N_5047,N_2915,N_2296);
nand U5048 (N_5048,N_2791,N_3949);
xor U5049 (N_5049,N_2671,N_2705);
xor U5050 (N_5050,N_2665,N_2412);
nor U5051 (N_5051,N_3663,N_3370);
xnor U5052 (N_5052,N_2012,N_3472);
xnor U5053 (N_5053,N_2379,N_3073);
and U5054 (N_5054,N_2257,N_3938);
and U5055 (N_5055,N_3636,N_3177);
nor U5056 (N_5056,N_3270,N_2345);
or U5057 (N_5057,N_2590,N_3923);
or U5058 (N_5058,N_2446,N_2983);
and U5059 (N_5059,N_3560,N_3444);
nor U5060 (N_5060,N_2107,N_3805);
nor U5061 (N_5061,N_2759,N_2274);
nor U5062 (N_5062,N_2523,N_2272);
xor U5063 (N_5063,N_3244,N_2639);
nor U5064 (N_5064,N_3045,N_3358);
nor U5065 (N_5065,N_3866,N_2052);
or U5066 (N_5066,N_2157,N_3135);
nand U5067 (N_5067,N_3284,N_2529);
nor U5068 (N_5068,N_2963,N_3449);
and U5069 (N_5069,N_2498,N_2741);
xnor U5070 (N_5070,N_3906,N_2996);
xnor U5071 (N_5071,N_2295,N_3071);
xnor U5072 (N_5072,N_2215,N_2077);
and U5073 (N_5073,N_2342,N_2732);
xnor U5074 (N_5074,N_2218,N_2622);
xor U5075 (N_5075,N_3237,N_2593);
or U5076 (N_5076,N_2255,N_3805);
xor U5077 (N_5077,N_3407,N_2411);
nand U5078 (N_5078,N_3653,N_2999);
nor U5079 (N_5079,N_2979,N_2689);
xor U5080 (N_5080,N_2197,N_2914);
or U5081 (N_5081,N_3095,N_2371);
nor U5082 (N_5082,N_2136,N_3497);
nor U5083 (N_5083,N_2908,N_2541);
and U5084 (N_5084,N_2944,N_3786);
and U5085 (N_5085,N_2948,N_2757);
and U5086 (N_5086,N_3087,N_3750);
and U5087 (N_5087,N_3039,N_3299);
xnor U5088 (N_5088,N_3135,N_2201);
xor U5089 (N_5089,N_3203,N_2445);
xnor U5090 (N_5090,N_3433,N_2830);
nand U5091 (N_5091,N_3996,N_3255);
nand U5092 (N_5092,N_3136,N_2612);
xnor U5093 (N_5093,N_2662,N_3273);
xnor U5094 (N_5094,N_2721,N_2676);
and U5095 (N_5095,N_2903,N_3567);
or U5096 (N_5096,N_2242,N_3636);
and U5097 (N_5097,N_2121,N_2477);
nor U5098 (N_5098,N_3943,N_3926);
nand U5099 (N_5099,N_2650,N_2942);
nor U5100 (N_5100,N_2989,N_2274);
xnor U5101 (N_5101,N_3846,N_2858);
or U5102 (N_5102,N_3052,N_3786);
or U5103 (N_5103,N_3340,N_2405);
and U5104 (N_5104,N_2913,N_3635);
xor U5105 (N_5105,N_3226,N_2374);
nand U5106 (N_5106,N_3721,N_3461);
nor U5107 (N_5107,N_3934,N_3002);
nand U5108 (N_5108,N_3325,N_2902);
or U5109 (N_5109,N_3003,N_3489);
xnor U5110 (N_5110,N_3020,N_3114);
and U5111 (N_5111,N_2458,N_2020);
and U5112 (N_5112,N_3185,N_3544);
xor U5113 (N_5113,N_2177,N_3223);
xor U5114 (N_5114,N_2421,N_2396);
xnor U5115 (N_5115,N_3555,N_2901);
or U5116 (N_5116,N_3209,N_3726);
and U5117 (N_5117,N_3965,N_2152);
or U5118 (N_5118,N_3574,N_2391);
and U5119 (N_5119,N_3715,N_2398);
nor U5120 (N_5120,N_3389,N_2783);
xnor U5121 (N_5121,N_3262,N_2175);
nand U5122 (N_5122,N_2159,N_3480);
xor U5123 (N_5123,N_3497,N_3926);
xor U5124 (N_5124,N_2202,N_2402);
nor U5125 (N_5125,N_3719,N_2605);
and U5126 (N_5126,N_3158,N_2175);
nor U5127 (N_5127,N_2870,N_2398);
or U5128 (N_5128,N_2236,N_2262);
nand U5129 (N_5129,N_2671,N_2222);
nand U5130 (N_5130,N_2614,N_3532);
xor U5131 (N_5131,N_3826,N_2732);
xor U5132 (N_5132,N_3405,N_2851);
xnor U5133 (N_5133,N_2328,N_2570);
xor U5134 (N_5134,N_2887,N_2822);
nor U5135 (N_5135,N_3818,N_3467);
and U5136 (N_5136,N_2477,N_2248);
nor U5137 (N_5137,N_2949,N_3417);
nand U5138 (N_5138,N_3852,N_3301);
nor U5139 (N_5139,N_3438,N_3608);
or U5140 (N_5140,N_3414,N_2299);
xor U5141 (N_5141,N_2940,N_2182);
and U5142 (N_5142,N_2651,N_2663);
nand U5143 (N_5143,N_2643,N_3231);
nand U5144 (N_5144,N_3392,N_2310);
nor U5145 (N_5145,N_3691,N_3959);
nor U5146 (N_5146,N_2117,N_2700);
or U5147 (N_5147,N_2913,N_2105);
nand U5148 (N_5148,N_3705,N_2274);
nor U5149 (N_5149,N_2684,N_3289);
xor U5150 (N_5150,N_3787,N_2623);
and U5151 (N_5151,N_2296,N_2274);
xor U5152 (N_5152,N_2191,N_2965);
nor U5153 (N_5153,N_3252,N_2774);
or U5154 (N_5154,N_2622,N_2263);
and U5155 (N_5155,N_2921,N_2622);
nand U5156 (N_5156,N_2598,N_2926);
or U5157 (N_5157,N_2023,N_2465);
and U5158 (N_5158,N_2367,N_2457);
or U5159 (N_5159,N_3381,N_2950);
nor U5160 (N_5160,N_3060,N_3248);
and U5161 (N_5161,N_2037,N_3499);
and U5162 (N_5162,N_2835,N_3997);
or U5163 (N_5163,N_2239,N_3133);
xor U5164 (N_5164,N_3124,N_2864);
and U5165 (N_5165,N_2277,N_2311);
and U5166 (N_5166,N_2620,N_3547);
or U5167 (N_5167,N_2798,N_3393);
nand U5168 (N_5168,N_3081,N_3226);
and U5169 (N_5169,N_2554,N_2904);
or U5170 (N_5170,N_2087,N_3789);
nand U5171 (N_5171,N_2703,N_3912);
and U5172 (N_5172,N_3404,N_2555);
and U5173 (N_5173,N_2403,N_2896);
and U5174 (N_5174,N_2675,N_2436);
nand U5175 (N_5175,N_3116,N_3728);
nand U5176 (N_5176,N_2059,N_2313);
nor U5177 (N_5177,N_2957,N_2011);
nand U5178 (N_5178,N_2238,N_3380);
or U5179 (N_5179,N_2676,N_2204);
nand U5180 (N_5180,N_3888,N_2962);
nor U5181 (N_5181,N_2101,N_3260);
or U5182 (N_5182,N_2142,N_3397);
and U5183 (N_5183,N_3254,N_2388);
or U5184 (N_5184,N_2688,N_2521);
and U5185 (N_5185,N_3118,N_2380);
nor U5186 (N_5186,N_3160,N_3778);
or U5187 (N_5187,N_3113,N_2054);
or U5188 (N_5188,N_2951,N_3650);
and U5189 (N_5189,N_2484,N_3764);
nor U5190 (N_5190,N_3813,N_3595);
nand U5191 (N_5191,N_3076,N_3887);
and U5192 (N_5192,N_2950,N_3219);
or U5193 (N_5193,N_2454,N_3268);
or U5194 (N_5194,N_3394,N_3736);
xnor U5195 (N_5195,N_3999,N_3209);
and U5196 (N_5196,N_3512,N_2590);
or U5197 (N_5197,N_2233,N_3033);
nor U5198 (N_5198,N_2515,N_3111);
nand U5199 (N_5199,N_2251,N_3189);
nor U5200 (N_5200,N_3617,N_2368);
and U5201 (N_5201,N_2622,N_3284);
or U5202 (N_5202,N_3954,N_2084);
and U5203 (N_5203,N_2166,N_3574);
xnor U5204 (N_5204,N_2764,N_2690);
xnor U5205 (N_5205,N_2402,N_2525);
and U5206 (N_5206,N_3490,N_3049);
or U5207 (N_5207,N_3106,N_2829);
nand U5208 (N_5208,N_3498,N_2222);
nand U5209 (N_5209,N_2500,N_2001);
and U5210 (N_5210,N_2431,N_3380);
xor U5211 (N_5211,N_2236,N_3810);
and U5212 (N_5212,N_3341,N_3151);
or U5213 (N_5213,N_3114,N_2034);
and U5214 (N_5214,N_3041,N_3867);
xnor U5215 (N_5215,N_3122,N_3378);
nor U5216 (N_5216,N_3237,N_3055);
xnor U5217 (N_5217,N_2884,N_3927);
nand U5218 (N_5218,N_2205,N_2882);
nand U5219 (N_5219,N_2231,N_2524);
nand U5220 (N_5220,N_3449,N_3452);
and U5221 (N_5221,N_3218,N_3342);
nor U5222 (N_5222,N_2987,N_2994);
or U5223 (N_5223,N_2546,N_3940);
xor U5224 (N_5224,N_2436,N_2658);
or U5225 (N_5225,N_3985,N_3664);
xnor U5226 (N_5226,N_3610,N_3045);
xnor U5227 (N_5227,N_3147,N_3247);
nand U5228 (N_5228,N_3793,N_2128);
nor U5229 (N_5229,N_2569,N_2335);
or U5230 (N_5230,N_3428,N_2843);
and U5231 (N_5231,N_2466,N_2053);
xor U5232 (N_5232,N_3180,N_3532);
nand U5233 (N_5233,N_3414,N_3610);
or U5234 (N_5234,N_2817,N_2774);
and U5235 (N_5235,N_2306,N_2728);
or U5236 (N_5236,N_3448,N_2272);
nand U5237 (N_5237,N_2060,N_3543);
xnor U5238 (N_5238,N_2758,N_2747);
or U5239 (N_5239,N_3287,N_3604);
nand U5240 (N_5240,N_2849,N_3877);
xnor U5241 (N_5241,N_3672,N_3155);
and U5242 (N_5242,N_2376,N_3104);
xor U5243 (N_5243,N_2276,N_2958);
or U5244 (N_5244,N_2249,N_2532);
or U5245 (N_5245,N_3783,N_2585);
xnor U5246 (N_5246,N_3001,N_3515);
xnor U5247 (N_5247,N_3265,N_3491);
nor U5248 (N_5248,N_3950,N_2710);
xnor U5249 (N_5249,N_2028,N_2053);
or U5250 (N_5250,N_2000,N_3052);
nand U5251 (N_5251,N_3012,N_3067);
nor U5252 (N_5252,N_3372,N_3742);
or U5253 (N_5253,N_2170,N_2741);
or U5254 (N_5254,N_3863,N_3827);
and U5255 (N_5255,N_3499,N_2797);
nor U5256 (N_5256,N_3611,N_2570);
xor U5257 (N_5257,N_2686,N_3159);
or U5258 (N_5258,N_2482,N_2101);
nor U5259 (N_5259,N_2249,N_3514);
and U5260 (N_5260,N_2653,N_3927);
or U5261 (N_5261,N_2485,N_3473);
xnor U5262 (N_5262,N_2568,N_2703);
xor U5263 (N_5263,N_2100,N_3816);
or U5264 (N_5264,N_3845,N_2663);
and U5265 (N_5265,N_2353,N_2661);
xnor U5266 (N_5266,N_2337,N_3297);
nand U5267 (N_5267,N_3260,N_2425);
nor U5268 (N_5268,N_2605,N_3600);
nor U5269 (N_5269,N_2226,N_2922);
nand U5270 (N_5270,N_2968,N_2652);
nand U5271 (N_5271,N_3320,N_2385);
nor U5272 (N_5272,N_2548,N_2153);
or U5273 (N_5273,N_3351,N_3180);
nor U5274 (N_5274,N_2272,N_2475);
nand U5275 (N_5275,N_2411,N_2671);
xor U5276 (N_5276,N_3475,N_3677);
or U5277 (N_5277,N_2417,N_3443);
xor U5278 (N_5278,N_2588,N_2373);
nor U5279 (N_5279,N_3482,N_3351);
nor U5280 (N_5280,N_3828,N_2684);
xor U5281 (N_5281,N_2681,N_2922);
or U5282 (N_5282,N_2005,N_3773);
nand U5283 (N_5283,N_3593,N_2330);
nor U5284 (N_5284,N_3873,N_3526);
or U5285 (N_5285,N_3143,N_3560);
and U5286 (N_5286,N_3625,N_3124);
or U5287 (N_5287,N_2573,N_3416);
or U5288 (N_5288,N_2825,N_2636);
and U5289 (N_5289,N_2308,N_2979);
nand U5290 (N_5290,N_3193,N_2228);
nand U5291 (N_5291,N_2563,N_3678);
or U5292 (N_5292,N_2768,N_2450);
nand U5293 (N_5293,N_2753,N_3113);
and U5294 (N_5294,N_3007,N_3728);
or U5295 (N_5295,N_3497,N_2082);
and U5296 (N_5296,N_2753,N_2471);
and U5297 (N_5297,N_3325,N_2878);
and U5298 (N_5298,N_2139,N_3889);
or U5299 (N_5299,N_2471,N_3235);
nand U5300 (N_5300,N_2646,N_3929);
nor U5301 (N_5301,N_3349,N_2179);
nor U5302 (N_5302,N_2788,N_3800);
or U5303 (N_5303,N_3620,N_3866);
xnor U5304 (N_5304,N_2417,N_3891);
or U5305 (N_5305,N_2554,N_2324);
and U5306 (N_5306,N_3160,N_3946);
and U5307 (N_5307,N_2269,N_2745);
xnor U5308 (N_5308,N_2367,N_2681);
nor U5309 (N_5309,N_3806,N_3737);
and U5310 (N_5310,N_2156,N_2771);
nor U5311 (N_5311,N_2245,N_3022);
nor U5312 (N_5312,N_2274,N_3904);
xor U5313 (N_5313,N_3139,N_3472);
nand U5314 (N_5314,N_2342,N_3374);
or U5315 (N_5315,N_3955,N_3055);
xnor U5316 (N_5316,N_3263,N_2750);
nor U5317 (N_5317,N_2099,N_2855);
nand U5318 (N_5318,N_3536,N_2791);
xnor U5319 (N_5319,N_3096,N_3355);
xor U5320 (N_5320,N_3457,N_3430);
nor U5321 (N_5321,N_2818,N_3835);
xnor U5322 (N_5322,N_2804,N_2259);
nor U5323 (N_5323,N_2457,N_2854);
xor U5324 (N_5324,N_3024,N_3085);
nor U5325 (N_5325,N_2087,N_2501);
nand U5326 (N_5326,N_3378,N_2943);
or U5327 (N_5327,N_3227,N_3556);
and U5328 (N_5328,N_3601,N_2202);
nor U5329 (N_5329,N_3117,N_2964);
and U5330 (N_5330,N_2248,N_3685);
nand U5331 (N_5331,N_2087,N_3408);
xor U5332 (N_5332,N_2337,N_3077);
nor U5333 (N_5333,N_2077,N_2270);
nor U5334 (N_5334,N_3377,N_3792);
and U5335 (N_5335,N_3898,N_2723);
or U5336 (N_5336,N_3375,N_2302);
nor U5337 (N_5337,N_3717,N_3958);
or U5338 (N_5338,N_3315,N_2259);
xnor U5339 (N_5339,N_3620,N_3156);
or U5340 (N_5340,N_3349,N_3458);
and U5341 (N_5341,N_2512,N_2426);
and U5342 (N_5342,N_2705,N_3303);
xor U5343 (N_5343,N_2087,N_3070);
and U5344 (N_5344,N_2379,N_3063);
nor U5345 (N_5345,N_2501,N_2972);
nor U5346 (N_5346,N_2620,N_3501);
nand U5347 (N_5347,N_2404,N_2550);
nor U5348 (N_5348,N_2132,N_3530);
xnor U5349 (N_5349,N_3831,N_2810);
nand U5350 (N_5350,N_3862,N_3827);
or U5351 (N_5351,N_3097,N_3539);
nor U5352 (N_5352,N_3174,N_3124);
nor U5353 (N_5353,N_3689,N_2537);
xnor U5354 (N_5354,N_3349,N_2198);
and U5355 (N_5355,N_2267,N_2153);
nand U5356 (N_5356,N_3432,N_2364);
and U5357 (N_5357,N_2651,N_2174);
nor U5358 (N_5358,N_2152,N_3854);
xor U5359 (N_5359,N_3559,N_2702);
and U5360 (N_5360,N_2114,N_3148);
xnor U5361 (N_5361,N_3892,N_3783);
xor U5362 (N_5362,N_3378,N_3388);
xor U5363 (N_5363,N_2077,N_3806);
nand U5364 (N_5364,N_3528,N_2641);
nand U5365 (N_5365,N_2755,N_3900);
nor U5366 (N_5366,N_3993,N_3197);
xor U5367 (N_5367,N_2835,N_2921);
xor U5368 (N_5368,N_2429,N_3896);
nor U5369 (N_5369,N_2115,N_2974);
nor U5370 (N_5370,N_3281,N_2116);
or U5371 (N_5371,N_2881,N_3982);
nand U5372 (N_5372,N_2743,N_3076);
and U5373 (N_5373,N_3540,N_3617);
and U5374 (N_5374,N_2259,N_2230);
or U5375 (N_5375,N_2050,N_3299);
nand U5376 (N_5376,N_3938,N_2920);
and U5377 (N_5377,N_3017,N_3278);
nand U5378 (N_5378,N_3394,N_3016);
or U5379 (N_5379,N_3675,N_2223);
xnor U5380 (N_5380,N_2471,N_2468);
nand U5381 (N_5381,N_3387,N_2813);
and U5382 (N_5382,N_2539,N_3842);
nor U5383 (N_5383,N_2176,N_3950);
or U5384 (N_5384,N_3357,N_2301);
nor U5385 (N_5385,N_2693,N_3528);
nand U5386 (N_5386,N_3556,N_3070);
and U5387 (N_5387,N_2729,N_2933);
or U5388 (N_5388,N_3411,N_3443);
xor U5389 (N_5389,N_2630,N_3495);
nand U5390 (N_5390,N_3932,N_2985);
and U5391 (N_5391,N_2454,N_2742);
nor U5392 (N_5392,N_3207,N_2951);
xor U5393 (N_5393,N_3631,N_2300);
or U5394 (N_5394,N_3866,N_2494);
or U5395 (N_5395,N_3148,N_2720);
and U5396 (N_5396,N_2788,N_2160);
nand U5397 (N_5397,N_2605,N_3439);
nand U5398 (N_5398,N_3982,N_2706);
or U5399 (N_5399,N_2923,N_3672);
nor U5400 (N_5400,N_2550,N_2027);
nor U5401 (N_5401,N_2213,N_2971);
nor U5402 (N_5402,N_2430,N_2354);
or U5403 (N_5403,N_3834,N_2173);
or U5404 (N_5404,N_2050,N_2648);
nand U5405 (N_5405,N_2121,N_2382);
xnor U5406 (N_5406,N_3638,N_3121);
and U5407 (N_5407,N_3767,N_3283);
or U5408 (N_5408,N_2172,N_2926);
nor U5409 (N_5409,N_3373,N_2959);
nand U5410 (N_5410,N_3593,N_2515);
nand U5411 (N_5411,N_2497,N_3297);
and U5412 (N_5412,N_2255,N_2064);
xnor U5413 (N_5413,N_2095,N_3320);
nor U5414 (N_5414,N_2375,N_2798);
and U5415 (N_5415,N_2602,N_3162);
nand U5416 (N_5416,N_3487,N_3438);
nand U5417 (N_5417,N_2303,N_2096);
and U5418 (N_5418,N_3783,N_3682);
or U5419 (N_5419,N_3357,N_3035);
nand U5420 (N_5420,N_2410,N_2780);
xor U5421 (N_5421,N_2966,N_3091);
and U5422 (N_5422,N_2100,N_2385);
nand U5423 (N_5423,N_3837,N_3396);
or U5424 (N_5424,N_3824,N_2185);
xor U5425 (N_5425,N_3244,N_3511);
or U5426 (N_5426,N_2736,N_2035);
and U5427 (N_5427,N_2528,N_3688);
nand U5428 (N_5428,N_3614,N_3031);
or U5429 (N_5429,N_3626,N_2557);
or U5430 (N_5430,N_2591,N_2421);
xnor U5431 (N_5431,N_3092,N_3203);
nand U5432 (N_5432,N_2359,N_2081);
nand U5433 (N_5433,N_2204,N_3141);
nand U5434 (N_5434,N_2894,N_2043);
nor U5435 (N_5435,N_2438,N_3645);
or U5436 (N_5436,N_3547,N_3334);
and U5437 (N_5437,N_2753,N_3727);
nor U5438 (N_5438,N_3280,N_3623);
and U5439 (N_5439,N_2741,N_3300);
nand U5440 (N_5440,N_3814,N_3032);
xnor U5441 (N_5441,N_2235,N_2923);
or U5442 (N_5442,N_3211,N_2140);
or U5443 (N_5443,N_2787,N_3998);
nor U5444 (N_5444,N_2947,N_3295);
or U5445 (N_5445,N_2433,N_2068);
xor U5446 (N_5446,N_2783,N_3565);
and U5447 (N_5447,N_2636,N_2275);
xnor U5448 (N_5448,N_3167,N_2648);
nor U5449 (N_5449,N_3179,N_2265);
nand U5450 (N_5450,N_2994,N_2969);
or U5451 (N_5451,N_2655,N_2772);
nand U5452 (N_5452,N_2660,N_2088);
nor U5453 (N_5453,N_2714,N_3159);
nor U5454 (N_5454,N_2131,N_3964);
nand U5455 (N_5455,N_3365,N_2554);
and U5456 (N_5456,N_3011,N_3569);
and U5457 (N_5457,N_2405,N_3876);
nand U5458 (N_5458,N_2682,N_3494);
or U5459 (N_5459,N_2057,N_2622);
and U5460 (N_5460,N_3399,N_3524);
nor U5461 (N_5461,N_3828,N_2752);
and U5462 (N_5462,N_3598,N_3715);
and U5463 (N_5463,N_3087,N_2753);
or U5464 (N_5464,N_3463,N_2818);
and U5465 (N_5465,N_2876,N_3277);
or U5466 (N_5466,N_2996,N_2401);
xnor U5467 (N_5467,N_3625,N_3395);
xor U5468 (N_5468,N_2064,N_3151);
or U5469 (N_5469,N_2471,N_2687);
nand U5470 (N_5470,N_3648,N_2290);
nor U5471 (N_5471,N_3995,N_3334);
nand U5472 (N_5472,N_3219,N_3577);
xnor U5473 (N_5473,N_3161,N_3917);
or U5474 (N_5474,N_2015,N_3090);
and U5475 (N_5475,N_2896,N_3896);
nand U5476 (N_5476,N_3189,N_2398);
xor U5477 (N_5477,N_3298,N_3202);
nor U5478 (N_5478,N_2770,N_2820);
and U5479 (N_5479,N_2815,N_3094);
and U5480 (N_5480,N_3996,N_2822);
xnor U5481 (N_5481,N_3158,N_2887);
nand U5482 (N_5482,N_3077,N_2078);
xor U5483 (N_5483,N_3882,N_3886);
and U5484 (N_5484,N_2321,N_2060);
xnor U5485 (N_5485,N_2701,N_3735);
nor U5486 (N_5486,N_3288,N_2469);
or U5487 (N_5487,N_3290,N_2214);
or U5488 (N_5488,N_2926,N_3122);
nor U5489 (N_5489,N_3557,N_3883);
xnor U5490 (N_5490,N_3914,N_3601);
or U5491 (N_5491,N_3181,N_2830);
nor U5492 (N_5492,N_3327,N_2435);
xnor U5493 (N_5493,N_3426,N_2578);
or U5494 (N_5494,N_2743,N_3591);
or U5495 (N_5495,N_2980,N_3157);
nor U5496 (N_5496,N_3591,N_2176);
xor U5497 (N_5497,N_2858,N_2442);
xor U5498 (N_5498,N_3248,N_2265);
or U5499 (N_5499,N_3837,N_3380);
nor U5500 (N_5500,N_2803,N_3578);
or U5501 (N_5501,N_3234,N_2967);
and U5502 (N_5502,N_2848,N_3216);
nor U5503 (N_5503,N_2455,N_2986);
xor U5504 (N_5504,N_2722,N_2808);
nand U5505 (N_5505,N_2185,N_2832);
or U5506 (N_5506,N_2099,N_2287);
and U5507 (N_5507,N_2705,N_2617);
and U5508 (N_5508,N_3856,N_3059);
or U5509 (N_5509,N_3192,N_3773);
and U5510 (N_5510,N_2490,N_2778);
nor U5511 (N_5511,N_2998,N_3916);
xnor U5512 (N_5512,N_3152,N_2393);
nor U5513 (N_5513,N_3236,N_3816);
and U5514 (N_5514,N_3860,N_3592);
and U5515 (N_5515,N_2290,N_2022);
nor U5516 (N_5516,N_2157,N_3532);
xor U5517 (N_5517,N_3522,N_2429);
nor U5518 (N_5518,N_2381,N_2202);
and U5519 (N_5519,N_3395,N_2087);
nand U5520 (N_5520,N_2584,N_3036);
xor U5521 (N_5521,N_2272,N_3384);
xnor U5522 (N_5522,N_2863,N_3077);
nand U5523 (N_5523,N_2705,N_3059);
and U5524 (N_5524,N_2606,N_2243);
or U5525 (N_5525,N_3901,N_2720);
or U5526 (N_5526,N_2480,N_3739);
xor U5527 (N_5527,N_3314,N_2047);
nor U5528 (N_5528,N_2180,N_3925);
nor U5529 (N_5529,N_3179,N_2394);
or U5530 (N_5530,N_3944,N_3455);
nand U5531 (N_5531,N_2426,N_3045);
or U5532 (N_5532,N_2973,N_2757);
nand U5533 (N_5533,N_3879,N_2910);
or U5534 (N_5534,N_2286,N_2999);
or U5535 (N_5535,N_2714,N_2502);
and U5536 (N_5536,N_3180,N_3158);
nor U5537 (N_5537,N_2832,N_3945);
or U5538 (N_5538,N_2988,N_2955);
nand U5539 (N_5539,N_2831,N_2887);
nand U5540 (N_5540,N_3593,N_2780);
or U5541 (N_5541,N_3522,N_2116);
xor U5542 (N_5542,N_2114,N_3234);
nor U5543 (N_5543,N_2761,N_2393);
or U5544 (N_5544,N_3653,N_3215);
nand U5545 (N_5545,N_3244,N_2618);
nor U5546 (N_5546,N_2984,N_3157);
and U5547 (N_5547,N_3889,N_3710);
xor U5548 (N_5548,N_2255,N_2167);
and U5549 (N_5549,N_2308,N_3334);
nand U5550 (N_5550,N_2536,N_3445);
and U5551 (N_5551,N_2324,N_2345);
and U5552 (N_5552,N_2715,N_2319);
and U5553 (N_5553,N_2890,N_3344);
and U5554 (N_5554,N_3629,N_3385);
xnor U5555 (N_5555,N_3641,N_3171);
and U5556 (N_5556,N_2755,N_3457);
or U5557 (N_5557,N_3126,N_2915);
xnor U5558 (N_5558,N_2819,N_3629);
xnor U5559 (N_5559,N_2352,N_3826);
xor U5560 (N_5560,N_3153,N_3938);
or U5561 (N_5561,N_2444,N_2217);
nor U5562 (N_5562,N_3802,N_2389);
and U5563 (N_5563,N_2065,N_3774);
and U5564 (N_5564,N_2036,N_2597);
nand U5565 (N_5565,N_2568,N_2767);
xor U5566 (N_5566,N_2352,N_2578);
xnor U5567 (N_5567,N_3240,N_2529);
xnor U5568 (N_5568,N_3491,N_2689);
or U5569 (N_5569,N_3404,N_2574);
nand U5570 (N_5570,N_3637,N_2079);
nand U5571 (N_5571,N_2871,N_3968);
xnor U5572 (N_5572,N_3044,N_2356);
nor U5573 (N_5573,N_3262,N_3212);
or U5574 (N_5574,N_3876,N_3424);
or U5575 (N_5575,N_3261,N_3435);
or U5576 (N_5576,N_2748,N_3108);
and U5577 (N_5577,N_3721,N_2980);
and U5578 (N_5578,N_3638,N_2040);
or U5579 (N_5579,N_3885,N_3688);
nand U5580 (N_5580,N_2577,N_3959);
nand U5581 (N_5581,N_2970,N_3470);
xor U5582 (N_5582,N_3677,N_3420);
nand U5583 (N_5583,N_2208,N_3014);
xor U5584 (N_5584,N_3089,N_2084);
and U5585 (N_5585,N_3423,N_3933);
or U5586 (N_5586,N_2207,N_3716);
xor U5587 (N_5587,N_3110,N_3856);
and U5588 (N_5588,N_3841,N_2209);
nand U5589 (N_5589,N_3825,N_3525);
and U5590 (N_5590,N_2950,N_2002);
or U5591 (N_5591,N_3984,N_3706);
and U5592 (N_5592,N_2938,N_2279);
or U5593 (N_5593,N_2220,N_3197);
nor U5594 (N_5594,N_2976,N_3380);
xnor U5595 (N_5595,N_3892,N_3739);
nand U5596 (N_5596,N_2683,N_2790);
or U5597 (N_5597,N_2961,N_2414);
nor U5598 (N_5598,N_3554,N_3615);
or U5599 (N_5599,N_2382,N_2594);
nand U5600 (N_5600,N_2559,N_2411);
nand U5601 (N_5601,N_2653,N_2459);
nor U5602 (N_5602,N_2817,N_3792);
and U5603 (N_5603,N_3816,N_2498);
nor U5604 (N_5604,N_3322,N_3928);
nand U5605 (N_5605,N_3079,N_3756);
nand U5606 (N_5606,N_3970,N_3150);
and U5607 (N_5607,N_3839,N_2976);
xnor U5608 (N_5608,N_3207,N_3651);
and U5609 (N_5609,N_3903,N_3329);
nor U5610 (N_5610,N_3477,N_3297);
xnor U5611 (N_5611,N_3359,N_3258);
nand U5612 (N_5612,N_2423,N_2473);
xnor U5613 (N_5613,N_2384,N_2826);
xnor U5614 (N_5614,N_3363,N_3310);
nor U5615 (N_5615,N_3824,N_3646);
and U5616 (N_5616,N_3076,N_3118);
nor U5617 (N_5617,N_3389,N_2393);
and U5618 (N_5618,N_2032,N_3085);
nand U5619 (N_5619,N_2926,N_3076);
nor U5620 (N_5620,N_2269,N_3007);
nor U5621 (N_5621,N_3948,N_3906);
or U5622 (N_5622,N_3375,N_3493);
nand U5623 (N_5623,N_2250,N_2435);
nand U5624 (N_5624,N_2168,N_2783);
or U5625 (N_5625,N_3213,N_3963);
xnor U5626 (N_5626,N_2113,N_3160);
or U5627 (N_5627,N_3150,N_2919);
and U5628 (N_5628,N_3261,N_2402);
and U5629 (N_5629,N_3535,N_2503);
nor U5630 (N_5630,N_2475,N_3367);
xnor U5631 (N_5631,N_2244,N_2542);
nor U5632 (N_5632,N_2507,N_3635);
nor U5633 (N_5633,N_3803,N_3920);
xnor U5634 (N_5634,N_2613,N_2402);
or U5635 (N_5635,N_3920,N_3655);
and U5636 (N_5636,N_2407,N_2596);
or U5637 (N_5637,N_3016,N_3419);
xnor U5638 (N_5638,N_3416,N_3327);
nand U5639 (N_5639,N_2365,N_2572);
nand U5640 (N_5640,N_2235,N_3143);
xor U5641 (N_5641,N_3199,N_2400);
and U5642 (N_5642,N_2550,N_2934);
and U5643 (N_5643,N_2565,N_2864);
xnor U5644 (N_5644,N_3464,N_3269);
nor U5645 (N_5645,N_2728,N_2378);
xor U5646 (N_5646,N_3030,N_3808);
and U5647 (N_5647,N_2419,N_2582);
or U5648 (N_5648,N_3717,N_3660);
or U5649 (N_5649,N_2326,N_2985);
xnor U5650 (N_5650,N_2834,N_2610);
and U5651 (N_5651,N_3577,N_3791);
nand U5652 (N_5652,N_2184,N_2251);
nor U5653 (N_5653,N_2863,N_2333);
xor U5654 (N_5654,N_2252,N_2225);
nand U5655 (N_5655,N_2781,N_3861);
nor U5656 (N_5656,N_2937,N_2156);
nor U5657 (N_5657,N_3738,N_2064);
or U5658 (N_5658,N_3909,N_2006);
nor U5659 (N_5659,N_2862,N_2430);
and U5660 (N_5660,N_2438,N_2350);
and U5661 (N_5661,N_2649,N_2312);
nand U5662 (N_5662,N_2751,N_3279);
xnor U5663 (N_5663,N_3754,N_2905);
nand U5664 (N_5664,N_2438,N_3136);
nor U5665 (N_5665,N_2522,N_3498);
xnor U5666 (N_5666,N_2692,N_3185);
or U5667 (N_5667,N_3226,N_2779);
or U5668 (N_5668,N_3916,N_2109);
and U5669 (N_5669,N_2715,N_2038);
nand U5670 (N_5670,N_3036,N_2779);
nand U5671 (N_5671,N_2133,N_2084);
or U5672 (N_5672,N_2063,N_3860);
and U5673 (N_5673,N_3157,N_3551);
nand U5674 (N_5674,N_2533,N_2965);
nor U5675 (N_5675,N_2853,N_2618);
nand U5676 (N_5676,N_2384,N_2999);
xor U5677 (N_5677,N_2904,N_2528);
and U5678 (N_5678,N_2437,N_3523);
nor U5679 (N_5679,N_2265,N_3395);
nand U5680 (N_5680,N_3230,N_2174);
xor U5681 (N_5681,N_3852,N_3510);
nand U5682 (N_5682,N_2381,N_3850);
or U5683 (N_5683,N_3941,N_2272);
nor U5684 (N_5684,N_2335,N_2620);
or U5685 (N_5685,N_2238,N_3041);
xor U5686 (N_5686,N_2614,N_2639);
nand U5687 (N_5687,N_3191,N_3237);
nand U5688 (N_5688,N_3949,N_3767);
or U5689 (N_5689,N_3124,N_2728);
nand U5690 (N_5690,N_2678,N_2661);
and U5691 (N_5691,N_2636,N_3495);
nand U5692 (N_5692,N_2884,N_2034);
or U5693 (N_5693,N_3429,N_2468);
and U5694 (N_5694,N_2800,N_2678);
or U5695 (N_5695,N_2706,N_2663);
or U5696 (N_5696,N_2096,N_3951);
and U5697 (N_5697,N_2988,N_2448);
nor U5698 (N_5698,N_2276,N_2943);
nand U5699 (N_5699,N_2641,N_3805);
nor U5700 (N_5700,N_3747,N_2927);
and U5701 (N_5701,N_2024,N_3546);
and U5702 (N_5702,N_3251,N_2382);
and U5703 (N_5703,N_2410,N_3088);
nand U5704 (N_5704,N_3851,N_3945);
or U5705 (N_5705,N_3998,N_3523);
nor U5706 (N_5706,N_2648,N_3206);
or U5707 (N_5707,N_2340,N_3294);
and U5708 (N_5708,N_3935,N_3938);
nand U5709 (N_5709,N_2094,N_3746);
xor U5710 (N_5710,N_3196,N_2674);
xnor U5711 (N_5711,N_2295,N_2545);
xor U5712 (N_5712,N_3924,N_3274);
nand U5713 (N_5713,N_3390,N_2757);
nand U5714 (N_5714,N_3006,N_3825);
nor U5715 (N_5715,N_3919,N_2280);
and U5716 (N_5716,N_2121,N_3002);
nand U5717 (N_5717,N_2003,N_2307);
nor U5718 (N_5718,N_3098,N_2985);
nor U5719 (N_5719,N_2688,N_3044);
or U5720 (N_5720,N_2092,N_2778);
and U5721 (N_5721,N_2883,N_2473);
or U5722 (N_5722,N_2964,N_2704);
or U5723 (N_5723,N_3447,N_2310);
xor U5724 (N_5724,N_2726,N_3611);
and U5725 (N_5725,N_2305,N_2081);
nand U5726 (N_5726,N_3851,N_2876);
nand U5727 (N_5727,N_2555,N_2960);
xor U5728 (N_5728,N_3533,N_2560);
nand U5729 (N_5729,N_2653,N_2554);
nor U5730 (N_5730,N_3610,N_2261);
nand U5731 (N_5731,N_3124,N_3719);
or U5732 (N_5732,N_2657,N_3617);
nor U5733 (N_5733,N_3640,N_2407);
or U5734 (N_5734,N_2925,N_3143);
and U5735 (N_5735,N_2406,N_3521);
or U5736 (N_5736,N_3625,N_2201);
xnor U5737 (N_5737,N_3291,N_3419);
xnor U5738 (N_5738,N_3369,N_2507);
nor U5739 (N_5739,N_3144,N_2859);
nand U5740 (N_5740,N_3954,N_3196);
or U5741 (N_5741,N_3980,N_3740);
nand U5742 (N_5742,N_3096,N_2318);
or U5743 (N_5743,N_3873,N_2875);
or U5744 (N_5744,N_2634,N_3024);
or U5745 (N_5745,N_2319,N_2760);
nand U5746 (N_5746,N_3900,N_2335);
xor U5747 (N_5747,N_2221,N_2493);
or U5748 (N_5748,N_2072,N_2709);
nor U5749 (N_5749,N_3117,N_3699);
or U5750 (N_5750,N_3121,N_2233);
or U5751 (N_5751,N_3553,N_3385);
and U5752 (N_5752,N_2181,N_2307);
and U5753 (N_5753,N_2494,N_2634);
xor U5754 (N_5754,N_2064,N_3382);
and U5755 (N_5755,N_2356,N_3915);
nor U5756 (N_5756,N_3317,N_2018);
xnor U5757 (N_5757,N_2115,N_3473);
nand U5758 (N_5758,N_3575,N_3526);
nand U5759 (N_5759,N_2436,N_2396);
nand U5760 (N_5760,N_2400,N_2303);
or U5761 (N_5761,N_3522,N_3694);
and U5762 (N_5762,N_2545,N_3609);
and U5763 (N_5763,N_3664,N_3061);
or U5764 (N_5764,N_2682,N_2647);
xor U5765 (N_5765,N_3903,N_2723);
or U5766 (N_5766,N_3189,N_2079);
and U5767 (N_5767,N_3300,N_2564);
and U5768 (N_5768,N_2238,N_2469);
or U5769 (N_5769,N_3826,N_2723);
and U5770 (N_5770,N_3712,N_3310);
xor U5771 (N_5771,N_3232,N_3518);
or U5772 (N_5772,N_3092,N_3926);
nor U5773 (N_5773,N_3046,N_3593);
nand U5774 (N_5774,N_2814,N_2319);
or U5775 (N_5775,N_3376,N_2303);
and U5776 (N_5776,N_2539,N_3387);
and U5777 (N_5777,N_2613,N_2835);
xnor U5778 (N_5778,N_2682,N_2098);
xor U5779 (N_5779,N_3282,N_3846);
xnor U5780 (N_5780,N_3919,N_3369);
nor U5781 (N_5781,N_2063,N_2538);
or U5782 (N_5782,N_2707,N_3778);
nand U5783 (N_5783,N_3023,N_2350);
nor U5784 (N_5784,N_2046,N_3289);
or U5785 (N_5785,N_2373,N_2247);
nand U5786 (N_5786,N_2110,N_2938);
nor U5787 (N_5787,N_2925,N_2331);
nor U5788 (N_5788,N_3254,N_2932);
nand U5789 (N_5789,N_2981,N_2496);
nand U5790 (N_5790,N_3047,N_3081);
or U5791 (N_5791,N_3663,N_2885);
or U5792 (N_5792,N_3371,N_3747);
nor U5793 (N_5793,N_2197,N_3511);
or U5794 (N_5794,N_2547,N_3771);
nand U5795 (N_5795,N_2803,N_3728);
or U5796 (N_5796,N_3306,N_2030);
xor U5797 (N_5797,N_3211,N_2927);
nor U5798 (N_5798,N_2528,N_3112);
xor U5799 (N_5799,N_3562,N_2185);
xnor U5800 (N_5800,N_3584,N_3017);
and U5801 (N_5801,N_3359,N_2723);
nand U5802 (N_5802,N_3095,N_2133);
xnor U5803 (N_5803,N_3692,N_2994);
and U5804 (N_5804,N_2772,N_3207);
xnor U5805 (N_5805,N_3178,N_3188);
nor U5806 (N_5806,N_2396,N_2515);
nor U5807 (N_5807,N_2753,N_2581);
nand U5808 (N_5808,N_2460,N_3765);
xnor U5809 (N_5809,N_3179,N_3340);
nor U5810 (N_5810,N_2236,N_2429);
xnor U5811 (N_5811,N_3899,N_2978);
nand U5812 (N_5812,N_3243,N_3854);
nand U5813 (N_5813,N_2647,N_3045);
nor U5814 (N_5814,N_2526,N_2771);
nand U5815 (N_5815,N_2876,N_2468);
and U5816 (N_5816,N_2210,N_3344);
xnor U5817 (N_5817,N_3389,N_3274);
or U5818 (N_5818,N_2321,N_2879);
xnor U5819 (N_5819,N_2034,N_3606);
nor U5820 (N_5820,N_2979,N_3853);
and U5821 (N_5821,N_3248,N_3271);
nand U5822 (N_5822,N_3351,N_3446);
nand U5823 (N_5823,N_3741,N_3740);
xor U5824 (N_5824,N_3184,N_3239);
nor U5825 (N_5825,N_2817,N_2955);
nor U5826 (N_5826,N_3423,N_3141);
nor U5827 (N_5827,N_3630,N_3927);
xnor U5828 (N_5828,N_3619,N_2132);
nor U5829 (N_5829,N_3694,N_2636);
and U5830 (N_5830,N_2168,N_2508);
nor U5831 (N_5831,N_3835,N_2407);
and U5832 (N_5832,N_2373,N_2161);
xnor U5833 (N_5833,N_3942,N_2878);
xor U5834 (N_5834,N_2477,N_2118);
xor U5835 (N_5835,N_2616,N_2889);
xor U5836 (N_5836,N_2234,N_3370);
and U5837 (N_5837,N_3990,N_3355);
nand U5838 (N_5838,N_2406,N_3906);
xor U5839 (N_5839,N_2376,N_2021);
xnor U5840 (N_5840,N_3854,N_3597);
nor U5841 (N_5841,N_3151,N_2494);
nor U5842 (N_5842,N_3193,N_2274);
nor U5843 (N_5843,N_3189,N_3074);
nor U5844 (N_5844,N_3570,N_2490);
and U5845 (N_5845,N_2425,N_3893);
nand U5846 (N_5846,N_3162,N_3243);
nand U5847 (N_5847,N_2363,N_3765);
xor U5848 (N_5848,N_3398,N_2707);
xnor U5849 (N_5849,N_3974,N_2190);
and U5850 (N_5850,N_3256,N_3333);
xor U5851 (N_5851,N_3909,N_3645);
and U5852 (N_5852,N_2174,N_2875);
xor U5853 (N_5853,N_3751,N_2146);
xor U5854 (N_5854,N_3313,N_3675);
xnor U5855 (N_5855,N_3132,N_3756);
nor U5856 (N_5856,N_2690,N_3358);
or U5857 (N_5857,N_2822,N_2137);
nand U5858 (N_5858,N_3511,N_3773);
xnor U5859 (N_5859,N_2882,N_3127);
nor U5860 (N_5860,N_2288,N_3337);
nor U5861 (N_5861,N_2685,N_3942);
nand U5862 (N_5862,N_3320,N_2694);
and U5863 (N_5863,N_2060,N_2807);
and U5864 (N_5864,N_2542,N_3740);
xnor U5865 (N_5865,N_3808,N_3922);
nor U5866 (N_5866,N_2221,N_2905);
nor U5867 (N_5867,N_2455,N_2985);
or U5868 (N_5868,N_2708,N_2690);
or U5869 (N_5869,N_2131,N_2774);
xnor U5870 (N_5870,N_3067,N_3934);
and U5871 (N_5871,N_2979,N_3973);
nor U5872 (N_5872,N_3186,N_2008);
xor U5873 (N_5873,N_3573,N_3062);
nor U5874 (N_5874,N_3074,N_3503);
xor U5875 (N_5875,N_2381,N_2920);
nand U5876 (N_5876,N_3138,N_2888);
xor U5877 (N_5877,N_3750,N_3141);
or U5878 (N_5878,N_3520,N_2560);
nand U5879 (N_5879,N_2774,N_2809);
nor U5880 (N_5880,N_2380,N_3233);
and U5881 (N_5881,N_3456,N_2735);
nor U5882 (N_5882,N_3622,N_2742);
xor U5883 (N_5883,N_2461,N_2185);
or U5884 (N_5884,N_3564,N_2665);
and U5885 (N_5885,N_2539,N_2147);
nand U5886 (N_5886,N_2973,N_3563);
or U5887 (N_5887,N_3379,N_3844);
nor U5888 (N_5888,N_2555,N_2485);
and U5889 (N_5889,N_2943,N_3825);
nor U5890 (N_5890,N_3585,N_2412);
nand U5891 (N_5891,N_2957,N_3487);
nand U5892 (N_5892,N_3437,N_2431);
xnor U5893 (N_5893,N_2855,N_2525);
and U5894 (N_5894,N_3486,N_2799);
or U5895 (N_5895,N_3015,N_2313);
xor U5896 (N_5896,N_2370,N_2630);
and U5897 (N_5897,N_2231,N_2740);
or U5898 (N_5898,N_3287,N_2474);
xor U5899 (N_5899,N_2013,N_2362);
nor U5900 (N_5900,N_3188,N_2548);
xor U5901 (N_5901,N_2426,N_2179);
nor U5902 (N_5902,N_3732,N_2710);
nand U5903 (N_5903,N_3734,N_2339);
nor U5904 (N_5904,N_2694,N_2070);
nor U5905 (N_5905,N_2778,N_2444);
nor U5906 (N_5906,N_2659,N_3566);
nand U5907 (N_5907,N_2442,N_3289);
nor U5908 (N_5908,N_2814,N_3109);
nor U5909 (N_5909,N_2102,N_2197);
and U5910 (N_5910,N_2782,N_2841);
and U5911 (N_5911,N_2567,N_2017);
nor U5912 (N_5912,N_2848,N_3791);
or U5913 (N_5913,N_3828,N_2584);
and U5914 (N_5914,N_3458,N_2687);
and U5915 (N_5915,N_3875,N_3810);
nand U5916 (N_5916,N_2431,N_3036);
xor U5917 (N_5917,N_3827,N_3134);
or U5918 (N_5918,N_2100,N_2057);
or U5919 (N_5919,N_3469,N_3276);
xor U5920 (N_5920,N_3532,N_3047);
nor U5921 (N_5921,N_2596,N_2314);
and U5922 (N_5922,N_2110,N_2621);
xnor U5923 (N_5923,N_3805,N_3878);
or U5924 (N_5924,N_3667,N_2467);
nor U5925 (N_5925,N_2697,N_3776);
or U5926 (N_5926,N_2772,N_2205);
and U5927 (N_5927,N_2174,N_2097);
nand U5928 (N_5928,N_2998,N_2867);
nor U5929 (N_5929,N_3958,N_2742);
nand U5930 (N_5930,N_3783,N_3828);
or U5931 (N_5931,N_3588,N_2883);
nor U5932 (N_5932,N_2943,N_3469);
nand U5933 (N_5933,N_2687,N_2426);
and U5934 (N_5934,N_3039,N_3987);
nand U5935 (N_5935,N_2965,N_2861);
nor U5936 (N_5936,N_3808,N_2357);
or U5937 (N_5937,N_2889,N_3114);
and U5938 (N_5938,N_2259,N_3277);
or U5939 (N_5939,N_2762,N_3427);
and U5940 (N_5940,N_2557,N_2835);
nand U5941 (N_5941,N_3877,N_3999);
or U5942 (N_5942,N_2755,N_2175);
and U5943 (N_5943,N_2939,N_3152);
nor U5944 (N_5944,N_2837,N_2158);
or U5945 (N_5945,N_3318,N_3935);
nand U5946 (N_5946,N_3884,N_3619);
nand U5947 (N_5947,N_3850,N_2881);
or U5948 (N_5948,N_2799,N_2738);
xor U5949 (N_5949,N_3851,N_2576);
or U5950 (N_5950,N_2707,N_3377);
xnor U5951 (N_5951,N_3664,N_2729);
or U5952 (N_5952,N_3511,N_2601);
xor U5953 (N_5953,N_2197,N_2999);
xnor U5954 (N_5954,N_3097,N_3025);
or U5955 (N_5955,N_2908,N_3125);
or U5956 (N_5956,N_2926,N_3352);
xnor U5957 (N_5957,N_3113,N_3095);
nand U5958 (N_5958,N_2499,N_2404);
or U5959 (N_5959,N_2520,N_3895);
or U5960 (N_5960,N_2493,N_2022);
xor U5961 (N_5961,N_2774,N_3082);
nor U5962 (N_5962,N_2218,N_3203);
nor U5963 (N_5963,N_3595,N_2211);
nand U5964 (N_5964,N_3705,N_3674);
and U5965 (N_5965,N_2454,N_3752);
or U5966 (N_5966,N_3889,N_3354);
nor U5967 (N_5967,N_2894,N_3849);
and U5968 (N_5968,N_3811,N_3494);
nand U5969 (N_5969,N_3455,N_3120);
nand U5970 (N_5970,N_2276,N_3075);
nand U5971 (N_5971,N_2524,N_3981);
or U5972 (N_5972,N_3460,N_3603);
nor U5973 (N_5973,N_2747,N_3307);
and U5974 (N_5974,N_3059,N_2844);
or U5975 (N_5975,N_2812,N_3269);
and U5976 (N_5976,N_3896,N_3796);
xor U5977 (N_5977,N_3105,N_2335);
nor U5978 (N_5978,N_2137,N_3111);
nor U5979 (N_5979,N_2059,N_3284);
and U5980 (N_5980,N_2679,N_2865);
nor U5981 (N_5981,N_2648,N_2324);
nand U5982 (N_5982,N_2644,N_3084);
or U5983 (N_5983,N_3221,N_2754);
xnor U5984 (N_5984,N_2347,N_2994);
and U5985 (N_5985,N_2484,N_2022);
xor U5986 (N_5986,N_2089,N_3194);
nand U5987 (N_5987,N_2991,N_2418);
nand U5988 (N_5988,N_3999,N_3738);
or U5989 (N_5989,N_2146,N_3316);
nand U5990 (N_5990,N_2917,N_3944);
xor U5991 (N_5991,N_3948,N_2138);
nand U5992 (N_5992,N_2558,N_3668);
nor U5993 (N_5993,N_3622,N_3659);
nor U5994 (N_5994,N_2246,N_2479);
and U5995 (N_5995,N_3334,N_2093);
or U5996 (N_5996,N_3472,N_2246);
xnor U5997 (N_5997,N_3982,N_3780);
or U5998 (N_5998,N_2154,N_3571);
or U5999 (N_5999,N_3497,N_2195);
and U6000 (N_6000,N_4904,N_4571);
or U6001 (N_6001,N_4573,N_5995);
nand U6002 (N_6002,N_4444,N_5348);
nand U6003 (N_6003,N_5085,N_4323);
nor U6004 (N_6004,N_5349,N_5471);
xor U6005 (N_6005,N_4868,N_5793);
and U6006 (N_6006,N_5087,N_5785);
nand U6007 (N_6007,N_4273,N_5727);
nand U6008 (N_6008,N_4471,N_4024);
xor U6009 (N_6009,N_4641,N_5812);
xnor U6010 (N_6010,N_4971,N_5177);
nor U6011 (N_6011,N_5514,N_5998);
xor U6012 (N_6012,N_5126,N_4239);
nor U6013 (N_6013,N_5970,N_4330);
and U6014 (N_6014,N_5778,N_4990);
xor U6015 (N_6015,N_4418,N_5212);
nor U6016 (N_6016,N_4317,N_5508);
xnor U6017 (N_6017,N_4059,N_4790);
nand U6018 (N_6018,N_5066,N_5566);
xnor U6019 (N_6019,N_4335,N_5516);
and U6020 (N_6020,N_5927,N_5216);
nand U6021 (N_6021,N_5930,N_4111);
or U6022 (N_6022,N_4257,N_5546);
xnor U6023 (N_6023,N_5574,N_5284);
and U6024 (N_6024,N_4823,N_4566);
nor U6025 (N_6025,N_4159,N_5657);
or U6026 (N_6026,N_5338,N_4707);
nand U6027 (N_6027,N_4163,N_4483);
and U6028 (N_6028,N_5450,N_5015);
or U6029 (N_6029,N_5726,N_5773);
nor U6030 (N_6030,N_4120,N_4093);
or U6031 (N_6031,N_4950,N_4071);
or U6032 (N_6032,N_4194,N_5115);
and U6033 (N_6033,N_5913,N_5867);
or U6034 (N_6034,N_5013,N_5201);
xnor U6035 (N_6035,N_5491,N_5571);
or U6036 (N_6036,N_5905,N_4073);
nand U6037 (N_6037,N_5709,N_5360);
xnor U6038 (N_6038,N_4352,N_5889);
nor U6039 (N_6039,N_4495,N_4425);
nor U6040 (N_6040,N_5440,N_4067);
nand U6041 (N_6041,N_4396,N_5534);
nand U6042 (N_6042,N_4362,N_5781);
and U6043 (N_6043,N_4388,N_5005);
nor U6044 (N_6044,N_4004,N_4781);
nand U6045 (N_6045,N_4989,N_5277);
or U6046 (N_6046,N_5044,N_5073);
nor U6047 (N_6047,N_5553,N_4786);
xor U6048 (N_6048,N_4065,N_4215);
or U6049 (N_6049,N_5486,N_4162);
and U6050 (N_6050,N_5819,N_5313);
nand U6051 (N_6051,N_5267,N_4360);
or U6052 (N_6052,N_5862,N_4896);
and U6053 (N_6053,N_5039,N_5760);
nand U6054 (N_6054,N_5092,N_5842);
or U6055 (N_6055,N_4520,N_4445);
xnor U6056 (N_6056,N_4910,N_4898);
nand U6057 (N_6057,N_5231,N_5679);
nor U6058 (N_6058,N_5991,N_5869);
or U6059 (N_6059,N_5958,N_4176);
xor U6060 (N_6060,N_4985,N_5114);
xor U6061 (N_6061,N_4413,N_5499);
nor U6062 (N_6062,N_5725,N_5462);
or U6063 (N_6063,N_4730,N_5170);
nor U6064 (N_6064,N_5314,N_4166);
nor U6065 (N_6065,N_4408,N_4490);
or U6066 (N_6066,N_5703,N_5558);
or U6067 (N_6067,N_5274,N_5503);
nand U6068 (N_6068,N_4652,N_5856);
nor U6069 (N_6069,N_4694,N_5505);
nand U6070 (N_6070,N_4683,N_4438);
nor U6071 (N_6071,N_5208,N_5756);
nand U6072 (N_6072,N_5433,N_5006);
or U6073 (N_6073,N_4554,N_4243);
or U6074 (N_6074,N_4563,N_4959);
nor U6075 (N_6075,N_4552,N_4881);
or U6076 (N_6076,N_4010,N_4252);
xnor U6077 (N_6077,N_5506,N_4502);
and U6078 (N_6078,N_4091,N_4744);
or U6079 (N_6079,N_5938,N_5003);
nand U6080 (N_6080,N_4969,N_4605);
and U6081 (N_6081,N_5105,N_5149);
nor U6082 (N_6082,N_5630,N_5384);
and U6083 (N_6083,N_5780,N_5899);
nand U6084 (N_6084,N_4801,N_5838);
nand U6085 (N_6085,N_5108,N_5205);
nor U6086 (N_6086,N_5189,N_4721);
nor U6087 (N_6087,N_4521,N_5960);
or U6088 (N_6088,N_4003,N_5064);
xor U6089 (N_6089,N_4364,N_5861);
and U6090 (N_6090,N_4871,N_5653);
or U6091 (N_6091,N_5366,N_4991);
nor U6092 (N_6092,N_5548,N_5902);
or U6093 (N_6093,N_5145,N_4556);
and U6094 (N_6094,N_4633,N_5391);
and U6095 (N_6095,N_4015,N_4079);
nand U6096 (N_6096,N_4547,N_4232);
nand U6097 (N_6097,N_4347,N_4892);
xnor U6098 (N_6098,N_4443,N_5196);
nor U6099 (N_6099,N_4596,N_4285);
xor U6100 (N_6100,N_4442,N_4642);
nand U6101 (N_6101,N_4584,N_4157);
nor U6102 (N_6102,N_5102,N_4706);
xor U6103 (N_6103,N_4934,N_5501);
or U6104 (N_6104,N_5786,N_5569);
or U6105 (N_6105,N_4979,N_4765);
nand U6106 (N_6106,N_5772,N_5042);
xor U6107 (N_6107,N_4929,N_4837);
and U6108 (N_6108,N_5833,N_4283);
nor U6109 (N_6109,N_4265,N_5178);
nand U6110 (N_6110,N_4613,N_4282);
xnor U6111 (N_6111,N_4245,N_5831);
nand U6112 (N_6112,N_5748,N_4307);
xor U6113 (N_6113,N_5129,N_5376);
and U6114 (N_6114,N_4489,N_4378);
or U6115 (N_6115,N_5155,N_4462);
or U6116 (N_6116,N_5942,N_4729);
nor U6117 (N_6117,N_5174,N_5230);
nand U6118 (N_6118,N_4090,N_5853);
nor U6119 (N_6119,N_5561,N_4623);
and U6120 (N_6120,N_4419,N_5002);
xnor U6121 (N_6121,N_4296,N_5879);
nor U6122 (N_6122,N_4062,N_5807);
and U6123 (N_6123,N_4716,N_4710);
and U6124 (N_6124,N_4133,N_4741);
nor U6125 (N_6125,N_4855,N_4188);
and U6126 (N_6126,N_4274,N_5148);
and U6127 (N_6127,N_4536,N_5487);
or U6128 (N_6128,N_4369,N_5575);
and U6129 (N_6129,N_4937,N_4263);
or U6130 (N_6130,N_4873,N_5568);
nor U6131 (N_6131,N_5700,N_4535);
nor U6132 (N_6132,N_5962,N_4705);
or U6133 (N_6133,N_5413,N_4349);
and U6134 (N_6134,N_4545,N_5482);
nor U6135 (N_6135,N_5556,N_5400);
and U6136 (N_6136,N_5636,N_5083);
and U6137 (N_6137,N_4051,N_4621);
nand U6138 (N_6138,N_5969,N_5020);
nor U6139 (N_6139,N_4280,N_4509);
nand U6140 (N_6140,N_4504,N_5410);
and U6141 (N_6141,N_5635,N_5454);
nand U6142 (N_6142,N_5933,N_5398);
and U6143 (N_6143,N_4875,N_5086);
nor U6144 (N_6144,N_5164,N_4175);
and U6145 (N_6145,N_4465,N_4410);
nor U6146 (N_6146,N_5300,N_5423);
nor U6147 (N_6147,N_5891,N_5967);
xnor U6148 (N_6148,N_4591,N_5791);
nand U6149 (N_6149,N_5478,N_5359);
or U6150 (N_6150,N_5881,N_5870);
nor U6151 (N_6151,N_4049,N_5301);
and U6152 (N_6152,N_5077,N_4763);
xnor U6153 (N_6153,N_4619,N_5777);
nor U6154 (N_6154,N_5874,N_4013);
and U6155 (N_6155,N_4261,N_4310);
nand U6156 (N_6156,N_5744,N_4997);
xnor U6157 (N_6157,N_4412,N_5082);
xor U6158 (N_6158,N_4662,N_5517);
or U6159 (N_6159,N_4774,N_5993);
nand U6160 (N_6160,N_4519,N_5522);
nand U6161 (N_6161,N_5597,N_4286);
or U6162 (N_6162,N_5934,N_5612);
xor U6163 (N_6163,N_5901,N_4397);
nand U6164 (N_6164,N_5587,N_4686);
nand U6165 (N_6165,N_4404,N_5183);
xor U6166 (N_6166,N_4912,N_5715);
nor U6167 (N_6167,N_4850,N_4788);
nor U6168 (N_6168,N_5334,N_4382);
or U6169 (N_6169,N_4319,N_4271);
nor U6170 (N_6170,N_4949,N_5627);
and U6171 (N_6171,N_4551,N_4451);
xor U6172 (N_6172,N_4034,N_5695);
nand U6173 (N_6173,N_4544,N_5303);
nand U6174 (N_6174,N_5792,N_4860);
nor U6175 (N_6175,N_5661,N_5676);
or U6176 (N_6176,N_4754,N_4312);
and U6177 (N_6177,N_4513,N_4399);
or U6178 (N_6178,N_4085,N_5908);
and U6179 (N_6179,N_4758,N_5437);
nor U6180 (N_6180,N_5825,N_5882);
nand U6181 (N_6181,N_4210,N_4316);
nand U6182 (N_6182,N_5296,N_4935);
xnor U6183 (N_6183,N_5974,N_4909);
or U6184 (N_6184,N_5062,N_5428);
and U6185 (N_6185,N_4607,N_5886);
or U6186 (N_6186,N_4759,N_5733);
nor U6187 (N_6187,N_4485,N_4262);
nand U6188 (N_6188,N_5241,N_5917);
nand U6189 (N_6189,N_4344,N_4392);
nor U6190 (N_6190,N_4762,N_4432);
nand U6191 (N_6191,N_5918,N_5751);
xnor U6192 (N_6192,N_4129,N_4039);
xnor U6193 (N_6193,N_5139,N_5144);
xnor U6194 (N_6194,N_5452,N_5382);
nand U6195 (N_6195,N_4200,N_4919);
nand U6196 (N_6196,N_5670,N_4588);
nor U6197 (N_6197,N_4565,N_5146);
nand U6198 (N_6198,N_4576,N_4427);
nand U6199 (N_6199,N_4191,N_5288);
nand U6200 (N_6200,N_5147,N_4528);
or U6201 (N_6201,N_5099,N_4785);
or U6202 (N_6202,N_4831,N_5941);
nand U6203 (N_6203,N_5192,N_5477);
nor U6204 (N_6204,N_4944,N_5841);
and U6205 (N_6205,N_5061,N_5112);
or U6206 (N_6206,N_5010,N_5684);
nor U6207 (N_6207,N_5816,N_5541);
or U6208 (N_6208,N_4530,N_5403);
nor U6209 (N_6209,N_5065,N_5690);
nor U6210 (N_6210,N_4632,N_4247);
or U6211 (N_6211,N_4322,N_4858);
xor U6212 (N_6212,N_5463,N_5798);
nor U6213 (N_6213,N_5260,N_5426);
or U6214 (N_6214,N_5762,N_5213);
xnor U6215 (N_6215,N_4231,N_5949);
and U6216 (N_6216,N_5176,N_4724);
or U6217 (N_6217,N_5988,N_4911);
or U6218 (N_6218,N_5181,N_4301);
nor U6219 (N_6219,N_4685,N_5321);
nor U6220 (N_6220,N_5855,N_4250);
or U6221 (N_6221,N_5259,N_5362);
xnor U6222 (N_6222,N_5240,N_5909);
and U6223 (N_6223,N_5127,N_5312);
and U6224 (N_6224,N_5672,N_4830);
xor U6225 (N_6225,N_5417,N_4383);
nand U6226 (N_6226,N_5251,N_5686);
and U6227 (N_6227,N_4776,N_4030);
xnor U6228 (N_6228,N_4720,N_4279);
or U6229 (N_6229,N_4867,N_4928);
nand U6230 (N_6230,N_5776,N_5666);
or U6231 (N_6231,N_5030,N_4077);
nand U6232 (N_6232,N_5675,N_5134);
nor U6233 (N_6233,N_5716,N_4311);
xnor U6234 (N_6234,N_4506,N_5219);
xor U6235 (N_6235,N_4201,N_4154);
nor U6236 (N_6236,N_5957,N_4204);
and U6237 (N_6237,N_5734,N_5894);
and U6238 (N_6238,N_5973,N_4138);
nor U6239 (N_6239,N_4165,N_4784);
nor U6240 (N_6240,N_5641,N_5950);
xor U6241 (N_6241,N_5720,N_5782);
xor U6242 (N_6242,N_5797,N_4075);
or U6243 (N_6243,N_4006,N_5618);
nand U6244 (N_6244,N_4488,N_4821);
xnor U6245 (N_6245,N_5591,N_5947);
nor U6246 (N_6246,N_4518,N_5775);
xnor U6247 (N_6247,N_4648,N_4113);
or U6248 (N_6248,N_5677,N_4523);
nor U6249 (N_6249,N_4818,N_4052);
xor U6250 (N_6250,N_4532,N_5755);
nand U6251 (N_6251,N_4481,N_5943);
and U6252 (N_6252,N_5451,N_4604);
nor U6253 (N_6253,N_4476,N_5429);
xnor U6254 (N_6254,N_5570,N_4167);
or U6255 (N_6255,N_5784,N_4844);
nor U6256 (N_6256,N_5954,N_5788);
and U6257 (N_6257,N_4889,N_5502);
or U6258 (N_6258,N_4691,N_4853);
or U6259 (N_6259,N_5399,N_5924);
xnor U6260 (N_6260,N_4331,N_4223);
xor U6261 (N_6261,N_5693,N_5158);
xnor U6262 (N_6262,N_4186,N_5204);
and U6263 (N_6263,N_4738,N_5848);
or U6264 (N_6264,N_5252,N_4233);
or U6265 (N_6265,N_4696,N_4882);
nor U6266 (N_6266,N_4125,N_5154);
nand U6267 (N_6267,N_5560,N_4149);
and U6268 (N_6268,N_5054,N_4346);
nand U6269 (N_6269,N_5774,N_5804);
nor U6270 (N_6270,N_5713,N_4760);
and U6271 (N_6271,N_5536,N_5436);
xnor U6272 (N_6272,N_5904,N_5826);
nor U6273 (N_6273,N_5047,N_5122);
and U6274 (N_6274,N_4647,N_5352);
or U6275 (N_6275,N_4241,N_5735);
and U6276 (N_6276,N_4592,N_4491);
and U6277 (N_6277,N_5599,N_5538);
nand U6278 (N_6278,N_5465,N_4514);
xor U6279 (N_6279,N_5221,N_5070);
nand U6280 (N_6280,N_4893,N_4766);
or U6281 (N_6281,N_4127,N_5717);
and U6282 (N_6282,N_4505,N_5868);
xor U6283 (N_6283,N_4865,N_4612);
nor U6284 (N_6284,N_5585,N_5787);
or U6285 (N_6285,N_5320,N_5658);
xnor U6286 (N_6286,N_4297,N_4456);
nand U6287 (N_6287,N_5012,N_4208);
nor U6288 (N_6288,N_4816,N_4468);
and U6289 (N_6289,N_4925,N_5443);
nor U6290 (N_6290,N_4862,N_4742);
xor U6291 (N_6291,N_4812,N_5238);
xor U6292 (N_6292,N_5632,N_5009);
nand U6293 (N_6293,N_4531,N_4040);
xnor U6294 (N_6294,N_4938,N_4511);
xnor U6295 (N_6295,N_5202,N_4081);
nor U6296 (N_6296,N_4423,N_5237);
and U6297 (N_6297,N_5235,N_4048);
and U6298 (N_6298,N_5997,N_4061);
xnor U6299 (N_6299,N_4022,N_4190);
nor U6300 (N_6300,N_4680,N_5014);
and U6301 (N_6301,N_4601,N_4731);
nand U6302 (N_6302,N_4439,N_5691);
and U6303 (N_6303,N_5412,N_4883);
xnor U6304 (N_6304,N_5416,N_4042);
nor U6305 (N_6305,N_4338,N_4735);
or U6306 (N_6306,N_5628,N_5515);
nand U6307 (N_6307,N_5509,N_4224);
xor U6308 (N_6308,N_4209,N_5031);
xor U6309 (N_6309,N_4849,N_4541);
and U6310 (N_6310,N_5959,N_4747);
nand U6311 (N_6311,N_4666,N_5222);
xnor U6312 (N_6312,N_4214,N_5393);
and U6313 (N_6313,N_4320,N_4023);
and U6314 (N_6314,N_4975,N_5381);
xor U6315 (N_6315,N_4230,N_5101);
nand U6316 (N_6316,N_4597,N_5718);
and U6317 (N_6317,N_4060,N_4089);
or U6318 (N_6318,N_4082,N_5165);
nor U6319 (N_6319,N_5660,N_5021);
nand U6320 (N_6320,N_4140,N_4806);
and U6321 (N_6321,N_4074,N_5863);
and U6322 (N_6322,N_5298,N_4318);
nor U6323 (N_6323,N_5912,N_5888);
or U6324 (N_6324,N_5371,N_4645);
or U6325 (N_6325,N_5810,N_5866);
nand U6326 (N_6326,N_5109,N_5217);
or U6327 (N_6327,N_4288,N_4907);
or U6328 (N_6328,N_5493,N_4072);
nand U6329 (N_6329,N_4562,N_4585);
and U6330 (N_6330,N_4945,N_4328);
xnor U6331 (N_6331,N_4764,N_4834);
xnor U6332 (N_6332,N_5964,N_4473);
nor U6333 (N_6333,N_5769,N_5581);
and U6334 (N_6334,N_5851,N_4461);
or U6335 (N_6335,N_4259,N_4863);
or U6336 (N_6336,N_4646,N_5602);
nand U6337 (N_6337,N_5152,N_5357);
nor U6338 (N_6338,N_5479,N_4942);
or U6339 (N_6339,N_4007,N_4906);
and U6340 (N_6340,N_5318,N_5601);
and U6341 (N_6341,N_4102,N_5837);
nand U6342 (N_6342,N_5552,N_4792);
nor U6343 (N_6343,N_5453,N_5223);
nor U6344 (N_6344,N_5840,N_5186);
nor U6345 (N_6345,N_4527,N_4580);
or U6346 (N_6346,N_5759,N_4508);
xor U6347 (N_6347,N_5519,N_5307);
or U6348 (N_6348,N_4824,N_5405);
or U6349 (N_6349,N_5972,N_4510);
nand U6350 (N_6350,N_4430,N_5537);
and U6351 (N_6351,N_5681,N_4128);
and U6352 (N_6352,N_4878,N_4248);
xor U6353 (N_6353,N_5771,N_5871);
nand U6354 (N_6354,N_4044,N_4832);
and U6355 (N_6355,N_5642,N_5704);
and U6356 (N_6356,N_4570,N_4417);
nor U6357 (N_6357,N_5072,N_4943);
and U6358 (N_6358,N_5282,N_4001);
nor U6359 (N_6359,N_5276,N_4973);
or U6360 (N_6360,N_5119,N_5008);
nor U6361 (N_6361,N_5257,N_4953);
nor U6362 (N_6362,N_5940,N_5356);
and U6363 (N_6363,N_5374,N_4630);
or U6364 (N_6364,N_4579,N_4558);
nor U6365 (N_6365,N_5944,N_5038);
and U6366 (N_6366,N_4936,N_4926);
nor U6367 (N_6367,N_4032,N_4092);
and U6368 (N_6368,N_5996,N_4054);
nor U6369 (N_6369,N_4284,N_4105);
and U6370 (N_6370,N_5233,N_4228);
nand U6371 (N_6371,N_4329,N_4679);
and U6372 (N_6372,N_5279,N_4045);
and U6373 (N_6373,N_4711,N_4422);
or U6374 (N_6374,N_5422,N_4238);
xor U6375 (N_6375,N_4933,N_4891);
xnor U6376 (N_6376,N_5402,N_5929);
nor U6377 (N_6377,N_5449,N_4698);
or U6378 (N_6378,N_4315,N_4761);
or U6379 (N_6379,N_4857,N_5339);
xnor U6380 (N_6380,N_4804,N_4428);
xnor U6381 (N_6381,N_4314,N_4304);
nor U6382 (N_6382,N_5652,N_5169);
or U6383 (N_6383,N_5093,N_5689);
nor U6384 (N_6384,N_5032,N_4017);
nor U6385 (N_6385,N_4914,N_4281);
or U6386 (N_6386,N_4611,N_5529);
nand U6387 (N_6387,N_4507,N_5434);
nand U6388 (N_6388,N_5325,N_4433);
or U6389 (N_6389,N_5915,N_4753);
and U6390 (N_6390,N_4908,N_4348);
nor U6391 (N_6391,N_4515,N_5518);
xor U6392 (N_6392,N_5476,N_4885);
xor U6393 (N_6393,N_5275,N_4829);
xor U6394 (N_6394,N_4538,N_4174);
and U6395 (N_6395,N_5662,N_5135);
nor U6396 (N_6396,N_4389,N_5157);
and U6397 (N_6397,N_4540,N_4772);
nand U6398 (N_6398,N_4012,N_5378);
xnor U6399 (N_6399,N_5655,N_4293);
nand U6400 (N_6400,N_5111,N_5631);
and U6401 (N_6401,N_5712,N_4447);
and U6402 (N_6402,N_5355,N_4709);
nand U6403 (N_6403,N_4702,N_4407);
or U6404 (N_6404,N_4827,N_4977);
and U6405 (N_6405,N_4109,N_5035);
nand U6406 (N_6406,N_4112,N_5565);
nand U6407 (N_6407,N_4637,N_5557);
and U6408 (N_6408,N_4177,N_4748);
nand U6409 (N_6409,N_4380,N_4625);
nor U6410 (N_6410,N_5650,N_5567);
nand U6411 (N_6411,N_5156,N_4756);
and U6412 (N_6412,N_4367,N_5022);
nor U6413 (N_6413,N_4459,N_4826);
xnor U6414 (N_6414,N_5588,N_4843);
nand U6415 (N_6415,N_4599,N_4235);
nand U6416 (N_6416,N_4251,N_4014);
or U6417 (N_6417,N_5946,N_4542);
nand U6418 (N_6418,N_4036,N_4475);
or U6419 (N_6419,N_5395,N_4055);
nand U6420 (N_6420,N_4966,N_5132);
xor U6421 (N_6421,N_5875,N_5987);
or U6422 (N_6422,N_4198,N_5980);
or U6423 (N_6423,N_4463,N_5545);
nand U6424 (N_6424,N_4393,N_5615);
and U6425 (N_6425,N_5049,N_4659);
xor U6426 (N_6426,N_4663,N_5179);
and U6427 (N_6427,N_4681,N_4076);
nand U6428 (N_6428,N_5724,N_4025);
or U6429 (N_6429,N_5955,N_5019);
and U6430 (N_6430,N_5549,N_4939);
nand U6431 (N_6431,N_5024,N_5865);
and U6432 (N_6432,N_4008,N_5728);
xor U6433 (N_6433,N_4840,N_4905);
and U6434 (N_6434,N_4087,N_5461);
nor U6435 (N_6435,N_4080,N_5971);
xor U6436 (N_6436,N_4970,N_4110);
nand U6437 (N_6437,N_4290,N_5920);
nand U6438 (N_6438,N_4526,N_5121);
or U6439 (N_6439,N_4581,N_4689);
and U6440 (N_6440,N_4197,N_5694);
nor U6441 (N_6441,N_5467,N_4839);
or U6442 (N_6442,N_4861,N_4602);
and U6443 (N_6443,N_4494,N_4578);
xnor U6444 (N_6444,N_4021,N_5138);
or U6445 (N_6445,N_5163,N_5377);
nor U6446 (N_6446,N_5198,N_4657);
nand U6447 (N_6447,N_4887,N_4467);
or U6448 (N_6448,N_5872,N_4037);
xor U6449 (N_6449,N_4336,N_5058);
and U6450 (N_6450,N_4525,N_5071);
or U6451 (N_6451,N_4097,N_4142);
xor U6452 (N_6452,N_4366,N_5068);
and U6453 (N_6453,N_4751,N_5191);
nand U6454 (N_6454,N_5919,N_5332);
nand U6455 (N_6455,N_5975,N_4351);
nor U6456 (N_6456,N_5576,N_4141);
nor U6457 (N_6457,N_5103,N_4056);
or U6458 (N_6458,N_4416,N_5470);
nor U6459 (N_6459,N_5151,N_4118);
or U6460 (N_6460,N_4340,N_5687);
and U6461 (N_6461,N_5302,N_5779);
and U6462 (N_6462,N_4227,N_4358);
or U6463 (N_6463,N_5067,N_4644);
nor U6464 (N_6464,N_4847,N_4718);
and U6465 (N_6465,N_4582,N_4363);
or U6466 (N_6466,N_5811,N_5699);
and U6467 (N_6467,N_5698,N_5977);
xnor U6468 (N_6468,N_5730,N_4639);
and U6469 (N_6469,N_4126,N_5387);
nand U6470 (N_6470,N_5598,N_5128);
xnor U6471 (N_6471,N_5048,N_5324);
xnor U6472 (N_6472,N_5446,N_4294);
nand U6473 (N_6473,N_4406,N_4980);
or U6474 (N_6474,N_4341,N_4365);
or U6475 (N_6475,N_4559,N_5439);
nor U6476 (N_6476,N_5407,N_5609);
nand U6477 (N_6477,N_4253,N_5766);
nor U6478 (N_6478,N_4477,N_4722);
and U6479 (N_6479,N_5523,N_4187);
or U6480 (N_6480,N_4216,N_5843);
nor U6481 (N_6481,N_4295,N_5131);
nor U6482 (N_6482,N_5076,N_5401);
nand U6483 (N_6483,N_5297,N_4673);
xnor U6484 (N_6484,N_5963,N_4752);
or U6485 (N_6485,N_5821,N_5220);
nor U6486 (N_6486,N_5577,N_5263);
nand U6487 (N_6487,N_5258,N_5622);
and U6488 (N_6488,N_5488,N_4326);
nor U6489 (N_6489,N_5554,N_4610);
xor U6490 (N_6490,N_5794,N_4298);
nor U6491 (N_6491,N_4512,N_5364);
or U6492 (N_6492,N_4131,N_4117);
nand U6493 (N_6493,N_5380,N_5926);
xnor U6494 (N_6494,N_5027,N_4920);
nor U6495 (N_6495,N_4376,N_4940);
or U6496 (N_6496,N_5512,N_5864);
and U6497 (N_6497,N_5442,N_5629);
nor U6498 (N_6498,N_5824,N_4058);
nor U6499 (N_6499,N_4305,N_4650);
nand U6500 (N_6500,N_4237,N_4609);
nand U6501 (N_6501,N_5411,N_4794);
xor U6502 (N_6502,N_5372,N_5369);
nor U6503 (N_6503,N_5271,N_5669);
xor U6504 (N_6504,N_4994,N_4617);
xnor U6505 (N_6505,N_4543,N_5123);
or U6506 (N_6506,N_4915,N_5828);
or U6507 (N_6507,N_5424,N_4670);
nand U6508 (N_6508,N_4574,N_4916);
or U6509 (N_6509,N_5880,N_4205);
or U6510 (N_6510,N_4828,N_4395);
nand U6511 (N_6511,N_5559,N_4173);
and U6512 (N_6512,N_5634,N_4569);
nor U6513 (N_6513,N_4095,N_4289);
xnor U6514 (N_6514,N_4361,N_5025);
nor U6515 (N_6515,N_4627,N_5595);
and U6516 (N_6516,N_5555,N_5616);
and U6517 (N_6517,N_5043,N_5063);
xnor U6518 (N_6518,N_5337,N_5638);
or U6519 (N_6519,N_5928,N_4634);
and U6520 (N_6520,N_4734,N_4876);
and U6521 (N_6521,N_5053,N_5688);
nand U6522 (N_6522,N_5335,N_5823);
or U6523 (N_6523,N_4864,N_5768);
nand U6524 (N_6524,N_5765,N_4600);
nor U6525 (N_6525,N_5753,N_4615);
nand U6526 (N_6526,N_5564,N_4498);
nand U6527 (N_6527,N_5328,N_5903);
nand U6528 (N_6528,N_5857,N_5607);
and U6529 (N_6529,N_4682,N_5141);
xor U6530 (N_6530,N_5961,N_4811);
nor U6531 (N_6531,N_4805,N_4041);
and U6532 (N_6532,N_4675,N_5368);
and U6533 (N_6533,N_4888,N_5016);
and U6534 (N_6534,N_4493,N_4373);
nand U6535 (N_6535,N_5110,N_5211);
or U6536 (N_6536,N_5580,N_5834);
nand U6537 (N_6537,N_4963,N_4664);
nand U6538 (N_6538,N_4094,N_5767);
and U6539 (N_6539,N_4287,N_4851);
nor U6540 (N_6540,N_4446,N_5247);
or U6541 (N_6541,N_5351,N_5408);
or U6542 (N_6542,N_5140,N_5939);
nand U6543 (N_6543,N_4897,N_5409);
or U6544 (N_6544,N_5323,N_5890);
and U6545 (N_6545,N_4700,N_5827);
or U6546 (N_6546,N_4084,N_4394);
or U6547 (N_6547,N_5729,N_5603);
nor U6548 (N_6548,N_4773,N_5596);
and U6549 (N_6549,N_5990,N_5264);
or U6550 (N_6550,N_5224,N_5120);
nor U6551 (N_6551,N_4377,N_5921);
or U6552 (N_6552,N_5873,N_4086);
nand U6553 (N_6553,N_5427,N_4047);
xnor U6554 (N_6554,N_5540,N_5000);
nor U6555 (N_6555,N_4746,N_4132);
nand U6556 (N_6556,N_5968,N_4921);
nand U6557 (N_6557,N_4158,N_5069);
or U6558 (N_6558,N_5701,N_4822);
or U6559 (N_6559,N_4057,N_5893);
or U6560 (N_6560,N_5613,N_4561);
xor U6561 (N_6561,N_4192,N_4984);
nor U6562 (N_6562,N_4654,N_5878);
nand U6563 (N_6563,N_5175,N_5671);
and U6564 (N_6564,N_4780,N_4269);
and U6565 (N_6565,N_4218,N_4798);
or U6566 (N_6566,N_4189,N_4750);
xnor U6567 (N_6567,N_5136,N_5562);
xor U6568 (N_6568,N_5740,N_4684);
xnor U6569 (N_6569,N_4278,N_5084);
and U6570 (N_6570,N_5245,N_5783);
or U6571 (N_6571,N_5130,N_4846);
nor U6572 (N_6572,N_4808,N_5336);
xnor U6573 (N_6573,N_4068,N_4713);
nand U6574 (N_6574,N_4640,N_4454);
nand U6575 (N_6575,N_5579,N_5182);
nand U6576 (N_6576,N_5142,N_5592);
nand U6577 (N_6577,N_4217,N_4795);
or U6578 (N_6578,N_4031,N_4449);
and U6579 (N_6579,N_5542,N_4757);
nand U6580 (N_6580,N_5194,N_4181);
or U6581 (N_6581,N_5404,N_5820);
or U6582 (N_6582,N_5430,N_5897);
nor U6583 (N_6583,N_5593,N_5287);
xor U6584 (N_6584,N_5168,N_5342);
nand U6585 (N_6585,N_4768,N_5994);
nand U6586 (N_6586,N_5343,N_4927);
and U6587 (N_6587,N_5651,N_5589);
or U6588 (N_6588,N_4255,N_4254);
and U6589 (N_6589,N_4196,N_5383);
or U6590 (N_6590,N_5850,N_4590);
nor U6591 (N_6591,N_4987,N_4952);
nor U6592 (N_6592,N_5117,N_4767);
nor U6593 (N_6593,N_4387,N_4437);
nor U6594 (N_6594,N_4033,N_5209);
or U6595 (N_6595,N_5719,N_4420);
and U6596 (N_6596,N_4116,N_5721);
nand U6597 (N_6597,N_4739,N_5758);
xor U6598 (N_6598,N_5643,N_5829);
and U6599 (N_6599,N_4414,N_4123);
or U6600 (N_6600,N_4736,N_4183);
or U6601 (N_6601,N_4825,N_4638);
or U6602 (N_6602,N_5608,N_5742);
and U6603 (N_6603,N_5327,N_5333);
or U6604 (N_6604,N_5023,N_5839);
or U6605 (N_6605,N_5214,N_4219);
and U6606 (N_6606,N_5386,N_4070);
or U6607 (N_6607,N_4852,N_5484);
and U6608 (N_6608,N_5731,N_5415);
nand U6609 (N_6609,N_4771,N_4575);
and U6610 (N_6610,N_5654,N_5624);
and U6611 (N_6611,N_4020,N_5226);
nor U6612 (N_6612,N_4457,N_4671);
nand U6613 (N_6613,N_5234,N_5011);
and U6614 (N_6614,N_5583,N_5199);
or U6615 (N_6615,N_4567,N_4115);
nor U6616 (N_6616,N_5706,N_4564);
or U6617 (N_6617,N_5490,N_4948);
and U6618 (N_6618,N_5594,N_5373);
and U6619 (N_6619,N_5936,N_5800);
or U6620 (N_6620,N_4066,N_5854);
nand U6621 (N_6621,N_4168,N_5457);
xor U6622 (N_6622,N_4522,N_4699);
and U6623 (N_6623,N_5749,N_4027);
or U6624 (N_6624,N_4496,N_5159);
nand U6625 (N_6625,N_4401,N_4339);
or U6626 (N_6626,N_4913,N_5983);
nand U6627 (N_6627,N_5243,N_4434);
nor U6628 (N_6628,N_4947,N_5524);
nor U6629 (N_6629,N_5492,N_4107);
nand U6630 (N_6630,N_4688,N_4424);
or U6631 (N_6631,N_5860,N_5330);
or U6632 (N_6632,N_4104,N_5535);
and U6633 (N_6633,N_4337,N_5544);
xnor U6634 (N_6634,N_4717,N_5089);
and U6635 (N_6635,N_5600,N_5789);
or U6636 (N_6636,N_4169,N_4303);
and U6637 (N_6637,N_4815,N_5953);
and U6638 (N_6638,N_5711,N_4587);
nand U6639 (N_6639,N_5249,N_5268);
nor U6640 (N_6640,N_5531,N_5133);
and U6641 (N_6641,N_4783,N_5808);
nor U6642 (N_6642,N_5246,N_4359);
nand U6643 (N_6643,N_4484,N_5705);
nand U6644 (N_6644,N_4749,N_5532);
nor U6645 (N_6645,N_4005,N_5218);
or U6646 (N_6646,N_5883,N_5341);
nor U6647 (N_6647,N_5397,N_4614);
or U6648 (N_6648,N_4098,N_4807);
xor U6649 (N_6649,N_5137,N_4203);
or U6650 (N_6650,N_4787,N_4384);
and U6651 (N_6651,N_4137,N_4981);
or U6652 (N_6652,N_5326,N_4155);
and U6653 (N_6653,N_5272,N_5190);
xor U6654 (N_6654,N_5160,N_5228);
nand U6655 (N_6655,N_5388,N_5080);
and U6656 (N_6656,N_5185,N_5648);
nand U6657 (N_6657,N_4593,N_5796);
nor U6658 (N_6658,N_5184,N_4955);
or U6659 (N_6659,N_4620,N_4108);
and U6660 (N_6660,N_4343,N_5528);
nand U6661 (N_6661,N_4992,N_4737);
or U6662 (N_6662,N_4486,N_4035);
and U6663 (N_6663,N_4557,N_4182);
xnor U6664 (N_6664,N_5474,N_4838);
or U6665 (N_6665,N_4221,N_5707);
nand U6666 (N_6666,N_5250,N_4988);
nand U6667 (N_6667,N_5309,N_4665);
nor U6668 (N_6668,N_5815,N_5885);
or U6669 (N_6669,N_4354,N_5948);
xnor U6670 (N_6670,N_4130,N_5172);
and U6671 (N_6671,N_5925,N_5619);
nor U6672 (N_6672,N_4803,N_4452);
and U6673 (N_6673,N_5906,N_4078);
or U6674 (N_6674,N_5803,N_5664);
or U6675 (N_6675,N_4819,N_5458);
or U6676 (N_6676,N_5644,N_4869);
or U6677 (N_6677,N_4606,N_5746);
nand U6678 (N_6678,N_4353,N_4594);
xor U6679 (N_6679,N_5456,N_4313);
or U6680 (N_6680,N_5586,N_4678);
or U6681 (N_6681,N_5007,N_4667);
nand U6682 (N_6682,N_5074,N_5210);
nand U6683 (N_6683,N_4306,N_4577);
nand U6684 (N_6684,N_4649,N_4448);
or U6685 (N_6685,N_5747,N_4415);
nor U6686 (N_6686,N_4266,N_5459);
and U6687 (N_6687,N_5187,N_4256);
nor U6688 (N_6688,N_4160,N_4212);
and U6689 (N_6689,N_4299,N_5255);
nor U6690 (N_6690,N_5034,N_5830);
or U6691 (N_6691,N_4546,N_4371);
or U6692 (N_6692,N_4723,N_4833);
or U6693 (N_6693,N_5914,N_5448);
or U6694 (N_6694,N_5582,N_4516);
or U6695 (N_6695,N_4268,N_4946);
nand U6696 (N_6696,N_4595,N_5663);
xor U6697 (N_6697,N_4029,N_5420);
and U6698 (N_6698,N_5036,N_4961);
nor U6699 (N_6699,N_4789,N_5266);
xnor U6700 (N_6700,N_5345,N_5633);
nand U6701 (N_6701,N_4466,N_4598);
and U6702 (N_6702,N_4148,N_4267);
and U6703 (N_6703,N_5344,N_5283);
xnor U6704 (N_6704,N_4793,N_4026);
and U6705 (N_6705,N_5847,N_5945);
and U6706 (N_6706,N_4879,N_4470);
nor U6707 (N_6707,N_4986,N_4740);
or U6708 (N_6708,N_5096,N_4802);
and U6709 (N_6709,N_4622,N_5674);
and U6710 (N_6710,N_5500,N_5932);
xnor U6711 (N_6711,N_5590,N_5483);
xor U6712 (N_6712,N_4143,N_5236);
xnor U6713 (N_6713,N_4121,N_5640);
or U6714 (N_6714,N_5539,N_5331);
nor U6715 (N_6715,N_4450,N_5261);
or U6716 (N_6716,N_4292,N_4841);
xor U6717 (N_6717,N_5293,N_5375);
or U6718 (N_6718,N_5173,N_5951);
xor U6719 (N_6719,N_5738,N_5814);
xor U6720 (N_6720,N_5673,N_4553);
nor U6721 (N_6721,N_5059,N_5846);
xor U6722 (N_6722,N_5166,N_4469);
xnor U6723 (N_6723,N_5060,N_5858);
and U6724 (N_6724,N_4636,N_4206);
or U6725 (N_6725,N_4460,N_5028);
xor U6726 (N_6726,N_4550,N_4028);
nor U6727 (N_6727,N_4770,N_5965);
and U6728 (N_6728,N_4968,N_5835);
and U6729 (N_6729,N_5741,N_4809);
xor U6730 (N_6730,N_5308,N_4332);
or U6731 (N_6731,N_5033,N_4660);
or U6732 (N_6732,N_4618,N_4411);
nand U6733 (N_6733,N_4714,N_4492);
or U6734 (N_6734,N_4195,N_4119);
or U6735 (N_6735,N_5610,N_4122);
nand U6736 (N_6736,N_4324,N_4845);
and U6737 (N_6737,N_4375,N_4153);
nand U6738 (N_6738,N_5256,N_5041);
or U6739 (N_6739,N_4220,N_4147);
or U6740 (N_6740,N_4234,N_4405);
nand U6741 (N_6741,N_5285,N_4658);
and U6742 (N_6742,N_5876,N_4676);
and U6743 (N_6743,N_5480,N_5305);
and U6744 (N_6744,N_4213,N_4848);
nor U6745 (N_6745,N_4733,N_5392);
or U6746 (N_6746,N_5892,N_4134);
and U6747 (N_6747,N_5852,N_4229);
nand U6748 (N_6748,N_5078,N_4038);
nor U6749 (N_6749,N_5737,N_5495);
and U6750 (N_6750,N_5802,N_4479);
and U6751 (N_6751,N_4549,N_5306);
and U6752 (N_6752,N_4368,N_4400);
nand U6753 (N_6753,N_4302,N_4226);
nor U6754 (N_6754,N_4954,N_5620);
nor U6755 (N_6755,N_4960,N_5723);
nand U6756 (N_6756,N_5329,N_5678);
xor U6757 (N_6757,N_5167,N_4385);
xor U6758 (N_6758,N_5836,N_4172);
and U6759 (N_6759,N_4962,N_5898);
and U6760 (N_6760,N_5986,N_4441);
or U6761 (N_6761,N_4779,N_4529);
and U6762 (N_6762,N_5253,N_5052);
or U6763 (N_6763,N_5806,N_4957);
and U6764 (N_6764,N_4455,N_4136);
xnor U6765 (N_6765,N_5050,N_4325);
nand U6766 (N_6766,N_5817,N_5026);
xnor U6767 (N_6767,N_5750,N_5900);
or U6768 (N_6768,N_5193,N_4672);
nor U6769 (N_6769,N_5489,N_5525);
nor U6770 (N_6770,N_4100,N_5281);
or U6771 (N_6771,N_5273,N_5795);
nand U6772 (N_6772,N_4390,N_4842);
nand U6773 (N_6773,N_5319,N_4431);
nand U6774 (N_6774,N_5511,N_5354);
xnor U6775 (N_6775,N_4693,N_4011);
nor U6776 (N_6776,N_4193,N_5421);
nand U6777 (N_6777,N_4797,N_4886);
nand U6778 (N_6778,N_5708,N_5418);
nor U6779 (N_6779,N_5248,N_4769);
or U6780 (N_6780,N_5107,N_4624);
nor U6781 (N_6781,N_5849,N_4440);
nor U6782 (N_6782,N_5637,N_5125);
or U6783 (N_6783,N_5513,N_5745);
and U6784 (N_6784,N_4856,N_4778);
nand U6785 (N_6785,N_5625,N_5161);
xnor U6786 (N_6786,N_5907,N_5761);
or U6787 (N_6787,N_4480,N_5668);
xor U6788 (N_6788,N_5656,N_5195);
or U6789 (N_6789,N_4880,N_4555);
xnor U6790 (N_6790,N_4884,N_5347);
xnor U6791 (N_6791,N_5310,N_4817);
xor U6792 (N_6792,N_4161,N_4178);
nand U6793 (N_6793,N_5510,N_4482);
or U6794 (N_6794,N_5763,N_4890);
xnor U6795 (N_6795,N_4458,N_4171);
nor U6796 (N_6796,N_4941,N_4866);
nor U6797 (N_6797,N_4429,N_5229);
or U6798 (N_6798,N_5714,N_4918);
xnor U6799 (N_6799,N_4993,N_5805);
xor U6800 (N_6800,N_4009,N_5419);
and U6801 (N_6801,N_5414,N_5203);
nand U6802 (N_6802,N_5317,N_4403);
nand U6803 (N_6803,N_5088,N_5188);
or U6804 (N_6804,N_4260,N_4568);
xnor U6805 (N_6805,N_4499,N_5884);
and U6806 (N_6806,N_4668,N_4002);
nand U6807 (N_6807,N_5295,N_4240);
nand U6808 (N_6808,N_4053,N_4272);
or U6809 (N_6809,N_5358,N_4814);
xor U6810 (N_6810,N_4379,N_5460);
xnor U6811 (N_6811,N_5365,N_4472);
nand U6812 (N_6812,N_5001,N_5659);
nor U6813 (N_6813,N_5578,N_4894);
and U6814 (N_6814,N_5822,N_4083);
xor U6815 (N_6815,N_5051,N_4999);
or U6816 (N_6816,N_5004,N_5646);
xnor U6817 (N_6817,N_5494,N_4674);
xnor U6818 (N_6818,N_4932,N_5497);
and U6819 (N_6819,N_5563,N_4372);
or U6820 (N_6820,N_4677,N_5046);
nand U6821 (N_6821,N_5547,N_5045);
nor U6822 (N_6822,N_4923,N_4669);
or U6823 (N_6823,N_4421,N_4309);
nor U6824 (N_6824,N_4088,N_4180);
nand U6825 (N_6825,N_4589,N_4064);
or U6826 (N_6826,N_5090,N_5396);
xnor U6827 (N_6827,N_4381,N_4139);
or U6828 (N_6828,N_5530,N_4539);
or U6829 (N_6829,N_4043,N_5520);
nand U6830 (N_6830,N_5606,N_4958);
and U6831 (N_6831,N_4464,N_5278);
nor U6832 (N_6832,N_4951,N_5350);
xor U6833 (N_6833,N_4225,N_5507);
or U6834 (N_6834,N_5770,N_4583);
or U6835 (N_6835,N_4270,N_5743);
xor U6836 (N_6836,N_5106,N_5683);
or U6837 (N_6837,N_5171,N_4000);
xnor U6838 (N_6838,N_5029,N_5754);
nor U6839 (N_6839,N_5289,N_4164);
or U6840 (N_6840,N_4548,N_5270);
nand U6841 (N_6841,N_5896,N_5551);
nor U6842 (N_6842,N_5639,N_4202);
xnor U6843 (N_6843,N_5982,N_4870);
or U6844 (N_6844,N_4643,N_4983);
xnor U6845 (N_6845,N_4998,N_5844);
and U6846 (N_6846,N_4629,N_5290);
and U6847 (N_6847,N_4474,N_4974);
or U6848 (N_6848,N_5757,N_5017);
nor U6849 (N_6849,N_4517,N_4207);
nand U6850 (N_6850,N_4152,N_5265);
and U6851 (N_6851,N_5200,N_5647);
nand U6852 (N_6852,N_4106,N_4144);
nand U6853 (N_6853,N_4964,N_5466);
and U6854 (N_6854,N_4497,N_4264);
xor U6855 (N_6855,N_4922,N_4872);
nand U6856 (N_6856,N_5441,N_4628);
and U6857 (N_6857,N_4342,N_4016);
or U6858 (N_6858,N_4199,N_5150);
or U6859 (N_6859,N_4500,N_5572);
nand U6860 (N_6860,N_5180,N_5361);
and U6861 (N_6861,N_5294,N_5979);
xor U6862 (N_6862,N_4796,N_4096);
xor U6863 (N_6863,N_4965,N_4655);
or U6864 (N_6864,N_5040,N_4426);
xor U6865 (N_6865,N_4246,N_4656);
nor U6866 (N_6866,N_5611,N_5206);
xnor U6867 (N_6867,N_4063,N_5118);
nand U6868 (N_6868,N_4327,N_5225);
and U6869 (N_6869,N_5104,N_5353);
nor U6870 (N_6870,N_5455,N_4184);
and U6871 (N_6871,N_5227,N_4732);
nand U6872 (N_6872,N_4917,N_5304);
nor U6873 (N_6873,N_5764,N_5935);
nand U6874 (N_6874,N_5081,N_5911);
nand U6875 (N_6875,N_4626,N_5018);
nor U6876 (N_6876,N_5604,N_5091);
xor U6877 (N_6877,N_5473,N_5425);
or U6878 (N_6878,N_5239,N_5623);
or U6879 (N_6879,N_5094,N_4695);
nor U6880 (N_6880,N_5472,N_4103);
and U6881 (N_6881,N_4236,N_4146);
xnor U6882 (N_6882,N_4661,N_4321);
nor U6883 (N_6883,N_4895,N_4708);
xnor U6884 (N_6884,N_4743,N_5079);
nor U6885 (N_6885,N_4019,N_4703);
or U6886 (N_6886,N_4900,N_5573);
nor U6887 (N_6887,N_5162,N_5895);
nor U6888 (N_6888,N_5682,N_4050);
xnor U6889 (N_6889,N_5697,N_4931);
and U6890 (N_6890,N_5280,N_4727);
nor U6891 (N_6891,N_4967,N_4478);
and U6892 (N_6892,N_5394,N_4701);
nor U6893 (N_6893,N_5845,N_5262);
nor U6894 (N_6894,N_4501,N_4810);
xnor U6895 (N_6895,N_4631,N_5527);
or U6896 (N_6896,N_4813,N_5389);
nand U6897 (N_6897,N_4903,N_4755);
nor U6898 (N_6898,N_5859,N_4114);
and U6899 (N_6899,N_5665,N_4836);
nor U6900 (N_6900,N_5444,N_4726);
nor U6901 (N_6901,N_5550,N_4859);
or U6902 (N_6902,N_4603,N_4976);
and U6903 (N_6903,N_5667,N_5113);
and U6904 (N_6904,N_4687,N_4820);
nor U6905 (N_6905,N_4135,N_5346);
and U6906 (N_6906,N_4356,N_4242);
or U6907 (N_6907,N_4874,N_4586);
nand U6908 (N_6908,N_5736,N_4572);
nand U6909 (N_6909,N_5116,N_5316);
or U6910 (N_6910,N_5197,N_4503);
xor U6911 (N_6911,N_4854,N_5832);
or U6912 (N_6912,N_4901,N_4291);
nand U6913 (N_6913,N_5966,N_4300);
or U6914 (N_6914,N_4719,N_4924);
and U6915 (N_6915,N_5124,N_5702);
nand U6916 (N_6916,N_5242,N_5985);
or U6917 (N_6917,N_5605,N_5057);
and U6918 (N_6918,N_5299,N_4170);
xor U6919 (N_6919,N_4902,N_5475);
or U6920 (N_6920,N_5153,N_4258);
nand U6921 (N_6921,N_4899,N_5696);
or U6922 (N_6922,N_4996,N_5584);
nor U6923 (N_6923,N_5254,N_4930);
nor U6924 (N_6924,N_5431,N_5291);
and U6925 (N_6925,N_5543,N_5367);
or U6926 (N_6926,N_4101,N_4487);
and U6927 (N_6927,N_5614,N_4692);
nand U6928 (N_6928,N_4978,N_5445);
and U6929 (N_6929,N_4436,N_4635);
and U6930 (N_6930,N_5215,N_5385);
or U6931 (N_6931,N_5956,N_4357);
nor U6932 (N_6932,N_4982,N_5989);
xnor U6933 (N_6933,N_4435,N_5496);
nor U6934 (N_6934,N_5887,N_5207);
nand U6935 (N_6935,N_4728,N_5617);
nor U6936 (N_6936,N_4276,N_4537);
nor U6937 (N_6937,N_4653,N_5952);
xnor U6938 (N_6938,N_5923,N_4524);
xor U6939 (N_6939,N_5485,N_4211);
nor U6940 (N_6940,N_5435,N_5801);
or U6941 (N_6941,N_5406,N_5481);
nand U6942 (N_6942,N_5818,N_5722);
and U6943 (N_6943,N_5447,N_5685);
or U6944 (N_6944,N_4697,N_4799);
nand U6945 (N_6945,N_5981,N_4156);
nor U6946 (N_6946,N_5790,N_4150);
and U6947 (N_6947,N_4782,N_4275);
nand U6948 (N_6948,N_5799,N_4355);
xor U6949 (N_6949,N_4704,N_4608);
nor U6950 (N_6950,N_5649,N_4835);
nor U6951 (N_6951,N_4046,N_4386);
xnor U6952 (N_6952,N_4244,N_4185);
xor U6953 (N_6953,N_5910,N_5379);
or U6954 (N_6954,N_5937,N_5143);
or U6955 (N_6955,N_5526,N_4398);
xnor U6956 (N_6956,N_5037,N_5097);
and U6957 (N_6957,N_5390,N_5645);
and U6958 (N_6958,N_5075,N_5056);
nor U6959 (N_6959,N_4995,N_5626);
and U6960 (N_6960,N_4151,N_5469);
nor U6961 (N_6961,N_5621,N_5999);
nand U6962 (N_6962,N_4124,N_5464);
nand U6963 (N_6963,N_4533,N_5292);
or U6964 (N_6964,N_5098,N_4391);
and U6965 (N_6965,N_4956,N_5363);
xnor U6966 (N_6966,N_4308,N_4616);
xnor U6967 (N_6967,N_5978,N_5468);
or U6968 (N_6968,N_4277,N_4334);
nand U6969 (N_6969,N_4453,N_4775);
xnor U6970 (N_6970,N_5370,N_5739);
nand U6971 (N_6971,N_5813,N_4374);
xnor U6972 (N_6972,N_4402,N_5269);
nand U6973 (N_6973,N_5533,N_5340);
nor U6974 (N_6974,N_5732,N_4222);
xor U6975 (N_6975,N_5809,N_4069);
xnor U6976 (N_6976,N_4145,N_4877);
xor U6977 (N_6977,N_5286,N_5976);
xor U6978 (N_6978,N_4179,N_4690);
and U6979 (N_6979,N_4345,N_4712);
or U6980 (N_6980,N_5322,N_4745);
nand U6981 (N_6981,N_5432,N_5931);
and U6982 (N_6982,N_5095,N_5922);
and U6983 (N_6983,N_4249,N_5055);
xor U6984 (N_6984,N_4333,N_5680);
or U6985 (N_6985,N_4409,N_5498);
or U6986 (N_6986,N_5916,N_4777);
and U6987 (N_6987,N_4651,N_5984);
or U6988 (N_6988,N_5992,N_4099);
nor U6989 (N_6989,N_4350,N_5692);
or U6990 (N_6990,N_5752,N_5100);
or U6991 (N_6991,N_5232,N_5244);
nand U6992 (N_6992,N_4972,N_5521);
nor U6993 (N_6993,N_4800,N_4791);
and U6994 (N_6994,N_4560,N_4725);
and U6995 (N_6995,N_4370,N_5438);
or U6996 (N_6996,N_5877,N_5311);
or U6997 (N_6997,N_5710,N_5315);
or U6998 (N_6998,N_4715,N_4018);
and U6999 (N_6999,N_5504,N_4534);
or U7000 (N_7000,N_4853,N_4993);
nand U7001 (N_7001,N_4523,N_4394);
and U7002 (N_7002,N_5137,N_5922);
and U7003 (N_7003,N_4730,N_5816);
nor U7004 (N_7004,N_5723,N_5059);
nor U7005 (N_7005,N_4023,N_4422);
nand U7006 (N_7006,N_4564,N_4295);
xor U7007 (N_7007,N_5786,N_5869);
nand U7008 (N_7008,N_5082,N_5753);
and U7009 (N_7009,N_4303,N_4995);
nand U7010 (N_7010,N_5475,N_4904);
and U7011 (N_7011,N_5858,N_4031);
and U7012 (N_7012,N_4230,N_4454);
xor U7013 (N_7013,N_5961,N_4185);
xnor U7014 (N_7014,N_4323,N_5924);
nor U7015 (N_7015,N_5324,N_4695);
nand U7016 (N_7016,N_5151,N_5008);
or U7017 (N_7017,N_4474,N_4125);
and U7018 (N_7018,N_5368,N_5893);
nand U7019 (N_7019,N_5477,N_4265);
and U7020 (N_7020,N_4551,N_5441);
nor U7021 (N_7021,N_4916,N_5665);
nand U7022 (N_7022,N_5771,N_4817);
or U7023 (N_7023,N_5614,N_4169);
or U7024 (N_7024,N_4225,N_5653);
or U7025 (N_7025,N_4091,N_4564);
xor U7026 (N_7026,N_4043,N_5447);
xnor U7027 (N_7027,N_4547,N_5825);
nor U7028 (N_7028,N_5740,N_5001);
or U7029 (N_7029,N_4997,N_5928);
and U7030 (N_7030,N_5452,N_5308);
nor U7031 (N_7031,N_4383,N_4644);
xnor U7032 (N_7032,N_4350,N_5654);
and U7033 (N_7033,N_5704,N_5745);
nor U7034 (N_7034,N_5060,N_5083);
or U7035 (N_7035,N_4797,N_4370);
xnor U7036 (N_7036,N_5823,N_5051);
and U7037 (N_7037,N_5883,N_5983);
nor U7038 (N_7038,N_5000,N_5769);
or U7039 (N_7039,N_5824,N_4288);
xor U7040 (N_7040,N_5819,N_4582);
and U7041 (N_7041,N_5834,N_5887);
nand U7042 (N_7042,N_4069,N_5296);
xnor U7043 (N_7043,N_4097,N_4726);
nand U7044 (N_7044,N_4010,N_5549);
xor U7045 (N_7045,N_4898,N_4007);
and U7046 (N_7046,N_4107,N_4991);
nand U7047 (N_7047,N_5417,N_4498);
xnor U7048 (N_7048,N_5738,N_5499);
xor U7049 (N_7049,N_5767,N_4754);
nor U7050 (N_7050,N_4960,N_4566);
and U7051 (N_7051,N_5000,N_4947);
nor U7052 (N_7052,N_5002,N_4084);
and U7053 (N_7053,N_4156,N_4367);
nand U7054 (N_7054,N_5216,N_4078);
nor U7055 (N_7055,N_4406,N_4162);
nand U7056 (N_7056,N_4669,N_4447);
and U7057 (N_7057,N_4438,N_4958);
nor U7058 (N_7058,N_4198,N_5881);
or U7059 (N_7059,N_4456,N_5453);
xnor U7060 (N_7060,N_5609,N_4880);
and U7061 (N_7061,N_4198,N_4835);
xnor U7062 (N_7062,N_4538,N_4346);
nor U7063 (N_7063,N_5024,N_4393);
xnor U7064 (N_7064,N_5789,N_5412);
nor U7065 (N_7065,N_4317,N_5281);
or U7066 (N_7066,N_4003,N_5747);
nor U7067 (N_7067,N_4143,N_4808);
xnor U7068 (N_7068,N_5366,N_5154);
or U7069 (N_7069,N_4096,N_5010);
nor U7070 (N_7070,N_4122,N_4311);
xor U7071 (N_7071,N_4045,N_4472);
and U7072 (N_7072,N_5036,N_4726);
xnor U7073 (N_7073,N_4958,N_5733);
nand U7074 (N_7074,N_5177,N_4567);
and U7075 (N_7075,N_4958,N_4072);
nor U7076 (N_7076,N_4433,N_4888);
and U7077 (N_7077,N_4199,N_4697);
nor U7078 (N_7078,N_4109,N_5944);
nand U7079 (N_7079,N_5070,N_5703);
xor U7080 (N_7080,N_4817,N_5677);
nor U7081 (N_7081,N_4615,N_5830);
nand U7082 (N_7082,N_5574,N_4591);
nor U7083 (N_7083,N_4993,N_5626);
nor U7084 (N_7084,N_5770,N_4023);
nand U7085 (N_7085,N_4704,N_5673);
or U7086 (N_7086,N_5045,N_5986);
nand U7087 (N_7087,N_4323,N_4215);
and U7088 (N_7088,N_5051,N_5114);
nand U7089 (N_7089,N_5064,N_4976);
and U7090 (N_7090,N_4881,N_5253);
xnor U7091 (N_7091,N_4981,N_4962);
nor U7092 (N_7092,N_5832,N_4320);
xnor U7093 (N_7093,N_4758,N_4340);
xnor U7094 (N_7094,N_4028,N_5678);
nor U7095 (N_7095,N_4702,N_5404);
nor U7096 (N_7096,N_4339,N_5459);
nor U7097 (N_7097,N_4850,N_5387);
nand U7098 (N_7098,N_4703,N_5413);
nand U7099 (N_7099,N_4263,N_4059);
xnor U7100 (N_7100,N_4406,N_5729);
and U7101 (N_7101,N_4316,N_5555);
nor U7102 (N_7102,N_5739,N_5327);
nor U7103 (N_7103,N_4480,N_5468);
and U7104 (N_7104,N_4017,N_5583);
and U7105 (N_7105,N_5959,N_4357);
nand U7106 (N_7106,N_5121,N_4969);
nand U7107 (N_7107,N_4679,N_4434);
or U7108 (N_7108,N_4498,N_5842);
xor U7109 (N_7109,N_5625,N_4761);
xnor U7110 (N_7110,N_5909,N_5659);
nor U7111 (N_7111,N_5565,N_4364);
xor U7112 (N_7112,N_4722,N_4437);
nand U7113 (N_7113,N_4782,N_4920);
or U7114 (N_7114,N_4522,N_5605);
and U7115 (N_7115,N_5610,N_5858);
and U7116 (N_7116,N_4416,N_5108);
xor U7117 (N_7117,N_5916,N_5833);
nor U7118 (N_7118,N_5940,N_4071);
nand U7119 (N_7119,N_5281,N_5638);
nor U7120 (N_7120,N_4637,N_5637);
nor U7121 (N_7121,N_4195,N_5784);
nand U7122 (N_7122,N_4353,N_4537);
nor U7123 (N_7123,N_5636,N_5977);
xnor U7124 (N_7124,N_5026,N_4331);
and U7125 (N_7125,N_4926,N_5765);
and U7126 (N_7126,N_5177,N_4250);
nor U7127 (N_7127,N_5928,N_4088);
nand U7128 (N_7128,N_4453,N_4221);
or U7129 (N_7129,N_5899,N_5173);
and U7130 (N_7130,N_4331,N_4676);
nor U7131 (N_7131,N_4523,N_4707);
and U7132 (N_7132,N_5387,N_5275);
xnor U7133 (N_7133,N_5638,N_5530);
nand U7134 (N_7134,N_5566,N_5458);
and U7135 (N_7135,N_5167,N_5004);
xor U7136 (N_7136,N_4959,N_5774);
nor U7137 (N_7137,N_4322,N_5419);
or U7138 (N_7138,N_4468,N_5647);
nand U7139 (N_7139,N_4962,N_4441);
nand U7140 (N_7140,N_5000,N_4330);
nor U7141 (N_7141,N_5128,N_5845);
nor U7142 (N_7142,N_4329,N_5733);
nor U7143 (N_7143,N_5839,N_5345);
or U7144 (N_7144,N_5679,N_5995);
nor U7145 (N_7145,N_5935,N_5648);
nand U7146 (N_7146,N_5095,N_5384);
xor U7147 (N_7147,N_5146,N_4737);
nor U7148 (N_7148,N_4593,N_5846);
nand U7149 (N_7149,N_4729,N_5440);
nand U7150 (N_7150,N_4787,N_4843);
nor U7151 (N_7151,N_5206,N_5141);
nor U7152 (N_7152,N_5922,N_5793);
xnor U7153 (N_7153,N_4013,N_4446);
nor U7154 (N_7154,N_4453,N_4096);
or U7155 (N_7155,N_5058,N_4559);
xor U7156 (N_7156,N_4822,N_5080);
nor U7157 (N_7157,N_4253,N_5169);
nand U7158 (N_7158,N_4154,N_5825);
xor U7159 (N_7159,N_5682,N_5584);
xor U7160 (N_7160,N_5319,N_4733);
nand U7161 (N_7161,N_4485,N_5536);
nand U7162 (N_7162,N_4633,N_5131);
or U7163 (N_7163,N_5520,N_4323);
or U7164 (N_7164,N_5905,N_5980);
xor U7165 (N_7165,N_5905,N_4863);
nor U7166 (N_7166,N_5073,N_5776);
or U7167 (N_7167,N_4291,N_5175);
and U7168 (N_7168,N_5947,N_5166);
nor U7169 (N_7169,N_5021,N_4920);
nand U7170 (N_7170,N_4958,N_4754);
and U7171 (N_7171,N_5788,N_4094);
nor U7172 (N_7172,N_4108,N_5037);
or U7173 (N_7173,N_4666,N_4296);
nand U7174 (N_7174,N_4393,N_5278);
nor U7175 (N_7175,N_5182,N_4077);
nand U7176 (N_7176,N_4810,N_4920);
nor U7177 (N_7177,N_4735,N_4181);
nand U7178 (N_7178,N_5097,N_4041);
nor U7179 (N_7179,N_4107,N_5124);
and U7180 (N_7180,N_4518,N_5488);
nor U7181 (N_7181,N_4258,N_4085);
nor U7182 (N_7182,N_5307,N_4491);
or U7183 (N_7183,N_5522,N_5982);
nand U7184 (N_7184,N_5842,N_4300);
xnor U7185 (N_7185,N_4880,N_5750);
nor U7186 (N_7186,N_5213,N_4607);
and U7187 (N_7187,N_5625,N_5961);
nand U7188 (N_7188,N_4141,N_5148);
xor U7189 (N_7189,N_5785,N_4338);
or U7190 (N_7190,N_4165,N_4833);
xnor U7191 (N_7191,N_4628,N_4311);
xor U7192 (N_7192,N_5012,N_4778);
nand U7193 (N_7193,N_4824,N_5407);
nor U7194 (N_7194,N_5231,N_5523);
nand U7195 (N_7195,N_5073,N_4843);
or U7196 (N_7196,N_4036,N_4035);
nand U7197 (N_7197,N_4261,N_5849);
or U7198 (N_7198,N_4874,N_4944);
nor U7199 (N_7199,N_5661,N_5416);
nor U7200 (N_7200,N_4373,N_5153);
nor U7201 (N_7201,N_5574,N_5112);
xor U7202 (N_7202,N_4438,N_5616);
or U7203 (N_7203,N_4604,N_4907);
nand U7204 (N_7204,N_5795,N_5443);
nand U7205 (N_7205,N_5008,N_4711);
nor U7206 (N_7206,N_4368,N_5307);
xor U7207 (N_7207,N_5051,N_5230);
nor U7208 (N_7208,N_4694,N_5258);
xor U7209 (N_7209,N_5263,N_4057);
nand U7210 (N_7210,N_5589,N_5979);
xnor U7211 (N_7211,N_5402,N_4407);
and U7212 (N_7212,N_4682,N_4803);
and U7213 (N_7213,N_4690,N_4756);
and U7214 (N_7214,N_4986,N_4208);
xnor U7215 (N_7215,N_5135,N_5968);
nor U7216 (N_7216,N_5157,N_5533);
and U7217 (N_7217,N_5909,N_4844);
nand U7218 (N_7218,N_5400,N_4028);
and U7219 (N_7219,N_4479,N_5564);
nand U7220 (N_7220,N_4206,N_5203);
and U7221 (N_7221,N_5303,N_4403);
and U7222 (N_7222,N_5956,N_4735);
and U7223 (N_7223,N_4432,N_5926);
nor U7224 (N_7224,N_5393,N_4014);
nand U7225 (N_7225,N_5299,N_5907);
xor U7226 (N_7226,N_4607,N_5771);
xnor U7227 (N_7227,N_5218,N_5002);
or U7228 (N_7228,N_4576,N_5382);
nor U7229 (N_7229,N_4889,N_4710);
nor U7230 (N_7230,N_5639,N_5106);
nor U7231 (N_7231,N_5462,N_5922);
or U7232 (N_7232,N_5093,N_4066);
nor U7233 (N_7233,N_4773,N_4774);
nor U7234 (N_7234,N_4542,N_5280);
and U7235 (N_7235,N_4035,N_4224);
xnor U7236 (N_7236,N_4646,N_4993);
nor U7237 (N_7237,N_4318,N_5677);
nand U7238 (N_7238,N_4541,N_4674);
xnor U7239 (N_7239,N_5311,N_4939);
or U7240 (N_7240,N_4178,N_4763);
nor U7241 (N_7241,N_4501,N_4285);
nand U7242 (N_7242,N_4063,N_4561);
and U7243 (N_7243,N_4332,N_5087);
and U7244 (N_7244,N_5531,N_4501);
nand U7245 (N_7245,N_4994,N_4870);
or U7246 (N_7246,N_5642,N_4219);
and U7247 (N_7247,N_4758,N_4954);
nor U7248 (N_7248,N_4897,N_4269);
or U7249 (N_7249,N_4936,N_4944);
nor U7250 (N_7250,N_4395,N_4713);
nand U7251 (N_7251,N_4452,N_4287);
nand U7252 (N_7252,N_5620,N_4817);
nor U7253 (N_7253,N_4246,N_5923);
xnor U7254 (N_7254,N_4923,N_4399);
and U7255 (N_7255,N_5093,N_4116);
and U7256 (N_7256,N_5428,N_4022);
and U7257 (N_7257,N_5949,N_5759);
nor U7258 (N_7258,N_5768,N_4507);
or U7259 (N_7259,N_4999,N_5850);
xor U7260 (N_7260,N_4492,N_5867);
or U7261 (N_7261,N_4284,N_4216);
nor U7262 (N_7262,N_4750,N_4824);
nand U7263 (N_7263,N_5083,N_4509);
and U7264 (N_7264,N_4991,N_5612);
and U7265 (N_7265,N_5442,N_5435);
or U7266 (N_7266,N_5754,N_4599);
nand U7267 (N_7267,N_4038,N_4433);
and U7268 (N_7268,N_5885,N_5941);
xnor U7269 (N_7269,N_4273,N_4227);
nand U7270 (N_7270,N_5576,N_4479);
or U7271 (N_7271,N_4337,N_4468);
or U7272 (N_7272,N_5520,N_4131);
and U7273 (N_7273,N_5057,N_4804);
or U7274 (N_7274,N_5889,N_5119);
nor U7275 (N_7275,N_4306,N_5709);
or U7276 (N_7276,N_5322,N_4189);
and U7277 (N_7277,N_5423,N_5761);
xor U7278 (N_7278,N_4740,N_4621);
xnor U7279 (N_7279,N_4254,N_4645);
and U7280 (N_7280,N_5101,N_4825);
and U7281 (N_7281,N_5756,N_5401);
or U7282 (N_7282,N_4199,N_4816);
nand U7283 (N_7283,N_5159,N_4561);
nand U7284 (N_7284,N_5267,N_5646);
xor U7285 (N_7285,N_5425,N_4161);
nor U7286 (N_7286,N_4922,N_5582);
and U7287 (N_7287,N_5776,N_4435);
or U7288 (N_7288,N_5834,N_4602);
and U7289 (N_7289,N_4717,N_5618);
or U7290 (N_7290,N_4371,N_5482);
xor U7291 (N_7291,N_4381,N_5960);
or U7292 (N_7292,N_5790,N_4153);
xnor U7293 (N_7293,N_5636,N_4978);
nor U7294 (N_7294,N_5399,N_5380);
or U7295 (N_7295,N_4284,N_4815);
nor U7296 (N_7296,N_4181,N_5710);
nor U7297 (N_7297,N_5276,N_4150);
xor U7298 (N_7298,N_4698,N_5995);
nor U7299 (N_7299,N_5475,N_4799);
nor U7300 (N_7300,N_5063,N_4226);
nor U7301 (N_7301,N_5670,N_5594);
and U7302 (N_7302,N_5160,N_5814);
nand U7303 (N_7303,N_4766,N_4319);
and U7304 (N_7304,N_4694,N_5536);
or U7305 (N_7305,N_4649,N_5206);
and U7306 (N_7306,N_5673,N_4712);
and U7307 (N_7307,N_5956,N_4698);
and U7308 (N_7308,N_4543,N_5257);
nand U7309 (N_7309,N_5335,N_4105);
and U7310 (N_7310,N_4219,N_4677);
nand U7311 (N_7311,N_5237,N_5979);
nor U7312 (N_7312,N_4657,N_5798);
xor U7313 (N_7313,N_5030,N_4978);
and U7314 (N_7314,N_4518,N_5850);
nand U7315 (N_7315,N_5979,N_4808);
nand U7316 (N_7316,N_4897,N_4873);
nor U7317 (N_7317,N_4768,N_5109);
nor U7318 (N_7318,N_4357,N_5596);
or U7319 (N_7319,N_5115,N_4468);
nand U7320 (N_7320,N_4211,N_5490);
xor U7321 (N_7321,N_4960,N_4119);
nand U7322 (N_7322,N_5356,N_5814);
or U7323 (N_7323,N_4768,N_4070);
or U7324 (N_7324,N_5352,N_4528);
xor U7325 (N_7325,N_5538,N_4063);
nor U7326 (N_7326,N_4027,N_4666);
or U7327 (N_7327,N_4260,N_5264);
nor U7328 (N_7328,N_4835,N_4901);
or U7329 (N_7329,N_4017,N_5000);
xnor U7330 (N_7330,N_5508,N_5381);
nor U7331 (N_7331,N_5769,N_5327);
xor U7332 (N_7332,N_5499,N_5388);
or U7333 (N_7333,N_5909,N_5647);
nor U7334 (N_7334,N_5839,N_4939);
xnor U7335 (N_7335,N_5994,N_5407);
nand U7336 (N_7336,N_5940,N_5765);
xnor U7337 (N_7337,N_4698,N_4602);
xnor U7338 (N_7338,N_4651,N_4768);
nor U7339 (N_7339,N_5686,N_4625);
xor U7340 (N_7340,N_5209,N_5083);
or U7341 (N_7341,N_4475,N_4487);
nand U7342 (N_7342,N_5483,N_5876);
and U7343 (N_7343,N_5416,N_4990);
nand U7344 (N_7344,N_5646,N_5420);
nand U7345 (N_7345,N_4695,N_5386);
xnor U7346 (N_7346,N_5301,N_5691);
or U7347 (N_7347,N_5613,N_4667);
nor U7348 (N_7348,N_4635,N_5141);
nor U7349 (N_7349,N_4966,N_4660);
nand U7350 (N_7350,N_4763,N_5926);
or U7351 (N_7351,N_4086,N_5585);
nand U7352 (N_7352,N_5440,N_5129);
or U7353 (N_7353,N_5741,N_5277);
and U7354 (N_7354,N_5245,N_4975);
nor U7355 (N_7355,N_5734,N_4944);
nand U7356 (N_7356,N_4426,N_5668);
xor U7357 (N_7357,N_5111,N_4849);
nor U7358 (N_7358,N_5691,N_5907);
nor U7359 (N_7359,N_4989,N_5051);
and U7360 (N_7360,N_5726,N_5552);
nor U7361 (N_7361,N_4754,N_4250);
or U7362 (N_7362,N_5971,N_4584);
nor U7363 (N_7363,N_5765,N_5646);
and U7364 (N_7364,N_5972,N_5054);
xnor U7365 (N_7365,N_4918,N_5109);
nand U7366 (N_7366,N_5834,N_5793);
xnor U7367 (N_7367,N_5109,N_5456);
and U7368 (N_7368,N_5487,N_5865);
nor U7369 (N_7369,N_4737,N_4865);
nand U7370 (N_7370,N_5280,N_4614);
nor U7371 (N_7371,N_5992,N_4564);
nand U7372 (N_7372,N_5942,N_5800);
or U7373 (N_7373,N_5335,N_5876);
nor U7374 (N_7374,N_4502,N_4382);
xor U7375 (N_7375,N_5095,N_5566);
nand U7376 (N_7376,N_4007,N_4942);
nand U7377 (N_7377,N_4763,N_5273);
xor U7378 (N_7378,N_5365,N_5596);
xor U7379 (N_7379,N_5785,N_5582);
or U7380 (N_7380,N_5708,N_5738);
xor U7381 (N_7381,N_4031,N_4330);
xnor U7382 (N_7382,N_5560,N_4624);
nand U7383 (N_7383,N_5186,N_5503);
nor U7384 (N_7384,N_5766,N_4571);
xnor U7385 (N_7385,N_5855,N_5829);
or U7386 (N_7386,N_5686,N_4260);
xnor U7387 (N_7387,N_4455,N_4913);
xor U7388 (N_7388,N_4158,N_4454);
nor U7389 (N_7389,N_5346,N_4522);
or U7390 (N_7390,N_5948,N_4620);
nor U7391 (N_7391,N_5381,N_4993);
or U7392 (N_7392,N_4957,N_5783);
nand U7393 (N_7393,N_5293,N_4949);
xnor U7394 (N_7394,N_5020,N_4972);
nand U7395 (N_7395,N_4917,N_5568);
or U7396 (N_7396,N_5211,N_4217);
and U7397 (N_7397,N_4351,N_4991);
or U7398 (N_7398,N_4615,N_5100);
and U7399 (N_7399,N_4247,N_4595);
and U7400 (N_7400,N_4659,N_5533);
and U7401 (N_7401,N_5392,N_5302);
and U7402 (N_7402,N_5301,N_5289);
nand U7403 (N_7403,N_5119,N_5280);
nand U7404 (N_7404,N_4249,N_5815);
nor U7405 (N_7405,N_5560,N_4053);
and U7406 (N_7406,N_4769,N_5298);
and U7407 (N_7407,N_5713,N_4537);
or U7408 (N_7408,N_5646,N_4613);
or U7409 (N_7409,N_5784,N_5067);
xnor U7410 (N_7410,N_4627,N_4798);
or U7411 (N_7411,N_4476,N_4874);
or U7412 (N_7412,N_4010,N_4864);
and U7413 (N_7413,N_5488,N_4817);
xnor U7414 (N_7414,N_5546,N_4152);
nor U7415 (N_7415,N_4965,N_5879);
or U7416 (N_7416,N_4915,N_5420);
xor U7417 (N_7417,N_4151,N_4730);
xor U7418 (N_7418,N_5988,N_5033);
nand U7419 (N_7419,N_5866,N_4355);
or U7420 (N_7420,N_5050,N_4135);
nand U7421 (N_7421,N_4536,N_5850);
xor U7422 (N_7422,N_4508,N_4012);
xor U7423 (N_7423,N_5911,N_5974);
and U7424 (N_7424,N_5111,N_4356);
nand U7425 (N_7425,N_4372,N_4424);
or U7426 (N_7426,N_4744,N_5742);
or U7427 (N_7427,N_4602,N_5044);
or U7428 (N_7428,N_4273,N_5673);
or U7429 (N_7429,N_4402,N_4379);
or U7430 (N_7430,N_5240,N_5751);
xnor U7431 (N_7431,N_4459,N_4982);
xnor U7432 (N_7432,N_4139,N_4918);
or U7433 (N_7433,N_4309,N_4785);
or U7434 (N_7434,N_4493,N_4960);
nor U7435 (N_7435,N_4979,N_4679);
nor U7436 (N_7436,N_5972,N_5577);
and U7437 (N_7437,N_5721,N_4612);
nor U7438 (N_7438,N_4474,N_5762);
xnor U7439 (N_7439,N_4969,N_4994);
xnor U7440 (N_7440,N_4543,N_4388);
or U7441 (N_7441,N_5708,N_4388);
nand U7442 (N_7442,N_4788,N_4008);
nor U7443 (N_7443,N_5134,N_4523);
nor U7444 (N_7444,N_4582,N_5510);
xnor U7445 (N_7445,N_5345,N_4563);
and U7446 (N_7446,N_5497,N_5118);
or U7447 (N_7447,N_5886,N_4732);
or U7448 (N_7448,N_4884,N_5876);
nand U7449 (N_7449,N_4005,N_5136);
or U7450 (N_7450,N_4681,N_5502);
nor U7451 (N_7451,N_5594,N_5228);
and U7452 (N_7452,N_5737,N_5060);
and U7453 (N_7453,N_4576,N_5958);
nor U7454 (N_7454,N_4863,N_5157);
nand U7455 (N_7455,N_5809,N_4094);
or U7456 (N_7456,N_5601,N_5394);
and U7457 (N_7457,N_4055,N_5442);
and U7458 (N_7458,N_5238,N_5471);
nand U7459 (N_7459,N_5988,N_5690);
nor U7460 (N_7460,N_4559,N_4105);
nor U7461 (N_7461,N_5205,N_5901);
nand U7462 (N_7462,N_4634,N_4403);
xnor U7463 (N_7463,N_5842,N_5275);
nand U7464 (N_7464,N_4668,N_4306);
nor U7465 (N_7465,N_4767,N_4690);
and U7466 (N_7466,N_4926,N_5368);
and U7467 (N_7467,N_5716,N_5080);
nand U7468 (N_7468,N_5716,N_5444);
and U7469 (N_7469,N_4096,N_5593);
and U7470 (N_7470,N_5492,N_4221);
nand U7471 (N_7471,N_4638,N_5255);
nor U7472 (N_7472,N_5544,N_4467);
nor U7473 (N_7473,N_4908,N_4080);
nand U7474 (N_7474,N_5120,N_4015);
nor U7475 (N_7475,N_5508,N_4652);
or U7476 (N_7476,N_4614,N_5903);
nor U7477 (N_7477,N_4644,N_4295);
nor U7478 (N_7478,N_5743,N_4829);
nand U7479 (N_7479,N_5890,N_4812);
nand U7480 (N_7480,N_5673,N_5770);
xnor U7481 (N_7481,N_4846,N_4824);
or U7482 (N_7482,N_5359,N_5851);
and U7483 (N_7483,N_4922,N_4584);
or U7484 (N_7484,N_4419,N_4136);
nand U7485 (N_7485,N_5830,N_4540);
and U7486 (N_7486,N_5186,N_4101);
and U7487 (N_7487,N_4279,N_4594);
or U7488 (N_7488,N_5301,N_4026);
nand U7489 (N_7489,N_5548,N_5175);
xnor U7490 (N_7490,N_4536,N_5111);
and U7491 (N_7491,N_4771,N_4276);
or U7492 (N_7492,N_5544,N_4060);
or U7493 (N_7493,N_4547,N_5424);
nand U7494 (N_7494,N_4573,N_5623);
xor U7495 (N_7495,N_4923,N_5773);
or U7496 (N_7496,N_4298,N_5955);
xor U7497 (N_7497,N_4857,N_5938);
xnor U7498 (N_7498,N_5864,N_4427);
xnor U7499 (N_7499,N_4203,N_4123);
nand U7500 (N_7500,N_5959,N_5199);
xnor U7501 (N_7501,N_4555,N_5020);
xnor U7502 (N_7502,N_4285,N_5322);
xor U7503 (N_7503,N_5646,N_4562);
xor U7504 (N_7504,N_5658,N_4101);
and U7505 (N_7505,N_5797,N_5221);
xnor U7506 (N_7506,N_4945,N_4682);
and U7507 (N_7507,N_5112,N_5375);
xnor U7508 (N_7508,N_5282,N_5970);
nand U7509 (N_7509,N_4601,N_5186);
nand U7510 (N_7510,N_4827,N_4767);
or U7511 (N_7511,N_4974,N_4610);
xnor U7512 (N_7512,N_4818,N_4128);
nor U7513 (N_7513,N_5666,N_4433);
or U7514 (N_7514,N_4461,N_4578);
or U7515 (N_7515,N_5802,N_4010);
nor U7516 (N_7516,N_4378,N_4755);
nor U7517 (N_7517,N_5527,N_4787);
and U7518 (N_7518,N_4540,N_5189);
nand U7519 (N_7519,N_5375,N_4618);
or U7520 (N_7520,N_5630,N_5020);
and U7521 (N_7521,N_4072,N_4226);
xnor U7522 (N_7522,N_5901,N_5926);
nand U7523 (N_7523,N_5067,N_4737);
nor U7524 (N_7524,N_4537,N_4307);
nand U7525 (N_7525,N_5458,N_4533);
nor U7526 (N_7526,N_5894,N_5254);
nand U7527 (N_7527,N_5960,N_5904);
xor U7528 (N_7528,N_5397,N_4409);
or U7529 (N_7529,N_5757,N_4068);
and U7530 (N_7530,N_5774,N_4945);
nor U7531 (N_7531,N_5785,N_4016);
xor U7532 (N_7532,N_5340,N_5515);
or U7533 (N_7533,N_4965,N_4781);
xnor U7534 (N_7534,N_5032,N_4560);
or U7535 (N_7535,N_5721,N_5263);
and U7536 (N_7536,N_4257,N_5590);
nand U7537 (N_7537,N_4171,N_4378);
xnor U7538 (N_7538,N_4744,N_5153);
nand U7539 (N_7539,N_5523,N_4999);
nor U7540 (N_7540,N_4053,N_4649);
nor U7541 (N_7541,N_5740,N_4919);
or U7542 (N_7542,N_4617,N_5570);
nand U7543 (N_7543,N_5436,N_4534);
or U7544 (N_7544,N_5241,N_4507);
or U7545 (N_7545,N_5373,N_5284);
or U7546 (N_7546,N_5467,N_4805);
xor U7547 (N_7547,N_5504,N_4748);
nand U7548 (N_7548,N_4790,N_4020);
nor U7549 (N_7549,N_5346,N_4733);
nor U7550 (N_7550,N_4843,N_4859);
xnor U7551 (N_7551,N_4297,N_5626);
and U7552 (N_7552,N_5657,N_4203);
and U7553 (N_7553,N_4700,N_5076);
or U7554 (N_7554,N_5137,N_4855);
and U7555 (N_7555,N_4790,N_5693);
or U7556 (N_7556,N_5987,N_4085);
nand U7557 (N_7557,N_4252,N_5876);
and U7558 (N_7558,N_4087,N_4832);
xor U7559 (N_7559,N_5160,N_5703);
xnor U7560 (N_7560,N_5120,N_5213);
xnor U7561 (N_7561,N_5350,N_5818);
and U7562 (N_7562,N_4872,N_5496);
nor U7563 (N_7563,N_5817,N_4781);
nor U7564 (N_7564,N_4952,N_5987);
and U7565 (N_7565,N_4343,N_4655);
or U7566 (N_7566,N_4924,N_5820);
and U7567 (N_7567,N_4552,N_5500);
and U7568 (N_7568,N_5502,N_4625);
xor U7569 (N_7569,N_5514,N_5032);
or U7570 (N_7570,N_5817,N_4842);
nand U7571 (N_7571,N_4125,N_5453);
xnor U7572 (N_7572,N_4800,N_5749);
nand U7573 (N_7573,N_5873,N_4660);
nand U7574 (N_7574,N_4486,N_5970);
xnor U7575 (N_7575,N_4645,N_4812);
nor U7576 (N_7576,N_4262,N_5256);
and U7577 (N_7577,N_5719,N_4377);
or U7578 (N_7578,N_5354,N_4793);
nand U7579 (N_7579,N_5105,N_4766);
xnor U7580 (N_7580,N_4952,N_4299);
and U7581 (N_7581,N_4861,N_4553);
xnor U7582 (N_7582,N_4059,N_5342);
and U7583 (N_7583,N_4059,N_5837);
xnor U7584 (N_7584,N_4973,N_5093);
or U7585 (N_7585,N_4167,N_4761);
and U7586 (N_7586,N_4351,N_4745);
or U7587 (N_7587,N_4615,N_5222);
nand U7588 (N_7588,N_5320,N_5721);
nand U7589 (N_7589,N_5917,N_4672);
nand U7590 (N_7590,N_5316,N_5250);
nor U7591 (N_7591,N_5801,N_5111);
or U7592 (N_7592,N_4703,N_5383);
or U7593 (N_7593,N_5968,N_4978);
and U7594 (N_7594,N_4155,N_5144);
and U7595 (N_7595,N_4288,N_5817);
or U7596 (N_7596,N_4272,N_5704);
nand U7597 (N_7597,N_4975,N_4477);
or U7598 (N_7598,N_4727,N_5088);
or U7599 (N_7599,N_5866,N_4769);
nor U7600 (N_7600,N_4290,N_4140);
or U7601 (N_7601,N_4857,N_5695);
xor U7602 (N_7602,N_5514,N_5110);
or U7603 (N_7603,N_4235,N_4922);
nand U7604 (N_7604,N_5572,N_4967);
or U7605 (N_7605,N_5172,N_5564);
nand U7606 (N_7606,N_4474,N_5365);
or U7607 (N_7607,N_5406,N_5679);
nand U7608 (N_7608,N_5408,N_5574);
nand U7609 (N_7609,N_4027,N_5797);
and U7610 (N_7610,N_4424,N_4203);
nor U7611 (N_7611,N_5079,N_4680);
xor U7612 (N_7612,N_5227,N_5250);
nor U7613 (N_7613,N_4852,N_4419);
nand U7614 (N_7614,N_5356,N_5927);
and U7615 (N_7615,N_5499,N_5631);
or U7616 (N_7616,N_4597,N_5672);
or U7617 (N_7617,N_4683,N_5447);
nand U7618 (N_7618,N_5062,N_5104);
xnor U7619 (N_7619,N_4549,N_4875);
and U7620 (N_7620,N_5489,N_5527);
nor U7621 (N_7621,N_5862,N_4071);
nand U7622 (N_7622,N_5306,N_5940);
xor U7623 (N_7623,N_5387,N_5837);
xnor U7624 (N_7624,N_4590,N_5533);
or U7625 (N_7625,N_4265,N_4373);
or U7626 (N_7626,N_4426,N_4402);
and U7627 (N_7627,N_4710,N_4594);
and U7628 (N_7628,N_4717,N_4986);
or U7629 (N_7629,N_5070,N_4730);
or U7630 (N_7630,N_4001,N_4598);
xor U7631 (N_7631,N_4556,N_5613);
xor U7632 (N_7632,N_5593,N_5562);
nand U7633 (N_7633,N_4965,N_4860);
nand U7634 (N_7634,N_5125,N_5005);
xor U7635 (N_7635,N_4958,N_4016);
xnor U7636 (N_7636,N_5041,N_5106);
or U7637 (N_7637,N_5211,N_4428);
or U7638 (N_7638,N_5588,N_5143);
and U7639 (N_7639,N_5957,N_4818);
nand U7640 (N_7640,N_4175,N_5456);
xnor U7641 (N_7641,N_5368,N_4093);
and U7642 (N_7642,N_4970,N_4436);
nor U7643 (N_7643,N_4153,N_5796);
nor U7644 (N_7644,N_4363,N_4694);
or U7645 (N_7645,N_4765,N_5738);
nor U7646 (N_7646,N_4867,N_5574);
and U7647 (N_7647,N_5071,N_5016);
nor U7648 (N_7648,N_4805,N_5775);
xor U7649 (N_7649,N_4286,N_4574);
nor U7650 (N_7650,N_4791,N_4034);
or U7651 (N_7651,N_5673,N_5099);
nor U7652 (N_7652,N_5421,N_4522);
nor U7653 (N_7653,N_4061,N_5814);
or U7654 (N_7654,N_5595,N_5306);
nand U7655 (N_7655,N_5949,N_4394);
nand U7656 (N_7656,N_4843,N_4022);
and U7657 (N_7657,N_5604,N_4674);
xor U7658 (N_7658,N_4870,N_5970);
nor U7659 (N_7659,N_4832,N_4132);
nand U7660 (N_7660,N_4172,N_5736);
or U7661 (N_7661,N_4016,N_5546);
nor U7662 (N_7662,N_4839,N_4441);
and U7663 (N_7663,N_4297,N_4681);
nor U7664 (N_7664,N_4642,N_4252);
or U7665 (N_7665,N_4541,N_4710);
or U7666 (N_7666,N_5390,N_5099);
nand U7667 (N_7667,N_4872,N_5029);
xor U7668 (N_7668,N_4091,N_5738);
or U7669 (N_7669,N_4272,N_5877);
nor U7670 (N_7670,N_4484,N_5781);
or U7671 (N_7671,N_5313,N_5227);
and U7672 (N_7672,N_5582,N_4260);
nor U7673 (N_7673,N_4218,N_4610);
nor U7674 (N_7674,N_4062,N_4173);
or U7675 (N_7675,N_5318,N_4204);
and U7676 (N_7676,N_4189,N_5555);
xnor U7677 (N_7677,N_5038,N_5691);
xnor U7678 (N_7678,N_5576,N_5505);
nor U7679 (N_7679,N_5555,N_5930);
nand U7680 (N_7680,N_5300,N_4456);
and U7681 (N_7681,N_4008,N_5144);
nand U7682 (N_7682,N_5222,N_5041);
and U7683 (N_7683,N_4495,N_5952);
or U7684 (N_7684,N_5841,N_4993);
and U7685 (N_7685,N_4449,N_5672);
and U7686 (N_7686,N_5534,N_4594);
xor U7687 (N_7687,N_5523,N_5250);
and U7688 (N_7688,N_5518,N_4550);
and U7689 (N_7689,N_4865,N_4032);
or U7690 (N_7690,N_4043,N_5809);
nand U7691 (N_7691,N_5207,N_4622);
xor U7692 (N_7692,N_5230,N_4225);
xor U7693 (N_7693,N_5175,N_4716);
or U7694 (N_7694,N_5926,N_5905);
or U7695 (N_7695,N_4959,N_4702);
and U7696 (N_7696,N_5022,N_5652);
and U7697 (N_7697,N_5606,N_4757);
or U7698 (N_7698,N_5129,N_5436);
nor U7699 (N_7699,N_5143,N_4097);
and U7700 (N_7700,N_4535,N_5116);
xnor U7701 (N_7701,N_4379,N_4651);
nand U7702 (N_7702,N_5440,N_4500);
or U7703 (N_7703,N_5654,N_5421);
and U7704 (N_7704,N_5417,N_5303);
nand U7705 (N_7705,N_5639,N_5101);
or U7706 (N_7706,N_4950,N_5910);
nor U7707 (N_7707,N_4843,N_5475);
and U7708 (N_7708,N_5965,N_4154);
and U7709 (N_7709,N_5419,N_5220);
nand U7710 (N_7710,N_5497,N_5222);
or U7711 (N_7711,N_4346,N_5056);
xor U7712 (N_7712,N_5337,N_4065);
xnor U7713 (N_7713,N_5620,N_5481);
nor U7714 (N_7714,N_5555,N_5744);
nor U7715 (N_7715,N_5349,N_5675);
xor U7716 (N_7716,N_4099,N_4857);
or U7717 (N_7717,N_4351,N_4641);
xor U7718 (N_7718,N_4117,N_5425);
nand U7719 (N_7719,N_5007,N_5200);
nor U7720 (N_7720,N_5511,N_4798);
xnor U7721 (N_7721,N_5917,N_4989);
xnor U7722 (N_7722,N_4875,N_5355);
or U7723 (N_7723,N_4249,N_5041);
nor U7724 (N_7724,N_5081,N_4030);
or U7725 (N_7725,N_4608,N_5836);
nand U7726 (N_7726,N_5959,N_4732);
and U7727 (N_7727,N_4889,N_5283);
nand U7728 (N_7728,N_5519,N_5249);
and U7729 (N_7729,N_5694,N_5997);
nor U7730 (N_7730,N_5344,N_4155);
nor U7731 (N_7731,N_5884,N_5427);
nand U7732 (N_7732,N_5024,N_5013);
xnor U7733 (N_7733,N_4625,N_4956);
nor U7734 (N_7734,N_5766,N_4725);
nor U7735 (N_7735,N_4875,N_4820);
xor U7736 (N_7736,N_4282,N_4258);
nor U7737 (N_7737,N_4109,N_5633);
nand U7738 (N_7738,N_5165,N_5830);
and U7739 (N_7739,N_4069,N_4093);
and U7740 (N_7740,N_5740,N_5631);
or U7741 (N_7741,N_5666,N_5752);
or U7742 (N_7742,N_5586,N_4993);
and U7743 (N_7743,N_5858,N_5255);
or U7744 (N_7744,N_4955,N_5402);
or U7745 (N_7745,N_5044,N_5384);
and U7746 (N_7746,N_4849,N_5993);
xnor U7747 (N_7747,N_4201,N_4655);
nor U7748 (N_7748,N_4115,N_4482);
and U7749 (N_7749,N_5832,N_4903);
nand U7750 (N_7750,N_4303,N_5773);
nor U7751 (N_7751,N_5555,N_4136);
xor U7752 (N_7752,N_4421,N_4950);
or U7753 (N_7753,N_5224,N_5250);
nand U7754 (N_7754,N_4961,N_5921);
nand U7755 (N_7755,N_5987,N_5679);
nand U7756 (N_7756,N_4171,N_5873);
nor U7757 (N_7757,N_5418,N_5104);
xor U7758 (N_7758,N_4999,N_5660);
and U7759 (N_7759,N_5624,N_5376);
or U7760 (N_7760,N_4059,N_5729);
nand U7761 (N_7761,N_4664,N_4567);
nor U7762 (N_7762,N_4736,N_4430);
nor U7763 (N_7763,N_4668,N_4901);
or U7764 (N_7764,N_4651,N_4241);
nand U7765 (N_7765,N_5035,N_5924);
and U7766 (N_7766,N_5497,N_4908);
and U7767 (N_7767,N_5018,N_5915);
or U7768 (N_7768,N_4056,N_5060);
nor U7769 (N_7769,N_4549,N_5668);
or U7770 (N_7770,N_5865,N_4284);
and U7771 (N_7771,N_4695,N_4842);
nand U7772 (N_7772,N_4019,N_4426);
xor U7773 (N_7773,N_5177,N_4198);
nor U7774 (N_7774,N_5754,N_5034);
or U7775 (N_7775,N_5134,N_4473);
nand U7776 (N_7776,N_5659,N_4633);
and U7777 (N_7777,N_4199,N_5378);
nor U7778 (N_7778,N_4370,N_5050);
and U7779 (N_7779,N_5542,N_5103);
or U7780 (N_7780,N_5487,N_5991);
and U7781 (N_7781,N_4197,N_5272);
nor U7782 (N_7782,N_5878,N_5535);
xor U7783 (N_7783,N_4164,N_4163);
and U7784 (N_7784,N_4113,N_5344);
nor U7785 (N_7785,N_5599,N_4037);
and U7786 (N_7786,N_4971,N_5089);
and U7787 (N_7787,N_5394,N_5734);
nor U7788 (N_7788,N_5144,N_4767);
or U7789 (N_7789,N_4457,N_5564);
nor U7790 (N_7790,N_5769,N_4127);
and U7791 (N_7791,N_5139,N_5164);
nor U7792 (N_7792,N_4095,N_5924);
or U7793 (N_7793,N_4014,N_4191);
or U7794 (N_7794,N_4152,N_5585);
nor U7795 (N_7795,N_5472,N_5235);
or U7796 (N_7796,N_5990,N_4136);
and U7797 (N_7797,N_4711,N_5403);
nand U7798 (N_7798,N_4640,N_5545);
xnor U7799 (N_7799,N_5099,N_4286);
xnor U7800 (N_7800,N_4458,N_4478);
and U7801 (N_7801,N_5049,N_4995);
or U7802 (N_7802,N_5198,N_5594);
nand U7803 (N_7803,N_5010,N_5924);
nor U7804 (N_7804,N_5786,N_5811);
nand U7805 (N_7805,N_5035,N_5608);
and U7806 (N_7806,N_4246,N_4255);
nand U7807 (N_7807,N_5930,N_5881);
xor U7808 (N_7808,N_5484,N_5757);
and U7809 (N_7809,N_4142,N_4408);
or U7810 (N_7810,N_5329,N_4531);
nor U7811 (N_7811,N_4885,N_4652);
and U7812 (N_7812,N_5462,N_5161);
and U7813 (N_7813,N_4550,N_5907);
or U7814 (N_7814,N_4829,N_5124);
xor U7815 (N_7815,N_5391,N_4128);
and U7816 (N_7816,N_5763,N_5437);
nand U7817 (N_7817,N_5243,N_4683);
xnor U7818 (N_7818,N_4963,N_4020);
xnor U7819 (N_7819,N_5538,N_5128);
and U7820 (N_7820,N_5775,N_4537);
xor U7821 (N_7821,N_4531,N_5035);
xor U7822 (N_7822,N_5306,N_4135);
xnor U7823 (N_7823,N_4673,N_4758);
nand U7824 (N_7824,N_4070,N_5807);
nor U7825 (N_7825,N_4825,N_5610);
nor U7826 (N_7826,N_5145,N_4807);
and U7827 (N_7827,N_4952,N_4846);
nor U7828 (N_7828,N_5807,N_4488);
nor U7829 (N_7829,N_5737,N_5657);
nand U7830 (N_7830,N_4063,N_5811);
nor U7831 (N_7831,N_5808,N_5865);
or U7832 (N_7832,N_5412,N_4407);
and U7833 (N_7833,N_4146,N_4585);
nor U7834 (N_7834,N_5524,N_5222);
nor U7835 (N_7835,N_5359,N_5539);
and U7836 (N_7836,N_5763,N_5820);
nor U7837 (N_7837,N_5285,N_4412);
and U7838 (N_7838,N_5337,N_5866);
or U7839 (N_7839,N_4637,N_4835);
and U7840 (N_7840,N_5585,N_5679);
and U7841 (N_7841,N_4097,N_4387);
and U7842 (N_7842,N_5762,N_5305);
xnor U7843 (N_7843,N_4310,N_5278);
xnor U7844 (N_7844,N_4001,N_4399);
and U7845 (N_7845,N_4188,N_5000);
or U7846 (N_7846,N_5200,N_4850);
nor U7847 (N_7847,N_4802,N_4932);
or U7848 (N_7848,N_4764,N_5649);
and U7849 (N_7849,N_5337,N_5950);
and U7850 (N_7850,N_5966,N_4351);
nor U7851 (N_7851,N_5058,N_5954);
xor U7852 (N_7852,N_5737,N_5676);
or U7853 (N_7853,N_4655,N_4821);
xnor U7854 (N_7854,N_4859,N_5429);
nor U7855 (N_7855,N_4686,N_4306);
and U7856 (N_7856,N_5682,N_5199);
and U7857 (N_7857,N_5723,N_4471);
nand U7858 (N_7858,N_4440,N_4634);
or U7859 (N_7859,N_4432,N_4874);
nor U7860 (N_7860,N_5522,N_5224);
nand U7861 (N_7861,N_5170,N_5588);
and U7862 (N_7862,N_5287,N_5308);
and U7863 (N_7863,N_4710,N_4284);
nor U7864 (N_7864,N_4747,N_4063);
and U7865 (N_7865,N_4105,N_4643);
and U7866 (N_7866,N_4205,N_4479);
nor U7867 (N_7867,N_4536,N_4720);
and U7868 (N_7868,N_4667,N_5012);
nand U7869 (N_7869,N_4693,N_4850);
nor U7870 (N_7870,N_5149,N_4203);
nand U7871 (N_7871,N_4640,N_5427);
and U7872 (N_7872,N_5075,N_4152);
xor U7873 (N_7873,N_5683,N_5835);
nand U7874 (N_7874,N_5219,N_5758);
nand U7875 (N_7875,N_4308,N_4870);
or U7876 (N_7876,N_5334,N_5219);
and U7877 (N_7877,N_4267,N_4034);
and U7878 (N_7878,N_5229,N_4036);
or U7879 (N_7879,N_4834,N_4298);
nand U7880 (N_7880,N_4400,N_5899);
and U7881 (N_7881,N_4483,N_5380);
xor U7882 (N_7882,N_5912,N_4863);
nand U7883 (N_7883,N_4206,N_5216);
xor U7884 (N_7884,N_5214,N_4810);
and U7885 (N_7885,N_5764,N_5469);
or U7886 (N_7886,N_4255,N_5974);
nand U7887 (N_7887,N_4000,N_5318);
or U7888 (N_7888,N_4976,N_5251);
or U7889 (N_7889,N_5701,N_5199);
xnor U7890 (N_7890,N_4842,N_5081);
nand U7891 (N_7891,N_4081,N_4876);
nand U7892 (N_7892,N_4596,N_5581);
nand U7893 (N_7893,N_5962,N_4411);
or U7894 (N_7894,N_5651,N_4303);
xnor U7895 (N_7895,N_5165,N_5554);
and U7896 (N_7896,N_5461,N_4713);
and U7897 (N_7897,N_5327,N_4132);
xor U7898 (N_7898,N_4128,N_4234);
and U7899 (N_7899,N_4635,N_4849);
or U7900 (N_7900,N_4741,N_5636);
and U7901 (N_7901,N_4047,N_4817);
or U7902 (N_7902,N_5750,N_4985);
or U7903 (N_7903,N_4831,N_5857);
and U7904 (N_7904,N_4383,N_5440);
nand U7905 (N_7905,N_4075,N_4784);
or U7906 (N_7906,N_4862,N_5357);
and U7907 (N_7907,N_4517,N_5083);
nor U7908 (N_7908,N_4606,N_5076);
nand U7909 (N_7909,N_4293,N_4545);
nor U7910 (N_7910,N_4047,N_5546);
or U7911 (N_7911,N_4942,N_5865);
nor U7912 (N_7912,N_4337,N_4175);
or U7913 (N_7913,N_5831,N_4679);
nand U7914 (N_7914,N_4068,N_5097);
xnor U7915 (N_7915,N_5946,N_4821);
nand U7916 (N_7916,N_5017,N_4072);
or U7917 (N_7917,N_4698,N_4225);
nand U7918 (N_7918,N_5979,N_5611);
nand U7919 (N_7919,N_4926,N_4274);
nand U7920 (N_7920,N_4807,N_4569);
and U7921 (N_7921,N_5897,N_5603);
and U7922 (N_7922,N_4286,N_5435);
and U7923 (N_7923,N_5743,N_4912);
nor U7924 (N_7924,N_5769,N_4386);
nand U7925 (N_7925,N_4115,N_4991);
nor U7926 (N_7926,N_4089,N_5813);
or U7927 (N_7927,N_5039,N_4061);
and U7928 (N_7928,N_5598,N_5362);
nand U7929 (N_7929,N_5397,N_5930);
xor U7930 (N_7930,N_4474,N_4245);
or U7931 (N_7931,N_4556,N_4639);
nor U7932 (N_7932,N_5627,N_4380);
xor U7933 (N_7933,N_5470,N_5416);
nor U7934 (N_7934,N_4541,N_4662);
or U7935 (N_7935,N_5299,N_5242);
nand U7936 (N_7936,N_4628,N_5013);
xor U7937 (N_7937,N_4034,N_5169);
or U7938 (N_7938,N_4170,N_4397);
xnor U7939 (N_7939,N_5694,N_4870);
nor U7940 (N_7940,N_4684,N_4542);
and U7941 (N_7941,N_4197,N_4001);
xnor U7942 (N_7942,N_4476,N_4055);
nor U7943 (N_7943,N_5579,N_4405);
and U7944 (N_7944,N_4440,N_4829);
or U7945 (N_7945,N_4872,N_5192);
xnor U7946 (N_7946,N_5085,N_4562);
nor U7947 (N_7947,N_5713,N_5463);
nand U7948 (N_7948,N_5064,N_5978);
nor U7949 (N_7949,N_5528,N_4959);
nand U7950 (N_7950,N_4758,N_4111);
and U7951 (N_7951,N_5557,N_4534);
and U7952 (N_7952,N_4901,N_5766);
nand U7953 (N_7953,N_5406,N_5742);
nor U7954 (N_7954,N_5515,N_5469);
nand U7955 (N_7955,N_5177,N_4943);
or U7956 (N_7956,N_4635,N_4522);
or U7957 (N_7957,N_4999,N_5719);
nand U7958 (N_7958,N_4901,N_5337);
or U7959 (N_7959,N_5736,N_4870);
nor U7960 (N_7960,N_4570,N_4314);
and U7961 (N_7961,N_4358,N_5775);
xnor U7962 (N_7962,N_5716,N_5954);
nand U7963 (N_7963,N_5109,N_4315);
xnor U7964 (N_7964,N_5277,N_4296);
nand U7965 (N_7965,N_5035,N_5084);
or U7966 (N_7966,N_4132,N_5931);
nor U7967 (N_7967,N_4993,N_4226);
nand U7968 (N_7968,N_4664,N_5140);
nor U7969 (N_7969,N_5696,N_5094);
or U7970 (N_7970,N_4980,N_4188);
nor U7971 (N_7971,N_5602,N_5857);
or U7972 (N_7972,N_4870,N_4097);
and U7973 (N_7973,N_5047,N_5014);
nand U7974 (N_7974,N_4986,N_4745);
and U7975 (N_7975,N_5599,N_4656);
or U7976 (N_7976,N_4762,N_5597);
xnor U7977 (N_7977,N_5693,N_5600);
and U7978 (N_7978,N_4800,N_4677);
or U7979 (N_7979,N_5246,N_5936);
and U7980 (N_7980,N_5086,N_4351);
nor U7981 (N_7981,N_4505,N_4315);
nand U7982 (N_7982,N_5638,N_5789);
xor U7983 (N_7983,N_5328,N_5423);
xnor U7984 (N_7984,N_4079,N_4534);
xor U7985 (N_7985,N_5126,N_4949);
nor U7986 (N_7986,N_5436,N_5604);
xnor U7987 (N_7987,N_4802,N_5695);
xnor U7988 (N_7988,N_5165,N_5672);
nor U7989 (N_7989,N_4944,N_4153);
xnor U7990 (N_7990,N_5797,N_4684);
nand U7991 (N_7991,N_5093,N_5298);
xnor U7992 (N_7992,N_4556,N_4862);
or U7993 (N_7993,N_4845,N_4174);
or U7994 (N_7994,N_5567,N_5286);
nand U7995 (N_7995,N_4887,N_5035);
nor U7996 (N_7996,N_5046,N_5719);
xor U7997 (N_7997,N_4531,N_5867);
nand U7998 (N_7998,N_5275,N_5008);
nor U7999 (N_7999,N_5779,N_5909);
xnor U8000 (N_8000,N_6874,N_7561);
nand U8001 (N_8001,N_6551,N_7190);
and U8002 (N_8002,N_6878,N_6369);
nand U8003 (N_8003,N_6402,N_7503);
nand U8004 (N_8004,N_6965,N_6389);
xor U8005 (N_8005,N_7225,N_7095);
nor U8006 (N_8006,N_6920,N_6271);
or U8007 (N_8007,N_7722,N_6054);
nor U8008 (N_8008,N_7299,N_7821);
xnor U8009 (N_8009,N_6269,N_6562);
nand U8010 (N_8010,N_7264,N_7427);
nor U8011 (N_8011,N_7471,N_7271);
and U8012 (N_8012,N_7774,N_6118);
and U8013 (N_8013,N_7795,N_7495);
and U8014 (N_8014,N_7933,N_7813);
nand U8015 (N_8015,N_6895,N_6342);
and U8016 (N_8016,N_6711,N_6262);
nand U8017 (N_8017,N_6749,N_6891);
or U8018 (N_8018,N_6537,N_6468);
and U8019 (N_8019,N_6351,N_6481);
xor U8020 (N_8020,N_7882,N_7545);
xor U8021 (N_8021,N_6632,N_7581);
nor U8022 (N_8022,N_7684,N_7201);
nand U8023 (N_8023,N_7765,N_6638);
and U8024 (N_8024,N_7466,N_7219);
and U8025 (N_8025,N_7409,N_7000);
nor U8026 (N_8026,N_6970,N_6676);
and U8027 (N_8027,N_7686,N_7006);
xor U8028 (N_8028,N_7300,N_6267);
and U8029 (N_8029,N_6794,N_7407);
nand U8030 (N_8030,N_6786,N_6046);
xor U8031 (N_8031,N_6295,N_7568);
xnor U8032 (N_8032,N_7717,N_6339);
or U8033 (N_8033,N_7517,N_7314);
nand U8034 (N_8034,N_6502,N_6083);
and U8035 (N_8035,N_6792,N_6966);
and U8036 (N_8036,N_6325,N_7163);
or U8037 (N_8037,N_7158,N_7964);
nor U8038 (N_8038,N_6281,N_6958);
nand U8039 (N_8039,N_7560,N_6187);
nand U8040 (N_8040,N_6013,N_6565);
xnor U8041 (N_8041,N_7154,N_7856);
nor U8042 (N_8042,N_6388,N_7479);
or U8043 (N_8043,N_6020,N_7376);
and U8044 (N_8044,N_7824,N_6939);
or U8045 (N_8045,N_6748,N_7655);
xor U8046 (N_8046,N_6735,N_7372);
nor U8047 (N_8047,N_7507,N_6041);
nand U8048 (N_8048,N_6071,N_7604);
nor U8049 (N_8049,N_7391,N_7910);
and U8050 (N_8050,N_7249,N_6104);
xor U8051 (N_8051,N_6964,N_6807);
xor U8052 (N_8052,N_7513,N_6933);
xnor U8053 (N_8053,N_7962,N_7169);
and U8054 (N_8054,N_6961,N_7798);
nor U8055 (N_8055,N_6151,N_7067);
and U8056 (N_8056,N_7961,N_7605);
nor U8057 (N_8057,N_6882,N_6650);
nand U8058 (N_8058,N_7024,N_7540);
and U8059 (N_8059,N_6095,N_7834);
nand U8060 (N_8060,N_7414,N_6808);
nand U8061 (N_8061,N_7213,N_7452);
and U8062 (N_8062,N_6084,N_6226);
nand U8063 (N_8063,N_6304,N_6609);
xor U8064 (N_8064,N_7562,N_6854);
and U8065 (N_8065,N_7426,N_7442);
xor U8066 (N_8066,N_7701,N_7234);
xor U8067 (N_8067,N_7959,N_6330);
xnor U8068 (N_8068,N_7412,N_6985);
nand U8069 (N_8069,N_7385,N_7642);
xnor U8070 (N_8070,N_7504,N_7535);
or U8071 (N_8071,N_7853,N_6991);
nor U8072 (N_8072,N_7134,N_7886);
or U8073 (N_8073,N_7963,N_6288);
nor U8074 (N_8074,N_7901,N_7111);
or U8075 (N_8075,N_6706,N_6850);
and U8076 (N_8076,N_6908,N_6027);
or U8077 (N_8077,N_7999,N_6193);
nand U8078 (N_8078,N_7229,N_6012);
nor U8079 (N_8079,N_7100,N_6846);
nand U8080 (N_8080,N_7365,N_6873);
nand U8081 (N_8081,N_6513,N_6756);
or U8082 (N_8082,N_7913,N_7924);
xor U8083 (N_8083,N_7986,N_7761);
nand U8084 (N_8084,N_7051,N_7510);
and U8085 (N_8085,N_6040,N_7716);
or U8086 (N_8086,N_7070,N_7662);
nand U8087 (N_8087,N_7278,N_6941);
xor U8088 (N_8088,N_6441,N_6569);
xor U8089 (N_8089,N_6107,N_6254);
and U8090 (N_8090,N_6541,N_7773);
and U8091 (N_8091,N_6936,N_7081);
and U8092 (N_8092,N_6437,N_7152);
or U8093 (N_8093,N_6761,N_7073);
nand U8094 (N_8094,N_7596,N_7276);
nand U8095 (N_8095,N_7989,N_6762);
xnor U8096 (N_8096,N_6333,N_7671);
nand U8097 (N_8097,N_6345,N_7354);
nor U8098 (N_8098,N_6595,N_7657);
and U8099 (N_8099,N_7436,N_7832);
or U8100 (N_8100,N_7284,N_7666);
nor U8101 (N_8101,N_7233,N_6431);
nor U8102 (N_8102,N_6392,N_7810);
nor U8103 (N_8103,N_7392,N_7450);
nand U8104 (N_8104,N_6615,N_6772);
xnor U8105 (N_8105,N_6840,N_6935);
nor U8106 (N_8106,N_7970,N_7891);
and U8107 (N_8107,N_6172,N_6272);
nand U8108 (N_8108,N_6754,N_6539);
and U8109 (N_8109,N_7124,N_6328);
xnor U8110 (N_8110,N_7514,N_6015);
xnor U8111 (N_8111,N_7651,N_6899);
or U8112 (N_8112,N_6136,N_6394);
nand U8113 (N_8113,N_6930,N_6732);
and U8114 (N_8114,N_6278,N_6542);
or U8115 (N_8115,N_6633,N_7415);
nor U8116 (N_8116,N_6249,N_7681);
nor U8117 (N_8117,N_7413,N_6234);
and U8118 (N_8118,N_6209,N_6725);
and U8119 (N_8119,N_7456,N_7367);
nor U8120 (N_8120,N_7950,N_6386);
nand U8121 (N_8121,N_6062,N_6189);
or U8122 (N_8122,N_6163,N_7453);
nand U8123 (N_8123,N_6162,N_6750);
or U8124 (N_8124,N_6645,N_7746);
or U8125 (N_8125,N_7389,N_7439);
nand U8126 (N_8126,N_7378,N_6420);
xor U8127 (N_8127,N_6397,N_6098);
nand U8128 (N_8128,N_7350,N_6166);
nor U8129 (N_8129,N_7610,N_7240);
xor U8130 (N_8130,N_6309,N_6547);
xor U8131 (N_8131,N_7207,N_6666);
nand U8132 (N_8132,N_7335,N_7965);
nor U8133 (N_8133,N_7870,N_7725);
and U8134 (N_8134,N_6043,N_7622);
nand U8135 (N_8135,N_7929,N_6925);
xor U8136 (N_8136,N_6391,N_6023);
xnor U8137 (N_8137,N_7328,N_7546);
or U8138 (N_8138,N_6496,N_7862);
nor U8139 (N_8139,N_7630,N_6816);
or U8140 (N_8140,N_6212,N_7582);
xor U8141 (N_8141,N_7290,N_6485);
nand U8142 (N_8142,N_7098,N_7855);
nand U8143 (N_8143,N_7296,N_7358);
and U8144 (N_8144,N_7019,N_6717);
nand U8145 (N_8145,N_6753,N_7990);
or U8146 (N_8146,N_7789,N_7611);
xnor U8147 (N_8147,N_6948,N_7682);
or U8148 (N_8148,N_6892,N_6443);
nor U8149 (N_8149,N_6450,N_7735);
and U8150 (N_8150,N_6852,N_7160);
and U8151 (N_8151,N_6442,N_6059);
xnor U8152 (N_8152,N_7905,N_6553);
xor U8153 (N_8153,N_7659,N_7762);
and U8154 (N_8154,N_6463,N_6233);
nand U8155 (N_8155,N_7083,N_7275);
and U8156 (N_8156,N_7108,N_7748);
nand U8157 (N_8157,N_7036,N_6604);
or U8158 (N_8158,N_6406,N_7918);
xor U8159 (N_8159,N_6740,N_6960);
nand U8160 (N_8160,N_6672,N_7180);
nand U8161 (N_8161,N_7680,N_7629);
nand U8162 (N_8162,N_6310,N_6074);
or U8163 (N_8163,N_7008,N_7902);
nand U8164 (N_8164,N_7491,N_7723);
nand U8165 (N_8165,N_7068,N_6866);
xor U8166 (N_8166,N_7075,N_7114);
nand U8167 (N_8167,N_6837,N_7899);
nand U8168 (N_8168,N_7074,N_7281);
nand U8169 (N_8169,N_6584,N_7858);
xor U8170 (N_8170,N_7028,N_7884);
or U8171 (N_8171,N_7486,N_7548);
or U8172 (N_8172,N_7488,N_6683);
nand U8173 (N_8173,N_6534,N_6428);
or U8174 (N_8174,N_6824,N_7802);
xnor U8175 (N_8175,N_7836,N_6715);
nor U8176 (N_8176,N_6419,N_7565);
xnor U8177 (N_8177,N_7742,N_6952);
nand U8178 (N_8178,N_7804,N_6649);
nor U8179 (N_8179,N_7211,N_6188);
or U8180 (N_8180,N_6282,N_6275);
and U8181 (N_8181,N_7845,N_7643);
and U8182 (N_8182,N_7692,N_6779);
xor U8183 (N_8183,N_7032,N_6101);
or U8184 (N_8184,N_6079,N_6512);
or U8185 (N_8185,N_7338,N_7265);
nand U8186 (N_8186,N_7625,N_7975);
nor U8187 (N_8187,N_7112,N_6549);
nand U8188 (N_8188,N_6360,N_7880);
xnor U8189 (N_8189,N_6865,N_6993);
nor U8190 (N_8190,N_6917,N_7776);
nand U8191 (N_8191,N_6491,N_7307);
xnor U8192 (N_8192,N_6752,N_7137);
and U8193 (N_8193,N_6220,N_7731);
or U8194 (N_8194,N_7405,N_6603);
xnor U8195 (N_8195,N_6413,N_6247);
and U8196 (N_8196,N_6744,N_6287);
nor U8197 (N_8197,N_6540,N_7669);
and U8198 (N_8198,N_6456,N_7644);
nand U8199 (N_8199,N_7288,N_6144);
or U8200 (N_8200,N_6660,N_7595);
or U8201 (N_8201,N_7598,N_7472);
or U8202 (N_8202,N_7909,N_7697);
and U8203 (N_8203,N_7947,N_7764);
nor U8204 (N_8204,N_6962,N_7865);
nor U8205 (N_8205,N_7418,N_6938);
nand U8206 (N_8206,N_7958,N_7849);
xnor U8207 (N_8207,N_6574,N_7345);
or U8208 (N_8208,N_6704,N_6528);
nand U8209 (N_8209,N_6783,N_6670);
xor U8210 (N_8210,N_6695,N_6306);
and U8211 (N_8211,N_6769,N_6110);
nand U8212 (N_8212,N_7583,N_7529);
and U8213 (N_8213,N_7664,N_6257);
nand U8214 (N_8214,N_6289,N_6228);
or U8215 (N_8215,N_7547,N_7755);
and U8216 (N_8216,N_7976,N_6222);
or U8217 (N_8217,N_7474,N_7661);
or U8218 (N_8218,N_6208,N_7592);
nor U8219 (N_8219,N_7558,N_7734);
and U8220 (N_8220,N_7982,N_6698);
and U8221 (N_8221,N_6308,N_6571);
and U8222 (N_8222,N_7874,N_6346);
or U8223 (N_8223,N_7624,N_6157);
and U8224 (N_8224,N_6500,N_6980);
and U8225 (N_8225,N_7985,N_7291);
nand U8226 (N_8226,N_7030,N_7822);
and U8227 (N_8227,N_7919,N_7706);
nor U8228 (N_8228,N_6517,N_7317);
or U8229 (N_8229,N_7967,N_7770);
or U8230 (N_8230,N_7665,N_7041);
and U8231 (N_8231,N_6582,N_6694);
xor U8232 (N_8232,N_6489,N_7194);
or U8233 (N_8233,N_7347,N_6199);
nand U8234 (N_8234,N_7013,N_7612);
or U8235 (N_8235,N_6155,N_7091);
nand U8236 (N_8236,N_7104,N_7779);
or U8237 (N_8237,N_6021,N_7893);
nor U8238 (N_8238,N_6253,N_6176);
nor U8239 (N_8239,N_6826,N_7702);
nor U8240 (N_8240,N_7301,N_6194);
nand U8241 (N_8241,N_7873,N_7012);
xor U8242 (N_8242,N_7331,N_7839);
or U8243 (N_8243,N_7980,N_7386);
nor U8244 (N_8244,N_7177,N_6058);
nor U8245 (N_8245,N_6085,N_7071);
or U8246 (N_8246,N_7618,N_7519);
and U8247 (N_8247,N_7383,N_6529);
or U8248 (N_8248,N_6832,N_7241);
and U8249 (N_8249,N_7156,N_7210);
xnor U8250 (N_8250,N_6651,N_7903);
xnor U8251 (N_8251,N_7594,N_7401);
nor U8252 (N_8252,N_7628,N_7252);
nor U8253 (N_8253,N_6432,N_7876);
nand U8254 (N_8254,N_7232,N_7550);
xnor U8255 (N_8255,N_7732,N_6738);
nor U8256 (N_8256,N_7602,N_6094);
nor U8257 (N_8257,N_7228,N_6870);
nor U8258 (N_8258,N_7033,N_6474);
nor U8259 (N_8259,N_6338,N_6192);
nor U8260 (N_8260,N_6305,N_6904);
xnor U8261 (N_8261,N_7410,N_6602);
or U8262 (N_8262,N_6697,N_6108);
xnor U8263 (N_8263,N_7390,N_7621);
or U8264 (N_8264,N_6379,N_6567);
nand U8265 (N_8265,N_7733,N_7786);
xor U8266 (N_8266,N_6862,N_7946);
xor U8267 (N_8267,N_6376,N_6995);
nand U8268 (N_8268,N_7738,N_7841);
nor U8269 (N_8269,N_6037,N_7090);
xor U8270 (N_8270,N_7185,N_7448);
nand U8271 (N_8271,N_7772,N_6302);
nor U8272 (N_8272,N_6032,N_7174);
xor U8273 (N_8273,N_6374,N_6035);
xor U8274 (N_8274,N_6324,N_7193);
nand U8275 (N_8275,N_6230,N_6564);
or U8276 (N_8276,N_7783,N_7522);
nor U8277 (N_8277,N_6216,N_7775);
and U8278 (N_8278,N_6736,N_6909);
and U8279 (N_8279,N_7767,N_7343);
nor U8280 (N_8280,N_7586,N_7784);
xor U8281 (N_8281,N_6344,N_6130);
nand U8282 (N_8282,N_7246,N_6644);
or U8283 (N_8283,N_6906,N_6550);
nand U8284 (N_8284,N_6334,N_7147);
nor U8285 (N_8285,N_6703,N_7708);
nand U8286 (N_8286,N_7237,N_6025);
and U8287 (N_8287,N_6531,N_7633);
or U8288 (N_8288,N_6242,N_7992);
nand U8289 (N_8289,N_7266,N_7554);
nand U8290 (N_8290,N_6461,N_7653);
and U8291 (N_8291,N_7029,N_7741);
nand U8292 (N_8292,N_6219,N_6237);
nand U8293 (N_8293,N_6536,N_6781);
nor U8294 (N_8294,N_7105,N_6957);
or U8295 (N_8295,N_7502,N_7142);
xnor U8296 (N_8296,N_6579,N_7438);
or U8297 (N_8297,N_6987,N_7782);
or U8298 (N_8298,N_6169,N_7200);
nor U8299 (N_8299,N_6092,N_6818);
and U8300 (N_8300,N_6211,N_6538);
nand U8301 (N_8301,N_6598,N_6280);
nor U8302 (N_8302,N_7256,N_6853);
and U8303 (N_8303,N_6887,N_7212);
nand U8304 (N_8304,N_6778,N_6875);
nor U8305 (N_8305,N_6894,N_7601);
and U8306 (N_8306,N_7539,N_7167);
and U8307 (N_8307,N_6239,N_6950);
nor U8308 (N_8308,N_7854,N_6326);
or U8309 (N_8309,N_7875,N_7476);
and U8310 (N_8310,N_6712,N_7393);
nand U8311 (N_8311,N_6967,N_7805);
xor U8312 (N_8312,N_6469,N_6614);
xor U8313 (N_8313,N_6149,N_6066);
and U8314 (N_8314,N_6861,N_6733);
xnor U8315 (N_8315,N_7254,N_6998);
nand U8316 (N_8316,N_6024,N_6204);
xor U8317 (N_8317,N_7788,N_7205);
or U8318 (N_8318,N_7198,N_7058);
xor U8319 (N_8319,N_7316,N_7526);
or U8320 (N_8320,N_6544,N_7569);
xor U8321 (N_8321,N_6341,N_6440);
nor U8322 (N_8322,N_7370,N_7710);
nand U8323 (N_8323,N_6064,N_6116);
and U8324 (N_8324,N_6159,N_6659);
or U8325 (N_8325,N_7831,N_6809);
nor U8326 (N_8326,N_7458,N_6864);
and U8327 (N_8327,N_7750,N_6922);
or U8328 (N_8328,N_7261,N_6634);
xnor U8329 (N_8329,N_6820,N_6896);
or U8330 (N_8330,N_6273,N_7585);
xor U8331 (N_8331,N_7727,N_6364);
nand U8332 (N_8332,N_7340,N_6765);
xnor U8333 (N_8333,N_7400,N_7184);
or U8334 (N_8334,N_7110,N_7815);
xor U8335 (N_8335,N_6298,N_6158);
and U8336 (N_8336,N_6583,N_7294);
nand U8337 (N_8337,N_6708,N_7096);
nor U8338 (N_8338,N_6774,N_7923);
xor U8339 (N_8339,N_7803,N_7463);
and U8340 (N_8340,N_6625,N_6251);
or U8341 (N_8341,N_7530,N_6990);
or U8342 (N_8342,N_6884,N_6042);
xnor U8343 (N_8343,N_6924,N_6377);
xor U8344 (N_8344,N_6974,N_7286);
nor U8345 (N_8345,N_7675,N_7915);
or U8346 (N_8346,N_6841,N_6332);
nand U8347 (N_8347,N_6883,N_6051);
and U8348 (N_8348,N_7336,N_7082);
and U8349 (N_8349,N_7171,N_7660);
or U8350 (N_8350,N_6405,N_6353);
or U8351 (N_8351,N_6179,N_7217);
nand U8352 (N_8352,N_6102,N_6624);
nand U8353 (N_8353,N_6594,N_7878);
xor U8354 (N_8354,N_6438,N_7140);
and U8355 (N_8355,N_7640,N_7049);
nand U8356 (N_8356,N_6038,N_7189);
nand U8357 (N_8357,N_6331,N_7215);
nor U8358 (N_8358,N_7864,N_6642);
nor U8359 (N_8359,N_7079,N_7981);
or U8360 (N_8360,N_6141,N_6137);
xor U8361 (N_8361,N_6050,N_6823);
or U8362 (N_8362,N_6848,N_7443);
xnor U8363 (N_8363,N_7126,N_6857);
xnor U8364 (N_8364,N_7859,N_7149);
or U8365 (N_8365,N_6819,N_7144);
or U8366 (N_8366,N_6039,N_7120);
or U8367 (N_8367,N_6297,N_6073);
nor U8368 (N_8368,N_7176,N_6177);
xnor U8369 (N_8369,N_7801,N_6983);
and U8370 (N_8370,N_6727,N_7877);
or U8371 (N_8371,N_6688,N_6473);
nand U8372 (N_8372,N_7943,N_6398);
nor U8373 (N_8373,N_7785,N_7097);
and U8374 (N_8374,N_7850,N_7035);
and U8375 (N_8375,N_6843,N_7590);
nand U8376 (N_8376,N_6775,N_6975);
nor U8377 (N_8377,N_6718,N_7009);
or U8378 (N_8378,N_6476,N_6248);
nand U8379 (N_8379,N_6266,N_6796);
and U8380 (N_8380,N_6618,N_7753);
xor U8381 (N_8381,N_7465,N_6294);
xor U8382 (N_8382,N_7871,N_6689);
xnor U8383 (N_8383,N_6448,N_6019);
and U8384 (N_8384,N_6988,N_7066);
or U8385 (N_8385,N_6548,N_6655);
or U8386 (N_8386,N_7928,N_6396);
nor U8387 (N_8387,N_6480,N_6352);
nand U8388 (N_8388,N_6726,N_6347);
nor U8389 (N_8389,N_7224,N_7128);
xnor U8390 (N_8390,N_6293,N_7188);
and U8391 (N_8391,N_6673,N_6510);
xor U8392 (N_8392,N_6359,N_7253);
nand U8393 (N_8393,N_7652,N_7099);
and U8394 (N_8394,N_7258,N_7820);
nor U8395 (N_8395,N_7168,N_7969);
nand U8396 (N_8396,N_7809,N_6115);
nand U8397 (N_8397,N_7940,N_6773);
nor U8398 (N_8398,N_6362,N_7355);
and U8399 (N_8399,N_6466,N_7645);
nand U8400 (N_8400,N_6806,N_6343);
nand U8401 (N_8401,N_7883,N_7204);
or U8402 (N_8402,N_6103,N_7931);
nor U8403 (N_8403,N_6845,N_7305);
nand U8404 (N_8404,N_7221,N_6180);
or U8405 (N_8405,N_6368,N_6563);
or U8406 (N_8406,N_6949,N_6143);
xor U8407 (N_8407,N_6872,N_7777);
nor U8408 (N_8408,N_6488,N_7543);
or U8409 (N_8409,N_6764,N_6641);
xor U8410 (N_8410,N_7988,N_7216);
and U8411 (N_8411,N_6755,N_7183);
nand U8412 (N_8412,N_7306,N_7648);
nor U8413 (N_8413,N_6036,N_6812);
nand U8414 (N_8414,N_7457,N_7360);
and U8415 (N_8415,N_6462,N_7245);
and U8416 (N_8416,N_7942,N_7711);
and U8417 (N_8417,N_6099,N_7394);
nor U8418 (N_8418,N_6001,N_6145);
nor U8419 (N_8419,N_7040,N_6804);
nor U8420 (N_8420,N_7759,N_7792);
nor U8421 (N_8421,N_7363,N_7039);
xnor U8422 (N_8422,N_6006,N_6217);
or U8423 (N_8423,N_6395,N_6648);
nand U8424 (N_8424,N_6270,N_7283);
nand U8425 (N_8425,N_7896,N_6555);
or U8426 (N_8426,N_6014,N_7574);
and U8427 (N_8427,N_7182,N_7022);
nor U8428 (N_8428,N_7800,N_7889);
nand U8429 (N_8429,N_6955,N_7778);
nor U8430 (N_8430,N_7080,N_7869);
and U8431 (N_8431,N_7218,N_6514);
nand U8432 (N_8432,N_7699,N_6611);
nor U8433 (N_8433,N_7257,N_6525);
and U8434 (N_8434,N_7991,N_7117);
nand U8435 (N_8435,N_7084,N_7435);
nand U8436 (N_8436,N_6057,N_6913);
or U8437 (N_8437,N_6134,N_7911);
or U8438 (N_8438,N_6372,N_7106);
xnor U8439 (N_8439,N_6320,N_6373);
nand U8440 (N_8440,N_7556,N_6959);
and U8441 (N_8441,N_6838,N_7688);
nand U8442 (N_8442,N_6319,N_6411);
or U8443 (N_8443,N_7318,N_6465);
or U8444 (N_8444,N_7272,N_7103);
nand U8445 (N_8445,N_6508,N_7721);
nor U8446 (N_8446,N_6044,N_6327);
xnor U8447 (N_8447,N_7285,N_6365);
and U8448 (N_8448,N_6203,N_7004);
nand U8449 (N_8449,N_6526,N_6709);
and U8450 (N_8450,N_6447,N_7270);
nor U8451 (N_8451,N_7123,N_6161);
and U8452 (N_8452,N_7487,N_7818);
xnor U8453 (N_8453,N_7388,N_7749);
or U8454 (N_8454,N_7298,N_6232);
and U8455 (N_8455,N_7674,N_7957);
nor U8456 (N_8456,N_7002,N_7248);
xor U8457 (N_8457,N_6621,N_7446);
and U8458 (N_8458,N_7027,N_7542);
and U8459 (N_8459,N_6586,N_7380);
xor U8460 (N_8460,N_7906,N_7718);
nand U8461 (N_8461,N_6471,N_7553);
and U8462 (N_8462,N_7238,N_7763);
or U8463 (N_8463,N_6356,N_7374);
xor U8464 (N_8464,N_7289,N_7751);
and U8465 (N_8465,N_7698,N_7527);
or U8466 (N_8466,N_7373,N_6191);
or U8467 (N_8467,N_6453,N_7483);
xnor U8468 (N_8468,N_7485,N_6597);
and U8469 (N_8469,N_6307,N_6120);
or U8470 (N_8470,N_6106,N_6264);
and U8471 (N_8471,N_6125,N_6593);
or U8472 (N_8472,N_7088,N_7945);
xor U8473 (N_8473,N_7619,N_7321);
or U8474 (N_8474,N_7052,N_6119);
and U8475 (N_8475,N_6399,N_6989);
nor U8476 (N_8476,N_7138,N_6901);
xor U8477 (N_8477,N_6799,N_6560);
xnor U8478 (N_8478,N_7736,N_7279);
and U8479 (N_8479,N_6055,N_6197);
and U8480 (N_8480,N_6945,N_6026);
or U8481 (N_8481,N_7433,N_6449);
and U8482 (N_8482,N_7308,N_6700);
and U8483 (N_8483,N_6384,N_6429);
nor U8484 (N_8484,N_6122,N_7808);
xnor U8485 (N_8485,N_6075,N_6427);
nor U8486 (N_8486,N_7724,N_7536);
nand U8487 (N_8487,N_7847,N_7838);
or U8488 (N_8488,N_7627,N_7145);
xnor U8489 (N_8489,N_6943,N_7421);
nand U8490 (N_8490,N_7707,N_6000);
nand U8491 (N_8491,N_7251,N_7920);
and U8492 (N_8492,N_7533,N_7059);
or U8493 (N_8493,N_6366,N_6034);
and U8494 (N_8494,N_7968,N_7094);
nor U8495 (N_8495,N_6879,N_6830);
nor U8496 (N_8496,N_7334,N_6314);
nand U8497 (N_8497,N_7431,N_7277);
xnor U8498 (N_8498,N_7157,N_7324);
nand U8499 (N_8499,N_7326,N_6667);
nor U8500 (N_8500,N_6876,N_7055);
and U8501 (N_8501,N_6627,N_6265);
or U8502 (N_8502,N_7819,N_6205);
nor U8503 (N_8503,N_6680,N_6932);
or U8504 (N_8504,N_7015,N_6300);
nand U8505 (N_8505,N_6631,N_7987);
nor U8506 (N_8506,N_6422,N_7781);
nor U8507 (N_8507,N_7119,N_7646);
nand U8508 (N_8508,N_6256,N_7603);
xnor U8509 (N_8509,N_6070,N_7451);
or U8510 (N_8510,N_6608,N_7274);
or U8511 (N_8511,N_6575,N_6515);
and U8512 (N_8512,N_6530,N_7572);
and U8513 (N_8513,N_7694,N_6827);
nand U8514 (N_8514,N_7744,N_6113);
xor U8515 (N_8515,N_6868,N_7395);
and U8516 (N_8516,N_7037,N_7244);
nor U8517 (N_8517,N_7053,N_6782);
nand U8518 (N_8518,N_6928,N_7769);
xnor U8519 (N_8519,N_6665,N_6585);
or U8520 (N_8520,N_7890,N_6243);
xnor U8521 (N_8521,N_7017,N_7085);
nand U8522 (N_8522,N_6795,N_6229);
nand U8523 (N_8523,N_7837,N_7857);
or U8524 (N_8524,N_7464,N_7162);
nor U8525 (N_8525,N_7310,N_6147);
nand U8526 (N_8526,N_7806,N_6997);
nand U8527 (N_8527,N_6283,N_6724);
or U8528 (N_8528,N_6433,N_6707);
and U8529 (N_8529,N_6871,N_7580);
xor U8530 (N_8530,N_6412,N_6802);
and U8531 (N_8531,N_7835,N_7637);
nand U8532 (N_8532,N_7371,N_7678);
xnor U8533 (N_8533,N_6620,N_6619);
nor U8534 (N_8534,N_7528,N_6080);
nand U8535 (N_8535,N_6061,N_7826);
and U8536 (N_8536,N_6286,N_7399);
or U8537 (N_8537,N_7690,N_7613);
or U8538 (N_8538,N_6768,N_7320);
and U8539 (N_8539,N_6780,N_7926);
nor U8540 (N_8540,N_7007,N_6322);
and U8541 (N_8541,N_7501,N_7672);
and U8542 (N_8542,N_6185,N_6934);
xnor U8543 (N_8543,N_7209,N_6018);
xnor U8544 (N_8544,N_6671,N_6121);
xnor U8545 (N_8545,N_6223,N_6132);
nand U8546 (N_8546,N_6096,N_6898);
and U8547 (N_8547,N_6142,N_7922);
and U8548 (N_8548,N_7353,N_6643);
and U8549 (N_8549,N_6763,N_6646);
or U8550 (N_8550,N_6475,N_7615);
nand U8551 (N_8551,N_6669,N_6028);
nor U8552 (N_8552,N_6662,N_7369);
xor U8553 (N_8553,N_7866,N_6834);
xor U8554 (N_8554,N_7952,N_6757);
nand U8555 (N_8555,N_7506,N_6154);
nand U8556 (N_8556,N_6543,N_7898);
nor U8557 (N_8557,N_7676,N_7349);
nand U8558 (N_8558,N_6944,N_7424);
or U8559 (N_8559,N_7173,N_7518);
and U8560 (N_8560,N_6719,N_6977);
nor U8561 (N_8561,N_7861,N_7469);
and U8562 (N_8562,N_6607,N_6954);
or U8563 (N_8563,N_7578,N_6915);
nand U8564 (N_8564,N_6072,N_6246);
and U8565 (N_8565,N_6016,N_6801);
nor U8566 (N_8566,N_7045,N_6336);
nand U8567 (N_8567,N_6201,N_7983);
nor U8568 (N_8568,N_7740,N_7812);
nand U8569 (N_8569,N_7437,N_7243);
or U8570 (N_8570,N_6409,N_6464);
nand U8571 (N_8571,N_7571,N_6128);
nor U8572 (N_8572,N_6357,N_7937);
nor U8573 (N_8573,N_6052,N_7339);
nor U8574 (N_8574,N_6317,N_7292);
and U8575 (N_8575,N_6589,N_6065);
xor U8576 (N_8576,N_6244,N_7247);
xor U8577 (N_8577,N_6511,N_7014);
and U8578 (N_8578,N_6111,N_6777);
and U8579 (N_8579,N_6390,N_6495);
nand U8580 (N_8580,N_6160,N_7842);
nand U8581 (N_8581,N_7018,N_7823);
nand U8582 (N_8582,N_6681,N_6410);
or U8583 (N_8583,N_6546,N_7327);
nand U8584 (N_8584,N_6045,N_6606);
nand U8585 (N_8585,N_6181,N_6255);
xor U8586 (N_8586,N_6573,N_6408);
nand U8587 (N_8587,N_6831,N_6973);
nand U8588 (N_8588,N_7364,N_6815);
nand U8589 (N_8589,N_7576,N_7971);
xor U8590 (N_8590,N_6174,N_6140);
xor U8591 (N_8591,N_6183,N_6279);
and U8592 (N_8592,N_7631,N_7650);
nand U8593 (N_8593,N_6127,N_6927);
xnor U8594 (N_8594,N_7329,N_7579);
or U8595 (N_8595,N_7687,N_6747);
nor U8596 (N_8596,N_6123,N_6361);
xor U8597 (N_8597,N_7267,N_6063);
or U8598 (N_8598,N_6100,N_6482);
xnor U8599 (N_8599,N_6186,N_6213);
nand U8600 (N_8600,N_7817,N_6731);
and U8601 (N_8601,N_7760,N_7591);
and U8602 (N_8602,N_7852,N_6385);
or U8603 (N_8603,N_7745,N_7563);
nand U8604 (N_8604,N_6921,N_7121);
and U8605 (N_8605,N_7512,N_7384);
nor U8606 (N_8606,N_7076,N_6393);
nor U8607 (N_8607,N_7693,N_7375);
or U8608 (N_8608,N_7757,N_6519);
nor U8609 (N_8609,N_7811,N_6592);
nor U8610 (N_8610,N_7848,N_6238);
and U8611 (N_8611,N_7807,N_6787);
and U8612 (N_8612,N_6404,N_7411);
xor U8613 (N_8613,N_6436,N_6506);
nand U8614 (N_8614,N_7322,N_6504);
and U8615 (N_8615,N_6291,N_7500);
nor U8616 (N_8616,N_7044,N_7259);
or U8617 (N_8617,N_7181,N_6479);
or U8618 (N_8618,N_7996,N_6527);
nand U8619 (N_8619,N_6284,N_6767);
or U8620 (N_8620,N_6612,N_6049);
nand U8621 (N_8621,N_6942,N_6963);
nand U8622 (N_8622,N_7161,N_7302);
nor U8623 (N_8623,N_7282,N_6793);
nor U8624 (N_8624,N_7480,N_7127);
nand U8625 (N_8625,N_6138,N_6218);
xnor U8626 (N_8626,N_7043,N_6499);
nor U8627 (N_8627,N_7010,N_6828);
nor U8628 (N_8628,N_6093,N_7673);
or U8629 (N_8629,N_6350,N_7417);
xor U8630 (N_8630,N_6416,N_6492);
xnor U8631 (N_8631,N_6860,N_6078);
and U8632 (N_8632,N_6986,N_7700);
nor U8633 (N_8633,N_7273,N_6770);
nand U8634 (N_8634,N_6446,N_7220);
or U8635 (N_8635,N_6953,N_6148);
nand U8636 (N_8636,N_6533,N_6982);
xor U8637 (N_8637,N_6452,N_6600);
nand U8638 (N_8638,N_7575,N_6720);
and U8639 (N_8639,N_7186,N_6311);
nand U8640 (N_8640,N_6839,N_7166);
or U8641 (N_8641,N_7309,N_7493);
nor U8642 (N_8642,N_6912,N_7816);
and U8643 (N_8643,N_7691,N_7728);
xor U8644 (N_8644,N_6835,N_6658);
xor U8645 (N_8645,N_6292,N_6730);
and U8646 (N_8646,N_6556,N_6081);
nand U8647 (N_8647,N_7936,N_6914);
xor U8648 (N_8648,N_6033,N_7900);
xor U8649 (N_8649,N_6992,N_7829);
nand U8650 (N_8650,N_6863,N_7262);
nor U8651 (N_8651,N_6109,N_7050);
and U8652 (N_8652,N_7381,N_7552);
nand U8653 (N_8653,N_6903,N_6639);
nor U8654 (N_8654,N_7830,N_7206);
xor U8655 (N_8655,N_7523,N_6414);
nor U8656 (N_8656,N_6716,N_7250);
and U8657 (N_8657,N_6976,N_7481);
or U8658 (N_8658,N_7984,N_7478);
and U8659 (N_8659,N_6337,N_6518);
nor U8660 (N_8660,N_7230,N_6363);
nand U8661 (N_8661,N_6771,N_6316);
xnor U8662 (N_8662,N_7056,N_7925);
and U8663 (N_8663,N_7011,N_6969);
or U8664 (N_8664,N_6139,N_7887);
nor U8665 (N_8665,N_7564,N_7420);
or U8666 (N_8666,N_7078,N_6682);
nand U8667 (N_8667,N_7505,N_6599);
or U8668 (N_8668,N_6856,N_6198);
nand U8669 (N_8669,N_7143,N_6214);
nor U8670 (N_8670,N_7459,N_7475);
or U8671 (N_8671,N_7600,N_7796);
and U8672 (N_8672,N_7570,N_6114);
nand U8673 (N_8673,N_7607,N_7065);
and U8674 (N_8674,N_7165,N_6091);
nor U8675 (N_8675,N_7754,N_7705);
xnor U8676 (N_8676,N_7348,N_7509);
xnor U8677 (N_8677,N_7927,N_6616);
nor U8678 (N_8678,N_7917,N_6558);
and U8679 (N_8679,N_7712,N_6811);
and U8680 (N_8680,N_6004,N_7136);
or U8681 (N_8681,N_6022,N_7846);
nand U8682 (N_8682,N_7477,N_7544);
xnor U8683 (N_8683,N_7639,N_7566);
nor U8684 (N_8684,N_6805,N_6030);
nor U8685 (N_8685,N_6630,N_6507);
and U8686 (N_8686,N_6685,N_6501);
and U8687 (N_8687,N_7440,N_7454);
nand U8688 (N_8688,N_7658,N_6654);
nor U8689 (N_8689,N_6524,N_7492);
nor U8690 (N_8690,N_7403,N_6503);
or U8691 (N_8691,N_6675,N_6578);
and U8692 (N_8692,N_7953,N_6129);
nand U8693 (N_8693,N_6825,N_7141);
xor U8694 (N_8694,N_7408,N_6089);
or U8695 (N_8695,N_7685,N_7930);
nand U8696 (N_8696,N_7541,N_6684);
nor U8697 (N_8697,N_7346,N_6383);
xnor U8698 (N_8698,N_6354,N_6231);
and U8699 (N_8699,N_7397,N_6417);
nand U8700 (N_8700,N_7496,N_6206);
and U8701 (N_8701,N_6888,N_6734);
or U8702 (N_8702,N_6776,N_7130);
nor U8703 (N_8703,N_6687,N_6173);
nor U8704 (N_8704,N_6445,N_6800);
nand U8705 (N_8705,N_6318,N_7977);
xor U8706 (N_8706,N_7844,N_7061);
nand U8707 (N_8707,N_7146,N_7255);
nor U8708 (N_8708,N_7791,N_6742);
or U8709 (N_8709,N_6691,N_6535);
nand U8710 (N_8710,N_7932,N_7715);
nand U8711 (N_8711,N_6881,N_6371);
or U8712 (N_8712,N_6097,N_6696);
nand U8713 (N_8713,N_7623,N_6729);
xnor U8714 (N_8714,N_7191,N_6637);
nor U8715 (N_8715,N_7534,N_7235);
xor U8716 (N_8716,N_6919,N_7997);
nand U8717 (N_8717,N_6252,N_7978);
xnor U8718 (N_8718,N_6613,N_7620);
xor U8719 (N_8719,N_6493,N_6401);
and U8720 (N_8720,N_7102,N_6444);
nand U8721 (N_8721,N_7159,N_6002);
and U8722 (N_8722,N_7868,N_6067);
nand U8723 (N_8723,N_7129,N_7064);
xnor U8724 (N_8724,N_6557,N_6200);
nand U8725 (N_8725,N_6467,N_7949);
nand U8726 (N_8726,N_6175,N_7851);
nand U8727 (N_8727,N_7077,N_7311);
nor U8728 (N_8728,N_6126,N_7087);
nand U8729 (N_8729,N_6367,N_6923);
xor U8730 (N_8730,N_6916,N_7521);
or U8731 (N_8731,N_7872,N_7222);
xnor U8732 (N_8732,N_7609,N_7429);
or U8733 (N_8733,N_6554,N_7537);
nor U8734 (N_8734,N_6867,N_6714);
and U8735 (N_8735,N_6168,N_6153);
nand U8736 (N_8736,N_7197,N_7202);
xnor U8737 (N_8737,N_6008,N_7332);
nand U8738 (N_8738,N_7567,N_6068);
or U8739 (N_8739,N_7118,N_6215);
nand U8740 (N_8740,N_6146,N_6240);
or U8741 (N_8741,N_7888,N_6069);
xor U8742 (N_8742,N_6626,N_7170);
nand U8743 (N_8743,N_6739,N_7695);
xnor U8744 (N_8744,N_6117,N_6817);
xor U8745 (N_8745,N_6321,N_6387);
or U8746 (N_8746,N_6721,N_6060);
and U8747 (N_8747,N_7133,N_7827);
nor U8748 (N_8748,N_7714,N_7046);
nand U8749 (N_8749,N_7093,N_7904);
nor U8750 (N_8750,N_6164,N_7470);
nand U8751 (N_8751,N_7468,N_7236);
or U8752 (N_8752,N_7325,N_6590);
and U8753 (N_8753,N_6664,N_6077);
and U8754 (N_8754,N_6657,N_6577);
and U8755 (N_8755,N_6421,N_7497);
and U8756 (N_8756,N_6167,N_7153);
nand U8757 (N_8757,N_7489,N_7362);
and U8758 (N_8758,N_7461,N_6455);
xnor U8759 (N_8759,N_7979,N_7404);
nand U8760 (N_8760,N_6403,N_7960);
or U8761 (N_8761,N_6323,N_7148);
nand U8762 (N_8762,N_6048,N_7203);
or U8763 (N_8763,N_7626,N_7719);
and U8764 (N_8764,N_6737,N_7208);
nand U8765 (N_8765,N_6135,N_7799);
nor U8766 (N_8766,N_7293,N_6926);
nor U8767 (N_8767,N_6791,N_7944);
xnor U8768 (N_8768,N_7840,N_6329);
xnor U8769 (N_8769,N_7696,N_6378);
xor U8770 (N_8770,N_7406,N_7109);
xnor U8771 (N_8771,N_7532,N_6723);
or U8772 (N_8772,N_7538,N_7175);
and U8773 (N_8773,N_7730,N_7879);
xor U8774 (N_8774,N_7511,N_7107);
nand U8775 (N_8775,N_6581,N_7498);
nand U8776 (N_8776,N_6971,N_7092);
and U8777 (N_8777,N_6635,N_6784);
nand U8778 (N_8778,N_7897,N_6076);
and U8779 (N_8779,N_6224,N_7449);
nor U8780 (N_8780,N_6893,N_6902);
or U8781 (N_8781,N_7467,N_6312);
or U8782 (N_8782,N_6907,N_6190);
nand U8783 (N_8783,N_6522,N_6981);
nor U8784 (N_8784,N_7636,N_7825);
nor U8785 (N_8785,N_7908,N_7444);
nor U8786 (N_8786,N_6486,N_6210);
or U8787 (N_8787,N_7771,N_6929);
or U8788 (N_8788,N_6956,N_6505);
nor U8789 (N_8789,N_6498,N_7747);
nand U8790 (N_8790,N_7434,N_6423);
xnor U8791 (N_8791,N_6746,N_6947);
and U8792 (N_8792,N_7768,N_7551);
and U8793 (N_8793,N_6745,N_7679);
xnor U8794 (N_8794,N_7368,N_6227);
and U8795 (N_8795,N_7524,N_7597);
and U8796 (N_8796,N_6458,N_7520);
xnor U8797 (N_8797,N_6836,N_7214);
nor U8798 (N_8798,N_7242,N_7428);
nand U8799 (N_8799,N_6931,N_7295);
xor U8800 (N_8800,N_6559,N_7445);
nor U8801 (N_8801,N_6640,N_6897);
xor U8802 (N_8802,N_6679,N_6241);
and U8803 (N_8803,N_7313,N_7025);
nor U8804 (N_8804,N_7881,N_6497);
and U8805 (N_8805,N_6690,N_7268);
nor U8806 (N_8806,N_7072,N_6829);
or U8807 (N_8807,N_7139,N_6086);
nand U8808 (N_8808,N_7589,N_7752);
nor U8809 (N_8809,N_6918,N_6472);
or U8810 (N_8810,N_7584,N_6381);
nand U8811 (N_8811,N_6207,N_6859);
nor U8812 (N_8812,N_6946,N_6760);
xnor U8813 (N_8813,N_6591,N_6202);
xor U8814 (N_8814,N_6426,N_6221);
or U8815 (N_8815,N_7034,N_7398);
xnor U8816 (N_8816,N_7955,N_7914);
nand U8817 (N_8817,N_6087,N_6184);
nand U8818 (N_8818,N_7709,N_6382);
and U8819 (N_8819,N_7196,N_6978);
nand U8820 (N_8820,N_6290,N_7790);
nor U8821 (N_8821,N_7972,N_7303);
xor U8822 (N_8822,N_6424,N_7116);
xor U8823 (N_8823,N_6483,N_6968);
nor U8824 (N_8824,N_6833,N_7001);
and U8825 (N_8825,N_7713,N_7351);
or U8826 (N_8826,N_7387,N_7649);
and U8827 (N_8827,N_7164,N_7280);
xnor U8828 (N_8828,N_6335,N_6261);
and U8829 (N_8829,N_7756,N_7192);
nor U8830 (N_8830,N_6435,N_7047);
nand U8831 (N_8831,N_6131,N_7490);
nand U8832 (N_8832,N_7357,N_6610);
or U8833 (N_8833,N_7333,N_7089);
or U8834 (N_8834,N_7060,N_6263);
nand U8835 (N_8835,N_6810,N_7023);
nor U8836 (N_8836,N_7131,N_6552);
xor U8837 (N_8837,N_6889,N_7344);
nor U8838 (N_8838,N_7966,N_6743);
nor U8839 (N_8839,N_7616,N_6677);
nand U8840 (N_8840,N_7430,N_7559);
nor U8841 (N_8841,N_6728,N_6789);
nor U8842 (N_8842,N_6722,N_7263);
nor U8843 (N_8843,N_7608,N_6678);
or U8844 (N_8844,N_7743,N_7885);
or U8845 (N_8845,N_7312,N_7425);
xnor U8846 (N_8846,N_6532,N_7337);
xnor U8847 (N_8847,N_6605,N_7132);
or U8848 (N_8848,N_7113,N_7323);
and U8849 (N_8849,N_6009,N_6702);
xor U8850 (N_8850,N_6844,N_6520);
nor U8851 (N_8851,N_6629,N_6011);
and U8852 (N_8852,N_7179,N_6235);
xor U8853 (N_8853,N_6259,N_6766);
or U8854 (N_8854,N_6490,N_7341);
nor U8855 (N_8855,N_7416,N_7441);
xnor U8856 (N_8856,N_7086,N_6545);
nand U8857 (N_8857,N_6647,N_7287);
nor U8858 (N_8858,N_7614,N_6509);
nand U8859 (N_8859,N_7951,N_6105);
and U8860 (N_8860,N_7656,N_6487);
xor U8861 (N_8861,N_7402,N_6580);
xor U8862 (N_8862,N_7793,N_7973);
nand U8863 (N_8863,N_6124,N_7993);
xnor U8864 (N_8864,N_6751,N_6656);
or U8865 (N_8865,N_6858,N_7054);
xnor U8866 (N_8866,N_6803,N_7462);
or U8867 (N_8867,N_7423,N_6165);
and U8868 (N_8868,N_6112,N_7396);
and U8869 (N_8869,N_6705,N_7359);
or U8870 (N_8870,N_6674,N_7994);
nor U8871 (N_8871,N_7948,N_6951);
and U8872 (N_8872,N_7555,N_7525);
nor U8873 (N_8873,N_7726,N_6566);
and U8874 (N_8874,N_6561,N_6788);
and U8875 (N_8875,N_7115,N_6349);
nor U8876 (N_8876,N_7135,N_6088);
xor U8877 (N_8877,N_7780,N_7187);
xnor U8878 (N_8878,N_6375,N_7668);
or U8879 (N_8879,N_7038,N_7101);
nand U8880 (N_8880,N_7867,N_6434);
nand U8881 (N_8881,N_6274,N_6692);
or U8882 (N_8882,N_7995,N_7634);
nand U8883 (N_8883,N_6814,N_6470);
nor U8884 (N_8884,N_6182,N_6056);
nor U8885 (N_8885,N_7588,N_6459);
nand U8886 (N_8886,N_7366,N_6277);
nor U8887 (N_8887,N_7941,N_6790);
nand U8888 (N_8888,N_6236,N_6663);
nor U8889 (N_8889,N_7223,N_6999);
or U8890 (N_8890,N_6340,N_7057);
xnor U8891 (N_8891,N_6017,N_6686);
or U8892 (N_8892,N_6053,N_6358);
xnor U8893 (N_8893,N_7304,N_7494);
xor U8894 (N_8894,N_7689,N_7907);
nor U8895 (N_8895,N_7638,N_7954);
nand U8896 (N_8896,N_6890,N_7860);
nand U8897 (N_8897,N_7069,N_7935);
xnor U8898 (N_8898,N_6425,N_7432);
and U8899 (N_8899,N_6713,N_6905);
nor U8900 (N_8900,N_6276,N_7794);
and U8901 (N_8901,N_7021,N_7704);
nor U8902 (N_8902,N_6996,N_6516);
xnor U8903 (N_8903,N_7599,N_7670);
nor U8904 (N_8904,N_7737,N_6303);
nand U8905 (N_8905,N_7361,N_6196);
and U8906 (N_8906,N_6758,N_7319);
nor U8907 (N_8907,N_6250,N_6797);
or U8908 (N_8908,N_7814,N_7377);
xor U8909 (N_8909,N_7843,N_7683);
nor U8910 (N_8910,N_7419,N_7026);
or U8911 (N_8911,N_7379,N_6668);
nor U8912 (N_8912,N_6885,N_6082);
or U8913 (N_8913,N_7508,N_7916);
and U8914 (N_8914,N_6937,N_7062);
nor U8915 (N_8915,N_7894,N_7447);
and U8916 (N_8916,N_6031,N_6622);
nor U8917 (N_8917,N_7484,N_7641);
xnor U8918 (N_8918,N_6880,N_7151);
nor U8919 (N_8919,N_6821,N_7482);
and U8920 (N_8920,N_6523,N_6798);
or U8921 (N_8921,N_7260,N_6478);
xnor U8922 (N_8922,N_6568,N_6152);
nor U8923 (N_8923,N_7231,N_6661);
and U8924 (N_8924,N_6260,N_6457);
nor U8925 (N_8925,N_7758,N_7042);
nand U8926 (N_8926,N_7617,N_7178);
and U8927 (N_8927,N_7226,N_6296);
nand U8928 (N_8928,N_7199,N_6979);
or U8929 (N_8929,N_6699,N_6348);
nor U8930 (N_8930,N_7938,N_6047);
nand U8931 (N_8931,N_7647,N_6418);
nand U8932 (N_8932,N_6090,N_7048);
and U8933 (N_8933,N_6370,N_7315);
nor U8934 (N_8934,N_6007,N_6940);
and U8935 (N_8935,N_7956,N_6576);
xor U8936 (N_8936,N_6439,N_6693);
nor U8937 (N_8937,N_6570,N_7125);
nor U8938 (N_8938,N_7352,N_6572);
and U8939 (N_8939,N_7227,N_6851);
xnor U8940 (N_8940,N_6877,N_7667);
and U8941 (N_8941,N_7016,N_7122);
nor U8942 (N_8942,N_6400,N_6003);
nand U8943 (N_8943,N_7005,N_6886);
xnor U8944 (N_8944,N_7297,N_6849);
or U8945 (N_8945,N_7895,N_6170);
and U8946 (N_8946,N_6245,N_7330);
or U8947 (N_8947,N_6477,N_7635);
nand U8948 (N_8948,N_7934,N_7382);
nor U8949 (N_8949,N_6430,N_7020);
xor U8950 (N_8950,N_7516,N_6587);
or U8951 (N_8951,N_6171,N_6178);
nand U8952 (N_8952,N_6653,N_6315);
xor U8953 (N_8953,N_6355,N_7172);
xnor U8954 (N_8954,N_6313,N_6847);
nand U8955 (N_8955,N_6301,N_7739);
xnor U8956 (N_8956,N_6636,N_7422);
xor U8957 (N_8957,N_6225,N_7557);
and U8958 (N_8958,N_7797,N_7239);
or U8959 (N_8959,N_7342,N_6133);
or U8960 (N_8960,N_6451,N_6741);
or U8961 (N_8961,N_7549,N_7577);
nand U8962 (N_8962,N_6407,N_7356);
and U8963 (N_8963,N_6710,N_7573);
nor U8964 (N_8964,N_7766,N_6842);
xor U8965 (N_8965,N_6156,N_7269);
and U8966 (N_8966,N_6195,N_7921);
nand U8967 (N_8967,N_6822,N_6415);
and U8968 (N_8968,N_6268,N_7515);
and U8969 (N_8969,N_7195,N_7473);
nor U8970 (N_8970,N_7587,N_7031);
and U8971 (N_8971,N_6029,N_6869);
xnor U8972 (N_8972,N_7632,N_7531);
xnor U8973 (N_8973,N_7939,N_6460);
or U8974 (N_8974,N_6299,N_7593);
or U8975 (N_8975,N_6285,N_6900);
nor U8976 (N_8976,N_7828,N_6813);
or U8977 (N_8977,N_6701,N_7892);
and U8978 (N_8978,N_7974,N_7787);
xor U8979 (N_8979,N_7460,N_6911);
nor U8980 (N_8980,N_7863,N_7606);
nand U8981 (N_8981,N_7150,N_7912);
nand U8982 (N_8982,N_6910,N_6494);
xor U8983 (N_8983,N_6628,N_6005);
or U8984 (N_8984,N_6617,N_6623);
or U8985 (N_8985,N_7720,N_7663);
and U8986 (N_8986,N_6596,N_6258);
and U8987 (N_8987,N_7729,N_7833);
nand U8988 (N_8988,N_6484,N_6855);
or U8989 (N_8989,N_6994,N_6588);
and U8990 (N_8990,N_6521,N_7998);
xnor U8991 (N_8991,N_7654,N_6972);
nor U8992 (N_8992,N_7155,N_6380);
and U8993 (N_8993,N_7703,N_6150);
nor U8994 (N_8994,N_6984,N_6010);
nand U8995 (N_8995,N_6759,N_7455);
nand U8996 (N_8996,N_6652,N_7003);
nand U8997 (N_8997,N_6785,N_6454);
and U8998 (N_8998,N_6601,N_7063);
xor U8999 (N_8999,N_7499,N_7677);
xnor U9000 (N_9000,N_6915,N_6643);
and U9001 (N_9001,N_6098,N_6212);
nand U9002 (N_9002,N_7204,N_6678);
and U9003 (N_9003,N_6802,N_7415);
nand U9004 (N_9004,N_7274,N_6059);
nand U9005 (N_9005,N_6603,N_7201);
xor U9006 (N_9006,N_7144,N_7917);
and U9007 (N_9007,N_6960,N_7924);
xnor U9008 (N_9008,N_7138,N_7831);
and U9009 (N_9009,N_7954,N_6702);
or U9010 (N_9010,N_6199,N_7947);
nor U9011 (N_9011,N_6268,N_6230);
nor U9012 (N_9012,N_6247,N_6843);
and U9013 (N_9013,N_6412,N_6908);
nand U9014 (N_9014,N_6567,N_7558);
nor U9015 (N_9015,N_7585,N_6832);
xor U9016 (N_9016,N_6493,N_6680);
nand U9017 (N_9017,N_6716,N_6576);
and U9018 (N_9018,N_6653,N_6901);
nand U9019 (N_9019,N_6199,N_6160);
nor U9020 (N_9020,N_6201,N_6924);
nor U9021 (N_9021,N_7211,N_7054);
xor U9022 (N_9022,N_6689,N_6756);
nor U9023 (N_9023,N_6540,N_6780);
nor U9024 (N_9024,N_6030,N_7481);
xor U9025 (N_9025,N_7721,N_6783);
nor U9026 (N_9026,N_7529,N_7438);
xnor U9027 (N_9027,N_6605,N_6944);
nor U9028 (N_9028,N_6555,N_7495);
nand U9029 (N_9029,N_6486,N_7058);
nor U9030 (N_9030,N_6406,N_6641);
or U9031 (N_9031,N_6357,N_7763);
and U9032 (N_9032,N_7742,N_7971);
and U9033 (N_9033,N_7750,N_7299);
xnor U9034 (N_9034,N_7511,N_6617);
nor U9035 (N_9035,N_6877,N_6431);
nand U9036 (N_9036,N_7857,N_6062);
or U9037 (N_9037,N_7671,N_6355);
and U9038 (N_9038,N_6105,N_7769);
or U9039 (N_9039,N_7190,N_6169);
and U9040 (N_9040,N_7150,N_6955);
nand U9041 (N_9041,N_7052,N_6218);
or U9042 (N_9042,N_6357,N_6969);
nand U9043 (N_9043,N_6487,N_7766);
or U9044 (N_9044,N_6695,N_6911);
xnor U9045 (N_9045,N_6883,N_7001);
nor U9046 (N_9046,N_7542,N_6017);
nor U9047 (N_9047,N_6913,N_6599);
and U9048 (N_9048,N_6723,N_7150);
xnor U9049 (N_9049,N_7307,N_6265);
and U9050 (N_9050,N_7009,N_7699);
nand U9051 (N_9051,N_6138,N_6061);
and U9052 (N_9052,N_6508,N_7399);
nand U9053 (N_9053,N_6545,N_7458);
and U9054 (N_9054,N_6168,N_6450);
xnor U9055 (N_9055,N_6700,N_6362);
nand U9056 (N_9056,N_7481,N_6928);
nor U9057 (N_9057,N_7867,N_6908);
nor U9058 (N_9058,N_6021,N_6251);
nand U9059 (N_9059,N_6996,N_6186);
nand U9060 (N_9060,N_6050,N_7180);
or U9061 (N_9061,N_6738,N_6735);
nor U9062 (N_9062,N_7753,N_6096);
nand U9063 (N_9063,N_6696,N_7967);
xnor U9064 (N_9064,N_6559,N_7797);
nand U9065 (N_9065,N_7918,N_7245);
xnor U9066 (N_9066,N_6615,N_7283);
and U9067 (N_9067,N_6596,N_7083);
nand U9068 (N_9068,N_6549,N_6522);
and U9069 (N_9069,N_6643,N_7721);
and U9070 (N_9070,N_6571,N_6882);
and U9071 (N_9071,N_7205,N_6704);
and U9072 (N_9072,N_6659,N_6758);
nand U9073 (N_9073,N_7622,N_7906);
nand U9074 (N_9074,N_6079,N_6305);
or U9075 (N_9075,N_7974,N_7005);
nand U9076 (N_9076,N_7899,N_6213);
and U9077 (N_9077,N_7508,N_7767);
xnor U9078 (N_9078,N_7189,N_7234);
nor U9079 (N_9079,N_6314,N_6736);
and U9080 (N_9080,N_6303,N_6293);
nand U9081 (N_9081,N_6370,N_6253);
nor U9082 (N_9082,N_6251,N_6246);
and U9083 (N_9083,N_7820,N_7014);
xor U9084 (N_9084,N_6944,N_7705);
nor U9085 (N_9085,N_7998,N_7211);
nand U9086 (N_9086,N_6414,N_6354);
xor U9087 (N_9087,N_7183,N_6647);
and U9088 (N_9088,N_7616,N_7638);
nor U9089 (N_9089,N_6213,N_6755);
nor U9090 (N_9090,N_6618,N_7256);
nand U9091 (N_9091,N_7925,N_7673);
xor U9092 (N_9092,N_6266,N_6791);
nor U9093 (N_9093,N_7024,N_6820);
nand U9094 (N_9094,N_6791,N_7243);
xor U9095 (N_9095,N_7885,N_6451);
nand U9096 (N_9096,N_6275,N_6011);
and U9097 (N_9097,N_7606,N_6768);
or U9098 (N_9098,N_6137,N_7412);
xnor U9099 (N_9099,N_7922,N_7947);
and U9100 (N_9100,N_6765,N_6662);
or U9101 (N_9101,N_7376,N_7414);
nor U9102 (N_9102,N_7281,N_7920);
nand U9103 (N_9103,N_6314,N_6503);
nor U9104 (N_9104,N_6945,N_7886);
xnor U9105 (N_9105,N_7210,N_7256);
nor U9106 (N_9106,N_6649,N_6523);
and U9107 (N_9107,N_7438,N_6736);
or U9108 (N_9108,N_6201,N_6709);
nor U9109 (N_9109,N_6340,N_6722);
and U9110 (N_9110,N_7302,N_6041);
xnor U9111 (N_9111,N_6974,N_7733);
and U9112 (N_9112,N_7213,N_6921);
or U9113 (N_9113,N_6365,N_7654);
nand U9114 (N_9114,N_7343,N_6676);
xnor U9115 (N_9115,N_7548,N_7631);
xnor U9116 (N_9116,N_6849,N_7619);
or U9117 (N_9117,N_6109,N_6668);
and U9118 (N_9118,N_7565,N_6331);
and U9119 (N_9119,N_6789,N_7947);
nand U9120 (N_9120,N_7797,N_7837);
and U9121 (N_9121,N_6833,N_7821);
nor U9122 (N_9122,N_6853,N_6784);
nand U9123 (N_9123,N_7372,N_7057);
nand U9124 (N_9124,N_6954,N_7781);
xnor U9125 (N_9125,N_7389,N_6942);
and U9126 (N_9126,N_6546,N_6192);
nor U9127 (N_9127,N_7626,N_6649);
and U9128 (N_9128,N_7290,N_6322);
xor U9129 (N_9129,N_6282,N_7336);
or U9130 (N_9130,N_6429,N_7254);
nand U9131 (N_9131,N_6293,N_7262);
nor U9132 (N_9132,N_6996,N_6873);
nor U9133 (N_9133,N_7531,N_7913);
and U9134 (N_9134,N_7283,N_7766);
or U9135 (N_9135,N_6860,N_7706);
nor U9136 (N_9136,N_7714,N_7971);
and U9137 (N_9137,N_7880,N_6284);
nor U9138 (N_9138,N_6262,N_7008);
and U9139 (N_9139,N_7780,N_6963);
and U9140 (N_9140,N_6681,N_7687);
or U9141 (N_9141,N_7143,N_6062);
nand U9142 (N_9142,N_7079,N_6846);
and U9143 (N_9143,N_6351,N_7626);
or U9144 (N_9144,N_6116,N_7363);
xor U9145 (N_9145,N_6045,N_6122);
and U9146 (N_9146,N_6719,N_7544);
xnor U9147 (N_9147,N_7057,N_7605);
nand U9148 (N_9148,N_7767,N_7251);
nand U9149 (N_9149,N_7635,N_6084);
nand U9150 (N_9150,N_7397,N_7430);
xor U9151 (N_9151,N_6713,N_6185);
xor U9152 (N_9152,N_7176,N_6330);
nor U9153 (N_9153,N_6260,N_7822);
nor U9154 (N_9154,N_6898,N_6785);
and U9155 (N_9155,N_7573,N_6890);
or U9156 (N_9156,N_6693,N_7212);
nand U9157 (N_9157,N_7301,N_6677);
xnor U9158 (N_9158,N_6274,N_7361);
or U9159 (N_9159,N_6978,N_7915);
xnor U9160 (N_9160,N_7946,N_7024);
or U9161 (N_9161,N_6465,N_7427);
and U9162 (N_9162,N_7596,N_6564);
and U9163 (N_9163,N_7543,N_6070);
nor U9164 (N_9164,N_7717,N_6029);
xor U9165 (N_9165,N_6805,N_6048);
nor U9166 (N_9166,N_6873,N_6106);
nor U9167 (N_9167,N_6830,N_7778);
xor U9168 (N_9168,N_7632,N_7405);
and U9169 (N_9169,N_7917,N_7537);
and U9170 (N_9170,N_6902,N_6374);
xnor U9171 (N_9171,N_6014,N_7579);
nand U9172 (N_9172,N_6643,N_7717);
nor U9173 (N_9173,N_7378,N_6304);
xnor U9174 (N_9174,N_7038,N_7516);
nor U9175 (N_9175,N_6538,N_7639);
xnor U9176 (N_9176,N_7455,N_6712);
nor U9177 (N_9177,N_7771,N_7218);
or U9178 (N_9178,N_7970,N_6283);
nor U9179 (N_9179,N_7583,N_7360);
nor U9180 (N_9180,N_6081,N_7947);
and U9181 (N_9181,N_6583,N_7752);
and U9182 (N_9182,N_7034,N_7596);
and U9183 (N_9183,N_6904,N_7356);
and U9184 (N_9184,N_6742,N_7703);
and U9185 (N_9185,N_7119,N_6254);
and U9186 (N_9186,N_7343,N_6222);
or U9187 (N_9187,N_7858,N_7651);
and U9188 (N_9188,N_6012,N_6797);
nand U9189 (N_9189,N_6167,N_7699);
xor U9190 (N_9190,N_7869,N_7972);
xnor U9191 (N_9191,N_7859,N_7233);
xnor U9192 (N_9192,N_6840,N_6707);
nor U9193 (N_9193,N_6802,N_7927);
and U9194 (N_9194,N_7707,N_6465);
nor U9195 (N_9195,N_7067,N_7182);
or U9196 (N_9196,N_7249,N_7652);
nand U9197 (N_9197,N_6087,N_7674);
and U9198 (N_9198,N_6330,N_7018);
nor U9199 (N_9199,N_7485,N_6982);
nor U9200 (N_9200,N_7681,N_6407);
nor U9201 (N_9201,N_6428,N_6871);
xnor U9202 (N_9202,N_7855,N_7253);
or U9203 (N_9203,N_6887,N_6634);
nand U9204 (N_9204,N_7657,N_6438);
nand U9205 (N_9205,N_6541,N_6108);
or U9206 (N_9206,N_7627,N_7849);
nand U9207 (N_9207,N_7576,N_6888);
nor U9208 (N_9208,N_7492,N_7501);
or U9209 (N_9209,N_6127,N_7499);
xnor U9210 (N_9210,N_7342,N_6944);
or U9211 (N_9211,N_6431,N_7265);
or U9212 (N_9212,N_7315,N_6418);
xor U9213 (N_9213,N_6971,N_6829);
or U9214 (N_9214,N_7310,N_6831);
and U9215 (N_9215,N_7895,N_7578);
or U9216 (N_9216,N_7205,N_7488);
nand U9217 (N_9217,N_6846,N_6884);
or U9218 (N_9218,N_7754,N_7690);
xnor U9219 (N_9219,N_7146,N_6682);
xor U9220 (N_9220,N_6921,N_7044);
nor U9221 (N_9221,N_7174,N_7117);
or U9222 (N_9222,N_6074,N_6901);
and U9223 (N_9223,N_6399,N_6201);
nor U9224 (N_9224,N_7408,N_6662);
xor U9225 (N_9225,N_6032,N_6171);
and U9226 (N_9226,N_6965,N_7888);
xor U9227 (N_9227,N_6782,N_6308);
xor U9228 (N_9228,N_7052,N_7487);
xor U9229 (N_9229,N_7877,N_7084);
nor U9230 (N_9230,N_7804,N_6219);
or U9231 (N_9231,N_7851,N_6736);
and U9232 (N_9232,N_6601,N_7543);
and U9233 (N_9233,N_6355,N_6788);
and U9234 (N_9234,N_7233,N_6290);
and U9235 (N_9235,N_7545,N_7305);
or U9236 (N_9236,N_6541,N_6311);
nand U9237 (N_9237,N_7244,N_6596);
xnor U9238 (N_9238,N_6743,N_6819);
xnor U9239 (N_9239,N_6741,N_7219);
and U9240 (N_9240,N_6031,N_7106);
nor U9241 (N_9241,N_6938,N_7249);
nor U9242 (N_9242,N_7201,N_6942);
xnor U9243 (N_9243,N_7232,N_6215);
nand U9244 (N_9244,N_6701,N_7043);
nand U9245 (N_9245,N_6246,N_6436);
and U9246 (N_9246,N_7108,N_7309);
nand U9247 (N_9247,N_6708,N_6749);
and U9248 (N_9248,N_6574,N_7678);
and U9249 (N_9249,N_7584,N_6949);
nor U9250 (N_9250,N_6631,N_6843);
and U9251 (N_9251,N_6523,N_7172);
nor U9252 (N_9252,N_6930,N_6286);
nor U9253 (N_9253,N_6191,N_7172);
xnor U9254 (N_9254,N_6258,N_6744);
nand U9255 (N_9255,N_7777,N_6034);
xor U9256 (N_9256,N_7310,N_7519);
nor U9257 (N_9257,N_7534,N_6042);
nor U9258 (N_9258,N_6676,N_6447);
nand U9259 (N_9259,N_6655,N_7380);
nand U9260 (N_9260,N_6269,N_7826);
and U9261 (N_9261,N_7550,N_7143);
and U9262 (N_9262,N_7507,N_7714);
and U9263 (N_9263,N_7856,N_6770);
xnor U9264 (N_9264,N_7277,N_6220);
xnor U9265 (N_9265,N_6824,N_6990);
or U9266 (N_9266,N_7761,N_7169);
and U9267 (N_9267,N_6152,N_7429);
and U9268 (N_9268,N_7224,N_6433);
xor U9269 (N_9269,N_7180,N_7522);
nand U9270 (N_9270,N_6102,N_7617);
nand U9271 (N_9271,N_7506,N_6585);
nand U9272 (N_9272,N_7109,N_7395);
or U9273 (N_9273,N_7514,N_7069);
or U9274 (N_9274,N_7895,N_6021);
xor U9275 (N_9275,N_7295,N_7506);
nand U9276 (N_9276,N_7076,N_7634);
or U9277 (N_9277,N_7704,N_6416);
xnor U9278 (N_9278,N_6184,N_6595);
nand U9279 (N_9279,N_6123,N_7104);
xnor U9280 (N_9280,N_7840,N_6227);
and U9281 (N_9281,N_6728,N_7511);
or U9282 (N_9282,N_6377,N_7578);
nor U9283 (N_9283,N_6509,N_7893);
or U9284 (N_9284,N_7851,N_6798);
nand U9285 (N_9285,N_7737,N_6275);
xnor U9286 (N_9286,N_6266,N_6363);
xnor U9287 (N_9287,N_6888,N_7191);
and U9288 (N_9288,N_7469,N_7472);
nand U9289 (N_9289,N_6217,N_7248);
xor U9290 (N_9290,N_6066,N_7579);
and U9291 (N_9291,N_6485,N_6055);
nor U9292 (N_9292,N_7902,N_7268);
xor U9293 (N_9293,N_6785,N_6954);
nand U9294 (N_9294,N_7211,N_7606);
nor U9295 (N_9295,N_7730,N_7045);
xor U9296 (N_9296,N_7785,N_7693);
or U9297 (N_9297,N_6912,N_6968);
and U9298 (N_9298,N_7947,N_6145);
xnor U9299 (N_9299,N_7532,N_7996);
or U9300 (N_9300,N_7312,N_7867);
and U9301 (N_9301,N_6260,N_7641);
and U9302 (N_9302,N_7992,N_6007);
nor U9303 (N_9303,N_6962,N_7556);
and U9304 (N_9304,N_7856,N_7776);
and U9305 (N_9305,N_6138,N_6001);
nor U9306 (N_9306,N_6835,N_6151);
nor U9307 (N_9307,N_6192,N_7789);
nor U9308 (N_9308,N_6746,N_7903);
nor U9309 (N_9309,N_7280,N_6189);
or U9310 (N_9310,N_6851,N_6669);
and U9311 (N_9311,N_7687,N_7682);
and U9312 (N_9312,N_7786,N_6139);
nor U9313 (N_9313,N_7583,N_7833);
xnor U9314 (N_9314,N_6695,N_7634);
or U9315 (N_9315,N_6979,N_6777);
or U9316 (N_9316,N_6885,N_6557);
or U9317 (N_9317,N_6262,N_6049);
or U9318 (N_9318,N_6264,N_7797);
nand U9319 (N_9319,N_7042,N_7517);
nor U9320 (N_9320,N_6842,N_6881);
or U9321 (N_9321,N_7161,N_7522);
nor U9322 (N_9322,N_7375,N_7756);
and U9323 (N_9323,N_7503,N_7403);
nor U9324 (N_9324,N_6027,N_6394);
nor U9325 (N_9325,N_6294,N_6691);
nand U9326 (N_9326,N_6784,N_7186);
or U9327 (N_9327,N_6949,N_6635);
nor U9328 (N_9328,N_7875,N_7787);
nand U9329 (N_9329,N_7978,N_6377);
xor U9330 (N_9330,N_7815,N_6469);
xnor U9331 (N_9331,N_6223,N_7347);
or U9332 (N_9332,N_6751,N_6457);
nor U9333 (N_9333,N_6631,N_6363);
or U9334 (N_9334,N_6100,N_6636);
xor U9335 (N_9335,N_7937,N_7711);
xnor U9336 (N_9336,N_7670,N_6209);
and U9337 (N_9337,N_7418,N_7316);
and U9338 (N_9338,N_6642,N_7487);
and U9339 (N_9339,N_6091,N_7321);
or U9340 (N_9340,N_6442,N_7044);
xor U9341 (N_9341,N_7044,N_6940);
nand U9342 (N_9342,N_6661,N_6081);
nor U9343 (N_9343,N_7494,N_7533);
nor U9344 (N_9344,N_7657,N_6207);
nor U9345 (N_9345,N_7703,N_7325);
nor U9346 (N_9346,N_6995,N_6762);
or U9347 (N_9347,N_6952,N_7047);
and U9348 (N_9348,N_6125,N_6641);
and U9349 (N_9349,N_7436,N_6155);
and U9350 (N_9350,N_7774,N_7328);
nor U9351 (N_9351,N_7796,N_6679);
nor U9352 (N_9352,N_7585,N_6197);
nand U9353 (N_9353,N_6593,N_7007);
nand U9354 (N_9354,N_6551,N_6579);
nor U9355 (N_9355,N_6920,N_7965);
or U9356 (N_9356,N_7399,N_7180);
nor U9357 (N_9357,N_7889,N_6496);
nand U9358 (N_9358,N_7429,N_7593);
nand U9359 (N_9359,N_7855,N_6469);
nor U9360 (N_9360,N_6573,N_7281);
nor U9361 (N_9361,N_6839,N_6286);
nand U9362 (N_9362,N_6025,N_6894);
nand U9363 (N_9363,N_7795,N_6414);
nand U9364 (N_9364,N_6787,N_6747);
or U9365 (N_9365,N_6782,N_6891);
nand U9366 (N_9366,N_7949,N_6391);
and U9367 (N_9367,N_6972,N_7125);
and U9368 (N_9368,N_7967,N_7045);
or U9369 (N_9369,N_7673,N_7626);
nand U9370 (N_9370,N_7800,N_7715);
nand U9371 (N_9371,N_7460,N_6464);
xor U9372 (N_9372,N_6198,N_7135);
xnor U9373 (N_9373,N_6893,N_6705);
xnor U9374 (N_9374,N_6649,N_7195);
nand U9375 (N_9375,N_6531,N_6495);
or U9376 (N_9376,N_6825,N_7477);
nand U9377 (N_9377,N_7958,N_7667);
nor U9378 (N_9378,N_6395,N_7512);
xor U9379 (N_9379,N_7607,N_6389);
or U9380 (N_9380,N_6677,N_6981);
nand U9381 (N_9381,N_6650,N_6748);
nor U9382 (N_9382,N_6705,N_7755);
and U9383 (N_9383,N_7305,N_7497);
nand U9384 (N_9384,N_7328,N_7444);
or U9385 (N_9385,N_6637,N_6964);
nor U9386 (N_9386,N_7984,N_6537);
nand U9387 (N_9387,N_7025,N_7506);
nor U9388 (N_9388,N_6259,N_6533);
or U9389 (N_9389,N_6909,N_7205);
nor U9390 (N_9390,N_6118,N_7591);
nand U9391 (N_9391,N_6201,N_6215);
nor U9392 (N_9392,N_6871,N_6811);
nand U9393 (N_9393,N_7853,N_6522);
xor U9394 (N_9394,N_6708,N_6134);
or U9395 (N_9395,N_7083,N_6888);
nor U9396 (N_9396,N_6640,N_6968);
or U9397 (N_9397,N_7730,N_6568);
or U9398 (N_9398,N_6750,N_7889);
or U9399 (N_9399,N_6952,N_6096);
nand U9400 (N_9400,N_6497,N_7517);
xnor U9401 (N_9401,N_6346,N_7895);
or U9402 (N_9402,N_7027,N_6357);
xnor U9403 (N_9403,N_7597,N_6599);
xnor U9404 (N_9404,N_6169,N_6866);
nor U9405 (N_9405,N_6622,N_7598);
nor U9406 (N_9406,N_6806,N_6178);
nor U9407 (N_9407,N_7972,N_6335);
and U9408 (N_9408,N_6389,N_7284);
or U9409 (N_9409,N_6062,N_6717);
xor U9410 (N_9410,N_7591,N_7690);
xor U9411 (N_9411,N_7214,N_7108);
nor U9412 (N_9412,N_6742,N_6338);
nor U9413 (N_9413,N_6015,N_7797);
nand U9414 (N_9414,N_6397,N_7648);
nor U9415 (N_9415,N_6748,N_6612);
and U9416 (N_9416,N_6687,N_6304);
xor U9417 (N_9417,N_7891,N_7731);
and U9418 (N_9418,N_6150,N_6890);
xor U9419 (N_9419,N_7687,N_7010);
or U9420 (N_9420,N_6121,N_6903);
xnor U9421 (N_9421,N_7482,N_7463);
and U9422 (N_9422,N_6075,N_7361);
or U9423 (N_9423,N_6136,N_6678);
nor U9424 (N_9424,N_6647,N_7046);
and U9425 (N_9425,N_7602,N_7465);
or U9426 (N_9426,N_7381,N_6629);
nand U9427 (N_9427,N_7293,N_6505);
xnor U9428 (N_9428,N_7548,N_6341);
or U9429 (N_9429,N_6087,N_7354);
or U9430 (N_9430,N_6364,N_7237);
and U9431 (N_9431,N_6231,N_6049);
xnor U9432 (N_9432,N_7287,N_7294);
xnor U9433 (N_9433,N_7622,N_6261);
nand U9434 (N_9434,N_6221,N_6570);
xnor U9435 (N_9435,N_7921,N_6191);
xnor U9436 (N_9436,N_6695,N_6316);
or U9437 (N_9437,N_6038,N_6747);
nor U9438 (N_9438,N_6957,N_6768);
nor U9439 (N_9439,N_6450,N_7290);
and U9440 (N_9440,N_7218,N_7405);
xnor U9441 (N_9441,N_7806,N_6381);
nor U9442 (N_9442,N_6638,N_6746);
and U9443 (N_9443,N_6895,N_7396);
nand U9444 (N_9444,N_6589,N_6614);
xnor U9445 (N_9445,N_6853,N_7414);
and U9446 (N_9446,N_7495,N_6192);
nor U9447 (N_9447,N_7317,N_6280);
xor U9448 (N_9448,N_7776,N_6403);
xnor U9449 (N_9449,N_7533,N_6815);
nor U9450 (N_9450,N_6465,N_7198);
or U9451 (N_9451,N_7459,N_7629);
or U9452 (N_9452,N_7994,N_7106);
or U9453 (N_9453,N_6889,N_7670);
nand U9454 (N_9454,N_7723,N_7457);
or U9455 (N_9455,N_6191,N_6053);
and U9456 (N_9456,N_6828,N_7205);
xnor U9457 (N_9457,N_7372,N_7570);
and U9458 (N_9458,N_7564,N_6040);
or U9459 (N_9459,N_6124,N_6380);
and U9460 (N_9460,N_7433,N_6900);
or U9461 (N_9461,N_7052,N_7408);
or U9462 (N_9462,N_7759,N_6337);
nor U9463 (N_9463,N_7878,N_7495);
nor U9464 (N_9464,N_7043,N_7574);
nor U9465 (N_9465,N_7863,N_6995);
and U9466 (N_9466,N_6166,N_7323);
xor U9467 (N_9467,N_6608,N_7976);
and U9468 (N_9468,N_6177,N_6002);
nand U9469 (N_9469,N_6823,N_6149);
nor U9470 (N_9470,N_7914,N_7247);
nor U9471 (N_9471,N_6055,N_6691);
xor U9472 (N_9472,N_7746,N_7251);
or U9473 (N_9473,N_7177,N_7898);
xor U9474 (N_9474,N_6847,N_7293);
nor U9475 (N_9475,N_6620,N_6667);
or U9476 (N_9476,N_7698,N_7116);
and U9477 (N_9477,N_6029,N_6471);
xor U9478 (N_9478,N_6191,N_6903);
nor U9479 (N_9479,N_7218,N_7552);
nor U9480 (N_9480,N_6520,N_7840);
or U9481 (N_9481,N_7194,N_6897);
xnor U9482 (N_9482,N_7783,N_6593);
nor U9483 (N_9483,N_7848,N_6903);
nand U9484 (N_9484,N_6691,N_6137);
or U9485 (N_9485,N_6029,N_7605);
or U9486 (N_9486,N_7352,N_7302);
and U9487 (N_9487,N_6389,N_7271);
nor U9488 (N_9488,N_7681,N_6492);
or U9489 (N_9489,N_7906,N_7658);
and U9490 (N_9490,N_7297,N_7977);
nand U9491 (N_9491,N_6180,N_7778);
xor U9492 (N_9492,N_6075,N_6490);
nand U9493 (N_9493,N_7007,N_6938);
nor U9494 (N_9494,N_7763,N_7038);
nand U9495 (N_9495,N_6384,N_7543);
and U9496 (N_9496,N_6522,N_7024);
xnor U9497 (N_9497,N_7092,N_7388);
nor U9498 (N_9498,N_6610,N_6723);
xor U9499 (N_9499,N_7225,N_6490);
nand U9500 (N_9500,N_7597,N_6292);
xnor U9501 (N_9501,N_7619,N_6744);
xnor U9502 (N_9502,N_7965,N_6114);
or U9503 (N_9503,N_7433,N_6141);
or U9504 (N_9504,N_7260,N_6917);
nand U9505 (N_9505,N_7850,N_6287);
xor U9506 (N_9506,N_7885,N_7167);
or U9507 (N_9507,N_6098,N_6155);
nand U9508 (N_9508,N_6458,N_7720);
and U9509 (N_9509,N_7068,N_6837);
and U9510 (N_9510,N_7324,N_7469);
or U9511 (N_9511,N_6688,N_7668);
or U9512 (N_9512,N_7598,N_7735);
or U9513 (N_9513,N_7249,N_6870);
nand U9514 (N_9514,N_6741,N_6644);
nand U9515 (N_9515,N_6888,N_7160);
nor U9516 (N_9516,N_7541,N_7538);
or U9517 (N_9517,N_7361,N_6694);
nor U9518 (N_9518,N_7585,N_6260);
xnor U9519 (N_9519,N_6159,N_7074);
xor U9520 (N_9520,N_6057,N_7876);
or U9521 (N_9521,N_6759,N_6525);
nand U9522 (N_9522,N_7943,N_6429);
xor U9523 (N_9523,N_7898,N_6791);
xor U9524 (N_9524,N_6999,N_6569);
nor U9525 (N_9525,N_7840,N_6919);
or U9526 (N_9526,N_7289,N_6695);
nand U9527 (N_9527,N_7233,N_6910);
or U9528 (N_9528,N_7896,N_6983);
or U9529 (N_9529,N_6902,N_7547);
or U9530 (N_9530,N_7285,N_7768);
and U9531 (N_9531,N_7386,N_7804);
nand U9532 (N_9532,N_7888,N_7496);
and U9533 (N_9533,N_7072,N_6498);
nand U9534 (N_9534,N_7570,N_7472);
nand U9535 (N_9535,N_6973,N_7238);
nor U9536 (N_9536,N_7324,N_7394);
nand U9537 (N_9537,N_7412,N_6400);
xnor U9538 (N_9538,N_7905,N_7669);
and U9539 (N_9539,N_7890,N_6120);
xnor U9540 (N_9540,N_7668,N_7660);
nor U9541 (N_9541,N_7894,N_7409);
nor U9542 (N_9542,N_7900,N_7803);
nor U9543 (N_9543,N_6854,N_6713);
xor U9544 (N_9544,N_7757,N_7885);
xnor U9545 (N_9545,N_7494,N_7999);
or U9546 (N_9546,N_7639,N_6094);
nand U9547 (N_9547,N_6741,N_7615);
nand U9548 (N_9548,N_6440,N_6424);
xnor U9549 (N_9549,N_7402,N_6763);
and U9550 (N_9550,N_6269,N_7485);
and U9551 (N_9551,N_6820,N_7215);
nor U9552 (N_9552,N_7979,N_7828);
and U9553 (N_9553,N_7193,N_6719);
xor U9554 (N_9554,N_7930,N_7543);
xnor U9555 (N_9555,N_7568,N_6560);
or U9556 (N_9556,N_7807,N_6450);
xor U9557 (N_9557,N_6492,N_6088);
nand U9558 (N_9558,N_7121,N_6019);
nand U9559 (N_9559,N_7679,N_6504);
and U9560 (N_9560,N_7104,N_7975);
xor U9561 (N_9561,N_7581,N_7181);
nand U9562 (N_9562,N_6755,N_6535);
nand U9563 (N_9563,N_7518,N_7269);
and U9564 (N_9564,N_7040,N_6182);
or U9565 (N_9565,N_7585,N_7012);
nand U9566 (N_9566,N_6657,N_6362);
nand U9567 (N_9567,N_7343,N_7030);
nor U9568 (N_9568,N_7806,N_7887);
or U9569 (N_9569,N_7857,N_6410);
and U9570 (N_9570,N_7152,N_6766);
xnor U9571 (N_9571,N_7185,N_6592);
nand U9572 (N_9572,N_6083,N_7146);
or U9573 (N_9573,N_7554,N_6100);
or U9574 (N_9574,N_6755,N_7867);
nand U9575 (N_9575,N_7448,N_6021);
xnor U9576 (N_9576,N_6833,N_7794);
xor U9577 (N_9577,N_6187,N_7392);
and U9578 (N_9578,N_6886,N_6580);
nand U9579 (N_9579,N_7849,N_7663);
xnor U9580 (N_9580,N_6565,N_7256);
and U9581 (N_9581,N_6981,N_6279);
or U9582 (N_9582,N_6846,N_7507);
xnor U9583 (N_9583,N_7992,N_7437);
nor U9584 (N_9584,N_7019,N_6515);
or U9585 (N_9585,N_6200,N_7014);
and U9586 (N_9586,N_6976,N_6741);
xnor U9587 (N_9587,N_7523,N_7811);
or U9588 (N_9588,N_7674,N_6582);
and U9589 (N_9589,N_7479,N_6511);
xor U9590 (N_9590,N_6956,N_7265);
nand U9591 (N_9591,N_6074,N_7193);
xnor U9592 (N_9592,N_7443,N_6363);
nor U9593 (N_9593,N_7480,N_6431);
xnor U9594 (N_9594,N_7336,N_7153);
and U9595 (N_9595,N_6216,N_6885);
and U9596 (N_9596,N_6239,N_6993);
nand U9597 (N_9597,N_7026,N_6299);
xnor U9598 (N_9598,N_7012,N_7945);
and U9599 (N_9599,N_7517,N_7326);
or U9600 (N_9600,N_7031,N_6858);
and U9601 (N_9601,N_6805,N_6992);
nand U9602 (N_9602,N_6052,N_6085);
nor U9603 (N_9603,N_6701,N_6644);
nand U9604 (N_9604,N_7858,N_7088);
nor U9605 (N_9605,N_7217,N_7096);
nand U9606 (N_9606,N_7590,N_6348);
xor U9607 (N_9607,N_6605,N_7486);
nor U9608 (N_9608,N_6194,N_7123);
and U9609 (N_9609,N_6675,N_6672);
nand U9610 (N_9610,N_6811,N_7388);
nand U9611 (N_9611,N_7956,N_7470);
xor U9612 (N_9612,N_6081,N_6794);
nand U9613 (N_9613,N_6060,N_6792);
and U9614 (N_9614,N_6620,N_6047);
nand U9615 (N_9615,N_7558,N_7836);
nand U9616 (N_9616,N_6882,N_7653);
or U9617 (N_9617,N_7260,N_7484);
and U9618 (N_9618,N_7328,N_6296);
and U9619 (N_9619,N_7506,N_6989);
nand U9620 (N_9620,N_6261,N_6918);
xor U9621 (N_9621,N_7241,N_7976);
and U9622 (N_9622,N_7884,N_7512);
xnor U9623 (N_9623,N_6718,N_7169);
nor U9624 (N_9624,N_7564,N_7098);
xnor U9625 (N_9625,N_7268,N_7065);
xnor U9626 (N_9626,N_6384,N_6382);
and U9627 (N_9627,N_7510,N_7126);
or U9628 (N_9628,N_6177,N_7674);
nand U9629 (N_9629,N_7120,N_7809);
or U9630 (N_9630,N_7053,N_6484);
xnor U9631 (N_9631,N_6726,N_7618);
xnor U9632 (N_9632,N_7156,N_7214);
nor U9633 (N_9633,N_6819,N_6275);
xnor U9634 (N_9634,N_6123,N_6695);
xor U9635 (N_9635,N_7434,N_7030);
nor U9636 (N_9636,N_6480,N_7850);
nor U9637 (N_9637,N_6536,N_6859);
or U9638 (N_9638,N_7975,N_6173);
or U9639 (N_9639,N_6523,N_7523);
xor U9640 (N_9640,N_6037,N_6653);
and U9641 (N_9641,N_6926,N_6849);
and U9642 (N_9642,N_7657,N_6471);
xnor U9643 (N_9643,N_7069,N_7269);
xor U9644 (N_9644,N_6765,N_6979);
nand U9645 (N_9645,N_7742,N_7995);
and U9646 (N_9646,N_7471,N_7841);
nor U9647 (N_9647,N_7574,N_7178);
nor U9648 (N_9648,N_6902,N_6235);
or U9649 (N_9649,N_6057,N_7609);
xor U9650 (N_9650,N_7211,N_7766);
and U9651 (N_9651,N_7822,N_6172);
xor U9652 (N_9652,N_6782,N_7609);
nor U9653 (N_9653,N_7413,N_7192);
or U9654 (N_9654,N_7005,N_6530);
and U9655 (N_9655,N_6015,N_7264);
or U9656 (N_9656,N_6404,N_7282);
xnor U9657 (N_9657,N_7548,N_7989);
or U9658 (N_9658,N_7661,N_6147);
nand U9659 (N_9659,N_6569,N_6184);
xnor U9660 (N_9660,N_7064,N_6786);
or U9661 (N_9661,N_6572,N_7717);
and U9662 (N_9662,N_6472,N_7238);
xnor U9663 (N_9663,N_6631,N_6346);
nand U9664 (N_9664,N_7680,N_6574);
nand U9665 (N_9665,N_6989,N_7618);
nand U9666 (N_9666,N_6345,N_7097);
and U9667 (N_9667,N_6775,N_6655);
and U9668 (N_9668,N_6454,N_6583);
nand U9669 (N_9669,N_6848,N_6276);
or U9670 (N_9670,N_7641,N_6560);
xnor U9671 (N_9671,N_7128,N_6513);
nor U9672 (N_9672,N_6822,N_6503);
and U9673 (N_9673,N_6398,N_7586);
xor U9674 (N_9674,N_6922,N_6898);
and U9675 (N_9675,N_7714,N_6858);
nand U9676 (N_9676,N_6871,N_6990);
or U9677 (N_9677,N_7927,N_7524);
nand U9678 (N_9678,N_7409,N_7146);
xor U9679 (N_9679,N_6350,N_6944);
and U9680 (N_9680,N_7058,N_7268);
xor U9681 (N_9681,N_6502,N_6397);
or U9682 (N_9682,N_7984,N_6152);
nor U9683 (N_9683,N_6716,N_7469);
and U9684 (N_9684,N_7810,N_6554);
nor U9685 (N_9685,N_6128,N_7675);
or U9686 (N_9686,N_7808,N_7912);
or U9687 (N_9687,N_7210,N_6035);
or U9688 (N_9688,N_7573,N_7763);
xor U9689 (N_9689,N_7693,N_7951);
nor U9690 (N_9690,N_7787,N_6243);
and U9691 (N_9691,N_6257,N_6871);
or U9692 (N_9692,N_7151,N_6441);
and U9693 (N_9693,N_6848,N_6670);
nand U9694 (N_9694,N_6507,N_6731);
nand U9695 (N_9695,N_6563,N_6186);
nand U9696 (N_9696,N_6043,N_7976);
or U9697 (N_9697,N_7451,N_6141);
or U9698 (N_9698,N_6794,N_6067);
nor U9699 (N_9699,N_6232,N_7190);
xnor U9700 (N_9700,N_6968,N_6177);
or U9701 (N_9701,N_7315,N_7578);
and U9702 (N_9702,N_7591,N_7426);
nand U9703 (N_9703,N_7734,N_7575);
xor U9704 (N_9704,N_7825,N_6178);
or U9705 (N_9705,N_7500,N_7997);
and U9706 (N_9706,N_6716,N_7226);
xor U9707 (N_9707,N_6121,N_6297);
or U9708 (N_9708,N_7083,N_7027);
nor U9709 (N_9709,N_7968,N_7312);
or U9710 (N_9710,N_6347,N_7410);
and U9711 (N_9711,N_7139,N_6142);
nand U9712 (N_9712,N_7582,N_7387);
or U9713 (N_9713,N_6818,N_7804);
nand U9714 (N_9714,N_6398,N_7276);
nor U9715 (N_9715,N_6415,N_7347);
and U9716 (N_9716,N_6312,N_7445);
or U9717 (N_9717,N_6633,N_7330);
nor U9718 (N_9718,N_7902,N_6902);
or U9719 (N_9719,N_6218,N_6028);
nor U9720 (N_9720,N_7199,N_6145);
nor U9721 (N_9721,N_7034,N_6449);
nor U9722 (N_9722,N_6381,N_7019);
and U9723 (N_9723,N_6836,N_7418);
nor U9724 (N_9724,N_6952,N_6117);
and U9725 (N_9725,N_6823,N_6274);
nor U9726 (N_9726,N_7864,N_6016);
nand U9727 (N_9727,N_7332,N_6334);
and U9728 (N_9728,N_6707,N_6970);
nor U9729 (N_9729,N_6005,N_6584);
nand U9730 (N_9730,N_7238,N_6915);
nand U9731 (N_9731,N_6626,N_6656);
nand U9732 (N_9732,N_6118,N_6192);
nand U9733 (N_9733,N_7767,N_7012);
or U9734 (N_9734,N_6655,N_7127);
xor U9735 (N_9735,N_6349,N_7003);
nor U9736 (N_9736,N_6973,N_7149);
and U9737 (N_9737,N_6253,N_7442);
nor U9738 (N_9738,N_7596,N_6871);
or U9739 (N_9739,N_7917,N_7427);
xor U9740 (N_9740,N_7415,N_7339);
and U9741 (N_9741,N_7635,N_7977);
xor U9742 (N_9742,N_7540,N_7377);
nor U9743 (N_9743,N_7897,N_6252);
nand U9744 (N_9744,N_6549,N_7091);
nand U9745 (N_9745,N_6869,N_7629);
xor U9746 (N_9746,N_7239,N_7028);
xnor U9747 (N_9747,N_6302,N_6924);
nand U9748 (N_9748,N_6044,N_6490);
or U9749 (N_9749,N_6116,N_6028);
nand U9750 (N_9750,N_7718,N_6393);
nand U9751 (N_9751,N_7946,N_6801);
nor U9752 (N_9752,N_7446,N_6014);
nand U9753 (N_9753,N_7036,N_6193);
nor U9754 (N_9754,N_6915,N_6317);
nor U9755 (N_9755,N_7260,N_6511);
xor U9756 (N_9756,N_6383,N_7043);
nor U9757 (N_9757,N_7103,N_7991);
or U9758 (N_9758,N_6053,N_7016);
nand U9759 (N_9759,N_6594,N_6216);
or U9760 (N_9760,N_7104,N_6417);
nand U9761 (N_9761,N_7229,N_6448);
nand U9762 (N_9762,N_6384,N_6653);
or U9763 (N_9763,N_7771,N_6211);
and U9764 (N_9764,N_7980,N_6547);
or U9765 (N_9765,N_6004,N_7886);
nor U9766 (N_9766,N_7777,N_6598);
xnor U9767 (N_9767,N_7868,N_6340);
nor U9768 (N_9768,N_7500,N_7811);
nor U9769 (N_9769,N_6173,N_6485);
or U9770 (N_9770,N_6378,N_6898);
or U9771 (N_9771,N_6842,N_7173);
nor U9772 (N_9772,N_7338,N_6246);
and U9773 (N_9773,N_6008,N_7688);
or U9774 (N_9774,N_7190,N_7890);
nand U9775 (N_9775,N_6908,N_7066);
or U9776 (N_9776,N_6862,N_7591);
nor U9777 (N_9777,N_6316,N_7988);
nor U9778 (N_9778,N_6672,N_7647);
and U9779 (N_9779,N_7624,N_6483);
xor U9780 (N_9780,N_6476,N_7714);
and U9781 (N_9781,N_7156,N_7473);
xnor U9782 (N_9782,N_6746,N_7212);
or U9783 (N_9783,N_7737,N_6962);
nand U9784 (N_9784,N_7754,N_7627);
or U9785 (N_9785,N_7267,N_7651);
or U9786 (N_9786,N_6521,N_7616);
xnor U9787 (N_9787,N_7203,N_6020);
or U9788 (N_9788,N_7574,N_6786);
or U9789 (N_9789,N_6183,N_6308);
and U9790 (N_9790,N_6149,N_6914);
xor U9791 (N_9791,N_7632,N_7307);
and U9792 (N_9792,N_6502,N_6327);
or U9793 (N_9793,N_7150,N_7624);
and U9794 (N_9794,N_7028,N_6600);
and U9795 (N_9795,N_7924,N_6606);
xnor U9796 (N_9796,N_6979,N_6917);
nand U9797 (N_9797,N_7867,N_7741);
nor U9798 (N_9798,N_7437,N_6826);
xnor U9799 (N_9799,N_7314,N_6022);
or U9800 (N_9800,N_6717,N_7214);
and U9801 (N_9801,N_7840,N_6255);
and U9802 (N_9802,N_7146,N_6348);
nand U9803 (N_9803,N_7867,N_7219);
xor U9804 (N_9804,N_7896,N_7085);
xor U9805 (N_9805,N_7135,N_7100);
and U9806 (N_9806,N_6572,N_7158);
and U9807 (N_9807,N_7703,N_7165);
or U9808 (N_9808,N_6274,N_7458);
xor U9809 (N_9809,N_7590,N_6874);
nor U9810 (N_9810,N_7375,N_6388);
nand U9811 (N_9811,N_7251,N_7015);
and U9812 (N_9812,N_7381,N_6483);
xnor U9813 (N_9813,N_7659,N_7137);
xnor U9814 (N_9814,N_7711,N_7748);
and U9815 (N_9815,N_7828,N_6234);
nor U9816 (N_9816,N_6842,N_6373);
and U9817 (N_9817,N_6837,N_6739);
and U9818 (N_9818,N_6601,N_6426);
xor U9819 (N_9819,N_6339,N_7565);
xnor U9820 (N_9820,N_6316,N_6396);
xor U9821 (N_9821,N_6898,N_7260);
or U9822 (N_9822,N_7961,N_7023);
nand U9823 (N_9823,N_6955,N_7545);
nand U9824 (N_9824,N_7074,N_7061);
and U9825 (N_9825,N_6970,N_7363);
nand U9826 (N_9826,N_7065,N_6239);
xnor U9827 (N_9827,N_7294,N_7363);
or U9828 (N_9828,N_7405,N_6756);
and U9829 (N_9829,N_6920,N_7052);
and U9830 (N_9830,N_6916,N_7628);
nand U9831 (N_9831,N_6409,N_6654);
xor U9832 (N_9832,N_7754,N_7541);
and U9833 (N_9833,N_6188,N_6993);
or U9834 (N_9834,N_7224,N_6687);
xnor U9835 (N_9835,N_7569,N_6800);
and U9836 (N_9836,N_7274,N_6036);
and U9837 (N_9837,N_7177,N_7633);
nor U9838 (N_9838,N_7275,N_7374);
nand U9839 (N_9839,N_7824,N_6475);
or U9840 (N_9840,N_6773,N_6791);
nor U9841 (N_9841,N_7091,N_6394);
nand U9842 (N_9842,N_6514,N_7300);
xnor U9843 (N_9843,N_6281,N_6914);
nand U9844 (N_9844,N_6855,N_6728);
and U9845 (N_9845,N_7331,N_7018);
nor U9846 (N_9846,N_7192,N_6374);
nand U9847 (N_9847,N_6482,N_6379);
nor U9848 (N_9848,N_7685,N_7618);
and U9849 (N_9849,N_7584,N_7833);
nand U9850 (N_9850,N_6710,N_6771);
nor U9851 (N_9851,N_6206,N_6566);
nand U9852 (N_9852,N_7893,N_7621);
nand U9853 (N_9853,N_7464,N_6640);
and U9854 (N_9854,N_6392,N_6465);
nor U9855 (N_9855,N_7284,N_6652);
and U9856 (N_9856,N_7091,N_6412);
and U9857 (N_9857,N_6163,N_6677);
and U9858 (N_9858,N_6117,N_6112);
and U9859 (N_9859,N_7661,N_7267);
xnor U9860 (N_9860,N_7369,N_7590);
or U9861 (N_9861,N_7397,N_6747);
and U9862 (N_9862,N_6650,N_6340);
or U9863 (N_9863,N_6250,N_6599);
and U9864 (N_9864,N_7187,N_6068);
nor U9865 (N_9865,N_6815,N_7898);
and U9866 (N_9866,N_7374,N_6475);
and U9867 (N_9867,N_6910,N_7614);
nand U9868 (N_9868,N_7784,N_7096);
nand U9869 (N_9869,N_7599,N_6092);
xnor U9870 (N_9870,N_6958,N_6338);
nand U9871 (N_9871,N_7927,N_6756);
nand U9872 (N_9872,N_6672,N_7352);
nand U9873 (N_9873,N_6242,N_6018);
xor U9874 (N_9874,N_6045,N_6198);
and U9875 (N_9875,N_7790,N_7168);
nand U9876 (N_9876,N_7820,N_7621);
and U9877 (N_9877,N_7404,N_7392);
nand U9878 (N_9878,N_7262,N_7540);
and U9879 (N_9879,N_7896,N_6584);
nand U9880 (N_9880,N_6495,N_7907);
nor U9881 (N_9881,N_6866,N_6120);
nor U9882 (N_9882,N_7623,N_7987);
nand U9883 (N_9883,N_7063,N_6534);
or U9884 (N_9884,N_6304,N_6937);
nor U9885 (N_9885,N_6499,N_7335);
nor U9886 (N_9886,N_6713,N_7667);
nor U9887 (N_9887,N_6439,N_7693);
nand U9888 (N_9888,N_7772,N_7739);
nand U9889 (N_9889,N_6727,N_6582);
nor U9890 (N_9890,N_6260,N_6114);
nor U9891 (N_9891,N_6262,N_6623);
nor U9892 (N_9892,N_7629,N_6261);
xor U9893 (N_9893,N_7533,N_6620);
xnor U9894 (N_9894,N_6196,N_6778);
nor U9895 (N_9895,N_6211,N_7895);
nand U9896 (N_9896,N_7885,N_7175);
nand U9897 (N_9897,N_7650,N_7557);
nor U9898 (N_9898,N_7695,N_7975);
or U9899 (N_9899,N_7864,N_6540);
nor U9900 (N_9900,N_7744,N_6456);
xor U9901 (N_9901,N_6322,N_6548);
nor U9902 (N_9902,N_7795,N_6562);
nor U9903 (N_9903,N_6516,N_6904);
xor U9904 (N_9904,N_7778,N_7753);
nand U9905 (N_9905,N_6118,N_7664);
nand U9906 (N_9906,N_7484,N_6102);
nor U9907 (N_9907,N_6936,N_6066);
and U9908 (N_9908,N_6045,N_7609);
or U9909 (N_9909,N_6689,N_7398);
xnor U9910 (N_9910,N_7865,N_7435);
and U9911 (N_9911,N_6845,N_6437);
or U9912 (N_9912,N_7551,N_7150);
xor U9913 (N_9913,N_7608,N_6359);
or U9914 (N_9914,N_6139,N_6595);
and U9915 (N_9915,N_6191,N_6979);
nand U9916 (N_9916,N_6282,N_6320);
nor U9917 (N_9917,N_7850,N_7596);
or U9918 (N_9918,N_7591,N_7918);
and U9919 (N_9919,N_6171,N_7519);
nand U9920 (N_9920,N_6372,N_7364);
nor U9921 (N_9921,N_6288,N_6073);
xnor U9922 (N_9922,N_6134,N_7521);
or U9923 (N_9923,N_6733,N_6252);
xor U9924 (N_9924,N_7577,N_6077);
nand U9925 (N_9925,N_6624,N_7995);
or U9926 (N_9926,N_7861,N_7642);
nand U9927 (N_9927,N_6570,N_7690);
nand U9928 (N_9928,N_7320,N_7442);
nand U9929 (N_9929,N_7851,N_6695);
nor U9930 (N_9930,N_7393,N_7124);
nand U9931 (N_9931,N_6563,N_7871);
xor U9932 (N_9932,N_7538,N_6841);
or U9933 (N_9933,N_6292,N_7362);
and U9934 (N_9934,N_6048,N_7446);
or U9935 (N_9935,N_7765,N_7091);
nand U9936 (N_9936,N_7885,N_6058);
nor U9937 (N_9937,N_7109,N_6087);
and U9938 (N_9938,N_6232,N_7629);
xor U9939 (N_9939,N_7405,N_7401);
xnor U9940 (N_9940,N_7667,N_6308);
xnor U9941 (N_9941,N_6152,N_7852);
nand U9942 (N_9942,N_7233,N_7846);
nor U9943 (N_9943,N_6229,N_7389);
nor U9944 (N_9944,N_6678,N_7028);
nand U9945 (N_9945,N_7792,N_6900);
and U9946 (N_9946,N_7098,N_7857);
xor U9947 (N_9947,N_6312,N_6139);
or U9948 (N_9948,N_7591,N_7455);
or U9949 (N_9949,N_7332,N_7215);
xnor U9950 (N_9950,N_6101,N_7015);
xnor U9951 (N_9951,N_7150,N_7270);
nor U9952 (N_9952,N_7653,N_6267);
nand U9953 (N_9953,N_6552,N_7482);
or U9954 (N_9954,N_6699,N_6885);
nand U9955 (N_9955,N_6855,N_6425);
and U9956 (N_9956,N_6730,N_6355);
or U9957 (N_9957,N_7828,N_7550);
and U9958 (N_9958,N_7221,N_7240);
or U9959 (N_9959,N_7667,N_6165);
nand U9960 (N_9960,N_7049,N_7267);
or U9961 (N_9961,N_7182,N_6858);
xnor U9962 (N_9962,N_7286,N_6633);
xor U9963 (N_9963,N_7666,N_7728);
and U9964 (N_9964,N_7902,N_7405);
and U9965 (N_9965,N_6135,N_6586);
or U9966 (N_9966,N_7365,N_6726);
nor U9967 (N_9967,N_6265,N_7097);
or U9968 (N_9968,N_6065,N_6582);
and U9969 (N_9969,N_6241,N_6997);
nor U9970 (N_9970,N_7425,N_7451);
nor U9971 (N_9971,N_6078,N_7821);
xnor U9972 (N_9972,N_7955,N_7371);
and U9973 (N_9973,N_6355,N_6396);
and U9974 (N_9974,N_6106,N_7496);
xor U9975 (N_9975,N_7095,N_6887);
and U9976 (N_9976,N_6774,N_6620);
nor U9977 (N_9977,N_6149,N_6762);
and U9978 (N_9978,N_7325,N_7358);
xor U9979 (N_9979,N_6301,N_7259);
or U9980 (N_9980,N_7281,N_6152);
and U9981 (N_9981,N_6901,N_6825);
nor U9982 (N_9982,N_6811,N_6462);
nor U9983 (N_9983,N_7606,N_6850);
or U9984 (N_9984,N_6045,N_6474);
nand U9985 (N_9985,N_7298,N_6147);
xor U9986 (N_9986,N_6511,N_7718);
nand U9987 (N_9987,N_6281,N_7668);
xor U9988 (N_9988,N_6917,N_7979);
and U9989 (N_9989,N_7271,N_7874);
and U9990 (N_9990,N_6368,N_7942);
and U9991 (N_9991,N_6097,N_7079);
xnor U9992 (N_9992,N_7662,N_6868);
or U9993 (N_9993,N_6858,N_6950);
nand U9994 (N_9994,N_7884,N_7168);
nand U9995 (N_9995,N_6380,N_6464);
and U9996 (N_9996,N_7719,N_7678);
or U9997 (N_9997,N_7167,N_7298);
nor U9998 (N_9998,N_6800,N_7507);
and U9999 (N_9999,N_6586,N_7446);
xnor U10000 (N_10000,N_8128,N_9804);
nor U10001 (N_10001,N_8436,N_9624);
or U10002 (N_10002,N_9473,N_9150);
or U10003 (N_10003,N_9651,N_9011);
or U10004 (N_10004,N_9870,N_9723);
and U10005 (N_10005,N_9288,N_9520);
nand U10006 (N_10006,N_9866,N_9340);
or U10007 (N_10007,N_9951,N_9964);
nand U10008 (N_10008,N_8832,N_8684);
and U10009 (N_10009,N_9675,N_9263);
xor U10010 (N_10010,N_9072,N_9500);
or U10011 (N_10011,N_8857,N_8715);
nand U10012 (N_10012,N_8126,N_9111);
nand U10013 (N_10013,N_8762,N_9927);
or U10014 (N_10014,N_9602,N_9930);
xnor U10015 (N_10015,N_8936,N_8217);
nand U10016 (N_10016,N_8879,N_8340);
nand U10017 (N_10017,N_8183,N_9643);
or U10018 (N_10018,N_8500,N_9060);
nor U10019 (N_10019,N_9338,N_9783);
or U10020 (N_10020,N_8804,N_8605);
nand U10021 (N_10021,N_9911,N_9204);
or U10022 (N_10022,N_8945,N_9616);
xnor U10023 (N_10023,N_8694,N_9026);
xnor U10024 (N_10024,N_9317,N_9403);
xnor U10025 (N_10025,N_9692,N_8142);
nor U10026 (N_10026,N_9115,N_9016);
nor U10027 (N_10027,N_8344,N_8181);
nor U10028 (N_10028,N_8711,N_9640);
nor U10029 (N_10029,N_8134,N_8251);
and U10030 (N_10030,N_8587,N_9428);
and U10031 (N_10031,N_9599,N_9265);
xnor U10032 (N_10032,N_8187,N_8488);
xnor U10033 (N_10033,N_9537,N_9677);
or U10034 (N_10034,N_9375,N_9237);
nand U10035 (N_10035,N_8039,N_8652);
xnor U10036 (N_10036,N_8678,N_8428);
nand U10037 (N_10037,N_8672,N_9733);
nor U10038 (N_10038,N_9841,N_9147);
nor U10039 (N_10039,N_9541,N_8115);
nand U10040 (N_10040,N_8537,N_9736);
nand U10041 (N_10041,N_8974,N_9515);
nor U10042 (N_10042,N_9716,N_9217);
and U10043 (N_10043,N_9769,N_9580);
xnor U10044 (N_10044,N_9626,N_8151);
nand U10045 (N_10045,N_8878,N_9853);
nand U10046 (N_10046,N_8314,N_8411);
nand U10047 (N_10047,N_9314,N_9980);
and U10048 (N_10048,N_8498,N_8419);
and U10049 (N_10049,N_9835,N_8139);
nor U10050 (N_10050,N_8862,N_8267);
nand U10051 (N_10051,N_8642,N_9944);
and U10052 (N_10052,N_8035,N_9482);
xor U10053 (N_10053,N_8268,N_8797);
xor U10054 (N_10054,N_8746,N_8034);
xor U10055 (N_10055,N_8273,N_8552);
nand U10056 (N_10056,N_8095,N_9421);
nor U10057 (N_10057,N_9502,N_8310);
nor U10058 (N_10058,N_9195,N_9591);
nor U10059 (N_10059,N_8157,N_8303);
or U10060 (N_10060,N_9902,N_8438);
nand U10061 (N_10061,N_9724,N_9793);
xnor U10062 (N_10062,N_9499,N_9647);
or U10063 (N_10063,N_8640,N_8188);
and U10064 (N_10064,N_9846,N_8019);
nand U10065 (N_10065,N_9109,N_9123);
nand U10066 (N_10066,N_9874,N_8688);
xnor U10067 (N_10067,N_8647,N_9734);
xnor U10068 (N_10068,N_8466,N_8323);
xnor U10069 (N_10069,N_8673,N_8405);
and U10070 (N_10070,N_9729,N_9711);
or U10071 (N_10071,N_9255,N_8546);
nand U10072 (N_10072,N_9176,N_8225);
nand U10073 (N_10073,N_8734,N_9884);
nor U10074 (N_10074,N_8534,N_9518);
nor U10075 (N_10075,N_9100,N_8830);
nand U10076 (N_10076,N_9023,N_8901);
nand U10077 (N_10077,N_8088,N_8713);
and U10078 (N_10078,N_8368,N_9277);
and U10079 (N_10079,N_8686,N_8728);
and U10080 (N_10080,N_8279,N_8361);
nor U10081 (N_10081,N_8881,N_8121);
xor U10082 (N_10082,N_9781,N_9452);
or U10083 (N_10083,N_9092,N_9068);
nor U10084 (N_10084,N_9410,N_8621);
nor U10085 (N_10085,N_8650,N_9654);
xnor U10086 (N_10086,N_9311,N_9163);
xor U10087 (N_10087,N_8433,N_8698);
and U10088 (N_10088,N_8743,N_8401);
nor U10089 (N_10089,N_8031,N_8471);
nor U10090 (N_10090,N_8275,N_8493);
xnor U10091 (N_10091,N_9230,N_9800);
nand U10092 (N_10092,N_9384,N_8354);
nor U10093 (N_10093,N_9212,N_9046);
and U10094 (N_10094,N_8767,N_9628);
nand U10095 (N_10095,N_9620,N_9069);
xor U10096 (N_10096,N_9064,N_9320);
and U10097 (N_10097,N_8016,N_8150);
xor U10098 (N_10098,N_9462,N_8021);
or U10099 (N_10099,N_9858,N_9519);
xnor U10100 (N_10100,N_9816,N_9094);
nor U10101 (N_10101,N_9083,N_9810);
nand U10102 (N_10102,N_9901,N_9666);
and U10103 (N_10103,N_9778,N_8331);
and U10104 (N_10104,N_9637,N_9169);
or U10105 (N_10105,N_9514,N_9638);
nor U10106 (N_10106,N_9946,N_8210);
xnor U10107 (N_10107,N_8547,N_9542);
nor U10108 (N_10108,N_8302,N_9659);
nor U10109 (N_10109,N_8064,N_9942);
nor U10110 (N_10110,N_8330,N_8001);
or U10111 (N_10111,N_8192,N_9743);
and U10112 (N_10112,N_8564,N_8292);
nand U10113 (N_10113,N_9074,N_9614);
or U10114 (N_10114,N_8399,N_9306);
or U10115 (N_10115,N_8083,N_8998);
and U10116 (N_10116,N_9528,N_9243);
and U10117 (N_10117,N_9059,N_9272);
xor U10118 (N_10118,N_9012,N_9594);
xnor U10119 (N_10119,N_9553,N_8750);
nand U10120 (N_10120,N_9814,N_8925);
or U10121 (N_10121,N_8404,N_8172);
nand U10122 (N_10122,N_8844,N_8449);
xnor U10123 (N_10123,N_9408,N_9953);
xnor U10124 (N_10124,N_9044,N_8032);
or U10125 (N_10125,N_8165,N_8924);
xor U10126 (N_10126,N_8696,N_8730);
nand U10127 (N_10127,N_9075,N_8784);
or U10128 (N_10128,N_9376,N_8620);
and U10129 (N_10129,N_8484,N_9106);
and U10130 (N_10130,N_8699,N_9459);
xor U10131 (N_10131,N_8491,N_9439);
xor U10132 (N_10132,N_9360,N_9685);
nor U10133 (N_10133,N_8478,N_8232);
nand U10134 (N_10134,N_9973,N_8148);
nand U10135 (N_10135,N_8934,N_8381);
and U10136 (N_10136,N_8454,N_9895);
xnor U10137 (N_10137,N_9903,N_8495);
or U10138 (N_10138,N_9291,N_8635);
or U10139 (N_10139,N_8507,N_8984);
or U10140 (N_10140,N_9621,N_8004);
nand U10141 (N_10141,N_8231,N_8006);
nor U10142 (N_10142,N_8780,N_9513);
and U10143 (N_10143,N_9406,N_9251);
nand U10144 (N_10144,N_8072,N_8884);
nand U10145 (N_10145,N_8068,N_9374);
nand U10146 (N_10146,N_9145,N_9142);
xor U10147 (N_10147,N_8983,N_9921);
xor U10148 (N_10148,N_8062,N_8946);
nand U10149 (N_10149,N_9290,N_8972);
nand U10150 (N_10150,N_9745,N_9777);
nand U10151 (N_10151,N_9129,N_8332);
nor U10152 (N_10152,N_9947,N_9907);
and U10153 (N_10153,N_8837,N_8918);
nor U10154 (N_10154,N_9538,N_9674);
nand U10155 (N_10155,N_8420,N_8362);
nor U10156 (N_10156,N_8350,N_9160);
xor U10157 (N_10157,N_9448,N_8453);
nor U10158 (N_10158,N_8113,N_9008);
and U10159 (N_10159,N_9573,N_8245);
nor U10160 (N_10160,N_9634,N_9357);
xor U10161 (N_10161,N_9019,N_9371);
nor U10162 (N_10162,N_9052,N_9885);
nor U10163 (N_10163,N_8586,N_9707);
and U10164 (N_10164,N_9367,N_9209);
or U10165 (N_10165,N_9605,N_8900);
xor U10166 (N_10166,N_9969,N_8732);
nand U10167 (N_10167,N_9632,N_9863);
nor U10168 (N_10168,N_8477,N_9372);
and U10169 (N_10169,N_8395,N_9557);
and U10170 (N_10170,N_8549,N_9709);
and U10171 (N_10171,N_9655,N_8435);
nand U10172 (N_10172,N_9569,N_9466);
and U10173 (N_10173,N_9154,N_9429);
xor U10174 (N_10174,N_9896,N_8515);
nor U10175 (N_10175,N_8705,N_9963);
xnor U10176 (N_10176,N_9388,N_9392);
or U10177 (N_10177,N_9050,N_9323);
xnor U10178 (N_10178,N_9919,N_8197);
and U10179 (N_10179,N_8511,N_8682);
or U10180 (N_10180,N_8342,N_8882);
nand U10181 (N_10181,N_9307,N_9104);
and U10182 (N_10182,N_9970,N_9764);
or U10183 (N_10183,N_8608,N_8423);
and U10184 (N_10184,N_8770,N_8513);
nor U10185 (N_10185,N_8313,N_8677);
or U10186 (N_10186,N_8297,N_9236);
xnor U10187 (N_10187,N_8845,N_9521);
and U10188 (N_10188,N_8927,N_8379);
or U10189 (N_10189,N_8285,N_8056);
nor U10190 (N_10190,N_9268,N_9547);
and U10191 (N_10191,N_8129,N_9292);
nand U10192 (N_10192,N_9344,N_9840);
and U10193 (N_10193,N_9164,N_8645);
nand U10194 (N_10194,N_9425,N_8123);
nor U10195 (N_10195,N_9713,N_8893);
nor U10196 (N_10196,N_8080,N_9890);
and U10197 (N_10197,N_9319,N_8262);
and U10198 (N_10198,N_9939,N_9631);
nor U10199 (N_10199,N_9759,N_9775);
nor U10200 (N_10200,N_8809,N_9641);
and U10201 (N_10201,N_9510,N_9281);
xnor U10202 (N_10202,N_8124,N_8013);
and U10203 (N_10203,N_8207,N_8119);
nand U10204 (N_10204,N_9851,N_8270);
nand U10205 (N_10205,N_9447,N_9022);
nor U10206 (N_10206,N_9394,N_9586);
and U10207 (N_10207,N_8191,N_9102);
xnor U10208 (N_10208,N_9107,N_8982);
xor U10209 (N_10209,N_8400,N_9414);
or U10210 (N_10210,N_9161,N_9167);
nand U10211 (N_10211,N_8445,N_9181);
xor U10212 (N_10212,N_9952,N_9994);
and U10213 (N_10213,N_8753,N_9999);
or U10214 (N_10214,N_9219,N_8514);
xnor U10215 (N_10215,N_8667,N_9125);
nand U10216 (N_10216,N_8594,N_9748);
and U10217 (N_10217,N_9278,N_8458);
nand U10218 (N_10218,N_8196,N_9198);
and U10219 (N_10219,N_9561,N_9047);
and U10220 (N_10220,N_8920,N_9303);
or U10221 (N_10221,N_8108,N_9279);
or U10222 (N_10222,N_8014,N_9875);
or U10223 (N_10223,N_9861,N_9527);
nand U10224 (N_10224,N_8455,N_9691);
xnor U10225 (N_10225,N_9043,N_9218);
nand U10226 (N_10226,N_9923,N_9078);
nor U10227 (N_10227,N_9006,N_9767);
or U10228 (N_10228,N_8193,N_9752);
and U10229 (N_10229,N_8280,N_9451);
or U10230 (N_10230,N_8120,N_9698);
xor U10231 (N_10231,N_8931,N_9868);
nor U10232 (N_10232,N_9088,N_9787);
xnor U10233 (N_10233,N_9049,N_9289);
xor U10234 (N_10234,N_9581,N_9152);
nor U10235 (N_10235,N_8364,N_8155);
nand U10236 (N_10236,N_9472,N_8200);
and U10237 (N_10237,N_9828,N_9113);
and U10238 (N_10238,N_9133,N_8276);
and U10239 (N_10239,N_8289,N_8363);
nand U10240 (N_10240,N_8629,N_9475);
xor U10241 (N_10241,N_9867,N_9048);
and U10242 (N_10242,N_9487,N_8066);
xor U10243 (N_10243,N_9501,N_8567);
and U10244 (N_10244,N_9131,N_9393);
nor U10245 (N_10245,N_8973,N_9132);
xor U10246 (N_10246,N_8863,N_9757);
nand U10247 (N_10247,N_9018,N_9928);
or U10248 (N_10248,N_8136,N_8177);
and U10249 (N_10249,N_8287,N_8539);
xnor U10250 (N_10250,N_9997,N_8295);
nand U10251 (N_10251,N_9996,N_9668);
and U10252 (N_10252,N_8359,N_9894);
or U10253 (N_10253,N_9409,N_8530);
nand U10254 (N_10254,N_9812,N_8706);
or U10255 (N_10255,N_9080,N_8798);
nor U10256 (N_10256,N_9266,N_8748);
nor U10257 (N_10257,N_8990,N_8560);
or U10258 (N_10258,N_8503,N_8729);
xor U10259 (N_10259,N_9465,N_8612);
and U10260 (N_10260,N_8710,N_8131);
and U10261 (N_10261,N_9207,N_8456);
and U10262 (N_10262,N_8545,N_9968);
or U10263 (N_10263,N_8459,N_9180);
or U10264 (N_10264,N_9456,N_8649);
nor U10265 (N_10265,N_9979,N_8548);
nor U10266 (N_10266,N_9534,N_8130);
and U10267 (N_10267,N_9546,N_8074);
nor U10268 (N_10268,N_9956,N_9837);
and U10269 (N_10269,N_9054,N_8807);
nor U10270 (N_10270,N_8348,N_9672);
xor U10271 (N_10271,N_8860,N_8833);
and U10272 (N_10272,N_9726,N_8956);
nor U10273 (N_10273,N_8628,N_8389);
or U10274 (N_10274,N_9108,N_9784);
nand U10275 (N_10275,N_8087,N_8308);
nand U10276 (N_10276,N_9995,N_9438);
nor U10277 (N_10277,N_9248,N_9187);
and U10278 (N_10278,N_9583,N_9157);
xnor U10279 (N_10279,N_9938,N_8749);
nand U10280 (N_10280,N_9335,N_8570);
nor U10281 (N_10281,N_8194,N_9873);
and U10282 (N_10282,N_8542,N_8446);
xnor U10283 (N_10283,N_8300,N_9765);
and U10284 (N_10284,N_9084,N_8333);
nor U10285 (N_10285,N_8106,N_8334);
xnor U10286 (N_10286,N_8992,N_9441);
and U10287 (N_10287,N_9257,N_9240);
or U10288 (N_10288,N_8215,N_8818);
xnor U10289 (N_10289,N_9790,N_8853);
nand U10290 (N_10290,N_8100,N_9474);
nor U10291 (N_10291,N_8221,N_8049);
nor U10292 (N_10292,N_9305,N_8601);
xnor U10293 (N_10293,N_9315,N_9378);
nor U10294 (N_10294,N_8098,N_8376);
nor U10295 (N_10295,N_9639,N_9860);
nand U10296 (N_10296,N_9433,N_8665);
or U10297 (N_10297,N_9168,N_9398);
nor U10298 (N_10298,N_9854,N_9916);
and U10299 (N_10299,N_8718,N_8854);
and U10300 (N_10300,N_9227,N_8025);
nor U10301 (N_10301,N_8864,N_9313);
and U10302 (N_10302,N_9975,N_8581);
or U10303 (N_10303,N_9101,N_9222);
xor U10304 (N_10304,N_9238,N_9509);
xor U10305 (N_10305,N_8774,N_9066);
nor U10306 (N_10306,N_9029,N_8916);
nor U10307 (N_10307,N_9269,N_9937);
nor U10308 (N_10308,N_8464,N_9865);
nor U10309 (N_10309,N_8159,N_8712);
and U10310 (N_10310,N_8805,N_8906);
and U10311 (N_10311,N_8257,N_8182);
and U10312 (N_10312,N_8583,N_9690);
and U10313 (N_10313,N_8265,N_9912);
or U10314 (N_10314,N_8380,N_9780);
nand U10315 (N_10315,N_8573,N_8737);
and U10316 (N_10316,N_9663,N_8761);
xnor U10317 (N_10317,N_8917,N_9330);
xor U10318 (N_10318,N_9548,N_9529);
and U10319 (N_10319,N_9427,N_8700);
nor U10320 (N_10320,N_8084,N_8063);
or U10321 (N_10321,N_9119,N_8460);
xnor U10322 (N_10322,N_9401,N_9310);
xnor U10323 (N_10323,N_8118,N_9485);
nor U10324 (N_10324,N_8271,N_9040);
nor U10325 (N_10325,N_8434,N_8824);
nor U10326 (N_10326,N_8790,N_8681);
or U10327 (N_10327,N_9091,N_8887);
nand U10328 (N_10328,N_8429,N_8637);
and U10329 (N_10329,N_8747,N_8768);
xnor U10330 (N_10330,N_8791,N_9825);
or U10331 (N_10331,N_8950,N_9214);
or U10332 (N_10332,N_9194,N_9366);
xor U10333 (N_10333,N_8969,N_9977);
nor U10334 (N_10334,N_9116,N_8377);
nand U10335 (N_10335,N_8226,N_9353);
and U10336 (N_10336,N_8885,N_8632);
nor U10337 (N_10337,N_8859,N_8209);
or U10338 (N_10338,N_9706,N_9223);
xnor U10339 (N_10339,N_8024,N_9817);
xnor U10340 (N_10340,N_8141,N_8625);
or U10341 (N_10341,N_8851,N_8995);
nor U10342 (N_10342,N_8352,N_8501);
or U10343 (N_10343,N_9680,N_8284);
nor U10344 (N_10344,N_8028,N_9185);
nand U10345 (N_10345,N_8373,N_9148);
and U10346 (N_10346,N_8994,N_8961);
nand U10347 (N_10347,N_8759,N_9823);
nand U10348 (N_10348,N_9796,N_9516);
nand U10349 (N_10349,N_8259,N_9244);
xor U10350 (N_10350,N_8651,N_9191);
xor U10351 (N_10351,N_9717,N_8913);
and U10352 (N_10352,N_8962,N_9124);
nand U10353 (N_10353,N_9559,N_9146);
or U10354 (N_10354,N_8687,N_8840);
nand U10355 (N_10355,N_8258,N_9241);
xnor U10356 (N_10356,N_9683,N_9171);
nor U10357 (N_10357,N_8942,N_8320);
nand U10358 (N_10358,N_9792,N_8092);
nor U10359 (N_10359,N_8050,N_9824);
xor U10360 (N_10360,N_9629,N_8657);
nand U10361 (N_10361,N_9155,N_8149);
nor U10362 (N_10362,N_9469,N_9574);
xnor U10363 (N_10363,N_8216,N_9089);
nor U10364 (N_10364,N_9431,N_8075);
nand U10365 (N_10365,N_8988,N_9434);
nand U10366 (N_10366,N_8921,N_9976);
xor U10367 (N_10367,N_8926,N_9972);
nor U10368 (N_10368,N_8133,N_9962);
and U10369 (N_10369,N_8058,N_9028);
or U10370 (N_10370,N_9369,N_8356);
xnor U10371 (N_10371,N_9551,N_8494);
xnor U10372 (N_10372,N_9387,N_8538);
and U10373 (N_10373,N_8152,N_9750);
or U10374 (N_10374,N_9261,N_8481);
xnor U10375 (N_10375,N_9184,N_8264);
nor U10376 (N_10376,N_8427,N_9373);
nor U10377 (N_10377,N_8042,N_8079);
nor U10378 (N_10378,N_8073,N_8071);
or U10379 (N_10379,N_8755,N_9785);
or U10380 (N_10380,N_9768,N_9437);
or U10381 (N_10381,N_8440,N_9036);
and U10382 (N_10382,N_9522,N_9460);
and U10383 (N_10383,N_8590,N_8680);
xnor U10384 (N_10384,N_8848,N_9199);
or U10385 (N_10385,N_8451,N_9596);
or U10386 (N_10386,N_9200,N_8236);
nor U10387 (N_10387,N_9495,N_9924);
or U10388 (N_10388,N_8958,N_8817);
and U10389 (N_10389,N_8283,N_9744);
nor U10390 (N_10390,N_8278,N_8843);
or U10391 (N_10391,N_9694,N_9604);
or U10392 (N_10392,N_9014,N_9983);
nor U10393 (N_10393,N_8140,N_9235);
or U10394 (N_10394,N_9253,N_8967);
nor U10395 (N_10395,N_8989,N_9929);
xor U10396 (N_10396,N_8529,N_9267);
nor U10397 (N_10397,N_9887,N_9440);
xor U10398 (N_10398,N_9359,N_8229);
or U10399 (N_10399,N_8002,N_8358);
nor U10400 (N_10400,N_8815,N_9280);
xnor U10401 (N_10401,N_8987,N_9332);
or U10402 (N_10402,N_8568,N_9159);
or U10403 (N_10403,N_8383,N_8899);
nand U10404 (N_10404,N_9355,N_9662);
nor U10405 (N_10405,N_8430,N_8574);
nand U10406 (N_10406,N_9749,N_9284);
nand U10407 (N_10407,N_9153,N_8369);
and U10408 (N_10408,N_8668,N_9435);
or U10409 (N_10409,N_8146,N_9779);
xnor U10410 (N_10410,N_9705,N_9708);
nor U10411 (N_10411,N_9611,N_8611);
nor U10412 (N_10412,N_8719,N_8374);
nor U10413 (N_10413,N_8658,N_8971);
nand U10414 (N_10414,N_8431,N_8528);
nand U10415 (N_10415,N_9216,N_9587);
nor U10416 (N_10416,N_9318,N_9986);
and U10417 (N_10417,N_8085,N_9943);
xor U10418 (N_10418,N_9467,N_8822);
or U10419 (N_10419,N_8644,N_8442);
nor U10420 (N_10420,N_9888,N_9714);
nand U10421 (N_10421,N_9170,N_8486);
nand U10422 (N_10422,N_8029,N_8007);
xnor U10423 (N_10423,N_8469,N_9966);
or U10424 (N_10424,N_8826,N_9037);
or U10425 (N_10425,N_9525,N_9879);
and U10426 (N_10426,N_9543,N_8518);
xnor U10427 (N_10427,N_9051,N_8892);
xnor U10428 (N_10428,N_8615,N_9117);
and U10429 (N_10429,N_8609,N_9772);
or U10430 (N_10430,N_9090,N_8089);
xnor U10431 (N_10431,N_8010,N_8889);
or U10432 (N_10432,N_8444,N_9606);
and U10433 (N_10433,N_9991,N_8891);
nand U10434 (N_10434,N_8597,N_9166);
xor U10435 (N_10435,N_9678,N_8653);
nand U10436 (N_10436,N_8160,N_8298);
nand U10437 (N_10437,N_9661,N_9085);
nand U10438 (N_10438,N_9601,N_8536);
nor U10439 (N_10439,N_8145,N_9815);
nand U10440 (N_10440,N_9762,N_8555);
or U10441 (N_10441,N_8170,N_8163);
nand U10442 (N_10442,N_8041,N_9880);
xnor U10443 (N_10443,N_8877,N_8318);
nor U10444 (N_10444,N_9489,N_9498);
xor U10445 (N_10445,N_8616,N_8269);
nor U10446 (N_10446,N_9756,N_8388);
nor U10447 (N_10447,N_9576,N_8669);
xnor U10448 (N_10448,N_8742,N_8102);
or U10449 (N_10449,N_8156,N_9789);
nor U10450 (N_10450,N_9301,N_9595);
nor U10451 (N_10451,N_9417,N_8176);
xor U10452 (N_10452,N_9635,N_9915);
nand U10453 (N_10453,N_8964,N_9354);
and U10454 (N_10454,N_9886,N_9533);
xor U10455 (N_10455,N_9883,N_8046);
xor U10456 (N_10456,N_8252,N_8497);
or U10457 (N_10457,N_8094,N_9827);
nand U10458 (N_10458,N_9327,N_8527);
xor U10459 (N_10459,N_9897,N_9177);
nand U10460 (N_10460,N_8949,N_9038);
nor U10461 (N_10461,N_9331,N_8296);
nand U10462 (N_10462,N_8099,N_8544);
xor U10463 (N_10463,N_9656,N_8754);
nor U10464 (N_10464,N_9343,N_9712);
or U10465 (N_10465,N_8836,N_9027);
nand U10466 (N_10466,N_9847,N_8968);
nand U10467 (N_10467,N_9348,N_9377);
nand U10468 (N_10468,N_9247,N_8726);
or U10469 (N_10469,N_9249,N_9696);
xor U10470 (N_10470,N_9258,N_9099);
xnor U10471 (N_10471,N_8322,N_9494);
or U10472 (N_10472,N_8000,N_9562);
and U10473 (N_10473,N_9741,N_9282);
nor U10474 (N_10474,N_8841,N_9245);
and U10475 (N_10475,N_8109,N_9458);
nand U10476 (N_10476,N_9660,N_9881);
nand U10477 (N_10477,N_8201,N_8474);
or U10478 (N_10478,N_8592,N_9558);
or U10479 (N_10479,N_8143,N_9203);
nand U10480 (N_10480,N_9623,N_8230);
nand U10481 (N_10481,N_8222,N_9312);
or U10482 (N_10482,N_9383,N_9933);
nor U10483 (N_10483,N_9517,N_8397);
and U10484 (N_10484,N_9096,N_9560);
or U10485 (N_10485,N_8787,N_8896);
or U10486 (N_10486,N_9957,N_8239);
nor U10487 (N_10487,N_8935,N_9162);
or U10488 (N_10488,N_9000,N_8476);
or U10489 (N_10489,N_9889,N_9552);
and U10490 (N_10490,N_9001,N_9761);
xor U10491 (N_10491,N_9567,N_8965);
xor U10492 (N_10492,N_9192,N_9188);
nor U10493 (N_10493,N_9718,N_9411);
and U10494 (N_10494,N_8852,N_9336);
xnor U10495 (N_10495,N_9206,N_9165);
or U10496 (N_10496,N_8387,N_9644);
xor U10497 (N_10497,N_8919,N_8472);
nand U10498 (N_10498,N_8490,N_8867);
xnor U10499 (N_10499,N_9855,N_8689);
nor U10500 (N_10500,N_8873,N_8059);
and U10501 (N_10501,N_8091,N_8773);
nand U10502 (N_10502,N_8237,N_9544);
or U10503 (N_10503,N_8421,N_9610);
nand U10504 (N_10504,N_9843,N_8939);
or U10505 (N_10505,N_8329,N_9086);
xnor U10506 (N_10506,N_9555,N_9370);
nor U10507 (N_10507,N_8186,N_9004);
nand U10508 (N_10508,N_9954,N_8272);
and U10509 (N_10509,N_8664,N_9721);
and U10510 (N_10510,N_8572,N_8316);
xor U10511 (N_10511,N_8757,N_9294);
and U10512 (N_10512,N_9405,N_9234);
or U10513 (N_10513,N_9321,N_9464);
xor U10514 (N_10514,N_8247,N_9524);
xor U10515 (N_10515,N_9598,N_8508);
nor U10516 (N_10516,N_8426,N_9917);
xor U10517 (N_10517,N_9189,N_8510);
xor U10518 (N_10518,N_9140,N_9404);
nor U10519 (N_10519,N_9492,N_9877);
nand U10520 (N_10520,N_9839,N_9455);
nand U10521 (N_10521,N_8915,N_8299);
nand U10522 (N_10522,N_8872,N_8351);
or U10523 (N_10523,N_9144,N_9922);
nor U10524 (N_10524,N_9337,N_8654);
xor U10525 (N_10525,N_9097,N_9295);
nor U10526 (N_10526,N_8521,N_9490);
nor U10527 (N_10527,N_8606,N_8943);
xnor U10528 (N_10528,N_9893,N_9424);
xnor U10529 (N_10529,N_8602,N_8985);
and U10530 (N_10530,N_8450,N_9532);
nor U10531 (N_10531,N_8540,N_9719);
xor U10532 (N_10532,N_9728,N_8077);
and U10533 (N_10533,N_9770,N_8496);
or U10534 (N_10534,N_9720,N_9974);
nor U10535 (N_10535,N_9483,N_9681);
and U10536 (N_10536,N_9110,N_9613);
nand U10537 (N_10537,N_9570,N_9095);
nand U10538 (N_10538,N_9987,N_9183);
and U10539 (N_10539,N_9009,N_9730);
and U10540 (N_10540,N_8023,N_9530);
and U10541 (N_10541,N_8422,N_9228);
xnor U10542 (N_10542,N_8823,N_8418);
xnor U10543 (N_10543,N_8184,N_8116);
nand U10544 (N_10544,N_8849,N_8026);
or U10545 (N_10545,N_9687,N_9430);
nand U10546 (N_10546,N_8561,N_9454);
nor U10547 (N_10547,N_8202,N_8808);
xor U10548 (N_10548,N_9418,N_9413);
xor U10549 (N_10549,N_9584,N_8703);
and U10550 (N_10550,N_8960,N_8219);
xor U10551 (N_10551,N_8618,N_9368);
or U10552 (N_10552,N_8467,N_8489);
or U10553 (N_10553,N_9682,N_8828);
or U10554 (N_10554,N_9087,N_8439);
xnor U10555 (N_10555,N_8717,N_9871);
xor U10556 (N_10556,N_8293,N_8482);
or U10557 (N_10557,N_9339,N_9463);
nor U10558 (N_10558,N_8928,N_8462);
and U10559 (N_10559,N_8585,N_9925);
nand U10560 (N_10560,N_8691,N_8402);
nor U10561 (N_10561,N_8213,N_8693);
nor U10562 (N_10562,N_9420,N_9746);
and U10563 (N_10563,N_8970,N_8656);
nand U10564 (N_10564,N_8576,N_8067);
and U10565 (N_10565,N_8519,N_8783);
nor U10566 (N_10566,N_8357,N_9503);
nor U10567 (N_10567,N_9797,N_8312);
and U10568 (N_10568,N_9173,N_9504);
or U10569 (N_10569,N_8171,N_8414);
or U10570 (N_10570,N_9057,N_9385);
and U10571 (N_10571,N_8321,N_9609);
and U10572 (N_10572,N_8241,N_9931);
and U10573 (N_10573,N_8307,N_9347);
nand U10574 (N_10574,N_8775,N_8281);
or U10575 (N_10575,N_8479,N_8048);
xnor U10576 (N_10576,N_9645,N_8214);
xor U10577 (N_10577,N_9710,N_8324);
nor U10578 (N_10578,N_9082,N_8627);
and U10579 (N_10579,N_9017,N_9423);
xnor U10580 (N_10580,N_8745,N_8952);
nand U10581 (N_10581,N_8337,N_9801);
or U10582 (N_10582,N_9130,N_8779);
xor U10583 (N_10583,N_8012,N_9055);
nor U10584 (N_10584,N_8242,N_9412);
xor U10585 (N_10585,N_8255,N_9852);
or U10586 (N_10586,N_8909,N_9892);
and U10587 (N_10587,N_8741,N_9864);
xnor U10588 (N_10588,N_8282,N_9067);
and U10589 (N_10589,N_8722,N_8856);
or U10590 (N_10590,N_9480,N_8579);
and U10591 (N_10591,N_8487,N_9891);
nor U10592 (N_10592,N_8437,N_9549);
nand U10593 (N_10593,N_9579,N_8335);
nor U10594 (N_10594,N_8850,N_9809);
nand U10595 (N_10595,N_9293,N_8532);
and U10596 (N_10596,N_8829,N_8020);
and U10597 (N_10597,N_8051,N_9484);
xnor U10598 (N_10598,N_8336,N_8558);
or U10599 (N_10599,N_9127,N_8203);
nor U10600 (N_10600,N_8846,N_8189);
and U10601 (N_10601,N_9273,N_8328);
and U10602 (N_10602,N_8930,N_9093);
or U10603 (N_10603,N_9172,N_8765);
or U10604 (N_10604,N_9042,N_9686);
nand U10605 (N_10605,N_8744,N_8557);
and U10606 (N_10606,N_8256,N_9156);
and U10607 (N_10607,N_8008,N_9210);
nor U10608 (N_10608,N_8343,N_8932);
xor U10609 (N_10609,N_9380,N_9618);
nor U10610 (N_10610,N_9960,N_9600);
or U10611 (N_10611,N_8223,N_8655);
nand U10612 (N_10612,N_8875,N_8551);
and U10613 (N_10613,N_8166,N_9232);
or U10614 (N_10614,N_8175,N_9507);
and U10615 (N_10615,N_9590,N_8076);
xnor U10616 (N_10616,N_8813,N_8671);
xor U10617 (N_10617,N_8403,N_8263);
xor U10618 (N_10618,N_9264,N_8724);
and U10619 (N_10619,N_8976,N_8347);
nand U10620 (N_10620,N_8061,N_8506);
xor U10621 (N_10621,N_8512,N_8533);
or U10622 (N_10622,N_9324,N_8731);
nor U10623 (N_10623,N_9114,N_9112);
xnor U10624 (N_10624,N_9593,N_9842);
nand U10625 (N_10625,N_8205,N_8317);
nor U10626 (N_10626,N_8866,N_8135);
nor U10627 (N_10627,N_9992,N_9688);
and U10628 (N_10628,N_9565,N_9262);
xor U10629 (N_10629,N_8505,N_8392);
nor U10630 (N_10630,N_8721,N_8986);
nor U10631 (N_10631,N_8288,N_9316);
nor U10632 (N_10632,N_8365,N_9798);
and U10633 (N_10633,N_8441,N_9178);
xor U10634 (N_10634,N_8360,N_8168);
nor U10635 (N_10635,N_9136,N_8834);
nand U10636 (N_10636,N_9617,N_9808);
nand U10637 (N_10637,N_8164,N_9829);
or U10638 (N_10638,N_9478,N_9731);
xor U10639 (N_10639,N_9285,N_9575);
xnor U10640 (N_10640,N_9665,N_8338);
nor U10641 (N_10641,N_8593,N_8543);
nand U10642 (N_10642,N_8782,N_9913);
nand U10643 (N_10643,N_9568,N_8114);
nor U10644 (N_10644,N_9914,N_9649);
and U10645 (N_10645,N_9419,N_9773);
xnor U10646 (N_10646,N_9676,N_8997);
nand U10647 (N_10647,N_9149,N_8180);
or U10648 (N_10648,N_8410,N_8898);
or U10649 (N_10649,N_9356,N_9664);
nand U10650 (N_10650,N_8470,N_8228);
or U10651 (N_10651,N_9821,N_8277);
xor U10652 (N_10652,N_9309,N_9386);
or U10653 (N_10653,N_8820,N_8821);
and U10654 (N_10654,N_9908,N_9190);
or U10655 (N_10655,N_8858,N_8874);
nand U10656 (N_10656,N_8888,N_9722);
and U10657 (N_10657,N_8492,N_9328);
and U10658 (N_10658,N_9231,N_8036);
xnor U10659 (N_10659,N_9572,N_9899);
nor U10660 (N_10660,N_8078,N_8894);
nor U10661 (N_10661,N_9577,N_8910);
and U10662 (N_10662,N_8763,N_9007);
nor U10663 (N_10663,N_8725,N_8802);
nand U10664 (N_10664,N_9834,N_8117);
or U10665 (N_10665,N_8553,N_8090);
and U10666 (N_10666,N_8954,N_8132);
xnor U10667 (N_10667,N_8897,N_8250);
xor U10668 (N_10668,N_9822,N_8125);
or U10669 (N_10669,N_8274,N_8525);
and U10670 (N_10670,N_9477,N_8756);
nand U10671 (N_10671,N_8375,N_8390);
or U10672 (N_10672,N_9563,N_8738);
nor U10673 (N_10673,N_9753,N_9622);
xor U10674 (N_10674,N_9679,N_8127);
nor U10675 (N_10675,N_8122,N_9174);
and U10676 (N_10676,N_8584,N_8516);
and U10677 (N_10677,N_9506,N_9540);
or U10678 (N_10678,N_8382,N_8517);
and U10679 (N_10679,N_8912,N_8167);
or U10680 (N_10680,N_9832,N_9539);
and U10681 (N_10681,N_9693,N_9197);
xor U10682 (N_10682,N_8465,N_9182);
xor U10683 (N_10683,N_9802,N_9260);
xnor U10684 (N_10684,N_8473,N_8600);
xor U10685 (N_10685,N_9755,N_9684);
nor U10686 (N_10686,N_9497,N_8598);
nand U10687 (N_10687,N_8301,N_8550);
nor U10688 (N_10688,N_9242,N_8009);
or U10689 (N_10689,N_8786,N_8947);
or U10690 (N_10690,N_8610,N_8636);
or U10691 (N_10691,N_8614,N_9612);
and U10692 (N_10692,N_8015,N_9869);
nand U10693 (N_10693,N_9302,N_8599);
xor U10694 (N_10694,N_8211,N_8883);
and U10695 (N_10695,N_9984,N_8996);
or U10696 (N_10696,N_9945,N_8224);
xor U10697 (N_10697,N_9121,N_9603);
and U10698 (N_10698,N_8038,N_8624);
nand U10699 (N_10699,N_9196,N_8941);
or U10700 (N_10700,N_8714,N_8795);
nor U10701 (N_10701,N_9934,N_9807);
and U10702 (N_10702,N_9045,N_9950);
xnor U10703 (N_10703,N_8659,N_8260);
nand U10704 (N_10704,N_9740,N_8249);
and U10705 (N_10705,N_8670,N_9642);
xor U10706 (N_10706,N_8760,N_9442);
nor U10707 (N_10707,N_8785,N_9030);
or U10708 (N_10708,N_9699,N_8457);
xnor U10709 (N_10709,N_8243,N_8793);
xor U10710 (N_10710,N_9481,N_9461);
or U10711 (N_10711,N_8886,N_8880);
or U10712 (N_10712,N_9143,N_9493);
xnor U10713 (N_10713,N_9379,N_9021);
nand U10714 (N_10714,N_9653,N_9081);
xor U10715 (N_10715,N_8037,N_8695);
nand U10716 (N_10716,N_9646,N_9508);
nand U10717 (N_10717,N_9704,N_8144);
and U10718 (N_10718,N_9215,N_9274);
nor U10719 (N_10719,N_9003,N_8349);
xor U10720 (N_10720,N_9450,N_9224);
nand U10721 (N_10721,N_8979,N_8847);
or U10722 (N_10722,N_9588,N_8541);
or U10723 (N_10723,N_9326,N_9760);
and U10724 (N_10724,N_9479,N_9955);
xnor U10725 (N_10725,N_8154,N_8701);
nor U10726 (N_10726,N_9138,N_9550);
xor U10727 (N_10727,N_8060,N_8953);
xor U10728 (N_10728,N_9103,N_9669);
and U10729 (N_10729,N_8739,N_8461);
nand U10730 (N_10730,N_9118,N_9689);
nand U10731 (N_10731,N_8933,N_8812);
xnor U10732 (N_10732,N_9820,N_9175);
nand U10733 (N_10733,N_8661,N_8311);
xor U10734 (N_10734,N_8955,N_9512);
or U10735 (N_10735,N_8407,N_9033);
nor U10736 (N_10736,N_9220,N_8626);
xnor U10737 (N_10737,N_8027,N_8346);
xor U10738 (N_10738,N_9592,N_8769);
xor U10739 (N_10739,N_9056,N_8504);
nand U10740 (N_10740,N_9299,N_9625);
xnor U10741 (N_10741,N_9358,N_8294);
nor U10742 (N_10742,N_8876,N_9936);
nand U10743 (N_10743,N_8777,N_9342);
xor U10744 (N_10744,N_8185,N_8663);
and U10745 (N_10745,N_9608,N_9122);
and U10746 (N_10746,N_9445,N_8803);
xnor U10747 (N_10747,N_9819,N_8030);
and U10748 (N_10748,N_9959,N_9031);
nor U10749 (N_10749,N_9831,N_8398);
nand U10750 (N_10750,N_8178,N_8869);
nand U10751 (N_10751,N_8069,N_8070);
xnor U10752 (N_10752,N_9186,N_8417);
and U10753 (N_10753,N_9918,N_9298);
and U10754 (N_10754,N_8622,N_9700);
nand U10755 (N_10755,N_8341,N_9453);
and U10756 (N_10756,N_8385,N_9811);
nand U10757 (N_10757,N_8792,N_9578);
nand U10758 (N_10758,N_9856,N_8524);
or U10759 (N_10759,N_8977,N_9619);
nor U10760 (N_10760,N_8198,N_9402);
xor U10761 (N_10761,N_8604,N_8697);
or U10762 (N_10762,N_9010,N_9566);
nand U10763 (N_10763,N_8235,N_9848);
nand U10764 (N_10764,N_8633,N_8816);
nand U10765 (N_10765,N_8033,N_9905);
or U10766 (N_10766,N_9878,N_8443);
and U10767 (N_10767,N_9732,N_9967);
nor U10768 (N_10768,N_8842,N_8396);
or U10769 (N_10769,N_9589,N_9225);
nor U10770 (N_10770,N_8179,N_9671);
or U10771 (N_10771,N_9833,N_8758);
nand U10772 (N_10772,N_9754,N_8589);
nand U10773 (N_10773,N_8811,N_8827);
and U10774 (N_10774,N_9582,N_9491);
nor U10775 (N_10775,N_9158,N_9774);
nand U10776 (N_10776,N_8531,N_8096);
xnor U10777 (N_10777,N_8993,N_8017);
and U10778 (N_10778,N_9941,N_9283);
and U10779 (N_10779,N_8617,N_8662);
nand U10780 (N_10780,N_8448,N_8290);
xnor U10781 (N_10781,N_8937,N_8607);
xnor U10782 (N_10782,N_8707,N_8978);
and U10783 (N_10783,N_9032,N_8675);
xor U10784 (N_10784,N_9511,N_8929);
and U10785 (N_10785,N_8353,N_8502);
nand U10786 (N_10786,N_9297,N_8619);
nor U10787 (N_10787,N_9763,N_9391);
nand U10788 (N_10788,N_9695,N_9876);
and U10789 (N_10789,N_8679,N_8565);
xor U10790 (N_10790,N_9213,N_8153);
xor U10791 (N_10791,N_8520,N_9910);
nor U10792 (N_10792,N_9926,N_8902);
and U10793 (N_10793,N_9782,N_8716);
nor U10794 (N_10794,N_8327,N_8372);
xor U10795 (N_10795,N_8147,N_8218);
and U10796 (N_10796,N_9426,N_9120);
and U10797 (N_10797,N_8204,N_8325);
or U10798 (N_10798,N_8923,N_9351);
xor U10799 (N_10799,N_8309,N_9862);
xnor U10800 (N_10800,N_8796,N_8261);
nand U10801 (N_10801,N_9486,N_9395);
xor U10802 (N_10802,N_8975,N_9556);
nor U10803 (N_10803,N_8463,N_9053);
and U10804 (N_10804,N_9341,N_9545);
nor U10805 (N_10805,N_9202,N_9673);
nand U10806 (N_10806,N_9449,N_8174);
or U10807 (N_10807,N_9444,N_8424);
nand U10808 (N_10808,N_9468,N_8304);
nor U10809 (N_10809,N_8234,N_8603);
or U10810 (N_10810,N_8771,N_8819);
or U10811 (N_10811,N_8690,N_8173);
nand U10812 (N_10812,N_9989,N_9407);
nor U10813 (N_10813,N_9961,N_8799);
xor U10814 (N_10814,N_9015,N_8111);
or U10815 (N_10815,N_8169,N_8233);
xnor U10816 (N_10816,N_9794,N_9076);
nor U10817 (N_10817,N_8057,N_9352);
xor U10818 (N_10818,N_9776,N_8588);
nor U10819 (N_10819,N_9803,N_8367);
or U10820 (N_10820,N_8107,N_9898);
nor U10821 (N_10821,N_9422,N_8660);
or U10822 (N_10822,N_9535,N_8648);
xnor U10823 (N_10823,N_8468,N_9758);
nand U10824 (N_10824,N_8578,N_9271);
nand U10825 (N_10825,N_9276,N_8053);
xnor U10826 (N_10826,N_8904,N_9457);
xnor U10827 (N_10827,N_8509,N_9287);
nand U10828 (N_10828,N_9838,N_9636);
and U10829 (N_10829,N_8814,N_8286);
and U10830 (N_10830,N_9920,N_8595);
or U10831 (N_10831,N_8253,N_9471);
and U10832 (N_10832,N_9151,N_9399);
xor U10833 (N_10833,N_9098,N_9965);
nand U10834 (N_10834,N_9949,N_9571);
and U10835 (N_10835,N_8093,N_9211);
nand U10836 (N_10836,N_9063,N_9226);
or U10837 (N_10837,N_8559,N_9727);
or U10838 (N_10838,N_8047,N_9988);
or U10839 (N_10839,N_8702,N_8907);
nor U10840 (N_10840,N_8708,N_8966);
xnor U10841 (N_10841,N_8623,N_8138);
nor U10842 (N_10842,N_8190,N_8086);
or U10843 (N_10843,N_9079,N_9564);
nand U10844 (N_10844,N_9134,N_9766);
nand U10845 (N_10845,N_9436,N_9308);
and U10846 (N_10846,N_9526,N_9751);
nor U10847 (N_10847,N_8634,N_9788);
and U10848 (N_10848,N_8776,N_8801);
nand U10849 (N_10849,N_9221,N_9909);
and U10850 (N_10850,N_8839,N_9737);
xor U10851 (N_10851,N_8522,N_9872);
and U10852 (N_10852,N_8055,N_9126);
and U10853 (N_10853,N_9795,N_8951);
and U10854 (N_10854,N_8208,N_8735);
xnor U10855 (N_10855,N_8097,N_9286);
or U10856 (N_10856,N_8081,N_9845);
or U10857 (N_10857,N_9252,N_9382);
nand U10858 (N_10858,N_9818,N_9020);
or U10859 (N_10859,N_9259,N_9697);
or U10860 (N_10860,N_9739,N_9208);
nor U10861 (N_10861,N_8905,N_9735);
nand U10862 (N_10862,N_8112,N_8789);
nor U10863 (N_10863,N_8727,N_8391);
nor U10864 (N_10864,N_8254,N_8195);
or U10865 (N_10865,N_9844,N_9034);
or U10866 (N_10866,N_9334,N_8772);
nor U10867 (N_10867,N_8563,N_8371);
nor U10868 (N_10868,N_8162,N_9065);
nor U10869 (N_10869,N_8022,N_8082);
nor U10870 (N_10870,N_8483,N_9771);
and U10871 (N_10871,N_9364,N_9836);
nor U10872 (N_10872,N_9813,N_8794);
or U10873 (N_10873,N_8052,N_8526);
nand U10874 (N_10874,N_8709,N_9135);
xor U10875 (N_10875,N_9906,N_8266);
nor U10876 (N_10876,N_9002,N_8105);
nor U10877 (N_10877,N_9476,N_9857);
xor U10878 (N_10878,N_8315,N_8914);
nand U10879 (N_10879,N_8999,N_9993);
nand U10880 (N_10880,N_9035,N_9139);
xnor U10881 (N_10881,N_9747,N_9024);
xor U10882 (N_10882,N_9799,N_8366);
and U10883 (N_10883,N_8158,N_9849);
or U10884 (N_10884,N_8104,N_8416);
xnor U10885 (N_10885,N_9702,N_8447);
nand U10886 (N_10886,N_8452,N_8005);
and U10887 (N_10887,N_8674,N_9345);
nand U10888 (N_10888,N_8206,N_8838);
nor U10889 (N_10889,N_8326,N_8810);
and U10890 (N_10890,N_9361,N_9981);
nand U10891 (N_10891,N_9073,N_8868);
nand U10892 (N_10892,N_9985,N_8571);
nand U10893 (N_10893,N_9432,N_8638);
xnor U10894 (N_10894,N_9062,N_9982);
xor U10895 (N_10895,N_9805,N_9496);
nor U10896 (N_10896,N_9254,N_8413);
nand U10897 (N_10897,N_9648,N_9650);
or U10898 (N_10898,N_8733,N_9350);
xnor U10899 (N_10899,N_9488,N_9300);
or U10900 (N_10900,N_8103,N_9137);
or U10901 (N_10901,N_9141,N_9071);
nand U10902 (N_10902,N_8045,N_8238);
xnor U10903 (N_10903,N_8940,N_8244);
xnor U10904 (N_10904,N_8800,N_9128);
nor U10905 (N_10905,N_9932,N_8991);
or U10906 (N_10906,N_8957,N_8556);
and U10907 (N_10907,N_8161,N_8948);
xor U10908 (N_10908,N_8393,N_8566);
or U10909 (N_10909,N_8751,N_8040);
nand U10910 (N_10910,N_9179,N_9990);
xnor U10911 (N_10911,N_9859,N_8412);
nand U10912 (N_10912,N_8683,N_8865);
or U10913 (N_10913,N_8764,N_9397);
xnor U10914 (N_10914,N_8692,N_9470);
and U10915 (N_10915,N_8394,N_9742);
nand U10916 (N_10916,N_8938,N_8825);
or U10917 (N_10917,N_8569,N_8831);
nand U10918 (N_10918,N_9978,N_9627);
or U10919 (N_10919,N_8778,N_8246);
nor U10920 (N_10920,N_9349,N_9246);
nand U10921 (N_10921,N_9270,N_8003);
xor U10922 (N_10922,N_8944,N_9998);
xnor U10923 (N_10923,N_8220,N_9304);
nor U10924 (N_10924,N_8980,N_8011);
xnor U10925 (N_10925,N_9275,N_8723);
nor U10926 (N_10926,N_9971,N_9025);
xor U10927 (N_10927,N_9554,N_8355);
nand U10928 (N_10928,N_8485,N_8890);
nor U10929 (N_10929,N_8596,N_9958);
or U10930 (N_10930,N_9233,N_9505);
nand U10931 (N_10931,N_9585,N_9205);
xnor U10932 (N_10932,N_8861,N_8582);
nand U10933 (N_10933,N_8781,N_8499);
nand U10934 (N_10934,N_9333,N_8575);
and U10935 (N_10935,N_9389,N_9362);
and U10936 (N_10936,N_9415,N_8137);
nand U10937 (N_10937,N_9396,N_8908);
or U10938 (N_10938,N_9940,N_8406);
nand U10939 (N_10939,N_9900,N_9882);
and U10940 (N_10940,N_9077,N_8704);
or U10941 (N_10941,N_8639,N_8630);
and U10942 (N_10942,N_8646,N_8740);
and U10943 (N_10943,N_8736,N_9597);
xor U10944 (N_10944,N_9416,N_9229);
and U10945 (N_10945,N_8631,N_9443);
nand U10946 (N_10946,N_9201,N_9806);
xnor U10947 (N_10947,N_9446,N_8240);
and U10948 (N_10948,N_9400,N_9791);
nand U10949 (N_10949,N_8963,N_8580);
and U10950 (N_10950,N_9039,N_8835);
nor U10951 (N_10951,N_9239,N_9630);
nand U10952 (N_10952,N_8720,N_8199);
nand U10953 (N_10953,N_8227,N_9346);
and U10954 (N_10954,N_8370,N_9826);
and U10955 (N_10955,N_8425,N_9329);
nand U10956 (N_10956,N_9296,N_8043);
nand U10957 (N_10957,N_8306,N_8959);
nand U10958 (N_10958,N_8054,N_9058);
nor U10959 (N_10959,N_8666,N_8384);
or U10960 (N_10960,N_8591,N_8480);
nand U10961 (N_10961,N_8409,N_8339);
and U10962 (N_10962,N_9948,N_8855);
nand U10963 (N_10963,N_9193,N_8562);
or U10964 (N_10964,N_8345,N_9652);
nor U10965 (N_10965,N_8378,N_8248);
nor U10966 (N_10966,N_8475,N_8613);
nor U10967 (N_10967,N_8577,N_9325);
xor U10968 (N_10968,N_8523,N_8685);
nor U10969 (N_10969,N_9904,N_9536);
xor U10970 (N_10970,N_9061,N_8319);
nor U10971 (N_10971,N_9523,N_8535);
nand U10972 (N_10972,N_8386,N_8752);
xor U10973 (N_10973,N_8065,N_9830);
xnor U10974 (N_10974,N_9670,N_8101);
nor U10975 (N_10975,N_9013,N_9005);
nor U10976 (N_10976,N_8018,N_9531);
or U10977 (N_10977,N_8922,N_9633);
and U10978 (N_10978,N_9715,N_8044);
nand U10979 (N_10979,N_8305,N_9738);
and U10980 (N_10980,N_9615,N_8415);
nand U10981 (N_10981,N_9322,N_8641);
nand U10982 (N_10982,N_8554,N_8911);
and U10983 (N_10983,N_9657,N_8981);
xnor U10984 (N_10984,N_9041,N_9935);
nor U10985 (N_10985,N_8788,N_8432);
xor U10986 (N_10986,N_9658,N_9070);
and U10987 (N_10987,N_8766,N_9667);
and U10988 (N_10988,N_9607,N_8871);
or U10989 (N_10989,N_8212,N_8643);
nand U10990 (N_10990,N_8408,N_9703);
or U10991 (N_10991,N_8903,N_9250);
nand U10992 (N_10992,N_9256,N_9850);
or U10993 (N_10993,N_9105,N_9390);
nand U10994 (N_10994,N_8870,N_9363);
xor U10995 (N_10995,N_8110,N_8291);
or U10996 (N_10996,N_9725,N_9365);
nor U10997 (N_10997,N_8895,N_9381);
or U10998 (N_10998,N_8676,N_9786);
or U10999 (N_10999,N_9701,N_8806);
or U11000 (N_11000,N_9310,N_9998);
nand U11001 (N_11001,N_9436,N_8811);
and U11002 (N_11002,N_8817,N_8622);
and U11003 (N_11003,N_9726,N_8049);
or U11004 (N_11004,N_9972,N_9165);
xnor U11005 (N_11005,N_9838,N_8942);
nand U11006 (N_11006,N_9389,N_8811);
and U11007 (N_11007,N_9424,N_8144);
and U11008 (N_11008,N_9738,N_9154);
xnor U11009 (N_11009,N_9606,N_8515);
nand U11010 (N_11010,N_8066,N_9311);
and U11011 (N_11011,N_8121,N_8234);
nand U11012 (N_11012,N_8670,N_8486);
nor U11013 (N_11013,N_9245,N_9757);
xor U11014 (N_11014,N_9180,N_8471);
nor U11015 (N_11015,N_8398,N_9052);
xor U11016 (N_11016,N_9034,N_8191);
or U11017 (N_11017,N_8681,N_9673);
or U11018 (N_11018,N_9828,N_8730);
nand U11019 (N_11019,N_9584,N_9035);
xor U11020 (N_11020,N_8093,N_9137);
and U11021 (N_11021,N_8518,N_8274);
and U11022 (N_11022,N_9041,N_8925);
nor U11023 (N_11023,N_9048,N_9312);
and U11024 (N_11024,N_8938,N_9753);
and U11025 (N_11025,N_8470,N_9993);
or U11026 (N_11026,N_9690,N_9599);
nor U11027 (N_11027,N_8512,N_9651);
and U11028 (N_11028,N_9921,N_9854);
or U11029 (N_11029,N_9054,N_9826);
or U11030 (N_11030,N_8248,N_8739);
or U11031 (N_11031,N_9917,N_8589);
and U11032 (N_11032,N_9297,N_8225);
xnor U11033 (N_11033,N_9558,N_9477);
nand U11034 (N_11034,N_9831,N_8095);
xor U11035 (N_11035,N_9310,N_9892);
nand U11036 (N_11036,N_9361,N_9719);
nand U11037 (N_11037,N_9936,N_9402);
nor U11038 (N_11038,N_8081,N_8580);
nor U11039 (N_11039,N_8604,N_9013);
or U11040 (N_11040,N_9394,N_9360);
xnor U11041 (N_11041,N_8311,N_9713);
nand U11042 (N_11042,N_8865,N_9509);
and U11043 (N_11043,N_8456,N_8160);
nor U11044 (N_11044,N_8481,N_8109);
nand U11045 (N_11045,N_9409,N_8387);
nand U11046 (N_11046,N_8185,N_9753);
nor U11047 (N_11047,N_9932,N_9885);
nor U11048 (N_11048,N_8765,N_9195);
xor U11049 (N_11049,N_9351,N_8286);
nor U11050 (N_11050,N_8754,N_8076);
xnor U11051 (N_11051,N_9396,N_8932);
nor U11052 (N_11052,N_8868,N_8413);
and U11053 (N_11053,N_8432,N_8700);
and U11054 (N_11054,N_9179,N_9009);
xor U11055 (N_11055,N_8273,N_8290);
xnor U11056 (N_11056,N_8485,N_9987);
nand U11057 (N_11057,N_9998,N_8226);
or U11058 (N_11058,N_9663,N_8705);
nor U11059 (N_11059,N_8870,N_9646);
nand U11060 (N_11060,N_8499,N_8676);
xor U11061 (N_11061,N_8659,N_9037);
and U11062 (N_11062,N_9383,N_8281);
or U11063 (N_11063,N_8109,N_8140);
xnor U11064 (N_11064,N_8899,N_8772);
xnor U11065 (N_11065,N_8996,N_8780);
nand U11066 (N_11066,N_8356,N_9839);
nor U11067 (N_11067,N_9290,N_9264);
or U11068 (N_11068,N_8367,N_9760);
or U11069 (N_11069,N_9420,N_8698);
xor U11070 (N_11070,N_9401,N_9162);
and U11071 (N_11071,N_8078,N_8730);
nor U11072 (N_11072,N_9109,N_9542);
or U11073 (N_11073,N_8841,N_9450);
nand U11074 (N_11074,N_9490,N_8148);
xor U11075 (N_11075,N_8720,N_9225);
or U11076 (N_11076,N_8997,N_9760);
xor U11077 (N_11077,N_8635,N_8378);
and U11078 (N_11078,N_9006,N_8641);
or U11079 (N_11079,N_8066,N_9433);
nor U11080 (N_11080,N_9562,N_9471);
xnor U11081 (N_11081,N_8812,N_9307);
or U11082 (N_11082,N_8997,N_9865);
xor U11083 (N_11083,N_9295,N_9682);
and U11084 (N_11084,N_9933,N_9848);
xnor U11085 (N_11085,N_8928,N_8785);
and U11086 (N_11086,N_8198,N_8330);
or U11087 (N_11087,N_8395,N_8100);
nand U11088 (N_11088,N_9665,N_9291);
and U11089 (N_11089,N_8643,N_9882);
and U11090 (N_11090,N_9511,N_9201);
nand U11091 (N_11091,N_9893,N_9193);
xor U11092 (N_11092,N_8913,N_9281);
or U11093 (N_11093,N_9204,N_9873);
nand U11094 (N_11094,N_8465,N_8765);
nand U11095 (N_11095,N_9743,N_9699);
and U11096 (N_11096,N_8381,N_8231);
or U11097 (N_11097,N_9199,N_8635);
nand U11098 (N_11098,N_9554,N_9714);
or U11099 (N_11099,N_9321,N_8905);
or U11100 (N_11100,N_8128,N_8908);
or U11101 (N_11101,N_8532,N_8137);
and U11102 (N_11102,N_8114,N_9935);
and U11103 (N_11103,N_9310,N_9423);
and U11104 (N_11104,N_8618,N_8540);
xnor U11105 (N_11105,N_9761,N_8152);
and U11106 (N_11106,N_9479,N_9114);
nor U11107 (N_11107,N_9352,N_9823);
nor U11108 (N_11108,N_9106,N_8715);
or U11109 (N_11109,N_8855,N_9956);
nand U11110 (N_11110,N_8963,N_8265);
and U11111 (N_11111,N_9848,N_8434);
nor U11112 (N_11112,N_8753,N_8856);
xor U11113 (N_11113,N_8976,N_9338);
or U11114 (N_11114,N_9725,N_9126);
and U11115 (N_11115,N_8442,N_9305);
xnor U11116 (N_11116,N_8203,N_8787);
or U11117 (N_11117,N_8638,N_8508);
nand U11118 (N_11118,N_9427,N_9371);
nor U11119 (N_11119,N_8172,N_9752);
or U11120 (N_11120,N_9892,N_9544);
nand U11121 (N_11121,N_8936,N_8288);
and U11122 (N_11122,N_8300,N_8564);
and U11123 (N_11123,N_9046,N_9275);
nor U11124 (N_11124,N_8565,N_9612);
nand U11125 (N_11125,N_9500,N_8425);
nand U11126 (N_11126,N_8578,N_9256);
and U11127 (N_11127,N_8404,N_8636);
and U11128 (N_11128,N_9602,N_9800);
and U11129 (N_11129,N_8459,N_8933);
or U11130 (N_11130,N_8421,N_9227);
nor U11131 (N_11131,N_8002,N_8521);
nor U11132 (N_11132,N_8030,N_9447);
nand U11133 (N_11133,N_8546,N_9724);
and U11134 (N_11134,N_9447,N_9538);
xnor U11135 (N_11135,N_9444,N_8854);
xnor U11136 (N_11136,N_9071,N_9344);
and U11137 (N_11137,N_9216,N_8516);
xnor U11138 (N_11138,N_9992,N_8279);
nor U11139 (N_11139,N_8769,N_9087);
or U11140 (N_11140,N_8901,N_8566);
nand U11141 (N_11141,N_9270,N_8755);
nand U11142 (N_11142,N_9843,N_9508);
nand U11143 (N_11143,N_8157,N_9368);
nand U11144 (N_11144,N_9373,N_9083);
nand U11145 (N_11145,N_9112,N_9741);
nor U11146 (N_11146,N_8814,N_9202);
nand U11147 (N_11147,N_9413,N_8933);
xnor U11148 (N_11148,N_8465,N_8861);
xor U11149 (N_11149,N_8349,N_9995);
nand U11150 (N_11150,N_9680,N_8804);
nor U11151 (N_11151,N_8045,N_8885);
or U11152 (N_11152,N_9728,N_9760);
nor U11153 (N_11153,N_9645,N_9111);
or U11154 (N_11154,N_8880,N_8095);
xor U11155 (N_11155,N_9080,N_9337);
xor U11156 (N_11156,N_8831,N_8672);
nand U11157 (N_11157,N_9684,N_8302);
or U11158 (N_11158,N_9381,N_8128);
nor U11159 (N_11159,N_8448,N_8791);
nor U11160 (N_11160,N_9162,N_9927);
or U11161 (N_11161,N_8977,N_8290);
and U11162 (N_11162,N_9415,N_8544);
and U11163 (N_11163,N_8862,N_9630);
and U11164 (N_11164,N_9827,N_8618);
nand U11165 (N_11165,N_8086,N_9001);
and U11166 (N_11166,N_8090,N_9790);
nor U11167 (N_11167,N_9469,N_9117);
and U11168 (N_11168,N_9248,N_9296);
and U11169 (N_11169,N_8760,N_9325);
and U11170 (N_11170,N_8381,N_8590);
xnor U11171 (N_11171,N_9976,N_8536);
or U11172 (N_11172,N_9456,N_9827);
and U11173 (N_11173,N_8977,N_9837);
xnor U11174 (N_11174,N_8998,N_8702);
xnor U11175 (N_11175,N_8552,N_8752);
xnor U11176 (N_11176,N_8629,N_9169);
or U11177 (N_11177,N_8043,N_9526);
and U11178 (N_11178,N_9273,N_9571);
nor U11179 (N_11179,N_8199,N_8894);
or U11180 (N_11180,N_8486,N_8317);
xor U11181 (N_11181,N_9034,N_9619);
nand U11182 (N_11182,N_9998,N_8612);
nor U11183 (N_11183,N_9788,N_8088);
nor U11184 (N_11184,N_9637,N_9383);
nor U11185 (N_11185,N_8778,N_8925);
and U11186 (N_11186,N_9134,N_9822);
or U11187 (N_11187,N_8489,N_9981);
and U11188 (N_11188,N_9484,N_8863);
or U11189 (N_11189,N_8984,N_9826);
nor U11190 (N_11190,N_9133,N_8521);
nand U11191 (N_11191,N_8482,N_8540);
and U11192 (N_11192,N_8720,N_9809);
xor U11193 (N_11193,N_8722,N_9549);
nor U11194 (N_11194,N_9999,N_8564);
nand U11195 (N_11195,N_9558,N_9546);
nand U11196 (N_11196,N_9444,N_8567);
nor U11197 (N_11197,N_9464,N_8376);
or U11198 (N_11198,N_9423,N_9676);
and U11199 (N_11199,N_9614,N_8465);
xnor U11200 (N_11200,N_8346,N_8494);
or U11201 (N_11201,N_8372,N_9168);
or U11202 (N_11202,N_8360,N_9655);
and U11203 (N_11203,N_9484,N_9312);
nor U11204 (N_11204,N_8098,N_8087);
nand U11205 (N_11205,N_9283,N_9572);
nor U11206 (N_11206,N_9292,N_9304);
nor U11207 (N_11207,N_9176,N_8539);
or U11208 (N_11208,N_8850,N_8466);
and U11209 (N_11209,N_9023,N_8205);
nand U11210 (N_11210,N_9005,N_9783);
nor U11211 (N_11211,N_9025,N_8264);
nand U11212 (N_11212,N_8442,N_9513);
xnor U11213 (N_11213,N_9803,N_9194);
and U11214 (N_11214,N_9243,N_8499);
nor U11215 (N_11215,N_9897,N_9707);
nand U11216 (N_11216,N_9385,N_9722);
and U11217 (N_11217,N_8521,N_8594);
or U11218 (N_11218,N_8676,N_8627);
or U11219 (N_11219,N_9035,N_9905);
nand U11220 (N_11220,N_8545,N_8073);
xor U11221 (N_11221,N_8182,N_8521);
nor U11222 (N_11222,N_9735,N_8606);
or U11223 (N_11223,N_9559,N_8946);
xnor U11224 (N_11224,N_8306,N_8617);
nor U11225 (N_11225,N_9009,N_9361);
nor U11226 (N_11226,N_8908,N_8941);
or U11227 (N_11227,N_8775,N_9543);
and U11228 (N_11228,N_9563,N_8028);
nor U11229 (N_11229,N_9825,N_8743);
nand U11230 (N_11230,N_8135,N_8188);
nand U11231 (N_11231,N_8346,N_8871);
nand U11232 (N_11232,N_8761,N_8647);
nor U11233 (N_11233,N_9796,N_9860);
nand U11234 (N_11234,N_9985,N_9355);
and U11235 (N_11235,N_8404,N_8820);
xnor U11236 (N_11236,N_8140,N_9268);
xnor U11237 (N_11237,N_8150,N_9119);
or U11238 (N_11238,N_9820,N_8738);
and U11239 (N_11239,N_8161,N_8850);
nor U11240 (N_11240,N_9988,N_9628);
xor U11241 (N_11241,N_9234,N_8159);
nor U11242 (N_11242,N_9524,N_9408);
and U11243 (N_11243,N_9936,N_9016);
nor U11244 (N_11244,N_8329,N_9769);
nor U11245 (N_11245,N_8396,N_8706);
nor U11246 (N_11246,N_9829,N_8062);
nand U11247 (N_11247,N_9254,N_8689);
nand U11248 (N_11248,N_8490,N_8033);
nor U11249 (N_11249,N_9477,N_9161);
nand U11250 (N_11250,N_9038,N_9411);
nor U11251 (N_11251,N_9339,N_8197);
xnor U11252 (N_11252,N_8190,N_8028);
nand U11253 (N_11253,N_9617,N_9350);
and U11254 (N_11254,N_9668,N_9741);
or U11255 (N_11255,N_8950,N_8091);
nor U11256 (N_11256,N_9805,N_8289);
or U11257 (N_11257,N_8720,N_8366);
xnor U11258 (N_11258,N_9878,N_9632);
and U11259 (N_11259,N_9574,N_9005);
nor U11260 (N_11260,N_9693,N_9289);
or U11261 (N_11261,N_8163,N_9637);
nor U11262 (N_11262,N_8444,N_9170);
xnor U11263 (N_11263,N_8401,N_8855);
or U11264 (N_11264,N_8242,N_8014);
nor U11265 (N_11265,N_8743,N_9493);
xnor U11266 (N_11266,N_8923,N_8920);
and U11267 (N_11267,N_9809,N_8383);
nand U11268 (N_11268,N_9090,N_9933);
or U11269 (N_11269,N_9433,N_9770);
xnor U11270 (N_11270,N_8311,N_8959);
or U11271 (N_11271,N_9082,N_9506);
nor U11272 (N_11272,N_9761,N_9402);
and U11273 (N_11273,N_8048,N_9892);
nor U11274 (N_11274,N_8301,N_8817);
nand U11275 (N_11275,N_8152,N_8172);
or U11276 (N_11276,N_8962,N_9697);
nand U11277 (N_11277,N_9148,N_9435);
or U11278 (N_11278,N_8055,N_8448);
and U11279 (N_11279,N_9178,N_8836);
or U11280 (N_11280,N_8342,N_8265);
nand U11281 (N_11281,N_8792,N_8038);
nor U11282 (N_11282,N_9864,N_8869);
nand U11283 (N_11283,N_8861,N_8004);
and U11284 (N_11284,N_8880,N_9349);
and U11285 (N_11285,N_8672,N_9972);
nor U11286 (N_11286,N_9530,N_9161);
xor U11287 (N_11287,N_9983,N_9038);
or U11288 (N_11288,N_8429,N_8037);
or U11289 (N_11289,N_9349,N_9556);
or U11290 (N_11290,N_8084,N_8456);
nor U11291 (N_11291,N_8953,N_9130);
nor U11292 (N_11292,N_8151,N_8631);
nand U11293 (N_11293,N_9206,N_9025);
and U11294 (N_11294,N_9700,N_8583);
nand U11295 (N_11295,N_8212,N_8360);
or U11296 (N_11296,N_9386,N_9137);
or U11297 (N_11297,N_8739,N_9548);
or U11298 (N_11298,N_9847,N_8014);
and U11299 (N_11299,N_8545,N_8972);
nor U11300 (N_11300,N_8633,N_8738);
nor U11301 (N_11301,N_8849,N_9051);
xor U11302 (N_11302,N_8410,N_9867);
nand U11303 (N_11303,N_9669,N_9310);
and U11304 (N_11304,N_8251,N_9823);
nor U11305 (N_11305,N_8368,N_9761);
nand U11306 (N_11306,N_9161,N_9754);
xnor U11307 (N_11307,N_8255,N_9229);
or U11308 (N_11308,N_9516,N_9255);
xnor U11309 (N_11309,N_9421,N_9904);
nor U11310 (N_11310,N_9932,N_8068);
or U11311 (N_11311,N_8984,N_8735);
or U11312 (N_11312,N_8146,N_8065);
xnor U11313 (N_11313,N_8727,N_9392);
nor U11314 (N_11314,N_8021,N_8797);
nor U11315 (N_11315,N_8212,N_8118);
xnor U11316 (N_11316,N_8383,N_8628);
or U11317 (N_11317,N_8201,N_9174);
or U11318 (N_11318,N_8766,N_9006);
xnor U11319 (N_11319,N_9171,N_8312);
nand U11320 (N_11320,N_8393,N_9333);
xor U11321 (N_11321,N_8205,N_9314);
nand U11322 (N_11322,N_9857,N_9145);
nand U11323 (N_11323,N_8551,N_9989);
or U11324 (N_11324,N_9594,N_8394);
xnor U11325 (N_11325,N_9603,N_9621);
nand U11326 (N_11326,N_9094,N_8940);
and U11327 (N_11327,N_9087,N_9889);
nand U11328 (N_11328,N_8130,N_9961);
or U11329 (N_11329,N_8118,N_9523);
or U11330 (N_11330,N_8493,N_8142);
and U11331 (N_11331,N_8421,N_8208);
nand U11332 (N_11332,N_8476,N_8576);
nor U11333 (N_11333,N_9541,N_9009);
nor U11334 (N_11334,N_9718,N_8712);
xnor U11335 (N_11335,N_9454,N_8053);
xor U11336 (N_11336,N_8654,N_9184);
or U11337 (N_11337,N_8015,N_8362);
and U11338 (N_11338,N_8114,N_8864);
or U11339 (N_11339,N_9315,N_8844);
and U11340 (N_11340,N_9735,N_9803);
nand U11341 (N_11341,N_8525,N_8569);
xnor U11342 (N_11342,N_8689,N_9448);
nand U11343 (N_11343,N_8517,N_9377);
or U11344 (N_11344,N_8931,N_8210);
xor U11345 (N_11345,N_9607,N_8362);
nand U11346 (N_11346,N_8434,N_8454);
xnor U11347 (N_11347,N_8735,N_9845);
or U11348 (N_11348,N_8920,N_9584);
xnor U11349 (N_11349,N_8616,N_8964);
nor U11350 (N_11350,N_8062,N_9788);
xnor U11351 (N_11351,N_8094,N_8718);
xnor U11352 (N_11352,N_9648,N_8103);
and U11353 (N_11353,N_9512,N_9110);
nor U11354 (N_11354,N_9464,N_9448);
nor U11355 (N_11355,N_8493,N_9257);
xnor U11356 (N_11356,N_9094,N_8583);
nand U11357 (N_11357,N_9260,N_9791);
or U11358 (N_11358,N_9237,N_9008);
nand U11359 (N_11359,N_9388,N_8165);
nand U11360 (N_11360,N_9497,N_9835);
or U11361 (N_11361,N_9007,N_9806);
nand U11362 (N_11362,N_8867,N_8495);
nor U11363 (N_11363,N_8309,N_9212);
nand U11364 (N_11364,N_9664,N_8858);
nand U11365 (N_11365,N_9911,N_8393);
nor U11366 (N_11366,N_9040,N_9034);
or U11367 (N_11367,N_8349,N_8360);
nand U11368 (N_11368,N_8557,N_9771);
xnor U11369 (N_11369,N_9894,N_9571);
or U11370 (N_11370,N_8291,N_8734);
xor U11371 (N_11371,N_9102,N_8480);
xor U11372 (N_11372,N_8223,N_9283);
xnor U11373 (N_11373,N_8667,N_8457);
and U11374 (N_11374,N_8758,N_9031);
and U11375 (N_11375,N_9059,N_8751);
or U11376 (N_11376,N_9739,N_8578);
nor U11377 (N_11377,N_8851,N_8951);
nor U11378 (N_11378,N_8938,N_8739);
nand U11379 (N_11379,N_8712,N_9758);
nor U11380 (N_11380,N_9373,N_9706);
xnor U11381 (N_11381,N_9321,N_8400);
nand U11382 (N_11382,N_9516,N_9215);
xor U11383 (N_11383,N_8544,N_8646);
or U11384 (N_11384,N_8794,N_9947);
nand U11385 (N_11385,N_9642,N_8794);
or U11386 (N_11386,N_8952,N_9506);
xor U11387 (N_11387,N_9528,N_8983);
nand U11388 (N_11388,N_8337,N_8682);
xnor U11389 (N_11389,N_9644,N_9373);
nor U11390 (N_11390,N_9668,N_8324);
or U11391 (N_11391,N_9645,N_8247);
xor U11392 (N_11392,N_9295,N_9986);
and U11393 (N_11393,N_8991,N_8827);
nor U11394 (N_11394,N_9751,N_8964);
xnor U11395 (N_11395,N_9926,N_9562);
or U11396 (N_11396,N_8397,N_9705);
or U11397 (N_11397,N_8607,N_8782);
xnor U11398 (N_11398,N_8436,N_8375);
nand U11399 (N_11399,N_9065,N_9791);
xnor U11400 (N_11400,N_9319,N_8316);
xnor U11401 (N_11401,N_8375,N_8050);
nor U11402 (N_11402,N_9897,N_9708);
nand U11403 (N_11403,N_8574,N_9193);
xor U11404 (N_11404,N_9389,N_9929);
and U11405 (N_11405,N_8507,N_8350);
nor U11406 (N_11406,N_9699,N_8496);
nor U11407 (N_11407,N_8810,N_8733);
or U11408 (N_11408,N_8052,N_9214);
xnor U11409 (N_11409,N_9796,N_8524);
nor U11410 (N_11410,N_8297,N_9503);
nand U11411 (N_11411,N_9823,N_9905);
and U11412 (N_11412,N_9304,N_9016);
nand U11413 (N_11413,N_8718,N_8833);
nand U11414 (N_11414,N_8851,N_9019);
or U11415 (N_11415,N_8548,N_9255);
xor U11416 (N_11416,N_9324,N_8564);
nand U11417 (N_11417,N_8985,N_9732);
and U11418 (N_11418,N_9088,N_8941);
and U11419 (N_11419,N_9883,N_9824);
xnor U11420 (N_11420,N_8689,N_9816);
nand U11421 (N_11421,N_8017,N_9143);
and U11422 (N_11422,N_8385,N_8388);
or U11423 (N_11423,N_8114,N_8808);
and U11424 (N_11424,N_8484,N_8957);
nand U11425 (N_11425,N_8810,N_8879);
or U11426 (N_11426,N_9402,N_9129);
and U11427 (N_11427,N_9786,N_9553);
nor U11428 (N_11428,N_9874,N_9353);
or U11429 (N_11429,N_8661,N_9232);
nand U11430 (N_11430,N_8799,N_9512);
nand U11431 (N_11431,N_9879,N_9616);
nand U11432 (N_11432,N_8149,N_8058);
nor U11433 (N_11433,N_8361,N_8897);
xnor U11434 (N_11434,N_9658,N_8023);
nor U11435 (N_11435,N_8291,N_9991);
nor U11436 (N_11436,N_8682,N_8549);
and U11437 (N_11437,N_8724,N_9061);
and U11438 (N_11438,N_8159,N_9577);
xor U11439 (N_11439,N_8710,N_9992);
nand U11440 (N_11440,N_9388,N_9914);
nor U11441 (N_11441,N_9632,N_8616);
and U11442 (N_11442,N_8165,N_9243);
and U11443 (N_11443,N_8286,N_9855);
xor U11444 (N_11444,N_9955,N_8512);
or U11445 (N_11445,N_8006,N_8019);
and U11446 (N_11446,N_9496,N_8337);
xor U11447 (N_11447,N_8427,N_8684);
or U11448 (N_11448,N_9497,N_9793);
nor U11449 (N_11449,N_9387,N_9863);
xnor U11450 (N_11450,N_8807,N_9400);
nor U11451 (N_11451,N_8966,N_9131);
nor U11452 (N_11452,N_8475,N_9216);
and U11453 (N_11453,N_8116,N_9099);
nor U11454 (N_11454,N_9394,N_8136);
or U11455 (N_11455,N_9114,N_9765);
xor U11456 (N_11456,N_8179,N_9726);
nand U11457 (N_11457,N_8152,N_9958);
and U11458 (N_11458,N_9076,N_9655);
or U11459 (N_11459,N_8085,N_8099);
xnor U11460 (N_11460,N_8438,N_9659);
nand U11461 (N_11461,N_8803,N_9442);
or U11462 (N_11462,N_9275,N_8125);
nand U11463 (N_11463,N_8845,N_8025);
or U11464 (N_11464,N_8599,N_9463);
or U11465 (N_11465,N_9065,N_8864);
and U11466 (N_11466,N_9643,N_8162);
nand U11467 (N_11467,N_8925,N_9644);
and U11468 (N_11468,N_9719,N_9812);
nand U11469 (N_11469,N_9680,N_9967);
nor U11470 (N_11470,N_8603,N_9902);
xor U11471 (N_11471,N_9645,N_8634);
xnor U11472 (N_11472,N_8161,N_9749);
and U11473 (N_11473,N_9093,N_9771);
nand U11474 (N_11474,N_8921,N_9997);
xor U11475 (N_11475,N_8900,N_9412);
and U11476 (N_11476,N_9566,N_8198);
or U11477 (N_11477,N_9492,N_8118);
xor U11478 (N_11478,N_9634,N_9563);
nor U11479 (N_11479,N_9861,N_8872);
nor U11480 (N_11480,N_9030,N_9995);
xor U11481 (N_11481,N_8198,N_8502);
or U11482 (N_11482,N_8689,N_9712);
nand U11483 (N_11483,N_8262,N_9837);
nand U11484 (N_11484,N_9756,N_9638);
and U11485 (N_11485,N_9326,N_9626);
xor U11486 (N_11486,N_9062,N_8361);
or U11487 (N_11487,N_8577,N_9406);
nor U11488 (N_11488,N_9446,N_8845);
nor U11489 (N_11489,N_8248,N_9025);
and U11490 (N_11490,N_9561,N_8868);
nand U11491 (N_11491,N_9687,N_9689);
xnor U11492 (N_11492,N_9045,N_8803);
xnor U11493 (N_11493,N_9709,N_8380);
xnor U11494 (N_11494,N_8912,N_8965);
and U11495 (N_11495,N_9452,N_8046);
nor U11496 (N_11496,N_9003,N_8187);
nor U11497 (N_11497,N_9395,N_9751);
and U11498 (N_11498,N_8792,N_9072);
xor U11499 (N_11499,N_9159,N_9168);
or U11500 (N_11500,N_8097,N_8275);
xnor U11501 (N_11501,N_9981,N_8307);
xor U11502 (N_11502,N_9065,N_8773);
xnor U11503 (N_11503,N_9817,N_8971);
or U11504 (N_11504,N_8304,N_8479);
or U11505 (N_11505,N_8545,N_9516);
and U11506 (N_11506,N_8437,N_8804);
nor U11507 (N_11507,N_8749,N_8804);
nor U11508 (N_11508,N_8280,N_8594);
or U11509 (N_11509,N_9799,N_8223);
nor U11510 (N_11510,N_8953,N_8010);
xor U11511 (N_11511,N_9216,N_8128);
nand U11512 (N_11512,N_9336,N_9010);
nand U11513 (N_11513,N_9759,N_8379);
and U11514 (N_11514,N_9041,N_9664);
xnor U11515 (N_11515,N_8698,N_9351);
nor U11516 (N_11516,N_9416,N_9503);
nand U11517 (N_11517,N_9567,N_8307);
and U11518 (N_11518,N_8505,N_9110);
nand U11519 (N_11519,N_8448,N_9735);
and U11520 (N_11520,N_9434,N_9519);
and U11521 (N_11521,N_8836,N_9224);
nand U11522 (N_11522,N_8109,N_8304);
and U11523 (N_11523,N_9016,N_8272);
xor U11524 (N_11524,N_8709,N_9946);
xnor U11525 (N_11525,N_9058,N_9956);
and U11526 (N_11526,N_9554,N_8032);
nand U11527 (N_11527,N_9672,N_9111);
and U11528 (N_11528,N_9257,N_9913);
or U11529 (N_11529,N_9350,N_9273);
and U11530 (N_11530,N_8315,N_8105);
nand U11531 (N_11531,N_9320,N_9522);
nor U11532 (N_11532,N_8504,N_8068);
xor U11533 (N_11533,N_9530,N_9872);
xnor U11534 (N_11534,N_9698,N_9082);
and U11535 (N_11535,N_9520,N_8946);
and U11536 (N_11536,N_8891,N_8783);
xor U11537 (N_11537,N_9952,N_9340);
nand U11538 (N_11538,N_9735,N_9536);
nor U11539 (N_11539,N_9022,N_9665);
or U11540 (N_11540,N_8204,N_9765);
or U11541 (N_11541,N_8106,N_8623);
and U11542 (N_11542,N_9508,N_8638);
and U11543 (N_11543,N_8059,N_8670);
nand U11544 (N_11544,N_9349,N_9182);
nor U11545 (N_11545,N_8417,N_8836);
or U11546 (N_11546,N_8923,N_8124);
xor U11547 (N_11547,N_8090,N_8417);
nand U11548 (N_11548,N_8507,N_9045);
xnor U11549 (N_11549,N_8448,N_9612);
or U11550 (N_11550,N_8404,N_8143);
xor U11551 (N_11551,N_8357,N_9241);
and U11552 (N_11552,N_8457,N_8308);
xnor U11553 (N_11553,N_8417,N_9600);
and U11554 (N_11554,N_9675,N_9243);
and U11555 (N_11555,N_8723,N_8808);
and U11556 (N_11556,N_8486,N_9579);
nand U11557 (N_11557,N_8769,N_8582);
and U11558 (N_11558,N_8949,N_9461);
or U11559 (N_11559,N_9103,N_8044);
nand U11560 (N_11560,N_9904,N_9635);
and U11561 (N_11561,N_8434,N_9762);
nor U11562 (N_11562,N_9724,N_8570);
nand U11563 (N_11563,N_8589,N_8242);
nor U11564 (N_11564,N_9006,N_8445);
and U11565 (N_11565,N_8265,N_9003);
nor U11566 (N_11566,N_8889,N_8509);
nand U11567 (N_11567,N_9303,N_9000);
nand U11568 (N_11568,N_8630,N_8193);
xor U11569 (N_11569,N_8055,N_8226);
nor U11570 (N_11570,N_9364,N_9118);
nor U11571 (N_11571,N_8706,N_9666);
and U11572 (N_11572,N_9915,N_9801);
xnor U11573 (N_11573,N_8471,N_8727);
and U11574 (N_11574,N_8331,N_8017);
or U11575 (N_11575,N_9287,N_8256);
xnor U11576 (N_11576,N_9998,N_8212);
and U11577 (N_11577,N_9475,N_8312);
or U11578 (N_11578,N_8573,N_9814);
and U11579 (N_11579,N_8856,N_9224);
or U11580 (N_11580,N_9429,N_9800);
and U11581 (N_11581,N_8510,N_8914);
nand U11582 (N_11582,N_9312,N_9371);
or U11583 (N_11583,N_8389,N_9811);
nor U11584 (N_11584,N_8456,N_9776);
or U11585 (N_11585,N_9296,N_9227);
xnor U11586 (N_11586,N_8996,N_9449);
and U11587 (N_11587,N_8355,N_8504);
nor U11588 (N_11588,N_8840,N_8780);
and U11589 (N_11589,N_9406,N_8020);
or U11590 (N_11590,N_8363,N_8361);
nor U11591 (N_11591,N_9580,N_8697);
or U11592 (N_11592,N_8637,N_8722);
nor U11593 (N_11593,N_8762,N_9334);
nor U11594 (N_11594,N_9696,N_9909);
or U11595 (N_11595,N_8774,N_9486);
or U11596 (N_11596,N_8935,N_9510);
xnor U11597 (N_11597,N_8573,N_8727);
or U11598 (N_11598,N_9859,N_8160);
and U11599 (N_11599,N_9555,N_8185);
nand U11600 (N_11600,N_8280,N_9919);
nand U11601 (N_11601,N_8764,N_9315);
xnor U11602 (N_11602,N_9870,N_9942);
or U11603 (N_11603,N_9585,N_8381);
nor U11604 (N_11604,N_9342,N_8001);
or U11605 (N_11605,N_9006,N_9100);
xor U11606 (N_11606,N_8733,N_9811);
and U11607 (N_11607,N_9690,N_9509);
and U11608 (N_11608,N_8780,N_9262);
and U11609 (N_11609,N_9491,N_9205);
or U11610 (N_11610,N_8254,N_8041);
or U11611 (N_11611,N_8927,N_9829);
and U11612 (N_11612,N_8977,N_8006);
or U11613 (N_11613,N_9921,N_8141);
nor U11614 (N_11614,N_9482,N_8533);
nand U11615 (N_11615,N_9887,N_9980);
xnor U11616 (N_11616,N_9196,N_9891);
or U11617 (N_11617,N_8308,N_8154);
nand U11618 (N_11618,N_8720,N_9763);
nand U11619 (N_11619,N_9008,N_8152);
nand U11620 (N_11620,N_8005,N_8197);
nand U11621 (N_11621,N_9014,N_9614);
nand U11622 (N_11622,N_8045,N_9560);
nand U11623 (N_11623,N_8052,N_8844);
xor U11624 (N_11624,N_8951,N_9766);
nor U11625 (N_11625,N_8432,N_8615);
and U11626 (N_11626,N_8202,N_9309);
nor U11627 (N_11627,N_9223,N_8023);
xnor U11628 (N_11628,N_8810,N_8449);
nand U11629 (N_11629,N_8975,N_9421);
nand U11630 (N_11630,N_8775,N_9941);
xnor U11631 (N_11631,N_8568,N_8516);
or U11632 (N_11632,N_8558,N_9084);
nor U11633 (N_11633,N_8986,N_8389);
or U11634 (N_11634,N_9244,N_8889);
nand U11635 (N_11635,N_9868,N_9360);
and U11636 (N_11636,N_8508,N_9155);
nand U11637 (N_11637,N_8615,N_8006);
nand U11638 (N_11638,N_8564,N_9992);
nand U11639 (N_11639,N_9592,N_9226);
nor U11640 (N_11640,N_9543,N_8439);
xor U11641 (N_11641,N_8451,N_9528);
nor U11642 (N_11642,N_9933,N_8128);
nor U11643 (N_11643,N_9120,N_9789);
or U11644 (N_11644,N_8184,N_9095);
nand U11645 (N_11645,N_9615,N_9456);
nand U11646 (N_11646,N_9238,N_9627);
and U11647 (N_11647,N_9874,N_9749);
xnor U11648 (N_11648,N_8260,N_8544);
nand U11649 (N_11649,N_8512,N_8371);
and U11650 (N_11650,N_9435,N_9674);
nor U11651 (N_11651,N_8527,N_8917);
nand U11652 (N_11652,N_8766,N_8778);
xor U11653 (N_11653,N_9323,N_8953);
and U11654 (N_11654,N_8777,N_9507);
and U11655 (N_11655,N_8304,N_9246);
nand U11656 (N_11656,N_9510,N_8191);
and U11657 (N_11657,N_8529,N_8995);
or U11658 (N_11658,N_8528,N_8678);
nor U11659 (N_11659,N_9687,N_8730);
and U11660 (N_11660,N_8733,N_9010);
and U11661 (N_11661,N_9585,N_8619);
and U11662 (N_11662,N_8690,N_8359);
and U11663 (N_11663,N_9892,N_9001);
nand U11664 (N_11664,N_9675,N_9951);
xnor U11665 (N_11665,N_8972,N_9600);
nand U11666 (N_11666,N_8718,N_9234);
nand U11667 (N_11667,N_9747,N_8136);
nand U11668 (N_11668,N_9909,N_9657);
nand U11669 (N_11669,N_8948,N_8991);
nand U11670 (N_11670,N_8401,N_9411);
and U11671 (N_11671,N_8401,N_9386);
nor U11672 (N_11672,N_9971,N_8421);
nand U11673 (N_11673,N_8517,N_8867);
and U11674 (N_11674,N_8743,N_8364);
xnor U11675 (N_11675,N_8785,N_8535);
and U11676 (N_11676,N_8008,N_9186);
nand U11677 (N_11677,N_9467,N_9016);
nor U11678 (N_11678,N_9162,N_9682);
nand U11679 (N_11679,N_8879,N_9078);
nand U11680 (N_11680,N_8324,N_9817);
nand U11681 (N_11681,N_8492,N_9242);
nor U11682 (N_11682,N_9862,N_9930);
and U11683 (N_11683,N_8748,N_8821);
xnor U11684 (N_11684,N_9734,N_9740);
nor U11685 (N_11685,N_8334,N_8819);
or U11686 (N_11686,N_8210,N_8137);
or U11687 (N_11687,N_8498,N_8980);
xnor U11688 (N_11688,N_9093,N_9257);
and U11689 (N_11689,N_8194,N_9699);
nor U11690 (N_11690,N_9097,N_9540);
nor U11691 (N_11691,N_9599,N_9364);
xnor U11692 (N_11692,N_9798,N_8622);
xnor U11693 (N_11693,N_9996,N_8563);
nor U11694 (N_11694,N_8281,N_8038);
or U11695 (N_11695,N_8110,N_9965);
nand U11696 (N_11696,N_8848,N_8032);
or U11697 (N_11697,N_8581,N_8425);
or U11698 (N_11698,N_8686,N_9857);
and U11699 (N_11699,N_8517,N_9524);
nand U11700 (N_11700,N_9475,N_8706);
nand U11701 (N_11701,N_8877,N_9684);
or U11702 (N_11702,N_9499,N_8561);
xnor U11703 (N_11703,N_8972,N_9349);
xnor U11704 (N_11704,N_9430,N_9103);
xor U11705 (N_11705,N_9469,N_9275);
nor U11706 (N_11706,N_9820,N_8214);
nand U11707 (N_11707,N_8680,N_8040);
xnor U11708 (N_11708,N_9202,N_8390);
nand U11709 (N_11709,N_9265,N_9463);
xnor U11710 (N_11710,N_8908,N_9412);
nor U11711 (N_11711,N_9241,N_9691);
xor U11712 (N_11712,N_8407,N_8251);
or U11713 (N_11713,N_9385,N_8523);
or U11714 (N_11714,N_8048,N_9091);
xnor U11715 (N_11715,N_9392,N_8215);
or U11716 (N_11716,N_8749,N_8440);
nand U11717 (N_11717,N_9726,N_9360);
or U11718 (N_11718,N_8134,N_9080);
and U11719 (N_11719,N_9784,N_8363);
xor U11720 (N_11720,N_9744,N_8565);
or U11721 (N_11721,N_9717,N_8887);
and U11722 (N_11722,N_8072,N_9474);
nand U11723 (N_11723,N_8654,N_8022);
xor U11724 (N_11724,N_8930,N_8702);
and U11725 (N_11725,N_8733,N_8490);
xnor U11726 (N_11726,N_8890,N_9281);
nor U11727 (N_11727,N_8033,N_8851);
or U11728 (N_11728,N_9797,N_9167);
xor U11729 (N_11729,N_9938,N_9134);
xor U11730 (N_11730,N_9966,N_9180);
nand U11731 (N_11731,N_8140,N_8693);
and U11732 (N_11732,N_8848,N_9646);
or U11733 (N_11733,N_8123,N_9139);
nand U11734 (N_11734,N_9653,N_9100);
nor U11735 (N_11735,N_8115,N_8211);
xnor U11736 (N_11736,N_9430,N_8588);
nand U11737 (N_11737,N_8748,N_9470);
and U11738 (N_11738,N_9029,N_9386);
nand U11739 (N_11739,N_9124,N_9529);
nor U11740 (N_11740,N_8218,N_9716);
xor U11741 (N_11741,N_8556,N_9372);
nand U11742 (N_11742,N_8497,N_8230);
nor U11743 (N_11743,N_9170,N_8674);
xor U11744 (N_11744,N_9541,N_8130);
xnor U11745 (N_11745,N_8097,N_9606);
or U11746 (N_11746,N_8607,N_9476);
and U11747 (N_11747,N_9939,N_8279);
nand U11748 (N_11748,N_8171,N_8207);
nor U11749 (N_11749,N_9557,N_8762);
and U11750 (N_11750,N_8632,N_9128);
nor U11751 (N_11751,N_9314,N_8614);
xor U11752 (N_11752,N_8752,N_8911);
xor U11753 (N_11753,N_8489,N_8406);
nor U11754 (N_11754,N_8841,N_9907);
xor U11755 (N_11755,N_8330,N_8975);
nor U11756 (N_11756,N_9861,N_8225);
or U11757 (N_11757,N_8932,N_9332);
or U11758 (N_11758,N_8898,N_8888);
nor U11759 (N_11759,N_8607,N_8330);
nand U11760 (N_11760,N_9525,N_9887);
nand U11761 (N_11761,N_9904,N_9914);
nand U11762 (N_11762,N_9662,N_8964);
nand U11763 (N_11763,N_9539,N_8766);
xor U11764 (N_11764,N_8329,N_9975);
xnor U11765 (N_11765,N_9522,N_8685);
nor U11766 (N_11766,N_9295,N_9920);
nor U11767 (N_11767,N_9556,N_8461);
xor U11768 (N_11768,N_8423,N_9695);
xnor U11769 (N_11769,N_9160,N_9751);
and U11770 (N_11770,N_9378,N_8456);
nand U11771 (N_11771,N_9068,N_8846);
and U11772 (N_11772,N_9092,N_9491);
and U11773 (N_11773,N_9311,N_8720);
nor U11774 (N_11774,N_8364,N_9800);
nor U11775 (N_11775,N_9427,N_8566);
xor U11776 (N_11776,N_9517,N_9734);
nor U11777 (N_11777,N_9726,N_9003);
or U11778 (N_11778,N_8040,N_8531);
xnor U11779 (N_11779,N_9504,N_8263);
and U11780 (N_11780,N_8218,N_8711);
and U11781 (N_11781,N_8305,N_8000);
nand U11782 (N_11782,N_9475,N_8490);
nand U11783 (N_11783,N_8439,N_8725);
or U11784 (N_11784,N_9287,N_9098);
xnor U11785 (N_11785,N_9026,N_8915);
or U11786 (N_11786,N_8886,N_8172);
and U11787 (N_11787,N_8703,N_9743);
nand U11788 (N_11788,N_9266,N_8830);
xnor U11789 (N_11789,N_9810,N_8564);
nor U11790 (N_11790,N_8514,N_9002);
nor U11791 (N_11791,N_9372,N_8176);
nand U11792 (N_11792,N_8046,N_9160);
and U11793 (N_11793,N_8952,N_9231);
and U11794 (N_11794,N_9954,N_9734);
nand U11795 (N_11795,N_8231,N_9427);
and U11796 (N_11796,N_9170,N_8101);
and U11797 (N_11797,N_8487,N_9121);
nand U11798 (N_11798,N_8948,N_9829);
xnor U11799 (N_11799,N_9462,N_9860);
or U11800 (N_11800,N_8482,N_8705);
or U11801 (N_11801,N_9598,N_8537);
or U11802 (N_11802,N_9188,N_8889);
nand U11803 (N_11803,N_8403,N_9248);
or U11804 (N_11804,N_9115,N_9940);
nor U11805 (N_11805,N_8819,N_8651);
or U11806 (N_11806,N_9760,N_9265);
xnor U11807 (N_11807,N_9697,N_8989);
xnor U11808 (N_11808,N_9078,N_9296);
nor U11809 (N_11809,N_9883,N_8362);
or U11810 (N_11810,N_9962,N_9842);
xnor U11811 (N_11811,N_9062,N_8485);
nand U11812 (N_11812,N_9286,N_9633);
or U11813 (N_11813,N_8918,N_8117);
or U11814 (N_11814,N_9821,N_8665);
nor U11815 (N_11815,N_8772,N_9610);
and U11816 (N_11816,N_8668,N_9039);
and U11817 (N_11817,N_8004,N_9697);
nor U11818 (N_11818,N_9156,N_8496);
or U11819 (N_11819,N_8242,N_9418);
and U11820 (N_11820,N_8138,N_8184);
nand U11821 (N_11821,N_9112,N_8866);
or U11822 (N_11822,N_8535,N_9100);
xnor U11823 (N_11823,N_9308,N_9369);
nor U11824 (N_11824,N_9791,N_9884);
nand U11825 (N_11825,N_8888,N_8785);
and U11826 (N_11826,N_9587,N_9790);
and U11827 (N_11827,N_9286,N_9671);
and U11828 (N_11828,N_9455,N_8322);
xor U11829 (N_11829,N_8012,N_9572);
or U11830 (N_11830,N_9315,N_8579);
nand U11831 (N_11831,N_8348,N_8390);
and U11832 (N_11832,N_8003,N_9844);
and U11833 (N_11833,N_8767,N_8553);
and U11834 (N_11834,N_8466,N_9456);
and U11835 (N_11835,N_8210,N_9555);
or U11836 (N_11836,N_9855,N_9028);
nor U11837 (N_11837,N_9070,N_9945);
nand U11838 (N_11838,N_9687,N_8910);
nor U11839 (N_11839,N_8355,N_8889);
xnor U11840 (N_11840,N_8399,N_8254);
or U11841 (N_11841,N_8480,N_8246);
or U11842 (N_11842,N_8269,N_9948);
or U11843 (N_11843,N_9273,N_8779);
nor U11844 (N_11844,N_9285,N_8765);
and U11845 (N_11845,N_9169,N_8119);
or U11846 (N_11846,N_9352,N_9119);
nor U11847 (N_11847,N_8236,N_9372);
xor U11848 (N_11848,N_8376,N_9688);
nand U11849 (N_11849,N_9705,N_8124);
nand U11850 (N_11850,N_8679,N_9474);
nor U11851 (N_11851,N_8948,N_8324);
xor U11852 (N_11852,N_9560,N_8178);
xor U11853 (N_11853,N_8870,N_8697);
xnor U11854 (N_11854,N_8741,N_8588);
xor U11855 (N_11855,N_8171,N_9197);
xor U11856 (N_11856,N_9352,N_9954);
and U11857 (N_11857,N_9384,N_9704);
xnor U11858 (N_11858,N_8644,N_9802);
or U11859 (N_11859,N_9056,N_8798);
xnor U11860 (N_11860,N_9415,N_8912);
and U11861 (N_11861,N_9018,N_8849);
xnor U11862 (N_11862,N_8955,N_8296);
nor U11863 (N_11863,N_8578,N_8892);
nor U11864 (N_11864,N_8315,N_8606);
and U11865 (N_11865,N_9686,N_8275);
xnor U11866 (N_11866,N_9976,N_8336);
and U11867 (N_11867,N_9126,N_8791);
xor U11868 (N_11868,N_8524,N_9386);
and U11869 (N_11869,N_8350,N_9859);
xor U11870 (N_11870,N_9357,N_8435);
xor U11871 (N_11871,N_9765,N_8206);
nor U11872 (N_11872,N_9409,N_9687);
xnor U11873 (N_11873,N_9877,N_8538);
or U11874 (N_11874,N_8551,N_8785);
xnor U11875 (N_11875,N_9112,N_8719);
xnor U11876 (N_11876,N_9082,N_8687);
nor U11877 (N_11877,N_8119,N_9575);
nand U11878 (N_11878,N_8997,N_8901);
nand U11879 (N_11879,N_8650,N_8773);
nor U11880 (N_11880,N_9188,N_8547);
or U11881 (N_11881,N_8690,N_8005);
nand U11882 (N_11882,N_8125,N_8179);
nor U11883 (N_11883,N_8839,N_8749);
or U11884 (N_11884,N_9485,N_9063);
nand U11885 (N_11885,N_8521,N_8676);
or U11886 (N_11886,N_8426,N_8478);
nand U11887 (N_11887,N_8699,N_8754);
nor U11888 (N_11888,N_8651,N_9050);
nor U11889 (N_11889,N_8980,N_9686);
nand U11890 (N_11890,N_8702,N_8437);
nand U11891 (N_11891,N_8351,N_8533);
nand U11892 (N_11892,N_8072,N_9300);
or U11893 (N_11893,N_9125,N_8072);
and U11894 (N_11894,N_9445,N_8135);
and U11895 (N_11895,N_9769,N_9930);
or U11896 (N_11896,N_8581,N_9718);
or U11897 (N_11897,N_8052,N_8466);
nand U11898 (N_11898,N_8127,N_9950);
or U11899 (N_11899,N_8433,N_8483);
or U11900 (N_11900,N_8263,N_8894);
and U11901 (N_11901,N_9771,N_8705);
nand U11902 (N_11902,N_8164,N_9156);
nand U11903 (N_11903,N_8804,N_8475);
or U11904 (N_11904,N_8127,N_8979);
nand U11905 (N_11905,N_8290,N_9262);
or U11906 (N_11906,N_9480,N_8696);
and U11907 (N_11907,N_8893,N_9427);
nor U11908 (N_11908,N_9964,N_8910);
or U11909 (N_11909,N_9749,N_9702);
xnor U11910 (N_11910,N_8578,N_9016);
or U11911 (N_11911,N_9124,N_9815);
xnor U11912 (N_11912,N_8692,N_8808);
and U11913 (N_11913,N_8870,N_8696);
nand U11914 (N_11914,N_9622,N_8629);
nand U11915 (N_11915,N_9651,N_9945);
or U11916 (N_11916,N_9959,N_9196);
nor U11917 (N_11917,N_8624,N_9585);
nand U11918 (N_11918,N_9776,N_8162);
xnor U11919 (N_11919,N_8581,N_9957);
nor U11920 (N_11920,N_8449,N_8792);
nand U11921 (N_11921,N_8853,N_9272);
or U11922 (N_11922,N_9600,N_8565);
xor U11923 (N_11923,N_8388,N_8299);
xnor U11924 (N_11924,N_9704,N_9294);
nand U11925 (N_11925,N_8383,N_8850);
and U11926 (N_11926,N_8306,N_8281);
and U11927 (N_11927,N_9759,N_9395);
or U11928 (N_11928,N_8708,N_9248);
or U11929 (N_11929,N_9675,N_9079);
or U11930 (N_11930,N_8127,N_8279);
nor U11931 (N_11931,N_8732,N_8394);
xor U11932 (N_11932,N_8510,N_9687);
nor U11933 (N_11933,N_9822,N_8079);
and U11934 (N_11934,N_8708,N_9762);
nand U11935 (N_11935,N_9755,N_9893);
nor U11936 (N_11936,N_8352,N_9350);
or U11937 (N_11937,N_9419,N_9426);
xnor U11938 (N_11938,N_9223,N_9518);
and U11939 (N_11939,N_8451,N_8492);
nor U11940 (N_11940,N_9224,N_9019);
or U11941 (N_11941,N_8240,N_9098);
xnor U11942 (N_11942,N_8008,N_9683);
xnor U11943 (N_11943,N_8999,N_8720);
and U11944 (N_11944,N_9286,N_9455);
nor U11945 (N_11945,N_8864,N_9998);
or U11946 (N_11946,N_8359,N_9725);
and U11947 (N_11947,N_9303,N_9628);
or U11948 (N_11948,N_8040,N_9341);
and U11949 (N_11949,N_9556,N_9888);
nor U11950 (N_11950,N_8373,N_9380);
or U11951 (N_11951,N_9508,N_8948);
nor U11952 (N_11952,N_9904,N_9094);
nand U11953 (N_11953,N_8320,N_9743);
and U11954 (N_11954,N_8959,N_9370);
or U11955 (N_11955,N_8958,N_9665);
xnor U11956 (N_11956,N_9037,N_9508);
xnor U11957 (N_11957,N_8281,N_8816);
or U11958 (N_11958,N_8096,N_8245);
and U11959 (N_11959,N_9524,N_9068);
nand U11960 (N_11960,N_9536,N_9416);
nand U11961 (N_11961,N_8050,N_8494);
nand U11962 (N_11962,N_9822,N_8848);
or U11963 (N_11963,N_8519,N_9859);
xor U11964 (N_11964,N_9855,N_9729);
and U11965 (N_11965,N_8595,N_9577);
xnor U11966 (N_11966,N_9673,N_9894);
xnor U11967 (N_11967,N_8801,N_8864);
and U11968 (N_11968,N_8222,N_8456);
xnor U11969 (N_11969,N_8951,N_9906);
or U11970 (N_11970,N_9417,N_8596);
or U11971 (N_11971,N_9923,N_8694);
nand U11972 (N_11972,N_9842,N_9599);
xnor U11973 (N_11973,N_9392,N_8512);
and U11974 (N_11974,N_8883,N_9528);
and U11975 (N_11975,N_8410,N_9874);
and U11976 (N_11976,N_8333,N_8268);
xor U11977 (N_11977,N_9900,N_8864);
and U11978 (N_11978,N_9248,N_8339);
and U11979 (N_11979,N_8591,N_9908);
or U11980 (N_11980,N_8525,N_8487);
nor U11981 (N_11981,N_9437,N_8547);
xor U11982 (N_11982,N_8834,N_8683);
xnor U11983 (N_11983,N_8758,N_8902);
nand U11984 (N_11984,N_8040,N_9988);
xor U11985 (N_11985,N_8719,N_9240);
nor U11986 (N_11986,N_9152,N_8595);
nand U11987 (N_11987,N_9404,N_8749);
nor U11988 (N_11988,N_8222,N_9440);
nor U11989 (N_11989,N_8800,N_8804);
or U11990 (N_11990,N_8670,N_9293);
and U11991 (N_11991,N_9311,N_8549);
nor U11992 (N_11992,N_9251,N_9689);
nor U11993 (N_11993,N_9830,N_8124);
xor U11994 (N_11994,N_9469,N_9845);
xnor U11995 (N_11995,N_9693,N_9654);
and U11996 (N_11996,N_9428,N_9668);
nor U11997 (N_11997,N_9562,N_9013);
xor U11998 (N_11998,N_8818,N_9454);
xnor U11999 (N_11999,N_8858,N_8080);
nand U12000 (N_12000,N_11920,N_10369);
nand U12001 (N_12001,N_10697,N_10184);
or U12002 (N_12002,N_10969,N_10037);
or U12003 (N_12003,N_10512,N_10457);
or U12004 (N_12004,N_10963,N_10667);
or U12005 (N_12005,N_11618,N_10953);
and U12006 (N_12006,N_11680,N_11347);
or U12007 (N_12007,N_10873,N_10065);
or U12008 (N_12008,N_11393,N_11874);
nand U12009 (N_12009,N_10533,N_10284);
xor U12010 (N_12010,N_11947,N_10487);
and U12011 (N_12011,N_11610,N_10246);
or U12012 (N_12012,N_11217,N_10332);
xor U12013 (N_12013,N_11853,N_11536);
xnor U12014 (N_12014,N_11132,N_10554);
nand U12015 (N_12015,N_10991,N_10053);
or U12016 (N_12016,N_10012,N_11923);
nor U12017 (N_12017,N_11272,N_11230);
xnor U12018 (N_12018,N_11053,N_11124);
nor U12019 (N_12019,N_10608,N_11940);
xor U12020 (N_12020,N_11142,N_11390);
nand U12021 (N_12021,N_10511,N_10627);
xor U12022 (N_12022,N_10919,N_10326);
nand U12023 (N_12023,N_11308,N_10148);
nand U12024 (N_12024,N_11577,N_10207);
and U12025 (N_12025,N_10222,N_11777);
nor U12026 (N_12026,N_10147,N_10474);
or U12027 (N_12027,N_10894,N_11741);
or U12028 (N_12028,N_11918,N_11461);
xnor U12029 (N_12029,N_11269,N_10164);
nor U12030 (N_12030,N_11520,N_10393);
xor U12031 (N_12031,N_11103,N_10019);
and U12032 (N_12032,N_11973,N_10643);
nand U12033 (N_12033,N_10906,N_11411);
nor U12034 (N_12034,N_11449,N_11114);
nand U12035 (N_12035,N_10550,N_11740);
xor U12036 (N_12036,N_11842,N_11025);
or U12037 (N_12037,N_10366,N_11098);
nor U12038 (N_12038,N_10816,N_11589);
nand U12039 (N_12039,N_10997,N_11956);
or U12040 (N_12040,N_11338,N_11678);
nor U12041 (N_12041,N_10327,N_11819);
nand U12042 (N_12042,N_10276,N_10224);
and U12043 (N_12043,N_10828,N_10417);
and U12044 (N_12044,N_10678,N_10005);
and U12045 (N_12045,N_11910,N_10617);
nand U12046 (N_12046,N_10820,N_11993);
nor U12047 (N_12047,N_11070,N_10806);
xor U12048 (N_12048,N_11800,N_11722);
xnor U12049 (N_12049,N_10647,N_11454);
nand U12050 (N_12050,N_10600,N_10239);
nand U12051 (N_12051,N_10582,N_11609);
xnor U12052 (N_12052,N_11962,N_10888);
nand U12053 (N_12053,N_11882,N_11681);
and U12054 (N_12054,N_10498,N_11653);
or U12055 (N_12055,N_11541,N_11106);
nor U12056 (N_12056,N_11237,N_10572);
nor U12057 (N_12057,N_10435,N_11789);
xor U12058 (N_12058,N_10934,N_10334);
nand U12059 (N_12059,N_11959,N_10022);
and U12060 (N_12060,N_10928,N_11167);
or U12061 (N_12061,N_10531,N_11251);
and U12062 (N_12062,N_10350,N_11188);
xnor U12063 (N_12063,N_11970,N_11847);
and U12064 (N_12064,N_11627,N_11136);
and U12065 (N_12065,N_11265,N_10030);
and U12066 (N_12066,N_10727,N_11805);
xor U12067 (N_12067,N_11259,N_11340);
xor U12068 (N_12068,N_10559,N_10154);
or U12069 (N_12069,N_10416,N_11359);
nand U12070 (N_12070,N_11138,N_11643);
or U12071 (N_12071,N_11456,N_10201);
and U12072 (N_12072,N_11603,N_11980);
nand U12073 (N_12073,N_11398,N_10268);
xnor U12074 (N_12074,N_10557,N_10578);
nor U12075 (N_12075,N_11987,N_10931);
xnor U12076 (N_12076,N_11109,N_11650);
xor U12077 (N_12077,N_11858,N_11864);
nor U12078 (N_12078,N_10419,N_11171);
nand U12079 (N_12079,N_11943,N_10293);
and U12080 (N_12080,N_11620,N_11074);
and U12081 (N_12081,N_10981,N_11691);
and U12082 (N_12082,N_10575,N_10169);
nor U12083 (N_12083,N_11976,N_11424);
nand U12084 (N_12084,N_11538,N_10846);
or U12085 (N_12085,N_11032,N_11255);
nand U12086 (N_12086,N_10792,N_10176);
nand U12087 (N_12087,N_10145,N_10886);
and U12088 (N_12088,N_11231,N_11991);
nor U12089 (N_12089,N_11688,N_10493);
xor U12090 (N_12090,N_11376,N_11008);
nand U12091 (N_12091,N_10616,N_10236);
nand U12092 (N_12092,N_11952,N_10372);
xnor U12093 (N_12093,N_10755,N_10687);
xor U12094 (N_12094,N_10871,N_11178);
or U12095 (N_12095,N_11838,N_10129);
or U12096 (N_12096,N_11739,N_11222);
nand U12097 (N_12097,N_11969,N_11915);
xnor U12098 (N_12098,N_11556,N_10014);
xor U12099 (N_12099,N_11857,N_10759);
or U12100 (N_12100,N_10321,N_11594);
and U12101 (N_12101,N_10543,N_10202);
xnor U12102 (N_12102,N_10860,N_11082);
or U12103 (N_12103,N_11247,N_10814);
xor U12104 (N_12104,N_10371,N_11601);
or U12105 (N_12105,N_11825,N_10944);
or U12106 (N_12106,N_10445,N_10093);
nand U12107 (N_12107,N_10714,N_10349);
and U12108 (N_12108,N_11661,N_10181);
nor U12109 (N_12109,N_10982,N_11254);
nand U12110 (N_12110,N_11914,N_10866);
nor U12111 (N_12111,N_11563,N_11561);
xor U12112 (N_12112,N_11671,N_10735);
or U12113 (N_12113,N_10618,N_10206);
nand U12114 (N_12114,N_11266,N_11704);
xor U12115 (N_12115,N_10355,N_10116);
nor U12116 (N_12116,N_10933,N_10249);
xnor U12117 (N_12117,N_10753,N_10441);
xor U12118 (N_12118,N_10943,N_11094);
xnor U12119 (N_12119,N_10291,N_11925);
nand U12120 (N_12120,N_10825,N_10298);
and U12121 (N_12121,N_11723,N_11139);
xnor U12122 (N_12122,N_11485,N_11472);
nor U12123 (N_12123,N_11227,N_10604);
nand U12124 (N_12124,N_10706,N_11768);
or U12125 (N_12125,N_10320,N_11406);
and U12126 (N_12126,N_11089,N_11043);
nor U12127 (N_12127,N_11159,N_10813);
nand U12128 (N_12128,N_11913,N_11718);
xnor U12129 (N_12129,N_10345,N_11870);
nor U12130 (N_12130,N_10035,N_11083);
nand U12131 (N_12131,N_10168,N_10266);
nor U12132 (N_12132,N_10672,N_11007);
nand U12133 (N_12133,N_10044,N_11125);
nor U12134 (N_12134,N_11960,N_11885);
xnor U12135 (N_12135,N_10177,N_10704);
nor U12136 (N_12136,N_10950,N_11889);
nand U12137 (N_12137,N_10397,N_10640);
nor U12138 (N_12138,N_11558,N_10270);
and U12139 (N_12139,N_10862,N_11386);
and U12140 (N_12140,N_10954,N_11896);
xnor U12141 (N_12141,N_10114,N_10278);
xnor U12142 (N_12142,N_10252,N_10167);
xor U12143 (N_12143,N_10395,N_10898);
nor U12144 (N_12144,N_10175,N_11513);
or U12145 (N_12145,N_11154,N_11489);
nand U12146 (N_12146,N_10107,N_11562);
or U12147 (N_12147,N_10700,N_11758);
and U12148 (N_12148,N_11281,N_11782);
nand U12149 (N_12149,N_10884,N_11963);
nand U12150 (N_12150,N_10624,N_11057);
or U12151 (N_12151,N_11371,N_10213);
nand U12152 (N_12152,N_10485,N_11286);
and U12153 (N_12153,N_10516,N_10054);
xnor U12154 (N_12154,N_10221,N_11431);
or U12155 (N_12155,N_11719,N_11039);
nand U12156 (N_12156,N_10635,N_10446);
and U12157 (N_12157,N_10021,N_11937);
and U12158 (N_12158,N_10563,N_10621);
or U12159 (N_12159,N_10583,N_11994);
nor U12160 (N_12160,N_10243,N_10108);
or U12161 (N_12161,N_10212,N_10240);
nand U12162 (N_12162,N_10570,N_10799);
xnor U12163 (N_12163,N_10002,N_10318);
nand U12164 (N_12164,N_11771,N_11023);
or U12165 (N_12165,N_10805,N_10070);
xor U12166 (N_12166,N_10833,N_11897);
xnor U12167 (N_12167,N_11900,N_11717);
nand U12168 (N_12168,N_10936,N_11588);
and U12169 (N_12169,N_10786,N_11599);
nor U12170 (N_12170,N_11193,N_11555);
nand U12171 (N_12171,N_10089,N_11645);
and U12172 (N_12172,N_10074,N_11133);
and U12173 (N_12173,N_10962,N_10957);
nor U12174 (N_12174,N_11968,N_10025);
nand U12175 (N_12175,N_10602,N_10453);
nand U12176 (N_12176,N_11699,N_10245);
or U12177 (N_12177,N_10692,N_11370);
nand U12178 (N_12178,N_10673,N_10705);
xor U12179 (N_12179,N_11027,N_10426);
nor U12180 (N_12180,N_11773,N_11880);
and U12181 (N_12181,N_10679,N_10849);
nand U12182 (N_12182,N_10540,N_10254);
or U12183 (N_12183,N_11336,N_10132);
nand U12184 (N_12184,N_11835,N_10724);
or U12185 (N_12185,N_11426,N_10611);
xor U12186 (N_12186,N_10889,N_11774);
xor U12187 (N_12187,N_10845,N_10768);
nand U12188 (N_12188,N_11238,N_11614);
and U12189 (N_12189,N_10674,N_10102);
or U12190 (N_12190,N_11997,N_10058);
or U12191 (N_12191,N_11232,N_11236);
and U12192 (N_12192,N_10960,N_10762);
nor U12193 (N_12193,N_11213,N_10411);
nand U12194 (N_12194,N_11047,N_10425);
nor U12195 (N_12195,N_10096,N_10682);
nand U12196 (N_12196,N_11088,N_11930);
xnor U12197 (N_12197,N_10277,N_11743);
xnor U12198 (N_12198,N_10381,N_10171);
or U12199 (N_12199,N_10377,N_11625);
nor U12200 (N_12200,N_10358,N_11146);
xor U12201 (N_12201,N_11045,N_10351);
xnor U12202 (N_12202,N_10987,N_11097);
nand U12203 (N_12203,N_10402,N_11184);
nor U12204 (N_12204,N_11784,N_11294);
nor U12205 (N_12205,N_10439,N_11420);
xor U12206 (N_12206,N_11388,N_10086);
nor U12207 (N_12207,N_11175,N_10522);
or U12208 (N_12208,N_10297,N_10194);
nor U12209 (N_12209,N_11600,N_10091);
and U12210 (N_12210,N_10574,N_10269);
or U12211 (N_12211,N_10885,N_11587);
nand U12212 (N_12212,N_10422,N_11892);
nor U12213 (N_12213,N_11615,N_10784);
xnor U12214 (N_12214,N_11333,N_11462);
nand U12215 (N_12215,N_10219,N_10496);
or U12216 (N_12216,N_11715,N_10754);
nand U12217 (N_12217,N_11380,N_11433);
nand U12218 (N_12218,N_11831,N_10788);
nand U12219 (N_12219,N_11516,N_11651);
nand U12220 (N_12220,N_10923,N_10110);
nor U12221 (N_12221,N_10357,N_10447);
or U12222 (N_12222,N_10904,N_10038);
nor U12223 (N_12223,N_11760,N_10659);
nand U12224 (N_12224,N_11046,N_10189);
nand U12225 (N_12225,N_11612,N_10598);
nor U12226 (N_12226,N_10980,N_10782);
nand U12227 (N_12227,N_11578,N_11071);
or U12228 (N_12228,N_11355,N_11669);
xor U12229 (N_12229,N_10192,N_10015);
nand U12230 (N_12230,N_11644,N_10263);
or U12231 (N_12231,N_11826,N_10549);
xnor U12232 (N_12232,N_11697,N_10490);
or U12233 (N_12233,N_11078,N_10296);
and U12234 (N_12234,N_10329,N_10112);
nor U12235 (N_12235,N_11321,N_10289);
or U12236 (N_12236,N_10031,N_11529);
nand U12237 (N_12237,N_11324,N_11545);
nor U12238 (N_12238,N_10195,N_10795);
nor U12239 (N_12239,N_10551,N_10257);
xnor U12240 (N_12240,N_11730,N_10662);
nand U12241 (N_12241,N_11596,N_10527);
or U12242 (N_12242,N_10039,N_11537);
nand U12243 (N_12243,N_11099,N_11102);
xnor U12244 (N_12244,N_11938,N_11451);
and U12245 (N_12245,N_10890,N_11040);
and U12246 (N_12246,N_10737,N_10119);
nand U12247 (N_12247,N_11067,N_11873);
and U12248 (N_12248,N_10907,N_11817);
nor U12249 (N_12249,N_10810,N_10227);
nand U12250 (N_12250,N_11002,N_10769);
or U12251 (N_12251,N_11483,N_10279);
or U12252 (N_12252,N_10536,N_10363);
xor U12253 (N_12253,N_11328,N_11048);
nor U12254 (N_12254,N_11157,N_11063);
xor U12255 (N_12255,N_11244,N_11246);
or U12256 (N_12256,N_11158,N_10712);
or U12257 (N_12257,N_10275,N_10644);
and U12258 (N_12258,N_10558,N_11534);
xor U12259 (N_12259,N_11170,N_11341);
and U12260 (N_12260,N_10178,N_11539);
nor U12261 (N_12261,N_11110,N_11945);
nand U12262 (N_12262,N_10793,N_10838);
and U12263 (N_12263,N_11497,N_11482);
xnor U12264 (N_12264,N_11095,N_11313);
xor U12265 (N_12265,N_10491,N_11381);
nor U12266 (N_12266,N_10354,N_10681);
nand U12267 (N_12267,N_10095,N_11279);
xor U12268 (N_12268,N_11983,N_11278);
nor U12269 (N_12269,N_10566,N_11665);
nand U12270 (N_12270,N_11323,N_10580);
nor U12271 (N_12271,N_10314,N_10859);
or U12272 (N_12272,N_10316,N_10568);
nor U12273 (N_12273,N_11495,N_10218);
or U12274 (N_12274,N_10916,N_11827);
nor U12275 (N_12275,N_10995,N_10390);
xnor U12276 (N_12276,N_10478,N_11844);
xnor U12277 (N_12277,N_10630,N_10658);
or U12278 (N_12278,N_11107,N_11590);
or U12279 (N_12279,N_11392,N_10779);
or U12280 (N_12280,N_10949,N_11405);
and U12281 (N_12281,N_10143,N_10826);
nand U12282 (N_12282,N_10896,N_11385);
xor U12283 (N_12283,N_11734,N_10250);
xnor U12284 (N_12284,N_11121,N_11469);
and U12285 (N_12285,N_11573,N_10521);
xor U12286 (N_12286,N_10761,N_11737);
or U12287 (N_12287,N_11004,N_10106);
xor U12288 (N_12288,N_11458,N_11069);
xor U12289 (N_12289,N_11985,N_10695);
or U12290 (N_12290,N_10908,N_11149);
xnor U12291 (N_12291,N_11978,N_10688);
nand U12292 (N_12292,N_10292,N_11092);
or U12293 (N_12293,N_11367,N_11169);
or U12294 (N_12294,N_10383,N_11260);
or U12295 (N_12295,N_11394,N_11830);
or U12296 (N_12296,N_10313,N_10514);
nor U12297 (N_12297,N_11794,N_10398);
nand U12298 (N_12298,N_10821,N_11905);
xnor U12299 (N_12299,N_11037,N_11929);
or U12300 (N_12300,N_11856,N_10128);
nand U12301 (N_12301,N_11126,N_11443);
nor U12302 (N_12302,N_10046,N_11814);
xnor U12303 (N_12303,N_11346,N_10698);
xor U12304 (N_12304,N_11877,N_10264);
and U12305 (N_12305,N_11631,N_11434);
or U12306 (N_12306,N_11018,N_10396);
xor U12307 (N_12307,N_10994,N_11862);
or U12308 (N_12308,N_10481,N_11571);
or U12309 (N_12309,N_11508,N_10940);
or U12310 (N_12310,N_10310,N_10752);
nand U12311 (N_12311,N_11716,N_10707);
xnor U12312 (N_12312,N_10034,N_11626);
nand U12313 (N_12313,N_10857,N_11064);
and U12314 (N_12314,N_10475,N_11478);
nand U12315 (N_12315,N_10140,N_10160);
or U12316 (N_12316,N_10587,N_11944);
and U12317 (N_12317,N_10385,N_10099);
or U12318 (N_12318,N_10092,N_10599);
and U12319 (N_12319,N_11559,N_10626);
nand U12320 (N_12320,N_10946,N_11014);
and U12321 (N_12321,N_11453,N_10758);
and U12322 (N_12322,N_10083,N_11177);
xnor U12323 (N_12323,N_10651,N_10430);
xnor U12324 (N_12324,N_11641,N_10466);
nor U12325 (N_12325,N_10454,N_11635);
nor U12326 (N_12326,N_11711,N_10412);
nor U12327 (N_12327,N_10469,N_10448);
or U12328 (N_12328,N_10051,N_11179);
and U12329 (N_12329,N_11554,N_10852);
nand U12330 (N_12330,N_10556,N_11989);
and U12331 (N_12331,N_10855,N_11764);
nor U12332 (N_12332,N_10636,N_10338);
or U12333 (N_12333,N_10503,N_11696);
and U12334 (N_12334,N_11153,N_11242);
nand U12335 (N_12335,N_10130,N_11253);
or U12336 (N_12336,N_11274,N_11720);
nand U12337 (N_12337,N_11423,N_10376);
and U12338 (N_12338,N_11576,N_10449);
nand U12339 (N_12339,N_11506,N_11954);
nand U12340 (N_12340,N_10348,N_10042);
nand U12341 (N_12341,N_10080,N_10302);
nor U12342 (N_12342,N_11565,N_10879);
nand U12343 (N_12343,N_10062,N_11769);
or U12344 (N_12344,N_11331,N_11709);
nand U12345 (N_12345,N_10229,N_11505);
nand U12346 (N_12346,N_10591,N_10965);
xor U12347 (N_12347,N_10978,N_11310);
xnor U12348 (N_12348,N_10488,N_11019);
and U12349 (N_12349,N_10063,N_11387);
and U12350 (N_12350,N_11372,N_10166);
and U12351 (N_12351,N_11668,N_10186);
nor U12352 (N_12352,N_11912,N_10586);
or U12353 (N_12353,N_10328,N_11339);
or U12354 (N_12354,N_10897,N_11619);
or U12355 (N_12355,N_10592,N_11686);
nand U12356 (N_12356,N_11223,N_10356);
and U12357 (N_12357,N_11130,N_10473);
xor U12358 (N_12358,N_11654,N_10476);
and U12359 (N_12359,N_10585,N_11235);
nor U12360 (N_12360,N_10024,N_11942);
nor U12361 (N_12361,N_11195,N_10406);
nor U12362 (N_12362,N_11772,N_10492);
and U12363 (N_12363,N_10625,N_10122);
nor U12364 (N_12364,N_11417,N_10920);
nor U12365 (N_12365,N_11872,N_11318);
and U12366 (N_12366,N_11438,N_11250);
or U12367 (N_12367,N_11374,N_10217);
nand U12368 (N_12368,N_11904,N_11172);
and U12369 (N_12369,N_10341,N_10529);
nand U12370 (N_12370,N_10840,N_10507);
nand U12371 (N_12371,N_11593,N_11186);
and U12372 (N_12372,N_11721,N_11868);
xnor U12373 (N_12373,N_10751,N_11778);
nor U12374 (N_12374,N_10501,N_11068);
xor U12375 (N_12375,N_10827,N_10770);
nor U12376 (N_12376,N_11448,N_11893);
xnor U12377 (N_12377,N_10374,N_10418);
and U12378 (N_12378,N_11248,N_10209);
or U12379 (N_12379,N_10708,N_11334);
nor U12380 (N_12380,N_10938,N_11833);
nor U12381 (N_12381,N_11181,N_11519);
nor U12382 (N_12382,N_10156,N_11551);
xor U12383 (N_12383,N_11442,N_11163);
nor U12384 (N_12384,N_11304,N_10780);
nor U12385 (N_12385,N_10026,N_10103);
or U12386 (N_12386,N_10670,N_10979);
nand U12387 (N_12387,N_10620,N_11401);
nor U12388 (N_12388,N_10520,N_10922);
nand U12389 (N_12389,N_10016,N_11028);
nor U12390 (N_12390,N_10282,N_10502);
nand U12391 (N_12391,N_10807,N_10842);
or U12392 (N_12392,N_11876,N_10388);
and U12393 (N_12393,N_11271,N_10861);
nor U12394 (N_12394,N_11807,N_11036);
or U12395 (N_12395,N_11792,N_10094);
nand U12396 (N_12396,N_10389,N_10011);
nand U12397 (N_12397,N_10100,N_10652);
and U12398 (N_12398,N_11343,N_11957);
nor U12399 (N_12399,N_10403,N_10200);
xnor U12400 (N_12400,N_10961,N_11790);
and U12401 (N_12401,N_11510,N_11640);
and U12402 (N_12402,N_10346,N_11081);
nand U12403 (N_12403,N_11682,N_11672);
and U12404 (N_12404,N_11639,N_11818);
and U12405 (N_12405,N_10691,N_10596);
or U12406 (N_12406,N_11473,N_11560);
or U12407 (N_12407,N_11127,N_11086);
nand U12408 (N_12408,N_10258,N_10149);
nor U12409 (N_12409,N_11487,N_11292);
or U12410 (N_12410,N_11552,N_11305);
xor U12411 (N_12411,N_10135,N_11252);
nor U12412 (N_12412,N_10220,N_11958);
nor U12413 (N_12413,N_10500,N_10379);
nand U12414 (N_12414,N_11974,N_11349);
and U12415 (N_12415,N_10120,N_10665);
or U12416 (N_12416,N_11585,N_11779);
xnor U12417 (N_12417,N_11821,N_10548);
nand U12418 (N_12418,N_10226,N_10087);
nor U12419 (N_12419,N_11646,N_11525);
or U12420 (N_12420,N_10992,N_10368);
nor U12421 (N_12421,N_10937,N_11907);
or U12422 (N_12422,N_11141,N_10524);
nand U12423 (N_12423,N_10900,N_11982);
nor U12424 (N_12424,N_11113,N_11058);
or U12425 (N_12425,N_11311,N_10560);
nand U12426 (N_12426,N_11137,N_10050);
and U12427 (N_12427,N_10959,N_11753);
xor U12428 (N_12428,N_11834,N_11861);
nor U12429 (N_12429,N_10082,N_11926);
xor U12430 (N_12430,N_10942,N_11147);
and U12431 (N_12431,N_11330,N_10832);
nand U12432 (N_12432,N_10639,N_11636);
and U12433 (N_12433,N_11013,N_11895);
xnor U12434 (N_12434,N_10434,N_11972);
xnor U12435 (N_12435,N_11581,N_11233);
nand U12436 (N_12436,N_11574,N_11592);
xnor U12437 (N_12437,N_10028,N_10460);
nand U12438 (N_12438,N_10047,N_10459);
nor U12439 (N_12439,N_11815,N_11161);
nor U12440 (N_12440,N_10131,N_11724);
nand U12441 (N_12441,N_11979,N_11775);
and U12442 (N_12442,N_10935,N_10125);
or U12443 (N_12443,N_11403,N_10683);
nand U12444 (N_12444,N_11878,N_10072);
nor U12445 (N_12445,N_10274,N_11580);
or U12446 (N_12446,N_10834,N_11084);
and U12447 (N_12447,N_10101,N_10191);
nor U12448 (N_12448,N_11791,N_11738);
and U12449 (N_12449,N_10711,N_10068);
or U12450 (N_12450,N_10251,N_11542);
or U12451 (N_12451,N_11396,N_10456);
nor U12452 (N_12452,N_11445,N_10150);
or U12453 (N_12453,N_10510,N_10676);
nor U12454 (N_12454,N_10489,N_10528);
or U12455 (N_12455,N_10465,N_10734);
xnor U12456 (N_12456,N_10073,N_10399);
xnor U12457 (N_12457,N_10664,N_11350);
nor U12458 (N_12458,N_11140,N_11378);
and U12459 (N_12459,N_10594,N_11984);
or U12460 (N_12460,N_10174,N_10428);
xor U12461 (N_12461,N_10882,N_11630);
and U12462 (N_12462,N_11005,N_11368);
or U12463 (N_12463,N_11463,N_11700);
nor U12464 (N_12464,N_10000,N_11634);
and U12465 (N_12465,N_11303,N_10305);
xor U12466 (N_12466,N_10634,N_11884);
nor U12467 (N_12467,N_11632,N_11129);
nor U12468 (N_12468,N_11591,N_10455);
nor U12469 (N_12469,N_10188,N_10800);
xnor U12470 (N_12470,N_11117,N_11429);
and U12471 (N_12471,N_11091,N_11267);
or U12472 (N_12472,N_11933,N_11898);
or U12473 (N_12473,N_10079,N_11909);
xor U12474 (N_12474,N_11312,N_10391);
nand U12475 (N_12475,N_10464,N_10948);
and U12476 (N_12476,N_11264,N_11795);
xnor U12477 (N_12477,N_10610,N_10253);
or U12478 (N_12478,N_10774,N_10287);
or U12479 (N_12479,N_11888,N_11452);
xnor U12480 (N_12480,N_11356,N_11515);
xor U12481 (N_12481,N_11781,N_10941);
and U12482 (N_12482,N_11345,N_10956);
nand U12483 (N_12483,N_10539,N_10384);
nand U12484 (N_12484,N_10631,N_10179);
nor U12485 (N_12485,N_10836,N_10027);
and U12486 (N_12486,N_11622,N_10699);
nor U12487 (N_12487,N_10869,N_10360);
and U12488 (N_12488,N_10077,N_11362);
and U12489 (N_12489,N_10421,N_10165);
nor U12490 (N_12490,N_11637,N_10043);
xnor U12491 (N_12491,N_11421,N_10370);
nor U12492 (N_12492,N_10424,N_11490);
nor U12493 (N_12493,N_10579,N_11295);
nand U12494 (N_12494,N_10470,N_11301);
nor U12495 (N_12495,N_10415,N_11762);
xnor U12496 (N_12496,N_11761,N_11360);
xor U12497 (N_12497,N_10153,N_11531);
and U12498 (N_12498,N_11553,N_10367);
or U12499 (N_12499,N_11547,N_10715);
or U12500 (N_12500,N_10892,N_11220);
xnor U12501 (N_12501,N_11702,N_11852);
or U12502 (N_12502,N_10760,N_11754);
or U12503 (N_12503,N_11801,N_11948);
and U12504 (N_12504,N_11832,N_11257);
xor U12505 (N_12505,N_10713,N_11747);
nand U12506 (N_12506,N_11052,N_11206);
xor U12507 (N_12507,N_11932,N_11621);
nor U12508 (N_12508,N_10914,N_11501);
and U12509 (N_12509,N_11262,N_11494);
nor U12510 (N_12510,N_10158,N_10525);
nand U12511 (N_12511,N_10060,N_10364);
and U12512 (N_12512,N_10309,N_10538);
nor U12513 (N_12513,N_10835,N_10378);
nor U12514 (N_12514,N_11111,N_10420);
and U12515 (N_12515,N_11072,N_11733);
and U12516 (N_12516,N_10505,N_10286);
nand U12517 (N_12517,N_11470,N_10144);
or U12518 (N_12518,N_11353,N_11093);
nor U12519 (N_12519,N_11604,N_10067);
nor U12520 (N_12520,N_11075,N_11384);
nor U12521 (N_12521,N_11759,N_10561);
or U12522 (N_12522,N_11729,N_10504);
and U12523 (N_12523,N_10117,N_11010);
nor U12524 (N_12524,N_10461,N_11629);
nor U12525 (N_12525,N_10661,N_10623);
or U12526 (N_12526,N_10650,N_11517);
and U12527 (N_12527,N_10686,N_10818);
xor U12528 (N_12528,N_10637,N_10265);
or U12529 (N_12529,N_11316,N_11981);
or U12530 (N_12530,N_11191,N_10951);
nor U12531 (N_12531,N_10552,N_10105);
and U12532 (N_12532,N_11408,N_11457);
nor U12533 (N_12533,N_10482,N_11751);
nand U12534 (N_12534,N_11812,N_10562);
nor U12535 (N_12535,N_10947,N_10571);
xor U12536 (N_12536,N_11901,N_10317);
or U12537 (N_12537,N_10032,N_10055);
xor U12538 (N_12538,N_10064,N_10766);
xnor U12539 (N_12539,N_11908,N_10127);
xor U12540 (N_12540,N_10577,N_10789);
or U12541 (N_12541,N_11887,N_11329);
nor U12542 (N_12542,N_11911,N_11820);
xor U12543 (N_12543,N_10183,N_11056);
nor U12544 (N_12544,N_10427,N_11361);
and U12545 (N_12545,N_10613,N_11413);
nand U12546 (N_12546,N_10796,N_11243);
nor U12547 (N_12547,N_10812,N_11755);
and U12548 (N_12548,N_11667,N_10205);
xor U12549 (N_12549,N_11208,N_10241);
nor U12550 (N_12550,N_10300,N_10573);
and U12551 (N_12551,N_11710,N_11003);
and U12552 (N_12552,N_10663,N_11992);
nand U12553 (N_12553,N_11572,N_11535);
nor U12554 (N_12554,N_11288,N_10872);
or U12555 (N_12555,N_10917,N_10155);
and U12556 (N_12556,N_11694,N_10040);
and U12557 (N_12557,N_11846,N_11021);
xnor U12558 (N_12558,N_10646,N_11532);
and U12559 (N_12559,N_10359,N_11679);
nor U12560 (N_12560,N_11090,N_10020);
and U12561 (N_12561,N_11066,N_11291);
and U12562 (N_12562,N_10392,N_10113);
xnor U12563 (N_12563,N_11750,N_10023);
and U12564 (N_12564,N_10976,N_11509);
or U12565 (N_12565,N_11026,N_10008);
or U12566 (N_12566,N_11767,N_11055);
and U12567 (N_12567,N_10856,N_10233);
nor U12568 (N_12568,N_11961,N_10085);
and U12569 (N_12569,N_10208,N_11602);
xor U12570 (N_12570,N_10151,N_10124);
and U12571 (N_12571,N_11215,N_11986);
nor U12572 (N_12572,N_10903,N_11258);
or U12573 (N_12573,N_10535,N_11836);
xnor U12574 (N_12574,N_11297,N_11647);
and U12575 (N_12575,N_11224,N_10036);
or U12576 (N_12576,N_10876,N_10437);
nand U12577 (N_12577,N_11168,N_10731);
and U12578 (N_12578,N_11030,N_10983);
xor U12579 (N_12579,N_10353,N_10677);
or U12580 (N_12580,N_11152,N_10701);
or U12581 (N_12581,N_10052,N_11379);
nand U12582 (N_12582,N_11863,N_10290);
nor U12583 (N_12583,N_11466,N_10506);
or U12584 (N_12584,N_10971,N_11798);
or U12585 (N_12585,N_11488,N_10546);
nand U12586 (N_12586,N_11879,N_11412);
nand U12587 (N_12587,N_11471,N_10405);
and U12588 (N_12588,N_10401,N_10394);
xnor U12589 (N_12589,N_10765,N_10875);
and U12590 (N_12590,N_11101,N_10049);
nor U12591 (N_12591,N_11162,N_11616);
or U12592 (N_12592,N_11397,N_10984);
nor U12593 (N_12593,N_11809,N_11756);
nor U12594 (N_12594,N_10729,N_11060);
xnor U12595 (N_12595,N_10237,N_10654);
and U12596 (N_12596,N_10771,N_11732);
xnor U12597 (N_12597,N_10271,N_11924);
nor U12598 (N_12598,N_11218,N_10773);
nand U12599 (N_12599,N_10312,N_10718);
or U12600 (N_12600,N_10532,N_11674);
xor U12601 (N_12601,N_11810,N_11624);
xor U12602 (N_12602,N_10743,N_10451);
and U12603 (N_12603,N_11659,N_10337);
nor U12604 (N_12604,N_11492,N_11366);
xnor U12605 (N_12605,N_11319,N_11684);
nor U12606 (N_12606,N_11673,N_11804);
and U12607 (N_12607,N_11033,N_10881);
xnor U12608 (N_12608,N_10738,N_10939);
or U12609 (N_12609,N_11249,N_10605);
nor U12610 (N_12610,N_11617,N_11953);
xor U12611 (N_12611,N_10137,N_10696);
or U12612 (N_12612,N_10895,N_10214);
nor U12613 (N_12613,N_11939,N_10576);
xor U12614 (N_12614,N_10172,N_11802);
and U12615 (N_12615,N_10361,N_10104);
xnor U12616 (N_12616,N_11207,N_10952);
or U12617 (N_12617,N_11173,N_11692);
nor U12618 (N_12618,N_11797,N_11450);
xor U12619 (N_12619,N_11557,N_10985);
and U12620 (N_12620,N_10141,N_10438);
xor U12621 (N_12621,N_11428,N_10854);
or U12622 (N_12622,N_10003,N_10720);
nand U12623 (N_12623,N_10918,N_10858);
nand U12624 (N_12624,N_11706,N_11183);
xor U12625 (N_12625,N_10733,N_11080);
xnor U12626 (N_12626,N_11185,N_10615);
and U12627 (N_12627,N_10781,N_11034);
nand U12628 (N_12628,N_11916,N_10336);
xnor U12629 (N_12629,N_11239,N_11714);
nor U12630 (N_12630,N_11848,N_10228);
or U12631 (N_12631,N_10612,N_11415);
or U12632 (N_12632,N_10555,N_11284);
nor U12633 (N_12633,N_10638,N_10614);
or U12634 (N_12634,N_11486,N_11670);
nor U12635 (N_12635,N_11481,N_10685);
and U12636 (N_12636,N_10878,N_10443);
and U12637 (N_12637,N_11439,N_10671);
and U12638 (N_12638,N_11648,N_11364);
xnor U12639 (N_12639,N_11786,N_11787);
and U12640 (N_12640,N_10544,N_11854);
or U12641 (N_12641,N_11763,N_10606);
xnor U12642 (N_12642,N_10433,N_10442);
nand U12643 (N_12643,N_10910,N_10078);
xnor U12644 (N_12644,N_11214,N_10811);
and U12645 (N_12645,N_11951,N_11352);
nor U12646 (N_12646,N_11402,N_10182);
and U12647 (N_12647,N_11418,N_10911);
xor U12648 (N_12648,N_10716,N_10719);
nand U12649 (N_12649,N_10139,N_11182);
nor U12650 (N_12650,N_11633,N_10468);
nor U12651 (N_12651,N_10534,N_11212);
and U12652 (N_12652,N_11296,N_11871);
and U12653 (N_12653,N_10772,N_11703);
xnor U12654 (N_12654,N_10170,N_11568);
nand U12655 (N_12655,N_10084,N_10185);
nor U12656 (N_12656,N_10870,N_11584);
and U12657 (N_12657,N_10929,N_11205);
nand U12658 (N_12658,N_10197,N_11446);
xor U12659 (N_12659,N_10990,N_11031);
and U12660 (N_12660,N_11845,N_10847);
nand U12661 (N_12661,N_11727,N_10066);
and U12662 (N_12662,N_10157,N_10330);
nand U12663 (N_12663,N_11156,N_10517);
nand U12664 (N_12664,N_11165,N_11176);
xnor U12665 (N_12665,N_10499,N_10234);
nand U12666 (N_12666,N_10819,N_11708);
or U12667 (N_12667,N_11270,N_10537);
xnor U12668 (N_12668,N_11029,N_11166);
nand U12669 (N_12669,N_11228,N_11409);
xnor U12670 (N_12670,N_11282,N_10123);
nor U12671 (N_12671,N_10776,N_11320);
nor U12672 (N_12672,N_11300,N_11234);
xnor U12673 (N_12673,N_11062,N_10333);
xnor U12674 (N_12674,N_11204,N_11998);
nand U12675 (N_12675,N_11883,N_11038);
or U12676 (N_12676,N_10619,N_10463);
nor U12677 (N_12677,N_11919,N_11315);
nor U12678 (N_12678,N_10645,N_10877);
and U12679 (N_12679,N_10211,N_11677);
xnor U12680 (N_12680,N_11964,N_10993);
nor U12681 (N_12681,N_11839,N_10486);
nor U12682 (N_12682,N_11476,N_11200);
xor U12683 (N_12683,N_11261,N_11135);
nor U12684 (N_12684,N_11575,N_10693);
and U12685 (N_12685,N_10802,N_10088);
xor U12686 (N_12686,N_11073,N_10530);
nand U12687 (N_12687,N_10564,N_11290);
and U12688 (N_12688,N_10844,N_11496);
xnor U12689 (N_12689,N_11869,N_10423);
and U12690 (N_12690,N_11293,N_10955);
or U12691 (N_12691,N_10764,N_10215);
xnor U12692 (N_12692,N_11225,N_10452);
nor U12693 (N_12693,N_11946,N_11118);
nand U12694 (N_12694,N_11685,N_10958);
and U12695 (N_12695,N_11725,N_11736);
nor U12696 (N_12696,N_10924,N_11766);
nor U12697 (N_12697,N_10893,N_11941);
and U12698 (N_12698,N_10542,N_11342);
nand U12699 (N_12699,N_10553,N_10767);
nor U12700 (N_12700,N_10018,N_10967);
xnor U12701 (N_12701,N_11283,N_11484);
nor U12702 (N_12702,N_11540,N_10817);
nor U12703 (N_12703,N_11822,N_10745);
and U12704 (N_12704,N_11675,N_10584);
or U12705 (N_12705,N_10744,N_10232);
and U12706 (N_12706,N_11526,N_11076);
xnor U12707 (N_12707,N_11504,N_10162);
nor U12708 (N_12708,N_10675,N_10891);
nand U12709 (N_12709,N_10648,N_11322);
or U12710 (N_12710,N_10134,N_11765);
nand U12711 (N_12711,N_10013,N_11757);
nor U12712 (N_12712,N_11407,N_10115);
xnor U12713 (N_12713,N_11358,N_10121);
or U12714 (N_12714,N_10996,N_11550);
or U12715 (N_12715,N_11285,N_10479);
nand U12716 (N_12716,N_10547,N_11841);
nor U12717 (N_12717,N_10235,N_11414);
and U12718 (N_12718,N_10472,N_11607);
nor U12719 (N_12719,N_10915,N_11865);
xnor U12720 (N_12720,N_11383,N_10747);
or U12721 (N_12721,N_10710,N_11922);
nand U12722 (N_12722,N_10966,N_10071);
and U12723 (N_12723,N_10294,N_10261);
and U12724 (N_12724,N_11011,N_11521);
nor U12725 (N_12725,N_10925,N_11975);
or U12726 (N_12726,N_11276,N_10323);
xnor U12727 (N_12727,N_11363,N_10588);
nor U12728 (N_12728,N_11049,N_10343);
xnor U12729 (N_12729,N_11799,N_10375);
and U12730 (N_12730,N_10244,N_11666);
or U12731 (N_12731,N_10680,N_11015);
nand U12732 (N_12732,N_10839,N_11425);
nand U12733 (N_12733,N_11586,N_10429);
nand U12734 (N_12734,N_11275,N_11744);
or U12735 (N_12735,N_11606,N_11112);
nand U12736 (N_12736,N_11849,N_10098);
or U12737 (N_12737,N_10216,N_10732);
and U12738 (N_12738,N_11229,N_11134);
and U12739 (N_12739,N_11160,N_11145);
or U12740 (N_12740,N_10998,N_10797);
nor U12741 (N_12741,N_10303,N_11902);
xor U12742 (N_12742,N_11499,N_10335);
xor U12743 (N_12743,N_10004,N_10622);
and U12744 (N_12744,N_10666,N_11855);
nor U12745 (N_12745,N_10815,N_11306);
nor U12746 (N_12746,N_10829,N_11523);
nand U12747 (N_12747,N_10331,N_11999);
nor U12748 (N_12748,N_11144,N_11566);
xor U12749 (N_12749,N_10975,N_11967);
nand U12750 (N_12750,N_10097,N_10380);
xnor U12751 (N_12751,N_11894,N_11199);
xor U12752 (N_12752,N_10324,N_10777);
xnor U12753 (N_12753,N_11087,N_10986);
nand U12754 (N_12754,N_10927,N_10508);
nor U12755 (N_12755,N_10198,N_10386);
or U12756 (N_12756,N_10790,N_11712);
and U12757 (N_12757,N_11410,N_11148);
and U12758 (N_12758,N_11464,N_11108);
and U12759 (N_12759,N_10809,N_11155);
xor U12760 (N_12760,N_11245,N_10382);
nor U12761 (N_12761,N_11808,N_11611);
xor U12762 (N_12762,N_10668,N_10730);
nand U12763 (N_12763,N_11404,N_11437);
or U12764 (N_12764,N_10210,N_10256);
and U12765 (N_12765,N_10410,N_10932);
nand U12766 (N_12766,N_10649,N_10905);
or U12767 (N_12767,N_10319,N_10440);
nor U12768 (N_12768,N_11468,N_10803);
and U12769 (N_12769,N_11638,N_11000);
nor U12770 (N_12770,N_10717,N_10848);
xnor U12771 (N_12771,N_11419,N_10133);
and U12772 (N_12772,N_11548,N_10495);
xnor U12773 (N_12773,N_11377,N_11203);
nand U12774 (N_12774,N_10843,N_11749);
or U12775 (N_12775,N_11325,N_11444);
nand U12776 (N_12776,N_11427,N_11524);
nand U12777 (N_12777,N_11391,N_11660);
nor U12778 (N_12778,N_11001,N_11528);
nor U12779 (N_12779,N_11077,N_11530);
or U12780 (N_12780,N_11054,N_10785);
nand U12781 (N_12781,N_11180,N_10173);
and U12782 (N_12782,N_10921,N_11859);
nor U12783 (N_12783,N_10262,N_10629);
nor U12784 (N_12784,N_10069,N_10146);
or U12785 (N_12785,N_11309,N_10190);
and U12786 (N_12786,N_11447,N_11507);
or U12787 (N_12787,N_10238,N_10823);
xnor U12788 (N_12788,N_11860,N_10199);
nand U12789 (N_12789,N_10344,N_11664);
and U12790 (N_12790,N_10204,N_10739);
nand U12791 (N_12791,N_11079,N_10726);
nand U12792 (N_12792,N_10887,N_10864);
and U12793 (N_12793,N_10590,N_11201);
xor U12794 (N_12794,N_10841,N_11268);
or U12795 (N_12795,N_11051,N_11009);
nor U12796 (N_12796,N_10259,N_11731);
nand U12797 (N_12797,N_10404,N_11151);
xnor U12798 (N_12798,N_10161,N_10281);
or U12799 (N_12799,N_10883,N_10048);
xnor U12800 (N_12800,N_11917,N_11189);
and U12801 (N_12801,N_11511,N_11022);
or U12802 (N_12802,N_11477,N_11867);
xnor U12803 (N_12803,N_10193,N_11299);
nand U12804 (N_12804,N_11752,N_10798);
nor U12805 (N_12805,N_10830,N_11544);
or U12806 (N_12806,N_10041,N_10519);
or U12807 (N_12807,N_10462,N_11475);
xor U12808 (N_12808,N_10307,N_11512);
xnor U12809 (N_12809,N_11289,N_11829);
nor U12810 (N_12810,N_10703,N_11745);
xor U12811 (N_12811,N_11480,N_10138);
or U12812 (N_12812,N_11012,N_11354);
and U12813 (N_12813,N_11240,N_10007);
nor U12814 (N_12814,N_11811,N_10709);
xor U12815 (N_12815,N_11382,N_11662);
nand U12816 (N_12816,N_10930,N_11687);
nor U12817 (N_12817,N_10746,N_11656);
nand U12818 (N_12818,N_10778,N_11623);
xnor U12819 (N_12819,N_10628,N_10247);
xor U12820 (N_12820,N_10484,N_11931);
nor U12821 (N_12821,N_10010,N_10763);
xor U12822 (N_12822,N_11886,N_10180);
xor U12823 (N_12823,N_11105,N_11823);
and U12824 (N_12824,N_11059,N_10653);
or U12825 (N_12825,N_11657,N_10660);
or U12826 (N_12826,N_11683,N_11713);
nand U12827 (N_12827,N_11164,N_11570);
and U12828 (N_12828,N_11061,N_10851);
nor U12829 (N_12829,N_10081,N_11192);
nand U12830 (N_12830,N_11041,N_11263);
and U12831 (N_12831,N_11150,N_11196);
and U12832 (N_12832,N_10159,N_11816);
or U12833 (N_12833,N_11198,N_10196);
nor U12834 (N_12834,N_10824,N_10299);
nor U12835 (N_12835,N_11197,N_10690);
nor U12836 (N_12836,N_10945,N_11676);
xor U12837 (N_12837,N_10497,N_11351);
nor U12838 (N_12838,N_11307,N_10045);
nor U12839 (N_12839,N_11806,N_11006);
xor U12840 (N_12840,N_10632,N_11746);
nand U12841 (N_12841,N_10076,N_11399);
xnor U12842 (N_12842,N_10308,N_11564);
xnor U12843 (N_12843,N_11608,N_11017);
nor U12844 (N_12844,N_11256,N_11850);
or U12845 (N_12845,N_10301,N_11988);
and U12846 (N_12846,N_10513,N_10111);
or U12847 (N_12847,N_11881,N_11851);
nand U12848 (N_12848,N_10009,N_10518);
and U12849 (N_12849,N_10899,N_10061);
or U12850 (N_12850,N_11123,N_10432);
nor U12851 (N_12851,N_10223,N_11949);
xor U12852 (N_12852,N_11569,N_11474);
and U12853 (N_12853,N_10387,N_10059);
and U12854 (N_12854,N_10603,N_10655);
and U12855 (N_12855,N_11642,N_10322);
and U12856 (N_12856,N_11977,N_10867);
nor U12857 (N_12857,N_11210,N_10702);
nor U12858 (N_12858,N_11143,N_10999);
nor U12859 (N_12859,N_10748,N_11337);
xnor U12860 (N_12860,N_11302,N_11652);
xnor U12861 (N_12861,N_10365,N_11597);
nor U12862 (N_12862,N_10657,N_10593);
and U12863 (N_12863,N_10315,N_10471);
and U12864 (N_12864,N_11793,N_11843);
nand U12865 (N_12865,N_10721,N_11327);
nor U12866 (N_12866,N_11965,N_11104);
xnor U12867 (N_12867,N_10742,N_10595);
or U12868 (N_12868,N_11467,N_11280);
or U12869 (N_12869,N_11202,N_10831);
and U12870 (N_12870,N_11921,N_10775);
and U12871 (N_12871,N_10203,N_11190);
or U12872 (N_12872,N_11927,N_11131);
nand U12873 (N_12873,N_10756,N_10581);
and U12874 (N_12874,N_10749,N_10288);
and U12875 (N_12875,N_11273,N_10436);
or U12876 (N_12876,N_11435,N_11995);
and U12877 (N_12877,N_11065,N_10669);
or U12878 (N_12878,N_11375,N_10750);
and U12879 (N_12879,N_10029,N_11096);
nand U12880 (N_12880,N_10340,N_11546);
or U12881 (N_12881,N_10413,N_11748);
nand U12882 (N_12882,N_11016,N_11899);
nor U12883 (N_12883,N_11436,N_11788);
or U12884 (N_12884,N_10642,N_11116);
and U12885 (N_12885,N_10656,N_10230);
nor U12886 (N_12886,N_10225,N_10515);
nand U12887 (N_12887,N_11776,N_11287);
nand U12888 (N_12888,N_11707,N_10407);
nand U12889 (N_12889,N_11785,N_11024);
xor U12890 (N_12890,N_11595,N_10126);
nor U12891 (N_12891,N_11373,N_11100);
and U12892 (N_12892,N_11219,N_10973);
nand U12893 (N_12893,N_11803,N_10757);
nor U12894 (N_12894,N_11649,N_11430);
nand U12895 (N_12895,N_10090,N_10863);
and U12896 (N_12896,N_10902,N_11395);
nand U12897 (N_12897,N_11936,N_11690);
nor U12898 (N_12898,N_10801,N_10431);
xor U12899 (N_12899,N_11432,N_11120);
nand U12900 (N_12900,N_11211,N_11050);
xnor U12901 (N_12901,N_11579,N_11422);
or U12902 (N_12902,N_11824,N_10352);
nand U12903 (N_12903,N_10311,N_11317);
nand U12904 (N_12904,N_10968,N_11122);
and U12905 (N_12905,N_11465,N_11085);
xnor U12906 (N_12906,N_10874,N_10970);
nor U12907 (N_12907,N_10033,N_11628);
or U12908 (N_12908,N_10467,N_10912);
nand U12909 (N_12909,N_10791,N_11543);
xnor U12910 (N_12910,N_11934,N_10804);
nor U12911 (N_12911,N_11655,N_11783);
xor U12912 (N_12912,N_10977,N_11115);
nand U12913 (N_12913,N_10740,N_11241);
or U12914 (N_12914,N_11701,N_10822);
nor U12915 (N_12915,N_11335,N_11955);
nand U12916 (N_12916,N_10880,N_10163);
and U12917 (N_12917,N_10974,N_10118);
nor U12918 (N_12918,N_10260,N_11459);
nor U12919 (N_12919,N_10868,N_10865);
or U12920 (N_12920,N_11990,N_10901);
nand U12921 (N_12921,N_10913,N_11605);
and U12922 (N_12922,N_10694,N_11583);
nor U12923 (N_12923,N_10597,N_10325);
or U12924 (N_12924,N_10267,N_10001);
or U12925 (N_12925,N_11689,N_11828);
and U12926 (N_12926,N_11549,N_10741);
nand U12927 (N_12927,N_11728,N_10306);
nand U12928 (N_12928,N_11705,N_11042);
nor U12929 (N_12929,N_10339,N_11357);
nand U12930 (N_12930,N_10850,N_11613);
and U12931 (N_12931,N_10808,N_11493);
nand U12932 (N_12932,N_10444,N_10187);
nand U12933 (N_12933,N_10304,N_11514);
and U12934 (N_12934,N_10480,N_10152);
nor U12935 (N_12935,N_11455,N_10342);
xor U12936 (N_12936,N_11796,N_11348);
xnor U12937 (N_12937,N_10248,N_10722);
and U12938 (N_12938,N_10569,N_10641);
nand U12939 (N_12939,N_11389,N_10633);
nand U12940 (N_12940,N_11582,N_11950);
nand U12941 (N_12941,N_11598,N_11891);
and U12942 (N_12942,N_11780,N_10255);
nor U12943 (N_12943,N_11277,N_10988);
and U12944 (N_12944,N_10136,N_11044);
nand U12945 (N_12945,N_10609,N_10280);
nor U12946 (N_12946,N_11020,N_11128);
or U12947 (N_12947,N_11416,N_10787);
nor U12948 (N_12948,N_11906,N_11866);
xnor U12949 (N_12949,N_11491,N_11035);
xnor U12950 (N_12950,N_11216,N_10684);
nand U12951 (N_12951,N_11326,N_10926);
and U12952 (N_12952,N_11837,N_10017);
nor U12953 (N_12953,N_10057,N_10964);
nand U12954 (N_12954,N_11440,N_11119);
nor U12955 (N_12955,N_11971,N_11996);
nor U12956 (N_12956,N_11527,N_10794);
or U12957 (N_12957,N_10689,N_10523);
xnor U12958 (N_12958,N_11344,N_10607);
nand U12959 (N_12959,N_10728,N_11369);
nand U12960 (N_12960,N_10142,N_11928);
xor U12961 (N_12961,N_10736,N_11735);
and U12962 (N_12962,N_11875,N_10972);
or U12963 (N_12963,N_11695,N_11226);
xnor U12964 (N_12964,N_10989,N_10242);
or U12965 (N_12965,N_11518,N_10526);
and U12966 (N_12966,N_11479,N_11903);
or U12967 (N_12967,N_11522,N_10567);
nand U12968 (N_12968,N_11400,N_11533);
nand U12969 (N_12969,N_10273,N_11813);
nor U12970 (N_12970,N_10362,N_11187);
or U12971 (N_12971,N_10285,N_11663);
or U12972 (N_12972,N_11194,N_10400);
or U12973 (N_12973,N_10725,N_10494);
nor U12974 (N_12974,N_11693,N_10075);
and U12975 (N_12975,N_11502,N_10414);
xnor U12976 (N_12976,N_10347,N_10109);
or U12977 (N_12977,N_10409,N_11498);
or U12978 (N_12978,N_11935,N_10231);
nand U12979 (N_12979,N_10601,N_11174);
and U12980 (N_12980,N_10283,N_11698);
or U12981 (N_12981,N_10483,N_10295);
xnor U12982 (N_12982,N_11365,N_11221);
nand U12983 (N_12983,N_11890,N_11500);
and U12984 (N_12984,N_10509,N_11460);
xor U12985 (N_12985,N_11966,N_10056);
xor U12986 (N_12986,N_10373,N_11441);
nand U12987 (N_12987,N_11298,N_10853);
nor U12988 (N_12988,N_10458,N_10589);
xnor U12989 (N_12989,N_10783,N_10541);
or U12990 (N_12990,N_10545,N_10450);
and U12991 (N_12991,N_11770,N_10565);
xnor U12992 (N_12992,N_11503,N_11567);
and U12993 (N_12993,N_10408,N_11726);
and U12994 (N_12994,N_10006,N_10909);
or U12995 (N_12995,N_11209,N_11658);
nand U12996 (N_12996,N_11332,N_11840);
nor U12997 (N_12997,N_11314,N_10723);
nor U12998 (N_12998,N_10272,N_11742);
and U12999 (N_12999,N_10477,N_10837);
nor U13000 (N_13000,N_10312,N_10359);
or U13001 (N_13001,N_11161,N_11989);
and U13002 (N_13002,N_11896,N_10257);
xnor U13003 (N_13003,N_11200,N_10392);
nand U13004 (N_13004,N_10609,N_10675);
xor U13005 (N_13005,N_11677,N_11013);
or U13006 (N_13006,N_11209,N_11347);
or U13007 (N_13007,N_10304,N_10588);
nor U13008 (N_13008,N_10359,N_10349);
nor U13009 (N_13009,N_10493,N_11039);
nand U13010 (N_13010,N_11509,N_10395);
xnor U13011 (N_13011,N_11931,N_10170);
nand U13012 (N_13012,N_11341,N_11721);
xnor U13013 (N_13013,N_10266,N_11948);
or U13014 (N_13014,N_11782,N_10709);
and U13015 (N_13015,N_11359,N_10705);
nand U13016 (N_13016,N_10741,N_10583);
and U13017 (N_13017,N_10886,N_10276);
nand U13018 (N_13018,N_11266,N_10098);
nor U13019 (N_13019,N_11973,N_10002);
or U13020 (N_13020,N_10145,N_10581);
xor U13021 (N_13021,N_11781,N_11816);
and U13022 (N_13022,N_10060,N_11072);
nand U13023 (N_13023,N_10111,N_10534);
nand U13024 (N_13024,N_11531,N_11342);
or U13025 (N_13025,N_11802,N_10952);
and U13026 (N_13026,N_10426,N_10604);
xnor U13027 (N_13027,N_11068,N_11604);
nor U13028 (N_13028,N_10024,N_10494);
xnor U13029 (N_13029,N_11527,N_10102);
nand U13030 (N_13030,N_10473,N_11155);
nand U13031 (N_13031,N_10918,N_10857);
nor U13032 (N_13032,N_11271,N_11239);
nand U13033 (N_13033,N_11571,N_10980);
nand U13034 (N_13034,N_11424,N_11804);
xnor U13035 (N_13035,N_10243,N_11409);
nand U13036 (N_13036,N_11358,N_10822);
nand U13037 (N_13037,N_10840,N_10715);
nand U13038 (N_13038,N_11395,N_10435);
nor U13039 (N_13039,N_11275,N_11645);
nand U13040 (N_13040,N_10975,N_10399);
or U13041 (N_13041,N_10839,N_10556);
nor U13042 (N_13042,N_10522,N_11744);
xor U13043 (N_13043,N_11587,N_10858);
and U13044 (N_13044,N_11361,N_10149);
and U13045 (N_13045,N_10676,N_10746);
nand U13046 (N_13046,N_10315,N_10158);
nand U13047 (N_13047,N_11689,N_11365);
nor U13048 (N_13048,N_10103,N_10741);
nor U13049 (N_13049,N_10362,N_10627);
nor U13050 (N_13050,N_10064,N_11179);
nand U13051 (N_13051,N_10561,N_11480);
nor U13052 (N_13052,N_10129,N_10052);
nand U13053 (N_13053,N_11267,N_10587);
nand U13054 (N_13054,N_10355,N_11203);
nor U13055 (N_13055,N_11765,N_11311);
nor U13056 (N_13056,N_11692,N_11104);
nand U13057 (N_13057,N_11292,N_10026);
xor U13058 (N_13058,N_11961,N_10527);
nand U13059 (N_13059,N_10696,N_10839);
nor U13060 (N_13060,N_10519,N_11803);
or U13061 (N_13061,N_11311,N_11186);
xnor U13062 (N_13062,N_10930,N_11357);
and U13063 (N_13063,N_11619,N_10047);
nor U13064 (N_13064,N_10406,N_11244);
and U13065 (N_13065,N_10493,N_10169);
xnor U13066 (N_13066,N_11113,N_10854);
nor U13067 (N_13067,N_11295,N_11836);
and U13068 (N_13068,N_10248,N_10850);
nand U13069 (N_13069,N_10605,N_11457);
nand U13070 (N_13070,N_10470,N_11122);
xnor U13071 (N_13071,N_11981,N_10305);
nor U13072 (N_13072,N_11322,N_10934);
or U13073 (N_13073,N_11632,N_10704);
nor U13074 (N_13074,N_10877,N_11954);
and U13075 (N_13075,N_11178,N_11003);
or U13076 (N_13076,N_10077,N_10398);
xnor U13077 (N_13077,N_10060,N_10606);
and U13078 (N_13078,N_11128,N_11695);
and U13079 (N_13079,N_11569,N_11458);
xnor U13080 (N_13080,N_10026,N_10556);
or U13081 (N_13081,N_11012,N_11620);
nor U13082 (N_13082,N_11592,N_11254);
and U13083 (N_13083,N_11637,N_10035);
nand U13084 (N_13084,N_10003,N_10219);
nor U13085 (N_13085,N_11069,N_11339);
nand U13086 (N_13086,N_10871,N_11181);
and U13087 (N_13087,N_11887,N_11413);
and U13088 (N_13088,N_11331,N_10088);
and U13089 (N_13089,N_10705,N_11586);
nand U13090 (N_13090,N_11265,N_10122);
xnor U13091 (N_13091,N_10104,N_10640);
and U13092 (N_13092,N_11693,N_10195);
or U13093 (N_13093,N_10989,N_10045);
nor U13094 (N_13094,N_11757,N_11758);
and U13095 (N_13095,N_10439,N_11150);
or U13096 (N_13096,N_11581,N_11777);
nand U13097 (N_13097,N_11229,N_10335);
nand U13098 (N_13098,N_10422,N_11702);
nand U13099 (N_13099,N_10918,N_10169);
nor U13100 (N_13100,N_10075,N_11073);
or U13101 (N_13101,N_11594,N_10049);
or U13102 (N_13102,N_10600,N_10041);
nor U13103 (N_13103,N_10812,N_10755);
nor U13104 (N_13104,N_10988,N_11685);
nand U13105 (N_13105,N_11094,N_11426);
nor U13106 (N_13106,N_11545,N_10071);
xnor U13107 (N_13107,N_11723,N_11052);
xnor U13108 (N_13108,N_10299,N_11280);
and U13109 (N_13109,N_10475,N_10784);
nor U13110 (N_13110,N_11260,N_10411);
xnor U13111 (N_13111,N_10705,N_10952);
or U13112 (N_13112,N_11326,N_10942);
and U13113 (N_13113,N_11562,N_10242);
or U13114 (N_13114,N_10849,N_11081);
and U13115 (N_13115,N_11235,N_10476);
or U13116 (N_13116,N_10497,N_11717);
and U13117 (N_13117,N_10347,N_10372);
nand U13118 (N_13118,N_10484,N_10203);
nor U13119 (N_13119,N_11038,N_11903);
or U13120 (N_13120,N_10997,N_11905);
xnor U13121 (N_13121,N_11555,N_10018);
and U13122 (N_13122,N_10322,N_11389);
nand U13123 (N_13123,N_10424,N_10368);
nor U13124 (N_13124,N_11634,N_11640);
xor U13125 (N_13125,N_10224,N_11245);
or U13126 (N_13126,N_10332,N_10166);
nor U13127 (N_13127,N_10867,N_10862);
and U13128 (N_13128,N_10205,N_11197);
nand U13129 (N_13129,N_11712,N_11322);
nor U13130 (N_13130,N_11939,N_11841);
or U13131 (N_13131,N_11608,N_11962);
nand U13132 (N_13132,N_10847,N_11545);
nand U13133 (N_13133,N_11993,N_11756);
xnor U13134 (N_13134,N_10762,N_11058);
nand U13135 (N_13135,N_10689,N_11249);
nand U13136 (N_13136,N_10942,N_10243);
and U13137 (N_13137,N_10825,N_10838);
or U13138 (N_13138,N_11402,N_10248);
or U13139 (N_13139,N_11097,N_11186);
nand U13140 (N_13140,N_10694,N_10705);
or U13141 (N_13141,N_10900,N_10109);
or U13142 (N_13142,N_11847,N_10004);
and U13143 (N_13143,N_10021,N_11674);
nor U13144 (N_13144,N_10998,N_10780);
xor U13145 (N_13145,N_10550,N_11472);
and U13146 (N_13146,N_11923,N_10510);
nand U13147 (N_13147,N_10099,N_10629);
and U13148 (N_13148,N_11127,N_11736);
and U13149 (N_13149,N_10448,N_10764);
nand U13150 (N_13150,N_11495,N_11773);
xnor U13151 (N_13151,N_11391,N_11214);
xnor U13152 (N_13152,N_10595,N_11352);
or U13153 (N_13153,N_10696,N_11259);
and U13154 (N_13154,N_10333,N_10267);
xor U13155 (N_13155,N_10466,N_10656);
xnor U13156 (N_13156,N_11534,N_11853);
nand U13157 (N_13157,N_10506,N_10433);
nand U13158 (N_13158,N_11783,N_11065);
nor U13159 (N_13159,N_10295,N_10213);
nand U13160 (N_13160,N_10087,N_10147);
nor U13161 (N_13161,N_10578,N_11668);
nor U13162 (N_13162,N_11792,N_10474);
and U13163 (N_13163,N_11206,N_10909);
and U13164 (N_13164,N_10714,N_11248);
and U13165 (N_13165,N_10966,N_10166);
nor U13166 (N_13166,N_11370,N_11391);
and U13167 (N_13167,N_11082,N_11629);
and U13168 (N_13168,N_10522,N_11279);
or U13169 (N_13169,N_10045,N_10222);
nand U13170 (N_13170,N_11415,N_11358);
or U13171 (N_13171,N_11533,N_10785);
nor U13172 (N_13172,N_11623,N_11333);
nand U13173 (N_13173,N_10748,N_10534);
nor U13174 (N_13174,N_11085,N_10317);
nor U13175 (N_13175,N_11647,N_10158);
and U13176 (N_13176,N_11344,N_11887);
nor U13177 (N_13177,N_10483,N_10811);
nor U13178 (N_13178,N_11457,N_10937);
or U13179 (N_13179,N_10801,N_10148);
xnor U13180 (N_13180,N_11413,N_10969);
and U13181 (N_13181,N_10505,N_11103);
xnor U13182 (N_13182,N_11291,N_10405);
nor U13183 (N_13183,N_10401,N_11486);
and U13184 (N_13184,N_10266,N_11119);
nand U13185 (N_13185,N_11893,N_11374);
nand U13186 (N_13186,N_10174,N_10855);
nand U13187 (N_13187,N_11986,N_10893);
nor U13188 (N_13188,N_10229,N_11667);
and U13189 (N_13189,N_11611,N_11794);
xnor U13190 (N_13190,N_11411,N_10092);
and U13191 (N_13191,N_10367,N_11565);
nand U13192 (N_13192,N_10204,N_10141);
nand U13193 (N_13193,N_10225,N_10045);
or U13194 (N_13194,N_10280,N_11041);
nor U13195 (N_13195,N_10927,N_10534);
nand U13196 (N_13196,N_11352,N_10196);
or U13197 (N_13197,N_11794,N_10704);
nor U13198 (N_13198,N_11501,N_10756);
nand U13199 (N_13199,N_10044,N_11606);
or U13200 (N_13200,N_11946,N_11092);
nor U13201 (N_13201,N_11309,N_11858);
nand U13202 (N_13202,N_10447,N_10538);
or U13203 (N_13203,N_10358,N_10733);
xor U13204 (N_13204,N_11831,N_11533);
xnor U13205 (N_13205,N_10475,N_10994);
nand U13206 (N_13206,N_11056,N_10383);
xnor U13207 (N_13207,N_11243,N_11055);
and U13208 (N_13208,N_10505,N_10803);
or U13209 (N_13209,N_11723,N_11885);
and U13210 (N_13210,N_11217,N_10377);
nand U13211 (N_13211,N_11369,N_11850);
nand U13212 (N_13212,N_10499,N_10909);
nand U13213 (N_13213,N_11990,N_10108);
xnor U13214 (N_13214,N_10159,N_11948);
and U13215 (N_13215,N_11230,N_11356);
nor U13216 (N_13216,N_11321,N_10744);
nor U13217 (N_13217,N_11906,N_11167);
nand U13218 (N_13218,N_10176,N_11553);
and U13219 (N_13219,N_10923,N_11209);
or U13220 (N_13220,N_11487,N_11482);
nand U13221 (N_13221,N_10873,N_10807);
nand U13222 (N_13222,N_10777,N_10044);
xor U13223 (N_13223,N_11645,N_11582);
and U13224 (N_13224,N_10063,N_11598);
xnor U13225 (N_13225,N_11841,N_11711);
nor U13226 (N_13226,N_11849,N_10978);
or U13227 (N_13227,N_11235,N_10125);
nor U13228 (N_13228,N_10535,N_11866);
and U13229 (N_13229,N_10265,N_10159);
and U13230 (N_13230,N_11170,N_10140);
or U13231 (N_13231,N_10964,N_10406);
xor U13232 (N_13232,N_11950,N_11107);
or U13233 (N_13233,N_10849,N_10603);
nand U13234 (N_13234,N_10745,N_11634);
and U13235 (N_13235,N_10653,N_10502);
nand U13236 (N_13236,N_10388,N_11755);
and U13237 (N_13237,N_10061,N_11002);
and U13238 (N_13238,N_10153,N_11254);
or U13239 (N_13239,N_11238,N_11716);
nor U13240 (N_13240,N_11511,N_11507);
nor U13241 (N_13241,N_10673,N_10962);
xnor U13242 (N_13242,N_11638,N_10892);
nand U13243 (N_13243,N_11283,N_10204);
and U13244 (N_13244,N_11425,N_11432);
and U13245 (N_13245,N_10993,N_11518);
nor U13246 (N_13246,N_10409,N_10936);
nor U13247 (N_13247,N_10572,N_10891);
xnor U13248 (N_13248,N_11873,N_11269);
and U13249 (N_13249,N_11288,N_10096);
xnor U13250 (N_13250,N_10428,N_10182);
or U13251 (N_13251,N_10060,N_11275);
nand U13252 (N_13252,N_11996,N_11751);
nor U13253 (N_13253,N_11456,N_11376);
xor U13254 (N_13254,N_11210,N_10902);
nand U13255 (N_13255,N_10505,N_11899);
or U13256 (N_13256,N_10983,N_11055);
nand U13257 (N_13257,N_11462,N_11530);
and U13258 (N_13258,N_10586,N_10832);
or U13259 (N_13259,N_11008,N_11548);
or U13260 (N_13260,N_10637,N_10841);
and U13261 (N_13261,N_10334,N_10084);
xnor U13262 (N_13262,N_11586,N_11831);
nor U13263 (N_13263,N_10896,N_11171);
nor U13264 (N_13264,N_11870,N_10374);
xnor U13265 (N_13265,N_10746,N_10657);
xor U13266 (N_13266,N_10172,N_10774);
and U13267 (N_13267,N_11994,N_11491);
xnor U13268 (N_13268,N_11518,N_11100);
nand U13269 (N_13269,N_11700,N_11318);
nor U13270 (N_13270,N_10734,N_10025);
nor U13271 (N_13271,N_10149,N_11314);
nor U13272 (N_13272,N_11193,N_11693);
nor U13273 (N_13273,N_11445,N_11182);
xor U13274 (N_13274,N_10438,N_11817);
xor U13275 (N_13275,N_10238,N_11687);
and U13276 (N_13276,N_11210,N_10395);
and U13277 (N_13277,N_11288,N_11686);
nor U13278 (N_13278,N_11205,N_10946);
xor U13279 (N_13279,N_10893,N_10453);
and U13280 (N_13280,N_11443,N_10758);
xnor U13281 (N_13281,N_11841,N_11022);
nor U13282 (N_13282,N_11381,N_11104);
and U13283 (N_13283,N_11723,N_11933);
and U13284 (N_13284,N_11079,N_10127);
and U13285 (N_13285,N_11635,N_10391);
nand U13286 (N_13286,N_10467,N_10757);
nand U13287 (N_13287,N_11235,N_11191);
nand U13288 (N_13288,N_11107,N_11579);
xnor U13289 (N_13289,N_10144,N_10071);
nand U13290 (N_13290,N_10717,N_10676);
nor U13291 (N_13291,N_11121,N_10007);
xnor U13292 (N_13292,N_11418,N_10201);
xnor U13293 (N_13293,N_11867,N_11321);
and U13294 (N_13294,N_11974,N_10314);
and U13295 (N_13295,N_11699,N_11854);
nand U13296 (N_13296,N_10354,N_10202);
and U13297 (N_13297,N_11125,N_10210);
and U13298 (N_13298,N_10312,N_11174);
nor U13299 (N_13299,N_11461,N_11043);
nor U13300 (N_13300,N_10755,N_11727);
and U13301 (N_13301,N_10632,N_11036);
nor U13302 (N_13302,N_10973,N_11110);
nand U13303 (N_13303,N_10116,N_11559);
or U13304 (N_13304,N_10144,N_10198);
nor U13305 (N_13305,N_10265,N_11790);
nand U13306 (N_13306,N_10213,N_10207);
nand U13307 (N_13307,N_10405,N_10237);
or U13308 (N_13308,N_11075,N_11011);
nand U13309 (N_13309,N_10580,N_10192);
nor U13310 (N_13310,N_11468,N_11756);
xor U13311 (N_13311,N_10030,N_10903);
nand U13312 (N_13312,N_10266,N_11717);
and U13313 (N_13313,N_10784,N_11771);
or U13314 (N_13314,N_11629,N_10564);
nor U13315 (N_13315,N_11248,N_10485);
nor U13316 (N_13316,N_11464,N_11958);
nor U13317 (N_13317,N_10518,N_10882);
xor U13318 (N_13318,N_11346,N_11667);
nand U13319 (N_13319,N_11592,N_11739);
and U13320 (N_13320,N_11722,N_10610);
xor U13321 (N_13321,N_11546,N_10148);
nand U13322 (N_13322,N_10627,N_10920);
or U13323 (N_13323,N_10338,N_11989);
nand U13324 (N_13324,N_10248,N_10319);
nor U13325 (N_13325,N_11830,N_11391);
nor U13326 (N_13326,N_10817,N_10494);
nor U13327 (N_13327,N_11675,N_11777);
or U13328 (N_13328,N_11167,N_11697);
xor U13329 (N_13329,N_11392,N_11306);
nand U13330 (N_13330,N_11730,N_10462);
nor U13331 (N_13331,N_11064,N_10251);
xnor U13332 (N_13332,N_11091,N_11831);
xnor U13333 (N_13333,N_10649,N_11869);
nor U13334 (N_13334,N_11470,N_11923);
nand U13335 (N_13335,N_10048,N_11341);
nand U13336 (N_13336,N_11709,N_11714);
and U13337 (N_13337,N_11544,N_11951);
xor U13338 (N_13338,N_10670,N_10390);
xor U13339 (N_13339,N_10923,N_11112);
and U13340 (N_13340,N_11021,N_10938);
and U13341 (N_13341,N_11939,N_11242);
nor U13342 (N_13342,N_11876,N_11580);
and U13343 (N_13343,N_10250,N_10098);
xnor U13344 (N_13344,N_11595,N_11100);
nor U13345 (N_13345,N_11732,N_11099);
nand U13346 (N_13346,N_10537,N_11741);
or U13347 (N_13347,N_10439,N_11979);
nand U13348 (N_13348,N_10892,N_11531);
or U13349 (N_13349,N_10172,N_11428);
and U13350 (N_13350,N_10144,N_11151);
or U13351 (N_13351,N_10254,N_11818);
nor U13352 (N_13352,N_10399,N_11289);
xor U13353 (N_13353,N_11850,N_11675);
xor U13354 (N_13354,N_10883,N_11210);
nor U13355 (N_13355,N_11979,N_10556);
nand U13356 (N_13356,N_10858,N_10241);
and U13357 (N_13357,N_11820,N_10851);
nor U13358 (N_13358,N_10733,N_11179);
or U13359 (N_13359,N_11352,N_11970);
nand U13360 (N_13360,N_11294,N_10930);
nor U13361 (N_13361,N_11437,N_10125);
nand U13362 (N_13362,N_11369,N_10853);
nand U13363 (N_13363,N_10615,N_10372);
xor U13364 (N_13364,N_10985,N_11449);
xnor U13365 (N_13365,N_10466,N_10897);
and U13366 (N_13366,N_10400,N_11552);
nor U13367 (N_13367,N_10763,N_11596);
nand U13368 (N_13368,N_11851,N_11924);
or U13369 (N_13369,N_11924,N_11610);
or U13370 (N_13370,N_11366,N_11579);
or U13371 (N_13371,N_10298,N_10241);
nor U13372 (N_13372,N_11687,N_10089);
and U13373 (N_13373,N_11842,N_10969);
nand U13374 (N_13374,N_11909,N_10287);
xor U13375 (N_13375,N_11241,N_10217);
nand U13376 (N_13376,N_11846,N_11908);
and U13377 (N_13377,N_10564,N_11540);
nand U13378 (N_13378,N_10487,N_11565);
xor U13379 (N_13379,N_11452,N_10629);
nor U13380 (N_13380,N_10568,N_11046);
xnor U13381 (N_13381,N_11036,N_10368);
or U13382 (N_13382,N_10498,N_10354);
xnor U13383 (N_13383,N_11657,N_11730);
or U13384 (N_13384,N_10468,N_11922);
or U13385 (N_13385,N_10805,N_11844);
nor U13386 (N_13386,N_11222,N_10812);
or U13387 (N_13387,N_11349,N_11329);
and U13388 (N_13388,N_11062,N_10495);
nor U13389 (N_13389,N_10651,N_11963);
nor U13390 (N_13390,N_11212,N_10814);
and U13391 (N_13391,N_10235,N_10284);
nor U13392 (N_13392,N_10900,N_11960);
nor U13393 (N_13393,N_10318,N_11746);
or U13394 (N_13394,N_11872,N_11092);
or U13395 (N_13395,N_11479,N_10467);
nor U13396 (N_13396,N_11818,N_11205);
or U13397 (N_13397,N_11496,N_10978);
nor U13398 (N_13398,N_11818,N_10875);
and U13399 (N_13399,N_10861,N_11846);
nor U13400 (N_13400,N_10110,N_11747);
nor U13401 (N_13401,N_11268,N_10070);
xor U13402 (N_13402,N_10116,N_10205);
nand U13403 (N_13403,N_10638,N_11295);
and U13404 (N_13404,N_10447,N_11820);
nor U13405 (N_13405,N_10354,N_11601);
xnor U13406 (N_13406,N_11844,N_11551);
xnor U13407 (N_13407,N_10317,N_11426);
nand U13408 (N_13408,N_11356,N_10065);
nand U13409 (N_13409,N_10626,N_11800);
or U13410 (N_13410,N_11036,N_10847);
and U13411 (N_13411,N_11726,N_10936);
xor U13412 (N_13412,N_10547,N_10596);
or U13413 (N_13413,N_10057,N_11405);
nor U13414 (N_13414,N_10404,N_11457);
nor U13415 (N_13415,N_11527,N_11277);
nor U13416 (N_13416,N_11392,N_11348);
and U13417 (N_13417,N_10022,N_11729);
xor U13418 (N_13418,N_11882,N_10393);
and U13419 (N_13419,N_10046,N_10676);
nand U13420 (N_13420,N_10839,N_10508);
nor U13421 (N_13421,N_11128,N_11660);
or U13422 (N_13422,N_11248,N_11385);
nor U13423 (N_13423,N_11232,N_11093);
xor U13424 (N_13424,N_11333,N_11610);
nand U13425 (N_13425,N_10455,N_10266);
xnor U13426 (N_13426,N_10453,N_11170);
or U13427 (N_13427,N_10481,N_10470);
or U13428 (N_13428,N_11445,N_10654);
nand U13429 (N_13429,N_10576,N_10905);
nand U13430 (N_13430,N_10359,N_10108);
or U13431 (N_13431,N_11543,N_11575);
nand U13432 (N_13432,N_11827,N_10542);
xnor U13433 (N_13433,N_10885,N_11514);
xor U13434 (N_13434,N_11336,N_11438);
nor U13435 (N_13435,N_11609,N_10778);
or U13436 (N_13436,N_11954,N_10466);
nor U13437 (N_13437,N_11484,N_10577);
nand U13438 (N_13438,N_11361,N_11523);
and U13439 (N_13439,N_10164,N_11409);
xor U13440 (N_13440,N_10615,N_11407);
or U13441 (N_13441,N_10922,N_10122);
or U13442 (N_13442,N_11200,N_11428);
nand U13443 (N_13443,N_10559,N_10006);
xor U13444 (N_13444,N_10434,N_10492);
and U13445 (N_13445,N_10874,N_11342);
xor U13446 (N_13446,N_10487,N_11153);
nor U13447 (N_13447,N_11207,N_11619);
nor U13448 (N_13448,N_10436,N_10974);
and U13449 (N_13449,N_10880,N_11815);
nor U13450 (N_13450,N_11523,N_11217);
nor U13451 (N_13451,N_10546,N_11943);
nor U13452 (N_13452,N_11396,N_11596);
xnor U13453 (N_13453,N_10705,N_11470);
xnor U13454 (N_13454,N_11692,N_10750);
or U13455 (N_13455,N_10689,N_11647);
xnor U13456 (N_13456,N_10039,N_11339);
nand U13457 (N_13457,N_11178,N_10083);
nand U13458 (N_13458,N_10127,N_11357);
nor U13459 (N_13459,N_11509,N_11678);
xnor U13460 (N_13460,N_11293,N_11121);
nand U13461 (N_13461,N_10294,N_11672);
nand U13462 (N_13462,N_10674,N_10523);
nor U13463 (N_13463,N_10719,N_10490);
xnor U13464 (N_13464,N_10788,N_11822);
nor U13465 (N_13465,N_10550,N_10560);
nand U13466 (N_13466,N_10475,N_11356);
nand U13467 (N_13467,N_11996,N_11266);
or U13468 (N_13468,N_11596,N_11711);
nor U13469 (N_13469,N_10937,N_10720);
nand U13470 (N_13470,N_10636,N_10505);
nand U13471 (N_13471,N_10187,N_11550);
and U13472 (N_13472,N_11859,N_10944);
nand U13473 (N_13473,N_11699,N_11724);
and U13474 (N_13474,N_10849,N_11190);
nor U13475 (N_13475,N_11252,N_11899);
and U13476 (N_13476,N_10634,N_10763);
or U13477 (N_13477,N_11595,N_11485);
nand U13478 (N_13478,N_11005,N_11657);
nand U13479 (N_13479,N_11660,N_11191);
nand U13480 (N_13480,N_10218,N_11534);
nand U13481 (N_13481,N_11869,N_10396);
or U13482 (N_13482,N_11930,N_10964);
xnor U13483 (N_13483,N_10370,N_11088);
nand U13484 (N_13484,N_11763,N_10328);
and U13485 (N_13485,N_10525,N_10109);
and U13486 (N_13486,N_10965,N_11249);
nand U13487 (N_13487,N_11107,N_11420);
and U13488 (N_13488,N_10612,N_10674);
xnor U13489 (N_13489,N_10709,N_10863);
xnor U13490 (N_13490,N_11717,N_10257);
xnor U13491 (N_13491,N_10232,N_11237);
or U13492 (N_13492,N_10797,N_11083);
and U13493 (N_13493,N_11658,N_11899);
nor U13494 (N_13494,N_11535,N_10035);
xnor U13495 (N_13495,N_10794,N_10028);
or U13496 (N_13496,N_11943,N_10493);
and U13497 (N_13497,N_10646,N_11959);
and U13498 (N_13498,N_11357,N_10507);
and U13499 (N_13499,N_10868,N_11024);
or U13500 (N_13500,N_10755,N_11207);
nand U13501 (N_13501,N_11401,N_11774);
or U13502 (N_13502,N_10928,N_11837);
xnor U13503 (N_13503,N_11290,N_10250);
nor U13504 (N_13504,N_10337,N_10561);
or U13505 (N_13505,N_11340,N_11755);
nor U13506 (N_13506,N_10721,N_10606);
xor U13507 (N_13507,N_10525,N_11600);
or U13508 (N_13508,N_10068,N_11177);
and U13509 (N_13509,N_10229,N_11266);
and U13510 (N_13510,N_11002,N_10602);
nand U13511 (N_13511,N_11499,N_10914);
and U13512 (N_13512,N_11436,N_10374);
or U13513 (N_13513,N_10584,N_11320);
and U13514 (N_13514,N_10846,N_10392);
and U13515 (N_13515,N_11933,N_11226);
nor U13516 (N_13516,N_10185,N_10443);
nand U13517 (N_13517,N_11177,N_10988);
nand U13518 (N_13518,N_10586,N_11237);
or U13519 (N_13519,N_11442,N_10271);
or U13520 (N_13520,N_11802,N_11356);
or U13521 (N_13521,N_11426,N_10649);
and U13522 (N_13522,N_10894,N_10026);
or U13523 (N_13523,N_10144,N_11128);
or U13524 (N_13524,N_10154,N_11826);
nor U13525 (N_13525,N_10095,N_11201);
xnor U13526 (N_13526,N_10043,N_10836);
xnor U13527 (N_13527,N_10706,N_10667);
nand U13528 (N_13528,N_10368,N_10881);
and U13529 (N_13529,N_10940,N_11312);
nor U13530 (N_13530,N_11901,N_10784);
nor U13531 (N_13531,N_10187,N_10990);
or U13532 (N_13532,N_10287,N_10922);
and U13533 (N_13533,N_10582,N_11417);
nor U13534 (N_13534,N_11249,N_10440);
or U13535 (N_13535,N_11314,N_11023);
nand U13536 (N_13536,N_11565,N_10827);
xor U13537 (N_13537,N_10931,N_10928);
nor U13538 (N_13538,N_11131,N_11278);
nand U13539 (N_13539,N_11804,N_11907);
nor U13540 (N_13540,N_10195,N_10474);
xor U13541 (N_13541,N_10465,N_11205);
nand U13542 (N_13542,N_11401,N_10619);
and U13543 (N_13543,N_10269,N_10096);
xnor U13544 (N_13544,N_11988,N_11153);
nor U13545 (N_13545,N_10549,N_10604);
nand U13546 (N_13546,N_10301,N_11986);
and U13547 (N_13547,N_11208,N_11059);
nand U13548 (N_13548,N_10112,N_10015);
nand U13549 (N_13549,N_10770,N_10894);
and U13550 (N_13550,N_11982,N_10338);
nor U13551 (N_13551,N_11307,N_10582);
xor U13552 (N_13552,N_11604,N_11098);
xnor U13553 (N_13553,N_11588,N_10838);
nand U13554 (N_13554,N_11644,N_11766);
nor U13555 (N_13555,N_10438,N_10539);
nor U13556 (N_13556,N_11821,N_11525);
nand U13557 (N_13557,N_10629,N_11284);
nand U13558 (N_13558,N_11002,N_11532);
xor U13559 (N_13559,N_11415,N_10578);
or U13560 (N_13560,N_11963,N_11654);
nor U13561 (N_13561,N_10695,N_11619);
nor U13562 (N_13562,N_10956,N_10024);
nor U13563 (N_13563,N_10139,N_10918);
nor U13564 (N_13564,N_10947,N_11338);
or U13565 (N_13565,N_10374,N_10856);
nor U13566 (N_13566,N_11182,N_10064);
or U13567 (N_13567,N_10241,N_10490);
nand U13568 (N_13568,N_11198,N_10046);
and U13569 (N_13569,N_11370,N_10260);
or U13570 (N_13570,N_11772,N_10768);
xnor U13571 (N_13571,N_11248,N_10844);
or U13572 (N_13572,N_11048,N_11285);
nor U13573 (N_13573,N_11859,N_11313);
or U13574 (N_13574,N_11759,N_11094);
xor U13575 (N_13575,N_10005,N_11489);
and U13576 (N_13576,N_11259,N_10155);
or U13577 (N_13577,N_10800,N_11791);
or U13578 (N_13578,N_10698,N_10496);
or U13579 (N_13579,N_11140,N_10196);
nand U13580 (N_13580,N_11681,N_11756);
and U13581 (N_13581,N_10336,N_10027);
xnor U13582 (N_13582,N_10448,N_11019);
nand U13583 (N_13583,N_10203,N_10026);
or U13584 (N_13584,N_11740,N_11279);
nand U13585 (N_13585,N_11070,N_11629);
xnor U13586 (N_13586,N_10364,N_11589);
or U13587 (N_13587,N_11526,N_11517);
nor U13588 (N_13588,N_10785,N_10254);
and U13589 (N_13589,N_10222,N_11659);
or U13590 (N_13590,N_10220,N_11821);
nor U13591 (N_13591,N_10946,N_10465);
or U13592 (N_13592,N_11475,N_11033);
or U13593 (N_13593,N_10759,N_11856);
and U13594 (N_13594,N_10687,N_10299);
nand U13595 (N_13595,N_10075,N_11334);
nor U13596 (N_13596,N_10631,N_10780);
and U13597 (N_13597,N_10548,N_11013);
xnor U13598 (N_13598,N_11793,N_10728);
nand U13599 (N_13599,N_10855,N_11714);
xor U13600 (N_13600,N_11620,N_10268);
xnor U13601 (N_13601,N_10709,N_10619);
nor U13602 (N_13602,N_10464,N_10255);
and U13603 (N_13603,N_10095,N_10253);
and U13604 (N_13604,N_11375,N_10599);
xnor U13605 (N_13605,N_11521,N_11094);
xor U13606 (N_13606,N_11007,N_10062);
and U13607 (N_13607,N_10104,N_11565);
nand U13608 (N_13608,N_10499,N_10379);
and U13609 (N_13609,N_10688,N_10081);
or U13610 (N_13610,N_11609,N_11363);
and U13611 (N_13611,N_11435,N_11270);
xnor U13612 (N_13612,N_11604,N_10092);
nor U13613 (N_13613,N_10427,N_10717);
nor U13614 (N_13614,N_11673,N_11246);
xnor U13615 (N_13615,N_11055,N_10515);
nor U13616 (N_13616,N_11636,N_10981);
xnor U13617 (N_13617,N_11382,N_11022);
nor U13618 (N_13618,N_11659,N_11040);
nand U13619 (N_13619,N_11505,N_11909);
nor U13620 (N_13620,N_10931,N_10894);
xnor U13621 (N_13621,N_11160,N_10672);
nor U13622 (N_13622,N_11731,N_10593);
xor U13623 (N_13623,N_10918,N_10147);
nand U13624 (N_13624,N_10837,N_10441);
nor U13625 (N_13625,N_11537,N_11622);
xnor U13626 (N_13626,N_10216,N_11182);
and U13627 (N_13627,N_10013,N_11595);
nand U13628 (N_13628,N_10745,N_11731);
xnor U13629 (N_13629,N_11903,N_11829);
xnor U13630 (N_13630,N_11388,N_11530);
and U13631 (N_13631,N_10565,N_11008);
nand U13632 (N_13632,N_10290,N_11646);
xnor U13633 (N_13633,N_10607,N_11336);
nand U13634 (N_13634,N_11135,N_11009);
nor U13635 (N_13635,N_10517,N_11468);
and U13636 (N_13636,N_10837,N_10442);
and U13637 (N_13637,N_11588,N_11199);
xnor U13638 (N_13638,N_11412,N_11960);
nand U13639 (N_13639,N_11740,N_11619);
nand U13640 (N_13640,N_10029,N_11583);
xor U13641 (N_13641,N_10105,N_11853);
nand U13642 (N_13642,N_11164,N_11001);
xor U13643 (N_13643,N_10290,N_11889);
nand U13644 (N_13644,N_11087,N_10046);
and U13645 (N_13645,N_10061,N_11920);
nand U13646 (N_13646,N_11707,N_10783);
xnor U13647 (N_13647,N_11215,N_11238);
nor U13648 (N_13648,N_10949,N_10880);
and U13649 (N_13649,N_10248,N_10904);
and U13650 (N_13650,N_10920,N_11802);
xnor U13651 (N_13651,N_10752,N_10792);
nand U13652 (N_13652,N_11364,N_11868);
xor U13653 (N_13653,N_10399,N_11923);
xor U13654 (N_13654,N_11375,N_11050);
and U13655 (N_13655,N_11586,N_11817);
and U13656 (N_13656,N_10536,N_10185);
xor U13657 (N_13657,N_10861,N_10484);
xor U13658 (N_13658,N_11647,N_10655);
xnor U13659 (N_13659,N_11716,N_10634);
nor U13660 (N_13660,N_10106,N_10513);
nand U13661 (N_13661,N_10953,N_11763);
nor U13662 (N_13662,N_10981,N_11302);
nor U13663 (N_13663,N_10699,N_10009);
nor U13664 (N_13664,N_11512,N_11330);
xor U13665 (N_13665,N_11801,N_11051);
nand U13666 (N_13666,N_10109,N_11150);
nand U13667 (N_13667,N_10442,N_11733);
xor U13668 (N_13668,N_10988,N_10091);
or U13669 (N_13669,N_10303,N_10126);
or U13670 (N_13670,N_11704,N_11352);
and U13671 (N_13671,N_10500,N_11994);
nor U13672 (N_13672,N_10534,N_10767);
and U13673 (N_13673,N_11717,N_10733);
xor U13674 (N_13674,N_10557,N_11976);
or U13675 (N_13675,N_10067,N_11519);
or U13676 (N_13676,N_11474,N_10901);
nor U13677 (N_13677,N_11962,N_10595);
and U13678 (N_13678,N_11911,N_10989);
or U13679 (N_13679,N_11956,N_11966);
nand U13680 (N_13680,N_11474,N_11163);
or U13681 (N_13681,N_11020,N_10112);
nor U13682 (N_13682,N_11281,N_11942);
nor U13683 (N_13683,N_10296,N_10655);
or U13684 (N_13684,N_11209,N_11230);
or U13685 (N_13685,N_11070,N_11014);
or U13686 (N_13686,N_11528,N_11482);
or U13687 (N_13687,N_10771,N_10065);
or U13688 (N_13688,N_10789,N_10059);
nand U13689 (N_13689,N_10686,N_11965);
nand U13690 (N_13690,N_11640,N_11703);
nor U13691 (N_13691,N_10386,N_11132);
and U13692 (N_13692,N_10300,N_10657);
and U13693 (N_13693,N_11564,N_10206);
nor U13694 (N_13694,N_10411,N_11433);
nand U13695 (N_13695,N_11734,N_10391);
nand U13696 (N_13696,N_10261,N_11169);
nor U13697 (N_13697,N_11837,N_11583);
or U13698 (N_13698,N_11246,N_10194);
or U13699 (N_13699,N_11540,N_10071);
nand U13700 (N_13700,N_10349,N_11509);
and U13701 (N_13701,N_11006,N_10308);
nand U13702 (N_13702,N_11409,N_10236);
and U13703 (N_13703,N_11622,N_11030);
and U13704 (N_13704,N_11731,N_10340);
nand U13705 (N_13705,N_10008,N_10299);
xor U13706 (N_13706,N_11109,N_10388);
xnor U13707 (N_13707,N_10443,N_10423);
xnor U13708 (N_13708,N_10657,N_10599);
nand U13709 (N_13709,N_11945,N_11389);
xor U13710 (N_13710,N_11569,N_10310);
and U13711 (N_13711,N_10445,N_11194);
xnor U13712 (N_13712,N_10951,N_10709);
or U13713 (N_13713,N_11064,N_10817);
nand U13714 (N_13714,N_10841,N_11536);
nor U13715 (N_13715,N_10599,N_10936);
nor U13716 (N_13716,N_10075,N_11012);
nand U13717 (N_13717,N_10321,N_11898);
xnor U13718 (N_13718,N_11173,N_11982);
xor U13719 (N_13719,N_10574,N_10320);
or U13720 (N_13720,N_11905,N_11309);
xor U13721 (N_13721,N_10625,N_10028);
and U13722 (N_13722,N_11051,N_10042);
xor U13723 (N_13723,N_11197,N_11934);
and U13724 (N_13724,N_11417,N_11380);
nand U13725 (N_13725,N_11609,N_10471);
or U13726 (N_13726,N_10845,N_11996);
xor U13727 (N_13727,N_10521,N_11523);
nand U13728 (N_13728,N_10309,N_10190);
nand U13729 (N_13729,N_10230,N_11255);
nand U13730 (N_13730,N_11498,N_11684);
xor U13731 (N_13731,N_10221,N_11907);
nand U13732 (N_13732,N_10469,N_11258);
and U13733 (N_13733,N_10120,N_11783);
and U13734 (N_13734,N_10076,N_10560);
nand U13735 (N_13735,N_10229,N_11262);
or U13736 (N_13736,N_10073,N_11578);
xor U13737 (N_13737,N_10633,N_11282);
or U13738 (N_13738,N_11352,N_10254);
nor U13739 (N_13739,N_11378,N_11153);
or U13740 (N_13740,N_10970,N_10551);
nand U13741 (N_13741,N_10823,N_11042);
and U13742 (N_13742,N_11699,N_11162);
nor U13743 (N_13743,N_10213,N_11826);
and U13744 (N_13744,N_11135,N_11971);
nor U13745 (N_13745,N_10953,N_11867);
nor U13746 (N_13746,N_11541,N_11009);
or U13747 (N_13747,N_10926,N_11154);
or U13748 (N_13748,N_10431,N_10674);
nor U13749 (N_13749,N_11533,N_11108);
nor U13750 (N_13750,N_10240,N_11861);
nand U13751 (N_13751,N_11995,N_11635);
or U13752 (N_13752,N_10994,N_10160);
and U13753 (N_13753,N_10165,N_10259);
nand U13754 (N_13754,N_11918,N_11258);
nand U13755 (N_13755,N_10361,N_11094);
or U13756 (N_13756,N_10571,N_10193);
nor U13757 (N_13757,N_11227,N_11919);
nor U13758 (N_13758,N_10502,N_10380);
or U13759 (N_13759,N_11821,N_10931);
nor U13760 (N_13760,N_11448,N_10443);
nor U13761 (N_13761,N_11102,N_11761);
nor U13762 (N_13762,N_11142,N_11778);
nand U13763 (N_13763,N_10377,N_10203);
or U13764 (N_13764,N_11631,N_10828);
and U13765 (N_13765,N_11356,N_11695);
nand U13766 (N_13766,N_11861,N_10881);
and U13767 (N_13767,N_10001,N_10299);
and U13768 (N_13768,N_10442,N_11735);
and U13769 (N_13769,N_11987,N_10598);
or U13770 (N_13770,N_11635,N_11686);
or U13771 (N_13771,N_10453,N_11756);
or U13772 (N_13772,N_11106,N_10004);
xor U13773 (N_13773,N_11664,N_10784);
nor U13774 (N_13774,N_10361,N_11621);
and U13775 (N_13775,N_10156,N_10713);
xor U13776 (N_13776,N_10504,N_11934);
nand U13777 (N_13777,N_11865,N_10222);
nor U13778 (N_13778,N_10797,N_10059);
or U13779 (N_13779,N_11254,N_11573);
or U13780 (N_13780,N_10045,N_11515);
and U13781 (N_13781,N_11709,N_11344);
or U13782 (N_13782,N_10354,N_10284);
nand U13783 (N_13783,N_11933,N_10842);
nand U13784 (N_13784,N_10408,N_10768);
xor U13785 (N_13785,N_10424,N_10714);
nand U13786 (N_13786,N_10451,N_11067);
nand U13787 (N_13787,N_10414,N_11808);
and U13788 (N_13788,N_10785,N_10922);
and U13789 (N_13789,N_11870,N_10831);
or U13790 (N_13790,N_10308,N_11798);
or U13791 (N_13791,N_10289,N_11572);
nand U13792 (N_13792,N_11194,N_11450);
and U13793 (N_13793,N_10752,N_10948);
nand U13794 (N_13794,N_10640,N_11864);
nor U13795 (N_13795,N_11921,N_11464);
xnor U13796 (N_13796,N_10326,N_10256);
xnor U13797 (N_13797,N_10042,N_11864);
nand U13798 (N_13798,N_11056,N_10830);
nand U13799 (N_13799,N_11867,N_10467);
nor U13800 (N_13800,N_11276,N_10141);
nor U13801 (N_13801,N_10279,N_11867);
nand U13802 (N_13802,N_11951,N_10069);
and U13803 (N_13803,N_10348,N_10248);
and U13804 (N_13804,N_11252,N_10485);
xnor U13805 (N_13805,N_11565,N_11582);
or U13806 (N_13806,N_11384,N_10453);
or U13807 (N_13807,N_10089,N_10696);
nand U13808 (N_13808,N_11714,N_11582);
nor U13809 (N_13809,N_10191,N_11605);
xor U13810 (N_13810,N_10739,N_10232);
nor U13811 (N_13811,N_10084,N_10919);
and U13812 (N_13812,N_11782,N_10437);
xnor U13813 (N_13813,N_10494,N_11878);
or U13814 (N_13814,N_10610,N_11148);
and U13815 (N_13815,N_10365,N_11035);
xnor U13816 (N_13816,N_11431,N_11420);
nand U13817 (N_13817,N_11676,N_10962);
and U13818 (N_13818,N_10417,N_11903);
nand U13819 (N_13819,N_11806,N_11339);
nor U13820 (N_13820,N_11372,N_11486);
or U13821 (N_13821,N_10432,N_10482);
nor U13822 (N_13822,N_10236,N_11349);
xor U13823 (N_13823,N_11691,N_11548);
nor U13824 (N_13824,N_10455,N_11183);
nand U13825 (N_13825,N_10435,N_10397);
nand U13826 (N_13826,N_11814,N_11459);
nor U13827 (N_13827,N_10533,N_10405);
nand U13828 (N_13828,N_11058,N_10838);
or U13829 (N_13829,N_10201,N_10739);
or U13830 (N_13830,N_10481,N_10275);
or U13831 (N_13831,N_10906,N_11283);
nor U13832 (N_13832,N_10011,N_10740);
or U13833 (N_13833,N_10788,N_10454);
or U13834 (N_13834,N_10073,N_11674);
xnor U13835 (N_13835,N_11377,N_10812);
and U13836 (N_13836,N_10631,N_10184);
nand U13837 (N_13837,N_11495,N_10056);
nand U13838 (N_13838,N_11624,N_11400);
nor U13839 (N_13839,N_10157,N_11090);
nor U13840 (N_13840,N_11017,N_10014);
xor U13841 (N_13841,N_11956,N_11060);
and U13842 (N_13842,N_11342,N_11303);
nand U13843 (N_13843,N_11129,N_10597);
xnor U13844 (N_13844,N_11712,N_10600);
and U13845 (N_13845,N_10050,N_11334);
nor U13846 (N_13846,N_11088,N_10808);
xnor U13847 (N_13847,N_11717,N_11280);
nor U13848 (N_13848,N_11459,N_10388);
nand U13849 (N_13849,N_10591,N_10021);
xor U13850 (N_13850,N_10616,N_10439);
nor U13851 (N_13851,N_11803,N_11810);
and U13852 (N_13852,N_10516,N_10055);
nor U13853 (N_13853,N_10797,N_10267);
and U13854 (N_13854,N_11898,N_11784);
nand U13855 (N_13855,N_10422,N_10477);
xor U13856 (N_13856,N_11152,N_11879);
or U13857 (N_13857,N_10912,N_10192);
and U13858 (N_13858,N_11602,N_10627);
nor U13859 (N_13859,N_10195,N_11742);
or U13860 (N_13860,N_10535,N_10448);
xnor U13861 (N_13861,N_11186,N_10154);
xor U13862 (N_13862,N_10471,N_11085);
and U13863 (N_13863,N_10183,N_10705);
nand U13864 (N_13864,N_11283,N_10418);
nor U13865 (N_13865,N_10306,N_11472);
or U13866 (N_13866,N_10053,N_11950);
xnor U13867 (N_13867,N_10165,N_10577);
nand U13868 (N_13868,N_11162,N_10230);
nand U13869 (N_13869,N_11501,N_11550);
xor U13870 (N_13870,N_10470,N_11761);
nand U13871 (N_13871,N_11737,N_11187);
nand U13872 (N_13872,N_11695,N_11362);
nand U13873 (N_13873,N_10954,N_11277);
xnor U13874 (N_13874,N_10993,N_10427);
nor U13875 (N_13875,N_11413,N_10808);
and U13876 (N_13876,N_11616,N_10492);
and U13877 (N_13877,N_10660,N_11949);
nor U13878 (N_13878,N_10796,N_10151);
and U13879 (N_13879,N_10648,N_11176);
nor U13880 (N_13880,N_10484,N_11420);
and U13881 (N_13881,N_10303,N_10478);
or U13882 (N_13882,N_10716,N_10973);
nor U13883 (N_13883,N_10185,N_10133);
and U13884 (N_13884,N_11573,N_10295);
xnor U13885 (N_13885,N_10598,N_11833);
nand U13886 (N_13886,N_10297,N_10713);
and U13887 (N_13887,N_10469,N_10174);
nand U13888 (N_13888,N_11225,N_11329);
xor U13889 (N_13889,N_10464,N_10512);
nand U13890 (N_13890,N_10040,N_10602);
or U13891 (N_13891,N_11949,N_10028);
or U13892 (N_13892,N_11875,N_11959);
or U13893 (N_13893,N_11963,N_11081);
or U13894 (N_13894,N_11568,N_10740);
nor U13895 (N_13895,N_11191,N_10307);
nand U13896 (N_13896,N_10861,N_10289);
nor U13897 (N_13897,N_10123,N_11911);
nor U13898 (N_13898,N_10812,N_10386);
or U13899 (N_13899,N_10030,N_10386);
nor U13900 (N_13900,N_11074,N_10331);
nand U13901 (N_13901,N_11281,N_11334);
and U13902 (N_13902,N_10459,N_10085);
nand U13903 (N_13903,N_10802,N_10930);
or U13904 (N_13904,N_10703,N_10909);
nand U13905 (N_13905,N_11052,N_10878);
or U13906 (N_13906,N_10182,N_11132);
nand U13907 (N_13907,N_10315,N_11841);
nand U13908 (N_13908,N_11904,N_10237);
xnor U13909 (N_13909,N_10249,N_10710);
nor U13910 (N_13910,N_10662,N_11745);
xnor U13911 (N_13911,N_10045,N_11297);
nand U13912 (N_13912,N_10734,N_11467);
nor U13913 (N_13913,N_11125,N_11045);
or U13914 (N_13914,N_10072,N_11396);
nor U13915 (N_13915,N_11419,N_11560);
nand U13916 (N_13916,N_11905,N_10672);
or U13917 (N_13917,N_10728,N_10344);
nor U13918 (N_13918,N_11408,N_11414);
xnor U13919 (N_13919,N_11217,N_11629);
xnor U13920 (N_13920,N_10801,N_10645);
xor U13921 (N_13921,N_11745,N_11969);
nand U13922 (N_13922,N_11949,N_11740);
nor U13923 (N_13923,N_11105,N_11652);
nor U13924 (N_13924,N_11545,N_11872);
and U13925 (N_13925,N_11023,N_11252);
nand U13926 (N_13926,N_11963,N_11819);
nand U13927 (N_13927,N_10128,N_10340);
nand U13928 (N_13928,N_11092,N_11268);
nor U13929 (N_13929,N_10602,N_11588);
or U13930 (N_13930,N_11261,N_10211);
and U13931 (N_13931,N_11449,N_11555);
nor U13932 (N_13932,N_11571,N_10814);
nand U13933 (N_13933,N_11305,N_11102);
or U13934 (N_13934,N_10560,N_10379);
and U13935 (N_13935,N_11267,N_10972);
nand U13936 (N_13936,N_10021,N_11951);
nor U13937 (N_13937,N_11931,N_10424);
or U13938 (N_13938,N_11740,N_11976);
nor U13939 (N_13939,N_10343,N_11663);
xor U13940 (N_13940,N_11956,N_10929);
nand U13941 (N_13941,N_11855,N_10775);
and U13942 (N_13942,N_11544,N_11465);
or U13943 (N_13943,N_10836,N_11701);
nand U13944 (N_13944,N_10216,N_10495);
and U13945 (N_13945,N_11371,N_10541);
or U13946 (N_13946,N_11448,N_10059);
and U13947 (N_13947,N_10772,N_10505);
and U13948 (N_13948,N_11298,N_10628);
nor U13949 (N_13949,N_11982,N_11998);
and U13950 (N_13950,N_11564,N_10243);
and U13951 (N_13951,N_11048,N_10419);
nand U13952 (N_13952,N_10020,N_11001);
or U13953 (N_13953,N_10383,N_10910);
xnor U13954 (N_13954,N_10990,N_10863);
nand U13955 (N_13955,N_11521,N_10579);
nor U13956 (N_13956,N_10061,N_10070);
xnor U13957 (N_13957,N_11511,N_10907);
nor U13958 (N_13958,N_11260,N_11641);
nor U13959 (N_13959,N_10848,N_11969);
xor U13960 (N_13960,N_11207,N_11892);
nand U13961 (N_13961,N_10726,N_10648);
nand U13962 (N_13962,N_10021,N_10079);
nor U13963 (N_13963,N_11823,N_10066);
or U13964 (N_13964,N_10899,N_10356);
nor U13965 (N_13965,N_11107,N_11859);
or U13966 (N_13966,N_11416,N_11428);
or U13967 (N_13967,N_10536,N_10701);
nand U13968 (N_13968,N_10056,N_10208);
xnor U13969 (N_13969,N_11733,N_11002);
or U13970 (N_13970,N_10844,N_10652);
and U13971 (N_13971,N_10136,N_10768);
xnor U13972 (N_13972,N_11399,N_10006);
xor U13973 (N_13973,N_10164,N_10889);
nor U13974 (N_13974,N_11830,N_10800);
nor U13975 (N_13975,N_11962,N_10065);
or U13976 (N_13976,N_10591,N_10113);
nand U13977 (N_13977,N_11723,N_11461);
nand U13978 (N_13978,N_11581,N_11005);
or U13979 (N_13979,N_11941,N_11795);
nand U13980 (N_13980,N_11549,N_11760);
nor U13981 (N_13981,N_11052,N_10367);
xnor U13982 (N_13982,N_11597,N_11093);
xor U13983 (N_13983,N_10431,N_11407);
nand U13984 (N_13984,N_11362,N_10614);
and U13985 (N_13985,N_11224,N_10961);
nand U13986 (N_13986,N_10710,N_10697);
nor U13987 (N_13987,N_11080,N_11877);
xnor U13988 (N_13988,N_11111,N_11917);
nand U13989 (N_13989,N_11765,N_10580);
xor U13990 (N_13990,N_10308,N_11731);
nand U13991 (N_13991,N_11023,N_10504);
nor U13992 (N_13992,N_11340,N_10170);
xnor U13993 (N_13993,N_10804,N_11918);
and U13994 (N_13994,N_11965,N_11346);
xor U13995 (N_13995,N_11248,N_10330);
nor U13996 (N_13996,N_11896,N_11488);
nor U13997 (N_13997,N_11187,N_11122);
and U13998 (N_13998,N_10958,N_11068);
xor U13999 (N_13999,N_11663,N_10051);
xor U14000 (N_14000,N_13759,N_13041);
nand U14001 (N_14001,N_12547,N_12363);
nor U14002 (N_14002,N_12713,N_13931);
nor U14003 (N_14003,N_13833,N_13127);
nand U14004 (N_14004,N_12633,N_12059);
or U14005 (N_14005,N_12744,N_12045);
nand U14006 (N_14006,N_13923,N_13550);
xnor U14007 (N_14007,N_12806,N_13251);
nor U14008 (N_14008,N_12188,N_13319);
nand U14009 (N_14009,N_13510,N_12338);
and U14010 (N_14010,N_12126,N_13365);
nand U14011 (N_14011,N_12628,N_12864);
nand U14012 (N_14012,N_12025,N_12056);
and U14013 (N_14013,N_12588,N_13695);
nand U14014 (N_14014,N_13117,N_13873);
xnor U14015 (N_14015,N_12106,N_12478);
nand U14016 (N_14016,N_13414,N_13920);
xor U14017 (N_14017,N_13123,N_13140);
nor U14018 (N_14018,N_13783,N_12417);
and U14019 (N_14019,N_12399,N_12233);
nand U14020 (N_14020,N_13522,N_13216);
xnor U14021 (N_14021,N_13625,N_12248);
nand U14022 (N_14022,N_12447,N_12603);
or U14023 (N_14023,N_13806,N_13858);
and U14024 (N_14024,N_12510,N_12245);
xor U14025 (N_14025,N_13582,N_13932);
nor U14026 (N_14026,N_13190,N_13683);
or U14027 (N_14027,N_12961,N_12630);
nor U14028 (N_14028,N_13684,N_12142);
nand U14029 (N_14029,N_13405,N_12115);
nor U14030 (N_14030,N_13372,N_13142);
nand U14031 (N_14031,N_13407,N_12214);
nand U14032 (N_14032,N_12232,N_13347);
xnor U14033 (N_14033,N_13993,N_12169);
nand U14034 (N_14034,N_12272,N_12033);
or U14035 (N_14035,N_13616,N_12261);
xnor U14036 (N_14036,N_13348,N_13781);
and U14037 (N_14037,N_12640,N_13902);
nor U14038 (N_14038,N_13072,N_13831);
nor U14039 (N_14039,N_12354,N_13176);
and U14040 (N_14040,N_12515,N_13740);
xnor U14041 (N_14041,N_12830,N_12611);
nand U14042 (N_14042,N_12449,N_12181);
xnor U14043 (N_14043,N_12645,N_12779);
and U14044 (N_14044,N_12790,N_13069);
nor U14045 (N_14045,N_12884,N_13020);
and U14046 (N_14046,N_13776,N_12010);
nor U14047 (N_14047,N_13571,N_13496);
or U14048 (N_14048,N_12189,N_12937);
nor U14049 (N_14049,N_12255,N_12632);
nor U14050 (N_14050,N_12287,N_12361);
xor U14051 (N_14051,N_12737,N_13549);
nor U14052 (N_14052,N_12296,N_13475);
xnor U14053 (N_14053,N_12845,N_13434);
xnor U14054 (N_14054,N_12027,N_13480);
and U14055 (N_14055,N_13904,N_12266);
or U14056 (N_14056,N_13188,N_12557);
xnor U14057 (N_14057,N_12583,N_12860);
xnor U14058 (N_14058,N_12306,N_12295);
nand U14059 (N_14059,N_12317,N_13247);
and U14060 (N_14060,N_12765,N_12899);
xor U14061 (N_14061,N_12065,N_13563);
xor U14062 (N_14062,N_12176,N_13681);
and U14063 (N_14063,N_12007,N_12999);
nor U14064 (N_14064,N_13599,N_12279);
nor U14065 (N_14065,N_13311,N_12568);
and U14066 (N_14066,N_13736,N_13044);
and U14067 (N_14067,N_12532,N_13560);
nor U14068 (N_14068,N_13918,N_13099);
or U14069 (N_14069,N_12320,N_12822);
nor U14070 (N_14070,N_12225,N_12163);
nand U14071 (N_14071,N_13864,N_12170);
xnor U14072 (N_14072,N_12664,N_12504);
or U14073 (N_14073,N_12271,N_12308);
nand U14074 (N_14074,N_12331,N_12876);
nand U14075 (N_14075,N_13997,N_13274);
nand U14076 (N_14076,N_13441,N_12259);
xnor U14077 (N_14077,N_12959,N_13402);
or U14078 (N_14078,N_13789,N_12647);
nand U14079 (N_14079,N_12008,N_13258);
nor U14080 (N_14080,N_13682,N_12000);
nand U14081 (N_14081,N_13323,N_13288);
nand U14082 (N_14082,N_12618,N_13087);
and U14083 (N_14083,N_12955,N_12373);
and U14084 (N_14084,N_13276,N_13284);
or U14085 (N_14085,N_12337,N_13824);
nand U14086 (N_14086,N_12843,N_13185);
and U14087 (N_14087,N_12511,N_13801);
and U14088 (N_14088,N_12817,N_13792);
xor U14089 (N_14089,N_12850,N_13903);
and U14090 (N_14090,N_13883,N_13114);
nand U14091 (N_14091,N_13063,N_13081);
or U14092 (N_14092,N_13653,N_13652);
and U14093 (N_14093,N_12122,N_12656);
and U14094 (N_14094,N_12253,N_13690);
xor U14095 (N_14095,N_12997,N_13233);
nor U14096 (N_14096,N_12362,N_13723);
and U14097 (N_14097,N_13969,N_13587);
and U14098 (N_14098,N_12401,N_13760);
nor U14099 (N_14099,N_12523,N_13772);
xor U14100 (N_14100,N_12680,N_13203);
or U14101 (N_14101,N_13881,N_13906);
nor U14102 (N_14102,N_12151,N_13228);
nand U14103 (N_14103,N_12996,N_12521);
and U14104 (N_14104,N_12671,N_13335);
and U14105 (N_14105,N_13548,N_12453);
nor U14106 (N_14106,N_12629,N_12587);
xnor U14107 (N_14107,N_13602,N_12727);
xnor U14108 (N_14108,N_12646,N_13054);
xor U14109 (N_14109,N_13011,N_12638);
or U14110 (N_14110,N_12152,N_12082);
xnor U14111 (N_14111,N_12741,N_12528);
nand U14112 (N_14112,N_12116,N_12692);
and U14113 (N_14113,N_13463,N_13147);
nor U14114 (N_14114,N_12856,N_13905);
nand U14115 (N_14115,N_12683,N_12834);
or U14116 (N_14116,N_12653,N_13568);
nor U14117 (N_14117,N_13397,N_12085);
nand U14118 (N_14118,N_13609,N_12762);
and U14119 (N_14119,N_13161,N_13950);
nor U14120 (N_14120,N_12626,N_12662);
xor U14121 (N_14121,N_12435,N_13915);
and U14122 (N_14122,N_12672,N_13248);
and U14123 (N_14123,N_13083,N_12734);
nor U14124 (N_14124,N_12851,N_13492);
and U14125 (N_14125,N_12702,N_12930);
nand U14126 (N_14126,N_13930,N_13473);
nor U14127 (N_14127,N_12965,N_13565);
and U14128 (N_14128,N_12358,N_12198);
xnor U14129 (N_14129,N_13564,N_13380);
nor U14130 (N_14130,N_13738,N_13673);
xnor U14131 (N_14131,N_12828,N_13882);
xor U14132 (N_14132,N_13674,N_12813);
or U14133 (N_14133,N_12303,N_12659);
and U14134 (N_14134,N_13192,N_12885);
and U14135 (N_14135,N_12440,N_12346);
nand U14136 (N_14136,N_12015,N_12263);
and U14137 (N_14137,N_12313,N_13495);
nor U14138 (N_14138,N_12668,N_13164);
nor U14139 (N_14139,N_12284,N_12250);
nor U14140 (N_14140,N_12601,N_13057);
or U14141 (N_14141,N_12578,N_13913);
nor U14142 (N_14142,N_13502,N_13922);
nand U14143 (N_14143,N_12658,N_13221);
and U14144 (N_14144,N_12751,N_13384);
nor U14145 (N_14145,N_12458,N_12757);
nand U14146 (N_14146,N_13927,N_13045);
nor U14147 (N_14147,N_13659,N_12254);
nor U14148 (N_14148,N_13014,N_13416);
nand U14149 (N_14149,N_12770,N_13229);
nor U14150 (N_14150,N_13635,N_13369);
nand U14151 (N_14151,N_13572,N_12068);
xor U14152 (N_14152,N_13462,N_13240);
nand U14153 (N_14153,N_13805,N_13758);
nor U14154 (N_14154,N_13977,N_12782);
or U14155 (N_14155,N_12058,N_12912);
nand U14156 (N_14156,N_13937,N_12404);
nor U14157 (N_14157,N_12565,N_12446);
and U14158 (N_14158,N_12372,N_12720);
xnor U14159 (N_14159,N_13437,N_12969);
xor U14160 (N_14160,N_12552,N_13254);
or U14161 (N_14161,N_13614,N_13677);
xor U14162 (N_14162,N_12732,N_13692);
xnor U14163 (N_14163,N_13711,N_13082);
nand U14164 (N_14164,N_12904,N_12767);
nand U14165 (N_14165,N_13191,N_13113);
nor U14166 (N_14166,N_13489,N_12690);
nor U14167 (N_14167,N_13068,N_12215);
nor U14168 (N_14168,N_13012,N_13158);
nor U14169 (N_14169,N_12073,N_12740);
nand U14170 (N_14170,N_13699,N_13660);
and U14171 (N_14171,N_12479,N_12108);
and U14172 (N_14172,N_12242,N_12725);
xor U14173 (N_14173,N_13004,N_12132);
or U14174 (N_14174,N_13753,N_13184);
xor U14175 (N_14175,N_12766,N_13137);
xnor U14176 (N_14176,N_12219,N_12156);
or U14177 (N_14177,N_12950,N_12335);
nand U14178 (N_14178,N_12875,N_12429);
or U14179 (N_14179,N_13961,N_13090);
nand U14180 (N_14180,N_13938,N_12839);
xor U14181 (N_14181,N_13654,N_12759);
and U14182 (N_14182,N_13048,N_12061);
nand U14183 (N_14183,N_12794,N_13398);
or U14184 (N_14184,N_13089,N_12009);
nand U14185 (N_14185,N_13351,N_12477);
xor U14186 (N_14186,N_13062,N_13947);
nor U14187 (N_14187,N_13367,N_12004);
nand U14188 (N_14188,N_12499,N_12125);
or U14189 (N_14189,N_13763,N_13962);
and U14190 (N_14190,N_12480,N_13601);
xnor U14191 (N_14191,N_13157,N_12311);
nor U14192 (N_14192,N_12957,N_12129);
xor U14193 (N_14193,N_12676,N_12482);
or U14194 (N_14194,N_12408,N_13138);
xnor U14195 (N_14195,N_12451,N_12795);
nand U14196 (N_14196,N_13166,N_13130);
and U14197 (N_14197,N_12369,N_13102);
nor U14198 (N_14198,N_13995,N_13576);
or U14199 (N_14199,N_13303,N_13454);
nand U14200 (N_14200,N_13154,N_13386);
or U14201 (N_14201,N_12634,N_12493);
nand U14202 (N_14202,N_12030,N_13640);
nor U14203 (N_14203,N_12003,N_12269);
xnor U14204 (N_14204,N_13717,N_13604);
nor U14205 (N_14205,N_13476,N_13612);
nand U14206 (N_14206,N_13889,N_13579);
and U14207 (N_14207,N_12090,N_13617);
nor U14208 (N_14208,N_12422,N_13837);
nand U14209 (N_14209,N_13131,N_12467);
or U14210 (N_14210,N_13958,N_13648);
xnor U14211 (N_14211,N_13461,N_13382);
or U14212 (N_14212,N_12079,N_13636);
or U14213 (N_14213,N_13427,N_12827);
nand U14214 (N_14214,N_13340,N_13773);
or U14215 (N_14215,N_12416,N_13867);
xor U14216 (N_14216,N_12909,N_13511);
nor U14217 (N_14217,N_13497,N_13213);
nor U14218 (N_14218,N_12643,N_12426);
or U14219 (N_14219,N_12536,N_12507);
or U14220 (N_14220,N_13500,N_12371);
or U14221 (N_14221,N_13201,N_12432);
nor U14222 (N_14222,N_12925,N_13622);
nor U14223 (N_14223,N_13728,N_12799);
nand U14224 (N_14224,N_13107,N_12312);
nor U14225 (N_14225,N_12699,N_12991);
and U14226 (N_14226,N_12877,N_12614);
xnor U14227 (N_14227,N_12973,N_12454);
nand U14228 (N_14228,N_12879,N_12836);
and U14229 (N_14229,N_12863,N_13182);
or U14230 (N_14230,N_13606,N_12605);
nor U14231 (N_14231,N_13940,N_13104);
or U14232 (N_14232,N_12677,N_12878);
and U14233 (N_14233,N_12141,N_12021);
or U14234 (N_14234,N_12694,N_13133);
or U14235 (N_14235,N_12841,N_13531);
xor U14236 (N_14236,N_13160,N_13440);
nor U14237 (N_14237,N_13028,N_13136);
nor U14238 (N_14238,N_13097,N_13862);
nor U14239 (N_14239,N_12336,N_13042);
nor U14240 (N_14240,N_13632,N_13916);
nand U14241 (N_14241,N_13212,N_13639);
nand U14242 (N_14242,N_12902,N_13729);
xor U14243 (N_14243,N_13523,N_13588);
or U14244 (N_14244,N_13125,N_12423);
nor U14245 (N_14245,N_13146,N_12724);
or U14246 (N_14246,N_13697,N_12260);
nand U14247 (N_14247,N_13735,N_12204);
nor U14248 (N_14248,N_13139,N_12410);
or U14249 (N_14249,N_12052,N_12310);
or U14250 (N_14250,N_12239,N_13408);
or U14251 (N_14251,N_13598,N_13071);
nor U14252 (N_14252,N_13009,N_13153);
nor U14253 (N_14253,N_12971,N_13261);
or U14254 (N_14254,N_12500,N_13413);
xor U14255 (N_14255,N_13945,N_12347);
nor U14256 (N_14256,N_13869,N_12915);
or U14257 (N_14257,N_12746,N_13269);
or U14258 (N_14258,N_13657,N_13939);
xor U14259 (N_14259,N_13442,N_13557);
or U14260 (N_14260,N_12203,N_13234);
xnor U14261 (N_14261,N_13016,N_13286);
nor U14262 (N_14262,N_13946,N_12342);
and U14263 (N_14263,N_13064,N_13030);
and U14264 (N_14264,N_12134,N_13845);
nor U14265 (N_14265,N_12436,N_12264);
or U14266 (N_14266,N_12905,N_13996);
and U14267 (N_14267,N_13836,N_12979);
and U14268 (N_14268,N_13393,N_12881);
or U14269 (N_14269,N_13394,N_13467);
nor U14270 (N_14270,N_12911,N_13449);
nand U14271 (N_14271,N_12838,N_13156);
and U14272 (N_14272,N_13051,N_13821);
nand U14273 (N_14273,N_12993,N_13508);
and U14274 (N_14274,N_12055,N_12434);
and U14275 (N_14275,N_12162,N_13168);
nand U14276 (N_14276,N_13332,N_13799);
nor U14277 (N_14277,N_12534,N_13235);
nor U14278 (N_14278,N_12600,N_12944);
and U14279 (N_14279,N_12484,N_13299);
nor U14280 (N_14280,N_12538,N_12926);
nor U14281 (N_14281,N_13651,N_13554);
or U14282 (N_14282,N_13032,N_12774);
nand U14283 (N_14283,N_13593,N_13756);
or U14284 (N_14284,N_12460,N_12622);
nand U14285 (N_14285,N_12921,N_12120);
or U14286 (N_14286,N_13387,N_13448);
xnor U14287 (N_14287,N_12764,N_13730);
nor U14288 (N_14288,N_12798,N_12067);
xnor U14289 (N_14289,N_12406,N_13360);
or U14290 (N_14290,N_13830,N_12199);
xor U14291 (N_14291,N_13315,N_13509);
nor U14292 (N_14292,N_13895,N_13985);
xor U14293 (N_14293,N_13871,N_12174);
and U14294 (N_14294,N_13003,N_13844);
or U14295 (N_14295,N_13892,N_13943);
xnor U14296 (N_14296,N_12470,N_13267);
and U14297 (N_14297,N_12707,N_12462);
or U14298 (N_14298,N_12339,N_13917);
or U14299 (N_14299,N_12608,N_13007);
nor U14300 (N_14300,N_13793,N_13159);
xnor U14301 (N_14301,N_13976,N_12596);
or U14302 (N_14302,N_13739,N_13953);
xnor U14303 (N_14303,N_13490,N_13465);
and U14304 (N_14304,N_13116,N_13768);
or U14305 (N_14305,N_13936,N_13630);
xnor U14306 (N_14306,N_13691,N_12772);
or U14307 (N_14307,N_12636,N_13714);
xor U14308 (N_14308,N_12220,N_12550);
xnor U14309 (N_14309,N_13325,N_12620);
xor U14310 (N_14310,N_13378,N_12270);
and U14311 (N_14311,N_13577,N_12655);
nand U14312 (N_14312,N_13525,N_13110);
nand U14313 (N_14313,N_13098,N_13443);
or U14314 (N_14314,N_13008,N_12154);
xnor U14315 (N_14315,N_12329,N_12598);
or U14316 (N_14316,N_12666,N_12402);
nor U14317 (N_14317,N_12854,N_13412);
nor U14318 (N_14318,N_12407,N_13470);
nand U14319 (N_14319,N_13298,N_12688);
nand U14320 (N_14320,N_12695,N_12962);
nand U14321 (N_14321,N_12252,N_13876);
nand U14322 (N_14322,N_13210,N_13177);
nand U14323 (N_14323,N_12869,N_12276);
nor U14324 (N_14324,N_12942,N_13162);
and U14325 (N_14325,N_13446,N_12022);
and U14326 (N_14326,N_13912,N_12865);
nor U14327 (N_14327,N_13151,N_12922);
xor U14328 (N_14328,N_12047,N_13350);
nor U14329 (N_14329,N_12903,N_13537);
and U14330 (N_14330,N_13921,N_13388);
and U14331 (N_14331,N_13747,N_13106);
nand U14332 (N_14332,N_13933,N_13574);
or U14333 (N_14333,N_13941,N_13732);
or U14334 (N_14334,N_12370,N_13757);
and U14335 (N_14335,N_13866,N_13929);
or U14336 (N_14336,N_12989,N_13310);
xor U14337 (N_14337,N_12826,N_12686);
nor U14338 (N_14338,N_12414,N_12716);
xnor U14339 (N_14339,N_13779,N_12442);
nand U14340 (N_14340,N_12044,N_12769);
and U14341 (N_14341,N_13239,N_12901);
nand U14342 (N_14342,N_13352,N_13059);
nand U14343 (N_14343,N_12071,N_13647);
nand U14344 (N_14344,N_13671,N_13460);
nand U14345 (N_14345,N_13383,N_13132);
nor U14346 (N_14346,N_13512,N_13033);
or U14347 (N_14347,N_12972,N_13152);
or U14348 (N_14348,N_13271,N_12831);
or U14349 (N_14349,N_13679,N_13944);
nor U14350 (N_14350,N_13861,N_13888);
nand U14351 (N_14351,N_12535,N_12590);
and U14352 (N_14352,N_12327,N_13974);
xnor U14353 (N_14353,N_13452,N_13477);
or U14354 (N_14354,N_12844,N_12114);
nand U14355 (N_14355,N_12392,N_12820);
nor U14356 (N_14356,N_13814,N_12334);
or U14357 (N_14357,N_12368,N_12191);
xor U14358 (N_14358,N_12314,N_12977);
xnor U14359 (N_14359,N_12315,N_12328);
or U14360 (N_14360,N_12006,N_12290);
nand U14361 (N_14361,N_12560,N_12353);
or U14362 (N_14362,N_12146,N_13965);
nand U14363 (N_14363,N_12882,N_13392);
and U14364 (N_14364,N_12807,N_12998);
xor U14365 (N_14365,N_12558,N_13581);
and U14366 (N_14366,N_12639,N_13709);
nand U14367 (N_14367,N_13029,N_12652);
and U14368 (N_14368,N_12119,N_12005);
nor U14369 (N_14369,N_13223,N_12210);
xor U14370 (N_14370,N_13676,N_12316);
and U14371 (N_14371,N_13037,N_13447);
or U14372 (N_14372,N_13293,N_12352);
nor U14373 (N_14373,N_12213,N_12136);
and U14374 (N_14374,N_13320,N_13620);
nand U14375 (N_14375,N_12032,N_12051);
nand U14376 (N_14376,N_12803,N_12145);
nand U14377 (N_14377,N_12456,N_13520);
or U14378 (N_14378,N_13205,N_13115);
or U14379 (N_14379,N_13257,N_12619);
nor U14380 (N_14380,N_12819,N_13270);
nor U14381 (N_14381,N_13956,N_13379);
nor U14382 (N_14382,N_13865,N_12137);
and U14383 (N_14383,N_12092,N_13942);
nand U14384 (N_14384,N_13466,N_12113);
nand U14385 (N_14385,N_12468,N_13959);
xnor U14386 (N_14386,N_13469,N_13748);
nor U14387 (N_14387,N_12028,N_12216);
or U14388 (N_14388,N_12332,N_13842);
nand U14389 (N_14389,N_12987,N_12566);
nor U14390 (N_14390,N_12140,N_13890);
or U14391 (N_14391,N_13591,N_13710);
nor U14392 (N_14392,N_12847,N_12821);
and U14393 (N_14393,N_13330,N_12700);
and U14394 (N_14394,N_13178,N_12512);
nor U14395 (N_14395,N_12249,N_13825);
nand U14396 (N_14396,N_12932,N_12262);
nand U14397 (N_14397,N_12274,N_13786);
or U14398 (N_14398,N_12307,N_13645);
or U14399 (N_14399,N_13245,N_13505);
nand U14400 (N_14400,N_13589,N_12094);
xor U14401 (N_14401,N_13187,N_12222);
or U14402 (N_14402,N_12964,N_12131);
or U14403 (N_14403,N_12224,N_13445);
or U14404 (N_14404,N_12529,N_12489);
nand U14405 (N_14405,N_13809,N_13459);
xnor U14406 (N_14406,N_12733,N_12087);
nand U14407 (N_14407,N_12709,N_12714);
nand U14408 (N_14408,N_13643,N_13928);
or U14409 (N_14409,N_12237,N_12551);
or U14410 (N_14410,N_12450,N_12425);
and U14411 (N_14411,N_12867,N_13040);
and U14412 (N_14412,N_13027,N_12981);
nor U14413 (N_14413,N_13409,N_12486);
and U14414 (N_14414,N_13658,N_13545);
nand U14415 (N_14415,N_13707,N_13410);
nand U14416 (N_14416,N_13001,N_13451);
or U14417 (N_14417,N_13353,N_13503);
nor U14418 (N_14418,N_12810,N_12503);
and U14419 (N_14419,N_12173,N_12545);
xor U14420 (N_14420,N_12427,N_12559);
and U14421 (N_14421,N_12920,N_12124);
or U14422 (N_14422,N_12235,N_13435);
and U14423 (N_14423,N_12445,N_13290);
nand U14424 (N_14424,N_12852,N_12104);
nand U14425 (N_14425,N_12459,N_13715);
xor U14426 (N_14426,N_13552,N_13291);
nor U14427 (N_14427,N_13278,N_12305);
nor U14428 (N_14428,N_12175,N_12978);
or U14429 (N_14429,N_13751,N_12096);
xnor U14430 (N_14430,N_13093,N_13268);
nand U14431 (N_14431,N_12914,N_12501);
nand U14432 (N_14432,N_13701,N_13242);
nor U14433 (N_14433,N_12781,N_13282);
and U14434 (N_14434,N_13058,N_12297);
xor U14435 (N_14435,N_13624,N_12103);
xnor U14436 (N_14436,N_13084,N_12650);
or U14437 (N_14437,N_12474,N_12660);
nor U14438 (N_14438,N_12654,N_12356);
xnor U14439 (N_14439,N_13052,N_12711);
xnor U14440 (N_14440,N_12367,N_13627);
or U14441 (N_14441,N_12193,N_12031);
xor U14442 (N_14442,N_13444,N_12595);
nor U14443 (N_14443,N_13428,N_12101);
xor U14444 (N_14444,N_13567,N_12064);
and U14445 (N_14445,N_12861,N_12455);
or U14446 (N_14446,N_12066,N_13669);
nor U14447 (N_14447,N_12579,N_13886);
nor U14448 (N_14448,N_13401,N_13406);
or U14449 (N_14449,N_12665,N_13094);
nor U14450 (N_14450,N_13706,N_12825);
nand U14451 (N_14451,N_12112,N_12498);
nand U14452 (N_14452,N_12789,N_12701);
nand U14453 (N_14453,N_13634,N_12567);
and U14454 (N_14454,N_13629,N_12742);
nor U14455 (N_14455,N_13126,N_13517);
and U14456 (N_14456,N_12615,N_13074);
or U14457 (N_14457,N_13243,N_12496);
nand U14458 (N_14458,N_13518,N_12376);
nand U14459 (N_14459,N_12100,N_12063);
xor U14460 (N_14460,N_12563,N_13433);
or U14461 (N_14461,N_13798,N_13501);
or U14462 (N_14462,N_12211,N_12548);
nor U14463 (N_14463,N_13731,N_13838);
nor U14464 (N_14464,N_12398,N_13065);
nand U14465 (N_14465,N_12967,N_12048);
nor U14466 (N_14466,N_12516,N_13200);
xnor U14467 (N_14467,N_12719,N_13199);
or U14468 (N_14468,N_12221,N_13661);
xor U14469 (N_14469,N_13766,N_13345);
xor U14470 (N_14470,N_12586,N_12684);
and U14471 (N_14471,N_13493,N_13371);
nand U14472 (N_14472,N_13536,N_12349);
or U14473 (N_14473,N_12083,N_13356);
or U14474 (N_14474,N_12669,N_13215);
xnor U14475 (N_14475,N_13145,N_13855);
nand U14476 (N_14476,N_13665,N_12657);
nor U14477 (N_14477,N_13426,N_13488);
nand U14478 (N_14478,N_12800,N_12393);
nand U14479 (N_14479,N_12687,N_13907);
nor U14480 (N_14480,N_13994,N_12357);
or U14481 (N_14481,N_13725,N_13078);
xnor U14482 (N_14482,N_13948,N_13219);
xnor U14483 (N_14483,N_13638,N_13124);
nand U14484 (N_14484,N_12582,N_12924);
nand U14485 (N_14485,N_12835,N_13105);
nand U14486 (N_14486,N_13484,N_12265);
nor U14487 (N_14487,N_12366,N_13237);
or U14488 (N_14488,N_13991,N_12537);
or U14489 (N_14489,N_12667,N_13578);
nand U14490 (N_14490,N_12050,N_13694);
and U14491 (N_14491,N_12958,N_13236);
nor U14492 (N_14492,N_12273,N_12913);
and U14493 (N_14493,N_12539,N_12350);
or U14494 (N_14494,N_13453,N_13275);
nand U14495 (N_14495,N_12076,N_13562);
nand U14496 (N_14496,N_13264,N_12562);
or U14497 (N_14497,N_12491,N_13812);
nand U14498 (N_14498,N_12299,N_13762);
or U14499 (N_14499,N_13852,N_12077);
and U14500 (N_14500,N_12444,N_13432);
or U14501 (N_14501,N_12570,N_12982);
nand U14502 (N_14502,N_12208,N_12775);
nor U14503 (N_14503,N_12728,N_12281);
or U14504 (N_14504,N_13478,N_13986);
or U14505 (N_14505,N_12602,N_13790);
nand U14506 (N_14506,N_12526,N_12948);
nor U14507 (N_14507,N_12802,N_12949);
or U14508 (N_14508,N_12606,N_12610);
nor U14509 (N_14509,N_13322,N_13770);
nand U14510 (N_14510,N_13294,N_12374);
and U14511 (N_14511,N_12020,N_12710);
nand U14512 (N_14512,N_13111,N_13121);
xnor U14513 (N_14513,N_12754,N_12832);
nand U14514 (N_14514,N_12738,N_12326);
or U14515 (N_14515,N_13086,N_12471);
nand U14516 (N_14516,N_12518,N_13289);
or U14517 (N_14517,N_13456,N_12763);
or U14518 (N_14518,N_12730,N_12275);
nor U14519 (N_14519,N_12466,N_13375);
or U14520 (N_14520,N_12355,N_12990);
and U14521 (N_14521,N_12756,N_13336);
xnor U14522 (N_14522,N_12938,N_13840);
nor U14523 (N_14523,N_13628,N_13256);
or U14524 (N_14524,N_12846,N_12097);
nor U14525 (N_14525,N_12824,N_13755);
nand U14526 (N_14526,N_12542,N_12375);
nand U14527 (N_14527,N_12593,N_13737);
xor U14528 (N_14528,N_13080,N_13542);
nor U14529 (N_14529,N_13486,N_13702);
nor U14530 (N_14530,N_12571,N_13746);
and U14531 (N_14531,N_12889,N_13761);
nand U14532 (N_14532,N_13043,N_12469);
nor U14533 (N_14533,N_12430,N_12592);
xor U14534 (N_14534,N_12974,N_12300);
nor U14535 (N_14535,N_12871,N_12673);
nor U14536 (N_14536,N_13540,N_13418);
and U14537 (N_14537,N_12786,N_12919);
nor U14538 (N_14538,N_12995,N_13422);
nand U14539 (N_14539,N_12042,N_13010);
xor U14540 (N_14540,N_13498,N_13436);
xor U14541 (N_14541,N_12906,N_12777);
xnor U14542 (N_14542,N_13491,N_13250);
xor U14543 (N_14543,N_12597,N_13795);
nor U14544 (N_14544,N_13118,N_13050);
nor U14545 (N_14545,N_13171,N_12894);
or U14546 (N_14546,N_13631,N_12012);
nand U14547 (N_14547,N_13521,N_13266);
xor U14548 (N_14548,N_13872,N_12758);
and U14549 (N_14549,N_12706,N_13155);
nor U14550 (N_14550,N_12787,N_13718);
and U14551 (N_14551,N_13527,N_12433);
nand U14552 (N_14552,N_12060,N_13769);
and U14553 (N_14553,N_12133,N_12023);
and U14554 (N_14554,N_13811,N_12627);
nor U14555 (N_14555,N_12391,N_13849);
nor U14556 (N_14556,N_13803,N_12387);
xnor U14557 (N_14557,N_12190,N_13524);
nor U14558 (N_14558,N_12377,N_13173);
and U14559 (N_14559,N_13875,N_13984);
nand U14560 (N_14560,N_13964,N_13366);
nand U14561 (N_14561,N_13479,N_12325);
or U14562 (N_14562,N_13053,N_12294);
and U14563 (N_14563,N_12848,N_12635);
or U14564 (N_14564,N_13823,N_13633);
xnor U14565 (N_14565,N_13313,N_12441);
and U14566 (N_14566,N_12038,N_12607);
or U14567 (N_14567,N_12286,N_12321);
and U14568 (N_14568,N_13283,N_12735);
nor U14569 (N_14569,N_13277,N_13642);
or U14570 (N_14570,N_12898,N_12708);
xnor U14571 (N_14571,N_13218,N_13334);
xnor U14572 (N_14572,N_13590,N_13305);
and U14573 (N_14573,N_13670,N_12522);
and U14574 (N_14574,N_13514,N_12014);
nand U14575 (N_14575,N_12613,N_12760);
or U14576 (N_14576,N_12309,N_13358);
and U14577 (N_14577,N_13822,N_13668);
and U14578 (N_14578,N_12916,N_12385);
or U14579 (N_14579,N_12975,N_13750);
nand U14580 (N_14580,N_12093,N_13800);
nor U14581 (N_14581,N_12929,N_12544);
nor U14582 (N_14582,N_13745,N_12497);
and U14583 (N_14583,N_12490,N_13487);
nor U14584 (N_14584,N_12703,N_13880);
or U14585 (N_14585,N_13302,N_13023);
xnor U14586 (N_14586,N_13038,N_13955);
xor U14587 (N_14587,N_13265,N_13935);
xnor U14588 (N_14588,N_12968,N_13324);
xor U14589 (N_14589,N_13077,N_13141);
nor U14590 (N_14590,N_13238,N_12918);
nor U14591 (N_14591,N_13304,N_13031);
xnor U14592 (N_14592,N_13924,N_12409);
xnor U14593 (N_14593,N_13070,N_12343);
xor U14594 (N_14594,N_12118,N_13967);
xnor U14595 (N_14595,N_12729,N_12715);
xor U14596 (N_14596,N_13963,N_13047);
nor U14597 (N_14597,N_12411,N_12318);
or U14598 (N_14598,N_13430,N_13686);
xnor U14599 (N_14599,N_12148,N_12054);
nand U14600 (N_14600,N_13396,N_13363);
xnor U14601 (N_14601,N_12752,N_13415);
and U14602 (N_14602,N_12301,N_13914);
xnor U14603 (N_14603,N_12837,N_12197);
nor U14604 (N_14604,N_13983,N_13120);
nand U14605 (N_14605,N_13559,N_12517);
xnor U14606 (N_14606,N_12415,N_13231);
nand U14607 (N_14607,N_12091,N_12546);
xor U14608 (N_14608,N_12581,N_13815);
or U14609 (N_14609,N_13280,N_13189);
nand U14610 (N_14610,N_12389,N_13349);
nor U14611 (N_14611,N_12888,N_12166);
xnor U14612 (N_14612,N_13878,N_12502);
xor U14613 (N_14613,N_13780,N_12718);
nor U14614 (N_14614,N_12788,N_13569);
and U14615 (N_14615,N_13847,N_13252);
xnor U14616 (N_14616,N_13129,N_13595);
or U14617 (N_14617,N_13966,N_12379);
or U14618 (N_14618,N_13618,N_12897);
or U14619 (N_14619,N_13217,N_13685);
nor U14620 (N_14620,N_13663,N_13112);
or U14621 (N_14621,N_12247,N_12182);
or U14622 (N_14622,N_12616,N_13225);
or U14623 (N_14623,N_13399,N_12394);
xor U14624 (N_14624,N_12229,N_13377);
xnor U14625 (N_14625,N_13839,N_13662);
nand U14626 (N_14626,N_13980,N_13108);
xor U14627 (N_14627,N_13893,N_13623);
xnor U14628 (N_14628,N_13207,N_12648);
or U14629 (N_14629,N_12749,N_13376);
nor U14630 (N_14630,N_13901,N_12508);
or U14631 (N_14631,N_13879,N_13988);
nor U14632 (N_14632,N_12555,N_12663);
nand U14633 (N_14633,N_12236,N_12691);
nor U14634 (N_14634,N_12288,N_13910);
nor U14635 (N_14635,N_12258,N_13741);
and U14636 (N_14636,N_12475,N_12412);
or U14637 (N_14637,N_13533,N_13926);
nor U14638 (N_14638,N_12519,N_12524);
or U14639 (N_14639,N_12792,N_13339);
nor U14640 (N_14640,N_12591,N_12946);
nand U14641 (N_14641,N_13220,N_13934);
nor U14642 (N_14642,N_13744,N_12492);
nand U14643 (N_14643,N_12858,N_12159);
nor U14644 (N_14644,N_12983,N_13835);
or U14645 (N_14645,N_12722,N_12934);
xnor U14646 (N_14646,N_12556,N_13224);
and U14647 (N_14647,N_13169,N_13056);
or U14648 (N_14648,N_13211,N_13018);
and U14649 (N_14649,N_12147,N_12057);
nor U14650 (N_14650,N_12577,N_12157);
nand U14651 (N_14651,N_13600,N_13226);
and U14652 (N_14652,N_13580,N_13088);
nor U14653 (N_14653,N_13850,N_12388);
nand U14654 (N_14654,N_13615,N_13513);
nand U14655 (N_14655,N_13230,N_13854);
or U14656 (N_14656,N_12853,N_12624);
or U14657 (N_14657,N_12483,N_13259);
xnor U14658 (N_14658,N_13100,N_12280);
nand U14659 (N_14659,N_12400,N_13555);
and U14660 (N_14660,N_12935,N_13982);
or U14661 (N_14661,N_12143,N_13232);
xnor U14662 (N_14662,N_13316,N_13034);
and U14663 (N_14663,N_13202,N_13989);
and U14664 (N_14664,N_13196,N_12256);
nand U14665 (N_14665,N_13573,N_13342);
nor U14666 (N_14666,N_13092,N_13025);
or U14667 (N_14667,N_13894,N_12985);
nand U14668 (N_14668,N_12525,N_12495);
or U14669 (N_14669,N_13186,N_13419);
and U14670 (N_14670,N_13816,N_12241);
nor U14671 (N_14671,N_12696,N_13128);
xor U14672 (N_14672,N_13898,N_13135);
nand U14673 (N_14673,N_12679,N_13700);
xor U14674 (N_14674,N_12231,N_12171);
nand U14675 (N_14675,N_12452,N_13343);
or U14676 (N_14676,N_12891,N_12323);
and U14677 (N_14677,N_13987,N_13925);
or U14678 (N_14678,N_13306,N_13832);
and U14679 (N_14679,N_12793,N_13666);
or U14680 (N_14680,N_12670,N_12024);
and U14681 (N_14681,N_13000,N_13650);
and U14682 (N_14682,N_12257,N_12554);
nor U14683 (N_14683,N_12481,N_12917);
and U14684 (N_14684,N_12900,N_12464);
and U14685 (N_14685,N_13626,N_12941);
nor U14686 (N_14686,N_12465,N_13782);
nor U14687 (N_14687,N_12783,N_12001);
and U14688 (N_14688,N_12661,N_13566);
xnor U14689 (N_14689,N_12956,N_13708);
or U14690 (N_14690,N_12283,N_13246);
nor U14691 (N_14691,N_12945,N_13227);
nand U14692 (N_14692,N_13857,N_13119);
or U14693 (N_14693,N_12771,N_13719);
and U14694 (N_14694,N_13919,N_12842);
xor U14695 (N_14695,N_12304,N_12268);
nand U14696 (N_14696,N_13499,N_13998);
nor U14697 (N_14697,N_13528,N_13834);
nor U14698 (N_14698,N_12179,N_12149);
and U14699 (N_14699,N_12731,N_12078);
xor U14700 (N_14700,N_12230,N_13181);
or U14701 (N_14701,N_13494,N_13317);
xnor U14702 (N_14702,N_12185,N_13979);
nand U14703 (N_14703,N_13036,N_12960);
nand U14704 (N_14704,N_13091,N_12200);
xnor U14705 (N_14705,N_13558,N_12234);
xnor U14706 (N_14706,N_12463,N_13417);
nand U14707 (N_14707,N_12923,N_12217);
nor U14708 (N_14708,N_13597,N_13727);
or U14709 (N_14709,N_13992,N_12105);
or U14710 (N_14710,N_13613,N_13532);
and U14711 (N_14711,N_13244,N_12963);
and U14712 (N_14712,N_12074,N_13693);
nor U14713 (N_14713,N_13175,N_13095);
xor U14714 (N_14714,N_13713,N_12698);
and U14715 (N_14715,N_12043,N_12644);
nand U14716 (N_14716,N_12623,N_12886);
nor U14717 (N_14717,N_12753,N_12099);
and U14718 (N_14718,N_13535,N_13172);
or U14719 (N_14719,N_13607,N_12893);
or U14720 (N_14720,N_12086,N_13308);
nor U14721 (N_14721,N_13680,N_12062);
nand U14722 (N_14722,N_12952,N_13272);
or U14723 (N_14723,N_12324,N_12791);
or U14724 (N_14724,N_12485,N_12599);
and U14725 (N_14725,N_13321,N_12195);
or U14726 (N_14726,N_12341,N_13314);
nor U14727 (N_14727,N_12609,N_12098);
or U14728 (N_14728,N_12209,N_12947);
nand U14729 (N_14729,N_13287,N_13703);
or U14730 (N_14730,N_12823,N_12386);
and U14731 (N_14731,N_13096,N_12285);
and U14732 (N_14732,N_13049,N_12574);
xnor U14733 (N_14733,N_12251,N_12035);
xnor U14734 (N_14734,N_13667,N_12202);
and U14735 (N_14735,N_12473,N_12514);
or U14736 (N_14736,N_13644,N_13170);
and U14737 (N_14737,N_12395,N_13561);
nand U14738 (N_14738,N_12026,N_12641);
or U14739 (N_14739,N_13420,N_12382);
nor U14740 (N_14740,N_13039,N_12282);
nand U14741 (N_14741,N_13716,N_13066);
xor U14742 (N_14742,N_13733,N_13843);
xor U14743 (N_14743,N_13870,N_12814);
and U14744 (N_14744,N_12953,N_12246);
and U14745 (N_14745,N_12418,N_12158);
or U14746 (N_14746,N_12866,N_12816);
nor U14747 (N_14747,N_13395,N_12155);
nand U14748 (N_14748,N_12153,N_13971);
xnor U14749 (N_14749,N_12212,N_12747);
nand U14750 (N_14750,N_12428,N_13586);
or U14751 (N_14751,N_12161,N_13592);
or U14752 (N_14752,N_13061,N_13752);
and U14753 (N_14753,N_13194,N_13556);
xor U14754 (N_14754,N_13326,N_12111);
or U14755 (N_14755,N_12564,N_13361);
nand U14756 (N_14756,N_12138,N_13364);
nor U14757 (N_14757,N_13688,N_12359);
nand U14758 (N_14758,N_13859,N_12365);
nor U14759 (N_14759,N_13678,N_12785);
nor U14760 (N_14760,N_12540,N_12381);
nor U14761 (N_14761,N_13262,N_13891);
and U14762 (N_14762,N_13829,N_13403);
and U14763 (N_14763,N_12238,N_12585);
nor U14764 (N_14764,N_12289,N_13183);
nand U14765 (N_14765,N_13076,N_13515);
and U14766 (N_14766,N_13019,N_13163);
nor U14767 (N_14767,N_13279,N_12682);
or U14768 (N_14768,N_13949,N_12561);
and U14769 (N_14769,N_13206,N_13055);
xnor U14770 (N_14770,N_12223,N_12380);
and U14771 (N_14771,N_13354,N_12018);
and U14772 (N_14772,N_13391,N_13848);
or U14773 (N_14773,N_12580,N_12494);
nand U14774 (N_14774,N_13198,N_12340);
xnor U14775 (N_14775,N_13877,N_13960);
nand U14776 (N_14776,N_13307,N_13804);
or U14777 (N_14777,N_13826,N_12487);
nor U14778 (N_14778,N_12488,N_13438);
nand U14779 (N_14779,N_12196,N_12172);
xor U14780 (N_14780,N_13810,N_12612);
nor U14781 (N_14781,N_12438,N_13594);
nor U14782 (N_14782,N_13975,N_12080);
or U14783 (N_14783,N_12576,N_13474);
nand U14784 (N_14784,N_12890,N_12784);
nor U14785 (N_14785,N_12319,N_13193);
or U14786 (N_14786,N_13002,N_12870);
or U14787 (N_14787,N_13851,N_12840);
nor U14788 (N_14788,N_12513,N_12980);
nor U14789 (N_14789,N_13797,N_12649);
xor U14790 (N_14790,N_13483,N_12705);
nand U14791 (N_14791,N_12240,N_13337);
nand U14792 (N_14792,N_13712,N_12575);
nand U14793 (N_14793,N_12292,N_13722);
nand U14794 (N_14794,N_13611,N_12674);
and U14795 (N_14795,N_13546,N_13726);
nor U14796 (N_14796,N_13134,N_12736);
nand U14797 (N_14797,N_13828,N_12019);
nor U14798 (N_14798,N_12693,N_12040);
xor U14799 (N_14799,N_12895,N_12127);
xnor U14800 (N_14800,N_13021,N_13721);
xor U14801 (N_14801,N_12988,N_13423);
xor U14802 (N_14802,N_12029,N_13373);
and U14803 (N_14803,N_13791,N_13619);
nor U14804 (N_14804,N_12095,N_12088);
nor U14805 (N_14805,N_13553,N_12396);
xor U14806 (N_14806,N_13672,N_13006);
xnor U14807 (N_14807,N_13374,N_13174);
xor U14808 (N_14808,N_12121,N_13900);
nor U14809 (N_14809,N_12184,N_12322);
nand U14810 (N_14810,N_12986,N_13362);
nor U14811 (N_14811,N_12070,N_13860);
xnor U14812 (N_14812,N_13468,N_13785);
and U14813 (N_14813,N_12443,N_12424);
nor U14814 (N_14814,N_13754,N_13013);
xnor U14815 (N_14815,N_13103,N_12390);
xnor U14816 (N_14816,N_13734,N_13897);
nor U14817 (N_14817,N_12013,N_12874);
nand U14818 (N_14818,N_13583,N_13655);
nand U14819 (N_14819,N_12594,N_12572);
nor U14820 (N_14820,N_12804,N_13649);
and U14821 (N_14821,N_12192,N_12278);
nor U14822 (N_14822,N_12036,N_12034);
or U14823 (N_14823,N_12351,N_13544);
xnor U14824 (N_14824,N_13749,N_13641);
nand U14825 (N_14825,N_13585,N_12117);
xor U14826 (N_14826,N_13807,N_13687);
and U14827 (N_14827,N_13610,N_13035);
and U14828 (N_14828,N_13209,N_13538);
nor U14829 (N_14829,N_13526,N_12201);
and U14830 (N_14830,N_13338,N_13085);
xor U14831 (N_14831,N_13425,N_13385);
or U14832 (N_14832,N_12855,N_12992);
nor U14833 (N_14833,N_13148,N_13079);
nand U14834 (N_14834,N_12604,N_13341);
xnor U14835 (N_14835,N_13344,N_13424);
and U14836 (N_14836,N_12139,N_12943);
and U14837 (N_14837,N_13720,N_12107);
or U14838 (N_14838,N_13400,N_13180);
or U14839 (N_14839,N_12243,N_13689);
or U14840 (N_14840,N_13765,N_12721);
xor U14841 (N_14841,N_12167,N_13547);
and U14842 (N_14842,N_12039,N_13764);
or U14843 (N_14843,N_13530,N_12939);
and U14844 (N_14844,N_13297,N_12589);
xnor U14845 (N_14845,N_12750,N_12951);
nor U14846 (N_14846,N_13309,N_12873);
xor U14847 (N_14847,N_12617,N_13664);
and U14848 (N_14848,N_13796,N_12748);
nor U14849 (N_14849,N_12037,N_13331);
or U14850 (N_14850,N_12075,N_13911);
nand U14851 (N_14851,N_13296,N_12069);
or U14852 (N_14852,N_13300,N_13481);
or U14853 (N_14853,N_13346,N_12811);
xnor U14854 (N_14854,N_12621,N_13285);
and U14855 (N_14855,N_13024,N_12678);
nor U14856 (N_14856,N_13260,N_13551);
or U14857 (N_14857,N_13208,N_12476);
xnor U14858 (N_14858,N_13197,N_13621);
and U14859 (N_14859,N_12857,N_12089);
and U14860 (N_14860,N_13605,N_12002);
nand U14861 (N_14861,N_13482,N_12954);
nor U14862 (N_14862,N_13485,N_13637);
and U14863 (N_14863,N_12726,N_13333);
or U14864 (N_14864,N_12081,N_12833);
xnor U14865 (N_14865,N_13705,N_13899);
and U14866 (N_14866,N_12776,N_13506);
nand U14867 (N_14867,N_12017,N_13368);
or U14868 (N_14868,N_13853,N_12859);
nand U14869 (N_14869,N_13519,N_12072);
and U14870 (N_14870,N_13370,N_13778);
xnor U14871 (N_14871,N_12413,N_13704);
nor U14872 (N_14872,N_13381,N_13389);
nor U14873 (N_14873,N_13787,N_12697);
and U14874 (N_14874,N_12165,N_13122);
and U14875 (N_14875,N_13421,N_12743);
nor U14876 (N_14876,N_12931,N_13458);
and U14877 (N_14877,N_13909,N_13249);
nor U14878 (N_14878,N_13999,N_13743);
xor U14879 (N_14879,N_12801,N_12970);
nor U14880 (N_14880,N_12205,N_12796);
nor U14881 (N_14881,N_13794,N_12102);
xnor U14882 (N_14882,N_12448,N_12293);
xor U14883 (N_14883,N_12364,N_13570);
nor U14884 (N_14884,N_12509,N_13281);
or U14885 (N_14885,N_12712,N_13253);
or U14886 (N_14886,N_12928,N_13698);
nand U14887 (N_14887,N_12631,N_13457);
xor U14888 (N_14888,N_13017,N_12829);
or U14889 (N_14889,N_13818,N_12437);
nor U14890 (N_14890,N_12984,N_13429);
nor U14891 (N_14891,N_12642,N_13150);
xor U14892 (N_14892,N_12739,N_12849);
xnor U14893 (N_14893,N_13015,N_13885);
xnor U14894 (N_14894,N_12302,N_13255);
nor U14895 (N_14895,N_13868,N_13472);
nor U14896 (N_14896,N_12439,N_12896);
or U14897 (N_14897,N_12130,N_13329);
or U14898 (N_14898,N_12206,N_13504);
xnor U14899 (N_14899,N_13411,N_12049);
nor U14900 (N_14900,N_12348,N_13951);
xnor U14901 (N_14901,N_13101,N_13327);
or U14902 (N_14902,N_12818,N_12378);
xor U14903 (N_14903,N_12892,N_12168);
nand U14904 (N_14904,N_12123,N_12291);
and U14905 (N_14905,N_13788,N_13292);
xor U14906 (N_14906,N_13970,N_13742);
and U14907 (N_14907,N_12226,N_12384);
and U14908 (N_14908,N_12383,N_13046);
nand U14909 (N_14909,N_13431,N_12160);
nor U14910 (N_14910,N_12360,N_13060);
nor U14911 (N_14911,N_12966,N_13820);
nor U14912 (N_14912,N_13846,N_13450);
nand U14913 (N_14913,N_13603,N_13841);
or U14914 (N_14914,N_13214,N_13067);
nor U14915 (N_14915,N_13109,N_12689);
or U14916 (N_14916,N_12194,N_13908);
or U14917 (N_14917,N_13404,N_12150);
nand U14918 (N_14918,N_13026,N_12755);
or U14919 (N_14919,N_12908,N_13981);
and U14920 (N_14920,N_13775,N_13968);
nor U14921 (N_14921,N_12505,N_13808);
nand U14922 (N_14922,N_12717,N_13543);
nand U14923 (N_14923,N_12681,N_13195);
nand U14924 (N_14924,N_12637,N_12651);
nand U14925 (N_14925,N_12183,N_13784);
nor U14926 (N_14926,N_12569,N_12549);
or U14927 (N_14927,N_12573,N_13802);
nor U14928 (N_14928,N_12207,N_12180);
and U14929 (N_14929,N_13646,N_13817);
or U14930 (N_14930,N_12704,N_13874);
and U14931 (N_14931,N_13863,N_13241);
nand U14932 (N_14932,N_12011,N_12805);
nor U14933 (N_14933,N_12345,N_13143);
or U14934 (N_14934,N_12527,N_12397);
nand U14935 (N_14935,N_12244,N_12868);
and U14936 (N_14936,N_13954,N_12178);
xnor U14937 (N_14937,N_13390,N_12403);
and U14938 (N_14938,N_13539,N_13273);
and U14939 (N_14939,N_12685,N_12277);
nand U14940 (N_14940,N_12135,N_12936);
xor U14941 (N_14941,N_13312,N_12531);
nand U14942 (N_14942,N_13827,N_13471);
nor U14943 (N_14943,N_12780,N_13464);
xnor U14944 (N_14944,N_12472,N_12457);
xnor U14945 (N_14945,N_12420,N_12109);
and U14946 (N_14946,N_12880,N_13813);
or U14947 (N_14947,N_13073,N_13696);
nand U14948 (N_14948,N_13896,N_12046);
nor U14949 (N_14949,N_12883,N_12625);
and U14950 (N_14950,N_12330,N_12461);
and U14951 (N_14951,N_13596,N_13973);
nand U14952 (N_14952,N_13005,N_12110);
nor U14953 (N_14953,N_12144,N_12431);
nor U14954 (N_14954,N_12267,N_12976);
xnor U14955 (N_14955,N_12675,N_12584);
xnor U14956 (N_14956,N_12041,N_13584);
xnor U14957 (N_14957,N_12506,N_13724);
and U14958 (N_14958,N_13534,N_13222);
nand U14959 (N_14959,N_12927,N_12520);
xor U14960 (N_14960,N_12940,N_12773);
or U14961 (N_14961,N_13541,N_12164);
nand U14962 (N_14962,N_12907,N_12862);
nor U14963 (N_14963,N_12128,N_12541);
or U14964 (N_14964,N_12808,N_12333);
nor U14965 (N_14965,N_12815,N_12053);
and U14966 (N_14966,N_13439,N_12344);
nand U14967 (N_14967,N_13774,N_13675);
and U14968 (N_14968,N_12778,N_13167);
or U14969 (N_14969,N_12530,N_13301);
xnor U14970 (N_14970,N_12809,N_13507);
nand U14971 (N_14971,N_13972,N_12812);
nor U14972 (N_14972,N_12186,N_13516);
xnor U14973 (N_14973,N_13165,N_13952);
nor U14974 (N_14974,N_13884,N_12910);
xor U14975 (N_14975,N_12768,N_12084);
nand U14976 (N_14976,N_13990,N_13144);
xor U14977 (N_14977,N_13455,N_13328);
nand U14978 (N_14978,N_13022,N_13295);
or U14979 (N_14979,N_13887,N_12797);
and U14980 (N_14980,N_12761,N_12228);
or U14981 (N_14981,N_12887,N_13179);
and U14982 (N_14982,N_13359,N_13204);
or U14983 (N_14983,N_13357,N_13608);
nor U14984 (N_14984,N_12553,N_13978);
and U14985 (N_14985,N_12218,N_12533);
and U14986 (N_14986,N_12994,N_12745);
nand U14987 (N_14987,N_13263,N_13957);
xor U14988 (N_14988,N_13656,N_12421);
nand U14989 (N_14989,N_12016,N_13149);
xor U14990 (N_14990,N_12177,N_13355);
nor U14991 (N_14991,N_13575,N_13075);
nand U14992 (N_14992,N_12933,N_12405);
nor U14993 (N_14993,N_13767,N_12872);
and U14994 (N_14994,N_13777,N_12543);
or U14995 (N_14995,N_12723,N_12419);
or U14996 (N_14996,N_13529,N_12187);
or U14997 (N_14997,N_13771,N_13819);
nand U14998 (N_14998,N_13856,N_12298);
nor U14999 (N_14999,N_13318,N_12227);
or U15000 (N_15000,N_12504,N_12849);
nor U15001 (N_15001,N_13496,N_13295);
nand U15002 (N_15002,N_13932,N_13995);
xor U15003 (N_15003,N_13045,N_12757);
nor U15004 (N_15004,N_13752,N_12217);
nor U15005 (N_15005,N_12920,N_13485);
or U15006 (N_15006,N_12642,N_12002);
nand U15007 (N_15007,N_13279,N_12481);
nor U15008 (N_15008,N_13250,N_12349);
and U15009 (N_15009,N_13032,N_13726);
nor U15010 (N_15010,N_12953,N_13319);
xnor U15011 (N_15011,N_13021,N_12702);
xnor U15012 (N_15012,N_12571,N_13971);
and U15013 (N_15013,N_13916,N_13727);
nor U15014 (N_15014,N_13682,N_12575);
xor U15015 (N_15015,N_12456,N_13463);
nor U15016 (N_15016,N_12003,N_13398);
xnor U15017 (N_15017,N_12072,N_12291);
nand U15018 (N_15018,N_12958,N_13140);
nand U15019 (N_15019,N_12086,N_13664);
nor U15020 (N_15020,N_13617,N_13376);
xnor U15021 (N_15021,N_12166,N_13486);
or U15022 (N_15022,N_13118,N_12539);
or U15023 (N_15023,N_12221,N_12688);
or U15024 (N_15024,N_13494,N_13260);
xnor U15025 (N_15025,N_12858,N_12567);
nor U15026 (N_15026,N_13404,N_12419);
and U15027 (N_15027,N_13632,N_13637);
or U15028 (N_15028,N_13476,N_13798);
and U15029 (N_15029,N_13008,N_13894);
nor U15030 (N_15030,N_13479,N_13707);
or U15031 (N_15031,N_12586,N_13177);
or U15032 (N_15032,N_13718,N_12094);
nor U15033 (N_15033,N_12488,N_13239);
and U15034 (N_15034,N_13060,N_13018);
nor U15035 (N_15035,N_13833,N_13621);
or U15036 (N_15036,N_12178,N_12831);
nor U15037 (N_15037,N_12144,N_12991);
nor U15038 (N_15038,N_12685,N_13805);
and U15039 (N_15039,N_12060,N_12967);
nand U15040 (N_15040,N_12735,N_13316);
nor U15041 (N_15041,N_12933,N_12469);
xor U15042 (N_15042,N_12544,N_12616);
nor U15043 (N_15043,N_13440,N_13130);
or U15044 (N_15044,N_13165,N_12952);
nor U15045 (N_15045,N_12764,N_13833);
xnor U15046 (N_15046,N_13719,N_13981);
nand U15047 (N_15047,N_13518,N_13086);
or U15048 (N_15048,N_13647,N_12008);
or U15049 (N_15049,N_12913,N_13348);
nor U15050 (N_15050,N_12098,N_13481);
or U15051 (N_15051,N_12009,N_13528);
nor U15052 (N_15052,N_12020,N_12188);
nand U15053 (N_15053,N_13046,N_13602);
xor U15054 (N_15054,N_12269,N_13438);
nor U15055 (N_15055,N_12975,N_12466);
xor U15056 (N_15056,N_12558,N_12981);
or U15057 (N_15057,N_13287,N_13809);
nor U15058 (N_15058,N_12900,N_12423);
or U15059 (N_15059,N_13330,N_12839);
and U15060 (N_15060,N_13771,N_12673);
nor U15061 (N_15061,N_12921,N_13124);
nor U15062 (N_15062,N_13551,N_13131);
and U15063 (N_15063,N_12457,N_12541);
and U15064 (N_15064,N_12497,N_12306);
xor U15065 (N_15065,N_12588,N_12746);
or U15066 (N_15066,N_12849,N_13150);
nor U15067 (N_15067,N_12959,N_13206);
or U15068 (N_15068,N_13346,N_13864);
nand U15069 (N_15069,N_13277,N_12083);
nand U15070 (N_15070,N_12916,N_13165);
or U15071 (N_15071,N_13806,N_13448);
nand U15072 (N_15072,N_12861,N_13776);
xor U15073 (N_15073,N_12088,N_13928);
and U15074 (N_15074,N_13048,N_13652);
nor U15075 (N_15075,N_13249,N_13131);
xor U15076 (N_15076,N_12373,N_13343);
nand U15077 (N_15077,N_12899,N_13316);
or U15078 (N_15078,N_12004,N_13506);
xor U15079 (N_15079,N_12222,N_12774);
and U15080 (N_15080,N_12601,N_13285);
nor U15081 (N_15081,N_12476,N_13590);
or U15082 (N_15082,N_13467,N_13334);
nand U15083 (N_15083,N_12913,N_13945);
and U15084 (N_15084,N_12554,N_12101);
nor U15085 (N_15085,N_13581,N_13977);
and U15086 (N_15086,N_12510,N_12947);
or U15087 (N_15087,N_13472,N_12782);
nand U15088 (N_15088,N_12191,N_13571);
nor U15089 (N_15089,N_12379,N_13208);
and U15090 (N_15090,N_12846,N_13758);
nor U15091 (N_15091,N_13114,N_12731);
and U15092 (N_15092,N_12508,N_12379);
xnor U15093 (N_15093,N_13208,N_13469);
and U15094 (N_15094,N_13261,N_13674);
nand U15095 (N_15095,N_13587,N_12824);
nand U15096 (N_15096,N_12734,N_13647);
or U15097 (N_15097,N_13257,N_12492);
nor U15098 (N_15098,N_12142,N_13124);
nand U15099 (N_15099,N_13804,N_12178);
nand U15100 (N_15100,N_13488,N_13696);
xnor U15101 (N_15101,N_12309,N_12840);
nand U15102 (N_15102,N_12872,N_13255);
or U15103 (N_15103,N_13512,N_13329);
or U15104 (N_15104,N_12790,N_13060);
or U15105 (N_15105,N_12508,N_12873);
or U15106 (N_15106,N_13165,N_13563);
and U15107 (N_15107,N_13385,N_13105);
nor U15108 (N_15108,N_13233,N_13133);
or U15109 (N_15109,N_12973,N_12314);
nor U15110 (N_15110,N_13359,N_13302);
xnor U15111 (N_15111,N_12721,N_12776);
or U15112 (N_15112,N_13498,N_12097);
nor U15113 (N_15113,N_12741,N_13043);
nor U15114 (N_15114,N_12914,N_13680);
nor U15115 (N_15115,N_12269,N_13163);
nor U15116 (N_15116,N_12790,N_13108);
and U15117 (N_15117,N_12308,N_12995);
nand U15118 (N_15118,N_12329,N_13637);
and U15119 (N_15119,N_12167,N_12902);
nand U15120 (N_15120,N_12164,N_12971);
or U15121 (N_15121,N_12287,N_12981);
and U15122 (N_15122,N_13298,N_13884);
nand U15123 (N_15123,N_12981,N_13419);
or U15124 (N_15124,N_12375,N_12120);
xnor U15125 (N_15125,N_13770,N_13477);
and U15126 (N_15126,N_13186,N_13192);
nand U15127 (N_15127,N_12605,N_12881);
or U15128 (N_15128,N_12487,N_13693);
and U15129 (N_15129,N_13223,N_13940);
nand U15130 (N_15130,N_12365,N_13870);
nand U15131 (N_15131,N_13652,N_13847);
xor U15132 (N_15132,N_13214,N_13253);
and U15133 (N_15133,N_13623,N_13495);
and U15134 (N_15134,N_12737,N_12330);
or U15135 (N_15135,N_13304,N_12128);
nand U15136 (N_15136,N_12753,N_13109);
xnor U15137 (N_15137,N_13681,N_13751);
and U15138 (N_15138,N_13063,N_12238);
nand U15139 (N_15139,N_13589,N_12584);
xnor U15140 (N_15140,N_13292,N_12662);
and U15141 (N_15141,N_12328,N_13252);
nor U15142 (N_15142,N_12993,N_12348);
or U15143 (N_15143,N_13535,N_13393);
xnor U15144 (N_15144,N_12915,N_12925);
or U15145 (N_15145,N_12624,N_13498);
xor U15146 (N_15146,N_12577,N_12398);
xnor U15147 (N_15147,N_13330,N_13743);
and U15148 (N_15148,N_12079,N_13429);
xnor U15149 (N_15149,N_12880,N_12438);
and U15150 (N_15150,N_12211,N_13814);
and U15151 (N_15151,N_12169,N_13568);
or U15152 (N_15152,N_13605,N_13128);
and U15153 (N_15153,N_12676,N_12477);
nor U15154 (N_15154,N_12870,N_12074);
nand U15155 (N_15155,N_13651,N_12241);
xor U15156 (N_15156,N_13601,N_12274);
xnor U15157 (N_15157,N_12498,N_13343);
nor U15158 (N_15158,N_12567,N_13051);
nand U15159 (N_15159,N_12636,N_13424);
or U15160 (N_15160,N_13304,N_12866);
or U15161 (N_15161,N_12121,N_13379);
and U15162 (N_15162,N_13508,N_12432);
or U15163 (N_15163,N_12857,N_13575);
nand U15164 (N_15164,N_13990,N_13135);
xnor U15165 (N_15165,N_13902,N_12771);
xnor U15166 (N_15166,N_13651,N_12572);
or U15167 (N_15167,N_12604,N_13520);
xor U15168 (N_15168,N_13574,N_12766);
xnor U15169 (N_15169,N_12517,N_12571);
nand U15170 (N_15170,N_12599,N_13969);
nor U15171 (N_15171,N_13388,N_13026);
and U15172 (N_15172,N_12519,N_13187);
or U15173 (N_15173,N_12115,N_12808);
or U15174 (N_15174,N_13217,N_12167);
nor U15175 (N_15175,N_13384,N_12729);
or U15176 (N_15176,N_13255,N_12243);
or U15177 (N_15177,N_13850,N_13246);
or U15178 (N_15178,N_12087,N_12664);
nand U15179 (N_15179,N_13049,N_12894);
xor U15180 (N_15180,N_13654,N_12266);
or U15181 (N_15181,N_12002,N_12228);
nand U15182 (N_15182,N_12923,N_13791);
nand U15183 (N_15183,N_13849,N_12989);
or U15184 (N_15184,N_13105,N_13668);
nand U15185 (N_15185,N_13505,N_12633);
nand U15186 (N_15186,N_12101,N_13370);
xor U15187 (N_15187,N_13182,N_13496);
or U15188 (N_15188,N_12086,N_12080);
nand U15189 (N_15189,N_12331,N_12504);
or U15190 (N_15190,N_12048,N_12542);
nand U15191 (N_15191,N_12209,N_12285);
nor U15192 (N_15192,N_13741,N_13451);
xnor U15193 (N_15193,N_13925,N_13043);
nand U15194 (N_15194,N_12361,N_12339);
or U15195 (N_15195,N_13205,N_13256);
and U15196 (N_15196,N_13506,N_13050);
and U15197 (N_15197,N_13679,N_13756);
nor U15198 (N_15198,N_13158,N_12258);
xnor U15199 (N_15199,N_13319,N_13908);
nand U15200 (N_15200,N_13783,N_12318);
nor U15201 (N_15201,N_12727,N_13586);
or U15202 (N_15202,N_12570,N_13262);
or U15203 (N_15203,N_12079,N_12425);
xnor U15204 (N_15204,N_13878,N_13110);
and U15205 (N_15205,N_12382,N_12010);
xor U15206 (N_15206,N_12450,N_13992);
nor U15207 (N_15207,N_13247,N_12116);
xor U15208 (N_15208,N_13189,N_12618);
and U15209 (N_15209,N_13189,N_12947);
nand U15210 (N_15210,N_12274,N_13200);
or U15211 (N_15211,N_12709,N_12645);
nor U15212 (N_15212,N_13533,N_13294);
nand U15213 (N_15213,N_13780,N_13466);
nor U15214 (N_15214,N_12253,N_13904);
nand U15215 (N_15215,N_12701,N_12174);
nor U15216 (N_15216,N_12005,N_12675);
nor U15217 (N_15217,N_12161,N_13124);
nand U15218 (N_15218,N_13579,N_13994);
or U15219 (N_15219,N_13584,N_12312);
and U15220 (N_15220,N_12877,N_13564);
xnor U15221 (N_15221,N_12686,N_12221);
or U15222 (N_15222,N_13438,N_12699);
and U15223 (N_15223,N_13353,N_13429);
nor U15224 (N_15224,N_12130,N_12498);
nor U15225 (N_15225,N_12633,N_12908);
nor U15226 (N_15226,N_12414,N_13168);
nor U15227 (N_15227,N_12411,N_13651);
nand U15228 (N_15228,N_12691,N_12135);
nor U15229 (N_15229,N_12941,N_13131);
nor U15230 (N_15230,N_13868,N_13072);
and U15231 (N_15231,N_12788,N_12774);
or U15232 (N_15232,N_12592,N_12421);
nor U15233 (N_15233,N_12849,N_12565);
or U15234 (N_15234,N_12824,N_12832);
nand U15235 (N_15235,N_12529,N_12763);
nor U15236 (N_15236,N_12865,N_12592);
and U15237 (N_15237,N_12100,N_12190);
nand U15238 (N_15238,N_13468,N_12611);
xor U15239 (N_15239,N_12373,N_12105);
or U15240 (N_15240,N_13899,N_12918);
nor U15241 (N_15241,N_13433,N_12414);
nor U15242 (N_15242,N_13208,N_12591);
or U15243 (N_15243,N_12708,N_12492);
nand U15244 (N_15244,N_12861,N_13227);
nand U15245 (N_15245,N_13009,N_12637);
nor U15246 (N_15246,N_12518,N_13518);
and U15247 (N_15247,N_13690,N_12298);
nand U15248 (N_15248,N_12941,N_12424);
and U15249 (N_15249,N_13532,N_12692);
or U15250 (N_15250,N_12945,N_13892);
nor U15251 (N_15251,N_13739,N_12306);
nor U15252 (N_15252,N_12588,N_13489);
nor U15253 (N_15253,N_12080,N_12743);
and U15254 (N_15254,N_13879,N_12665);
nand U15255 (N_15255,N_12963,N_12417);
xnor U15256 (N_15256,N_12146,N_13172);
xor U15257 (N_15257,N_13002,N_12533);
xor U15258 (N_15258,N_12710,N_12149);
nand U15259 (N_15259,N_12921,N_12101);
or U15260 (N_15260,N_13901,N_13361);
and U15261 (N_15261,N_13096,N_12790);
and U15262 (N_15262,N_12057,N_12931);
or U15263 (N_15263,N_13278,N_12699);
nor U15264 (N_15264,N_13083,N_13288);
nor U15265 (N_15265,N_12130,N_13185);
nor U15266 (N_15266,N_12374,N_13274);
xor U15267 (N_15267,N_13976,N_12686);
and U15268 (N_15268,N_12460,N_12588);
or U15269 (N_15269,N_13326,N_12619);
and U15270 (N_15270,N_13693,N_12125);
and U15271 (N_15271,N_12938,N_12597);
xor U15272 (N_15272,N_12091,N_12928);
and U15273 (N_15273,N_13230,N_12181);
and U15274 (N_15274,N_13840,N_12611);
or U15275 (N_15275,N_12639,N_13006);
and U15276 (N_15276,N_13672,N_13445);
or U15277 (N_15277,N_12889,N_12910);
xor U15278 (N_15278,N_13251,N_12223);
or U15279 (N_15279,N_13296,N_12519);
or U15280 (N_15280,N_12826,N_13122);
and U15281 (N_15281,N_13873,N_12136);
nand U15282 (N_15282,N_12750,N_12665);
or U15283 (N_15283,N_13469,N_13988);
or U15284 (N_15284,N_13844,N_13277);
or U15285 (N_15285,N_13717,N_12393);
and U15286 (N_15286,N_13681,N_13361);
nor U15287 (N_15287,N_12249,N_12614);
or U15288 (N_15288,N_12427,N_13072);
and U15289 (N_15289,N_13493,N_12525);
nand U15290 (N_15290,N_13097,N_13793);
and U15291 (N_15291,N_12198,N_12896);
nand U15292 (N_15292,N_13684,N_13955);
or U15293 (N_15293,N_12015,N_12134);
nand U15294 (N_15294,N_13854,N_12139);
and U15295 (N_15295,N_13765,N_13232);
nand U15296 (N_15296,N_13454,N_12774);
xor U15297 (N_15297,N_12702,N_12548);
nor U15298 (N_15298,N_12094,N_13103);
xnor U15299 (N_15299,N_13312,N_13721);
nand U15300 (N_15300,N_13837,N_13788);
xnor U15301 (N_15301,N_12911,N_13706);
nor U15302 (N_15302,N_13186,N_12963);
nor U15303 (N_15303,N_13151,N_13543);
xor U15304 (N_15304,N_13357,N_13146);
nand U15305 (N_15305,N_12530,N_13764);
xnor U15306 (N_15306,N_13968,N_13986);
xnor U15307 (N_15307,N_13688,N_12834);
nand U15308 (N_15308,N_13248,N_13404);
nand U15309 (N_15309,N_12690,N_12487);
or U15310 (N_15310,N_12520,N_13354);
nor U15311 (N_15311,N_13522,N_13786);
nand U15312 (N_15312,N_12881,N_13998);
nand U15313 (N_15313,N_12359,N_13647);
xor U15314 (N_15314,N_13018,N_13142);
or U15315 (N_15315,N_13143,N_12241);
or U15316 (N_15316,N_13580,N_13317);
xnor U15317 (N_15317,N_12931,N_13189);
xnor U15318 (N_15318,N_12646,N_12442);
nor U15319 (N_15319,N_12695,N_13863);
xor U15320 (N_15320,N_13694,N_13544);
nor U15321 (N_15321,N_12995,N_12604);
nand U15322 (N_15322,N_12149,N_12401);
and U15323 (N_15323,N_12885,N_12414);
and U15324 (N_15324,N_12579,N_12970);
or U15325 (N_15325,N_12821,N_12558);
nand U15326 (N_15326,N_13981,N_12490);
nor U15327 (N_15327,N_13544,N_12810);
or U15328 (N_15328,N_13153,N_12530);
xnor U15329 (N_15329,N_12803,N_12206);
nand U15330 (N_15330,N_12832,N_13456);
and U15331 (N_15331,N_13889,N_12535);
and U15332 (N_15332,N_12838,N_12840);
nand U15333 (N_15333,N_13973,N_13754);
nor U15334 (N_15334,N_12016,N_13905);
or U15335 (N_15335,N_12673,N_13739);
nor U15336 (N_15336,N_12454,N_12844);
nor U15337 (N_15337,N_12590,N_12572);
or U15338 (N_15338,N_12853,N_12401);
nor U15339 (N_15339,N_13675,N_12494);
xnor U15340 (N_15340,N_12768,N_12680);
and U15341 (N_15341,N_13350,N_13630);
or U15342 (N_15342,N_12540,N_12634);
nand U15343 (N_15343,N_12781,N_13335);
nor U15344 (N_15344,N_13606,N_13972);
nor U15345 (N_15345,N_12709,N_13214);
or U15346 (N_15346,N_12881,N_12355);
nand U15347 (N_15347,N_13175,N_12590);
nor U15348 (N_15348,N_12858,N_12284);
xor U15349 (N_15349,N_13065,N_12069);
nor U15350 (N_15350,N_12528,N_13111);
or U15351 (N_15351,N_12990,N_12607);
or U15352 (N_15352,N_12030,N_12007);
nand U15353 (N_15353,N_12879,N_12883);
nand U15354 (N_15354,N_13732,N_12834);
and U15355 (N_15355,N_12531,N_12223);
xnor U15356 (N_15356,N_13241,N_12079);
and U15357 (N_15357,N_12004,N_13304);
nand U15358 (N_15358,N_12399,N_12236);
or U15359 (N_15359,N_13474,N_13272);
or U15360 (N_15360,N_13638,N_12939);
xor U15361 (N_15361,N_12863,N_13153);
xnor U15362 (N_15362,N_12547,N_12226);
or U15363 (N_15363,N_13682,N_13119);
and U15364 (N_15364,N_13306,N_13837);
and U15365 (N_15365,N_13839,N_12502);
and U15366 (N_15366,N_12450,N_12678);
and U15367 (N_15367,N_13187,N_12320);
nand U15368 (N_15368,N_12505,N_12034);
nor U15369 (N_15369,N_12044,N_13180);
and U15370 (N_15370,N_12895,N_12223);
nor U15371 (N_15371,N_13882,N_12137);
and U15372 (N_15372,N_12541,N_13102);
and U15373 (N_15373,N_13216,N_13365);
nand U15374 (N_15374,N_13896,N_13498);
or U15375 (N_15375,N_13043,N_12936);
nand U15376 (N_15376,N_13878,N_13298);
or U15377 (N_15377,N_12126,N_12620);
nor U15378 (N_15378,N_13427,N_13474);
nand U15379 (N_15379,N_12234,N_12437);
or U15380 (N_15380,N_13293,N_13012);
nand U15381 (N_15381,N_13339,N_12681);
xor U15382 (N_15382,N_13069,N_13864);
or U15383 (N_15383,N_12547,N_12394);
xnor U15384 (N_15384,N_13956,N_13493);
nand U15385 (N_15385,N_12374,N_13831);
nand U15386 (N_15386,N_12498,N_13845);
or U15387 (N_15387,N_12387,N_13777);
or U15388 (N_15388,N_13995,N_13165);
and U15389 (N_15389,N_13214,N_13880);
xnor U15390 (N_15390,N_13822,N_12596);
nand U15391 (N_15391,N_13785,N_12220);
xnor U15392 (N_15392,N_12922,N_13813);
or U15393 (N_15393,N_13311,N_13602);
nor U15394 (N_15394,N_12388,N_12080);
xor U15395 (N_15395,N_13749,N_12509);
xnor U15396 (N_15396,N_13071,N_12843);
nand U15397 (N_15397,N_13457,N_13331);
xor U15398 (N_15398,N_12984,N_12992);
and U15399 (N_15399,N_12291,N_13082);
nor U15400 (N_15400,N_13402,N_13411);
nand U15401 (N_15401,N_13471,N_13648);
and U15402 (N_15402,N_13551,N_13168);
nor U15403 (N_15403,N_12281,N_12878);
nor U15404 (N_15404,N_13128,N_13040);
or U15405 (N_15405,N_12522,N_12749);
nand U15406 (N_15406,N_13124,N_12059);
or U15407 (N_15407,N_13591,N_12492);
xor U15408 (N_15408,N_13578,N_13428);
and U15409 (N_15409,N_13412,N_13183);
or U15410 (N_15410,N_12004,N_12863);
xor U15411 (N_15411,N_12230,N_13589);
nand U15412 (N_15412,N_13031,N_13864);
nand U15413 (N_15413,N_13013,N_13962);
nand U15414 (N_15414,N_13726,N_12042);
or U15415 (N_15415,N_12933,N_12312);
nand U15416 (N_15416,N_12238,N_13249);
or U15417 (N_15417,N_12753,N_13202);
and U15418 (N_15418,N_13235,N_13878);
and U15419 (N_15419,N_13663,N_12689);
and U15420 (N_15420,N_12320,N_12641);
nand U15421 (N_15421,N_13582,N_12093);
and U15422 (N_15422,N_13278,N_12159);
and U15423 (N_15423,N_12602,N_12226);
nor U15424 (N_15424,N_13690,N_12381);
nand U15425 (N_15425,N_13149,N_12340);
xnor U15426 (N_15426,N_12559,N_12571);
and U15427 (N_15427,N_12191,N_13063);
or U15428 (N_15428,N_12715,N_12299);
nor U15429 (N_15429,N_12768,N_12284);
xor U15430 (N_15430,N_13992,N_12465);
and U15431 (N_15431,N_13223,N_13849);
or U15432 (N_15432,N_12583,N_12646);
nand U15433 (N_15433,N_12822,N_13649);
nand U15434 (N_15434,N_13353,N_12916);
and U15435 (N_15435,N_13183,N_12324);
or U15436 (N_15436,N_13272,N_13895);
and U15437 (N_15437,N_13524,N_13558);
nand U15438 (N_15438,N_13538,N_12918);
xor U15439 (N_15439,N_13824,N_12041);
nand U15440 (N_15440,N_12997,N_12741);
and U15441 (N_15441,N_12336,N_12915);
xor U15442 (N_15442,N_13966,N_12430);
xor U15443 (N_15443,N_13070,N_12825);
xor U15444 (N_15444,N_12842,N_12086);
nor U15445 (N_15445,N_13204,N_12234);
and U15446 (N_15446,N_12408,N_13165);
nor U15447 (N_15447,N_12410,N_12927);
and U15448 (N_15448,N_13873,N_13111);
and U15449 (N_15449,N_12848,N_12656);
or U15450 (N_15450,N_13782,N_13359);
nand U15451 (N_15451,N_12685,N_13271);
nor U15452 (N_15452,N_13588,N_13251);
nor U15453 (N_15453,N_12506,N_12276);
nand U15454 (N_15454,N_13451,N_13426);
or U15455 (N_15455,N_13026,N_13919);
xnor U15456 (N_15456,N_13031,N_12416);
nor U15457 (N_15457,N_13795,N_13638);
and U15458 (N_15458,N_12230,N_13896);
nand U15459 (N_15459,N_13934,N_12796);
xor U15460 (N_15460,N_12593,N_13466);
nor U15461 (N_15461,N_12278,N_13206);
xnor U15462 (N_15462,N_13547,N_13031);
nor U15463 (N_15463,N_13149,N_13285);
and U15464 (N_15464,N_13865,N_12758);
and U15465 (N_15465,N_12883,N_13320);
nand U15466 (N_15466,N_12632,N_12063);
and U15467 (N_15467,N_12918,N_12710);
and U15468 (N_15468,N_13824,N_13382);
nand U15469 (N_15469,N_12229,N_13968);
or U15470 (N_15470,N_12334,N_12197);
nand U15471 (N_15471,N_12737,N_13853);
and U15472 (N_15472,N_13219,N_12827);
or U15473 (N_15473,N_12119,N_12850);
and U15474 (N_15474,N_13904,N_12627);
nand U15475 (N_15475,N_13954,N_12025);
or U15476 (N_15476,N_13196,N_12028);
nor U15477 (N_15477,N_12145,N_12031);
and U15478 (N_15478,N_12536,N_13494);
nand U15479 (N_15479,N_13837,N_12593);
and U15480 (N_15480,N_12111,N_13696);
nor U15481 (N_15481,N_13314,N_12663);
xor U15482 (N_15482,N_13762,N_12513);
and U15483 (N_15483,N_12348,N_12124);
and U15484 (N_15484,N_13165,N_13933);
nand U15485 (N_15485,N_12270,N_13757);
nand U15486 (N_15486,N_13327,N_13224);
xnor U15487 (N_15487,N_12980,N_13655);
xor U15488 (N_15488,N_13460,N_12442);
xor U15489 (N_15489,N_13816,N_12361);
nor U15490 (N_15490,N_12146,N_12100);
nor U15491 (N_15491,N_12461,N_13418);
xor U15492 (N_15492,N_13360,N_13014);
nor U15493 (N_15493,N_13463,N_12294);
nor U15494 (N_15494,N_12713,N_12487);
nor U15495 (N_15495,N_13691,N_12482);
nand U15496 (N_15496,N_12412,N_13757);
and U15497 (N_15497,N_12294,N_12307);
nor U15498 (N_15498,N_13534,N_13490);
or U15499 (N_15499,N_13689,N_12426);
and U15500 (N_15500,N_12008,N_13484);
and U15501 (N_15501,N_13279,N_12426);
xor U15502 (N_15502,N_13383,N_12607);
nor U15503 (N_15503,N_13869,N_13461);
and U15504 (N_15504,N_12722,N_13573);
nor U15505 (N_15505,N_12185,N_13279);
nand U15506 (N_15506,N_13557,N_12642);
nand U15507 (N_15507,N_13773,N_12082);
or U15508 (N_15508,N_12325,N_12528);
nand U15509 (N_15509,N_12927,N_13906);
nor U15510 (N_15510,N_12117,N_13199);
xor U15511 (N_15511,N_12829,N_12385);
or U15512 (N_15512,N_13607,N_13831);
xnor U15513 (N_15513,N_13398,N_13360);
xnor U15514 (N_15514,N_12841,N_13350);
or U15515 (N_15515,N_12294,N_12613);
nand U15516 (N_15516,N_13749,N_13308);
nor U15517 (N_15517,N_13879,N_13808);
or U15518 (N_15518,N_13103,N_12715);
nand U15519 (N_15519,N_13688,N_13506);
or U15520 (N_15520,N_13069,N_12018);
and U15521 (N_15521,N_12891,N_12390);
and U15522 (N_15522,N_12529,N_12039);
nor U15523 (N_15523,N_13790,N_12760);
nand U15524 (N_15524,N_12271,N_12229);
and U15525 (N_15525,N_12255,N_13883);
nor U15526 (N_15526,N_13859,N_12110);
or U15527 (N_15527,N_13884,N_12804);
nand U15528 (N_15528,N_13416,N_13626);
xnor U15529 (N_15529,N_12688,N_12651);
nand U15530 (N_15530,N_13899,N_13781);
xnor U15531 (N_15531,N_12048,N_13086);
xnor U15532 (N_15532,N_13845,N_13478);
or U15533 (N_15533,N_12174,N_12945);
or U15534 (N_15534,N_12407,N_13890);
and U15535 (N_15535,N_12940,N_12727);
or U15536 (N_15536,N_13896,N_12842);
xnor U15537 (N_15537,N_13225,N_12775);
xnor U15538 (N_15538,N_13027,N_13631);
or U15539 (N_15539,N_12114,N_13707);
and U15540 (N_15540,N_13995,N_13785);
nor U15541 (N_15541,N_12812,N_13748);
nor U15542 (N_15542,N_12304,N_13694);
and U15543 (N_15543,N_12454,N_12007);
and U15544 (N_15544,N_13628,N_13555);
and U15545 (N_15545,N_12318,N_13276);
nor U15546 (N_15546,N_13477,N_13315);
nor U15547 (N_15547,N_13642,N_13567);
nand U15548 (N_15548,N_13920,N_12664);
nor U15549 (N_15549,N_13601,N_13511);
xnor U15550 (N_15550,N_13206,N_13660);
xor U15551 (N_15551,N_13136,N_12468);
nand U15552 (N_15552,N_12124,N_12423);
and U15553 (N_15553,N_12518,N_13614);
nand U15554 (N_15554,N_13745,N_12643);
xor U15555 (N_15555,N_12830,N_13065);
and U15556 (N_15556,N_13522,N_13353);
xor U15557 (N_15557,N_13229,N_13416);
or U15558 (N_15558,N_12110,N_12229);
xnor U15559 (N_15559,N_12118,N_13555);
nor U15560 (N_15560,N_13621,N_12312);
xor U15561 (N_15561,N_12518,N_13592);
or U15562 (N_15562,N_13855,N_13583);
xnor U15563 (N_15563,N_12528,N_13961);
and U15564 (N_15564,N_13498,N_13550);
nand U15565 (N_15565,N_12290,N_13342);
xnor U15566 (N_15566,N_13029,N_12682);
and U15567 (N_15567,N_12787,N_12117);
and U15568 (N_15568,N_12281,N_13567);
and U15569 (N_15569,N_12566,N_12837);
nor U15570 (N_15570,N_13012,N_13501);
nor U15571 (N_15571,N_12746,N_12912);
or U15572 (N_15572,N_13241,N_12687);
or U15573 (N_15573,N_12768,N_12157);
xnor U15574 (N_15574,N_12043,N_12990);
and U15575 (N_15575,N_12874,N_12158);
nand U15576 (N_15576,N_13734,N_12916);
xor U15577 (N_15577,N_12791,N_12842);
xor U15578 (N_15578,N_13364,N_12033);
and U15579 (N_15579,N_13165,N_12949);
xnor U15580 (N_15580,N_13640,N_13922);
or U15581 (N_15581,N_13312,N_13791);
or U15582 (N_15582,N_13013,N_12105);
nand U15583 (N_15583,N_13493,N_12406);
xor U15584 (N_15584,N_13378,N_13080);
or U15585 (N_15585,N_13561,N_12836);
nor U15586 (N_15586,N_13059,N_13901);
and U15587 (N_15587,N_12278,N_12323);
nand U15588 (N_15588,N_12813,N_13632);
nor U15589 (N_15589,N_12309,N_13506);
and U15590 (N_15590,N_12833,N_13360);
nand U15591 (N_15591,N_12245,N_12491);
xnor U15592 (N_15592,N_12833,N_13847);
nor U15593 (N_15593,N_13309,N_12416);
and U15594 (N_15594,N_13010,N_13604);
nor U15595 (N_15595,N_12450,N_12936);
nor U15596 (N_15596,N_13402,N_13393);
nor U15597 (N_15597,N_13769,N_13011);
and U15598 (N_15598,N_13520,N_13420);
and U15599 (N_15599,N_13005,N_13042);
xor U15600 (N_15600,N_12267,N_13540);
and U15601 (N_15601,N_12889,N_13306);
nand U15602 (N_15602,N_13375,N_12031);
xor U15603 (N_15603,N_12411,N_13056);
and U15604 (N_15604,N_13110,N_13100);
or U15605 (N_15605,N_12075,N_13971);
or U15606 (N_15606,N_13247,N_13347);
nor U15607 (N_15607,N_12538,N_12663);
xor U15608 (N_15608,N_13405,N_12147);
nor U15609 (N_15609,N_12326,N_12691);
xnor U15610 (N_15610,N_13310,N_12820);
xnor U15611 (N_15611,N_12214,N_12479);
nor U15612 (N_15612,N_13834,N_12516);
nand U15613 (N_15613,N_12893,N_12290);
or U15614 (N_15614,N_12596,N_12148);
nor U15615 (N_15615,N_12754,N_12015);
xnor U15616 (N_15616,N_13139,N_13768);
nand U15617 (N_15617,N_13498,N_12290);
and U15618 (N_15618,N_13479,N_13175);
and U15619 (N_15619,N_13727,N_13592);
and U15620 (N_15620,N_12335,N_12195);
nor U15621 (N_15621,N_13411,N_12524);
nand U15622 (N_15622,N_13858,N_12356);
or U15623 (N_15623,N_13751,N_13165);
or U15624 (N_15624,N_13227,N_12493);
and U15625 (N_15625,N_12731,N_13504);
nor U15626 (N_15626,N_13525,N_12947);
nand U15627 (N_15627,N_13822,N_12655);
or U15628 (N_15628,N_13683,N_13818);
nand U15629 (N_15629,N_12413,N_13366);
and U15630 (N_15630,N_12800,N_13758);
nand U15631 (N_15631,N_13022,N_12908);
nor U15632 (N_15632,N_13983,N_13803);
nor U15633 (N_15633,N_12664,N_12461);
and U15634 (N_15634,N_12896,N_12055);
xor U15635 (N_15635,N_12326,N_12780);
nor U15636 (N_15636,N_13578,N_13702);
or U15637 (N_15637,N_13861,N_12190);
xnor U15638 (N_15638,N_13106,N_13286);
nand U15639 (N_15639,N_12098,N_12790);
and U15640 (N_15640,N_13050,N_12768);
and U15641 (N_15641,N_13196,N_12575);
xnor U15642 (N_15642,N_13546,N_12826);
xor U15643 (N_15643,N_12977,N_12614);
nor U15644 (N_15644,N_13517,N_13504);
xor U15645 (N_15645,N_12925,N_12513);
and U15646 (N_15646,N_13448,N_13815);
xor U15647 (N_15647,N_12134,N_12832);
nand U15648 (N_15648,N_13442,N_12102);
xnor U15649 (N_15649,N_13738,N_13177);
xnor U15650 (N_15650,N_12324,N_13893);
and U15651 (N_15651,N_13567,N_13769);
xor U15652 (N_15652,N_13282,N_13798);
and U15653 (N_15653,N_13256,N_12072);
and U15654 (N_15654,N_13774,N_13245);
or U15655 (N_15655,N_13259,N_12656);
or U15656 (N_15656,N_12762,N_13452);
and U15657 (N_15657,N_12594,N_12787);
xnor U15658 (N_15658,N_13946,N_13203);
or U15659 (N_15659,N_12129,N_13905);
or U15660 (N_15660,N_13893,N_13326);
xnor U15661 (N_15661,N_12910,N_13787);
and U15662 (N_15662,N_12611,N_12886);
nor U15663 (N_15663,N_13718,N_12547);
nor U15664 (N_15664,N_13628,N_13258);
and U15665 (N_15665,N_12704,N_13156);
nand U15666 (N_15666,N_12872,N_12205);
nor U15667 (N_15667,N_12998,N_13005);
nor U15668 (N_15668,N_13580,N_13050);
nand U15669 (N_15669,N_12078,N_13482);
and U15670 (N_15670,N_12536,N_12314);
and U15671 (N_15671,N_12394,N_13116);
xor U15672 (N_15672,N_13563,N_12764);
nor U15673 (N_15673,N_13655,N_12080);
xnor U15674 (N_15674,N_12958,N_12739);
nand U15675 (N_15675,N_13453,N_12805);
nor U15676 (N_15676,N_13913,N_12590);
xor U15677 (N_15677,N_12052,N_12774);
xnor U15678 (N_15678,N_13272,N_12278);
nand U15679 (N_15679,N_12989,N_13901);
nand U15680 (N_15680,N_12816,N_12777);
and U15681 (N_15681,N_12415,N_12063);
nand U15682 (N_15682,N_12951,N_12079);
nand U15683 (N_15683,N_12122,N_12493);
and U15684 (N_15684,N_13545,N_12855);
or U15685 (N_15685,N_13415,N_12400);
nand U15686 (N_15686,N_13572,N_12054);
xnor U15687 (N_15687,N_13723,N_13163);
xor U15688 (N_15688,N_13526,N_13323);
xnor U15689 (N_15689,N_12705,N_13160);
xnor U15690 (N_15690,N_12762,N_12878);
or U15691 (N_15691,N_12217,N_12400);
xor U15692 (N_15692,N_12286,N_12304);
nand U15693 (N_15693,N_12685,N_12156);
xnor U15694 (N_15694,N_13446,N_13576);
nor U15695 (N_15695,N_13756,N_13455);
and U15696 (N_15696,N_12992,N_13783);
nand U15697 (N_15697,N_13199,N_13123);
xnor U15698 (N_15698,N_12166,N_12199);
nand U15699 (N_15699,N_13480,N_12492);
and U15700 (N_15700,N_13796,N_12168);
or U15701 (N_15701,N_12406,N_13166);
or U15702 (N_15702,N_12334,N_12980);
nor U15703 (N_15703,N_13033,N_13561);
xor U15704 (N_15704,N_13346,N_12287);
nor U15705 (N_15705,N_13112,N_12259);
nor U15706 (N_15706,N_13619,N_13034);
and U15707 (N_15707,N_12582,N_12454);
or U15708 (N_15708,N_13845,N_13603);
and U15709 (N_15709,N_12293,N_13268);
or U15710 (N_15710,N_12679,N_12636);
xnor U15711 (N_15711,N_13346,N_13414);
xnor U15712 (N_15712,N_13466,N_12144);
nor U15713 (N_15713,N_12413,N_12164);
nor U15714 (N_15714,N_12369,N_13575);
nor U15715 (N_15715,N_12475,N_13490);
nand U15716 (N_15716,N_12649,N_12302);
xor U15717 (N_15717,N_13725,N_12346);
and U15718 (N_15718,N_13829,N_12264);
nand U15719 (N_15719,N_13946,N_13078);
xnor U15720 (N_15720,N_13659,N_12206);
nor U15721 (N_15721,N_13520,N_12121);
xnor U15722 (N_15722,N_12782,N_12131);
nor U15723 (N_15723,N_12771,N_13433);
nor U15724 (N_15724,N_12576,N_13603);
or U15725 (N_15725,N_13100,N_12371);
nand U15726 (N_15726,N_12796,N_12541);
xor U15727 (N_15727,N_12992,N_12908);
xnor U15728 (N_15728,N_13167,N_13858);
and U15729 (N_15729,N_12278,N_13760);
or U15730 (N_15730,N_13228,N_12650);
and U15731 (N_15731,N_13794,N_12841);
nor U15732 (N_15732,N_13665,N_13115);
nand U15733 (N_15733,N_13901,N_12478);
or U15734 (N_15734,N_12847,N_13968);
xor U15735 (N_15735,N_12716,N_12689);
nand U15736 (N_15736,N_13363,N_13427);
xor U15737 (N_15737,N_12909,N_13744);
and U15738 (N_15738,N_13835,N_13240);
and U15739 (N_15739,N_12697,N_13220);
and U15740 (N_15740,N_13077,N_13135);
and U15741 (N_15741,N_12560,N_13989);
nand U15742 (N_15742,N_13178,N_12965);
nand U15743 (N_15743,N_12884,N_13128);
and U15744 (N_15744,N_12897,N_13955);
xnor U15745 (N_15745,N_12528,N_13380);
xnor U15746 (N_15746,N_13831,N_12022);
xnor U15747 (N_15747,N_12627,N_13450);
nand U15748 (N_15748,N_13966,N_13347);
nand U15749 (N_15749,N_13435,N_13451);
nand U15750 (N_15750,N_12739,N_12437);
and U15751 (N_15751,N_13841,N_12134);
xnor U15752 (N_15752,N_12579,N_12745);
xnor U15753 (N_15753,N_13283,N_13648);
nor U15754 (N_15754,N_13081,N_12202);
xnor U15755 (N_15755,N_13149,N_13259);
xnor U15756 (N_15756,N_13504,N_13767);
and U15757 (N_15757,N_12790,N_13782);
nor U15758 (N_15758,N_12320,N_13531);
and U15759 (N_15759,N_12341,N_13913);
or U15760 (N_15760,N_13253,N_12915);
xnor U15761 (N_15761,N_13150,N_13369);
or U15762 (N_15762,N_12003,N_12129);
or U15763 (N_15763,N_13740,N_12031);
or U15764 (N_15764,N_13841,N_12193);
and U15765 (N_15765,N_12473,N_13094);
nand U15766 (N_15766,N_13580,N_13888);
nor U15767 (N_15767,N_13253,N_13597);
and U15768 (N_15768,N_13008,N_12297);
or U15769 (N_15769,N_12211,N_12245);
nand U15770 (N_15770,N_13576,N_13275);
xnor U15771 (N_15771,N_13224,N_13255);
xor U15772 (N_15772,N_12422,N_13538);
xor U15773 (N_15773,N_13381,N_13247);
and U15774 (N_15774,N_13448,N_12751);
xnor U15775 (N_15775,N_12999,N_12150);
and U15776 (N_15776,N_13316,N_13341);
and U15777 (N_15777,N_13945,N_13643);
and U15778 (N_15778,N_12415,N_13675);
nor U15779 (N_15779,N_12173,N_13496);
nor U15780 (N_15780,N_12234,N_12902);
xor U15781 (N_15781,N_13233,N_13903);
nand U15782 (N_15782,N_13820,N_12239);
and U15783 (N_15783,N_12822,N_12577);
nand U15784 (N_15784,N_12790,N_13442);
nor U15785 (N_15785,N_13900,N_12405);
nand U15786 (N_15786,N_12391,N_13039);
nand U15787 (N_15787,N_12246,N_12596);
or U15788 (N_15788,N_12053,N_13596);
and U15789 (N_15789,N_12410,N_13580);
nand U15790 (N_15790,N_13027,N_13455);
and U15791 (N_15791,N_13153,N_12700);
xor U15792 (N_15792,N_12093,N_12069);
nor U15793 (N_15793,N_12649,N_12444);
or U15794 (N_15794,N_12942,N_13690);
xor U15795 (N_15795,N_13443,N_12425);
nor U15796 (N_15796,N_12297,N_12665);
xnor U15797 (N_15797,N_13484,N_13709);
nor U15798 (N_15798,N_13049,N_12568);
or U15799 (N_15799,N_12556,N_12230);
nor U15800 (N_15800,N_13610,N_13444);
and U15801 (N_15801,N_13503,N_13249);
nand U15802 (N_15802,N_12822,N_12476);
and U15803 (N_15803,N_13583,N_13561);
nand U15804 (N_15804,N_12806,N_12299);
xnor U15805 (N_15805,N_12058,N_12299);
and U15806 (N_15806,N_12361,N_12227);
nor U15807 (N_15807,N_13673,N_12632);
and U15808 (N_15808,N_12308,N_13383);
or U15809 (N_15809,N_13934,N_13142);
and U15810 (N_15810,N_13366,N_12724);
nand U15811 (N_15811,N_12100,N_12292);
xor U15812 (N_15812,N_13328,N_13714);
nand U15813 (N_15813,N_12904,N_12445);
nand U15814 (N_15814,N_12495,N_12269);
nor U15815 (N_15815,N_13207,N_12745);
and U15816 (N_15816,N_12694,N_12621);
nor U15817 (N_15817,N_13693,N_13689);
xnor U15818 (N_15818,N_12094,N_12727);
or U15819 (N_15819,N_12669,N_12892);
nand U15820 (N_15820,N_13327,N_12633);
and U15821 (N_15821,N_12084,N_12323);
xnor U15822 (N_15822,N_13799,N_13488);
nor U15823 (N_15823,N_12276,N_12032);
nand U15824 (N_15824,N_12074,N_12152);
nand U15825 (N_15825,N_13275,N_12073);
nand U15826 (N_15826,N_12239,N_12280);
xnor U15827 (N_15827,N_13653,N_12185);
nand U15828 (N_15828,N_13909,N_13132);
nand U15829 (N_15829,N_13676,N_13140);
nand U15830 (N_15830,N_13371,N_12123);
nor U15831 (N_15831,N_13678,N_13167);
or U15832 (N_15832,N_13093,N_12943);
and U15833 (N_15833,N_13463,N_12038);
xnor U15834 (N_15834,N_13951,N_13537);
and U15835 (N_15835,N_13161,N_13719);
nor U15836 (N_15836,N_13877,N_12762);
and U15837 (N_15837,N_12092,N_12668);
or U15838 (N_15838,N_13761,N_13692);
and U15839 (N_15839,N_12968,N_12288);
nand U15840 (N_15840,N_13205,N_12522);
xor U15841 (N_15841,N_13334,N_12952);
or U15842 (N_15842,N_12607,N_13877);
nand U15843 (N_15843,N_12529,N_12118);
nor U15844 (N_15844,N_13529,N_12152);
or U15845 (N_15845,N_12457,N_12952);
xnor U15846 (N_15846,N_13559,N_13223);
and U15847 (N_15847,N_12220,N_12164);
and U15848 (N_15848,N_12787,N_13541);
and U15849 (N_15849,N_13046,N_13896);
nor U15850 (N_15850,N_12572,N_12803);
and U15851 (N_15851,N_12348,N_12251);
nor U15852 (N_15852,N_13755,N_12217);
or U15853 (N_15853,N_12948,N_13472);
and U15854 (N_15854,N_12497,N_13335);
nor U15855 (N_15855,N_13817,N_13643);
or U15856 (N_15856,N_12481,N_13193);
nand U15857 (N_15857,N_13823,N_12904);
xnor U15858 (N_15858,N_12250,N_13145);
and U15859 (N_15859,N_13502,N_12359);
or U15860 (N_15860,N_12811,N_13893);
or U15861 (N_15861,N_13233,N_13193);
nor U15862 (N_15862,N_13960,N_12772);
and U15863 (N_15863,N_13921,N_13641);
or U15864 (N_15864,N_12416,N_12551);
nor U15865 (N_15865,N_13412,N_12391);
nand U15866 (N_15866,N_13643,N_13350);
or U15867 (N_15867,N_13797,N_12053);
or U15868 (N_15868,N_12436,N_13038);
nor U15869 (N_15869,N_13785,N_13930);
or U15870 (N_15870,N_13970,N_12483);
nor U15871 (N_15871,N_12762,N_12621);
xor U15872 (N_15872,N_12560,N_12213);
nand U15873 (N_15873,N_13798,N_13194);
xor U15874 (N_15874,N_13459,N_13290);
nor U15875 (N_15875,N_13136,N_13012);
nand U15876 (N_15876,N_13548,N_13295);
or U15877 (N_15877,N_13525,N_13561);
xor U15878 (N_15878,N_12402,N_12541);
or U15879 (N_15879,N_13560,N_13939);
and U15880 (N_15880,N_12539,N_13453);
and U15881 (N_15881,N_12767,N_12867);
and U15882 (N_15882,N_13874,N_13918);
and U15883 (N_15883,N_13659,N_12335);
or U15884 (N_15884,N_13767,N_13947);
xnor U15885 (N_15885,N_13656,N_12469);
nor U15886 (N_15886,N_13978,N_13293);
or U15887 (N_15887,N_13222,N_12465);
and U15888 (N_15888,N_12338,N_13780);
nor U15889 (N_15889,N_13500,N_13739);
nor U15890 (N_15890,N_12157,N_13996);
or U15891 (N_15891,N_12744,N_13344);
nand U15892 (N_15892,N_13679,N_13787);
nor U15893 (N_15893,N_13947,N_12886);
nor U15894 (N_15894,N_13877,N_12193);
nand U15895 (N_15895,N_13848,N_12208);
xnor U15896 (N_15896,N_13882,N_12532);
nor U15897 (N_15897,N_12017,N_13854);
nand U15898 (N_15898,N_12958,N_13485);
nand U15899 (N_15899,N_13146,N_12730);
nor U15900 (N_15900,N_12007,N_13912);
xnor U15901 (N_15901,N_12137,N_12345);
and U15902 (N_15902,N_13330,N_13126);
xor U15903 (N_15903,N_12917,N_12786);
nor U15904 (N_15904,N_12047,N_12015);
nand U15905 (N_15905,N_12488,N_13198);
nand U15906 (N_15906,N_13069,N_12603);
xnor U15907 (N_15907,N_13109,N_13584);
xnor U15908 (N_15908,N_13731,N_13110);
xor U15909 (N_15909,N_13335,N_12714);
and U15910 (N_15910,N_12171,N_12948);
nor U15911 (N_15911,N_13428,N_12523);
nor U15912 (N_15912,N_12024,N_13026);
nor U15913 (N_15913,N_13422,N_13507);
nand U15914 (N_15914,N_12543,N_13232);
and U15915 (N_15915,N_13953,N_13493);
xor U15916 (N_15916,N_13618,N_12822);
and U15917 (N_15917,N_12824,N_12467);
and U15918 (N_15918,N_13464,N_13495);
nor U15919 (N_15919,N_12610,N_12336);
or U15920 (N_15920,N_13643,N_12817);
or U15921 (N_15921,N_12546,N_12814);
and U15922 (N_15922,N_12344,N_13703);
or U15923 (N_15923,N_13476,N_13525);
xor U15924 (N_15924,N_12600,N_13189);
or U15925 (N_15925,N_13493,N_13351);
xnor U15926 (N_15926,N_12903,N_12924);
or U15927 (N_15927,N_12560,N_13364);
or U15928 (N_15928,N_13260,N_13902);
or U15929 (N_15929,N_12151,N_13861);
nor U15930 (N_15930,N_13111,N_13062);
nand U15931 (N_15931,N_13982,N_12082);
nand U15932 (N_15932,N_12017,N_13743);
and U15933 (N_15933,N_12648,N_13495);
nor U15934 (N_15934,N_12709,N_13791);
xor U15935 (N_15935,N_12119,N_13026);
nor U15936 (N_15936,N_12010,N_12297);
nor U15937 (N_15937,N_12264,N_12565);
and U15938 (N_15938,N_12583,N_12684);
nand U15939 (N_15939,N_13302,N_13679);
and U15940 (N_15940,N_13137,N_13430);
and U15941 (N_15941,N_12785,N_12266);
or U15942 (N_15942,N_12289,N_13084);
nor U15943 (N_15943,N_12296,N_12160);
and U15944 (N_15944,N_12911,N_12252);
or U15945 (N_15945,N_13574,N_12827);
xnor U15946 (N_15946,N_12129,N_13090);
nor U15947 (N_15947,N_13344,N_13433);
or U15948 (N_15948,N_12479,N_13448);
or U15949 (N_15949,N_13947,N_13923);
and U15950 (N_15950,N_13984,N_12679);
and U15951 (N_15951,N_13540,N_13793);
nor U15952 (N_15952,N_13168,N_13045);
xor U15953 (N_15953,N_12975,N_13550);
or U15954 (N_15954,N_13102,N_12841);
xnor U15955 (N_15955,N_13677,N_12239);
and U15956 (N_15956,N_12451,N_13449);
and U15957 (N_15957,N_13946,N_12956);
or U15958 (N_15958,N_12892,N_12980);
nor U15959 (N_15959,N_13651,N_13644);
and U15960 (N_15960,N_13084,N_12366);
or U15961 (N_15961,N_13981,N_13177);
nor U15962 (N_15962,N_12169,N_12822);
xor U15963 (N_15963,N_13613,N_12455);
xor U15964 (N_15964,N_13025,N_13433);
xor U15965 (N_15965,N_12583,N_12980);
or U15966 (N_15966,N_13257,N_13758);
or U15967 (N_15967,N_13008,N_13599);
and U15968 (N_15968,N_12442,N_13033);
nor U15969 (N_15969,N_13903,N_12691);
or U15970 (N_15970,N_12402,N_12361);
or U15971 (N_15971,N_12872,N_13823);
or U15972 (N_15972,N_12581,N_12196);
and U15973 (N_15973,N_13670,N_12095);
nand U15974 (N_15974,N_12779,N_13573);
nor U15975 (N_15975,N_12090,N_13042);
and U15976 (N_15976,N_12400,N_12518);
and U15977 (N_15977,N_13966,N_13394);
and U15978 (N_15978,N_12003,N_12028);
xnor U15979 (N_15979,N_13618,N_13744);
and U15980 (N_15980,N_13844,N_12409);
xnor U15981 (N_15981,N_13933,N_13786);
nand U15982 (N_15982,N_12664,N_12855);
nor U15983 (N_15983,N_12423,N_12886);
and U15984 (N_15984,N_12996,N_12657);
nand U15985 (N_15985,N_12959,N_12836);
xnor U15986 (N_15986,N_12065,N_12423);
nor U15987 (N_15987,N_13482,N_12555);
and U15988 (N_15988,N_12153,N_13475);
nand U15989 (N_15989,N_12385,N_13854);
xor U15990 (N_15990,N_12592,N_12363);
nor U15991 (N_15991,N_13028,N_12123);
nand U15992 (N_15992,N_12939,N_13743);
or U15993 (N_15993,N_12906,N_12750);
and U15994 (N_15994,N_13299,N_13107);
and U15995 (N_15995,N_12679,N_13718);
nor U15996 (N_15996,N_12178,N_12935);
or U15997 (N_15997,N_12040,N_12891);
and U15998 (N_15998,N_13204,N_12006);
nand U15999 (N_15999,N_12220,N_12288);
and U16000 (N_16000,N_14143,N_15873);
nor U16001 (N_16001,N_14173,N_15583);
or U16002 (N_16002,N_14693,N_15530);
and U16003 (N_16003,N_15222,N_15684);
nor U16004 (N_16004,N_15192,N_14784);
or U16005 (N_16005,N_15842,N_15307);
and U16006 (N_16006,N_15831,N_14115);
nor U16007 (N_16007,N_14222,N_15113);
and U16008 (N_16008,N_14291,N_14783);
and U16009 (N_16009,N_14395,N_14365);
nand U16010 (N_16010,N_15762,N_15754);
xnor U16011 (N_16011,N_14512,N_15341);
nand U16012 (N_16012,N_15701,N_14994);
nand U16013 (N_16013,N_14877,N_15315);
and U16014 (N_16014,N_15330,N_14073);
nand U16015 (N_16015,N_15248,N_15058);
or U16016 (N_16016,N_14789,N_14747);
nor U16017 (N_16017,N_14769,N_15279);
nor U16018 (N_16018,N_14616,N_15561);
nor U16019 (N_16019,N_15263,N_14581);
and U16020 (N_16020,N_14309,N_15476);
xor U16021 (N_16021,N_15952,N_14806);
nor U16022 (N_16022,N_14562,N_14648);
xor U16023 (N_16023,N_15611,N_15992);
nand U16024 (N_16024,N_14728,N_15888);
xnor U16025 (N_16025,N_15857,N_14958);
or U16026 (N_16026,N_14154,N_15344);
nor U16027 (N_16027,N_14987,N_14129);
nand U16028 (N_16028,N_14638,N_14724);
nand U16029 (N_16029,N_14428,N_14217);
and U16030 (N_16030,N_15678,N_14518);
nand U16031 (N_16031,N_14766,N_15062);
nor U16032 (N_16032,N_15598,N_14553);
nand U16033 (N_16033,N_15221,N_15320);
nand U16034 (N_16034,N_15504,N_14849);
and U16035 (N_16035,N_14011,N_14328);
nor U16036 (N_16036,N_14055,N_15464);
or U16037 (N_16037,N_14280,N_14490);
or U16038 (N_16038,N_14897,N_14458);
xor U16039 (N_16039,N_15675,N_14070);
nand U16040 (N_16040,N_14271,N_15358);
and U16041 (N_16041,N_15158,N_14858);
or U16042 (N_16042,N_15397,N_14618);
or U16043 (N_16043,N_15503,N_14252);
nor U16044 (N_16044,N_14606,N_15288);
and U16045 (N_16045,N_14323,N_14653);
nand U16046 (N_16046,N_14077,N_15318);
nand U16047 (N_16047,N_14098,N_15081);
nor U16048 (N_16048,N_15702,N_14669);
and U16049 (N_16049,N_15946,N_14981);
nand U16050 (N_16050,N_15989,N_15859);
or U16051 (N_16051,N_14378,N_14471);
xnor U16052 (N_16052,N_14611,N_15641);
or U16053 (N_16053,N_15170,N_14548);
nand U16054 (N_16054,N_14583,N_14937);
nor U16055 (N_16055,N_15677,N_14408);
or U16056 (N_16056,N_15496,N_14838);
nor U16057 (N_16057,N_15132,N_14692);
nand U16058 (N_16058,N_14145,N_15046);
or U16059 (N_16059,N_15932,N_15384);
xor U16060 (N_16060,N_15563,N_14713);
xor U16061 (N_16061,N_15841,N_14028);
and U16062 (N_16062,N_15198,N_14053);
xor U16063 (N_16063,N_14915,N_14676);
xor U16064 (N_16064,N_15728,N_14592);
and U16065 (N_16065,N_15412,N_14570);
and U16066 (N_16066,N_14110,N_15973);
nand U16067 (N_16067,N_15400,N_14440);
and U16068 (N_16068,N_15259,N_15087);
nor U16069 (N_16069,N_14199,N_14847);
and U16070 (N_16070,N_15945,N_15162);
and U16071 (N_16071,N_14060,N_14332);
xnor U16072 (N_16072,N_14065,N_14454);
nor U16073 (N_16073,N_14599,N_15238);
or U16074 (N_16074,N_14739,N_15974);
or U16075 (N_16075,N_15615,N_14141);
nor U16076 (N_16076,N_15981,N_15824);
and U16077 (N_16077,N_15159,N_15997);
xnor U16078 (N_16078,N_14863,N_15930);
nor U16079 (N_16079,N_15001,N_15582);
or U16080 (N_16080,N_14233,N_14084);
and U16081 (N_16081,N_15371,N_14759);
and U16082 (N_16082,N_15217,N_14696);
nand U16083 (N_16083,N_15699,N_15780);
xnor U16084 (N_16084,N_14008,N_14804);
xor U16085 (N_16085,N_14536,N_14552);
nand U16086 (N_16086,N_15244,N_15720);
nor U16087 (N_16087,N_14930,N_14468);
nand U16088 (N_16088,N_14284,N_14232);
nand U16089 (N_16089,N_14620,N_15525);
nor U16090 (N_16090,N_14164,N_14111);
nor U16091 (N_16091,N_15168,N_14515);
xor U16092 (N_16092,N_14615,N_14340);
xor U16093 (N_16093,N_14442,N_14314);
or U16094 (N_16094,N_15196,N_15127);
nor U16095 (N_16095,N_14373,N_15145);
nand U16096 (N_16096,N_14871,N_14659);
nor U16097 (N_16097,N_14596,N_15549);
or U16098 (N_16098,N_15486,N_14102);
nand U16099 (N_16099,N_15816,N_14444);
nor U16100 (N_16100,N_15529,N_15470);
nor U16101 (N_16101,N_15057,N_14758);
nor U16102 (N_16102,N_14630,N_15575);
nor U16103 (N_16103,N_15885,N_14338);
or U16104 (N_16104,N_14027,N_15018);
or U16105 (N_16105,N_14586,N_14076);
nor U16106 (N_16106,N_15960,N_14042);
xor U16107 (N_16107,N_14264,N_14159);
xnor U16108 (N_16108,N_14990,N_14350);
nor U16109 (N_16109,N_14067,N_15707);
nor U16110 (N_16110,N_15580,N_15241);
nand U16111 (N_16111,N_15505,N_15114);
and U16112 (N_16112,N_14075,N_14815);
xnor U16113 (N_16113,N_14526,N_15293);
or U16114 (N_16114,N_15017,N_14870);
and U16115 (N_16115,N_15480,N_14369);
or U16116 (N_16116,N_14297,N_15249);
xnor U16117 (N_16117,N_14014,N_14683);
nand U16118 (N_16118,N_14048,N_14698);
or U16119 (N_16119,N_14349,N_14272);
or U16120 (N_16120,N_14029,N_15578);
or U16121 (N_16121,N_14211,N_15312);
or U16122 (N_16122,N_15668,N_14206);
nor U16123 (N_16123,N_14470,N_15929);
and U16124 (N_16124,N_15370,N_15274);
or U16125 (N_16125,N_15676,N_14776);
or U16126 (N_16126,N_15793,N_14986);
xor U16127 (N_16127,N_14545,N_15447);
xnor U16128 (N_16128,N_15679,N_14608);
nor U16129 (N_16129,N_15513,N_15112);
xor U16130 (N_16130,N_14530,N_14384);
xor U16131 (N_16131,N_14820,N_14226);
nor U16132 (N_16132,N_14472,N_15534);
or U16133 (N_16133,N_15498,N_15009);
xnor U16134 (N_16134,N_14057,N_15607);
and U16135 (N_16135,N_14926,N_15423);
or U16136 (N_16136,N_15507,N_14887);
nor U16137 (N_16137,N_15354,N_15438);
xnor U16138 (N_16138,N_15352,N_15531);
nand U16139 (N_16139,N_15802,N_15305);
and U16140 (N_16140,N_15853,N_15011);
and U16141 (N_16141,N_15855,N_14868);
nor U16142 (N_16142,N_15373,N_15628);
and U16143 (N_16143,N_15581,N_15551);
nor U16144 (N_16144,N_14423,N_15418);
and U16145 (N_16145,N_15220,N_15794);
nor U16146 (N_16146,N_15807,N_15351);
nor U16147 (N_16147,N_15854,N_15879);
xor U16148 (N_16148,N_14017,N_15131);
nor U16149 (N_16149,N_14729,N_14992);
nand U16150 (N_16150,N_15030,N_14263);
and U16151 (N_16151,N_14749,N_15321);
nand U16152 (N_16152,N_14385,N_15382);
nand U16153 (N_16153,N_14100,N_14774);
xor U16154 (N_16154,N_15252,N_15410);
nor U16155 (N_16155,N_15367,N_14565);
and U16156 (N_16156,N_15200,N_14524);
nand U16157 (N_16157,N_15562,N_15008);
nor U16158 (N_16158,N_15253,N_15743);
nor U16159 (N_16159,N_14779,N_14318);
nor U16160 (N_16160,N_14337,N_14595);
nor U16161 (N_16161,N_15075,N_15823);
xor U16162 (N_16162,N_15478,N_14438);
xor U16163 (N_16163,N_15774,N_15887);
nand U16164 (N_16164,N_14517,N_15306);
or U16165 (N_16165,N_15079,N_15564);
or U16166 (N_16166,N_15991,N_15533);
or U16167 (N_16167,N_15124,N_15801);
nor U16168 (N_16168,N_14306,N_15752);
nand U16169 (N_16169,N_14906,N_15905);
and U16170 (N_16170,N_15738,N_14081);
and U16171 (N_16171,N_15744,N_15356);
nand U16172 (N_16172,N_14723,N_14203);
nand U16173 (N_16173,N_15181,N_14354);
xor U16174 (N_16174,N_15556,N_14096);
nor U16175 (N_16175,N_15299,N_14971);
or U16176 (N_16176,N_14273,N_14185);
and U16177 (N_16177,N_14624,N_15043);
or U16178 (N_16178,N_14922,N_15878);
and U16179 (N_16179,N_14507,N_15592);
and U16180 (N_16180,N_14605,N_15000);
nand U16181 (N_16181,N_15349,N_14965);
or U16182 (N_16182,N_15765,N_15800);
and U16183 (N_16183,N_14093,N_14920);
nand U16184 (N_16184,N_14845,N_15185);
xnor U16185 (N_16185,N_14092,N_15674);
xnor U16186 (N_16186,N_14686,N_15602);
nor U16187 (N_16187,N_14621,N_15789);
and U16188 (N_16188,N_14299,N_15023);
and U16189 (N_16189,N_14009,N_14560);
nand U16190 (N_16190,N_14654,N_15179);
xnor U16191 (N_16191,N_15240,N_15108);
and U16192 (N_16192,N_15390,N_14119);
nor U16193 (N_16193,N_15463,N_14039);
nor U16194 (N_16194,N_15117,N_14061);
or U16195 (N_16195,N_14223,N_14956);
nor U16196 (N_16196,N_15646,N_14329);
nor U16197 (N_16197,N_15041,N_14068);
nand U16198 (N_16198,N_14135,N_14945);
xnor U16199 (N_16199,N_14165,N_15385);
nor U16200 (N_16200,N_14695,N_14189);
or U16201 (N_16201,N_14801,N_14258);
xnor U16202 (N_16202,N_14492,N_15756);
or U16203 (N_16203,N_14033,N_15405);
nor U16204 (N_16204,N_14126,N_14546);
nand U16205 (N_16205,N_14416,N_15799);
nor U16206 (N_16206,N_15050,N_14106);
nor U16207 (N_16207,N_14549,N_15007);
nand U16208 (N_16208,N_15912,N_14940);
nor U16209 (N_16209,N_14667,N_15084);
xor U16210 (N_16210,N_14791,N_15022);
or U16211 (N_16211,N_15629,N_14647);
xor U16212 (N_16212,N_14445,N_14991);
or U16213 (N_16213,N_15353,N_15033);
nor U16214 (N_16214,N_15427,N_15931);
xnor U16215 (N_16215,N_15235,N_15663);
or U16216 (N_16216,N_15725,N_14032);
nor U16217 (N_16217,N_14679,N_14020);
xor U16218 (N_16218,N_15748,N_14089);
nor U16219 (N_16219,N_15261,N_15536);
nor U16220 (N_16220,N_14892,N_14368);
nand U16221 (N_16221,N_15559,N_14982);
nand U16222 (N_16222,N_14152,N_14513);
and U16223 (N_16223,N_14673,N_15956);
or U16224 (N_16224,N_15225,N_15610);
or U16225 (N_16225,N_15834,N_14274);
or U16226 (N_16226,N_15517,N_14483);
xor U16227 (N_16227,N_15784,N_15901);
or U16228 (N_16228,N_14382,N_14737);
xnor U16229 (N_16229,N_14699,N_15211);
nand U16230 (N_16230,N_14237,N_15746);
nand U16231 (N_16231,N_14425,N_14959);
xor U16232 (N_16232,N_14883,N_15941);
nand U16233 (N_16233,N_14256,N_14614);
and U16234 (N_16234,N_15500,N_15216);
nor U16235 (N_16235,N_14544,N_14054);
xnor U16236 (N_16236,N_14600,N_15488);
nand U16237 (N_16237,N_14805,N_15052);
xnor U16238 (N_16238,N_15983,N_14246);
nor U16239 (N_16239,N_14109,N_15817);
nor U16240 (N_16240,N_15369,N_15856);
or U16241 (N_16241,N_15361,N_15703);
nand U16242 (N_16242,N_14103,N_14025);
nand U16243 (N_16243,N_15543,N_15666);
xor U16244 (N_16244,N_15467,N_15515);
xnor U16245 (N_16245,N_15173,N_14666);
nand U16246 (N_16246,N_14862,N_14326);
xnor U16247 (N_16247,N_14631,N_15042);
and U16248 (N_16248,N_15366,N_14509);
nor U16249 (N_16249,N_15063,N_15798);
xor U16250 (N_16250,N_15979,N_14912);
xnor U16251 (N_16251,N_15540,N_15565);
nor U16252 (N_16252,N_14743,N_14617);
or U16253 (N_16253,N_14142,N_14215);
and U16254 (N_16254,N_14814,N_14910);
nor U16255 (N_16255,N_14276,N_15501);
or U16256 (N_16256,N_14234,N_15964);
and U16257 (N_16257,N_14591,N_15065);
nor U16258 (N_16258,N_14675,N_15612);
or U16259 (N_16259,N_15465,N_14363);
and U16260 (N_16260,N_15360,N_15411);
or U16261 (N_16261,N_14198,N_15048);
xor U16262 (N_16262,N_15828,N_15446);
nor U16263 (N_16263,N_15524,N_14422);
nor U16264 (N_16264,N_14829,N_15970);
nor U16265 (N_16265,N_15323,N_15242);
xnor U16266 (N_16266,N_15608,N_15922);
xnor U16267 (N_16267,N_15836,N_15589);
nand U16268 (N_16268,N_15039,N_14022);
nand U16269 (N_16269,N_14607,N_14827);
or U16270 (N_16270,N_14787,N_14316);
nor U16271 (N_16271,N_15419,N_14810);
or U16272 (N_16272,N_15335,N_14059);
and U16273 (N_16273,N_15566,N_14872);
and U16274 (N_16274,N_15118,N_14072);
nor U16275 (N_16275,N_14294,N_15276);
nand U16276 (N_16276,N_15440,N_14705);
or U16277 (N_16277,N_15616,N_14455);
and U16278 (N_16278,N_14213,N_14973);
or U16279 (N_16279,N_15100,N_15188);
xnor U16280 (N_16280,N_15790,N_14339);
nand U16281 (N_16281,N_14238,N_14220);
and U16282 (N_16282,N_15268,N_15571);
and U16283 (N_16283,N_15152,N_15685);
or U16284 (N_16284,N_14300,N_14816);
xnor U16285 (N_16285,N_15691,N_15285);
and U16286 (N_16286,N_14101,N_14852);
and U16287 (N_16287,N_14123,N_14936);
or U16288 (N_16288,N_14494,N_15333);
xor U16289 (N_16289,N_15205,N_15429);
nand U16290 (N_16290,N_15587,N_14050);
nor U16291 (N_16291,N_15636,N_14030);
or U16292 (N_16292,N_15437,N_15178);
and U16293 (N_16293,N_15004,N_15825);
xor U16294 (N_16294,N_14813,N_14114);
nor U16295 (N_16295,N_15938,N_14283);
and U16296 (N_16296,N_15758,N_15060);
nand U16297 (N_16297,N_14481,N_15839);
nor U16298 (N_16298,N_15896,N_14535);
nand U16299 (N_16299,N_14043,N_15135);
nor U16300 (N_16300,N_15586,N_15379);
or U16301 (N_16301,N_14998,N_14082);
and U16302 (N_16302,N_15771,N_14935);
xnor U16303 (N_16303,N_14037,N_15814);
or U16304 (N_16304,N_15136,N_14402);
xor U16305 (N_16305,N_15594,N_14904);
nand U16306 (N_16306,N_14094,N_15428);
xor U16307 (N_16307,N_14701,N_14367);
or U16308 (N_16308,N_15313,N_14431);
nand U16309 (N_16309,N_14304,N_15721);
or U16310 (N_16310,N_15325,N_15643);
nor U16311 (N_16311,N_14914,N_14436);
nor U16312 (N_16312,N_15708,N_15413);
nor U16313 (N_16313,N_15819,N_14661);
nand U16314 (N_16314,N_15545,N_14508);
xnor U16315 (N_16315,N_15694,N_14487);
nor U16316 (N_16316,N_14289,N_15404);
and U16317 (N_16317,N_15687,N_15479);
or U16318 (N_16318,N_14480,N_15422);
and U16319 (N_16319,N_14818,N_14225);
nor U16320 (N_16320,N_15346,N_15474);
and U16321 (N_16321,N_15426,N_15913);
nor U16322 (N_16322,N_15085,N_14196);
nor U16323 (N_16323,N_15747,N_14880);
xnor U16324 (N_16324,N_15454,N_15519);
or U16325 (N_16325,N_15891,N_15449);
nand U16326 (N_16326,N_14038,N_15271);
xor U16327 (N_16327,N_15713,N_15368);
xnor U16328 (N_16328,N_14275,N_15729);
or U16329 (N_16329,N_15742,N_14955);
nand U16330 (N_16330,N_14842,N_15680);
nand U16331 (N_16331,N_15852,N_15560);
nand U16332 (N_16332,N_15921,N_15634);
nand U16333 (N_16333,N_14125,N_14603);
xor U16334 (N_16334,N_14828,N_15441);
xnor U16335 (N_16335,N_14832,N_14356);
or U16336 (N_16336,N_14168,N_15209);
nand U16337 (N_16337,N_14551,N_15555);
or U16338 (N_16338,N_15664,N_14898);
nor U16339 (N_16339,N_14441,N_14850);
and U16340 (N_16340,N_14182,N_15201);
or U16341 (N_16341,N_14529,N_14325);
xor U16342 (N_16342,N_14505,N_14015);
or U16343 (N_16343,N_15055,N_15359);
or U16344 (N_16344,N_14456,N_15958);
nand U16345 (N_16345,N_14985,N_15648);
xor U16346 (N_16346,N_15134,N_15402);
xor U16347 (N_16347,N_14303,N_15709);
or U16348 (N_16348,N_14830,N_15254);
and U16349 (N_16349,N_14117,N_15626);
and U16350 (N_16350,N_14889,N_14171);
nor U16351 (N_16351,N_14243,N_14882);
nand U16352 (N_16352,N_15862,N_15767);
nand U16353 (N_16353,N_15133,N_14657);
and U16354 (N_16354,N_15212,N_14231);
or U16355 (N_16355,N_14978,N_14040);
nor U16356 (N_16356,N_15795,N_14878);
xnor U16357 (N_16357,N_14778,N_14269);
nor U16358 (N_16358,N_15980,N_15554);
xnor U16359 (N_16359,N_15881,N_15903);
nand U16360 (N_16360,N_15532,N_15657);
nand U16361 (N_16361,N_15154,N_14241);
and U16362 (N_16362,N_14960,N_15864);
nand U16363 (N_16363,N_15231,N_14194);
nand U16364 (N_16364,N_14939,N_14964);
xnor U16365 (N_16365,N_14873,N_14639);
xor U16366 (N_16366,N_14510,N_14023);
or U16367 (N_16367,N_15053,N_15420);
xnor U16368 (N_16368,N_14286,N_15697);
xor U16369 (N_16369,N_15355,N_15868);
and U16370 (N_16370,N_15787,N_14417);
and U16371 (N_16371,N_14799,N_15914);
nor U16372 (N_16372,N_15094,N_14523);
nor U16373 (N_16373,N_14802,N_15965);
or U16374 (N_16374,N_14166,N_14270);
nor U16375 (N_16375,N_14496,N_14684);
nor U16376 (N_16376,N_15189,N_15923);
nor U16377 (N_16377,N_14736,N_14181);
and U16378 (N_16378,N_15487,N_14645);
nand U16379 (N_16379,N_15658,N_14797);
xor U16380 (N_16380,N_14640,N_14954);
nand U16381 (N_16381,N_15755,N_15593);
and U16382 (N_16382,N_14671,N_15951);
nor U16383 (N_16383,N_15047,N_14907);
or U16384 (N_16384,N_15128,N_15090);
xnor U16385 (N_16385,N_15214,N_15255);
nand U16386 (N_16386,N_15073,N_15020);
or U16387 (N_16387,N_14561,N_14752);
nand U16388 (N_16388,N_15537,N_15967);
and U16389 (N_16389,N_14012,N_14765);
xor U16390 (N_16390,N_14690,N_15723);
or U16391 (N_16391,N_15494,N_14364);
xnor U16392 (N_16392,N_14970,N_14212);
nor U16393 (N_16393,N_15415,N_14909);
and U16394 (N_16394,N_14216,N_15387);
nand U16395 (N_16395,N_14137,N_15326);
nor U16396 (N_16396,N_14834,N_15844);
or U16397 (N_16397,N_15156,N_15781);
or U16398 (N_16398,N_15847,N_15064);
xor U16399 (N_16399,N_14157,N_15822);
nand U16400 (N_16400,N_14896,N_15750);
nand U16401 (N_16401,N_14254,N_14580);
or U16402 (N_16402,N_14178,N_14750);
and U16403 (N_16403,N_14755,N_15028);
nor U16404 (N_16404,N_15138,N_14559);
nor U16405 (N_16405,N_14687,N_15174);
xor U16406 (N_16406,N_15348,N_15630);
nand U16407 (N_16407,N_15682,N_14721);
or U16408 (N_16408,N_14228,N_14895);
nand U16409 (N_16409,N_14116,N_14622);
nand U16410 (N_16410,N_14148,N_14869);
and U16411 (N_16411,N_15683,N_14260);
nand U16412 (N_16412,N_15471,N_14511);
nand U16413 (N_16413,N_15227,N_14179);
and U16414 (N_16414,N_14360,N_15027);
xnor U16415 (N_16415,N_15871,N_15457);
xor U16416 (N_16416,N_14590,N_15870);
nor U16417 (N_16417,N_15432,N_14394);
nor U16418 (N_16418,N_15840,N_14346);
or U16419 (N_16419,N_14831,N_15792);
or U16420 (N_16420,N_15332,N_14812);
nor U16421 (N_16421,N_15727,N_15250);
or U16422 (N_16422,N_14372,N_14183);
nand U16423 (N_16423,N_14821,N_14680);
xnor U16424 (N_16424,N_15786,N_14477);
and U16425 (N_16425,N_15278,N_14533);
and U16426 (N_16426,N_14158,N_15267);
and U16427 (N_16427,N_14598,N_15003);
nor U16428 (N_16428,N_15775,N_14174);
and U16429 (N_16429,N_15233,N_14796);
xnor U16430 (N_16430,N_15761,N_14191);
xnor U16431 (N_16431,N_15074,N_15865);
or U16432 (N_16432,N_15876,N_14239);
nor U16433 (N_16433,N_15538,N_14634);
or U16434 (N_16434,N_15049,N_15130);
and U16435 (N_16435,N_14052,N_15576);
nand U16436 (N_16436,N_14412,N_14826);
and U16437 (N_16437,N_15906,N_15477);
xor U16438 (N_16438,N_15985,N_15187);
and U16439 (N_16439,N_14347,N_15489);
or U16440 (N_16440,N_14947,N_15431);
xnor U16441 (N_16441,N_14180,N_14041);
nor U16442 (N_16442,N_14036,N_15527);
or U16443 (N_16443,N_15948,N_15810);
and U16444 (N_16444,N_15547,N_14730);
nor U16445 (N_16445,N_14884,N_15393);
or U16446 (N_16446,N_14702,N_15652);
nor U16447 (N_16447,N_14780,N_14934);
and U16448 (N_16448,N_15329,N_15898);
and U16449 (N_16449,N_14968,N_15506);
nor U16450 (N_16450,N_15472,N_15161);
nand U16451 (N_16451,N_15199,N_14573);
nand U16452 (N_16452,N_15357,N_15749);
or U16453 (N_16453,N_14207,N_15229);
and U16454 (N_16454,N_14124,N_15882);
nor U16455 (N_16455,N_15462,N_14771);
or U16456 (N_16456,N_15877,N_14415);
xnor U16457 (N_16457,N_15889,N_14208);
xor U16458 (N_16458,N_14662,N_15088);
xor U16459 (N_16459,N_15640,N_15310);
and U16460 (N_16460,N_15025,N_15961);
nor U16461 (N_16461,N_14308,N_15791);
xor U16462 (N_16462,N_14162,N_15482);
and U16463 (N_16463,N_15553,N_15215);
nor U16464 (N_16464,N_15972,N_15649);
nor U16465 (N_16465,N_15191,N_14462);
nand U16466 (N_16466,N_14446,N_14835);
and U16467 (N_16467,N_15631,N_15518);
or U16468 (N_16468,N_14923,N_14761);
and U16469 (N_16469,N_14242,N_14609);
and U16470 (N_16470,N_14643,N_14642);
nand U16471 (N_16471,N_14482,N_14434);
nor U16472 (N_16472,N_15322,N_15491);
or U16473 (N_16473,N_14976,N_15021);
nor U16474 (N_16474,N_15104,N_15751);
nor U16475 (N_16475,N_14962,N_14219);
nand U16476 (N_16476,N_14649,N_14391);
and U16477 (N_16477,N_15510,N_15837);
nand U16478 (N_16478,N_15091,N_14265);
nor U16479 (N_16479,N_14694,N_14860);
xnor U16480 (N_16480,N_14476,N_14195);
or U16481 (N_16481,N_15975,N_15659);
and U16482 (N_16482,N_15275,N_14710);
nor U16483 (N_16483,N_15111,N_14432);
and U16484 (N_16484,N_14380,N_15202);
nand U16485 (N_16485,N_14353,N_14370);
and U16486 (N_16486,N_14227,N_15916);
and U16487 (N_16487,N_14933,N_14576);
or U16488 (N_16488,N_14379,N_14792);
nand U16489 (N_16489,N_14556,N_15436);
xnor U16490 (N_16490,N_14672,N_15095);
and U16491 (N_16491,N_14866,N_14656);
nand U16492 (N_16492,N_14249,N_14668);
nand U16493 (N_16493,N_15552,N_14034);
xor U16494 (N_16494,N_14277,N_14697);
xnor U16495 (N_16495,N_14646,N_15782);
nand U16496 (N_16496,N_14449,N_14578);
xnor U16497 (N_16497,N_15337,N_15895);
xnor U16498 (N_16498,N_15982,N_14295);
or U16499 (N_16499,N_15645,N_14594);
or U16500 (N_16500,N_15899,N_15497);
and U16501 (N_16501,N_14411,N_14230);
xor U16502 (N_16502,N_15971,N_15157);
nand U16503 (N_16503,N_15180,N_14450);
nor U16504 (N_16504,N_15194,N_15508);
and U16505 (N_16505,N_14543,N_14719);
and U16506 (N_16506,N_15123,N_15730);
nor U16507 (N_16507,N_15633,N_15511);
or U16508 (N_16508,N_15175,N_15509);
xnor U16509 (N_16509,N_15006,N_14993);
and U16510 (N_16510,N_15850,N_15942);
nor U16511 (N_16511,N_14756,N_14331);
nand U16512 (N_16512,N_15392,N_14388);
nor U16513 (N_16513,N_15918,N_15213);
nand U16514 (N_16514,N_15599,N_15040);
and U16515 (N_16515,N_15886,N_15298);
xnor U16516 (N_16516,N_15667,N_15714);
and U16517 (N_16517,N_15376,N_14825);
nor U16518 (N_16518,N_15998,N_15987);
or U16519 (N_16519,N_14567,N_15391);
nor U16520 (N_16520,N_15002,N_15732);
nand U16521 (N_16521,N_15141,N_15940);
and U16522 (N_16522,N_15226,N_15317);
nor U16523 (N_16523,N_14901,N_14469);
xor U16524 (N_16524,N_15716,N_15835);
xnor U16525 (N_16525,N_15395,N_14996);
nand U16526 (N_16526,N_14399,N_14785);
xor U16527 (N_16527,N_15093,N_15874);
nor U16528 (N_16528,N_14322,N_14995);
xor U16529 (N_16529,N_14931,N_14851);
nor U16530 (N_16530,N_14501,N_15019);
nor U16531 (N_16531,N_15944,N_15116);
or U16532 (N_16532,N_15848,N_14136);
xor U16533 (N_16533,N_14362,N_14969);
and U16534 (N_16534,N_14886,N_15861);
xor U16535 (N_16535,N_14823,N_14046);
and U16536 (N_16536,N_15502,N_14285);
nand U16537 (N_16537,N_15544,N_15089);
or U16538 (N_16538,N_14035,N_15984);
and U16539 (N_16539,N_14486,N_14540);
and U16540 (N_16540,N_15557,N_15439);
xor U16541 (N_16541,N_15270,N_15639);
and U16542 (N_16542,N_15148,N_14999);
nor U16543 (N_16543,N_15208,N_15803);
nor U16544 (N_16544,N_14405,N_14079);
nor U16545 (N_16545,N_14722,N_14809);
and U16546 (N_16546,N_14049,N_14613);
nand U16547 (N_16547,N_14604,N_14443);
and U16548 (N_16548,N_15069,N_14259);
nor U16549 (N_16549,N_14768,N_15045);
or U16550 (N_16550,N_15378,N_15172);
nand U16551 (N_16551,N_14874,N_15999);
xor U16552 (N_16552,N_14352,N_14400);
or U16553 (N_16553,N_15706,N_15796);
and U16554 (N_16554,N_15590,N_14674);
and U16555 (N_16555,N_14321,N_15588);
nor U16556 (N_16556,N_15469,N_14107);
xnor U16557 (N_16557,N_15818,N_15264);
nor U16558 (N_16558,N_15558,N_14636);
or U16559 (N_16559,N_15813,N_15336);
nand U16560 (N_16560,N_14893,N_15920);
or U16561 (N_16561,N_14112,N_15535);
and U16562 (N_16562,N_14980,N_14537);
nor U16563 (N_16563,N_15219,N_14344);
xnor U16564 (N_16564,N_14514,N_14840);
nor U16565 (N_16565,N_14268,N_14186);
and U16566 (N_16566,N_15722,N_15165);
and U16567 (N_16567,N_15377,N_15110);
nand U16568 (N_16568,N_15830,N_15097);
or U16569 (N_16569,N_14506,N_15160);
or U16570 (N_16570,N_15101,N_14740);
nand U16571 (N_16571,N_14612,N_14058);
nand U16572 (N_16572,N_15365,N_14188);
or U16573 (N_16573,N_14064,N_15204);
and U16574 (N_16574,N_15880,N_14160);
xnor U16575 (N_16575,N_14235,N_15012);
and U16576 (N_16576,N_15234,N_15955);
and U16577 (N_16577,N_14554,N_15651);
and U16578 (N_16578,N_14974,N_15342);
or U16579 (N_16579,N_15036,N_14952);
xor U16580 (N_16580,N_15038,N_15171);
and U16581 (N_16581,N_15808,N_15705);
and U16582 (N_16582,N_14734,N_15939);
or U16583 (N_16583,N_14626,N_14837);
and U16584 (N_16584,N_15031,N_14120);
and U16585 (N_16585,N_14932,N_14313);
nor U16586 (N_16586,N_15875,N_15363);
and U16587 (N_16587,N_14086,N_14885);
xnor U16588 (N_16588,N_15375,N_15236);
nand U16589 (N_16589,N_15327,N_15892);
or U16590 (N_16590,N_15256,N_15733);
or U16591 (N_16591,N_14335,N_14144);
xor U16592 (N_16592,N_14197,N_14464);
xnor U16593 (N_16593,N_14279,N_15228);
nand U16594 (N_16594,N_14499,N_15119);
nand U16595 (N_16595,N_14822,N_15067);
nand U16596 (N_16596,N_14421,N_14881);
or U16597 (N_16597,N_14296,N_15669);
and U16598 (N_16598,N_15289,N_15577);
or U16599 (N_16599,N_14288,N_15061);
xnor U16600 (N_16600,N_14000,N_14738);
or U16601 (N_16601,N_15362,N_15177);
xnor U16602 (N_16602,N_14150,N_15655);
nor U16603 (N_16603,N_14568,N_15456);
and U16604 (N_16604,N_15584,N_14292);
nor U16605 (N_16605,N_15977,N_15010);
nand U16606 (N_16606,N_14013,N_15297);
and U16607 (N_16607,N_14522,N_15035);
or U16608 (N_16608,N_15959,N_14290);
xnor U16609 (N_16609,N_15210,N_14593);
and U16610 (N_16610,N_14044,N_15237);
or U16611 (N_16611,N_15176,N_14807);
and U16612 (N_16612,N_15625,N_14310);
nor U16613 (N_16613,N_14474,N_15126);
or U16614 (N_16614,N_14833,N_14146);
and U16615 (N_16615,N_14045,N_15059);
or U16616 (N_16616,N_15670,N_14967);
nand U16617 (N_16617,N_14311,N_15417);
or U16618 (N_16618,N_14091,N_14374);
nand U16619 (N_16619,N_14966,N_14404);
nand U16620 (N_16620,N_14069,N_14341);
nand U16621 (N_16621,N_14879,N_14095);
xor U16622 (N_16622,N_14711,N_15295);
nor U16623 (N_16623,N_14224,N_14899);
nor U16624 (N_16624,N_14097,N_14278);
and U16625 (N_16625,N_15389,N_15269);
or U16626 (N_16626,N_14972,N_14201);
xnor U16627 (N_16627,N_14836,N_15239);
nor U16628 (N_16628,N_14016,N_14948);
and U16629 (N_16629,N_14193,N_14602);
or U16630 (N_16630,N_15146,N_15778);
nor U16631 (N_16631,N_15121,N_14413);
nand U16632 (N_16632,N_14210,N_15080);
and U16633 (N_16633,N_14005,N_15096);
xnor U16634 (N_16634,N_15169,N_15328);
or U16635 (N_16635,N_15394,N_15129);
nand U16636 (N_16636,N_15883,N_15224);
xnor U16637 (N_16637,N_15672,N_14754);
nor U16638 (N_16638,N_14571,N_15632);
nor U16639 (N_16639,N_15653,N_14018);
nand U16640 (N_16640,N_15186,N_14725);
xor U16641 (N_16641,N_14336,N_15693);
xnor U16642 (N_16642,N_15933,N_15386);
xor U16643 (N_16643,N_14155,N_14541);
or U16644 (N_16644,N_14760,N_14983);
and U16645 (N_16645,N_14927,N_14951);
or U16646 (N_16646,N_14418,N_15245);
or U16647 (N_16647,N_14641,N_14953);
nand U16648 (N_16648,N_14488,N_14420);
and U16649 (N_16649,N_15453,N_15140);
nand U16650 (N_16650,N_15151,N_15398);
nor U16651 (N_16651,N_14732,N_15071);
or U16652 (N_16652,N_15614,N_14677);
nor U16653 (N_16653,N_15860,N_14846);
nor U16654 (N_16654,N_15768,N_15115);
nor U16655 (N_16655,N_14865,N_14890);
or U16656 (N_16656,N_15772,N_15388);
nor U16657 (N_16657,N_14467,N_14714);
nor U16658 (N_16658,N_14921,N_15424);
nand U16659 (N_16659,N_15120,N_15627);
nor U16660 (N_16660,N_14855,N_14282);
or U16661 (N_16661,N_15995,N_15617);
and U16662 (N_16662,N_14848,N_15331);
xnor U16663 (N_16663,N_15724,N_14147);
nand U16664 (N_16664,N_15232,N_14169);
nor U16665 (N_16665,N_15303,N_15414);
xnor U16666 (N_16666,N_15430,N_14478);
nand U16667 (N_16667,N_14085,N_14727);
or U16668 (N_16668,N_14466,N_14876);
or U16669 (N_16669,N_15396,N_15711);
and U16670 (N_16670,N_15704,N_15206);
and U16671 (N_16671,N_15319,N_15757);
xnor U16672 (N_16672,N_15466,N_15686);
or U16673 (N_16673,N_15195,N_14798);
and U16674 (N_16674,N_15015,N_14572);
and U16675 (N_16675,N_15347,N_15143);
xnor U16676 (N_16676,N_14716,N_15448);
xor U16677 (N_16677,N_15719,N_15741);
xnor U16678 (N_16678,N_14495,N_15953);
nand U16679 (N_16679,N_15455,N_14118);
nand U16680 (N_16680,N_15475,N_14459);
nand U16681 (N_16681,N_14493,N_14867);
or U16682 (N_16682,N_15935,N_15978);
nor U16683 (N_16683,N_15766,N_15595);
nor U16684 (N_16684,N_14062,N_15826);
xor U16685 (N_16685,N_14078,N_15294);
or U16686 (N_16686,N_14063,N_14913);
or U16687 (N_16687,N_15805,N_14908);
or U16688 (N_16688,N_15994,N_14504);
nor U16689 (N_16689,N_14715,N_14782);
nor U16690 (N_16690,N_14963,N_14709);
and U16691 (N_16691,N_15277,N_14500);
nor U16692 (N_16692,N_15286,N_15737);
nor U16693 (N_16693,N_14843,N_14623);
or U16694 (N_16694,N_15144,N_14503);
and U16695 (N_16695,N_14733,N_15485);
nor U16696 (N_16696,N_15372,N_15603);
or U16697 (N_16697,N_14824,N_14393);
or U16698 (N_16698,N_14942,N_14139);
or U16699 (N_16699,N_14688,N_14202);
or U16700 (N_16700,N_14975,N_15092);
xor U16701 (N_16701,N_14547,N_15815);
and U16702 (N_16702,N_14997,N_14205);
xor U16703 (N_16703,N_15572,N_15829);
and U16704 (N_16704,N_15024,N_15656);
nand U16705 (N_16705,N_14128,N_14047);
and U16706 (N_16706,N_14475,N_14753);
nor U16707 (N_16707,N_15851,N_15715);
xor U16708 (N_16708,N_14704,N_14087);
or U16709 (N_16709,N_15712,N_15833);
nand U16710 (N_16710,N_14979,N_15218);
and U16711 (N_16711,N_15381,N_14247);
nor U16712 (N_16712,N_14628,N_14984);
or U16713 (N_16713,N_15153,N_14377);
and U16714 (N_16714,N_15163,N_15695);
or U16715 (N_16715,N_15620,N_14989);
nand U16716 (N_16716,N_14396,N_15407);
nand U16717 (N_16717,N_14320,N_15976);
nor U16718 (N_16718,N_14298,N_14651);
nor U16719 (N_16719,N_15434,N_14793);
or U16720 (N_16720,N_15183,N_14961);
xnor U16721 (N_16721,N_15710,N_15314);
nand U16722 (N_16722,N_15621,N_15689);
xor U16723 (N_16723,N_14333,N_15034);
and U16724 (N_16724,N_14266,N_14104);
xnor U16725 (N_16725,N_14917,N_15054);
nor U16726 (N_16726,N_15550,N_15444);
or U16727 (N_16727,N_15125,N_14463);
or U16728 (N_16728,N_14519,N_14664);
nor U16729 (N_16729,N_15812,N_14414);
nor U16730 (N_16730,N_14520,N_15573);
nand U16731 (N_16731,N_15911,N_15334);
and U16732 (N_16732,N_14190,N_15579);
or U16733 (N_16733,N_14527,N_14700);
and U16734 (N_16734,N_14941,N_15867);
nand U16735 (N_16735,N_15644,N_15866);
xor U16736 (N_16736,N_15283,N_15740);
nand U16737 (N_16737,N_14891,N_15696);
nor U16738 (N_16738,N_15613,N_14720);
and U16739 (N_16739,N_15339,N_14703);
nand U16740 (N_16740,N_14489,N_14589);
nor U16741 (N_16741,N_15910,N_14250);
or U16742 (N_16742,N_14542,N_14707);
or U16743 (N_16743,N_14330,N_15654);
and U16744 (N_16744,N_14502,N_15642);
nand U16745 (N_16745,N_15734,N_14019);
nor U16746 (N_16746,N_15207,N_15166);
and U16747 (N_16747,N_14392,N_14397);
xor U16748 (N_16748,N_14491,N_15863);
and U16749 (N_16749,N_14461,N_14448);
or U16750 (N_16750,N_14525,N_15421);
xor U16751 (N_16751,N_15493,N_15150);
nand U16752 (N_16752,N_15302,N_15460);
nand U16753 (N_16753,N_14577,N_15541);
nand U16754 (N_16754,N_15147,N_14138);
nor U16755 (N_16755,N_15452,N_14307);
nor U16756 (N_16756,N_15399,N_15484);
and U16757 (N_16757,N_14358,N_14001);
xor U16758 (N_16758,N_15514,N_14315);
nand U16759 (N_16759,N_14587,N_15528);
nor U16760 (N_16760,N_14127,N_14744);
or U16761 (N_16761,N_15443,N_14031);
xor U16762 (N_16762,N_15316,N_14426);
or U16763 (N_16763,N_14262,N_14864);
and U16764 (N_16764,N_14403,N_14437);
and U16765 (N_16765,N_14539,N_14447);
xor U16766 (N_16766,N_15499,N_15280);
and U16767 (N_16767,N_14343,N_14928);
or U16768 (N_16768,N_14655,N_14943);
xnor U16769 (N_16769,N_15673,N_15996);
or U16770 (N_16770,N_15759,N_14140);
or U16771 (N_16771,N_14433,N_14531);
or U16772 (N_16772,N_15849,N_15962);
nand U16773 (N_16773,N_14175,N_15492);
nand U16774 (N_16774,N_15260,N_14435);
xor U16775 (N_16775,N_15037,N_15343);
xor U16776 (N_16776,N_14944,N_15539);
or U16777 (N_16777,N_14176,N_15937);
nand U16778 (N_16778,N_15570,N_15606);
and U16779 (N_16779,N_14902,N_14248);
nand U16780 (N_16780,N_15601,N_15068);
nand U16781 (N_16781,N_14390,N_14903);
nor U16782 (N_16782,N_15770,N_14841);
nor U16783 (N_16783,N_14788,N_15350);
nor U16784 (N_16784,N_14663,N_14875);
xor U16785 (N_16785,N_15072,N_14071);
or U16786 (N_16786,N_14351,N_14281);
and U16787 (N_16787,N_14597,N_15005);
nand U16788 (N_16788,N_15900,N_14121);
or U16789 (N_16789,N_14427,N_14130);
nor U16790 (N_16790,N_15568,N_14773);
nand U16791 (N_16791,N_15445,N_15406);
xor U16792 (N_16792,N_14361,N_15139);
nor U16793 (N_16793,N_14113,N_15473);
xnor U16794 (N_16794,N_14327,N_15107);
xor U16795 (N_16795,N_14579,N_14163);
nor U16796 (N_16796,N_15243,N_14386);
and U16797 (N_16797,N_14149,N_15257);
and U16798 (N_16798,N_15928,N_14170);
nand U16799 (N_16799,N_14056,N_15523);
xor U16800 (N_16800,N_14861,N_14950);
nor U16801 (N_16801,N_15785,N_15618);
nor U16802 (N_16802,N_14949,N_14665);
xnor U16803 (N_16803,N_15635,N_15731);
and U16804 (N_16804,N_14652,N_14221);
xor U16805 (N_16805,N_14319,N_14460);
and U16806 (N_16806,N_14588,N_15512);
nand U16807 (N_16807,N_14401,N_14745);
nand U16808 (N_16808,N_15623,N_14888);
and U16809 (N_16809,N_14764,N_14083);
and U16810 (N_16810,N_15401,N_14670);
nand U16811 (N_16811,N_14484,N_14122);
nor U16812 (N_16812,N_14660,N_14808);
nor U16813 (N_16813,N_15908,N_15661);
and U16814 (N_16814,N_15692,N_14629);
nor U16815 (N_16815,N_15495,N_15647);
xnor U16816 (N_16816,N_15408,N_15609);
nand U16817 (N_16817,N_14633,N_14557);
and U16818 (N_16818,N_15164,N_15273);
xnor U16819 (N_16819,N_14564,N_14410);
nor U16820 (N_16820,N_15605,N_15308);
or U16821 (N_16821,N_15459,N_15380);
xor U16822 (N_16822,N_15301,N_15056);
and U16823 (N_16823,N_14635,N_14938);
and U16824 (N_16824,N_14708,N_14324);
or U16825 (N_16825,N_15567,N_14900);
nand U16826 (N_16826,N_14627,N_14007);
and U16827 (N_16827,N_14293,N_15934);
nand U16828 (N_16828,N_15776,N_14925);
nand U16829 (N_16829,N_15893,N_14528);
xor U16830 (N_16830,N_14348,N_14419);
nand U16831 (N_16831,N_15665,N_15282);
and U16832 (N_16832,N_14790,N_14905);
nor U16833 (N_16833,N_14726,N_14712);
xnor U16834 (N_16834,N_14498,N_14267);
or U16835 (N_16835,N_14786,N_14859);
and U16836 (N_16836,N_15246,N_14575);
and U16837 (N_16837,N_15290,N_14691);
and U16838 (N_16838,N_15926,N_15258);
nand U16839 (N_16839,N_15433,N_15155);
nand U16840 (N_16840,N_15542,N_14817);
and U16841 (N_16841,N_15600,N_14134);
or U16842 (N_16842,N_15490,N_15909);
nand U16843 (N_16843,N_14566,N_15103);
or U16844 (N_16844,N_14584,N_14929);
and U16845 (N_16845,N_14161,N_14800);
or U16846 (N_16846,N_14024,N_15843);
xnor U16847 (N_16847,N_15142,N_14803);
xnor U16848 (N_16848,N_14479,N_15099);
and U16849 (N_16849,N_14558,N_15622);
and U16850 (N_16850,N_14236,N_14151);
xnor U16851 (N_16851,N_14916,N_15735);
nor U16852 (N_16852,N_15409,N_15364);
or U16853 (N_16853,N_15016,N_14357);
and U16854 (N_16854,N_14582,N_14718);
nor U16855 (N_16855,N_14407,N_14555);
and U16856 (N_16856,N_14424,N_14839);
or U16857 (N_16857,N_14632,N_14601);
nor U16858 (N_16858,N_15838,N_15193);
nand U16859 (N_16859,N_14240,N_14371);
or U16860 (N_16860,N_14429,N_14255);
and U16861 (N_16861,N_14051,N_14658);
nor U16862 (N_16862,N_14132,N_14301);
and U16863 (N_16863,N_15266,N_15223);
or U16864 (N_16864,N_15340,N_15098);
xor U16865 (N_16865,N_14748,N_14619);
and U16866 (N_16866,N_15190,N_15044);
and U16867 (N_16867,N_14685,N_15029);
nor U16868 (N_16868,N_14376,N_14853);
nor U16869 (N_16869,N_14244,N_15739);
or U16870 (N_16870,N_14359,N_14021);
nor U16871 (N_16871,N_15569,N_14757);
nor U16872 (N_16872,N_14105,N_15671);
xor U16873 (N_16873,N_15917,N_15416);
nor U16874 (N_16874,N_14918,N_14066);
nor U16875 (N_16875,N_15884,N_14689);
nor U16876 (N_16876,N_14682,N_15968);
xnor U16877 (N_16877,N_15262,N_15300);
nor U16878 (N_16878,N_14473,N_15638);
nor U16879 (N_16879,N_15435,N_15915);
xor U16880 (N_16880,N_14777,N_14317);
or U16881 (N_16881,N_14977,N_15070);
nand U16882 (N_16882,N_14200,N_15943);
nor U16883 (N_16883,N_14746,N_15265);
and U16884 (N_16884,N_15650,N_14717);
and U16885 (N_16885,N_15788,N_15619);
and U16886 (N_16886,N_15309,N_15949);
nand U16887 (N_16887,N_15604,N_15548);
or U16888 (N_16888,N_15468,N_15820);
nand U16889 (N_16889,N_15718,N_14099);
nand U16890 (N_16890,N_15681,N_14781);
and U16891 (N_16891,N_14811,N_15804);
xnor U16892 (N_16892,N_14398,N_14957);
xnor U16893 (N_16893,N_14532,N_15821);
or U16894 (N_16894,N_15287,N_14006);
nand U16895 (N_16895,N_15442,N_15660);
and U16896 (N_16896,N_14156,N_15450);
nand U16897 (N_16897,N_14534,N_14177);
xnor U16898 (N_16898,N_14911,N_15597);
and U16899 (N_16899,N_15122,N_14406);
nand U16900 (N_16900,N_14770,N_14465);
or U16901 (N_16901,N_15105,N_14763);
nor U16902 (N_16902,N_15717,N_15203);
nor U16903 (N_16903,N_14497,N_14894);
or U16904 (N_16904,N_15291,N_14706);
or U16905 (N_16905,N_14854,N_15988);
or U16906 (N_16906,N_15251,N_15950);
or U16907 (N_16907,N_15963,N_14767);
nor U16908 (N_16908,N_15760,N_15082);
and U16909 (N_16909,N_15066,N_15296);
and U16910 (N_16910,N_15947,N_15451);
nor U16911 (N_16911,N_14762,N_14090);
xor U16912 (N_16912,N_14355,N_14026);
xor U16913 (N_16913,N_15574,N_15014);
nand U16914 (N_16914,N_14002,N_14088);
nor U16915 (N_16915,N_15516,N_14538);
nand U16916 (N_16916,N_15304,N_15924);
nor U16917 (N_16917,N_15521,N_15700);
nor U16918 (N_16918,N_15230,N_15109);
and U16919 (N_16919,N_15458,N_15764);
or U16920 (N_16920,N_14741,N_14650);
nor U16921 (N_16921,N_14919,N_15954);
nand U16922 (N_16922,N_14334,N_14819);
and U16923 (N_16923,N_15596,N_14305);
and U16924 (N_16924,N_15137,N_15324);
or U16925 (N_16925,N_14569,N_14251);
nand U16926 (N_16926,N_14004,N_15522);
nor U16927 (N_16927,N_14010,N_14187);
nand U16928 (N_16928,N_15585,N_14257);
nand U16929 (N_16929,N_14375,N_14453);
xnor U16930 (N_16930,N_15182,N_15846);
and U16931 (N_16931,N_15078,N_15966);
and U16932 (N_16932,N_15897,N_15546);
and U16933 (N_16933,N_14345,N_15936);
xor U16934 (N_16934,N_14637,N_15990);
nor U16935 (N_16935,N_15106,N_15662);
xor U16936 (N_16936,N_15149,N_15925);
nor U16937 (N_16937,N_14563,N_14409);
or U16938 (N_16938,N_14856,N_14133);
and U16939 (N_16939,N_14735,N_15520);
or U16940 (N_16940,N_15083,N_15827);
nand U16941 (N_16941,N_15184,N_14172);
or U16942 (N_16942,N_14080,N_15102);
and U16943 (N_16943,N_14153,N_15957);
xor U16944 (N_16944,N_15832,N_15872);
nor U16945 (N_16945,N_15745,N_15927);
nor U16946 (N_16946,N_14574,N_15247);
xor U16947 (N_16947,N_15637,N_14625);
xor U16948 (N_16948,N_15338,N_14245);
nand U16949 (N_16949,N_14550,N_15809);
nor U16950 (N_16950,N_15783,N_14452);
and U16951 (N_16951,N_15763,N_15902);
nand U16952 (N_16952,N_14204,N_14516);
and U16953 (N_16953,N_14946,N_15167);
xnor U16954 (N_16954,N_15272,N_15013);
nand U16955 (N_16955,N_15076,N_15690);
nand U16956 (N_16956,N_15483,N_15811);
xor U16957 (N_16957,N_14681,N_15526);
or U16958 (N_16958,N_14389,N_14521);
or U16959 (N_16959,N_15051,N_15736);
or U16960 (N_16960,N_14451,N_15481);
or U16961 (N_16961,N_15284,N_15086);
nand U16962 (N_16962,N_14218,N_15032);
xor U16963 (N_16963,N_15726,N_14795);
xor U16964 (N_16964,N_14485,N_14209);
nor U16965 (N_16965,N_14610,N_15806);
nor U16966 (N_16966,N_14214,N_14924);
nand U16967 (N_16967,N_14387,N_15688);
or U16968 (N_16968,N_14383,N_14342);
and U16969 (N_16969,N_14775,N_15425);
nand U16970 (N_16970,N_15894,N_15403);
xnor U16971 (N_16971,N_14184,N_14261);
and U16972 (N_16972,N_14312,N_14988);
and U16973 (N_16973,N_15904,N_15311);
xor U16974 (N_16974,N_15773,N_14253);
nor U16975 (N_16975,N_15993,N_14074);
nor U16976 (N_16976,N_15383,N_15769);
or U16977 (N_16977,N_15753,N_15777);
xor U16978 (N_16978,N_14457,N_14302);
nand U16979 (N_16979,N_15374,N_14366);
and U16980 (N_16980,N_15345,N_14772);
and U16981 (N_16981,N_15969,N_14439);
xor U16982 (N_16982,N_14794,N_14287);
nand U16983 (N_16983,N_15461,N_14003);
xnor U16984 (N_16984,N_14131,N_15591);
and U16985 (N_16985,N_15869,N_14167);
or U16986 (N_16986,N_15779,N_15907);
and U16987 (N_16987,N_14751,N_15986);
nor U16988 (N_16988,N_15292,N_15197);
xor U16989 (N_16989,N_14430,N_14381);
or U16990 (N_16990,N_14644,N_14731);
and U16991 (N_16991,N_15281,N_14678);
or U16992 (N_16992,N_15077,N_14192);
nand U16993 (N_16993,N_14229,N_14844);
nand U16994 (N_16994,N_15797,N_15026);
or U16995 (N_16995,N_15858,N_14742);
xnor U16996 (N_16996,N_14857,N_14108);
or U16997 (N_16997,N_15919,N_15624);
or U16998 (N_16998,N_15698,N_15845);
or U16999 (N_16999,N_14585,N_15890);
nor U17000 (N_17000,N_15264,N_14123);
or U17001 (N_17001,N_15264,N_15009);
nand U17002 (N_17002,N_14927,N_15099);
xnor U17003 (N_17003,N_15447,N_15849);
nor U17004 (N_17004,N_15198,N_15073);
and U17005 (N_17005,N_14903,N_15487);
nor U17006 (N_17006,N_14846,N_15822);
nand U17007 (N_17007,N_15203,N_15976);
nand U17008 (N_17008,N_15123,N_14410);
and U17009 (N_17009,N_14323,N_14088);
xnor U17010 (N_17010,N_14361,N_15424);
nor U17011 (N_17011,N_14140,N_14431);
and U17012 (N_17012,N_15479,N_14003);
xnor U17013 (N_17013,N_15064,N_14564);
and U17014 (N_17014,N_15176,N_14447);
or U17015 (N_17015,N_14661,N_14528);
and U17016 (N_17016,N_14162,N_14155);
and U17017 (N_17017,N_14398,N_14540);
nor U17018 (N_17018,N_14986,N_15113);
or U17019 (N_17019,N_15468,N_14792);
and U17020 (N_17020,N_14159,N_15356);
and U17021 (N_17021,N_14557,N_15648);
xnor U17022 (N_17022,N_14962,N_15024);
xnor U17023 (N_17023,N_14416,N_15683);
xnor U17024 (N_17024,N_15118,N_15330);
and U17025 (N_17025,N_15817,N_14748);
xor U17026 (N_17026,N_14217,N_15356);
nor U17027 (N_17027,N_14410,N_15202);
or U17028 (N_17028,N_15437,N_15210);
and U17029 (N_17029,N_14674,N_14530);
nand U17030 (N_17030,N_15644,N_15778);
and U17031 (N_17031,N_15314,N_15912);
or U17032 (N_17032,N_15703,N_14962);
nand U17033 (N_17033,N_15610,N_14953);
nor U17034 (N_17034,N_15640,N_15727);
nand U17035 (N_17035,N_14589,N_15176);
nand U17036 (N_17036,N_14154,N_14683);
and U17037 (N_17037,N_15814,N_15268);
nand U17038 (N_17038,N_14509,N_15508);
nor U17039 (N_17039,N_15427,N_14858);
and U17040 (N_17040,N_15320,N_14461);
or U17041 (N_17041,N_15203,N_14626);
nand U17042 (N_17042,N_15150,N_14250);
nand U17043 (N_17043,N_14478,N_14785);
nor U17044 (N_17044,N_14733,N_14378);
xor U17045 (N_17045,N_14618,N_14269);
or U17046 (N_17046,N_15717,N_14516);
and U17047 (N_17047,N_14031,N_15089);
nand U17048 (N_17048,N_14652,N_15428);
nor U17049 (N_17049,N_14856,N_14683);
nor U17050 (N_17050,N_15449,N_14020);
nand U17051 (N_17051,N_14813,N_15649);
xnor U17052 (N_17052,N_15596,N_14065);
or U17053 (N_17053,N_15512,N_14425);
and U17054 (N_17054,N_15841,N_15527);
xor U17055 (N_17055,N_14437,N_15648);
xor U17056 (N_17056,N_14370,N_14299);
xor U17057 (N_17057,N_14257,N_14852);
or U17058 (N_17058,N_15324,N_14190);
and U17059 (N_17059,N_15092,N_15609);
nor U17060 (N_17060,N_14847,N_15332);
nand U17061 (N_17061,N_14122,N_15558);
or U17062 (N_17062,N_14668,N_14456);
nor U17063 (N_17063,N_14555,N_14809);
and U17064 (N_17064,N_14204,N_15938);
or U17065 (N_17065,N_15928,N_14116);
or U17066 (N_17066,N_14276,N_14918);
or U17067 (N_17067,N_14267,N_14583);
and U17068 (N_17068,N_15047,N_14254);
xnor U17069 (N_17069,N_15600,N_15310);
xor U17070 (N_17070,N_15278,N_15642);
nor U17071 (N_17071,N_15681,N_15321);
nor U17072 (N_17072,N_15140,N_15306);
nand U17073 (N_17073,N_14690,N_14096);
xnor U17074 (N_17074,N_15946,N_15005);
nor U17075 (N_17075,N_14668,N_15406);
nand U17076 (N_17076,N_15561,N_15340);
xor U17077 (N_17077,N_14634,N_14806);
nor U17078 (N_17078,N_14866,N_14296);
nor U17079 (N_17079,N_15804,N_15638);
and U17080 (N_17080,N_15377,N_14873);
nor U17081 (N_17081,N_15990,N_14109);
and U17082 (N_17082,N_15858,N_14687);
nor U17083 (N_17083,N_14835,N_14592);
and U17084 (N_17084,N_15681,N_14017);
and U17085 (N_17085,N_15448,N_15065);
nand U17086 (N_17086,N_14242,N_14371);
nand U17087 (N_17087,N_14102,N_15650);
nor U17088 (N_17088,N_14373,N_14141);
nand U17089 (N_17089,N_14288,N_15212);
and U17090 (N_17090,N_14398,N_15632);
and U17091 (N_17091,N_15343,N_15464);
and U17092 (N_17092,N_14725,N_14864);
and U17093 (N_17093,N_15448,N_15454);
xnor U17094 (N_17094,N_15352,N_15241);
nor U17095 (N_17095,N_14209,N_15878);
or U17096 (N_17096,N_14496,N_15135);
xnor U17097 (N_17097,N_14152,N_15542);
or U17098 (N_17098,N_14066,N_15416);
xor U17099 (N_17099,N_14332,N_15388);
and U17100 (N_17100,N_15614,N_14231);
and U17101 (N_17101,N_15825,N_14336);
nor U17102 (N_17102,N_14347,N_15476);
or U17103 (N_17103,N_15081,N_14286);
nor U17104 (N_17104,N_15952,N_15168);
nor U17105 (N_17105,N_15829,N_15482);
nor U17106 (N_17106,N_14018,N_15117);
nor U17107 (N_17107,N_15213,N_14305);
nand U17108 (N_17108,N_15612,N_14525);
or U17109 (N_17109,N_15654,N_14992);
and U17110 (N_17110,N_14686,N_15789);
or U17111 (N_17111,N_14743,N_14486);
and U17112 (N_17112,N_15596,N_15573);
nor U17113 (N_17113,N_14912,N_14060);
nand U17114 (N_17114,N_14853,N_14285);
or U17115 (N_17115,N_15346,N_14123);
nand U17116 (N_17116,N_14168,N_15094);
or U17117 (N_17117,N_15869,N_14788);
or U17118 (N_17118,N_14364,N_14233);
nor U17119 (N_17119,N_15422,N_14186);
xnor U17120 (N_17120,N_15403,N_15101);
or U17121 (N_17121,N_15863,N_15338);
nand U17122 (N_17122,N_14788,N_14177);
nor U17123 (N_17123,N_14554,N_15771);
nand U17124 (N_17124,N_15070,N_14455);
and U17125 (N_17125,N_14307,N_15245);
xnor U17126 (N_17126,N_15943,N_15530);
nor U17127 (N_17127,N_15269,N_14347);
xnor U17128 (N_17128,N_14312,N_15876);
or U17129 (N_17129,N_15510,N_14000);
and U17130 (N_17130,N_14220,N_14783);
and U17131 (N_17131,N_14547,N_15688);
or U17132 (N_17132,N_15343,N_15432);
nor U17133 (N_17133,N_15742,N_15755);
nand U17134 (N_17134,N_14724,N_15641);
and U17135 (N_17135,N_15283,N_15515);
and U17136 (N_17136,N_14167,N_15730);
nor U17137 (N_17137,N_14162,N_15167);
xnor U17138 (N_17138,N_15192,N_14571);
nand U17139 (N_17139,N_15022,N_15932);
nor U17140 (N_17140,N_14934,N_15048);
and U17141 (N_17141,N_14519,N_15310);
nor U17142 (N_17142,N_15029,N_15340);
nand U17143 (N_17143,N_14979,N_14749);
and U17144 (N_17144,N_15333,N_14766);
xor U17145 (N_17145,N_15368,N_15721);
nor U17146 (N_17146,N_14347,N_14278);
nor U17147 (N_17147,N_15633,N_14195);
xor U17148 (N_17148,N_15876,N_15955);
nor U17149 (N_17149,N_14426,N_14955);
xnor U17150 (N_17150,N_15711,N_14237);
nor U17151 (N_17151,N_14860,N_14454);
or U17152 (N_17152,N_15611,N_15149);
and U17153 (N_17153,N_14603,N_15031);
xor U17154 (N_17154,N_14028,N_15706);
and U17155 (N_17155,N_14213,N_15023);
and U17156 (N_17156,N_15358,N_14620);
nand U17157 (N_17157,N_15291,N_14262);
xor U17158 (N_17158,N_14467,N_14367);
and U17159 (N_17159,N_15604,N_15259);
nor U17160 (N_17160,N_15347,N_14669);
xnor U17161 (N_17161,N_15031,N_14750);
xnor U17162 (N_17162,N_15102,N_15467);
nor U17163 (N_17163,N_14856,N_15633);
or U17164 (N_17164,N_14706,N_15367);
nand U17165 (N_17165,N_15331,N_14932);
xnor U17166 (N_17166,N_14247,N_14658);
xor U17167 (N_17167,N_15263,N_15887);
nand U17168 (N_17168,N_14286,N_14161);
or U17169 (N_17169,N_14234,N_14173);
and U17170 (N_17170,N_15301,N_15926);
nor U17171 (N_17171,N_14259,N_15434);
nand U17172 (N_17172,N_15083,N_15611);
nand U17173 (N_17173,N_15596,N_15229);
xnor U17174 (N_17174,N_15752,N_14817);
xnor U17175 (N_17175,N_14171,N_15257);
or U17176 (N_17176,N_14142,N_14712);
or U17177 (N_17177,N_15235,N_15163);
nand U17178 (N_17178,N_15949,N_14712);
nor U17179 (N_17179,N_14099,N_15791);
xor U17180 (N_17180,N_14164,N_15478);
and U17181 (N_17181,N_14085,N_14000);
nand U17182 (N_17182,N_15296,N_14930);
or U17183 (N_17183,N_15432,N_15700);
or U17184 (N_17184,N_14654,N_15431);
or U17185 (N_17185,N_14122,N_14185);
nand U17186 (N_17186,N_14790,N_15022);
or U17187 (N_17187,N_15404,N_15054);
xnor U17188 (N_17188,N_14367,N_15545);
nor U17189 (N_17189,N_15830,N_15603);
nor U17190 (N_17190,N_14554,N_14407);
nand U17191 (N_17191,N_15186,N_15090);
xnor U17192 (N_17192,N_14022,N_15507);
or U17193 (N_17193,N_14276,N_15758);
xnor U17194 (N_17194,N_15516,N_15133);
xor U17195 (N_17195,N_15474,N_14322);
nor U17196 (N_17196,N_15838,N_15758);
nand U17197 (N_17197,N_14426,N_14899);
nand U17198 (N_17198,N_15454,N_14267);
or U17199 (N_17199,N_14318,N_14938);
nor U17200 (N_17200,N_15223,N_15125);
nor U17201 (N_17201,N_15159,N_14220);
nand U17202 (N_17202,N_15598,N_14351);
nand U17203 (N_17203,N_15924,N_15996);
xnor U17204 (N_17204,N_14720,N_14823);
or U17205 (N_17205,N_14531,N_15041);
and U17206 (N_17206,N_15130,N_15964);
xor U17207 (N_17207,N_14055,N_15404);
and U17208 (N_17208,N_15278,N_14657);
nor U17209 (N_17209,N_15403,N_14982);
xnor U17210 (N_17210,N_15857,N_15608);
or U17211 (N_17211,N_14887,N_15923);
xor U17212 (N_17212,N_14351,N_15416);
or U17213 (N_17213,N_15468,N_15560);
nand U17214 (N_17214,N_14099,N_14148);
or U17215 (N_17215,N_15072,N_14738);
xor U17216 (N_17216,N_15677,N_15295);
or U17217 (N_17217,N_15346,N_14682);
nand U17218 (N_17218,N_14001,N_14534);
or U17219 (N_17219,N_14892,N_14232);
xnor U17220 (N_17220,N_15088,N_14037);
nand U17221 (N_17221,N_14367,N_14949);
nor U17222 (N_17222,N_14285,N_14660);
xnor U17223 (N_17223,N_15759,N_15103);
nand U17224 (N_17224,N_14442,N_14242);
or U17225 (N_17225,N_14707,N_15302);
xor U17226 (N_17226,N_15793,N_14675);
or U17227 (N_17227,N_14743,N_15063);
xnor U17228 (N_17228,N_14163,N_15035);
and U17229 (N_17229,N_15475,N_14241);
xnor U17230 (N_17230,N_15552,N_14814);
xnor U17231 (N_17231,N_14280,N_15386);
xnor U17232 (N_17232,N_14653,N_14161);
xor U17233 (N_17233,N_15621,N_15070);
and U17234 (N_17234,N_15539,N_14853);
nor U17235 (N_17235,N_14531,N_14504);
nor U17236 (N_17236,N_15796,N_14265);
xnor U17237 (N_17237,N_15311,N_14419);
nand U17238 (N_17238,N_15933,N_14381);
nor U17239 (N_17239,N_14946,N_15470);
and U17240 (N_17240,N_14567,N_15011);
and U17241 (N_17241,N_15932,N_15909);
and U17242 (N_17242,N_14301,N_15348);
xnor U17243 (N_17243,N_15775,N_14055);
nand U17244 (N_17244,N_14839,N_14627);
xor U17245 (N_17245,N_14695,N_15283);
or U17246 (N_17246,N_15976,N_14752);
nand U17247 (N_17247,N_14280,N_15716);
and U17248 (N_17248,N_15836,N_14772);
and U17249 (N_17249,N_14125,N_14153);
xnor U17250 (N_17250,N_15293,N_15125);
or U17251 (N_17251,N_15196,N_14143);
and U17252 (N_17252,N_14886,N_14241);
xnor U17253 (N_17253,N_15888,N_14221);
and U17254 (N_17254,N_15235,N_14178);
or U17255 (N_17255,N_14713,N_15316);
or U17256 (N_17256,N_15521,N_14702);
nand U17257 (N_17257,N_15088,N_14791);
or U17258 (N_17258,N_14640,N_14671);
nand U17259 (N_17259,N_14932,N_14363);
or U17260 (N_17260,N_14879,N_14064);
and U17261 (N_17261,N_15267,N_14142);
xor U17262 (N_17262,N_15645,N_15927);
xor U17263 (N_17263,N_14542,N_14253);
nand U17264 (N_17264,N_14766,N_15514);
nor U17265 (N_17265,N_14199,N_15930);
nor U17266 (N_17266,N_14480,N_14632);
nand U17267 (N_17267,N_15291,N_15597);
nand U17268 (N_17268,N_14389,N_15294);
nand U17269 (N_17269,N_15248,N_15222);
or U17270 (N_17270,N_14648,N_14876);
nand U17271 (N_17271,N_15469,N_15040);
xor U17272 (N_17272,N_14103,N_14892);
nand U17273 (N_17273,N_15278,N_14596);
and U17274 (N_17274,N_15334,N_14837);
nor U17275 (N_17275,N_15387,N_15128);
or U17276 (N_17276,N_14818,N_15956);
and U17277 (N_17277,N_15771,N_15280);
and U17278 (N_17278,N_14926,N_14660);
nor U17279 (N_17279,N_14919,N_15625);
xor U17280 (N_17280,N_15514,N_15149);
or U17281 (N_17281,N_14984,N_15529);
nand U17282 (N_17282,N_15812,N_15017);
nand U17283 (N_17283,N_14944,N_14524);
xor U17284 (N_17284,N_15883,N_15562);
xnor U17285 (N_17285,N_15892,N_15551);
nor U17286 (N_17286,N_15557,N_15078);
nor U17287 (N_17287,N_15255,N_15584);
nor U17288 (N_17288,N_15355,N_15661);
nand U17289 (N_17289,N_15748,N_15764);
nand U17290 (N_17290,N_14574,N_14783);
nor U17291 (N_17291,N_15587,N_14376);
or U17292 (N_17292,N_15493,N_15989);
and U17293 (N_17293,N_15521,N_15226);
and U17294 (N_17294,N_15755,N_15208);
nor U17295 (N_17295,N_14178,N_15859);
nand U17296 (N_17296,N_15591,N_14672);
and U17297 (N_17297,N_15835,N_15403);
or U17298 (N_17298,N_14599,N_15465);
nor U17299 (N_17299,N_15525,N_15539);
nand U17300 (N_17300,N_15262,N_14728);
or U17301 (N_17301,N_15134,N_14624);
nor U17302 (N_17302,N_15543,N_14052);
nor U17303 (N_17303,N_14793,N_14414);
nor U17304 (N_17304,N_14071,N_14096);
and U17305 (N_17305,N_14030,N_15567);
or U17306 (N_17306,N_14069,N_15711);
and U17307 (N_17307,N_14604,N_15195);
xor U17308 (N_17308,N_15878,N_15856);
nor U17309 (N_17309,N_14583,N_15085);
xor U17310 (N_17310,N_15395,N_15941);
nand U17311 (N_17311,N_15277,N_14776);
and U17312 (N_17312,N_15925,N_15152);
or U17313 (N_17313,N_15162,N_15930);
xnor U17314 (N_17314,N_14569,N_15937);
nand U17315 (N_17315,N_14436,N_15835);
or U17316 (N_17316,N_15685,N_14589);
xor U17317 (N_17317,N_15540,N_14451);
nand U17318 (N_17318,N_15868,N_15896);
xor U17319 (N_17319,N_14455,N_14188);
nand U17320 (N_17320,N_15397,N_15549);
and U17321 (N_17321,N_14408,N_15352);
nand U17322 (N_17322,N_14882,N_15559);
or U17323 (N_17323,N_15396,N_14687);
nor U17324 (N_17324,N_14884,N_15056);
xnor U17325 (N_17325,N_15626,N_14019);
nor U17326 (N_17326,N_14296,N_14630);
nand U17327 (N_17327,N_14669,N_15186);
nor U17328 (N_17328,N_15414,N_14342);
xnor U17329 (N_17329,N_14864,N_14619);
and U17330 (N_17330,N_14256,N_14900);
nand U17331 (N_17331,N_14967,N_14181);
or U17332 (N_17332,N_15774,N_14439);
nor U17333 (N_17333,N_15673,N_14670);
nor U17334 (N_17334,N_14685,N_15078);
or U17335 (N_17335,N_15650,N_14523);
nand U17336 (N_17336,N_14962,N_14653);
nor U17337 (N_17337,N_14737,N_14771);
and U17338 (N_17338,N_15251,N_15700);
xor U17339 (N_17339,N_15440,N_14914);
xor U17340 (N_17340,N_14993,N_14173);
or U17341 (N_17341,N_14499,N_14039);
xor U17342 (N_17342,N_14324,N_15648);
nand U17343 (N_17343,N_15863,N_14806);
or U17344 (N_17344,N_14286,N_15916);
or U17345 (N_17345,N_14297,N_15170);
nor U17346 (N_17346,N_14555,N_14926);
xor U17347 (N_17347,N_15591,N_15667);
xnor U17348 (N_17348,N_14319,N_15343);
nand U17349 (N_17349,N_15537,N_14837);
and U17350 (N_17350,N_14341,N_15568);
nor U17351 (N_17351,N_14527,N_15534);
and U17352 (N_17352,N_15617,N_14677);
and U17353 (N_17353,N_14736,N_14247);
or U17354 (N_17354,N_14250,N_14533);
xor U17355 (N_17355,N_15250,N_14622);
nor U17356 (N_17356,N_15040,N_14929);
or U17357 (N_17357,N_15013,N_15959);
nor U17358 (N_17358,N_15101,N_14316);
xnor U17359 (N_17359,N_15704,N_15071);
or U17360 (N_17360,N_14408,N_14421);
or U17361 (N_17361,N_14169,N_15016);
xnor U17362 (N_17362,N_14569,N_15558);
nor U17363 (N_17363,N_14663,N_15499);
nand U17364 (N_17364,N_15926,N_15047);
nand U17365 (N_17365,N_14339,N_15679);
xor U17366 (N_17366,N_14740,N_14540);
or U17367 (N_17367,N_14861,N_15489);
xor U17368 (N_17368,N_14319,N_15252);
nand U17369 (N_17369,N_15089,N_14035);
nand U17370 (N_17370,N_15990,N_15019);
nor U17371 (N_17371,N_14911,N_14015);
and U17372 (N_17372,N_15326,N_14934);
and U17373 (N_17373,N_14694,N_14664);
xnor U17374 (N_17374,N_15829,N_15624);
nor U17375 (N_17375,N_15307,N_14696);
nand U17376 (N_17376,N_15442,N_14863);
or U17377 (N_17377,N_15406,N_15530);
nand U17378 (N_17378,N_15267,N_15605);
xor U17379 (N_17379,N_14352,N_14024);
and U17380 (N_17380,N_14582,N_15800);
nor U17381 (N_17381,N_15653,N_14193);
xnor U17382 (N_17382,N_14114,N_15216);
nand U17383 (N_17383,N_15978,N_15009);
and U17384 (N_17384,N_15967,N_14039);
xnor U17385 (N_17385,N_14803,N_15963);
or U17386 (N_17386,N_15189,N_15661);
and U17387 (N_17387,N_14014,N_14363);
or U17388 (N_17388,N_14312,N_14202);
xnor U17389 (N_17389,N_15345,N_14504);
and U17390 (N_17390,N_15929,N_15487);
and U17391 (N_17391,N_15671,N_15819);
and U17392 (N_17392,N_14637,N_15483);
or U17393 (N_17393,N_15043,N_14335);
nor U17394 (N_17394,N_15741,N_15078);
or U17395 (N_17395,N_15565,N_14751);
nand U17396 (N_17396,N_14078,N_14188);
or U17397 (N_17397,N_15540,N_15283);
nand U17398 (N_17398,N_15889,N_14074);
nor U17399 (N_17399,N_14733,N_14825);
nor U17400 (N_17400,N_15918,N_15304);
nand U17401 (N_17401,N_14827,N_15429);
nand U17402 (N_17402,N_14174,N_14353);
or U17403 (N_17403,N_15136,N_15207);
nor U17404 (N_17404,N_15705,N_15132);
and U17405 (N_17405,N_14215,N_14546);
nor U17406 (N_17406,N_14316,N_15707);
nand U17407 (N_17407,N_14897,N_15392);
or U17408 (N_17408,N_14065,N_14417);
nand U17409 (N_17409,N_15986,N_15040);
xor U17410 (N_17410,N_15272,N_14973);
or U17411 (N_17411,N_15493,N_15969);
or U17412 (N_17412,N_15686,N_14081);
or U17413 (N_17413,N_15899,N_14446);
xnor U17414 (N_17414,N_14699,N_14692);
or U17415 (N_17415,N_15291,N_14817);
and U17416 (N_17416,N_14197,N_15653);
nand U17417 (N_17417,N_15549,N_15303);
and U17418 (N_17418,N_15731,N_14125);
nor U17419 (N_17419,N_15353,N_14108);
nand U17420 (N_17420,N_14472,N_15444);
and U17421 (N_17421,N_15680,N_15046);
nand U17422 (N_17422,N_14946,N_15700);
or U17423 (N_17423,N_15663,N_14249);
xor U17424 (N_17424,N_14174,N_15887);
nand U17425 (N_17425,N_15727,N_15493);
nand U17426 (N_17426,N_14305,N_14436);
nor U17427 (N_17427,N_15118,N_15652);
or U17428 (N_17428,N_15448,N_15051);
or U17429 (N_17429,N_15655,N_14003);
xnor U17430 (N_17430,N_14115,N_14255);
nand U17431 (N_17431,N_15342,N_14191);
nand U17432 (N_17432,N_15216,N_14255);
nor U17433 (N_17433,N_14134,N_14068);
or U17434 (N_17434,N_15857,N_15624);
nand U17435 (N_17435,N_15008,N_14271);
nand U17436 (N_17436,N_15888,N_14252);
nand U17437 (N_17437,N_14881,N_14026);
xnor U17438 (N_17438,N_15140,N_14223);
and U17439 (N_17439,N_14598,N_15937);
xnor U17440 (N_17440,N_14710,N_14355);
and U17441 (N_17441,N_15950,N_15510);
and U17442 (N_17442,N_14148,N_14284);
nand U17443 (N_17443,N_14757,N_15783);
nor U17444 (N_17444,N_15510,N_15827);
nand U17445 (N_17445,N_14527,N_15389);
xor U17446 (N_17446,N_15075,N_15158);
or U17447 (N_17447,N_15856,N_15711);
and U17448 (N_17448,N_14949,N_15909);
xor U17449 (N_17449,N_15133,N_14649);
or U17450 (N_17450,N_15264,N_14967);
and U17451 (N_17451,N_15995,N_15996);
xnor U17452 (N_17452,N_14411,N_14157);
nor U17453 (N_17453,N_14409,N_15698);
nor U17454 (N_17454,N_15075,N_15862);
or U17455 (N_17455,N_14293,N_15277);
nor U17456 (N_17456,N_14691,N_14926);
nand U17457 (N_17457,N_15739,N_14390);
or U17458 (N_17458,N_14602,N_14493);
xor U17459 (N_17459,N_15770,N_14547);
xnor U17460 (N_17460,N_15749,N_14703);
nor U17461 (N_17461,N_15999,N_14544);
nand U17462 (N_17462,N_15481,N_15936);
and U17463 (N_17463,N_15835,N_15326);
or U17464 (N_17464,N_14268,N_15719);
nand U17465 (N_17465,N_14688,N_14810);
nor U17466 (N_17466,N_14694,N_15578);
xor U17467 (N_17467,N_15971,N_14104);
nor U17468 (N_17468,N_14142,N_15106);
and U17469 (N_17469,N_14993,N_14470);
and U17470 (N_17470,N_15159,N_14724);
nand U17471 (N_17471,N_15158,N_14013);
nor U17472 (N_17472,N_14073,N_14309);
xor U17473 (N_17473,N_15219,N_14967);
and U17474 (N_17474,N_15758,N_14618);
or U17475 (N_17475,N_14418,N_15883);
xnor U17476 (N_17476,N_15287,N_14921);
xor U17477 (N_17477,N_14030,N_14458);
xnor U17478 (N_17478,N_14719,N_14178);
nand U17479 (N_17479,N_15912,N_15844);
or U17480 (N_17480,N_15931,N_15806);
or U17481 (N_17481,N_15525,N_15269);
nand U17482 (N_17482,N_15025,N_14976);
nor U17483 (N_17483,N_15140,N_14749);
and U17484 (N_17484,N_14139,N_14506);
or U17485 (N_17485,N_14965,N_15584);
nand U17486 (N_17486,N_15281,N_15792);
xor U17487 (N_17487,N_15061,N_15179);
nor U17488 (N_17488,N_14904,N_15636);
or U17489 (N_17489,N_15050,N_14767);
nor U17490 (N_17490,N_14118,N_14822);
xnor U17491 (N_17491,N_14521,N_15502);
xnor U17492 (N_17492,N_14749,N_14568);
or U17493 (N_17493,N_15813,N_14300);
xor U17494 (N_17494,N_14372,N_15289);
xor U17495 (N_17495,N_15588,N_14890);
and U17496 (N_17496,N_15555,N_15818);
xor U17497 (N_17497,N_15797,N_15940);
xor U17498 (N_17498,N_15078,N_15885);
xor U17499 (N_17499,N_14005,N_14562);
and U17500 (N_17500,N_14307,N_14729);
nand U17501 (N_17501,N_15886,N_14758);
xor U17502 (N_17502,N_14596,N_15126);
or U17503 (N_17503,N_14407,N_15981);
nand U17504 (N_17504,N_14705,N_14796);
or U17505 (N_17505,N_15667,N_15048);
xnor U17506 (N_17506,N_14536,N_14537);
nor U17507 (N_17507,N_14142,N_15841);
nor U17508 (N_17508,N_14642,N_15795);
nor U17509 (N_17509,N_15425,N_15909);
nor U17510 (N_17510,N_15618,N_15430);
xor U17511 (N_17511,N_15085,N_14331);
and U17512 (N_17512,N_14031,N_15916);
xor U17513 (N_17513,N_14236,N_14985);
xnor U17514 (N_17514,N_15382,N_15225);
and U17515 (N_17515,N_15350,N_15561);
nand U17516 (N_17516,N_15474,N_14897);
and U17517 (N_17517,N_14556,N_14053);
nand U17518 (N_17518,N_15400,N_15865);
and U17519 (N_17519,N_14769,N_14745);
nand U17520 (N_17520,N_15801,N_14913);
nor U17521 (N_17521,N_15375,N_15252);
nand U17522 (N_17522,N_14640,N_14677);
and U17523 (N_17523,N_15187,N_15106);
nand U17524 (N_17524,N_15911,N_14446);
nand U17525 (N_17525,N_15374,N_15090);
and U17526 (N_17526,N_15035,N_14284);
nand U17527 (N_17527,N_15834,N_15431);
or U17528 (N_17528,N_15916,N_15135);
or U17529 (N_17529,N_14615,N_14280);
nor U17530 (N_17530,N_14744,N_14479);
or U17531 (N_17531,N_14162,N_14935);
xnor U17532 (N_17532,N_15046,N_15056);
or U17533 (N_17533,N_14967,N_14909);
or U17534 (N_17534,N_14861,N_15807);
or U17535 (N_17535,N_14406,N_14926);
and U17536 (N_17536,N_14559,N_15550);
or U17537 (N_17537,N_15195,N_14152);
xor U17538 (N_17538,N_14870,N_14635);
xor U17539 (N_17539,N_14294,N_15087);
and U17540 (N_17540,N_15981,N_14436);
and U17541 (N_17541,N_15021,N_14062);
and U17542 (N_17542,N_15766,N_15744);
and U17543 (N_17543,N_14949,N_15357);
or U17544 (N_17544,N_14731,N_15378);
nor U17545 (N_17545,N_14039,N_14749);
xnor U17546 (N_17546,N_14291,N_14336);
nor U17547 (N_17547,N_14205,N_15883);
and U17548 (N_17548,N_14481,N_15717);
nor U17549 (N_17549,N_14507,N_15850);
or U17550 (N_17550,N_15640,N_14590);
or U17551 (N_17551,N_15675,N_15945);
nand U17552 (N_17552,N_15617,N_15050);
nor U17553 (N_17553,N_15403,N_15790);
and U17554 (N_17554,N_15549,N_15527);
and U17555 (N_17555,N_15350,N_15332);
and U17556 (N_17556,N_15557,N_15296);
xnor U17557 (N_17557,N_14563,N_14288);
or U17558 (N_17558,N_15266,N_14811);
or U17559 (N_17559,N_14695,N_15728);
xnor U17560 (N_17560,N_14198,N_15823);
xnor U17561 (N_17561,N_14347,N_14280);
or U17562 (N_17562,N_14014,N_14524);
nand U17563 (N_17563,N_14555,N_14474);
and U17564 (N_17564,N_14890,N_15434);
or U17565 (N_17565,N_15103,N_15216);
or U17566 (N_17566,N_15634,N_15614);
nor U17567 (N_17567,N_15719,N_14998);
nand U17568 (N_17568,N_14719,N_15550);
and U17569 (N_17569,N_15644,N_14051);
nor U17570 (N_17570,N_14565,N_15944);
xnor U17571 (N_17571,N_15871,N_14770);
nand U17572 (N_17572,N_15349,N_15751);
xnor U17573 (N_17573,N_14061,N_14354);
xor U17574 (N_17574,N_15941,N_15672);
nor U17575 (N_17575,N_14262,N_14925);
xnor U17576 (N_17576,N_15444,N_15819);
and U17577 (N_17577,N_14069,N_14658);
nand U17578 (N_17578,N_15906,N_14905);
or U17579 (N_17579,N_15952,N_15506);
nor U17580 (N_17580,N_15868,N_14296);
xor U17581 (N_17581,N_14774,N_14624);
nor U17582 (N_17582,N_15253,N_14318);
nand U17583 (N_17583,N_15798,N_14282);
nor U17584 (N_17584,N_14531,N_15520);
nand U17585 (N_17585,N_14867,N_14710);
or U17586 (N_17586,N_15773,N_14160);
and U17587 (N_17587,N_15119,N_14138);
nor U17588 (N_17588,N_15519,N_15470);
xnor U17589 (N_17589,N_15048,N_14622);
or U17590 (N_17590,N_15048,N_14703);
xnor U17591 (N_17591,N_15833,N_14417);
and U17592 (N_17592,N_14260,N_15367);
xnor U17593 (N_17593,N_15751,N_15608);
nor U17594 (N_17594,N_14445,N_14717);
and U17595 (N_17595,N_15691,N_15432);
and U17596 (N_17596,N_14994,N_15124);
or U17597 (N_17597,N_14912,N_15843);
and U17598 (N_17598,N_15454,N_15704);
xnor U17599 (N_17599,N_15773,N_14301);
xnor U17600 (N_17600,N_14416,N_14091);
and U17601 (N_17601,N_14218,N_15975);
nor U17602 (N_17602,N_15741,N_14782);
nor U17603 (N_17603,N_14933,N_14013);
xor U17604 (N_17604,N_14415,N_14640);
nor U17605 (N_17605,N_15520,N_15117);
nor U17606 (N_17606,N_14262,N_14003);
xnor U17607 (N_17607,N_15369,N_14696);
xnor U17608 (N_17608,N_15262,N_15087);
or U17609 (N_17609,N_14458,N_14313);
xor U17610 (N_17610,N_15722,N_14413);
and U17611 (N_17611,N_14530,N_14235);
nor U17612 (N_17612,N_14049,N_15355);
xnor U17613 (N_17613,N_14124,N_14147);
or U17614 (N_17614,N_15355,N_14961);
nor U17615 (N_17615,N_15510,N_14460);
nand U17616 (N_17616,N_15856,N_15824);
or U17617 (N_17617,N_15820,N_15576);
nor U17618 (N_17618,N_14495,N_15150);
xnor U17619 (N_17619,N_15858,N_15206);
xor U17620 (N_17620,N_15765,N_15475);
nand U17621 (N_17621,N_15715,N_15191);
or U17622 (N_17622,N_14658,N_14892);
nor U17623 (N_17623,N_14552,N_15710);
or U17624 (N_17624,N_15333,N_15427);
nor U17625 (N_17625,N_14445,N_14273);
nor U17626 (N_17626,N_15381,N_15434);
and U17627 (N_17627,N_15840,N_14416);
and U17628 (N_17628,N_15044,N_14978);
or U17629 (N_17629,N_14177,N_15248);
or U17630 (N_17630,N_15432,N_15087);
nor U17631 (N_17631,N_15021,N_15184);
xor U17632 (N_17632,N_14429,N_14590);
nor U17633 (N_17633,N_14621,N_14780);
and U17634 (N_17634,N_15276,N_14811);
xnor U17635 (N_17635,N_14028,N_15453);
or U17636 (N_17636,N_15443,N_15710);
or U17637 (N_17637,N_15277,N_14927);
and U17638 (N_17638,N_14162,N_15722);
and U17639 (N_17639,N_14209,N_15079);
xnor U17640 (N_17640,N_14251,N_15932);
xnor U17641 (N_17641,N_15570,N_14088);
xnor U17642 (N_17642,N_15396,N_14115);
or U17643 (N_17643,N_15707,N_14676);
or U17644 (N_17644,N_14375,N_15013);
nor U17645 (N_17645,N_14148,N_14429);
and U17646 (N_17646,N_15480,N_14083);
or U17647 (N_17647,N_15846,N_14547);
nor U17648 (N_17648,N_15413,N_14620);
xor U17649 (N_17649,N_15546,N_14561);
and U17650 (N_17650,N_14755,N_15014);
and U17651 (N_17651,N_14693,N_15856);
nor U17652 (N_17652,N_15331,N_14051);
xor U17653 (N_17653,N_14153,N_14139);
or U17654 (N_17654,N_14247,N_14364);
nand U17655 (N_17655,N_14885,N_15455);
xor U17656 (N_17656,N_15634,N_15494);
xnor U17657 (N_17657,N_15238,N_14407);
or U17658 (N_17658,N_15579,N_14968);
nor U17659 (N_17659,N_14548,N_14013);
nand U17660 (N_17660,N_14420,N_15830);
or U17661 (N_17661,N_15631,N_15986);
nor U17662 (N_17662,N_15838,N_14654);
xor U17663 (N_17663,N_14801,N_14346);
nand U17664 (N_17664,N_15592,N_15233);
and U17665 (N_17665,N_14210,N_14450);
or U17666 (N_17666,N_15125,N_15839);
xnor U17667 (N_17667,N_14465,N_15295);
or U17668 (N_17668,N_14855,N_15900);
nand U17669 (N_17669,N_15191,N_15308);
xnor U17670 (N_17670,N_15416,N_15423);
nand U17671 (N_17671,N_15739,N_15305);
or U17672 (N_17672,N_14954,N_15751);
xor U17673 (N_17673,N_14678,N_14878);
and U17674 (N_17674,N_15456,N_15113);
nand U17675 (N_17675,N_14011,N_15482);
nand U17676 (N_17676,N_15479,N_15085);
or U17677 (N_17677,N_14802,N_15869);
xor U17678 (N_17678,N_15676,N_15236);
xnor U17679 (N_17679,N_14326,N_15252);
and U17680 (N_17680,N_15581,N_15872);
xor U17681 (N_17681,N_14456,N_15884);
xnor U17682 (N_17682,N_14579,N_14831);
or U17683 (N_17683,N_15000,N_15445);
nand U17684 (N_17684,N_15165,N_14720);
nor U17685 (N_17685,N_14934,N_15696);
nor U17686 (N_17686,N_14412,N_14799);
or U17687 (N_17687,N_14890,N_14340);
and U17688 (N_17688,N_15608,N_15118);
xor U17689 (N_17689,N_15496,N_14403);
nor U17690 (N_17690,N_14222,N_14090);
or U17691 (N_17691,N_14300,N_15161);
nand U17692 (N_17692,N_15393,N_14573);
or U17693 (N_17693,N_15951,N_15330);
xnor U17694 (N_17694,N_15678,N_15371);
or U17695 (N_17695,N_15043,N_14513);
xor U17696 (N_17696,N_15564,N_15885);
nand U17697 (N_17697,N_14055,N_15584);
nand U17698 (N_17698,N_15298,N_14756);
xor U17699 (N_17699,N_15573,N_14251);
or U17700 (N_17700,N_15242,N_15518);
or U17701 (N_17701,N_14358,N_15168);
nor U17702 (N_17702,N_15179,N_14896);
xnor U17703 (N_17703,N_14195,N_14962);
or U17704 (N_17704,N_14713,N_15115);
or U17705 (N_17705,N_15094,N_15840);
and U17706 (N_17706,N_14344,N_14110);
xor U17707 (N_17707,N_14142,N_15397);
nor U17708 (N_17708,N_15364,N_14473);
xnor U17709 (N_17709,N_14092,N_15341);
or U17710 (N_17710,N_14498,N_14428);
nand U17711 (N_17711,N_15615,N_15191);
nand U17712 (N_17712,N_14335,N_14778);
or U17713 (N_17713,N_14878,N_15660);
nand U17714 (N_17714,N_15657,N_15283);
and U17715 (N_17715,N_14826,N_15228);
xor U17716 (N_17716,N_15403,N_15713);
or U17717 (N_17717,N_14168,N_14601);
or U17718 (N_17718,N_14575,N_15045);
nand U17719 (N_17719,N_14775,N_15704);
and U17720 (N_17720,N_15614,N_14688);
and U17721 (N_17721,N_15080,N_15961);
nand U17722 (N_17722,N_14948,N_14520);
xnor U17723 (N_17723,N_14684,N_14734);
nor U17724 (N_17724,N_15681,N_15677);
nor U17725 (N_17725,N_15575,N_14852);
nor U17726 (N_17726,N_14769,N_15015);
and U17727 (N_17727,N_14676,N_15486);
nand U17728 (N_17728,N_15254,N_15964);
nor U17729 (N_17729,N_15905,N_15079);
or U17730 (N_17730,N_14133,N_15882);
or U17731 (N_17731,N_14322,N_14746);
xnor U17732 (N_17732,N_15149,N_15805);
xor U17733 (N_17733,N_15077,N_15317);
nor U17734 (N_17734,N_14375,N_14992);
nor U17735 (N_17735,N_15113,N_15405);
xnor U17736 (N_17736,N_15464,N_14790);
and U17737 (N_17737,N_15461,N_15255);
nand U17738 (N_17738,N_14103,N_15591);
and U17739 (N_17739,N_14666,N_15250);
nor U17740 (N_17740,N_15200,N_15589);
xnor U17741 (N_17741,N_15034,N_15382);
nor U17742 (N_17742,N_14101,N_15309);
nor U17743 (N_17743,N_14166,N_14200);
or U17744 (N_17744,N_15387,N_15322);
or U17745 (N_17745,N_14347,N_14437);
and U17746 (N_17746,N_14220,N_14762);
nor U17747 (N_17747,N_14867,N_14834);
or U17748 (N_17748,N_14979,N_15262);
xnor U17749 (N_17749,N_14396,N_14809);
xnor U17750 (N_17750,N_15720,N_14189);
nand U17751 (N_17751,N_14654,N_15084);
and U17752 (N_17752,N_15643,N_14787);
and U17753 (N_17753,N_14435,N_14923);
nand U17754 (N_17754,N_14831,N_14503);
xor U17755 (N_17755,N_15859,N_15783);
and U17756 (N_17756,N_14995,N_14760);
xnor U17757 (N_17757,N_15050,N_15687);
nor U17758 (N_17758,N_15569,N_14865);
and U17759 (N_17759,N_15970,N_14596);
xor U17760 (N_17760,N_15605,N_14879);
and U17761 (N_17761,N_14064,N_15476);
nand U17762 (N_17762,N_15032,N_14820);
and U17763 (N_17763,N_14113,N_14356);
xor U17764 (N_17764,N_15045,N_14094);
and U17765 (N_17765,N_15600,N_14091);
or U17766 (N_17766,N_15183,N_15466);
xnor U17767 (N_17767,N_15764,N_14890);
or U17768 (N_17768,N_15696,N_15298);
or U17769 (N_17769,N_14708,N_15337);
and U17770 (N_17770,N_15175,N_14595);
nand U17771 (N_17771,N_14498,N_15667);
nor U17772 (N_17772,N_14935,N_14459);
or U17773 (N_17773,N_14370,N_15996);
nor U17774 (N_17774,N_14341,N_14191);
or U17775 (N_17775,N_14589,N_14991);
nand U17776 (N_17776,N_15744,N_15751);
and U17777 (N_17777,N_15513,N_15216);
nor U17778 (N_17778,N_15207,N_14603);
and U17779 (N_17779,N_14725,N_14330);
xnor U17780 (N_17780,N_14681,N_14669);
and U17781 (N_17781,N_14284,N_15033);
and U17782 (N_17782,N_15760,N_15984);
nand U17783 (N_17783,N_15195,N_15938);
nand U17784 (N_17784,N_15107,N_14616);
and U17785 (N_17785,N_14165,N_14071);
and U17786 (N_17786,N_14882,N_14152);
and U17787 (N_17787,N_14003,N_14596);
or U17788 (N_17788,N_14691,N_14935);
or U17789 (N_17789,N_14129,N_14018);
nor U17790 (N_17790,N_15626,N_15989);
nand U17791 (N_17791,N_14944,N_14174);
xnor U17792 (N_17792,N_15972,N_15540);
nand U17793 (N_17793,N_14139,N_15339);
or U17794 (N_17794,N_15412,N_15230);
nand U17795 (N_17795,N_15939,N_14093);
xnor U17796 (N_17796,N_14352,N_15992);
nor U17797 (N_17797,N_14107,N_14461);
or U17798 (N_17798,N_15966,N_14873);
nor U17799 (N_17799,N_15021,N_15473);
nand U17800 (N_17800,N_15538,N_14513);
and U17801 (N_17801,N_14457,N_14704);
nor U17802 (N_17802,N_15201,N_14538);
nor U17803 (N_17803,N_15972,N_15403);
or U17804 (N_17804,N_15622,N_14582);
and U17805 (N_17805,N_15617,N_14089);
nand U17806 (N_17806,N_15746,N_14295);
xor U17807 (N_17807,N_15135,N_15074);
and U17808 (N_17808,N_15715,N_14763);
nor U17809 (N_17809,N_15865,N_14645);
nor U17810 (N_17810,N_14990,N_14547);
nand U17811 (N_17811,N_15706,N_15172);
nand U17812 (N_17812,N_15549,N_15888);
or U17813 (N_17813,N_14351,N_14930);
xor U17814 (N_17814,N_14031,N_14235);
nand U17815 (N_17815,N_15499,N_15081);
xnor U17816 (N_17816,N_15735,N_15633);
and U17817 (N_17817,N_15306,N_14949);
xor U17818 (N_17818,N_15122,N_15833);
xor U17819 (N_17819,N_14601,N_15118);
nand U17820 (N_17820,N_14469,N_14976);
and U17821 (N_17821,N_14083,N_14646);
or U17822 (N_17822,N_15282,N_14837);
and U17823 (N_17823,N_15972,N_15877);
nor U17824 (N_17824,N_15786,N_15160);
nor U17825 (N_17825,N_14002,N_15781);
nand U17826 (N_17826,N_15453,N_14022);
nor U17827 (N_17827,N_14003,N_15168);
nand U17828 (N_17828,N_14842,N_14551);
nand U17829 (N_17829,N_15794,N_14328);
nor U17830 (N_17830,N_14462,N_15624);
or U17831 (N_17831,N_15517,N_15332);
nor U17832 (N_17832,N_15314,N_14309);
nand U17833 (N_17833,N_15508,N_15771);
xnor U17834 (N_17834,N_14354,N_15759);
or U17835 (N_17835,N_15189,N_14714);
nand U17836 (N_17836,N_14822,N_14012);
nor U17837 (N_17837,N_14269,N_14122);
and U17838 (N_17838,N_14348,N_14453);
nand U17839 (N_17839,N_15294,N_14650);
nor U17840 (N_17840,N_15296,N_14407);
and U17841 (N_17841,N_14278,N_15778);
nand U17842 (N_17842,N_14051,N_15321);
xor U17843 (N_17843,N_15840,N_15223);
nand U17844 (N_17844,N_15132,N_14240);
nor U17845 (N_17845,N_14789,N_15852);
or U17846 (N_17846,N_15467,N_15902);
or U17847 (N_17847,N_14574,N_14355);
or U17848 (N_17848,N_14606,N_15155);
or U17849 (N_17849,N_15958,N_15179);
and U17850 (N_17850,N_14708,N_15390);
or U17851 (N_17851,N_14671,N_15340);
or U17852 (N_17852,N_15662,N_14830);
xor U17853 (N_17853,N_14437,N_15381);
and U17854 (N_17854,N_14854,N_15229);
nand U17855 (N_17855,N_14235,N_15786);
xor U17856 (N_17856,N_15792,N_15120);
and U17857 (N_17857,N_14286,N_14572);
xor U17858 (N_17858,N_14231,N_14828);
xor U17859 (N_17859,N_14540,N_15452);
and U17860 (N_17860,N_14716,N_15989);
or U17861 (N_17861,N_14684,N_15778);
nor U17862 (N_17862,N_14911,N_15090);
nand U17863 (N_17863,N_14816,N_14083);
xor U17864 (N_17864,N_14102,N_14178);
xnor U17865 (N_17865,N_14783,N_14116);
xnor U17866 (N_17866,N_14207,N_14778);
or U17867 (N_17867,N_15462,N_15414);
nor U17868 (N_17868,N_14895,N_14101);
nor U17869 (N_17869,N_14166,N_14094);
nor U17870 (N_17870,N_14739,N_15427);
nand U17871 (N_17871,N_15317,N_15126);
nor U17872 (N_17872,N_15650,N_15981);
and U17873 (N_17873,N_15512,N_14132);
or U17874 (N_17874,N_15564,N_14429);
or U17875 (N_17875,N_14755,N_15174);
xor U17876 (N_17876,N_15669,N_14924);
xnor U17877 (N_17877,N_14893,N_14535);
nor U17878 (N_17878,N_14626,N_14316);
nand U17879 (N_17879,N_14731,N_15778);
or U17880 (N_17880,N_15166,N_14864);
nor U17881 (N_17881,N_15381,N_15683);
nand U17882 (N_17882,N_15162,N_14521);
nor U17883 (N_17883,N_14579,N_15151);
or U17884 (N_17884,N_14633,N_14753);
or U17885 (N_17885,N_15746,N_14012);
xnor U17886 (N_17886,N_15991,N_15530);
nand U17887 (N_17887,N_14807,N_14290);
xnor U17888 (N_17888,N_15794,N_15559);
or U17889 (N_17889,N_15746,N_14616);
xor U17890 (N_17890,N_14691,N_15887);
or U17891 (N_17891,N_15063,N_15242);
nand U17892 (N_17892,N_15049,N_15597);
or U17893 (N_17893,N_14681,N_15219);
nand U17894 (N_17894,N_14101,N_15660);
or U17895 (N_17895,N_14423,N_15928);
xnor U17896 (N_17896,N_14216,N_14037);
nor U17897 (N_17897,N_14110,N_14175);
or U17898 (N_17898,N_14970,N_15804);
and U17899 (N_17899,N_15147,N_14361);
nand U17900 (N_17900,N_15698,N_14607);
or U17901 (N_17901,N_14201,N_15149);
nand U17902 (N_17902,N_14775,N_14056);
or U17903 (N_17903,N_14358,N_14521);
or U17904 (N_17904,N_15546,N_14609);
nand U17905 (N_17905,N_14339,N_14887);
or U17906 (N_17906,N_15946,N_15690);
and U17907 (N_17907,N_15608,N_14885);
nor U17908 (N_17908,N_15834,N_15173);
nor U17909 (N_17909,N_15503,N_14193);
nor U17910 (N_17910,N_14754,N_14001);
or U17911 (N_17911,N_15569,N_15491);
nor U17912 (N_17912,N_14931,N_14968);
nand U17913 (N_17913,N_15195,N_15946);
nand U17914 (N_17914,N_14517,N_15262);
nand U17915 (N_17915,N_15191,N_14010);
nand U17916 (N_17916,N_15433,N_15127);
or U17917 (N_17917,N_14542,N_14302);
nor U17918 (N_17918,N_14118,N_15308);
and U17919 (N_17919,N_14732,N_15893);
nor U17920 (N_17920,N_14688,N_14588);
nand U17921 (N_17921,N_14913,N_15299);
xor U17922 (N_17922,N_15682,N_14691);
and U17923 (N_17923,N_14678,N_14779);
or U17924 (N_17924,N_14167,N_15277);
xnor U17925 (N_17925,N_15294,N_15693);
nor U17926 (N_17926,N_14565,N_14849);
xor U17927 (N_17927,N_15933,N_14295);
or U17928 (N_17928,N_14321,N_15029);
nor U17929 (N_17929,N_15693,N_14016);
or U17930 (N_17930,N_15529,N_14661);
and U17931 (N_17931,N_15946,N_14046);
nand U17932 (N_17932,N_15877,N_14002);
or U17933 (N_17933,N_14543,N_14202);
xnor U17934 (N_17934,N_14824,N_14913);
nand U17935 (N_17935,N_15998,N_15355);
xnor U17936 (N_17936,N_15740,N_15965);
or U17937 (N_17937,N_15804,N_15024);
or U17938 (N_17938,N_15495,N_14245);
nand U17939 (N_17939,N_15907,N_15162);
and U17940 (N_17940,N_15349,N_14893);
or U17941 (N_17941,N_15125,N_15113);
xor U17942 (N_17942,N_15795,N_15767);
nand U17943 (N_17943,N_14789,N_14028);
xnor U17944 (N_17944,N_14021,N_15218);
or U17945 (N_17945,N_15592,N_15131);
or U17946 (N_17946,N_15459,N_14187);
nand U17947 (N_17947,N_15380,N_15473);
nand U17948 (N_17948,N_14546,N_15665);
xnor U17949 (N_17949,N_14981,N_15299);
xor U17950 (N_17950,N_14281,N_15560);
or U17951 (N_17951,N_15141,N_14198);
xnor U17952 (N_17952,N_15971,N_15890);
and U17953 (N_17953,N_15684,N_15584);
and U17954 (N_17954,N_14579,N_15661);
nand U17955 (N_17955,N_15245,N_14088);
nor U17956 (N_17956,N_15270,N_14088);
nand U17957 (N_17957,N_15561,N_14109);
nor U17958 (N_17958,N_15175,N_15188);
and U17959 (N_17959,N_14440,N_15770);
xnor U17960 (N_17960,N_15313,N_14970);
or U17961 (N_17961,N_14587,N_15218);
xor U17962 (N_17962,N_15284,N_15316);
nand U17963 (N_17963,N_15105,N_14129);
or U17964 (N_17964,N_15052,N_15452);
nor U17965 (N_17965,N_14559,N_14586);
or U17966 (N_17966,N_15341,N_14311);
nand U17967 (N_17967,N_15514,N_15068);
nand U17968 (N_17968,N_14960,N_14810);
nand U17969 (N_17969,N_14192,N_14209);
xor U17970 (N_17970,N_15657,N_15981);
xor U17971 (N_17971,N_15346,N_15168);
and U17972 (N_17972,N_15603,N_15341);
or U17973 (N_17973,N_15333,N_14548);
or U17974 (N_17974,N_15492,N_15595);
or U17975 (N_17975,N_15208,N_15180);
xnor U17976 (N_17976,N_14207,N_15181);
nand U17977 (N_17977,N_15028,N_14304);
or U17978 (N_17978,N_14205,N_14006);
nor U17979 (N_17979,N_14318,N_14685);
nor U17980 (N_17980,N_15717,N_15124);
xnor U17981 (N_17981,N_15071,N_14207);
xor U17982 (N_17982,N_14833,N_14016);
or U17983 (N_17983,N_14634,N_15849);
xnor U17984 (N_17984,N_14867,N_14426);
nand U17985 (N_17985,N_14992,N_15532);
xor U17986 (N_17986,N_15259,N_14009);
or U17987 (N_17987,N_15767,N_15938);
nand U17988 (N_17988,N_14028,N_15550);
nor U17989 (N_17989,N_14190,N_14197);
xnor U17990 (N_17990,N_15947,N_15996);
or U17991 (N_17991,N_15339,N_14647);
and U17992 (N_17992,N_14101,N_15440);
nand U17993 (N_17993,N_15058,N_14994);
xor U17994 (N_17994,N_14116,N_14798);
nor U17995 (N_17995,N_14573,N_14499);
nand U17996 (N_17996,N_14337,N_15668);
and U17997 (N_17997,N_14579,N_14045);
xnor U17998 (N_17998,N_15652,N_14314);
nor U17999 (N_17999,N_15437,N_14669);
nor U18000 (N_18000,N_16031,N_16522);
nand U18001 (N_18001,N_17508,N_16207);
and U18002 (N_18002,N_16924,N_16110);
xor U18003 (N_18003,N_16988,N_16216);
nor U18004 (N_18004,N_17364,N_16663);
and U18005 (N_18005,N_16117,N_16621);
xor U18006 (N_18006,N_17278,N_17481);
nand U18007 (N_18007,N_16520,N_17395);
or U18008 (N_18008,N_16349,N_16135);
nor U18009 (N_18009,N_17532,N_16166);
and U18010 (N_18010,N_16125,N_16456);
nor U18011 (N_18011,N_16423,N_17429);
xnor U18012 (N_18012,N_16549,N_16259);
xnor U18013 (N_18013,N_16037,N_17277);
nor U18014 (N_18014,N_16703,N_16454);
and U18015 (N_18015,N_17403,N_16208);
or U18016 (N_18016,N_16393,N_16900);
or U18017 (N_18017,N_16251,N_17863);
and U18018 (N_18018,N_16396,N_17576);
nor U18019 (N_18019,N_17698,N_17566);
nand U18020 (N_18020,N_16333,N_17969);
or U18021 (N_18021,N_16075,N_16694);
xnor U18022 (N_18022,N_16679,N_16485);
nor U18023 (N_18023,N_16253,N_16690);
nand U18024 (N_18024,N_16504,N_17067);
nand U18025 (N_18025,N_16488,N_17703);
nor U18026 (N_18026,N_17693,N_16513);
nor U18027 (N_18027,N_17327,N_17011);
nor U18028 (N_18028,N_17785,N_16072);
nand U18029 (N_18029,N_17606,N_17548);
nand U18030 (N_18030,N_17183,N_16677);
nand U18031 (N_18031,N_17664,N_16081);
nor U18032 (N_18032,N_17255,N_16991);
nand U18033 (N_18033,N_17402,N_17153);
nand U18034 (N_18034,N_16726,N_17546);
nand U18035 (N_18035,N_16580,N_16569);
nand U18036 (N_18036,N_17462,N_16652);
or U18037 (N_18037,N_17887,N_16426);
and U18038 (N_18038,N_16821,N_16838);
or U18039 (N_18039,N_16002,N_17691);
nor U18040 (N_18040,N_16535,N_16752);
nor U18041 (N_18041,N_17600,N_17727);
nor U18042 (N_18042,N_16430,N_16360);
nor U18043 (N_18043,N_17227,N_17074);
or U18044 (N_18044,N_16243,N_17964);
or U18045 (N_18045,N_16944,N_17332);
nor U18046 (N_18046,N_16565,N_17810);
and U18047 (N_18047,N_17045,N_16671);
nand U18048 (N_18048,N_17545,N_17708);
nand U18049 (N_18049,N_17040,N_16477);
or U18050 (N_18050,N_17284,N_16296);
nor U18051 (N_18051,N_17145,N_17467);
and U18052 (N_18052,N_16270,N_17534);
xnor U18053 (N_18053,N_16280,N_16611);
nand U18054 (N_18054,N_17601,N_16312);
and U18055 (N_18055,N_17289,N_16894);
and U18056 (N_18056,N_17083,N_16297);
nand U18057 (N_18057,N_17497,N_16959);
nor U18058 (N_18058,N_16658,N_17109);
xnor U18059 (N_18059,N_17916,N_17578);
and U18060 (N_18060,N_16500,N_16509);
and U18061 (N_18061,N_17052,N_16661);
nand U18062 (N_18062,N_17550,N_16892);
or U18063 (N_18063,N_17054,N_16132);
xnor U18064 (N_18064,N_16700,N_16313);
xor U18065 (N_18065,N_17266,N_17742);
or U18066 (N_18066,N_17059,N_16647);
and U18067 (N_18067,N_16862,N_17437);
or U18068 (N_18068,N_16749,N_16965);
xor U18069 (N_18069,N_16790,N_16033);
nand U18070 (N_18070,N_17199,N_17769);
nand U18071 (N_18071,N_17347,N_16066);
and U18072 (N_18072,N_17082,N_17243);
nor U18073 (N_18073,N_17156,N_17700);
xor U18074 (N_18074,N_16142,N_17718);
nor U18075 (N_18075,N_16842,N_16226);
nand U18076 (N_18076,N_17860,N_16878);
nor U18077 (N_18077,N_17811,N_16058);
or U18078 (N_18078,N_17044,N_16763);
or U18079 (N_18079,N_17732,N_17316);
nand U18080 (N_18080,N_17895,N_16318);
nor U18081 (N_18081,N_17886,N_17956);
or U18082 (N_18082,N_17086,N_16936);
and U18083 (N_18083,N_17998,N_16641);
nor U18084 (N_18084,N_16219,N_16401);
and U18085 (N_18085,N_16152,N_16888);
nand U18086 (N_18086,N_17837,N_16350);
nor U18087 (N_18087,N_17671,N_16371);
nand U18088 (N_18088,N_16188,N_16566);
nor U18089 (N_18089,N_17107,N_16890);
nand U18090 (N_18090,N_16306,N_17959);
nor U18091 (N_18091,N_16738,N_17306);
and U18092 (N_18092,N_17979,N_16819);
nor U18093 (N_18093,N_16436,N_17207);
nor U18094 (N_18094,N_17373,N_16684);
and U18095 (N_18095,N_17817,N_16608);
xnor U18096 (N_18096,N_16521,N_17802);
nor U18097 (N_18097,N_17046,N_16692);
nand U18098 (N_18098,N_16215,N_17276);
and U18099 (N_18099,N_16537,N_17116);
nor U18100 (N_18100,N_16351,N_17999);
xnor U18101 (N_18101,N_17101,N_16265);
xor U18102 (N_18102,N_17588,N_17461);
and U18103 (N_18103,N_17220,N_17854);
or U18104 (N_18104,N_17791,N_17908);
nand U18105 (N_18105,N_16435,N_17981);
or U18106 (N_18106,N_16478,N_17166);
or U18107 (N_18107,N_17120,N_16914);
nand U18108 (N_18108,N_16499,N_16314);
nor U18109 (N_18109,N_16229,N_17222);
nand U18110 (N_18110,N_16996,N_17536);
nand U18111 (N_18111,N_17423,N_16281);
or U18112 (N_18112,N_17178,N_16344);
or U18113 (N_18113,N_17988,N_16833);
nand U18114 (N_18114,N_17911,N_17400);
or U18115 (N_18115,N_16856,N_17833);
nor U18116 (N_18116,N_16343,N_17361);
or U18117 (N_18117,N_17747,N_17454);
nand U18118 (N_18118,N_17517,N_16990);
xnor U18119 (N_18119,N_16585,N_16088);
nand U18120 (N_18120,N_17165,N_17917);
xor U18121 (N_18121,N_17650,N_17737);
and U18122 (N_18122,N_16626,N_17146);
nand U18123 (N_18123,N_17441,N_16116);
nor U18124 (N_18124,N_17203,N_17420);
nand U18125 (N_18125,N_16732,N_16332);
xnor U18126 (N_18126,N_17894,N_17591);
and U18127 (N_18127,N_17874,N_16258);
nor U18128 (N_18128,N_17341,N_17675);
nor U18129 (N_18129,N_17619,N_16015);
xnor U18130 (N_18130,N_17378,N_16859);
nand U18131 (N_18131,N_16788,N_16680);
nand U18132 (N_18132,N_17254,N_16262);
and U18133 (N_18133,N_17329,N_17762);
nand U18134 (N_18134,N_16645,N_17557);
nor U18135 (N_18135,N_17320,N_17063);
nand U18136 (N_18136,N_16712,N_16872);
and U18137 (N_18137,N_16861,N_16622);
or U18138 (N_18138,N_17186,N_16595);
and U18139 (N_18139,N_16880,N_17504);
xnor U18140 (N_18140,N_16736,N_16687);
nor U18141 (N_18141,N_16649,N_16307);
nor U18142 (N_18142,N_16552,N_17648);
and U18143 (N_18143,N_17013,N_17035);
xor U18144 (N_18144,N_16773,N_16204);
and U18145 (N_18145,N_17921,N_16505);
nand U18146 (N_18146,N_16616,N_16234);
and U18147 (N_18147,N_17972,N_16906);
or U18148 (N_18148,N_16852,N_16145);
and U18149 (N_18149,N_17089,N_17608);
nand U18150 (N_18150,N_16570,N_17724);
nor U18151 (N_18151,N_16173,N_16919);
nand U18152 (N_18152,N_17147,N_17585);
or U18153 (N_18153,N_16148,N_17980);
and U18154 (N_18154,N_16612,N_16836);
or U18155 (N_18155,N_16627,N_17855);
and U18156 (N_18156,N_17442,N_16330);
or U18157 (N_18157,N_16252,N_17626);
and U18158 (N_18158,N_16292,N_17899);
or U18159 (N_18159,N_16278,N_16363);
or U18160 (N_18160,N_16413,N_16986);
and U18161 (N_18161,N_17716,N_16650);
and U18162 (N_18162,N_17391,N_16723);
nand U18163 (N_18163,N_17880,N_17189);
xnor U18164 (N_18164,N_17336,N_17351);
and U18165 (N_18165,N_17846,N_17159);
nand U18166 (N_18166,N_17365,N_17503);
or U18167 (N_18167,N_17936,N_16766);
or U18168 (N_18168,N_17296,N_17405);
and U18169 (N_18169,N_16999,N_16448);
nor U18170 (N_18170,N_16779,N_16146);
nand U18171 (N_18171,N_16184,N_16567);
and U18172 (N_18172,N_16034,N_16795);
or U18173 (N_18173,N_17603,N_17009);
or U18174 (N_18174,N_17656,N_17502);
or U18175 (N_18175,N_16689,N_17131);
nor U18176 (N_18176,N_16941,N_16245);
or U18177 (N_18177,N_17715,N_17989);
or U18178 (N_18178,N_17438,N_16196);
nand U18179 (N_18179,N_17738,N_16972);
or U18180 (N_18180,N_16778,N_17864);
or U18181 (N_18181,N_17092,N_17132);
or U18182 (N_18182,N_17098,N_16047);
or U18183 (N_18183,N_16083,N_17741);
nand U18184 (N_18184,N_16004,N_16023);
nor U18185 (N_18185,N_17767,N_17531);
and U18186 (N_18186,N_16682,N_16701);
or U18187 (N_18187,N_17016,N_16961);
xor U18188 (N_18188,N_17629,N_17398);
xnor U18189 (N_18189,N_16378,N_17923);
xor U18190 (N_18190,N_17560,N_17645);
nor U18191 (N_18191,N_16932,N_16161);
xnor U18192 (N_18192,N_16171,N_16120);
xor U18193 (N_18193,N_17494,N_16642);
and U18194 (N_18194,N_16271,N_16489);
nor U18195 (N_18195,N_16238,N_17519);
or U18196 (N_18196,N_16809,N_16716);
nand U18197 (N_18197,N_17303,N_16847);
xor U18198 (N_18198,N_16098,N_16303);
xor U18199 (N_18199,N_17271,N_16370);
and U18200 (N_18200,N_17318,N_16929);
nand U18201 (N_18201,N_17300,N_16734);
and U18202 (N_18202,N_17260,N_17283);
nor U18203 (N_18203,N_17205,N_16839);
and U18204 (N_18204,N_17382,N_17196);
nand U18205 (N_18205,N_16619,N_17770);
and U18206 (N_18206,N_16040,N_17191);
nand U18207 (N_18207,N_17155,N_17056);
nor U18208 (N_18208,N_17012,N_17498);
nor U18209 (N_18209,N_17685,N_17847);
nand U18210 (N_18210,N_17910,N_16260);
and U18211 (N_18211,N_16434,N_16302);
or U18212 (N_18212,N_17334,N_17511);
xor U18213 (N_18213,N_17376,N_17031);
or U18214 (N_18214,N_17935,N_17931);
and U18215 (N_18215,N_16523,N_17579);
or U18216 (N_18216,N_16884,N_16870);
nand U18217 (N_18217,N_17929,N_17488);
and U18218 (N_18218,N_16147,N_17805);
or U18219 (N_18219,N_17726,N_16346);
or U18220 (N_18220,N_16904,N_17310);
nor U18221 (N_18221,N_16187,N_17478);
or U18222 (N_18222,N_16867,N_17134);
nand U18223 (N_18223,N_16432,N_16084);
nor U18224 (N_18224,N_16452,N_16966);
and U18225 (N_18225,N_17292,N_16976);
xor U18226 (N_18226,N_16978,N_17665);
and U18227 (N_18227,N_16741,N_16022);
nand U18228 (N_18228,N_17448,N_17256);
xor U18229 (N_18229,N_17623,N_17932);
and U18230 (N_18230,N_16143,N_16327);
xor U18231 (N_18231,N_17944,N_17851);
nor U18232 (N_18232,N_17514,N_17669);
and U18233 (N_18233,N_17386,N_17195);
or U18234 (N_18234,N_16206,N_16197);
and U18235 (N_18235,N_17294,N_16221);
xor U18236 (N_18236,N_16175,N_17028);
and U18237 (N_18237,N_17003,N_16637);
nor U18238 (N_18238,N_17942,N_16543);
nand U18239 (N_18239,N_16767,N_16273);
nand U18240 (N_18240,N_16848,N_17778);
nor U18241 (N_18241,N_16099,N_17712);
xor U18242 (N_18242,N_16877,N_16254);
nor U18243 (N_18243,N_17496,N_16104);
nor U18244 (N_18244,N_17471,N_16064);
nor U18245 (N_18245,N_16662,N_16028);
or U18246 (N_18246,N_17072,N_16406);
xnor U18247 (N_18247,N_16342,N_17048);
nand U18248 (N_18248,N_17433,N_17465);
nor U18249 (N_18249,N_17406,N_17314);
nor U18250 (N_18250,N_17414,N_16277);
and U18251 (N_18251,N_17934,N_16169);
nor U18252 (N_18252,N_16131,N_16902);
nor U18253 (N_18253,N_17676,N_17794);
and U18254 (N_18254,N_17862,N_16656);
nor U18255 (N_18255,N_17215,N_16157);
xor U18256 (N_18256,N_16475,N_17412);
nand U18257 (N_18257,N_17902,N_16174);
nor U18258 (N_18258,N_17041,N_16101);
nor U18259 (N_18259,N_16071,N_17635);
nor U18260 (N_18260,N_17477,N_17486);
or U18261 (N_18261,N_17723,N_17312);
nand U18262 (N_18262,N_16213,N_16304);
and U18263 (N_18263,N_16843,N_16823);
or U18264 (N_18264,N_17466,N_17135);
nand U18265 (N_18265,N_16531,N_17865);
or U18266 (N_18266,N_16471,N_17527);
and U18267 (N_18267,N_16151,N_16203);
or U18268 (N_18268,N_16695,N_16263);
nor U18269 (N_18269,N_16742,N_17080);
nand U18270 (N_18270,N_16511,N_16052);
and U18271 (N_18271,N_16782,N_17088);
nor U18272 (N_18272,N_17873,N_17963);
nand U18273 (N_18273,N_16053,N_16056);
and U18274 (N_18274,N_16740,N_17661);
nor U18275 (N_18275,N_17240,N_16538);
xor U18276 (N_18276,N_17211,N_16881);
or U18277 (N_18277,N_16283,N_16381);
nor U18278 (N_18278,N_16310,N_16705);
xor U18279 (N_18279,N_16607,N_17301);
xnor U18280 (N_18280,N_17628,N_17404);
nor U18281 (N_18281,N_16025,N_16728);
nor U18282 (N_18282,N_16268,N_17350);
xor U18283 (N_18283,N_17977,N_17396);
nand U18284 (N_18284,N_17813,N_17535);
xor U18285 (N_18285,N_17001,N_16640);
nand U18286 (N_18286,N_16225,N_16233);
nor U18287 (N_18287,N_17139,N_17225);
or U18288 (N_18288,N_16643,N_17385);
nand U18289 (N_18289,N_17960,N_17309);
nand U18290 (N_18290,N_16806,N_16074);
nand U18291 (N_18291,N_17286,N_17464);
xor U18292 (N_18292,N_17955,N_17815);
nand U18293 (N_18293,N_16793,N_17787);
xnor U18294 (N_18294,N_17662,N_17446);
or U18295 (N_18295,N_17549,N_16319);
or U18296 (N_18296,N_17752,N_17479);
xnor U18297 (N_18297,N_16722,N_17968);
xnor U18298 (N_18298,N_16810,N_16294);
or U18299 (N_18299,N_17912,N_17581);
and U18300 (N_18300,N_16460,N_17991);
and U18301 (N_18301,N_17389,N_17909);
nor U18302 (N_18302,N_17017,N_16453);
or U18303 (N_18303,N_17374,N_16560);
and U18304 (N_18304,N_17093,N_16963);
or U18305 (N_18305,N_16121,N_17951);
xor U18306 (N_18306,N_17328,N_16968);
xnor U18307 (N_18307,N_17354,N_16442);
xor U18308 (N_18308,N_16630,N_16797);
nand U18309 (N_18309,N_16541,N_17111);
and U18310 (N_18310,N_16091,N_17982);
xor U18311 (N_18311,N_17043,N_17812);
xor U18312 (N_18312,N_16122,N_17143);
or U18313 (N_18313,N_17105,N_16077);
nor U18314 (N_18314,N_17551,N_17005);
xor U18315 (N_18315,N_16449,N_17838);
nor U18316 (N_18316,N_17961,N_17797);
nor U18317 (N_18317,N_17188,N_16657);
and U18318 (N_18318,N_17268,N_17340);
nand U18319 (N_18319,N_17136,N_16411);
and U18320 (N_18320,N_16231,N_16284);
or U18321 (N_18321,N_16392,N_16461);
or U18322 (N_18322,N_16879,N_17200);
nor U18323 (N_18323,N_17680,N_16405);
and U18324 (N_18324,N_17983,N_16674);
and U18325 (N_18325,N_17439,N_16198);
nand U18326 (N_18326,N_16124,N_17226);
nand U18327 (N_18327,N_17524,N_17493);
nor U18328 (N_18328,N_17681,N_16372);
or U18329 (N_18329,N_16237,N_16492);
xor U18330 (N_18330,N_16130,N_16026);
nor U18331 (N_18331,N_16018,N_16618);
and U18332 (N_18332,N_17025,N_17369);
nand U18333 (N_18333,N_16764,N_16168);
xnor U18334 (N_18334,N_16648,N_17622);
xor U18335 (N_18335,N_16664,N_16447);
nand U18336 (N_18336,N_16581,N_16967);
or U18337 (N_18337,N_16118,N_17324);
or U18338 (N_18338,N_16753,N_16445);
and U18339 (N_18339,N_17021,N_16547);
and U18340 (N_18340,N_16871,N_17515);
xor U18341 (N_18341,N_16185,N_17777);
or U18342 (N_18342,N_17435,N_16554);
nand U18343 (N_18343,N_17940,N_17825);
nor U18344 (N_18344,N_17331,N_16711);
or U18345 (N_18345,N_17106,N_16938);
or U18346 (N_18346,N_16068,N_17257);
and U18347 (N_18347,N_16186,N_16339);
or U18348 (N_18348,N_17709,N_16236);
or U18349 (N_18349,N_16796,N_16975);
nand U18350 (N_18350,N_17876,N_16775);
nand U18351 (N_18351,N_17006,N_16338);
nor U18352 (N_18352,N_16247,N_16923);
nor U18353 (N_18353,N_16154,N_17209);
xnor U18354 (N_18354,N_17121,N_17710);
xnor U18355 (N_18355,N_16391,N_17599);
nand U18356 (N_18356,N_16309,N_16119);
nand U18357 (N_18357,N_17996,N_17231);
nand U18358 (N_18358,N_16737,N_16420);
nand U18359 (N_18359,N_16368,N_17858);
and U18360 (N_18360,N_16352,N_17714);
and U18361 (N_18361,N_17799,N_16421);
and U18362 (N_18362,N_17816,N_16336);
and U18363 (N_18363,N_17541,N_16159);
and U18364 (N_18364,N_17064,N_16887);
or U18365 (N_18365,N_16156,N_16160);
nor U18366 (N_18366,N_17450,N_17501);
xor U18367 (N_18367,N_17490,N_16127);
nor U18368 (N_18368,N_16670,N_17058);
nand U18369 (N_18369,N_16419,N_16386);
and U18370 (N_18370,N_16651,N_16558);
nand U18371 (N_18371,N_16710,N_17335);
and U18372 (N_18372,N_17687,N_16320);
nor U18373 (N_18373,N_17237,N_16224);
or U18374 (N_18374,N_17879,N_16365);
xnor U18375 (N_18375,N_16628,N_17224);
nor U18376 (N_18376,N_17142,N_17580);
nand U18377 (N_18377,N_16597,N_17239);
or U18378 (N_18378,N_16163,N_17452);
and U18379 (N_18379,N_16223,N_17353);
or U18380 (N_18380,N_17436,N_16718);
or U18381 (N_18381,N_16954,N_17945);
xor U18382 (N_18382,N_17282,N_17247);
xor U18383 (N_18383,N_16772,N_17213);
nor U18384 (N_18384,N_16592,N_17062);
and U18385 (N_18385,N_16745,N_16678);
nand U18386 (N_18386,N_17377,N_16472);
or U18387 (N_18387,N_17029,N_17828);
nand U18388 (N_18388,N_16542,N_16109);
and U18389 (N_18389,N_16379,N_17649);
and U18390 (N_18390,N_16355,N_16593);
or U18391 (N_18391,N_16189,N_16733);
and U18392 (N_18392,N_16831,N_16285);
xor U18393 (N_18393,N_17444,N_16623);
nor U18394 (N_18394,N_17674,N_17728);
xor U18395 (N_18395,N_16133,N_16586);
nand U18396 (N_18396,N_16688,N_16617);
nor U18397 (N_18397,N_16329,N_16389);
nor U18398 (N_18398,N_16340,N_16202);
xor U18399 (N_18399,N_17768,N_17250);
nor U18400 (N_18400,N_16707,N_16602);
and U18401 (N_18401,N_17636,N_16257);
or U18402 (N_18402,N_16080,N_16376);
xor U18403 (N_18403,N_17049,N_16050);
and U18404 (N_18404,N_16358,N_17157);
xor U18405 (N_18405,N_16212,N_16973);
or U18406 (N_18406,N_16761,N_17325);
nand U18407 (N_18407,N_17933,N_16668);
xnor U18408 (N_18408,N_16450,N_17866);
nand U18409 (N_18409,N_16780,N_17053);
nand U18410 (N_18410,N_17174,N_17896);
nand U18411 (N_18411,N_16427,N_17489);
nand U18412 (N_18412,N_17249,N_16041);
nand U18413 (N_18413,N_17824,N_17270);
nor U18414 (N_18414,N_17163,N_17753);
xnor U18415 (N_18415,N_17798,N_17843);
xor U18416 (N_18416,N_16964,N_17372);
and U18417 (N_18417,N_17678,N_17173);
or U18418 (N_18418,N_17459,N_16138);
or U18419 (N_18419,N_17238,N_16815);
xnor U18420 (N_18420,N_16113,N_16562);
xnor U18421 (N_18421,N_16463,N_17154);
xor U18422 (N_18422,N_17228,N_17458);
nor U18423 (N_18423,N_17647,N_16907);
or U18424 (N_18424,N_16743,N_16613);
nand U18425 (N_18425,N_17836,N_17590);
xor U18426 (N_18426,N_16889,N_17766);
nand U18427 (N_18427,N_17509,N_16899);
and U18428 (N_18428,N_17015,N_16498);
nand U18429 (N_18429,N_17133,N_17500);
nand U18430 (N_18430,N_17288,N_16503);
and U18431 (N_18431,N_17079,N_17904);
or U18432 (N_18432,N_17878,N_17516);
and U18433 (N_18433,N_16013,N_16786);
or U18434 (N_18434,N_16993,N_17850);
xnor U18435 (N_18435,N_16179,N_16055);
xnor U18436 (N_18436,N_17611,N_17589);
nand U18437 (N_18437,N_16334,N_16863);
nor U18438 (N_18438,N_16873,N_16719);
or U18439 (N_18439,N_17542,N_16012);
and U18440 (N_18440,N_16992,N_16359);
or U18441 (N_18441,N_16347,N_16624);
or U18442 (N_18442,N_16462,N_16242);
xor U18443 (N_18443,N_16931,N_16556);
and U18444 (N_18444,N_17949,N_16639);
nor U18445 (N_18445,N_16770,N_17469);
or U18446 (N_18446,N_16298,N_17537);
xor U18447 (N_18447,N_16905,N_16828);
nor U18448 (N_18448,N_17707,N_16027);
nand U18449 (N_18449,N_16162,N_16275);
and U18450 (N_18450,N_16007,N_17651);
or U18451 (N_18451,N_17598,N_17427);
xor U18452 (N_18452,N_16199,N_17010);
nor U18453 (N_18453,N_16844,N_16776);
or U18454 (N_18454,N_16123,N_16853);
nand U18455 (N_18455,N_16854,N_16735);
and U18456 (N_18456,N_17002,N_16955);
and U18457 (N_18457,N_17725,N_16006);
and U18458 (N_18458,N_16200,N_16096);
and U18459 (N_18459,N_17884,N_16059);
nor U18460 (N_18460,N_17388,N_17771);
xnor U18461 (N_18461,N_17612,N_16502);
and U18462 (N_18462,N_17686,N_16417);
nor U18463 (N_18463,N_17672,N_16410);
and U18464 (N_18464,N_17229,N_17966);
or U18465 (N_18465,N_16759,N_17482);
or U18466 (N_18466,N_16424,N_17954);
nor U18467 (N_18467,N_16194,N_16128);
and U18468 (N_18468,N_16514,N_16603);
and U18469 (N_18469,N_17171,N_16474);
and U18470 (N_18470,N_17024,N_16777);
or U18471 (N_18471,N_17317,N_16291);
nor U18472 (N_18472,N_16949,N_17938);
nand U18473 (N_18473,N_16416,N_17475);
nor U18474 (N_18474,N_17750,N_16079);
and U18475 (N_18475,N_17463,N_17366);
or U18476 (N_18476,N_16920,N_17652);
nor U18477 (N_18477,N_17822,N_17586);
or U18478 (N_18478,N_16491,N_17883);
and U18479 (N_18479,N_16898,N_17584);
xnor U18480 (N_18480,N_16362,N_16153);
xor U18481 (N_18481,N_16849,N_16942);
or U18482 (N_18482,N_17861,N_16882);
and U18483 (N_18483,N_16493,N_17460);
or U18484 (N_18484,N_17091,N_16137);
and U18485 (N_18485,N_17117,N_16846);
xor U18486 (N_18486,N_16308,N_16895);
xnor U18487 (N_18487,N_16183,N_16102);
nand U18488 (N_18488,N_16400,N_17216);
and U18489 (N_18489,N_17470,N_16561);
and U18490 (N_18490,N_17640,N_16606);
nor U18491 (N_18491,N_16459,N_16691);
xnor U18492 (N_18492,N_17180,N_17177);
nor U18493 (N_18493,N_17418,N_17841);
or U18494 (N_18494,N_16390,N_16129);
and U18495 (N_18495,N_16785,N_17162);
and U18496 (N_18496,N_16341,N_17272);
nand U18497 (N_18497,N_16572,N_17957);
and U18498 (N_18498,N_17543,N_16382);
xor U18499 (N_18499,N_16811,N_16095);
xnor U18500 (N_18500,N_16524,N_16532);
and U18501 (N_18501,N_16425,N_16575);
nand U18502 (N_18502,N_16655,N_16526);
nor U18503 (N_18503,N_17069,N_17941);
xor U18504 (N_18504,N_16087,N_17692);
nand U18505 (N_18505,N_16757,N_17995);
nor U18506 (N_18506,N_16227,N_16754);
or U18507 (N_18507,N_16654,N_16578);
xor U18508 (N_18508,N_17765,N_17042);
xor U18509 (N_18509,N_16693,N_16792);
and U18510 (N_18510,N_17337,N_17359);
and U18511 (N_18511,N_17763,N_16108);
nor U18512 (N_18512,N_16755,N_16858);
nand U18513 (N_18513,N_16495,N_17308);
nor U18514 (N_18514,N_16218,N_17345);
xnor U18515 (N_18515,N_16484,N_17773);
or U18516 (N_18516,N_17735,N_17447);
or U18517 (N_18517,N_17592,N_16791);
nor U18518 (N_18518,N_16666,N_17425);
or U18519 (N_18519,N_17974,N_16533);
or U18520 (N_18520,N_17814,N_17803);
nor U18521 (N_18521,N_17047,N_16353);
and U18522 (N_18522,N_17407,N_17889);
nor U18523 (N_18523,N_17533,N_16794);
xor U18524 (N_18524,N_17206,N_17809);
nand U18525 (N_18525,N_17682,N_16496);
or U18526 (N_18526,N_17559,N_16337);
nand U18527 (N_18527,N_17667,N_17233);
nor U18528 (N_18528,N_16771,N_17877);
or U18529 (N_18529,N_16322,N_16177);
nand U18530 (N_18530,N_16982,N_16093);
xnor U18531 (N_18531,N_16286,N_16114);
xnor U18532 (N_18532,N_17218,N_17161);
or U18533 (N_18533,N_17422,N_17018);
nand U18534 (N_18534,N_17319,N_17483);
nor U18535 (N_18535,N_17780,N_17633);
xor U18536 (N_18536,N_16660,N_16255);
and U18537 (N_18537,N_16164,N_16437);
xnor U18538 (N_18538,N_17907,N_16997);
and U18539 (N_18539,N_17164,N_16141);
nor U18540 (N_18540,N_17683,N_16945);
xor U18541 (N_18541,N_16295,N_16948);
nand U18542 (N_18542,N_17244,N_16576);
and U18543 (N_18543,N_16063,N_16272);
nand U18544 (N_18544,N_17212,N_17169);
nor U18545 (N_18545,N_17108,N_17019);
and U18546 (N_18546,N_16086,N_16172);
nor U18547 (N_18547,N_17520,N_17946);
and U18548 (N_18548,N_16629,N_16636);
or U18549 (N_18549,N_16675,N_17749);
xnor U18550 (N_18550,N_17291,N_17795);
nor U18551 (N_18551,N_16927,N_16596);
or U18552 (N_18552,N_16032,N_16364);
or U18553 (N_18553,N_17845,N_16913);
or U18554 (N_18554,N_16090,N_16891);
and U18555 (N_18555,N_17760,N_16325);
nor U18556 (N_18556,N_16044,N_16457);
nand U18557 (N_18557,N_17443,N_17563);
or U18558 (N_18558,N_17717,N_17118);
xnor U18559 (N_18559,N_17138,N_17736);
or U18560 (N_18560,N_16583,N_16540);
and U18561 (N_18561,N_17705,N_16165);
or U18562 (N_18562,N_17358,N_17241);
or U18563 (N_18563,N_16519,N_17745);
or U18564 (N_18564,N_17605,N_16910);
or U18565 (N_18565,N_16397,N_17823);
nand U18566 (N_18566,N_17744,N_17526);
or U18567 (N_18567,N_17970,N_16893);
nor U18568 (N_18568,N_16638,N_16813);
nand U18569 (N_18569,N_17616,N_17906);
xor U18570 (N_18570,N_16003,N_17037);
nand U18571 (N_18571,N_16274,N_17428);
nor U18572 (N_18572,N_17621,N_17431);
xor U18573 (N_18573,N_17095,N_16323);
nand U18574 (N_18574,N_16402,N_17641);
and U18575 (N_18575,N_16818,N_16876);
or U18576 (N_18576,N_16149,N_16250);
xnor U18577 (N_18577,N_16706,N_16357);
and U18578 (N_18578,N_17217,N_17918);
nor U18579 (N_18579,N_17066,N_17333);
nor U18580 (N_18580,N_17379,N_17182);
xnor U18581 (N_18581,N_17262,N_16201);
nand U18582 (N_18582,N_17060,N_17026);
xnor U18583 (N_18583,N_17617,N_17819);
nand U18584 (N_18584,N_16220,N_17832);
xor U18585 (N_18585,N_16431,N_16610);
nor U18586 (N_18586,N_17421,N_16486);
nor U18587 (N_18587,N_17706,N_17761);
nor U18588 (N_18588,N_17506,N_17528);
or U18589 (N_18589,N_16345,N_17657);
nand U18590 (N_18590,N_17684,N_16822);
nand U18591 (N_18591,N_17820,N_17513);
nor U18592 (N_18592,N_17654,N_16422);
or U18593 (N_18593,N_17870,N_17722);
and U18594 (N_18594,N_16326,N_17947);
or U18595 (N_18595,N_16490,N_17492);
xor U18596 (N_18596,N_17697,N_17399);
or U18597 (N_18597,N_16466,N_17141);
nand U18598 (N_18598,N_17572,N_16729);
and U18599 (N_18599,N_16958,N_17679);
nand U18600 (N_18600,N_16444,N_17187);
nor U18601 (N_18601,N_17655,N_17115);
nor U18602 (N_18602,N_17901,N_16317);
nor U18603 (N_18603,N_16713,N_17859);
and U18604 (N_18604,N_17793,N_16008);
xnor U18605 (N_18605,N_16399,N_17130);
nor U18606 (N_18606,N_17673,N_17445);
xnor U18607 (N_18607,N_17202,N_16774);
nor U18608 (N_18608,N_16646,N_16957);
xor U18609 (N_18609,N_17285,N_16747);
or U18610 (N_18610,N_16057,N_17562);
xnor U18611 (N_18611,N_17952,N_17349);
xnor U18612 (N_18612,N_17313,N_16506);
nand U18613 (N_18613,N_16293,N_17607);
nand U18614 (N_18614,N_16019,N_16439);
and U18615 (N_18615,N_17219,N_16940);
nor U18616 (N_18616,N_16515,N_16394);
and U18617 (N_18617,N_16483,N_17638);
and U18618 (N_18618,N_17057,N_17305);
and U18619 (N_18619,N_17539,N_17258);
nand U18620 (N_18620,N_16539,N_16758);
or U18621 (N_18621,N_16480,N_16935);
nor U18622 (N_18622,N_16106,N_17842);
and U18623 (N_18623,N_17711,N_16969);
and U18624 (N_18624,N_17898,N_17985);
or U18625 (N_18625,N_16686,N_17927);
nor U18626 (N_18626,N_17076,N_16126);
nand U18627 (N_18627,N_16769,N_16908);
and U18628 (N_18628,N_16190,N_16798);
or U18629 (N_18629,N_17279,N_17892);
or U18630 (N_18630,N_17801,N_16851);
nor U18631 (N_18631,N_17094,N_17644);
nor U18632 (N_18632,N_17758,N_16375);
and U18633 (N_18633,N_17393,N_17618);
xnor U18634 (N_18634,N_16868,N_16829);
nand U18635 (N_18635,N_16559,N_16469);
nor U18636 (N_18636,N_17610,N_16546);
or U18637 (N_18637,N_17126,N_17070);
or U18638 (N_18638,N_17759,N_17593);
or U18639 (N_18639,N_16748,N_16373);
xor U18640 (N_18640,N_17073,N_16527);
nor U18641 (N_18641,N_17529,N_17100);
nand U18642 (N_18642,N_17468,N_16267);
xnor U18643 (N_18643,N_17574,N_17848);
or U18644 (N_18644,N_17179,N_17302);
nand U18645 (N_18645,N_17694,N_17357);
nor U18646 (N_18646,N_16916,N_16625);
and U18647 (N_18647,N_16182,N_17577);
nand U18648 (N_18648,N_16407,N_16604);
or U18649 (N_18649,N_16762,N_17987);
or U18650 (N_18650,N_16014,N_16438);
and U18651 (N_18651,N_17004,N_16544);
nand U18652 (N_18652,N_17208,N_16210);
or U18653 (N_18653,N_17632,N_17627);
and U18654 (N_18654,N_17888,N_17782);
nand U18655 (N_18655,N_17129,N_17090);
and U18656 (N_18656,N_16441,N_16577);
xor U18657 (N_18657,N_16301,N_17835);
nor U18658 (N_18658,N_17235,N_17821);
and U18659 (N_18659,N_16299,N_16107);
nand U18660 (N_18660,N_16105,N_17204);
xnor U18661 (N_18661,N_16467,N_17127);
and U18662 (N_18662,N_17077,N_17844);
nand U18663 (N_18663,N_17007,N_16765);
or U18664 (N_18664,N_16653,N_16814);
nand U18665 (N_18665,N_16266,N_16100);
nand U18666 (N_18666,N_17784,N_17800);
xor U18667 (N_18667,N_17201,N_16615);
nor U18668 (N_18668,N_17387,N_16525);
nor U18669 (N_18669,N_17096,N_16170);
nor U18670 (N_18670,N_16590,N_16062);
nor U18671 (N_18671,N_17734,N_16140);
or U18672 (N_18672,N_16746,N_17913);
xor U18673 (N_18673,N_16950,N_16065);
nand U18674 (N_18674,N_17521,N_17781);
or U18675 (N_18675,N_16517,N_16835);
nor U18676 (N_18676,N_16614,N_16550);
xor U18677 (N_18677,N_17702,N_17808);
nor U18678 (N_18678,N_16802,N_17232);
and U18679 (N_18679,N_17948,N_16817);
nand U18680 (N_18680,N_16134,N_16812);
nor U18681 (N_18681,N_16097,N_16883);
or U18682 (N_18682,N_16699,N_16139);
xor U18683 (N_18683,N_16017,N_16176);
nor U18684 (N_18684,N_16799,N_16985);
nor U18685 (N_18685,N_16016,N_17253);
nor U18686 (N_18686,N_16832,N_17530);
nand U18687 (N_18687,N_17299,N_16584);
nand U18688 (N_18688,N_16568,N_17660);
nor U18689 (N_18689,N_17124,N_16896);
or U18690 (N_18690,N_16516,N_16787);
nor U18691 (N_18691,N_17295,N_17381);
nor U18692 (N_18692,N_16451,N_17476);
nand U18693 (N_18693,N_16563,N_17522);
nor U18694 (N_18694,N_16800,N_17190);
nor U18695 (N_18695,N_17152,N_16115);
and U18696 (N_18696,N_16952,N_16412);
or U18697 (N_18697,N_17326,N_17721);
or U18698 (N_18698,N_16903,N_17210);
nand U18699 (N_18699,N_16768,N_17455);
or U18700 (N_18700,N_16696,N_16054);
nor U18701 (N_18701,N_16937,N_16760);
xor U18702 (N_18702,N_17480,N_17367);
and U18703 (N_18703,N_17571,N_17355);
nor U18704 (N_18704,N_17248,N_16011);
or U18705 (N_18705,N_17356,N_17984);
xor U18706 (N_18706,N_17624,N_16249);
nor U18707 (N_18707,N_17167,N_17038);
or U18708 (N_18708,N_17034,N_16361);
or U18709 (N_18709,N_17642,N_16518);
nand U18710 (N_18710,N_16865,N_17290);
or U18711 (N_18711,N_16356,N_17993);
or U18712 (N_18712,N_16579,N_17344);
and U18713 (N_18713,N_17078,N_16409);
or U18714 (N_18714,N_17776,N_16446);
xnor U18715 (N_18715,N_17756,N_17754);
xor U18716 (N_18716,N_16886,N_17775);
and U18717 (N_18717,N_16669,N_17193);
nand U18718 (N_18718,N_17122,N_16348);
nand U18719 (N_18719,N_17699,N_16803);
or U18720 (N_18720,N_16721,N_17625);
nor U18721 (N_18721,N_16385,N_16594);
nand U18722 (N_18722,N_16067,N_16573);
or U18723 (N_18723,N_16901,N_17051);
nand U18724 (N_18724,N_17339,N_17125);
nand U18725 (N_18725,N_17417,N_17834);
nor U18726 (N_18726,N_17897,N_17273);
nor U18727 (N_18727,N_16983,N_16981);
nor U18728 (N_18728,N_16864,N_17583);
xor U18729 (N_18729,N_16473,N_17137);
xnor U18730 (N_18730,N_16953,N_17719);
xor U18731 (N_18731,N_17261,N_17620);
xnor U18732 (N_18732,N_17371,N_16497);
nand U18733 (N_18733,N_17348,N_17900);
nand U18734 (N_18734,N_17390,N_17830);
xnor U18735 (N_18735,N_16042,N_16970);
nor U18736 (N_18736,N_17099,N_17965);
and U18737 (N_18737,N_16875,N_16193);
or U18738 (N_18738,N_17926,N_16725);
or U18739 (N_18739,N_16820,N_17806);
nand U18740 (N_18740,N_16551,N_16974);
and U18741 (N_18741,N_17140,N_17410);
xnor U18742 (N_18742,N_16956,N_16915);
xor U18743 (N_18743,N_17287,N_17071);
and U18744 (N_18744,N_17856,N_17392);
nand U18745 (N_18745,N_17990,N_17739);
or U18746 (N_18746,N_17653,N_16367);
nand U18747 (N_18747,N_16943,N_17839);
nand U18748 (N_18748,N_16354,N_16951);
nor U18749 (N_18749,N_17330,N_16279);
and U18750 (N_18750,N_17362,N_16020);
nand U18751 (N_18751,N_17875,N_17994);
or U18752 (N_18752,N_16789,N_16264);
nand U18753 (N_18753,N_16501,N_16009);
nand U18754 (N_18754,N_16681,N_16979);
nand U18755 (N_18755,N_16739,N_16934);
or U18756 (N_18756,N_16545,N_16191);
xor U18757 (N_18757,N_16092,N_17604);
or U18758 (N_18758,N_16418,N_17594);
and U18759 (N_18759,N_16632,N_17055);
or U18760 (N_18760,N_17950,N_16962);
nand U18761 (N_18761,N_17905,N_17265);
xor U18762 (N_18762,N_17036,N_17323);
nand U18763 (N_18763,N_16667,N_16388);
xnor U18764 (N_18764,N_16155,N_17112);
and U18765 (N_18765,N_16001,N_17553);
nand U18766 (N_18766,N_17144,N_17197);
and U18767 (N_18767,N_17573,N_16926);
xor U18768 (N_18768,N_17540,N_16672);
and U18769 (N_18769,N_17185,N_17602);
and U18770 (N_18770,N_16807,N_16269);
nor U18771 (N_18771,N_17973,N_17755);
nor U18772 (N_18772,N_16824,N_16144);
nor U18773 (N_18773,N_16458,N_17690);
and U18774 (N_18774,N_17252,N_16971);
and U18775 (N_18775,N_16720,N_17867);
xor U18776 (N_18776,N_16178,N_16487);
xnor U18777 (N_18777,N_17677,N_17730);
nor U18778 (N_18778,N_17170,N_16324);
nor U18779 (N_18779,N_17796,N_16756);
nand U18780 (N_18780,N_17786,N_16676);
and U18781 (N_18781,N_17565,N_17236);
nand U18782 (N_18782,N_17558,N_16633);
and U18783 (N_18783,N_17434,N_16384);
or U18784 (N_18784,N_16414,N_16536);
nor U18785 (N_18785,N_16232,N_17432);
nor U18786 (N_18786,N_16804,N_16035);
and U18787 (N_18787,N_17587,N_17409);
nor U18788 (N_18788,N_16928,N_17790);
or U18789 (N_18789,N_16380,N_17720);
and U18790 (N_18790,N_16665,N_17595);
nand U18791 (N_18791,N_16195,N_16933);
and U18792 (N_18792,N_17783,N_16061);
nand U18793 (N_18793,N_16038,N_16103);
and U18794 (N_18794,N_17050,N_17788);
or U18795 (N_18795,N_17928,N_17192);
and U18796 (N_18796,N_16599,N_16046);
nand U18797 (N_18797,N_17772,N_17552);
xor U18798 (N_18798,N_17000,N_17176);
and U18799 (N_18799,N_17943,N_16730);
or U18800 (N_18800,N_17663,N_16398);
xnor U18801 (N_18801,N_16947,N_17413);
and U18802 (N_18802,N_17172,N_17751);
nor U18803 (N_18803,N_17554,N_17430);
xnor U18804 (N_18804,N_17829,N_16977);
nor U18805 (N_18805,N_16530,N_17380);
or U18806 (N_18806,N_16724,N_16897);
and U18807 (N_18807,N_17085,N_16082);
and U18808 (N_18808,N_17149,N_17868);
and U18809 (N_18809,N_17150,N_17807);
nand U18810 (N_18810,N_17251,N_16589);
or U18811 (N_18811,N_17953,N_16609);
or U18812 (N_18812,N_16366,N_17596);
and U18813 (N_18813,N_17637,N_16885);
or U18814 (N_18814,N_17882,N_16209);
xor U18815 (N_18815,N_16857,N_16918);
or U18816 (N_18816,N_17561,N_17792);
nor U18817 (N_18817,N_16049,N_17962);
and U18818 (N_18818,N_16415,N_16510);
nor U18819 (N_18819,N_16866,N_16801);
xor U18820 (N_18820,N_16909,N_16244);
and U18821 (N_18821,N_17242,N_17293);
nand U18822 (N_18822,N_17368,N_16548);
nor U18823 (N_18823,N_16930,N_17221);
or U18824 (N_18824,N_16288,N_17986);
nand U18825 (N_18825,N_16048,N_17871);
or U18826 (N_18826,N_17597,N_16850);
and U18827 (N_18827,N_16222,N_17505);
and U18828 (N_18828,N_17570,N_16464);
nand U18829 (N_18829,N_17670,N_17689);
xnor U18830 (N_18830,N_17615,N_17495);
nand U18831 (N_18831,N_17731,N_16377);
xnor U18832 (N_18832,N_17102,N_17614);
nor U18833 (N_18833,N_17924,N_17582);
and U18834 (N_18834,N_16702,N_16564);
or U18835 (N_18835,N_17696,N_17639);
nor U18836 (N_18836,N_16211,N_16246);
nand U18837 (N_18837,N_17397,N_17322);
xnor U18838 (N_18838,N_17297,N_16600);
and U18839 (N_18839,N_16634,N_17992);
and U18840 (N_18840,N_16587,N_17774);
xor U18841 (N_18841,N_16214,N_17748);
and U18842 (N_18842,N_16750,N_17491);
or U18843 (N_18843,N_16261,N_16697);
and U18844 (N_18844,N_16591,N_17740);
nor U18845 (N_18845,N_17487,N_17363);
and U18846 (N_18846,N_16256,N_17852);
or U18847 (N_18847,N_17087,N_16321);
and U18848 (N_18848,N_17457,N_16827);
nand U18849 (N_18849,N_17643,N_17818);
nor U18850 (N_18850,N_16781,N_17075);
or U18851 (N_18851,N_17779,N_16855);
nor U18852 (N_18852,N_16403,N_17922);
and U18853 (N_18853,N_16874,N_17872);
nor U18854 (N_18854,N_17885,N_16869);
nor U18855 (N_18855,N_16582,N_17831);
nor U18856 (N_18856,N_16290,N_17030);
nor U18857 (N_18857,N_17321,N_16939);
nor U18858 (N_18858,N_17181,N_16024);
and U18859 (N_18859,N_17032,N_17456);
or U18860 (N_18860,N_16094,N_17264);
and U18861 (N_18861,N_16840,N_16089);
or U18862 (N_18862,N_17523,N_17198);
and U18863 (N_18863,N_16476,N_16708);
nor U18864 (N_18864,N_16029,N_17424);
or U18865 (N_18865,N_17568,N_17473);
nor U18866 (N_18866,N_16825,N_16507);
nand U18867 (N_18867,N_16704,N_17757);
and U18868 (N_18868,N_16644,N_17245);
and U18869 (N_18869,N_17128,N_17827);
nand U18870 (N_18870,N_16841,N_17925);
xnor U18871 (N_18871,N_16429,N_16512);
or U18872 (N_18872,N_17033,N_17449);
xnor U18873 (N_18873,N_16481,N_17804);
nor U18874 (N_18874,N_16395,N_17510);
nor U18875 (N_18875,N_16717,N_17743);
nor U18876 (N_18876,N_17426,N_17103);
nand U18877 (N_18877,N_17958,N_16911);
or U18878 (N_18878,N_17370,N_17849);
nor U18879 (N_18879,N_17223,N_16989);
xnor U18880 (N_18880,N_17688,N_17569);
xor U18881 (N_18881,N_17113,N_16987);
xor U18882 (N_18882,N_17104,N_16922);
and U18883 (N_18883,N_17416,N_17544);
xnor U18884 (N_18884,N_17110,N_17474);
nand U18885 (N_18885,N_17097,N_16287);
xor U18886 (N_18886,N_17027,N_16111);
and U18887 (N_18887,N_17123,N_17275);
nand U18888 (N_18888,N_16239,N_16078);
nand U18889 (N_18889,N_16374,N_16408);
nor U18890 (N_18890,N_17564,N_16315);
xor U18891 (N_18891,N_16112,N_16571);
and U18892 (N_18892,N_17184,N_17383);
nor U18893 (N_18893,N_16150,N_16030);
nand U18894 (N_18894,N_17556,N_16043);
nor U18895 (N_18895,N_17214,N_16248);
nor U18896 (N_18896,N_17704,N_17315);
xnor U18897 (N_18897,N_17971,N_16228);
nor U18898 (N_18898,N_17634,N_17065);
or U18899 (N_18899,N_17484,N_16557);
and U18900 (N_18900,N_16783,N_16468);
or U18901 (N_18901,N_17668,N_16921);
or U18902 (N_18902,N_17903,N_17408);
or U18903 (N_18903,N_17346,N_16995);
and U18904 (N_18904,N_17342,N_16482);
nor U18905 (N_18905,N_16404,N_16685);
nand U18906 (N_18906,N_16300,N_17512);
nor U18907 (N_18907,N_16960,N_16010);
nand U18908 (N_18908,N_17613,N_17890);
and U18909 (N_18909,N_16830,N_16834);
and U18910 (N_18910,N_17789,N_17194);
and U18911 (N_18911,N_17914,N_16826);
or U18912 (N_18912,N_17975,N_17472);
and U18913 (N_18913,N_16289,N_16076);
and U18914 (N_18914,N_16282,N_17419);
xor U18915 (N_18915,N_16305,N_16731);
nand U18916 (N_18916,N_16751,N_16470);
xnor U18917 (N_18917,N_17840,N_16683);
nand U18918 (N_18918,N_17567,N_17263);
nand U18919 (N_18919,N_16816,N_16192);
nand U18920 (N_18920,N_17881,N_17609);
nor U18921 (N_18921,N_16073,N_17826);
or U18922 (N_18922,N_17547,N_17659);
nand U18923 (N_18923,N_16387,N_17151);
xor U18924 (N_18924,N_16659,N_16980);
nand U18925 (N_18925,N_16051,N_17893);
nand U18926 (N_18926,N_16440,N_17352);
or U18927 (N_18927,N_17246,N_17746);
nand U18928 (N_18928,N_16039,N_17160);
nand U18929 (N_18929,N_17338,N_16998);
nand U18930 (N_18930,N_16230,N_17701);
xor U18931 (N_18931,N_16534,N_16479);
nor U18932 (N_18932,N_16598,N_16069);
or U18933 (N_18933,N_16428,N_17976);
nor U18934 (N_18934,N_16601,N_17014);
and U18935 (N_18935,N_16605,N_17061);
or U18936 (N_18936,N_17274,N_16555);
nor U18937 (N_18937,N_17343,N_17008);
or U18938 (N_18938,N_16925,N_16369);
nor U18939 (N_18939,N_16217,N_16205);
xnor U18940 (N_18940,N_16508,N_17930);
nand U18941 (N_18941,N_17451,N_17411);
nor U18942 (N_18942,N_17658,N_17575);
and U18943 (N_18943,N_17267,N_17453);
nor U18944 (N_18944,N_17631,N_16433);
xnor U18945 (N_18945,N_16181,N_16167);
or U18946 (N_18946,N_17937,N_16311);
nand U18947 (N_18947,N_16494,N_17538);
or U18948 (N_18948,N_16553,N_16000);
nand U18949 (N_18949,N_17384,N_16837);
or U18950 (N_18950,N_16946,N_16784);
xor U18951 (N_18951,N_16845,N_17375);
or U18952 (N_18952,N_17401,N_17259);
or U18953 (N_18953,N_17695,N_17891);
or U18954 (N_18954,N_16715,N_17234);
nor U18955 (N_18955,N_17525,N_17869);
or U18956 (N_18956,N_17485,N_17168);
or U18957 (N_18957,N_17920,N_17039);
nand U18958 (N_18958,N_16036,N_17280);
or U18959 (N_18959,N_16045,N_16529);
and U18960 (N_18960,N_16994,N_16465);
nand U18961 (N_18961,N_17729,N_17555);
and U18962 (N_18962,N_16714,N_16060);
nand U18963 (N_18963,N_16383,N_16620);
nand U18964 (N_18964,N_16635,N_16158);
and U18965 (N_18965,N_17978,N_16673);
and U18966 (N_18966,N_17499,N_17394);
and U18967 (N_18967,N_17630,N_17230);
or U18968 (N_18968,N_16005,N_17175);
nand U18969 (N_18969,N_17311,N_17415);
xnor U18970 (N_18970,N_17666,N_16331);
and U18971 (N_18971,N_17939,N_16180);
xnor U18972 (N_18972,N_16574,N_17733);
xor U18973 (N_18973,N_16455,N_16085);
nor U18974 (N_18974,N_17020,N_17269);
nand U18975 (N_18975,N_17158,N_17360);
or U18976 (N_18976,N_16984,N_16698);
and U18977 (N_18977,N_17713,N_16235);
nand U18978 (N_18978,N_17919,N_16709);
and U18979 (N_18979,N_16727,N_17068);
and U18980 (N_18980,N_16276,N_17646);
and U18981 (N_18981,N_16070,N_17084);
nor U18982 (N_18982,N_17915,N_17440);
nand U18983 (N_18983,N_16744,N_17298);
and U18984 (N_18984,N_16808,N_17857);
nor U18985 (N_18985,N_17997,N_16917);
nand U18986 (N_18986,N_16443,N_16805);
xor U18987 (N_18987,N_16631,N_16241);
xnor U18988 (N_18988,N_17081,N_16021);
xnor U18989 (N_18989,N_17148,N_16240);
nand U18990 (N_18990,N_17119,N_16316);
nor U18991 (N_18991,N_17518,N_17507);
and U18992 (N_18992,N_16328,N_17853);
nand U18993 (N_18993,N_17023,N_17304);
or U18994 (N_18994,N_16335,N_17764);
xnor U18995 (N_18995,N_17022,N_17967);
nand U18996 (N_18996,N_16860,N_16588);
xnor U18997 (N_18997,N_16528,N_17307);
or U18998 (N_18998,N_17114,N_17281);
xnor U18999 (N_18999,N_16912,N_16136);
xor U19000 (N_19000,N_17573,N_16600);
nor U19001 (N_19001,N_17006,N_17977);
nor U19002 (N_19002,N_16335,N_17887);
and U19003 (N_19003,N_17852,N_16136);
xor U19004 (N_19004,N_16896,N_17574);
or U19005 (N_19005,N_16717,N_17720);
or U19006 (N_19006,N_17456,N_16444);
nor U19007 (N_19007,N_17295,N_16482);
nand U19008 (N_19008,N_17921,N_17654);
xnor U19009 (N_19009,N_16709,N_17255);
xnor U19010 (N_19010,N_16473,N_16289);
or U19011 (N_19011,N_16030,N_17528);
nor U19012 (N_19012,N_17159,N_17497);
nand U19013 (N_19013,N_17283,N_16504);
nor U19014 (N_19014,N_16174,N_16072);
xor U19015 (N_19015,N_16979,N_17214);
xnor U19016 (N_19016,N_17404,N_17763);
nor U19017 (N_19017,N_17713,N_16305);
or U19018 (N_19018,N_17768,N_17784);
xor U19019 (N_19019,N_17003,N_16690);
nor U19020 (N_19020,N_17956,N_17892);
and U19021 (N_19021,N_17808,N_16989);
or U19022 (N_19022,N_16560,N_17720);
and U19023 (N_19023,N_16176,N_17487);
and U19024 (N_19024,N_17004,N_17649);
xor U19025 (N_19025,N_17487,N_16908);
xor U19026 (N_19026,N_17281,N_17747);
nor U19027 (N_19027,N_17627,N_16427);
and U19028 (N_19028,N_17562,N_17005);
xnor U19029 (N_19029,N_17100,N_17002);
nand U19030 (N_19030,N_16087,N_16175);
nand U19031 (N_19031,N_17821,N_16463);
nand U19032 (N_19032,N_16124,N_16428);
and U19033 (N_19033,N_16998,N_16025);
or U19034 (N_19034,N_17597,N_16312);
and U19035 (N_19035,N_16969,N_17164);
and U19036 (N_19036,N_16343,N_16712);
and U19037 (N_19037,N_17445,N_16045);
xnor U19038 (N_19038,N_17838,N_16769);
nand U19039 (N_19039,N_17009,N_17114);
or U19040 (N_19040,N_17734,N_16297);
nand U19041 (N_19041,N_16890,N_16096);
and U19042 (N_19042,N_16829,N_17770);
or U19043 (N_19043,N_16505,N_17876);
nor U19044 (N_19044,N_16727,N_17807);
nand U19045 (N_19045,N_17819,N_17912);
xnor U19046 (N_19046,N_16040,N_17895);
nand U19047 (N_19047,N_17700,N_17089);
nand U19048 (N_19048,N_17165,N_17112);
nand U19049 (N_19049,N_17088,N_16352);
and U19050 (N_19050,N_17780,N_16452);
or U19051 (N_19051,N_16290,N_17162);
xor U19052 (N_19052,N_16337,N_17240);
and U19053 (N_19053,N_17349,N_16613);
xor U19054 (N_19054,N_16341,N_17363);
xnor U19055 (N_19055,N_16648,N_16091);
or U19056 (N_19056,N_16102,N_16223);
and U19057 (N_19057,N_16002,N_17699);
and U19058 (N_19058,N_17369,N_16459);
nand U19059 (N_19059,N_16626,N_16263);
xnor U19060 (N_19060,N_16979,N_16402);
or U19061 (N_19061,N_17319,N_17361);
or U19062 (N_19062,N_17684,N_16765);
xnor U19063 (N_19063,N_17566,N_17247);
or U19064 (N_19064,N_17798,N_16866);
xnor U19065 (N_19065,N_17889,N_16515);
nor U19066 (N_19066,N_16990,N_17845);
or U19067 (N_19067,N_16025,N_17667);
or U19068 (N_19068,N_17997,N_16363);
nand U19069 (N_19069,N_16490,N_17759);
nor U19070 (N_19070,N_16187,N_17002);
and U19071 (N_19071,N_17958,N_17290);
or U19072 (N_19072,N_16511,N_17400);
and U19073 (N_19073,N_16152,N_16478);
nor U19074 (N_19074,N_17658,N_16112);
and U19075 (N_19075,N_17809,N_16981);
and U19076 (N_19076,N_16853,N_16738);
or U19077 (N_19077,N_16392,N_17511);
xor U19078 (N_19078,N_16893,N_16652);
xor U19079 (N_19079,N_17643,N_16021);
or U19080 (N_19080,N_17681,N_17112);
nand U19081 (N_19081,N_17527,N_16084);
nor U19082 (N_19082,N_17240,N_16348);
xnor U19083 (N_19083,N_17036,N_16233);
xnor U19084 (N_19084,N_17974,N_17312);
xor U19085 (N_19085,N_17084,N_16222);
and U19086 (N_19086,N_16779,N_16004);
xnor U19087 (N_19087,N_17887,N_16010);
nand U19088 (N_19088,N_17910,N_16725);
nand U19089 (N_19089,N_16010,N_16722);
or U19090 (N_19090,N_16664,N_17427);
nand U19091 (N_19091,N_16716,N_16180);
nand U19092 (N_19092,N_16734,N_16830);
and U19093 (N_19093,N_16276,N_17217);
and U19094 (N_19094,N_17763,N_16276);
and U19095 (N_19095,N_16579,N_16611);
nand U19096 (N_19096,N_16015,N_16745);
and U19097 (N_19097,N_16676,N_16081);
and U19098 (N_19098,N_16637,N_16513);
or U19099 (N_19099,N_16312,N_16435);
nand U19100 (N_19100,N_17355,N_17108);
nand U19101 (N_19101,N_16173,N_17219);
nor U19102 (N_19102,N_16664,N_17992);
nand U19103 (N_19103,N_17800,N_16889);
xor U19104 (N_19104,N_16998,N_16535);
xnor U19105 (N_19105,N_17440,N_17566);
and U19106 (N_19106,N_17898,N_17308);
xor U19107 (N_19107,N_16815,N_16087);
or U19108 (N_19108,N_17387,N_17092);
xor U19109 (N_19109,N_16511,N_17273);
xor U19110 (N_19110,N_17372,N_16491);
or U19111 (N_19111,N_16498,N_17890);
or U19112 (N_19112,N_17999,N_17034);
or U19113 (N_19113,N_17980,N_17688);
nand U19114 (N_19114,N_17581,N_17872);
and U19115 (N_19115,N_17293,N_16980);
nor U19116 (N_19116,N_16340,N_17706);
and U19117 (N_19117,N_17710,N_16788);
or U19118 (N_19118,N_16777,N_16663);
nand U19119 (N_19119,N_17784,N_17648);
or U19120 (N_19120,N_17877,N_16462);
and U19121 (N_19121,N_16315,N_17458);
nand U19122 (N_19122,N_16106,N_17949);
xor U19123 (N_19123,N_16403,N_16296);
or U19124 (N_19124,N_16307,N_17017);
and U19125 (N_19125,N_16551,N_16439);
xor U19126 (N_19126,N_17617,N_16602);
and U19127 (N_19127,N_17465,N_16749);
xnor U19128 (N_19128,N_16110,N_16199);
and U19129 (N_19129,N_16182,N_16302);
and U19130 (N_19130,N_17894,N_17958);
or U19131 (N_19131,N_17816,N_17421);
nand U19132 (N_19132,N_16222,N_16859);
xor U19133 (N_19133,N_16594,N_17335);
or U19134 (N_19134,N_16494,N_16608);
nor U19135 (N_19135,N_16721,N_16517);
and U19136 (N_19136,N_17584,N_16435);
nand U19137 (N_19137,N_16230,N_17526);
xnor U19138 (N_19138,N_16628,N_16475);
or U19139 (N_19139,N_16735,N_16492);
and U19140 (N_19140,N_16668,N_17567);
nor U19141 (N_19141,N_17830,N_16666);
or U19142 (N_19142,N_16888,N_17879);
nand U19143 (N_19143,N_17333,N_16150);
xnor U19144 (N_19144,N_17880,N_16623);
nor U19145 (N_19145,N_16730,N_17325);
and U19146 (N_19146,N_16429,N_17220);
and U19147 (N_19147,N_16831,N_16601);
nand U19148 (N_19148,N_16037,N_17158);
nor U19149 (N_19149,N_17186,N_17708);
or U19150 (N_19150,N_16863,N_17917);
xor U19151 (N_19151,N_17943,N_16168);
xnor U19152 (N_19152,N_16843,N_16412);
and U19153 (N_19153,N_17268,N_16176);
nand U19154 (N_19154,N_17776,N_17620);
and U19155 (N_19155,N_17755,N_17437);
or U19156 (N_19156,N_16491,N_17738);
nand U19157 (N_19157,N_16997,N_16837);
or U19158 (N_19158,N_17201,N_17866);
xor U19159 (N_19159,N_16713,N_16756);
nor U19160 (N_19160,N_17720,N_16515);
xor U19161 (N_19161,N_17546,N_17609);
xor U19162 (N_19162,N_17420,N_17767);
or U19163 (N_19163,N_16968,N_17234);
xnor U19164 (N_19164,N_17608,N_17432);
nand U19165 (N_19165,N_16923,N_17535);
nand U19166 (N_19166,N_16986,N_17310);
nor U19167 (N_19167,N_17590,N_16881);
nor U19168 (N_19168,N_16247,N_17992);
and U19169 (N_19169,N_17114,N_16674);
and U19170 (N_19170,N_16436,N_16277);
xnor U19171 (N_19171,N_17614,N_17023);
xnor U19172 (N_19172,N_17306,N_16596);
xnor U19173 (N_19173,N_16777,N_17378);
nand U19174 (N_19174,N_17642,N_16030);
nor U19175 (N_19175,N_16358,N_16720);
and U19176 (N_19176,N_16413,N_17341);
xor U19177 (N_19177,N_16986,N_16724);
nor U19178 (N_19178,N_16354,N_17993);
nand U19179 (N_19179,N_16530,N_16159);
or U19180 (N_19180,N_16884,N_16001);
and U19181 (N_19181,N_16386,N_16533);
nand U19182 (N_19182,N_17519,N_16108);
or U19183 (N_19183,N_17776,N_16750);
nor U19184 (N_19184,N_16770,N_16633);
or U19185 (N_19185,N_16214,N_16377);
xnor U19186 (N_19186,N_16910,N_17524);
nor U19187 (N_19187,N_16005,N_16321);
nor U19188 (N_19188,N_17579,N_16011);
xnor U19189 (N_19189,N_17414,N_16928);
or U19190 (N_19190,N_16192,N_17312);
nand U19191 (N_19191,N_17048,N_17432);
xnor U19192 (N_19192,N_16535,N_16303);
or U19193 (N_19193,N_17273,N_17634);
xor U19194 (N_19194,N_16949,N_17867);
xnor U19195 (N_19195,N_16660,N_17218);
and U19196 (N_19196,N_17571,N_17648);
or U19197 (N_19197,N_16868,N_16299);
or U19198 (N_19198,N_17355,N_16858);
nor U19199 (N_19199,N_17391,N_17205);
nand U19200 (N_19200,N_16387,N_17981);
and U19201 (N_19201,N_16384,N_17825);
and U19202 (N_19202,N_16413,N_17856);
nand U19203 (N_19203,N_17558,N_17117);
xor U19204 (N_19204,N_16872,N_17929);
and U19205 (N_19205,N_16246,N_16568);
nor U19206 (N_19206,N_17457,N_16282);
nand U19207 (N_19207,N_17962,N_16240);
xnor U19208 (N_19208,N_16392,N_17588);
xor U19209 (N_19209,N_17256,N_17560);
nor U19210 (N_19210,N_16615,N_16110);
or U19211 (N_19211,N_16224,N_17842);
xnor U19212 (N_19212,N_16818,N_17164);
and U19213 (N_19213,N_17322,N_16832);
and U19214 (N_19214,N_16556,N_17112);
xnor U19215 (N_19215,N_17356,N_16544);
nand U19216 (N_19216,N_16375,N_16483);
nor U19217 (N_19217,N_17556,N_16424);
and U19218 (N_19218,N_17391,N_17591);
xnor U19219 (N_19219,N_17686,N_16010);
xor U19220 (N_19220,N_17596,N_17609);
or U19221 (N_19221,N_17012,N_17382);
and U19222 (N_19222,N_16789,N_17593);
or U19223 (N_19223,N_17594,N_16038);
or U19224 (N_19224,N_16307,N_16054);
nor U19225 (N_19225,N_17637,N_17156);
nand U19226 (N_19226,N_16974,N_16045);
xor U19227 (N_19227,N_16735,N_17544);
nand U19228 (N_19228,N_16055,N_16729);
nand U19229 (N_19229,N_16078,N_17239);
and U19230 (N_19230,N_17713,N_17112);
nor U19231 (N_19231,N_17351,N_16789);
nor U19232 (N_19232,N_16045,N_16783);
nor U19233 (N_19233,N_16421,N_17208);
nand U19234 (N_19234,N_16869,N_16442);
and U19235 (N_19235,N_16290,N_16262);
and U19236 (N_19236,N_16653,N_17687);
nand U19237 (N_19237,N_16198,N_17973);
xor U19238 (N_19238,N_16338,N_17472);
xnor U19239 (N_19239,N_17863,N_16839);
nor U19240 (N_19240,N_16232,N_16008);
or U19241 (N_19241,N_16237,N_17950);
and U19242 (N_19242,N_16786,N_16791);
xor U19243 (N_19243,N_17972,N_17729);
nand U19244 (N_19244,N_17868,N_17327);
nor U19245 (N_19245,N_17912,N_16071);
and U19246 (N_19246,N_17430,N_17948);
and U19247 (N_19247,N_16637,N_16058);
xor U19248 (N_19248,N_16085,N_16920);
and U19249 (N_19249,N_17830,N_16876);
and U19250 (N_19250,N_17812,N_16784);
nor U19251 (N_19251,N_17259,N_17826);
or U19252 (N_19252,N_17679,N_17148);
nor U19253 (N_19253,N_16725,N_17478);
xnor U19254 (N_19254,N_17440,N_16183);
nand U19255 (N_19255,N_16026,N_17573);
nor U19256 (N_19256,N_16682,N_16034);
xor U19257 (N_19257,N_16255,N_17971);
and U19258 (N_19258,N_17816,N_16478);
xor U19259 (N_19259,N_17652,N_17651);
nand U19260 (N_19260,N_17784,N_17578);
xnor U19261 (N_19261,N_16617,N_16214);
xor U19262 (N_19262,N_16310,N_17404);
nor U19263 (N_19263,N_16706,N_16517);
and U19264 (N_19264,N_16095,N_17092);
or U19265 (N_19265,N_17666,N_17982);
nor U19266 (N_19266,N_16313,N_17110);
xnor U19267 (N_19267,N_17221,N_16398);
or U19268 (N_19268,N_16304,N_17643);
nand U19269 (N_19269,N_17086,N_16105);
nor U19270 (N_19270,N_16487,N_16883);
nand U19271 (N_19271,N_17115,N_16356);
xor U19272 (N_19272,N_16071,N_17632);
nor U19273 (N_19273,N_16777,N_16487);
nor U19274 (N_19274,N_17168,N_17199);
nor U19275 (N_19275,N_16756,N_17218);
nor U19276 (N_19276,N_17893,N_16854);
nand U19277 (N_19277,N_16236,N_17380);
and U19278 (N_19278,N_17903,N_16902);
or U19279 (N_19279,N_17219,N_17292);
nand U19280 (N_19280,N_17796,N_17502);
xor U19281 (N_19281,N_16592,N_17309);
and U19282 (N_19282,N_17676,N_16437);
nand U19283 (N_19283,N_17259,N_17747);
nor U19284 (N_19284,N_17570,N_16828);
nor U19285 (N_19285,N_16570,N_17379);
and U19286 (N_19286,N_17408,N_16516);
nand U19287 (N_19287,N_16731,N_16601);
xor U19288 (N_19288,N_16796,N_16453);
xor U19289 (N_19289,N_17331,N_17751);
xnor U19290 (N_19290,N_16041,N_16463);
and U19291 (N_19291,N_17463,N_17395);
or U19292 (N_19292,N_17936,N_16077);
nand U19293 (N_19293,N_17592,N_16487);
nor U19294 (N_19294,N_16970,N_16960);
nor U19295 (N_19295,N_16541,N_17323);
nand U19296 (N_19296,N_17248,N_17364);
or U19297 (N_19297,N_16833,N_17866);
nor U19298 (N_19298,N_17724,N_16130);
nor U19299 (N_19299,N_17997,N_16453);
or U19300 (N_19300,N_16352,N_17386);
or U19301 (N_19301,N_17941,N_16988);
xnor U19302 (N_19302,N_16304,N_16686);
nor U19303 (N_19303,N_16248,N_16238);
and U19304 (N_19304,N_17498,N_16617);
and U19305 (N_19305,N_17706,N_17100);
or U19306 (N_19306,N_17009,N_17388);
xnor U19307 (N_19307,N_17753,N_16992);
and U19308 (N_19308,N_16403,N_17572);
or U19309 (N_19309,N_16010,N_16965);
nor U19310 (N_19310,N_16810,N_16391);
and U19311 (N_19311,N_17834,N_17000);
or U19312 (N_19312,N_17659,N_16525);
nand U19313 (N_19313,N_16317,N_16309);
nor U19314 (N_19314,N_16604,N_17418);
or U19315 (N_19315,N_17347,N_17301);
or U19316 (N_19316,N_17313,N_16149);
nand U19317 (N_19317,N_17613,N_16332);
nand U19318 (N_19318,N_16759,N_16585);
nor U19319 (N_19319,N_17085,N_17467);
nor U19320 (N_19320,N_16733,N_17845);
xnor U19321 (N_19321,N_16581,N_17246);
xnor U19322 (N_19322,N_17640,N_16642);
and U19323 (N_19323,N_16062,N_17538);
nand U19324 (N_19324,N_16942,N_16492);
nor U19325 (N_19325,N_16498,N_17685);
xor U19326 (N_19326,N_16432,N_17725);
or U19327 (N_19327,N_16100,N_16303);
nand U19328 (N_19328,N_17312,N_16162);
nor U19329 (N_19329,N_16076,N_16190);
and U19330 (N_19330,N_16756,N_17459);
nand U19331 (N_19331,N_17030,N_17416);
nand U19332 (N_19332,N_17695,N_17016);
or U19333 (N_19333,N_16318,N_17341);
or U19334 (N_19334,N_17324,N_17218);
nand U19335 (N_19335,N_17187,N_17913);
xor U19336 (N_19336,N_17437,N_17981);
nor U19337 (N_19337,N_16477,N_17353);
xnor U19338 (N_19338,N_17613,N_17195);
and U19339 (N_19339,N_17710,N_17874);
nand U19340 (N_19340,N_17908,N_17353);
nor U19341 (N_19341,N_16323,N_16151);
and U19342 (N_19342,N_17492,N_16377);
and U19343 (N_19343,N_17129,N_16560);
and U19344 (N_19344,N_16083,N_17584);
nor U19345 (N_19345,N_16506,N_17387);
or U19346 (N_19346,N_17961,N_16097);
nand U19347 (N_19347,N_16020,N_16070);
and U19348 (N_19348,N_16662,N_17045);
and U19349 (N_19349,N_17381,N_16677);
or U19350 (N_19350,N_16590,N_17678);
and U19351 (N_19351,N_16971,N_16375);
nor U19352 (N_19352,N_16404,N_16492);
and U19353 (N_19353,N_16542,N_16749);
nand U19354 (N_19354,N_17678,N_16487);
xor U19355 (N_19355,N_17574,N_17196);
nor U19356 (N_19356,N_16488,N_16583);
or U19357 (N_19357,N_17166,N_17887);
nor U19358 (N_19358,N_16307,N_17492);
xor U19359 (N_19359,N_16476,N_17992);
or U19360 (N_19360,N_17212,N_16300);
and U19361 (N_19361,N_17986,N_17579);
nor U19362 (N_19362,N_17924,N_16016);
or U19363 (N_19363,N_16190,N_16384);
nand U19364 (N_19364,N_17767,N_17876);
or U19365 (N_19365,N_17277,N_16529);
and U19366 (N_19366,N_16103,N_16382);
or U19367 (N_19367,N_16926,N_16663);
xor U19368 (N_19368,N_17534,N_16921);
nand U19369 (N_19369,N_17745,N_17502);
nor U19370 (N_19370,N_17206,N_17617);
and U19371 (N_19371,N_17448,N_16032);
xor U19372 (N_19372,N_17732,N_17700);
nor U19373 (N_19373,N_17951,N_16554);
and U19374 (N_19374,N_16120,N_16197);
nand U19375 (N_19375,N_16989,N_16214);
nand U19376 (N_19376,N_16787,N_16793);
nand U19377 (N_19377,N_17420,N_16060);
nor U19378 (N_19378,N_16918,N_17236);
or U19379 (N_19379,N_17519,N_17208);
nand U19380 (N_19380,N_16175,N_16845);
nor U19381 (N_19381,N_17624,N_17875);
nand U19382 (N_19382,N_16237,N_16886);
nand U19383 (N_19383,N_16712,N_17855);
and U19384 (N_19384,N_17050,N_16999);
or U19385 (N_19385,N_17815,N_16113);
and U19386 (N_19386,N_16043,N_17711);
nand U19387 (N_19387,N_16269,N_16317);
and U19388 (N_19388,N_17296,N_16545);
or U19389 (N_19389,N_17301,N_16426);
xnor U19390 (N_19390,N_17783,N_17296);
and U19391 (N_19391,N_17269,N_16738);
nand U19392 (N_19392,N_16258,N_17347);
nor U19393 (N_19393,N_16239,N_17034);
nor U19394 (N_19394,N_16671,N_17716);
nor U19395 (N_19395,N_17317,N_17495);
nor U19396 (N_19396,N_16144,N_17330);
nand U19397 (N_19397,N_17049,N_16783);
nor U19398 (N_19398,N_17585,N_16079);
nor U19399 (N_19399,N_16162,N_17954);
nor U19400 (N_19400,N_16852,N_17780);
or U19401 (N_19401,N_16351,N_16862);
xnor U19402 (N_19402,N_17953,N_16519);
and U19403 (N_19403,N_16240,N_16084);
nor U19404 (N_19404,N_17401,N_16420);
and U19405 (N_19405,N_16930,N_17406);
nor U19406 (N_19406,N_16600,N_16643);
nand U19407 (N_19407,N_17378,N_16387);
or U19408 (N_19408,N_17972,N_16170);
xor U19409 (N_19409,N_17927,N_17031);
nor U19410 (N_19410,N_16019,N_17929);
nand U19411 (N_19411,N_16834,N_16472);
nand U19412 (N_19412,N_17987,N_16286);
and U19413 (N_19413,N_17681,N_17648);
nand U19414 (N_19414,N_17000,N_16665);
nand U19415 (N_19415,N_16460,N_17298);
or U19416 (N_19416,N_16876,N_16830);
and U19417 (N_19417,N_17451,N_17129);
nand U19418 (N_19418,N_17371,N_17759);
or U19419 (N_19419,N_16844,N_16372);
nor U19420 (N_19420,N_17571,N_17887);
nand U19421 (N_19421,N_16512,N_17335);
nand U19422 (N_19422,N_17666,N_17035);
nor U19423 (N_19423,N_17973,N_17307);
nor U19424 (N_19424,N_17883,N_17612);
or U19425 (N_19425,N_16279,N_16275);
and U19426 (N_19426,N_17946,N_17996);
nand U19427 (N_19427,N_17661,N_17307);
nor U19428 (N_19428,N_16840,N_17756);
nand U19429 (N_19429,N_16793,N_17593);
xnor U19430 (N_19430,N_16620,N_16434);
and U19431 (N_19431,N_16831,N_16968);
xor U19432 (N_19432,N_17632,N_16884);
and U19433 (N_19433,N_17424,N_16148);
nand U19434 (N_19434,N_16970,N_17835);
nand U19435 (N_19435,N_16632,N_16434);
xor U19436 (N_19436,N_17429,N_17905);
xnor U19437 (N_19437,N_17152,N_17807);
nand U19438 (N_19438,N_17739,N_17023);
and U19439 (N_19439,N_17610,N_16544);
xnor U19440 (N_19440,N_17056,N_16175);
nand U19441 (N_19441,N_17369,N_17625);
or U19442 (N_19442,N_17880,N_17961);
and U19443 (N_19443,N_16632,N_17555);
or U19444 (N_19444,N_16982,N_16806);
or U19445 (N_19445,N_17778,N_16690);
nand U19446 (N_19446,N_17409,N_17709);
nor U19447 (N_19447,N_17955,N_16043);
xor U19448 (N_19448,N_17435,N_17498);
nor U19449 (N_19449,N_17905,N_16050);
or U19450 (N_19450,N_16078,N_17902);
nand U19451 (N_19451,N_16642,N_16529);
or U19452 (N_19452,N_17532,N_16428);
nor U19453 (N_19453,N_17597,N_17189);
xnor U19454 (N_19454,N_16158,N_17418);
and U19455 (N_19455,N_16103,N_17245);
and U19456 (N_19456,N_17978,N_17910);
nand U19457 (N_19457,N_16532,N_16659);
nand U19458 (N_19458,N_16311,N_17881);
and U19459 (N_19459,N_17849,N_16590);
nand U19460 (N_19460,N_17008,N_16378);
and U19461 (N_19461,N_17448,N_16932);
nand U19462 (N_19462,N_17985,N_16513);
and U19463 (N_19463,N_17009,N_17880);
xor U19464 (N_19464,N_17978,N_16336);
xor U19465 (N_19465,N_17378,N_16228);
xnor U19466 (N_19466,N_16955,N_17724);
and U19467 (N_19467,N_16104,N_17624);
and U19468 (N_19468,N_17983,N_17265);
xnor U19469 (N_19469,N_16423,N_16732);
nor U19470 (N_19470,N_16409,N_16347);
or U19471 (N_19471,N_16242,N_17617);
xnor U19472 (N_19472,N_17131,N_17295);
or U19473 (N_19473,N_17948,N_17861);
nor U19474 (N_19474,N_16816,N_16068);
nor U19475 (N_19475,N_16795,N_17074);
and U19476 (N_19476,N_17253,N_17877);
nor U19477 (N_19477,N_17615,N_16767);
or U19478 (N_19478,N_17645,N_16479);
xnor U19479 (N_19479,N_17048,N_16095);
and U19480 (N_19480,N_17877,N_17659);
xor U19481 (N_19481,N_16853,N_17302);
nand U19482 (N_19482,N_17517,N_17002);
nor U19483 (N_19483,N_16511,N_16681);
or U19484 (N_19484,N_17132,N_17423);
xor U19485 (N_19485,N_16219,N_17886);
nand U19486 (N_19486,N_16835,N_17186);
nand U19487 (N_19487,N_16601,N_17880);
or U19488 (N_19488,N_16367,N_16793);
nor U19489 (N_19489,N_17678,N_16129);
or U19490 (N_19490,N_16454,N_17895);
nor U19491 (N_19491,N_17294,N_17766);
nor U19492 (N_19492,N_16425,N_16654);
xor U19493 (N_19493,N_16577,N_16157);
xnor U19494 (N_19494,N_16399,N_17853);
nor U19495 (N_19495,N_16919,N_17548);
or U19496 (N_19496,N_16314,N_17634);
nand U19497 (N_19497,N_16653,N_16988);
xor U19498 (N_19498,N_16458,N_17258);
or U19499 (N_19499,N_16760,N_16177);
nand U19500 (N_19500,N_16817,N_17438);
and U19501 (N_19501,N_16223,N_16930);
or U19502 (N_19502,N_16732,N_17170);
nand U19503 (N_19503,N_17903,N_17246);
and U19504 (N_19504,N_17136,N_16495);
and U19505 (N_19505,N_16306,N_16948);
xor U19506 (N_19506,N_16850,N_16240);
and U19507 (N_19507,N_16330,N_17711);
and U19508 (N_19508,N_17707,N_17777);
xor U19509 (N_19509,N_16112,N_17933);
or U19510 (N_19510,N_16882,N_17235);
nand U19511 (N_19511,N_16178,N_16496);
xor U19512 (N_19512,N_17811,N_16606);
nor U19513 (N_19513,N_17904,N_16602);
or U19514 (N_19514,N_17951,N_16021);
or U19515 (N_19515,N_17544,N_17629);
nor U19516 (N_19516,N_17015,N_17899);
xor U19517 (N_19517,N_16745,N_16404);
nand U19518 (N_19518,N_16358,N_17628);
nand U19519 (N_19519,N_17099,N_16765);
nand U19520 (N_19520,N_16408,N_17812);
and U19521 (N_19521,N_16396,N_17418);
or U19522 (N_19522,N_16886,N_16570);
nor U19523 (N_19523,N_16171,N_16931);
nand U19524 (N_19524,N_17692,N_17002);
xor U19525 (N_19525,N_17878,N_17093);
or U19526 (N_19526,N_16439,N_16633);
xnor U19527 (N_19527,N_16121,N_16512);
or U19528 (N_19528,N_17702,N_16995);
and U19529 (N_19529,N_16716,N_17361);
nor U19530 (N_19530,N_17561,N_16472);
nand U19531 (N_19531,N_17475,N_16963);
xor U19532 (N_19532,N_17361,N_16794);
nor U19533 (N_19533,N_16793,N_16061);
xor U19534 (N_19534,N_16686,N_16698);
or U19535 (N_19535,N_16231,N_16803);
nand U19536 (N_19536,N_17435,N_17901);
or U19537 (N_19537,N_17161,N_17821);
nor U19538 (N_19538,N_17521,N_17971);
xnor U19539 (N_19539,N_17781,N_16674);
nand U19540 (N_19540,N_16299,N_17708);
and U19541 (N_19541,N_17478,N_16968);
nand U19542 (N_19542,N_17256,N_17455);
nor U19543 (N_19543,N_17230,N_16046);
xnor U19544 (N_19544,N_16988,N_17739);
and U19545 (N_19545,N_17553,N_17310);
nor U19546 (N_19546,N_17340,N_17284);
and U19547 (N_19547,N_17797,N_16433);
nor U19548 (N_19548,N_16734,N_16860);
nand U19549 (N_19549,N_16926,N_16402);
nand U19550 (N_19550,N_16626,N_16801);
xnor U19551 (N_19551,N_16093,N_17004);
or U19552 (N_19552,N_17355,N_16642);
or U19553 (N_19553,N_16844,N_16520);
or U19554 (N_19554,N_16502,N_16023);
nand U19555 (N_19555,N_17560,N_17818);
xnor U19556 (N_19556,N_17617,N_17640);
xnor U19557 (N_19557,N_16409,N_17021);
nor U19558 (N_19558,N_17357,N_17460);
nor U19559 (N_19559,N_17504,N_16242);
or U19560 (N_19560,N_16401,N_16952);
and U19561 (N_19561,N_16241,N_16706);
nand U19562 (N_19562,N_17283,N_16488);
or U19563 (N_19563,N_17638,N_17586);
and U19564 (N_19564,N_16898,N_16622);
and U19565 (N_19565,N_17542,N_17621);
xor U19566 (N_19566,N_17885,N_17621);
xor U19567 (N_19567,N_16276,N_17784);
and U19568 (N_19568,N_17280,N_16429);
and U19569 (N_19569,N_17552,N_17346);
xnor U19570 (N_19570,N_17518,N_16642);
nor U19571 (N_19571,N_16618,N_16135);
or U19572 (N_19572,N_17361,N_17632);
and U19573 (N_19573,N_16143,N_16454);
and U19574 (N_19574,N_17257,N_17513);
nor U19575 (N_19575,N_17461,N_16023);
and U19576 (N_19576,N_17783,N_17941);
nor U19577 (N_19577,N_16239,N_16388);
xor U19578 (N_19578,N_16365,N_17933);
nand U19579 (N_19579,N_17482,N_17970);
or U19580 (N_19580,N_17495,N_16653);
nor U19581 (N_19581,N_16914,N_17096);
xnor U19582 (N_19582,N_16561,N_17046);
and U19583 (N_19583,N_17239,N_16314);
xnor U19584 (N_19584,N_17274,N_16988);
or U19585 (N_19585,N_17032,N_17623);
or U19586 (N_19586,N_16598,N_16565);
or U19587 (N_19587,N_17326,N_17825);
xor U19588 (N_19588,N_17898,N_17648);
xor U19589 (N_19589,N_17787,N_16678);
nor U19590 (N_19590,N_17910,N_17877);
nor U19591 (N_19591,N_16267,N_17951);
nor U19592 (N_19592,N_16094,N_16929);
and U19593 (N_19593,N_16678,N_17977);
nor U19594 (N_19594,N_16969,N_16699);
nand U19595 (N_19595,N_17622,N_16927);
or U19596 (N_19596,N_16784,N_17841);
and U19597 (N_19597,N_16533,N_17486);
nand U19598 (N_19598,N_17995,N_17903);
xnor U19599 (N_19599,N_16719,N_17097);
or U19600 (N_19600,N_17131,N_16208);
nand U19601 (N_19601,N_16550,N_17680);
and U19602 (N_19602,N_16378,N_16132);
nand U19603 (N_19603,N_16395,N_17212);
nand U19604 (N_19604,N_16036,N_16489);
and U19605 (N_19605,N_16067,N_16055);
xor U19606 (N_19606,N_16799,N_17409);
nand U19607 (N_19607,N_17065,N_17929);
and U19608 (N_19608,N_16619,N_16257);
nor U19609 (N_19609,N_17186,N_17596);
and U19610 (N_19610,N_16389,N_17601);
or U19611 (N_19611,N_16431,N_17347);
nand U19612 (N_19612,N_17262,N_16822);
nand U19613 (N_19613,N_16678,N_17412);
xor U19614 (N_19614,N_17358,N_17637);
nor U19615 (N_19615,N_17925,N_16435);
nand U19616 (N_19616,N_16313,N_16962);
nor U19617 (N_19617,N_16201,N_17585);
or U19618 (N_19618,N_16941,N_17130);
nand U19619 (N_19619,N_17663,N_17965);
and U19620 (N_19620,N_17999,N_17523);
nor U19621 (N_19621,N_17930,N_16700);
or U19622 (N_19622,N_16830,N_17189);
nand U19623 (N_19623,N_16158,N_16513);
xor U19624 (N_19624,N_16113,N_16266);
nand U19625 (N_19625,N_16445,N_16874);
or U19626 (N_19626,N_16104,N_16157);
nand U19627 (N_19627,N_17129,N_16067);
nand U19628 (N_19628,N_16772,N_17646);
nand U19629 (N_19629,N_16841,N_17994);
nand U19630 (N_19630,N_17900,N_17362);
or U19631 (N_19631,N_17793,N_16121);
or U19632 (N_19632,N_16688,N_16068);
or U19633 (N_19633,N_16711,N_17512);
nand U19634 (N_19634,N_16163,N_17776);
xor U19635 (N_19635,N_16002,N_17195);
nand U19636 (N_19636,N_16534,N_16605);
xnor U19637 (N_19637,N_16155,N_16863);
and U19638 (N_19638,N_16819,N_17509);
xnor U19639 (N_19639,N_16234,N_17548);
xor U19640 (N_19640,N_16191,N_17719);
xnor U19641 (N_19641,N_16640,N_16793);
nor U19642 (N_19642,N_16942,N_16521);
xor U19643 (N_19643,N_16944,N_16082);
xor U19644 (N_19644,N_17178,N_17959);
nand U19645 (N_19645,N_17399,N_16670);
nor U19646 (N_19646,N_17044,N_16873);
xnor U19647 (N_19647,N_16921,N_16480);
and U19648 (N_19648,N_17330,N_16079);
nand U19649 (N_19649,N_16257,N_17174);
nor U19650 (N_19650,N_16725,N_17282);
or U19651 (N_19651,N_16504,N_17481);
nand U19652 (N_19652,N_16447,N_16621);
or U19653 (N_19653,N_16631,N_17329);
and U19654 (N_19654,N_16588,N_17375);
nand U19655 (N_19655,N_17004,N_17905);
xnor U19656 (N_19656,N_16492,N_16912);
nand U19657 (N_19657,N_17411,N_17796);
xnor U19658 (N_19658,N_17326,N_16657);
nor U19659 (N_19659,N_16564,N_17960);
nand U19660 (N_19660,N_16372,N_16885);
and U19661 (N_19661,N_16288,N_16926);
nand U19662 (N_19662,N_16848,N_17777);
nand U19663 (N_19663,N_16273,N_16731);
or U19664 (N_19664,N_17117,N_16951);
nand U19665 (N_19665,N_16397,N_17316);
and U19666 (N_19666,N_16692,N_16207);
xnor U19667 (N_19667,N_16638,N_16439);
xnor U19668 (N_19668,N_17782,N_16097);
or U19669 (N_19669,N_17739,N_17178);
and U19670 (N_19670,N_16084,N_17321);
nand U19671 (N_19671,N_16931,N_16839);
xor U19672 (N_19672,N_16481,N_16676);
nor U19673 (N_19673,N_16088,N_16889);
nand U19674 (N_19674,N_16220,N_16862);
and U19675 (N_19675,N_17079,N_16893);
xnor U19676 (N_19676,N_16044,N_16171);
and U19677 (N_19677,N_16228,N_17518);
or U19678 (N_19678,N_16677,N_17501);
nor U19679 (N_19679,N_16504,N_17931);
nand U19680 (N_19680,N_17660,N_16600);
nor U19681 (N_19681,N_17517,N_16574);
and U19682 (N_19682,N_16347,N_16962);
xnor U19683 (N_19683,N_17182,N_17103);
nand U19684 (N_19684,N_17994,N_17345);
xnor U19685 (N_19685,N_16720,N_16294);
xor U19686 (N_19686,N_16184,N_17273);
or U19687 (N_19687,N_17009,N_17795);
nor U19688 (N_19688,N_16373,N_16138);
and U19689 (N_19689,N_17721,N_16902);
nand U19690 (N_19690,N_17632,N_16657);
xnor U19691 (N_19691,N_16689,N_17667);
nor U19692 (N_19692,N_17804,N_17385);
xor U19693 (N_19693,N_16209,N_16886);
nand U19694 (N_19694,N_16010,N_17631);
xor U19695 (N_19695,N_16679,N_16080);
or U19696 (N_19696,N_17123,N_17740);
or U19697 (N_19697,N_17078,N_17858);
nand U19698 (N_19698,N_16725,N_17737);
or U19699 (N_19699,N_16760,N_16814);
or U19700 (N_19700,N_17634,N_16987);
or U19701 (N_19701,N_16613,N_17301);
xor U19702 (N_19702,N_17223,N_17196);
nor U19703 (N_19703,N_16568,N_17430);
nand U19704 (N_19704,N_16542,N_16496);
or U19705 (N_19705,N_17826,N_16803);
xor U19706 (N_19706,N_17450,N_17179);
nand U19707 (N_19707,N_16675,N_17521);
or U19708 (N_19708,N_16905,N_16877);
nand U19709 (N_19709,N_17907,N_16584);
and U19710 (N_19710,N_17493,N_17446);
and U19711 (N_19711,N_16663,N_16341);
or U19712 (N_19712,N_16361,N_16429);
xor U19713 (N_19713,N_16267,N_17102);
nand U19714 (N_19714,N_17931,N_17475);
and U19715 (N_19715,N_17825,N_16570);
and U19716 (N_19716,N_16351,N_16381);
nand U19717 (N_19717,N_17923,N_16574);
or U19718 (N_19718,N_17886,N_17869);
and U19719 (N_19719,N_16450,N_16194);
or U19720 (N_19720,N_16512,N_17580);
nand U19721 (N_19721,N_16762,N_16117);
nand U19722 (N_19722,N_17751,N_17540);
and U19723 (N_19723,N_16307,N_17511);
or U19724 (N_19724,N_17066,N_17683);
nor U19725 (N_19725,N_16570,N_17294);
or U19726 (N_19726,N_17134,N_17384);
xnor U19727 (N_19727,N_17478,N_17452);
and U19728 (N_19728,N_16532,N_16405);
xnor U19729 (N_19729,N_16069,N_16444);
nand U19730 (N_19730,N_17536,N_17565);
nor U19731 (N_19731,N_17988,N_17779);
and U19732 (N_19732,N_17232,N_16076);
and U19733 (N_19733,N_17009,N_16625);
or U19734 (N_19734,N_16806,N_17947);
nor U19735 (N_19735,N_16145,N_17125);
nand U19736 (N_19736,N_17111,N_16118);
nor U19737 (N_19737,N_17348,N_17620);
nor U19738 (N_19738,N_17362,N_16700);
or U19739 (N_19739,N_16278,N_17452);
or U19740 (N_19740,N_17025,N_16158);
nor U19741 (N_19741,N_17848,N_17357);
nor U19742 (N_19742,N_17557,N_16862);
nand U19743 (N_19743,N_17847,N_17584);
or U19744 (N_19744,N_16641,N_16266);
nand U19745 (N_19745,N_17586,N_17433);
or U19746 (N_19746,N_17591,N_16168);
xor U19747 (N_19747,N_16856,N_16918);
nor U19748 (N_19748,N_17218,N_17712);
nor U19749 (N_19749,N_16846,N_16712);
nand U19750 (N_19750,N_17995,N_16824);
and U19751 (N_19751,N_16420,N_16238);
nand U19752 (N_19752,N_17117,N_16646);
nor U19753 (N_19753,N_16923,N_17791);
nor U19754 (N_19754,N_17504,N_16888);
nand U19755 (N_19755,N_16370,N_17684);
and U19756 (N_19756,N_16835,N_16168);
nor U19757 (N_19757,N_16110,N_17619);
nor U19758 (N_19758,N_16456,N_16028);
xor U19759 (N_19759,N_16455,N_17412);
xnor U19760 (N_19760,N_16894,N_17795);
xor U19761 (N_19761,N_16898,N_17607);
and U19762 (N_19762,N_16088,N_17622);
or U19763 (N_19763,N_17258,N_17734);
and U19764 (N_19764,N_16020,N_16442);
or U19765 (N_19765,N_17781,N_16292);
xnor U19766 (N_19766,N_16487,N_16555);
or U19767 (N_19767,N_17204,N_16821);
and U19768 (N_19768,N_17558,N_17033);
xnor U19769 (N_19769,N_17272,N_16995);
or U19770 (N_19770,N_16870,N_16367);
and U19771 (N_19771,N_16212,N_17933);
nand U19772 (N_19772,N_16456,N_17648);
xor U19773 (N_19773,N_16652,N_16434);
xnor U19774 (N_19774,N_17905,N_17637);
or U19775 (N_19775,N_16802,N_16196);
nand U19776 (N_19776,N_16916,N_17004);
and U19777 (N_19777,N_16044,N_16861);
nor U19778 (N_19778,N_17029,N_17889);
and U19779 (N_19779,N_16789,N_17520);
or U19780 (N_19780,N_17754,N_16564);
or U19781 (N_19781,N_17513,N_16564);
nand U19782 (N_19782,N_17402,N_17550);
nor U19783 (N_19783,N_16120,N_16365);
and U19784 (N_19784,N_16371,N_16450);
and U19785 (N_19785,N_16664,N_17260);
and U19786 (N_19786,N_17695,N_17416);
nor U19787 (N_19787,N_16737,N_16220);
or U19788 (N_19788,N_17529,N_17546);
nor U19789 (N_19789,N_17541,N_16147);
and U19790 (N_19790,N_16473,N_17703);
nand U19791 (N_19791,N_16595,N_16184);
or U19792 (N_19792,N_16207,N_16434);
nand U19793 (N_19793,N_16335,N_17992);
nand U19794 (N_19794,N_17527,N_16242);
xor U19795 (N_19795,N_17302,N_16174);
or U19796 (N_19796,N_17413,N_17202);
or U19797 (N_19797,N_17003,N_17284);
nor U19798 (N_19798,N_16405,N_16004);
nor U19799 (N_19799,N_17768,N_17056);
nor U19800 (N_19800,N_17092,N_16306);
or U19801 (N_19801,N_17079,N_16766);
or U19802 (N_19802,N_17610,N_17515);
xnor U19803 (N_19803,N_17431,N_17672);
nor U19804 (N_19804,N_16516,N_16172);
xnor U19805 (N_19805,N_17337,N_17237);
or U19806 (N_19806,N_16812,N_16980);
xor U19807 (N_19807,N_17338,N_17646);
and U19808 (N_19808,N_16673,N_16550);
and U19809 (N_19809,N_17783,N_16135);
and U19810 (N_19810,N_16684,N_17202);
nand U19811 (N_19811,N_16356,N_17809);
nand U19812 (N_19812,N_17336,N_17027);
xnor U19813 (N_19813,N_17366,N_16847);
and U19814 (N_19814,N_16559,N_17528);
nand U19815 (N_19815,N_17480,N_16312);
and U19816 (N_19816,N_17451,N_16672);
nor U19817 (N_19817,N_16366,N_17759);
nand U19818 (N_19818,N_17917,N_16036);
xnor U19819 (N_19819,N_16972,N_17623);
xor U19820 (N_19820,N_17732,N_16625);
nor U19821 (N_19821,N_16769,N_16310);
nand U19822 (N_19822,N_17390,N_16111);
nand U19823 (N_19823,N_16841,N_16465);
nand U19824 (N_19824,N_17148,N_16807);
nor U19825 (N_19825,N_16091,N_16972);
nor U19826 (N_19826,N_17022,N_16329);
nand U19827 (N_19827,N_16497,N_17419);
or U19828 (N_19828,N_17459,N_17358);
nand U19829 (N_19829,N_17955,N_17724);
nand U19830 (N_19830,N_16033,N_17156);
xnor U19831 (N_19831,N_16139,N_17596);
and U19832 (N_19832,N_17267,N_16577);
nor U19833 (N_19833,N_17763,N_16244);
nor U19834 (N_19834,N_17938,N_17875);
and U19835 (N_19835,N_17002,N_16752);
nor U19836 (N_19836,N_17054,N_17132);
xnor U19837 (N_19837,N_16808,N_17100);
xor U19838 (N_19838,N_17713,N_16728);
xnor U19839 (N_19839,N_16378,N_16410);
nor U19840 (N_19840,N_16720,N_17056);
nand U19841 (N_19841,N_16292,N_17989);
nor U19842 (N_19842,N_16862,N_16679);
xor U19843 (N_19843,N_16194,N_16158);
xnor U19844 (N_19844,N_16126,N_16642);
or U19845 (N_19845,N_17384,N_16204);
and U19846 (N_19846,N_17782,N_17943);
or U19847 (N_19847,N_16176,N_16071);
nor U19848 (N_19848,N_16526,N_16797);
nor U19849 (N_19849,N_16915,N_16548);
or U19850 (N_19850,N_16746,N_17813);
or U19851 (N_19851,N_16512,N_16189);
nor U19852 (N_19852,N_16568,N_16937);
nand U19853 (N_19853,N_17532,N_16558);
nand U19854 (N_19854,N_16320,N_17092);
nor U19855 (N_19855,N_16595,N_17070);
nor U19856 (N_19856,N_17790,N_17851);
and U19857 (N_19857,N_17861,N_16612);
xnor U19858 (N_19858,N_16051,N_17423);
xnor U19859 (N_19859,N_17773,N_17431);
nand U19860 (N_19860,N_16353,N_17214);
xor U19861 (N_19861,N_16193,N_17173);
or U19862 (N_19862,N_16933,N_16967);
nor U19863 (N_19863,N_16583,N_17189);
and U19864 (N_19864,N_17562,N_17241);
or U19865 (N_19865,N_16279,N_16241);
nor U19866 (N_19866,N_17760,N_16982);
xor U19867 (N_19867,N_17122,N_17021);
or U19868 (N_19868,N_17037,N_16967);
or U19869 (N_19869,N_17101,N_16486);
xnor U19870 (N_19870,N_17147,N_17813);
or U19871 (N_19871,N_16367,N_17422);
nand U19872 (N_19872,N_17041,N_17288);
xor U19873 (N_19873,N_17751,N_17651);
and U19874 (N_19874,N_16893,N_16486);
xnor U19875 (N_19875,N_16177,N_16657);
and U19876 (N_19876,N_17128,N_17262);
or U19877 (N_19877,N_16122,N_16242);
nor U19878 (N_19878,N_17318,N_17162);
and U19879 (N_19879,N_16443,N_16826);
xnor U19880 (N_19880,N_16773,N_16703);
and U19881 (N_19881,N_17352,N_17909);
xnor U19882 (N_19882,N_16980,N_16899);
nor U19883 (N_19883,N_17542,N_16128);
nand U19884 (N_19884,N_17089,N_16925);
nor U19885 (N_19885,N_17113,N_16983);
nand U19886 (N_19886,N_16215,N_16866);
or U19887 (N_19887,N_16789,N_17062);
nor U19888 (N_19888,N_17938,N_17695);
nand U19889 (N_19889,N_16604,N_16817);
nor U19890 (N_19890,N_16674,N_16359);
nor U19891 (N_19891,N_16714,N_17583);
or U19892 (N_19892,N_17620,N_17397);
and U19893 (N_19893,N_16020,N_17735);
and U19894 (N_19894,N_16030,N_16716);
nand U19895 (N_19895,N_16761,N_16036);
nand U19896 (N_19896,N_17680,N_16866);
nor U19897 (N_19897,N_16555,N_16653);
nand U19898 (N_19898,N_16144,N_16680);
nor U19899 (N_19899,N_17420,N_16981);
nor U19900 (N_19900,N_16728,N_17358);
nand U19901 (N_19901,N_17150,N_16581);
xor U19902 (N_19902,N_16850,N_16588);
or U19903 (N_19903,N_17375,N_17469);
xor U19904 (N_19904,N_16624,N_16083);
nand U19905 (N_19905,N_17816,N_17967);
nor U19906 (N_19906,N_17984,N_16627);
or U19907 (N_19907,N_16739,N_17183);
or U19908 (N_19908,N_17367,N_16124);
xnor U19909 (N_19909,N_16147,N_17726);
xnor U19910 (N_19910,N_16317,N_16824);
or U19911 (N_19911,N_17163,N_17367);
nor U19912 (N_19912,N_16341,N_16352);
nor U19913 (N_19913,N_17271,N_16815);
or U19914 (N_19914,N_17973,N_17288);
nor U19915 (N_19915,N_17945,N_17627);
or U19916 (N_19916,N_16715,N_16776);
nor U19917 (N_19917,N_16598,N_17855);
and U19918 (N_19918,N_17916,N_16190);
and U19919 (N_19919,N_17582,N_17415);
nand U19920 (N_19920,N_16417,N_16634);
nand U19921 (N_19921,N_17749,N_17398);
nor U19922 (N_19922,N_17522,N_16370);
nand U19923 (N_19923,N_17723,N_17201);
xnor U19924 (N_19924,N_16765,N_17365);
xor U19925 (N_19925,N_16276,N_16565);
nor U19926 (N_19926,N_17312,N_16578);
and U19927 (N_19927,N_17706,N_17911);
nor U19928 (N_19928,N_16335,N_16569);
and U19929 (N_19929,N_16700,N_17058);
and U19930 (N_19930,N_17339,N_17351);
or U19931 (N_19931,N_16426,N_16850);
nor U19932 (N_19932,N_17419,N_16492);
xor U19933 (N_19933,N_17239,N_17449);
xor U19934 (N_19934,N_17686,N_16992);
xnor U19935 (N_19935,N_17842,N_16887);
xor U19936 (N_19936,N_17979,N_16122);
or U19937 (N_19937,N_17889,N_17930);
and U19938 (N_19938,N_17374,N_16938);
and U19939 (N_19939,N_17756,N_17985);
nor U19940 (N_19940,N_16479,N_16770);
nand U19941 (N_19941,N_16570,N_17290);
nor U19942 (N_19942,N_17955,N_16685);
nand U19943 (N_19943,N_17524,N_16562);
nor U19944 (N_19944,N_17974,N_17633);
nor U19945 (N_19945,N_17888,N_17611);
nor U19946 (N_19946,N_17628,N_16929);
nand U19947 (N_19947,N_17482,N_16325);
nor U19948 (N_19948,N_16495,N_17286);
or U19949 (N_19949,N_16157,N_17200);
nor U19950 (N_19950,N_17366,N_16533);
and U19951 (N_19951,N_16602,N_16094);
and U19952 (N_19952,N_17261,N_16378);
or U19953 (N_19953,N_16063,N_17374);
xor U19954 (N_19954,N_16497,N_16623);
nor U19955 (N_19955,N_16482,N_17385);
xnor U19956 (N_19956,N_16082,N_16982);
xor U19957 (N_19957,N_16990,N_16491);
or U19958 (N_19958,N_16404,N_17985);
xor U19959 (N_19959,N_16145,N_17327);
and U19960 (N_19960,N_17432,N_17931);
and U19961 (N_19961,N_16295,N_17119);
nand U19962 (N_19962,N_17448,N_16986);
nand U19963 (N_19963,N_16179,N_16005);
xnor U19964 (N_19964,N_17036,N_17805);
xnor U19965 (N_19965,N_17316,N_16813);
nor U19966 (N_19966,N_16078,N_16385);
or U19967 (N_19967,N_17001,N_17073);
nand U19968 (N_19968,N_17868,N_16322);
nor U19969 (N_19969,N_17977,N_16937);
nor U19970 (N_19970,N_16956,N_16115);
nor U19971 (N_19971,N_17826,N_16439);
nand U19972 (N_19972,N_16851,N_17439);
or U19973 (N_19973,N_16929,N_16082);
or U19974 (N_19974,N_16760,N_17914);
nor U19975 (N_19975,N_16050,N_16775);
nand U19976 (N_19976,N_17915,N_17181);
and U19977 (N_19977,N_17178,N_16084);
or U19978 (N_19978,N_17252,N_17025);
nor U19979 (N_19979,N_16585,N_17222);
nand U19980 (N_19980,N_16053,N_17835);
and U19981 (N_19981,N_17187,N_16772);
or U19982 (N_19982,N_17998,N_17962);
and U19983 (N_19983,N_16600,N_17632);
xnor U19984 (N_19984,N_17470,N_16481);
nor U19985 (N_19985,N_16050,N_16942);
xor U19986 (N_19986,N_17062,N_16309);
or U19987 (N_19987,N_16998,N_17494);
nand U19988 (N_19988,N_17443,N_17442);
or U19989 (N_19989,N_17147,N_17535);
nand U19990 (N_19990,N_16902,N_17658);
xnor U19991 (N_19991,N_16507,N_17978);
or U19992 (N_19992,N_16445,N_16988);
or U19993 (N_19993,N_16947,N_16919);
nand U19994 (N_19994,N_16810,N_16928);
nand U19995 (N_19995,N_16464,N_16083);
xor U19996 (N_19996,N_16468,N_17448);
and U19997 (N_19997,N_16709,N_17799);
nand U19998 (N_19998,N_16820,N_16856);
nand U19999 (N_19999,N_17192,N_17886);
nor U20000 (N_20000,N_18864,N_19893);
nand U20001 (N_20001,N_19763,N_19014);
nor U20002 (N_20002,N_19814,N_19576);
and U20003 (N_20003,N_18300,N_19647);
and U20004 (N_20004,N_18564,N_18678);
nand U20005 (N_20005,N_19206,N_18157);
nor U20006 (N_20006,N_19102,N_19913);
nor U20007 (N_20007,N_18266,N_19676);
xnor U20008 (N_20008,N_19830,N_18277);
xor U20009 (N_20009,N_19300,N_18137);
xnor U20010 (N_20010,N_19453,N_19817);
or U20011 (N_20011,N_19820,N_19862);
xnor U20012 (N_20012,N_18194,N_19500);
nand U20013 (N_20013,N_19897,N_19973);
and U20014 (N_20014,N_19509,N_19867);
nand U20015 (N_20015,N_19538,N_19465);
or U20016 (N_20016,N_18548,N_18090);
nor U20017 (N_20017,N_19038,N_18134);
nand U20018 (N_20018,N_18087,N_19727);
nor U20019 (N_20019,N_18707,N_18073);
or U20020 (N_20020,N_19164,N_18369);
xor U20021 (N_20021,N_18254,N_19156);
nand U20022 (N_20022,N_19725,N_19902);
nor U20023 (N_20023,N_18753,N_19226);
nor U20024 (N_20024,N_18488,N_19593);
nand U20025 (N_20025,N_18291,N_19209);
or U20026 (N_20026,N_18023,N_19436);
nand U20027 (N_20027,N_19493,N_18511);
xor U20028 (N_20028,N_18167,N_19578);
nor U20029 (N_20029,N_18032,N_19764);
or U20030 (N_20030,N_19675,N_18855);
nor U20031 (N_20031,N_18240,N_18725);
nand U20032 (N_20032,N_18734,N_19229);
xnor U20033 (N_20033,N_18785,N_19648);
and U20034 (N_20034,N_19200,N_19146);
or U20035 (N_20035,N_18402,N_18242);
nand U20036 (N_20036,N_19715,N_19400);
nand U20037 (N_20037,N_19688,N_19846);
nor U20038 (N_20038,N_19819,N_19935);
xnor U20039 (N_20039,N_19245,N_19418);
nor U20040 (N_20040,N_18462,N_18482);
nand U20041 (N_20041,N_18279,N_18133);
and U20042 (N_20042,N_18691,N_18780);
xor U20043 (N_20043,N_19505,N_18265);
xor U20044 (N_20044,N_18986,N_18508);
and U20045 (N_20045,N_18378,N_18628);
and U20046 (N_20046,N_19193,N_19099);
xnor U20047 (N_20047,N_19656,N_18316);
xnor U20048 (N_20048,N_19246,N_19285);
or U20049 (N_20049,N_18318,N_18064);
or U20050 (N_20050,N_19546,N_18322);
nor U20051 (N_20051,N_19704,N_18208);
xnor U20052 (N_20052,N_19249,N_19842);
or U20053 (N_20053,N_18321,N_19395);
nor U20054 (N_20054,N_19079,N_18372);
xor U20055 (N_20055,N_19690,N_18390);
and U20056 (N_20056,N_18722,N_19889);
nor U20057 (N_20057,N_19440,N_19225);
nand U20058 (N_20058,N_19899,N_19350);
xnor U20059 (N_20059,N_18455,N_19901);
and U20060 (N_20060,N_18703,N_18682);
xor U20061 (N_20061,N_18450,N_19622);
and U20062 (N_20062,N_18699,N_19398);
nand U20063 (N_20063,N_18719,N_18483);
nor U20064 (N_20064,N_18051,N_18422);
xor U20065 (N_20065,N_18163,N_19197);
nand U20066 (N_20066,N_19363,N_19953);
or U20067 (N_20067,N_19255,N_18355);
or U20068 (N_20068,N_18783,N_19644);
or U20069 (N_20069,N_19124,N_19729);
xnor U20070 (N_20070,N_18507,N_19416);
nand U20071 (N_20071,N_19766,N_18038);
nor U20072 (N_20072,N_19693,N_19222);
or U20073 (N_20073,N_19478,N_18463);
nor U20074 (N_20074,N_18037,N_18380);
or U20075 (N_20075,N_19134,N_19031);
nor U20076 (N_20076,N_19108,N_18210);
xnor U20077 (N_20077,N_19681,N_19734);
nand U20078 (N_20078,N_18563,N_18935);
nand U20079 (N_20079,N_18561,N_18795);
nand U20080 (N_20080,N_18968,N_19278);
and U20081 (N_20081,N_19822,N_19662);
xor U20082 (N_20082,N_19414,N_19908);
or U20083 (N_20083,N_19217,N_19745);
nor U20084 (N_20084,N_18216,N_19312);
nor U20085 (N_20085,N_19863,N_19275);
or U20086 (N_20086,N_19450,N_18312);
and U20087 (N_20087,N_19089,N_19488);
xnor U20088 (N_20088,N_18966,N_18035);
and U20089 (N_20089,N_18712,N_19941);
nor U20090 (N_20090,N_19887,N_18552);
nor U20091 (N_20091,N_19439,N_18826);
nand U20092 (N_20092,N_18130,N_19234);
and U20093 (N_20093,N_18579,N_19161);
and U20094 (N_20094,N_19857,N_19587);
and U20095 (N_20095,N_18184,N_18974);
xor U20096 (N_20096,N_19476,N_19351);
nand U20097 (N_20097,N_18782,N_19233);
nor U20098 (N_20098,N_19149,N_18962);
nor U20099 (N_20099,N_18146,N_19569);
nand U20100 (N_20100,N_19543,N_19349);
nand U20101 (N_20101,N_19267,N_18979);
xor U20102 (N_20102,N_19256,N_19288);
nor U20103 (N_20103,N_18152,N_18531);
xnor U20104 (N_20104,N_19265,N_18177);
nand U20105 (N_20105,N_19718,N_18195);
xnor U20106 (N_20106,N_19254,N_18001);
nand U20107 (N_20107,N_19599,N_19617);
or U20108 (N_20108,N_19402,N_19290);
or U20109 (N_20109,N_19748,N_18363);
xnor U20110 (N_20110,N_18614,N_19457);
nor U20111 (N_20111,N_19084,N_19631);
or U20112 (N_20112,N_18056,N_19043);
nand U20113 (N_20113,N_18804,N_19093);
nor U20114 (N_20114,N_19307,N_19282);
nor U20115 (N_20115,N_18245,N_19555);
or U20116 (N_20116,N_19213,N_19931);
or U20117 (N_20117,N_19366,N_18466);
nand U20118 (N_20118,N_18866,N_18768);
xnor U20119 (N_20119,N_19797,N_18438);
or U20120 (N_20120,N_19930,N_19419);
xnor U20121 (N_20121,N_19983,N_19507);
xnor U20122 (N_20122,N_18445,N_18283);
nor U20123 (N_20123,N_19284,N_19667);
and U20124 (N_20124,N_18863,N_19109);
nor U20125 (N_20125,N_19879,N_18924);
and U20126 (N_20126,N_18920,N_19774);
nand U20127 (N_20127,N_19968,N_18747);
and U20128 (N_20128,N_18621,N_19780);
xnor U20129 (N_20129,N_18250,N_18696);
and U20130 (N_20130,N_18995,N_18771);
nor U20131 (N_20131,N_18435,N_19218);
nor U20132 (N_20132,N_19105,N_18551);
or U20133 (N_20133,N_19484,N_18026);
xor U20134 (N_20134,N_18352,N_18350);
nor U20135 (N_20135,N_18083,N_18674);
or U20136 (N_20136,N_18952,N_18131);
or U20137 (N_20137,N_18406,N_19463);
or U20138 (N_20138,N_19322,N_18401);
nor U20139 (N_20139,N_18589,N_18207);
xnor U20140 (N_20140,N_19840,N_18166);
xor U20141 (N_20141,N_18097,N_18227);
xor U20142 (N_20142,N_18069,N_18325);
or U20143 (N_20143,N_18000,N_18758);
nand U20144 (N_20144,N_18259,N_18933);
and U20145 (N_20145,N_18368,N_19142);
nand U20146 (N_20146,N_19003,N_18870);
nand U20147 (N_20147,N_19785,N_18474);
or U20148 (N_20148,N_18904,N_19921);
xnor U20149 (N_20149,N_18084,N_18457);
xnor U20150 (N_20150,N_18764,N_19513);
and U20151 (N_20151,N_19701,N_19579);
and U20152 (N_20152,N_19020,N_18786);
nor U20153 (N_20153,N_19881,N_19449);
nand U20154 (N_20154,N_19553,N_18067);
and U20155 (N_20155,N_18324,N_19801);
nand U20156 (N_20156,N_19769,N_19974);
and U20157 (N_20157,N_19939,N_18066);
xnor U20158 (N_20158,N_18424,N_19558);
nor U20159 (N_20159,N_18244,N_18949);
xor U20160 (N_20160,N_19090,N_18713);
and U20161 (N_20161,N_19466,N_19654);
nor U20162 (N_20162,N_18900,N_19425);
or U20163 (N_20163,N_19344,N_19739);
nor U20164 (N_20164,N_18967,N_19030);
xor U20165 (N_20165,N_19746,N_18237);
or U20166 (N_20166,N_18102,N_18819);
nor U20167 (N_20167,N_19515,N_18007);
nor U20168 (N_20168,N_18268,N_18894);
nand U20169 (N_20169,N_18396,N_19260);
and U20170 (N_20170,N_19396,N_19577);
xnor U20171 (N_20171,N_18423,N_18046);
or U20172 (N_20172,N_19352,N_18295);
or U20173 (N_20173,N_18822,N_18761);
or U20174 (N_20174,N_19710,N_18540);
nor U20175 (N_20175,N_18088,N_18776);
nand U20176 (N_20176,N_18788,N_19682);
and U20177 (N_20177,N_19809,N_19266);
xnor U20178 (N_20178,N_18246,N_18486);
nand U20179 (N_20179,N_19504,N_19826);
nand U20180 (N_20180,N_18644,N_19182);
xor U20181 (N_20181,N_18711,N_18109);
xnor U20182 (N_20182,N_18730,N_18118);
nand U20183 (N_20183,N_18666,N_18387);
and U20184 (N_20184,N_18526,N_19582);
and U20185 (N_20185,N_18524,N_19337);
nand U20186 (N_20186,N_19520,N_19754);
xnor U20187 (N_20187,N_18701,N_18567);
nor U20188 (N_20188,N_18972,N_19499);
xor U20189 (N_20189,N_18777,N_19184);
and U20190 (N_20190,N_19121,N_19147);
nand U20191 (N_20191,N_18426,N_18476);
xnor U20192 (N_20192,N_18992,N_18969);
nor U20193 (N_20193,N_18055,N_18702);
or U20194 (N_20194,N_18351,N_18231);
or U20195 (N_20195,N_18105,N_19733);
nor U20196 (N_20196,N_19103,N_19318);
nand U20197 (N_20197,N_18065,N_18852);
or U20198 (N_20198,N_18489,N_19073);
and U20199 (N_20199,N_19160,N_18042);
and U20200 (N_20200,N_19037,N_18847);
nand U20201 (N_20201,N_18973,N_18304);
nor U20202 (N_20202,N_18182,N_18480);
or U20203 (N_20203,N_19835,N_19615);
nand U20204 (N_20204,N_19925,N_19660);
nand U20205 (N_20205,N_18191,N_19491);
and U20206 (N_20206,N_18584,N_18840);
and U20207 (N_20207,N_18880,N_19853);
nor U20208 (N_20208,N_19211,N_19023);
nor U20209 (N_20209,N_18262,N_18906);
xnor U20210 (N_20210,N_19742,N_19810);
or U20211 (N_20211,N_18779,N_18343);
xnor U20212 (N_20212,N_19972,N_18721);
or U20213 (N_20213,N_19354,N_19993);
nor U20214 (N_20214,N_19210,N_18305);
nand U20215 (N_20215,N_19987,N_18491);
and U20216 (N_20216,N_18781,N_19057);
or U20217 (N_20217,N_18835,N_18252);
and U20218 (N_20218,N_19977,N_18594);
and U20219 (N_20219,N_19198,N_18817);
or U20220 (N_20220,N_18763,N_18787);
or U20221 (N_20221,N_18175,N_18172);
or U20222 (N_20222,N_19315,N_18676);
xor U20223 (N_20223,N_19110,N_19871);
xnor U20224 (N_20224,N_19434,N_18243);
or U20225 (N_20225,N_18247,N_19635);
nor U20226 (N_20226,N_18796,N_19514);
nor U20227 (N_20227,N_18756,N_19286);
and U20228 (N_20228,N_19381,N_18190);
xnor U20229 (N_20229,N_18803,N_18848);
or U20230 (N_20230,N_18828,N_19750);
and U20231 (N_20231,N_18642,N_19013);
nor U20232 (N_20232,N_18834,N_18201);
or U20233 (N_20233,N_19503,N_18249);
or U20234 (N_20234,N_18873,N_19611);
xnor U20235 (N_20235,N_19944,N_19659);
and U20236 (N_20236,N_19825,N_18317);
nand U20237 (N_20237,N_18490,N_18695);
or U20238 (N_20238,N_18230,N_18140);
nand U20239 (N_20239,N_18641,N_19749);
nand U20240 (N_20240,N_18124,N_19461);
xnor U20241 (N_20241,N_18255,N_19651);
nand U20242 (N_20242,N_19757,N_18269);
or U20243 (N_20243,N_18532,N_19334);
and U20244 (N_20244,N_19329,N_18467);
nor U20245 (N_20245,N_19949,N_19298);
nand U20246 (N_20246,N_18911,N_19884);
nand U20247 (N_20247,N_18392,N_19613);
and U20248 (N_20248,N_18113,N_18500);
or U20249 (N_20249,N_18595,N_19995);
and U20250 (N_20250,N_19619,N_18586);
nor U20251 (N_20251,N_19951,N_18726);
nand U20252 (N_20252,N_18958,N_18668);
nand U20253 (N_20253,N_18444,N_19340);
nand U20254 (N_20254,N_18765,N_18465);
xor U20255 (N_20255,N_19410,N_19743);
nor U20256 (N_20256,N_19241,N_18058);
or U20257 (N_20257,N_19589,N_19860);
nor U20258 (N_20258,N_19095,N_19356);
nor U20259 (N_20259,N_18922,N_19097);
nand U20260 (N_20260,N_19303,N_18961);
nand U20261 (N_20261,N_18810,N_18484);
nor U20262 (N_20262,N_18050,N_19292);
and U20263 (N_20263,N_18882,N_19956);
and U20264 (N_20264,N_19741,N_18927);
nand U20265 (N_20265,N_19872,N_19737);
nor U20266 (N_20266,N_18650,N_19269);
and U20267 (N_20267,N_19692,N_18842);
and U20268 (N_20268,N_19088,N_19598);
nand U20269 (N_20269,N_18892,N_18141);
nand U20270 (N_20270,N_18741,N_18469);
or U20271 (N_20271,N_18613,N_18978);
and U20272 (N_20272,N_18419,N_18431);
and U20273 (N_20273,N_19320,N_18845);
or U20274 (N_20274,N_19890,N_19917);
or U20275 (N_20275,N_18149,N_19394);
nor U20276 (N_20276,N_19685,N_18213);
or U20277 (N_20277,N_19281,N_18222);
or U20278 (N_20278,N_18143,N_18400);
and U20279 (N_20279,N_19928,N_18662);
or U20280 (N_20280,N_19141,N_18253);
nor U20281 (N_20281,N_19534,N_18981);
xor U20282 (N_20282,N_19361,N_18769);
or U20283 (N_20283,N_19187,N_19755);
nand U20284 (N_20284,N_19768,N_19274);
and U20285 (N_20285,N_18068,N_19623);
nand U20286 (N_20286,N_18832,N_18720);
nand U20287 (N_20287,N_19427,N_19408);
nor U20288 (N_20288,N_18837,N_19824);
or U20289 (N_20289,N_18611,N_18329);
xor U20290 (N_20290,N_19091,N_19847);
nand U20291 (N_20291,N_18319,N_19783);
and U20292 (N_20292,N_18615,N_19247);
and U20293 (N_20293,N_18002,N_18204);
and U20294 (N_20294,N_19324,N_18774);
and U20295 (N_20295,N_18723,N_19458);
and U20296 (N_20296,N_19730,N_19678);
xor U20297 (N_20297,N_18938,N_19610);
nor U20298 (N_20298,N_19568,N_19294);
xnor U20299 (N_20299,N_18754,N_18330);
nor U20300 (N_20300,N_18394,N_19482);
xnor U20301 (N_20301,N_19524,N_19335);
and U20302 (N_20302,N_19405,N_19700);
nand U20303 (N_20303,N_19915,N_18142);
nand U20304 (N_20304,N_18784,N_19167);
nor U20305 (N_20305,N_18451,N_18126);
nor U20306 (N_20306,N_19709,N_19596);
nand U20307 (N_20307,N_18956,N_19002);
or U20308 (N_20308,N_19178,N_19898);
xnor U20309 (N_20309,N_19738,N_19521);
nor U20310 (N_20310,N_19536,N_19347);
nand U20311 (N_20311,N_18766,N_18030);
nand U20312 (N_20312,N_19698,N_18285);
nand U20313 (N_20313,N_18448,N_18085);
nand U20314 (N_20314,N_19882,N_19626);
xor U20315 (N_20315,N_19029,N_19072);
nand U20316 (N_20316,N_19495,N_18690);
xor U20317 (N_20317,N_19480,N_19861);
or U20318 (N_20318,N_19646,N_19443);
or U20319 (N_20319,N_18453,N_18820);
or U20320 (N_20320,N_19517,N_19032);
xnor U20321 (N_20321,N_18610,N_18775);
and U20322 (N_20322,N_18792,N_18461);
nor U20323 (N_20323,N_19816,N_19140);
and U20324 (N_20324,N_19954,N_19885);
nand U20325 (N_20325,N_18232,N_19502);
xor U20326 (N_20326,N_18331,N_19948);
or U20327 (N_20327,N_19195,N_18643);
and U20328 (N_20328,N_19638,N_19171);
xnor U20329 (N_20329,N_18953,N_18538);
nor U20330 (N_20330,N_18192,N_19771);
xnor U20331 (N_20331,N_19936,N_18186);
nand U20332 (N_20332,N_19670,N_18619);
xnor U20333 (N_20333,N_19833,N_19287);
nor U20334 (N_20334,N_18737,N_19852);
or U20335 (N_20335,N_18267,N_18012);
nand U20336 (N_20336,N_18150,N_18011);
xnor U20337 (N_20337,N_18694,N_19677);
and U20338 (N_20338,N_18744,N_19120);
nor U20339 (N_20339,N_18289,N_18773);
nand U20340 (N_20340,N_19485,N_19390);
nand U20341 (N_20341,N_18739,N_19855);
and U20342 (N_20342,N_19547,N_18442);
xnor U20343 (N_20343,N_18044,N_19680);
nand U20344 (N_20344,N_18223,N_18183);
or U20345 (N_20345,N_18506,N_18138);
nor U20346 (N_20346,N_19305,N_19650);
nand U20347 (N_20347,N_19444,N_19794);
nor U20348 (N_20348,N_19025,N_18959);
or U20349 (N_20349,N_19614,N_18566);
and U20350 (N_20350,N_19446,N_18336);
nand U20351 (N_20351,N_18313,N_19235);
or U20352 (N_20352,N_19726,N_19914);
nor U20353 (N_20353,N_19111,N_19201);
nor U20354 (N_20354,N_18248,N_18618);
nand U20355 (N_20355,N_18107,N_18637);
xor U20356 (N_20356,N_19959,N_19583);
xor U20357 (N_20357,N_18708,N_19236);
nand U20358 (N_20358,N_18333,N_18443);
and U20359 (N_20359,N_19173,N_19844);
xor U20360 (N_20360,N_18169,N_19049);
nor U20361 (N_20361,N_19238,N_19848);
xnor U20362 (N_20362,N_19788,N_19346);
and U20363 (N_20363,N_19412,N_18412);
nor U20364 (N_20364,N_18196,N_19736);
nand U20365 (N_20365,N_18361,N_19548);
and U20366 (N_20366,N_18573,N_19827);
and U20367 (N_20367,N_19214,N_18385);
nand U20368 (N_20368,N_18111,N_18576);
or U20369 (N_20369,N_19044,N_18170);
nand U20370 (N_20370,N_19906,N_19966);
nor U20371 (N_20371,N_18889,N_19572);
nand U20372 (N_20372,N_19085,N_18692);
and U20373 (N_20373,N_19026,N_19313);
nor U20374 (N_20374,N_18759,N_18179);
or U20375 (N_20375,N_19791,N_18609);
nor U20376 (N_20376,N_18257,N_19492);
or U20377 (N_20377,N_19903,N_18957);
nand U20378 (N_20378,N_19319,N_18094);
nor U20379 (N_20379,N_19336,N_19859);
and U20380 (N_20380,N_19063,N_18569);
and U20381 (N_20381,N_18509,N_18925);
nor U20382 (N_20382,N_19533,N_19665);
nand U20383 (N_20383,N_18556,N_19373);
xnor U20384 (N_20384,N_18799,N_19671);
nor U20385 (N_20385,N_18197,N_19433);
xnor U20386 (N_20386,N_18449,N_19015);
or U20387 (N_20387,N_18898,N_19919);
xnor U20388 (N_20388,N_19684,N_19148);
nand U20389 (N_20389,N_19838,N_18275);
or U20390 (N_20390,N_18178,N_19459);
xnor U20391 (N_20391,N_18153,N_19962);
and U20392 (N_20392,N_19960,N_18521);
xor U20393 (N_20393,N_19304,N_18127);
or U20394 (N_20394,N_19988,N_18399);
or U20395 (N_20395,N_18428,N_19712);
or U20396 (N_20396,N_19829,N_18272);
and U20397 (N_20397,N_19377,N_19168);
xor U20398 (N_20398,N_18063,N_18519);
nor U20399 (N_20399,N_18003,N_18420);
or U20400 (N_20400,N_19883,N_19793);
and U20401 (N_20401,N_18941,N_18757);
and U20402 (N_20402,N_19106,N_19188);
xnor U20403 (N_20403,N_19216,N_19557);
nand U20404 (N_20404,N_19083,N_19308);
or U20405 (N_20405,N_19912,N_18971);
xnor U20406 (N_20406,N_19909,N_19293);
nand U20407 (N_20407,N_19792,N_19230);
nor U20408 (N_20408,N_18332,N_19866);
nand U20409 (N_20409,N_19836,N_19343);
or U20410 (N_20410,N_18114,N_18629);
nor U20411 (N_20411,N_19309,N_19053);
and U20412 (N_20412,N_18871,N_18386);
nand U20413 (N_20413,N_18145,N_19523);
nor U20414 (N_20414,N_18108,N_19632);
and U20415 (N_20415,N_19258,N_19228);
and U20416 (N_20416,N_19666,N_18632);
nand U20417 (N_20417,N_18429,N_19474);
nor U20418 (N_20418,N_18663,N_18098);
nand U20419 (N_20419,N_18487,N_18673);
or U20420 (N_20420,N_18608,N_19052);
or U20421 (N_20421,N_18830,N_19937);
nand U20422 (N_20422,N_18980,N_19969);
or U20423 (N_20423,N_19018,N_19932);
nand U20424 (N_20424,N_19815,N_19181);
or U20425 (N_20425,N_19422,N_18057);
nor U20426 (N_20426,N_19054,N_18010);
nor U20427 (N_20427,N_19376,N_19702);
and U20428 (N_20428,N_18054,N_18926);
and U20429 (N_20429,N_18527,N_19460);
nand U20430 (N_20430,N_19082,N_19328);
or U20431 (N_20431,N_18339,N_19325);
nand U20432 (N_20432,N_19865,N_18539);
nor U20433 (N_20433,N_19027,N_18869);
and U20434 (N_20434,N_19464,N_19719);
nor U20435 (N_20435,N_19259,N_18858);
or U20436 (N_20436,N_19496,N_19122);
xnor U20437 (N_20437,N_19162,N_19971);
and U20438 (N_20438,N_18503,N_19904);
nand U20439 (N_20439,N_18851,N_18879);
xnor U20440 (N_20440,N_19165,N_18173);
and U20441 (N_20441,N_19289,N_19490);
xnor U20442 (N_20442,N_19098,N_18040);
and U20443 (N_20443,N_19744,N_18510);
or U20444 (N_20444,N_18314,N_18544);
xor U20445 (N_20445,N_18299,N_19905);
nor U20446 (N_20446,N_18298,N_19430);
nor U20447 (N_20447,N_18271,N_19649);
nand U20448 (N_20448,N_18502,N_18413);
nand U20449 (N_20449,N_18932,N_18593);
nand U20450 (N_20450,N_19455,N_19441);
or U20451 (N_20451,N_18872,N_18441);
xor U20452 (N_20452,N_18292,N_18121);
or U20453 (N_20453,N_19594,N_19800);
xor U20454 (N_20454,N_19934,N_18537);
xnor U20455 (N_20455,N_18988,N_18439);
nand U20456 (N_20456,N_18414,N_18464);
nand U20457 (N_20457,N_18534,N_18081);
xnor U20458 (N_20458,N_18748,N_18657);
nor U20459 (N_20459,N_18198,N_18543);
xnor U20460 (N_20460,N_19686,N_19843);
nor U20461 (N_20461,N_18542,N_19525);
and U20462 (N_20462,N_18373,N_18151);
and U20463 (N_20463,N_19886,N_19080);
and U20464 (N_20464,N_19409,N_18836);
nor U20465 (N_20465,N_19679,N_19805);
and U20466 (N_20466,N_19401,N_18616);
and U20467 (N_20467,N_19923,N_18742);
nand U20468 (N_20468,N_18393,N_18217);
and U20469 (N_20469,N_18342,N_19772);
or U20470 (N_20470,N_18171,N_19586);
nand U20471 (N_20471,N_18581,N_18047);
xor U20472 (N_20472,N_19077,N_19751);
nand U20473 (N_20473,N_18651,N_19802);
xor U20474 (N_20474,N_18472,N_19870);
xor U20475 (N_20475,N_19101,N_18309);
nor U20476 (N_20476,N_19896,N_19554);
xnor U20477 (N_20477,N_18125,N_18029);
nand U20478 (N_20478,N_18977,N_19628);
nor U20479 (N_20479,N_18923,N_18881);
and U20480 (N_20480,N_18646,N_19130);
or U20481 (N_20481,N_18280,N_19112);
xor U20482 (N_20482,N_18034,N_18590);
or U20483 (N_20483,N_19606,N_18028);
or U20484 (N_20484,N_19916,N_19240);
nand U20485 (N_20485,N_18808,N_18164);
and U20486 (N_20486,N_19874,N_18846);
or U20487 (N_20487,N_19573,N_18477);
nor U20488 (N_20488,N_19117,N_19642);
xor U20489 (N_20489,N_19609,N_18728);
and U20490 (N_20490,N_18752,N_18617);
xor U20491 (N_20491,N_18211,N_18261);
nand U20492 (N_20492,N_18278,N_18221);
nand U20493 (N_20493,N_18203,N_18705);
nor U20494 (N_20494,N_18071,N_18347);
xor U20495 (N_20495,N_19552,N_18416);
xnor U20496 (N_20496,N_18281,N_19470);
and U20497 (N_20497,N_18743,N_18370);
xor U20498 (N_20498,N_19404,N_18523);
and U20499 (N_20499,N_19722,N_18514);
nand U20500 (N_20500,N_19317,N_18717);
or U20501 (N_20501,N_18934,N_19563);
nor U20502 (N_20502,N_18154,N_19529);
nand U20503 (N_20503,N_18800,N_18640);
nor U20504 (N_20504,N_19511,N_18117);
nand U20505 (N_20505,N_18139,N_18824);
nand U20506 (N_20506,N_18485,N_18397);
and U20507 (N_20507,N_19125,N_19174);
nand U20508 (N_20508,N_19880,N_18340);
xnor U20509 (N_20509,N_19094,N_19131);
or U20510 (N_20510,N_18095,N_18492);
and U20511 (N_20511,N_18997,N_18404);
xnor U20512 (N_20512,N_18501,N_18493);
nor U20513 (N_20513,N_18843,N_19970);
and U20514 (N_20514,N_18155,N_19321);
or U20515 (N_20515,N_18345,N_19566);
nand U20516 (N_20516,N_18671,N_18860);
nand U20517 (N_20517,N_19575,N_18536);
or U20518 (N_20518,N_18120,N_19355);
or U20519 (N_20519,N_18425,N_19695);
or U20520 (N_20520,N_18896,N_19697);
nand U20521 (N_20521,N_18014,N_19311);
or U20522 (N_20522,N_18993,N_18680);
nor U20523 (N_20523,N_18129,N_18264);
nor U20524 (N_20524,N_18921,N_18943);
nor U20525 (N_20525,N_19139,N_18948);
xnor U20526 (N_20526,N_18122,N_19858);
or U20527 (N_20527,N_18517,N_18458);
nand U20528 (N_20528,N_19021,N_18174);
or U20529 (N_20529,N_18086,N_19775);
or U20530 (N_20530,N_18778,N_19545);
or U20531 (N_20531,N_18236,N_19323);
or U20532 (N_20532,N_19506,N_18887);
xnor U20533 (N_20533,N_19011,N_19588);
nand U20534 (N_20534,N_19627,N_18286);
nand U20535 (N_20535,N_18936,N_19279);
nand U20536 (N_20536,N_18061,N_18323);
nand U20537 (N_20537,N_18471,N_19519);
and U20538 (N_20538,N_19683,N_18273);
or U20539 (N_20539,N_19357,N_19542);
nand U20540 (N_20540,N_18365,N_19128);
nor U20541 (N_20541,N_18025,N_19839);
nor U20542 (N_20542,N_19560,N_18202);
or U20543 (N_20543,N_19481,N_18116);
and U20544 (N_20544,N_18516,N_18891);
nand U20545 (N_20545,N_19522,N_19873);
nor U20546 (N_20546,N_18999,N_18905);
and U20547 (N_20547,N_18496,N_19075);
and U20548 (N_20548,N_19624,N_19231);
xor U20549 (N_20549,N_18238,N_19982);
or U20550 (N_20550,N_18031,N_19981);
nor U20551 (N_20551,N_19639,N_19841);
nor U20552 (N_20552,N_18546,N_19447);
xnor U20553 (N_20553,N_19169,N_19371);
nand U20554 (N_20554,N_19732,N_18664);
or U20555 (N_20555,N_18520,N_18180);
nor U20556 (N_20556,N_19341,N_18407);
nand U20557 (N_20557,N_19227,N_18015);
or U20558 (N_20558,N_19192,N_19539);
or U20559 (N_20559,N_19986,N_19807);
xnor U20560 (N_20560,N_19877,N_19022);
nor U20561 (N_20561,N_18270,N_18652);
xnor U20562 (N_20562,N_19006,N_18653);
xnor U20563 (N_20563,N_19384,N_18103);
or U20564 (N_20564,N_19603,N_18639);
nand U20565 (N_20565,N_19584,N_19046);
xor U20566 (N_20566,N_18160,N_19854);
and U20567 (N_20567,N_19166,N_19431);
and U20568 (N_20568,N_18648,N_18356);
xnor U20569 (N_20569,N_19946,N_18079);
and U20570 (N_20570,N_18733,N_18901);
and U20571 (N_20571,N_18577,N_18515);
or U20572 (N_20572,N_18983,N_18415);
xnor U20573 (N_20573,N_18366,N_18998);
xor U20574 (N_20574,N_18187,N_18612);
or U20575 (N_20575,N_18867,N_18456);
xnor U20576 (N_20576,N_18917,N_19360);
xnor U20577 (N_20577,N_19918,N_18039);
or U20578 (N_20578,N_18638,N_19518);
xnor U20579 (N_20579,N_19276,N_18434);
nor U20580 (N_20580,N_18740,N_19876);
xnor U20581 (N_20581,N_19891,N_19765);
and U20582 (N_20582,N_19152,N_18410);
nand U20583 (N_20583,N_18346,N_18951);
and U20584 (N_20584,N_19849,N_19758);
nand U20585 (N_20585,N_18601,N_18877);
and U20586 (N_20586,N_19967,N_18602);
and U20587 (N_20587,N_18710,N_18381);
nand U20588 (N_20588,N_18376,N_18092);
xnor U20589 (N_20589,N_19922,N_18535);
nor U20590 (N_20590,N_18772,N_19607);
nand U20591 (N_20591,N_19428,N_18024);
or U20592 (N_20592,N_18942,N_18875);
nand U20593 (N_20593,N_19580,N_19268);
and U20594 (N_20594,N_18013,N_19468);
nand U20595 (N_20595,N_18371,N_19243);
nand U20596 (N_20596,N_18239,N_19508);
xor U20597 (N_20597,N_18645,N_19938);
nand U20598 (N_20598,N_19663,N_18022);
xnor U20599 (N_20599,N_19154,N_19251);
nor U20600 (N_20600,N_19796,N_19012);
nand U20601 (N_20601,N_19009,N_19042);
xor U20602 (N_20602,N_19530,N_18634);
nand U20603 (N_20603,N_19708,N_19237);
or U20604 (N_20604,N_18004,N_19812);
or U20605 (N_20605,N_18937,N_19224);
xor U20606 (N_20606,N_18334,N_19770);
nor U20607 (N_20607,N_19581,N_18931);
nand U20608 (N_20608,N_18403,N_19707);
or U20609 (N_20609,N_19674,N_19295);
and U20610 (N_20610,N_19717,N_18077);
nand U20611 (N_20611,N_18862,N_18437);
nor U20612 (N_20612,N_18854,N_19136);
nand U20613 (N_20613,N_18839,N_19048);
or U20614 (N_20614,N_18886,N_18693);
nor U20615 (N_20615,N_18290,N_18571);
and U20616 (N_20616,N_18233,N_19437);
xnor U20617 (N_20617,N_19203,N_18868);
nor U20618 (N_20618,N_18432,N_19432);
or U20619 (N_20619,N_18048,N_19961);
nand U20620 (N_20620,N_19358,N_18225);
and U20621 (N_20621,N_18954,N_18357);
nor U20622 (N_20622,N_18505,N_19991);
nand U20623 (N_20623,N_19980,N_18718);
xnor U20624 (N_20624,N_19668,N_19000);
and U20625 (N_20625,N_18320,N_19999);
xor U20626 (N_20626,N_18679,N_19270);
and U20627 (N_20627,N_19273,N_18575);
or U20628 (N_20628,N_18036,N_19472);
or U20629 (N_20629,N_18159,N_19990);
nor U20630 (N_20630,N_19779,N_19888);
or U20631 (N_20631,N_18165,N_19035);
xnor U20632 (N_20632,N_19571,N_19616);
and U20633 (N_20633,N_18389,N_18479);
nor U20634 (N_20634,N_18853,N_18970);
nand U20635 (N_20635,N_19633,N_18683);
xnor U20636 (N_20636,N_18557,N_19634);
and U20637 (N_20637,N_19512,N_18303);
or U20638 (N_20638,N_19205,N_18405);
nand U20639 (N_20639,N_18212,N_18812);
nor U20640 (N_20640,N_19947,N_18976);
nor U20641 (N_20641,N_19086,N_19705);
and U20642 (N_20642,N_18082,N_19590);
or U20643 (N_20643,N_19806,N_18989);
nor U20644 (N_20644,N_19151,N_18136);
nor U20645 (N_20645,N_18101,N_18053);
nand U20646 (N_20646,N_19926,N_19784);
xor U20647 (N_20647,N_18655,N_19291);
nand U20648 (N_20648,N_19028,N_19138);
nand U20649 (N_20649,N_19368,N_19979);
nor U20650 (N_20650,N_19636,N_19332);
xor U20651 (N_20651,N_18689,N_19747);
nand U20652 (N_20652,N_18494,N_18529);
or U20653 (N_20653,N_19721,N_19795);
nor U20654 (N_20654,N_19601,N_18685);
xnor U20655 (N_20655,N_18883,N_19735);
nor U20656 (N_20656,N_19630,N_19602);
nand U20657 (N_20657,N_18545,N_18660);
nand U20658 (N_20658,N_19976,N_18627);
nand U20659 (N_20659,N_18033,N_19723);
nand U20660 (N_20660,N_19661,N_19369);
nand U20661 (N_20661,N_18963,N_19372);
and U20662 (N_20662,N_19532,N_19196);
nand U20663 (N_20663,N_19731,N_19541);
nor U20664 (N_20664,N_18119,N_18687);
xor U20665 (N_20665,N_19232,N_19338);
nand U20666 (N_20666,N_19790,N_19248);
and U20667 (N_20667,N_18570,N_19811);
nand U20668 (N_20668,N_19950,N_18930);
xor U20669 (N_20669,N_19096,N_19875);
nor U20670 (N_20670,N_19045,N_18301);
xor U20671 (N_20671,N_18665,N_19263);
nor U20672 (N_20672,N_18789,N_18876);
or U20673 (N_20673,N_19501,N_19331);
and U20674 (N_20674,N_18512,N_19869);
nand U20675 (N_20675,N_18816,N_18688);
xor U20676 (N_20676,N_19510,N_18805);
nand U20677 (N_20677,N_19367,N_18647);
nor U20678 (N_20678,N_19526,N_19528);
or U20679 (N_20679,N_18547,N_18554);
or U20680 (N_20680,N_19019,N_19540);
nor U20681 (N_20681,N_18311,N_18670);
nor U20682 (N_20682,N_19001,N_18335);
and U20683 (N_20683,N_18226,N_19997);
xnor U20684 (N_20684,N_18991,N_19374);
nor U20685 (N_20685,N_18353,N_19957);
and U20686 (N_20686,N_19845,N_18633);
xor U20687 (N_20687,N_18224,N_19244);
xor U20688 (N_20688,N_18681,N_18189);
nand U20689 (N_20689,N_18809,N_19706);
or U20690 (N_20690,N_18328,N_19933);
or U20691 (N_20691,N_19985,N_19429);
or U20692 (N_20692,N_18865,N_18844);
xor U20693 (N_20693,N_18498,N_19143);
or U20694 (N_20694,N_18430,N_19864);
nand U20695 (N_20695,N_19215,N_18296);
xnor U20696 (N_20696,N_18344,N_19834);
nor U20697 (N_20697,N_19179,N_18878);
nor U20698 (N_20698,N_19475,N_18770);
or U20699 (N_20699,N_19943,N_18675);
or U20700 (N_20700,N_18409,N_19159);
or U20701 (N_20701,N_19223,N_18706);
nand U20702 (N_20702,N_18215,N_19426);
xor U20703 (N_20703,N_18985,N_19062);
xor U20704 (N_20704,N_18588,N_18398);
nor U20705 (N_20705,N_19144,N_19421);
nor U20706 (N_20706,N_18622,N_19393);
xnor U20707 (N_20707,N_19348,N_18874);
nor U20708 (N_20708,N_18110,N_19778);
xor U20709 (N_20709,N_19462,N_18550);
and U20710 (N_20710,N_18228,N_19942);
nand U20711 (N_20711,N_18755,N_18274);
or U20712 (N_20712,N_19920,N_18960);
or U20713 (N_20713,N_19306,N_19998);
and U20714 (N_20714,N_19669,N_18006);
xor U20715 (N_20715,N_18982,N_19387);
nor U20716 (N_20716,N_18797,N_19415);
or U20717 (N_20717,N_19116,N_19071);
or U20718 (N_20718,N_18630,N_19537);
and U20719 (N_20719,N_18070,N_18568);
nand U20720 (N_20720,N_18360,N_19637);
nor U20721 (N_20721,N_19442,N_18919);
or U20722 (N_20722,N_18760,N_18798);
and U20723 (N_20723,N_18909,N_19551);
xor U20724 (N_20724,N_19271,N_19039);
or U20725 (N_20725,N_18080,N_19544);
and U20726 (N_20726,N_19927,N_18338);
or U20727 (N_20727,N_18857,N_18624);
nand U20728 (N_20728,N_19185,N_18700);
nor U20729 (N_20729,N_19041,N_18027);
nand U20730 (N_20730,N_18732,N_18020);
or U20731 (N_20731,N_19145,N_19895);
or U20732 (N_20732,N_18849,N_18861);
xnor U20733 (N_20733,N_19994,N_19486);
nand U20734 (N_20734,N_19479,N_18468);
nand U20735 (N_20735,N_18677,N_18899);
and U20736 (N_20736,N_18893,N_19473);
xor U20737 (N_20737,N_18965,N_19137);
xor U20738 (N_20738,N_18104,N_18229);
and U20739 (N_20739,N_19004,N_18043);
and U20740 (N_20740,N_19672,N_18750);
nor U20741 (N_20741,N_18349,N_18603);
nand U20742 (N_20742,N_18162,N_19625);
xnor U20743 (N_20743,N_18572,N_18525);
nor U20744 (N_20744,N_19175,N_19894);
xnor U20745 (N_20745,N_18833,N_18156);
or U20746 (N_20746,N_19064,N_18897);
and U20747 (N_20747,N_19252,N_19386);
and U20748 (N_20748,N_19561,N_19114);
nand U20749 (N_20749,N_19699,N_18829);
xor U20750 (N_20750,N_18326,N_19591);
and U20751 (N_20751,N_19033,N_19498);
xor U20752 (N_20752,N_18017,N_18541);
xnor U20753 (N_20753,N_19996,N_19621);
nor U20754 (N_20754,N_18188,N_19658);
xnor U20755 (N_20755,N_19567,N_19061);
and U20756 (N_20756,N_19107,N_18821);
nand U20757 (N_20757,N_19250,N_18427);
nand U20758 (N_20758,N_19831,N_19158);
xnor U20759 (N_20759,N_19392,N_19333);
nor U20760 (N_20760,N_18859,N_18446);
nor U20761 (N_20761,N_19172,N_18470);
nand U20762 (N_20762,N_18205,N_18562);
xnor U20763 (N_20763,N_18106,N_18709);
nand U20764 (N_20764,N_19477,N_19759);
and U20765 (N_20765,N_19965,N_18574);
nand U20766 (N_20766,N_19067,N_19353);
or U20767 (N_20767,N_18850,N_19163);
xnor U20768 (N_20768,N_19958,N_18193);
xor U20769 (N_20769,N_19257,N_18185);
or U20770 (N_20770,N_18697,N_19955);
or U20771 (N_20771,N_19383,N_18635);
xor U20772 (N_20772,N_18667,N_18745);
nand U20773 (N_20773,N_19527,N_19087);
xnor U20774 (N_20774,N_18598,N_18288);
or U20775 (N_20775,N_18307,N_18604);
or U20776 (N_20776,N_19975,N_18234);
nand U20777 (N_20777,N_18597,N_18168);
xor U20778 (N_20778,N_18885,N_19516);
nor U20779 (N_20779,N_19424,N_19283);
or U20780 (N_20780,N_19720,N_18591);
nand U20781 (N_20781,N_19221,N_19804);
nor U20782 (N_20782,N_19411,N_19964);
or U20783 (N_20783,N_18945,N_18518);
or U20784 (N_20784,N_19940,N_18176);
nand U20785 (N_20785,N_19074,N_18890);
or U20786 (N_20786,N_19711,N_18802);
nor U20787 (N_20787,N_19612,N_19191);
nor U20788 (N_20788,N_18447,N_18746);
nand U20789 (N_20789,N_19762,N_18478);
or U20790 (N_20790,N_18135,N_19190);
nor U20791 (N_20791,N_18287,N_18888);
or U20792 (N_20792,N_18533,N_18219);
and U20793 (N_20793,N_18062,N_19406);
and U20794 (N_20794,N_18559,N_19454);
nand U20795 (N_20795,N_18649,N_18814);
and U20796 (N_20796,N_18684,N_19645);
and U20797 (N_20797,N_19302,N_19010);
nor U20798 (N_20798,N_18583,N_19092);
or U20799 (N_20799,N_18714,N_18388);
and U20800 (N_20800,N_18987,N_18475);
xor U20801 (N_20801,N_19391,N_18214);
and U20802 (N_20802,N_19316,N_18282);
nand U20803 (N_20803,N_19655,N_18297);
nand U20804 (N_20804,N_19629,N_19219);
nand U20805 (N_20805,N_18128,N_19535);
nand U20806 (N_20806,N_18497,N_18209);
nand U20807 (N_20807,N_18115,N_18391);
nor U20808 (N_20808,N_19060,N_19789);
nor U20809 (N_20809,N_18580,N_18767);
or U20810 (N_20810,N_18374,N_19299);
nand U20811 (N_20811,N_18582,N_18220);
xor U20812 (N_20812,N_18686,N_19050);
xnor U20813 (N_20813,N_18607,N_19438);
and U20814 (N_20814,N_19696,N_18382);
or U20815 (N_20815,N_19070,N_19242);
xnor U20816 (N_20816,N_19264,N_18377);
and U20817 (N_20817,N_19752,N_18738);
and U20818 (N_20818,N_18059,N_19691);
xnor U20819 (N_20819,N_18099,N_19310);
and U20820 (N_20820,N_18258,N_19066);
xnor U20821 (N_20821,N_19818,N_18751);
nand U20822 (N_20822,N_18975,N_19445);
xnor U20823 (N_20823,N_18016,N_19132);
and U20824 (N_20824,N_18009,N_18263);
or U20825 (N_20825,N_18008,N_19339);
nor U20826 (N_20826,N_19058,N_19456);
and U20827 (N_20827,N_18384,N_19652);
or U20828 (N_20828,N_18251,N_19714);
and U20829 (N_20829,N_18801,N_18294);
or U20830 (N_20830,N_19878,N_19868);
nor U20831 (N_20831,N_19643,N_19777);
nand U20832 (N_20832,N_19024,N_19786);
xor U20833 (N_20833,N_19420,N_18513);
xnor U20834 (N_20834,N_18418,N_18530);
nand U20835 (N_20835,N_18827,N_18856);
or U20836 (N_20836,N_19761,N_19359);
xnor U20837 (N_20837,N_18144,N_19129);
nand U20838 (N_20838,N_19657,N_18161);
or U20839 (N_20839,N_18348,N_19687);
or U20840 (N_20840,N_18553,N_18913);
nor U20841 (N_20841,N_19435,N_19565);
nand U20842 (N_20842,N_18256,N_19489);
xnor U20843 (N_20843,N_18815,N_19330);
nor U20844 (N_20844,N_18241,N_19798);
nor U20845 (N_20845,N_19673,N_19924);
xnor U20846 (N_20846,N_18606,N_18884);
or U20847 (N_20847,N_18041,N_18823);
and U20848 (N_20848,N_19407,N_19595);
nor U20849 (N_20849,N_19399,N_19945);
xnor U20850 (N_20850,N_18235,N_19135);
and U20851 (N_20851,N_19153,N_18359);
or U20852 (N_20852,N_19992,N_18605);
and U20853 (N_20853,N_18454,N_19007);
nor U20854 (N_20854,N_19370,N_18895);
nand U20855 (N_20855,N_19133,N_18731);
xor U20856 (N_20856,N_19277,N_19728);
or U20857 (N_20857,N_19497,N_19180);
nand U20858 (N_20858,N_18736,N_19385);
xnor U20859 (N_20859,N_19664,N_18549);
and U20860 (N_20860,N_19618,N_19653);
nand U20861 (N_20861,N_19115,N_18626);
nor U20862 (N_20862,N_18592,N_18495);
nand U20863 (N_20863,N_19076,N_18818);
and U20864 (N_20864,N_18528,N_18005);
nand U20865 (N_20865,N_19239,N_18395);
and U20866 (N_20866,N_18436,N_19963);
nand U20867 (N_20867,N_19008,N_19100);
nand U20868 (N_20868,N_18996,N_18914);
nor U20869 (N_20869,N_18994,N_19469);
xnor U20870 (N_20870,N_19837,N_19059);
or U20871 (N_20871,N_19379,N_19782);
nor U20872 (N_20872,N_19756,N_18794);
or U20873 (N_20873,N_18473,N_19767);
nor U20874 (N_20874,N_18729,N_19559);
or U20875 (N_20875,N_18481,N_18669);
nor U20876 (N_20876,N_18807,N_18918);
or U20877 (N_20877,N_19451,N_19113);
and U20878 (N_20878,N_19170,N_18019);
nor U20879 (N_20879,N_18793,N_19803);
xnor U20880 (N_20880,N_19823,N_18658);
and U20881 (N_20881,N_18724,N_18631);
nand U20882 (N_20882,N_18284,N_18555);
nor U20883 (N_20883,N_18459,N_19194);
nor U20884 (N_20884,N_18452,N_19397);
or U20885 (N_20885,N_19689,N_19850);
and U20886 (N_20886,N_18310,N_19056);
nand U20887 (N_20887,N_19005,N_19204);
or U20888 (N_20888,N_19549,N_19069);
nor U20889 (N_20889,N_18075,N_19952);
and U20890 (N_20890,N_18928,N_18716);
and U20891 (N_20891,N_19483,N_19220);
nor U20892 (N_20892,N_18838,N_19262);
nand U20893 (N_20893,N_19375,N_19984);
or U20894 (N_20894,N_19900,N_18625);
nor U20895 (N_20895,N_18940,N_19362);
and U20896 (N_20896,N_18218,N_19467);
and U20897 (N_20897,N_18199,N_18072);
and U20898 (N_20898,N_19081,N_18620);
nand U20899 (N_20899,N_18060,N_18460);
nand U20900 (N_20900,N_19452,N_18912);
and U20901 (N_20901,N_18955,N_19703);
nor U20902 (N_20902,N_18806,N_18749);
nor U20903 (N_20903,N_18947,N_18200);
nor U20904 (N_20904,N_19157,N_19126);
nand U20905 (N_20905,N_18623,N_19423);
xor U20906 (N_20906,N_19828,N_18052);
or U20907 (N_20907,N_18672,N_19448);
nor U20908 (N_20908,N_18929,N_18727);
or U20909 (N_20909,N_18315,N_18112);
xor U20910 (N_20910,N_19327,N_19055);
nand U20911 (N_20911,N_18293,N_18018);
and U20912 (N_20912,N_18522,N_18091);
nor U20913 (N_20913,N_19608,N_19989);
and U20914 (N_20914,N_18078,N_19910);
or U20915 (N_20915,N_18903,N_19123);
or U20916 (N_20916,N_19694,N_19911);
nand U20917 (N_20917,N_18440,N_18021);
nor U20918 (N_20918,N_19297,N_18600);
and U20919 (N_20919,N_18565,N_18964);
nand U20920 (N_20920,N_19380,N_19301);
nor U20921 (N_20921,N_19314,N_19017);
and U20922 (N_20922,N_19531,N_18076);
nor U20923 (N_20923,N_19342,N_19118);
nand U20924 (N_20924,N_19040,N_19574);
or U20925 (N_20925,N_19202,N_18337);
or U20926 (N_20926,N_19724,N_18916);
nand U20927 (N_20927,N_18341,N_18841);
nor U20928 (N_20928,N_18408,N_18560);
nor U20929 (N_20929,N_18910,N_18045);
xnor U20930 (N_20930,N_18811,N_18499);
nand U20931 (N_20931,N_19494,N_19713);
nor U20932 (N_20932,N_19929,N_19272);
nand U20933 (N_20933,N_19592,N_19620);
nand U20934 (N_20934,N_18096,N_18715);
nor U20935 (N_20935,N_19280,N_18984);
nor U20936 (N_20936,N_19378,N_19570);
xnor U20937 (N_20937,N_18587,N_19753);
and U20938 (N_20938,N_19199,N_19212);
xor U20939 (N_20939,N_18276,N_18358);
or U20940 (N_20940,N_18433,N_18147);
nor U20941 (N_20941,N_19597,N_18362);
and U20942 (N_20942,N_19604,N_19605);
and U20943 (N_20943,N_19907,N_19034);
nand U20944 (N_20944,N_19189,N_18417);
and U20945 (N_20945,N_18790,N_18558);
and U20946 (N_20946,N_19417,N_18950);
xor U20947 (N_20947,N_19799,N_18367);
nand U20948 (N_20948,N_19471,N_19345);
or U20949 (N_20949,N_19487,N_18148);
and U20950 (N_20950,N_18902,N_18132);
and U20951 (N_20951,N_19413,N_19892);
nand U20952 (N_20952,N_19065,N_19183);
and U20953 (N_20953,N_19155,N_18944);
nor U20954 (N_20954,N_18585,N_19978);
or U20955 (N_20955,N_18813,N_18636);
or U20956 (N_20956,N_19382,N_19716);
xnor U20957 (N_20957,N_19127,N_19177);
or U20958 (N_20958,N_18791,N_18354);
nor U20959 (N_20959,N_19261,N_19365);
and U20960 (N_20960,N_19208,N_18074);
and U20961 (N_20961,N_18308,N_19078);
and U20962 (N_20962,N_19036,N_19047);
nand U20963 (N_20963,N_19150,N_19740);
xnor U20964 (N_20964,N_19556,N_18704);
and U20965 (N_20965,N_19550,N_19207);
nor U20966 (N_20966,N_18698,N_18825);
nor U20967 (N_20967,N_18158,N_18946);
xor U20968 (N_20968,N_19389,N_19640);
nor U20969 (N_20969,N_18831,N_18093);
nor U20970 (N_20970,N_19186,N_19832);
nor U20971 (N_20971,N_19388,N_19104);
xor U20972 (N_20972,N_19787,N_19068);
nand U20973 (N_20973,N_19773,N_18915);
or U20974 (N_20974,N_18762,N_19253);
or U20975 (N_20975,N_18260,N_18206);
xnor U20976 (N_20976,N_18659,N_19051);
or U20977 (N_20977,N_18596,N_18661);
nor U20978 (N_20978,N_19296,N_18907);
and U20979 (N_20979,N_19364,N_18599);
or U20980 (N_20980,N_19781,N_18939);
nor U20981 (N_20981,N_18327,N_18181);
nand U20982 (N_20982,N_18383,N_18089);
nor U20983 (N_20983,N_18654,N_18375);
xnor U20984 (N_20984,N_19119,N_18421);
or U20985 (N_20985,N_18504,N_19403);
nor U20986 (N_20986,N_18379,N_19821);
nand U20987 (N_20987,N_18049,N_18306);
or U20988 (N_20988,N_19176,N_19641);
nor U20989 (N_20989,N_18735,N_19760);
and U20990 (N_20990,N_18364,N_18411);
or U20991 (N_20991,N_19851,N_19562);
nor U20992 (N_20992,N_19326,N_19856);
nor U20993 (N_20993,N_18100,N_18578);
nand U20994 (N_20994,N_18656,N_19600);
or U20995 (N_20995,N_18908,N_19776);
xnor U20996 (N_20996,N_19813,N_18123);
xor U20997 (N_20997,N_19564,N_19585);
nand U20998 (N_20998,N_19808,N_18990);
and U20999 (N_20999,N_18302,N_19016);
nor U21000 (N_21000,N_19130,N_19242);
xor U21001 (N_21001,N_18146,N_18697);
xnor U21002 (N_21002,N_18135,N_19516);
and U21003 (N_21003,N_19996,N_18770);
xnor U21004 (N_21004,N_19638,N_18686);
nand U21005 (N_21005,N_18347,N_19689);
nor U21006 (N_21006,N_19485,N_19172);
and U21007 (N_21007,N_19885,N_19660);
nor U21008 (N_21008,N_19696,N_19952);
nor U21009 (N_21009,N_18939,N_18152);
nand U21010 (N_21010,N_19485,N_18836);
xor U21011 (N_21011,N_19839,N_19829);
nand U21012 (N_21012,N_19782,N_18167);
or U21013 (N_21013,N_18228,N_19733);
xnor U21014 (N_21014,N_19675,N_18770);
xor U21015 (N_21015,N_19898,N_19864);
nand U21016 (N_21016,N_18712,N_18688);
xor U21017 (N_21017,N_18971,N_19942);
nor U21018 (N_21018,N_19357,N_18848);
and U21019 (N_21019,N_18585,N_19130);
xnor U21020 (N_21020,N_18993,N_19558);
and U21021 (N_21021,N_18139,N_19808);
nand U21022 (N_21022,N_18130,N_19021);
and U21023 (N_21023,N_18520,N_18797);
and U21024 (N_21024,N_18088,N_19668);
or U21025 (N_21025,N_18847,N_19769);
xor U21026 (N_21026,N_19660,N_18986);
xor U21027 (N_21027,N_19513,N_18715);
nand U21028 (N_21028,N_18595,N_19628);
and U21029 (N_21029,N_18013,N_19369);
nand U21030 (N_21030,N_18107,N_19057);
xnor U21031 (N_21031,N_19373,N_19096);
and U21032 (N_21032,N_19625,N_18211);
or U21033 (N_21033,N_18156,N_18059);
and U21034 (N_21034,N_18071,N_19778);
nand U21035 (N_21035,N_18323,N_18108);
nor U21036 (N_21036,N_19275,N_19211);
and U21037 (N_21037,N_19096,N_19433);
nand U21038 (N_21038,N_19348,N_19445);
and U21039 (N_21039,N_19332,N_18473);
nor U21040 (N_21040,N_18531,N_19343);
or U21041 (N_21041,N_18860,N_18416);
and U21042 (N_21042,N_18885,N_19747);
and U21043 (N_21043,N_18825,N_18604);
nor U21044 (N_21044,N_18673,N_18340);
nor U21045 (N_21045,N_19407,N_19342);
nor U21046 (N_21046,N_18771,N_19318);
and U21047 (N_21047,N_19999,N_19957);
xor U21048 (N_21048,N_19973,N_18497);
nor U21049 (N_21049,N_19410,N_18470);
nand U21050 (N_21050,N_18326,N_18339);
and U21051 (N_21051,N_19909,N_19215);
nor U21052 (N_21052,N_19711,N_19662);
nand U21053 (N_21053,N_18114,N_19042);
nor U21054 (N_21054,N_19059,N_19364);
or U21055 (N_21055,N_18129,N_18962);
and U21056 (N_21056,N_18001,N_18324);
or U21057 (N_21057,N_18337,N_18182);
nor U21058 (N_21058,N_18390,N_19385);
nor U21059 (N_21059,N_19364,N_18981);
nand U21060 (N_21060,N_18519,N_19058);
or U21061 (N_21061,N_19307,N_18354);
xor U21062 (N_21062,N_18705,N_18977);
xnor U21063 (N_21063,N_18564,N_18890);
nand U21064 (N_21064,N_18684,N_19293);
xor U21065 (N_21065,N_18659,N_18386);
nor U21066 (N_21066,N_18006,N_18087);
or U21067 (N_21067,N_19243,N_19767);
or U21068 (N_21068,N_18216,N_18743);
xnor U21069 (N_21069,N_18082,N_18229);
or U21070 (N_21070,N_19415,N_19046);
nor U21071 (N_21071,N_18863,N_19460);
nor U21072 (N_21072,N_18558,N_19487);
or U21073 (N_21073,N_18709,N_18982);
xor U21074 (N_21074,N_19763,N_18558);
nand U21075 (N_21075,N_18566,N_19108);
nor U21076 (N_21076,N_19611,N_18709);
nor U21077 (N_21077,N_19569,N_18814);
nand U21078 (N_21078,N_19671,N_18871);
nor U21079 (N_21079,N_18778,N_18576);
or U21080 (N_21080,N_19084,N_18847);
nor U21081 (N_21081,N_19184,N_19766);
xnor U21082 (N_21082,N_18975,N_19647);
nand U21083 (N_21083,N_18743,N_18571);
nand U21084 (N_21084,N_19463,N_18566);
and U21085 (N_21085,N_19705,N_19531);
and U21086 (N_21086,N_18902,N_19365);
nand U21087 (N_21087,N_18183,N_18884);
nor U21088 (N_21088,N_18450,N_18751);
and U21089 (N_21089,N_19828,N_19261);
or U21090 (N_21090,N_18051,N_18045);
nand U21091 (N_21091,N_18647,N_18654);
and U21092 (N_21092,N_18136,N_18390);
xnor U21093 (N_21093,N_19337,N_19291);
or U21094 (N_21094,N_19526,N_18677);
xnor U21095 (N_21095,N_18578,N_18122);
and U21096 (N_21096,N_19596,N_18455);
nand U21097 (N_21097,N_19701,N_19441);
and U21098 (N_21098,N_19032,N_18826);
and U21099 (N_21099,N_18735,N_19298);
or U21100 (N_21100,N_18395,N_18086);
or U21101 (N_21101,N_19122,N_18706);
and U21102 (N_21102,N_19986,N_18405);
and U21103 (N_21103,N_18184,N_18180);
xor U21104 (N_21104,N_19293,N_18691);
and U21105 (N_21105,N_18434,N_19246);
xnor U21106 (N_21106,N_18125,N_18368);
nor U21107 (N_21107,N_19521,N_18877);
nor U21108 (N_21108,N_19595,N_19178);
and U21109 (N_21109,N_19288,N_18446);
nand U21110 (N_21110,N_19158,N_19234);
or U21111 (N_21111,N_18956,N_19893);
and U21112 (N_21112,N_19231,N_18089);
nand U21113 (N_21113,N_18673,N_19812);
nor U21114 (N_21114,N_19535,N_18536);
or U21115 (N_21115,N_19322,N_19416);
or U21116 (N_21116,N_18148,N_18991);
nand U21117 (N_21117,N_19281,N_19954);
and U21118 (N_21118,N_18583,N_18788);
or U21119 (N_21119,N_18575,N_18492);
xnor U21120 (N_21120,N_19613,N_18523);
xor U21121 (N_21121,N_19066,N_18851);
nand U21122 (N_21122,N_18194,N_19383);
nor U21123 (N_21123,N_18676,N_18131);
nand U21124 (N_21124,N_19115,N_19001);
or U21125 (N_21125,N_18688,N_19937);
or U21126 (N_21126,N_18727,N_18188);
nand U21127 (N_21127,N_19454,N_18540);
xnor U21128 (N_21128,N_19434,N_19842);
xnor U21129 (N_21129,N_18171,N_18137);
nand U21130 (N_21130,N_19067,N_19947);
nor U21131 (N_21131,N_19014,N_18407);
xor U21132 (N_21132,N_18973,N_18781);
nand U21133 (N_21133,N_18516,N_19236);
and U21134 (N_21134,N_18437,N_19804);
and U21135 (N_21135,N_18784,N_19417);
xor U21136 (N_21136,N_18400,N_19974);
nand U21137 (N_21137,N_18022,N_19476);
and U21138 (N_21138,N_18607,N_19485);
and U21139 (N_21139,N_19583,N_18856);
or U21140 (N_21140,N_18316,N_19155);
or U21141 (N_21141,N_19445,N_19308);
nor U21142 (N_21142,N_19141,N_18848);
and U21143 (N_21143,N_18301,N_19570);
nand U21144 (N_21144,N_19794,N_19074);
nor U21145 (N_21145,N_18140,N_19764);
nand U21146 (N_21146,N_19869,N_19864);
or U21147 (N_21147,N_18049,N_19195);
or U21148 (N_21148,N_19460,N_18577);
xor U21149 (N_21149,N_19756,N_19132);
or U21150 (N_21150,N_18765,N_18653);
or U21151 (N_21151,N_18703,N_19778);
and U21152 (N_21152,N_18353,N_18450);
and U21153 (N_21153,N_19809,N_19675);
and U21154 (N_21154,N_19079,N_18508);
or U21155 (N_21155,N_19893,N_18795);
nor U21156 (N_21156,N_19964,N_19186);
nand U21157 (N_21157,N_18012,N_18988);
nor U21158 (N_21158,N_19228,N_18727);
nor U21159 (N_21159,N_19886,N_18237);
and U21160 (N_21160,N_18379,N_18912);
or U21161 (N_21161,N_19390,N_19557);
xor U21162 (N_21162,N_18794,N_19716);
or U21163 (N_21163,N_18812,N_18146);
nand U21164 (N_21164,N_18329,N_18080);
and U21165 (N_21165,N_18664,N_19201);
and U21166 (N_21166,N_18072,N_19925);
nor U21167 (N_21167,N_18038,N_19856);
and U21168 (N_21168,N_18267,N_18556);
nor U21169 (N_21169,N_18133,N_18217);
xor U21170 (N_21170,N_19570,N_18158);
nor U21171 (N_21171,N_19731,N_18338);
and U21172 (N_21172,N_19279,N_18184);
nor U21173 (N_21173,N_18922,N_19711);
or U21174 (N_21174,N_18537,N_18314);
xor U21175 (N_21175,N_18037,N_18546);
or U21176 (N_21176,N_19297,N_18824);
nor U21177 (N_21177,N_18702,N_19794);
and U21178 (N_21178,N_19581,N_18845);
or U21179 (N_21179,N_18076,N_19162);
nor U21180 (N_21180,N_18758,N_18098);
nand U21181 (N_21181,N_19885,N_19167);
nand U21182 (N_21182,N_19503,N_18259);
nor U21183 (N_21183,N_18225,N_18467);
and U21184 (N_21184,N_18782,N_19919);
nor U21185 (N_21185,N_18216,N_19595);
xor U21186 (N_21186,N_19394,N_19949);
nand U21187 (N_21187,N_19773,N_19846);
nor U21188 (N_21188,N_18137,N_19906);
xnor U21189 (N_21189,N_18923,N_19374);
xor U21190 (N_21190,N_18498,N_18169);
nor U21191 (N_21191,N_18057,N_19770);
or U21192 (N_21192,N_19430,N_18159);
or U21193 (N_21193,N_18626,N_19620);
nor U21194 (N_21194,N_18269,N_19849);
or U21195 (N_21195,N_19784,N_19428);
or U21196 (N_21196,N_18312,N_18361);
nand U21197 (N_21197,N_18805,N_18912);
and U21198 (N_21198,N_18825,N_19864);
and U21199 (N_21199,N_19575,N_18854);
or U21200 (N_21200,N_18121,N_18706);
nor U21201 (N_21201,N_18394,N_19995);
nand U21202 (N_21202,N_19661,N_18021);
xnor U21203 (N_21203,N_19353,N_19879);
nor U21204 (N_21204,N_18781,N_19358);
nand U21205 (N_21205,N_19967,N_19524);
and U21206 (N_21206,N_18990,N_19417);
and U21207 (N_21207,N_19619,N_18410);
xor U21208 (N_21208,N_19080,N_18249);
or U21209 (N_21209,N_18285,N_18897);
nand U21210 (N_21210,N_18133,N_19042);
nor U21211 (N_21211,N_18677,N_19733);
and U21212 (N_21212,N_19839,N_19457);
nand U21213 (N_21213,N_19682,N_19084);
or U21214 (N_21214,N_19537,N_18579);
xor U21215 (N_21215,N_19851,N_19672);
and U21216 (N_21216,N_19426,N_18104);
and U21217 (N_21217,N_19483,N_18171);
nor U21218 (N_21218,N_19665,N_18997);
nor U21219 (N_21219,N_18556,N_18839);
or U21220 (N_21220,N_19929,N_19286);
and U21221 (N_21221,N_19118,N_19801);
nor U21222 (N_21222,N_18340,N_19029);
or U21223 (N_21223,N_19966,N_18860);
xor U21224 (N_21224,N_18325,N_18443);
xnor U21225 (N_21225,N_19410,N_18097);
nor U21226 (N_21226,N_18704,N_19987);
nor U21227 (N_21227,N_18896,N_19687);
nand U21228 (N_21228,N_19035,N_18975);
nand U21229 (N_21229,N_19343,N_18990);
xor U21230 (N_21230,N_19272,N_18624);
or U21231 (N_21231,N_19146,N_18040);
or U21232 (N_21232,N_19923,N_18084);
nor U21233 (N_21233,N_18312,N_19875);
nor U21234 (N_21234,N_19043,N_18500);
or U21235 (N_21235,N_18485,N_18144);
xor U21236 (N_21236,N_19753,N_19217);
nand U21237 (N_21237,N_19834,N_18145);
or U21238 (N_21238,N_18125,N_18724);
and U21239 (N_21239,N_18662,N_19082);
and U21240 (N_21240,N_18417,N_18938);
nand U21241 (N_21241,N_19042,N_19154);
nand U21242 (N_21242,N_18482,N_19494);
nand U21243 (N_21243,N_18478,N_18010);
xor U21244 (N_21244,N_19807,N_19292);
and U21245 (N_21245,N_19596,N_18202);
nand U21246 (N_21246,N_19151,N_19888);
xnor U21247 (N_21247,N_19962,N_19464);
or U21248 (N_21248,N_18440,N_18275);
nor U21249 (N_21249,N_19541,N_18828);
nor U21250 (N_21250,N_19016,N_19911);
and U21251 (N_21251,N_18258,N_19875);
nand U21252 (N_21252,N_19742,N_18289);
or U21253 (N_21253,N_18842,N_18205);
nand U21254 (N_21254,N_18041,N_19082);
or U21255 (N_21255,N_19578,N_18462);
nor U21256 (N_21256,N_18390,N_18265);
or U21257 (N_21257,N_19093,N_18902);
nand U21258 (N_21258,N_19712,N_18360);
and U21259 (N_21259,N_19631,N_18696);
or U21260 (N_21260,N_19069,N_18727);
nand U21261 (N_21261,N_19686,N_18559);
nor U21262 (N_21262,N_19102,N_18224);
and U21263 (N_21263,N_19338,N_19153);
or U21264 (N_21264,N_18484,N_19928);
nand U21265 (N_21265,N_19997,N_18872);
or U21266 (N_21266,N_18899,N_18350);
xor U21267 (N_21267,N_19475,N_18075);
or U21268 (N_21268,N_19321,N_18903);
or U21269 (N_21269,N_18341,N_18618);
or U21270 (N_21270,N_18945,N_19584);
xor U21271 (N_21271,N_19212,N_18310);
nand U21272 (N_21272,N_19576,N_19260);
xor U21273 (N_21273,N_19848,N_19166);
nor U21274 (N_21274,N_18542,N_19596);
and U21275 (N_21275,N_18450,N_18037);
nand U21276 (N_21276,N_18201,N_18167);
and U21277 (N_21277,N_18784,N_18056);
and U21278 (N_21278,N_19792,N_19539);
xor U21279 (N_21279,N_18380,N_19893);
nand U21280 (N_21280,N_19802,N_18269);
or U21281 (N_21281,N_18178,N_19621);
xnor U21282 (N_21282,N_19055,N_18557);
nand U21283 (N_21283,N_18399,N_19701);
and U21284 (N_21284,N_19208,N_18401);
xor U21285 (N_21285,N_18645,N_18778);
nand U21286 (N_21286,N_19984,N_18434);
nand U21287 (N_21287,N_19731,N_19274);
nor U21288 (N_21288,N_19838,N_18201);
nand U21289 (N_21289,N_18501,N_19766);
xnor U21290 (N_21290,N_19665,N_19571);
and U21291 (N_21291,N_19305,N_18997);
xor U21292 (N_21292,N_18802,N_19983);
nor U21293 (N_21293,N_18949,N_18596);
nand U21294 (N_21294,N_18062,N_19789);
xnor U21295 (N_21295,N_19614,N_19849);
and U21296 (N_21296,N_18885,N_18787);
or U21297 (N_21297,N_19598,N_19991);
xor U21298 (N_21298,N_18119,N_18419);
xor U21299 (N_21299,N_19814,N_18978);
xnor U21300 (N_21300,N_19820,N_19451);
nand U21301 (N_21301,N_19827,N_19629);
and U21302 (N_21302,N_19667,N_19641);
and U21303 (N_21303,N_19868,N_18345);
and U21304 (N_21304,N_18365,N_19070);
xnor U21305 (N_21305,N_18296,N_19890);
nor U21306 (N_21306,N_19995,N_19581);
or U21307 (N_21307,N_18015,N_18058);
nand U21308 (N_21308,N_18595,N_19787);
or U21309 (N_21309,N_19239,N_18114);
nand U21310 (N_21310,N_18064,N_18926);
or U21311 (N_21311,N_19852,N_18263);
nand U21312 (N_21312,N_19089,N_19839);
xnor U21313 (N_21313,N_19121,N_18989);
or U21314 (N_21314,N_18639,N_18999);
nor U21315 (N_21315,N_19476,N_19130);
nor U21316 (N_21316,N_19093,N_18850);
nand U21317 (N_21317,N_18320,N_18103);
xor U21318 (N_21318,N_18076,N_18813);
nand U21319 (N_21319,N_19119,N_19681);
nand U21320 (N_21320,N_18497,N_19144);
and U21321 (N_21321,N_18495,N_18067);
nand U21322 (N_21322,N_18624,N_19726);
or U21323 (N_21323,N_19040,N_19263);
or U21324 (N_21324,N_19877,N_18595);
xor U21325 (N_21325,N_19322,N_19520);
or U21326 (N_21326,N_18065,N_19091);
nand U21327 (N_21327,N_18318,N_19530);
nor U21328 (N_21328,N_18143,N_19364);
nor U21329 (N_21329,N_19060,N_18845);
and U21330 (N_21330,N_19413,N_18179);
nor U21331 (N_21331,N_19602,N_18812);
and U21332 (N_21332,N_18971,N_18590);
or U21333 (N_21333,N_18446,N_18113);
nand U21334 (N_21334,N_18592,N_19190);
and U21335 (N_21335,N_19451,N_19722);
nor U21336 (N_21336,N_19289,N_18412);
xnor U21337 (N_21337,N_18405,N_19105);
xor U21338 (N_21338,N_19409,N_19384);
or U21339 (N_21339,N_18622,N_19195);
and U21340 (N_21340,N_19096,N_18717);
nand U21341 (N_21341,N_19397,N_18659);
or U21342 (N_21342,N_18905,N_19135);
nand U21343 (N_21343,N_19998,N_18347);
and U21344 (N_21344,N_18348,N_18047);
nor U21345 (N_21345,N_19104,N_19788);
nand U21346 (N_21346,N_18668,N_18605);
and U21347 (N_21347,N_18729,N_18494);
and U21348 (N_21348,N_19328,N_18788);
or U21349 (N_21349,N_19575,N_18334);
nor U21350 (N_21350,N_18862,N_18208);
or U21351 (N_21351,N_19954,N_18160);
xnor U21352 (N_21352,N_19793,N_19424);
nand U21353 (N_21353,N_18902,N_18593);
xor U21354 (N_21354,N_18942,N_18517);
or U21355 (N_21355,N_18959,N_19432);
and U21356 (N_21356,N_19418,N_19493);
and U21357 (N_21357,N_18046,N_19097);
and U21358 (N_21358,N_18872,N_18137);
and U21359 (N_21359,N_19340,N_18428);
and U21360 (N_21360,N_18254,N_19952);
xnor U21361 (N_21361,N_18018,N_19374);
and U21362 (N_21362,N_18360,N_18351);
nor U21363 (N_21363,N_19668,N_18328);
xor U21364 (N_21364,N_18108,N_18131);
xor U21365 (N_21365,N_19774,N_19336);
or U21366 (N_21366,N_18045,N_18971);
nand U21367 (N_21367,N_18893,N_18540);
nor U21368 (N_21368,N_19717,N_18097);
nand U21369 (N_21369,N_19177,N_18028);
or U21370 (N_21370,N_19062,N_19786);
or U21371 (N_21371,N_18048,N_18826);
and U21372 (N_21372,N_18069,N_19259);
nor U21373 (N_21373,N_18747,N_19509);
nor U21374 (N_21374,N_19254,N_18440);
or U21375 (N_21375,N_18304,N_19515);
and U21376 (N_21376,N_18145,N_19410);
nand U21377 (N_21377,N_19903,N_18373);
nand U21378 (N_21378,N_18191,N_19584);
and U21379 (N_21379,N_18297,N_19748);
or U21380 (N_21380,N_19134,N_18237);
nand U21381 (N_21381,N_18164,N_19240);
and U21382 (N_21382,N_18436,N_19776);
xnor U21383 (N_21383,N_18566,N_18719);
nand U21384 (N_21384,N_18438,N_18090);
nand U21385 (N_21385,N_19041,N_19011);
and U21386 (N_21386,N_18955,N_19852);
and U21387 (N_21387,N_19213,N_19760);
nor U21388 (N_21388,N_19683,N_19215);
nand U21389 (N_21389,N_19180,N_18678);
xor U21390 (N_21390,N_19465,N_19305);
or U21391 (N_21391,N_19651,N_19726);
nor U21392 (N_21392,N_19058,N_18091);
nor U21393 (N_21393,N_18471,N_18941);
nand U21394 (N_21394,N_18004,N_19704);
and U21395 (N_21395,N_18284,N_19516);
or U21396 (N_21396,N_18377,N_19751);
nand U21397 (N_21397,N_18042,N_18825);
nor U21398 (N_21398,N_18713,N_18095);
nor U21399 (N_21399,N_19583,N_18461);
nor U21400 (N_21400,N_19400,N_19237);
and U21401 (N_21401,N_18449,N_18164);
nor U21402 (N_21402,N_19973,N_19411);
or U21403 (N_21403,N_18961,N_18375);
and U21404 (N_21404,N_18558,N_18775);
and U21405 (N_21405,N_18101,N_19181);
and U21406 (N_21406,N_19667,N_18781);
nand U21407 (N_21407,N_19252,N_19006);
xor U21408 (N_21408,N_18679,N_18725);
xnor U21409 (N_21409,N_19169,N_19381);
nand U21410 (N_21410,N_19279,N_19327);
and U21411 (N_21411,N_18753,N_18132);
or U21412 (N_21412,N_19577,N_19819);
nand U21413 (N_21413,N_18534,N_18871);
nand U21414 (N_21414,N_18068,N_19764);
xnor U21415 (N_21415,N_19345,N_18296);
nand U21416 (N_21416,N_18271,N_18901);
and U21417 (N_21417,N_18976,N_18427);
nor U21418 (N_21418,N_18494,N_19514);
xnor U21419 (N_21419,N_18518,N_18979);
or U21420 (N_21420,N_19974,N_19958);
xnor U21421 (N_21421,N_18926,N_18254);
nand U21422 (N_21422,N_19324,N_18231);
or U21423 (N_21423,N_18707,N_18177);
xnor U21424 (N_21424,N_19590,N_18278);
nor U21425 (N_21425,N_19119,N_19648);
xor U21426 (N_21426,N_18916,N_19159);
xor U21427 (N_21427,N_19883,N_19689);
nand U21428 (N_21428,N_18540,N_19893);
and U21429 (N_21429,N_18798,N_18061);
or U21430 (N_21430,N_18161,N_19361);
nor U21431 (N_21431,N_19917,N_19100);
and U21432 (N_21432,N_18125,N_18077);
nor U21433 (N_21433,N_18530,N_19840);
nand U21434 (N_21434,N_19451,N_18171);
or U21435 (N_21435,N_19963,N_19010);
xor U21436 (N_21436,N_19521,N_18783);
nand U21437 (N_21437,N_19436,N_19535);
and U21438 (N_21438,N_18509,N_19685);
xor U21439 (N_21439,N_19959,N_19677);
nand U21440 (N_21440,N_19683,N_19431);
xnor U21441 (N_21441,N_19405,N_19091);
nor U21442 (N_21442,N_19167,N_19779);
and U21443 (N_21443,N_19454,N_19352);
nor U21444 (N_21444,N_18943,N_18482);
nor U21445 (N_21445,N_19424,N_19999);
and U21446 (N_21446,N_19831,N_19944);
nand U21447 (N_21447,N_19301,N_19626);
nor U21448 (N_21448,N_18157,N_18179);
or U21449 (N_21449,N_19543,N_18120);
nand U21450 (N_21450,N_19960,N_18595);
and U21451 (N_21451,N_18782,N_19607);
nor U21452 (N_21452,N_18685,N_18702);
nor U21453 (N_21453,N_19974,N_18030);
nor U21454 (N_21454,N_18053,N_18560);
or U21455 (N_21455,N_18396,N_18924);
nor U21456 (N_21456,N_19772,N_19037);
or U21457 (N_21457,N_18411,N_18174);
xor U21458 (N_21458,N_18584,N_18215);
nor U21459 (N_21459,N_18874,N_19327);
and U21460 (N_21460,N_19003,N_18126);
and U21461 (N_21461,N_18675,N_18741);
nor U21462 (N_21462,N_18236,N_18645);
xnor U21463 (N_21463,N_19062,N_19982);
nor U21464 (N_21464,N_19477,N_19706);
xnor U21465 (N_21465,N_19385,N_19824);
nand U21466 (N_21466,N_19787,N_18020);
and U21467 (N_21467,N_18845,N_19325);
nor U21468 (N_21468,N_18338,N_19297);
nor U21469 (N_21469,N_18306,N_19768);
xnor U21470 (N_21470,N_19834,N_18432);
and U21471 (N_21471,N_18685,N_18152);
xnor U21472 (N_21472,N_18387,N_19621);
and U21473 (N_21473,N_18085,N_19166);
and U21474 (N_21474,N_18536,N_18159);
nand U21475 (N_21475,N_18344,N_18973);
or U21476 (N_21476,N_18672,N_18601);
nand U21477 (N_21477,N_19330,N_19335);
and U21478 (N_21478,N_18262,N_18828);
and U21479 (N_21479,N_19225,N_18925);
nor U21480 (N_21480,N_19011,N_18867);
nand U21481 (N_21481,N_18625,N_19562);
nor U21482 (N_21482,N_18726,N_18633);
or U21483 (N_21483,N_19045,N_19072);
or U21484 (N_21484,N_18567,N_19272);
xor U21485 (N_21485,N_18807,N_19094);
nand U21486 (N_21486,N_18425,N_18837);
xnor U21487 (N_21487,N_18356,N_18002);
or U21488 (N_21488,N_19933,N_19538);
nand U21489 (N_21489,N_19791,N_18489);
or U21490 (N_21490,N_18989,N_18890);
xnor U21491 (N_21491,N_18883,N_19117);
xnor U21492 (N_21492,N_19342,N_18295);
or U21493 (N_21493,N_18901,N_18196);
xnor U21494 (N_21494,N_18808,N_19995);
or U21495 (N_21495,N_19862,N_18440);
or U21496 (N_21496,N_19746,N_18347);
or U21497 (N_21497,N_18424,N_18977);
or U21498 (N_21498,N_19341,N_19560);
nor U21499 (N_21499,N_19278,N_19632);
xor U21500 (N_21500,N_19001,N_18651);
and U21501 (N_21501,N_18964,N_19392);
xnor U21502 (N_21502,N_19767,N_19687);
or U21503 (N_21503,N_18461,N_19801);
and U21504 (N_21504,N_19411,N_19409);
or U21505 (N_21505,N_18922,N_18227);
nor U21506 (N_21506,N_18955,N_18677);
or U21507 (N_21507,N_19249,N_19718);
and U21508 (N_21508,N_19455,N_19999);
or U21509 (N_21509,N_19646,N_19598);
xor U21510 (N_21510,N_18193,N_18005);
and U21511 (N_21511,N_18234,N_18723);
or U21512 (N_21512,N_19502,N_18368);
nand U21513 (N_21513,N_19460,N_18219);
and U21514 (N_21514,N_18990,N_18908);
nor U21515 (N_21515,N_19375,N_18591);
or U21516 (N_21516,N_18572,N_18642);
and U21517 (N_21517,N_18575,N_19830);
xnor U21518 (N_21518,N_18576,N_19140);
xor U21519 (N_21519,N_18297,N_18830);
nand U21520 (N_21520,N_19997,N_18652);
and U21521 (N_21521,N_18329,N_18628);
nand U21522 (N_21522,N_19021,N_19845);
and U21523 (N_21523,N_19633,N_18048);
nor U21524 (N_21524,N_18334,N_19151);
xor U21525 (N_21525,N_18329,N_19341);
nor U21526 (N_21526,N_18946,N_18111);
nor U21527 (N_21527,N_19511,N_18664);
or U21528 (N_21528,N_18267,N_18230);
nor U21529 (N_21529,N_18850,N_18031);
or U21530 (N_21530,N_19577,N_18727);
or U21531 (N_21531,N_18007,N_19811);
nor U21532 (N_21532,N_19879,N_19982);
nand U21533 (N_21533,N_18513,N_18259);
xnor U21534 (N_21534,N_18381,N_19073);
and U21535 (N_21535,N_19441,N_19897);
nand U21536 (N_21536,N_19007,N_19439);
nand U21537 (N_21537,N_18718,N_19775);
and U21538 (N_21538,N_19045,N_18743);
nor U21539 (N_21539,N_19215,N_19373);
or U21540 (N_21540,N_19922,N_19952);
and U21541 (N_21541,N_19659,N_18778);
nor U21542 (N_21542,N_19985,N_19939);
nand U21543 (N_21543,N_19196,N_19082);
xnor U21544 (N_21544,N_18443,N_18326);
nor U21545 (N_21545,N_18836,N_18895);
nor U21546 (N_21546,N_18339,N_19865);
nand U21547 (N_21547,N_19671,N_19858);
xnor U21548 (N_21548,N_18264,N_19484);
nor U21549 (N_21549,N_19330,N_18909);
or U21550 (N_21550,N_19521,N_19515);
nor U21551 (N_21551,N_19545,N_19460);
or U21552 (N_21552,N_18124,N_18305);
or U21553 (N_21553,N_19716,N_18179);
nor U21554 (N_21554,N_19512,N_18136);
xnor U21555 (N_21555,N_18700,N_19436);
nand U21556 (N_21556,N_19209,N_18964);
xor U21557 (N_21557,N_18781,N_18159);
xor U21558 (N_21558,N_18553,N_18374);
nor U21559 (N_21559,N_19143,N_19222);
xnor U21560 (N_21560,N_19397,N_19119);
nor U21561 (N_21561,N_19899,N_18929);
nand U21562 (N_21562,N_18296,N_18574);
or U21563 (N_21563,N_19502,N_19462);
xnor U21564 (N_21564,N_19483,N_19395);
nand U21565 (N_21565,N_19860,N_19565);
xor U21566 (N_21566,N_19018,N_19822);
and U21567 (N_21567,N_19990,N_19226);
xor U21568 (N_21568,N_19847,N_18766);
xor U21569 (N_21569,N_18131,N_19326);
nor U21570 (N_21570,N_19966,N_19384);
xor U21571 (N_21571,N_19393,N_18629);
or U21572 (N_21572,N_19008,N_18691);
and U21573 (N_21573,N_19281,N_19730);
nor U21574 (N_21574,N_19776,N_18100);
and U21575 (N_21575,N_18770,N_18174);
or U21576 (N_21576,N_18142,N_18582);
or U21577 (N_21577,N_18978,N_19164);
or U21578 (N_21578,N_18589,N_18945);
xnor U21579 (N_21579,N_19720,N_18460);
or U21580 (N_21580,N_18687,N_18146);
nand U21581 (N_21581,N_18958,N_19889);
nand U21582 (N_21582,N_18851,N_18428);
nand U21583 (N_21583,N_18786,N_19839);
or U21584 (N_21584,N_18881,N_19869);
or U21585 (N_21585,N_19512,N_19097);
and U21586 (N_21586,N_18730,N_18918);
nand U21587 (N_21587,N_18945,N_18443);
nand U21588 (N_21588,N_19235,N_19488);
or U21589 (N_21589,N_19644,N_18460);
nand U21590 (N_21590,N_18033,N_18046);
and U21591 (N_21591,N_19831,N_19991);
nand U21592 (N_21592,N_18396,N_19076);
or U21593 (N_21593,N_19862,N_18858);
nor U21594 (N_21594,N_19568,N_18699);
and U21595 (N_21595,N_19659,N_18518);
xnor U21596 (N_21596,N_18180,N_19584);
xor U21597 (N_21597,N_18451,N_19381);
and U21598 (N_21598,N_19026,N_18922);
xor U21599 (N_21599,N_18710,N_19196);
nand U21600 (N_21600,N_18319,N_19806);
nand U21601 (N_21601,N_19413,N_18814);
nand U21602 (N_21602,N_18968,N_19973);
nand U21603 (N_21603,N_19207,N_19676);
nor U21604 (N_21604,N_19230,N_18804);
nand U21605 (N_21605,N_19148,N_18579);
nand U21606 (N_21606,N_18592,N_18166);
nor U21607 (N_21607,N_18078,N_18537);
or U21608 (N_21608,N_19839,N_18714);
xor U21609 (N_21609,N_18739,N_19134);
nand U21610 (N_21610,N_19334,N_19777);
nand U21611 (N_21611,N_19672,N_18732);
or U21612 (N_21612,N_19694,N_19649);
nor U21613 (N_21613,N_19376,N_18060);
nand U21614 (N_21614,N_18787,N_18212);
nand U21615 (N_21615,N_18650,N_19594);
nand U21616 (N_21616,N_19493,N_18724);
xnor U21617 (N_21617,N_18795,N_18530);
nor U21618 (N_21618,N_18257,N_18941);
nand U21619 (N_21619,N_18173,N_19538);
nor U21620 (N_21620,N_18201,N_19718);
and U21621 (N_21621,N_18486,N_18255);
nand U21622 (N_21622,N_18316,N_18533);
xor U21623 (N_21623,N_18044,N_19554);
nand U21624 (N_21624,N_19932,N_18384);
nor U21625 (N_21625,N_19886,N_18858);
xor U21626 (N_21626,N_18030,N_18613);
nor U21627 (N_21627,N_19743,N_19681);
and U21628 (N_21628,N_18739,N_18797);
nand U21629 (N_21629,N_19821,N_18394);
and U21630 (N_21630,N_19729,N_19358);
nor U21631 (N_21631,N_19007,N_19395);
xnor U21632 (N_21632,N_18749,N_18190);
xnor U21633 (N_21633,N_19642,N_19147);
nand U21634 (N_21634,N_19579,N_18547);
xnor U21635 (N_21635,N_19469,N_19942);
nand U21636 (N_21636,N_19805,N_18955);
nand U21637 (N_21637,N_18783,N_19477);
or U21638 (N_21638,N_18223,N_18321);
or U21639 (N_21639,N_19222,N_18939);
xor U21640 (N_21640,N_19863,N_18473);
and U21641 (N_21641,N_19603,N_19018);
nor U21642 (N_21642,N_18856,N_19348);
or U21643 (N_21643,N_19791,N_19096);
or U21644 (N_21644,N_18442,N_18042);
nand U21645 (N_21645,N_19383,N_18764);
and U21646 (N_21646,N_19936,N_18369);
xnor U21647 (N_21647,N_18503,N_18907);
or U21648 (N_21648,N_19510,N_19245);
xor U21649 (N_21649,N_19757,N_18500);
nand U21650 (N_21650,N_19154,N_18165);
xnor U21651 (N_21651,N_19555,N_18014);
xnor U21652 (N_21652,N_18355,N_19517);
or U21653 (N_21653,N_18744,N_19783);
nor U21654 (N_21654,N_19578,N_18265);
xor U21655 (N_21655,N_19603,N_18395);
nor U21656 (N_21656,N_18216,N_19340);
and U21657 (N_21657,N_18418,N_19175);
nor U21658 (N_21658,N_18997,N_19978);
or U21659 (N_21659,N_19548,N_19785);
nor U21660 (N_21660,N_18015,N_19814);
nor U21661 (N_21661,N_19639,N_18038);
nor U21662 (N_21662,N_19069,N_18014);
and U21663 (N_21663,N_19807,N_18921);
nor U21664 (N_21664,N_19588,N_19005);
and U21665 (N_21665,N_18908,N_19571);
or U21666 (N_21666,N_18659,N_19926);
nand U21667 (N_21667,N_18745,N_19614);
or U21668 (N_21668,N_18371,N_19303);
or U21669 (N_21669,N_19263,N_19031);
nor U21670 (N_21670,N_18169,N_19877);
xnor U21671 (N_21671,N_19674,N_19870);
xnor U21672 (N_21672,N_18728,N_18008);
and U21673 (N_21673,N_18307,N_18763);
and U21674 (N_21674,N_19885,N_18205);
and U21675 (N_21675,N_19768,N_19416);
and U21676 (N_21676,N_19594,N_18744);
nor U21677 (N_21677,N_18198,N_19157);
or U21678 (N_21678,N_19190,N_18112);
and U21679 (N_21679,N_18212,N_19768);
and U21680 (N_21680,N_19160,N_18284);
xor U21681 (N_21681,N_19927,N_18544);
and U21682 (N_21682,N_18881,N_19012);
nand U21683 (N_21683,N_18288,N_19736);
or U21684 (N_21684,N_19197,N_19509);
nand U21685 (N_21685,N_18317,N_19821);
and U21686 (N_21686,N_19217,N_19410);
xnor U21687 (N_21687,N_18751,N_19925);
xnor U21688 (N_21688,N_18272,N_19046);
nand U21689 (N_21689,N_19830,N_19715);
xnor U21690 (N_21690,N_19827,N_18751);
nand U21691 (N_21691,N_18741,N_19964);
nor U21692 (N_21692,N_18601,N_19467);
nor U21693 (N_21693,N_18759,N_19225);
and U21694 (N_21694,N_19911,N_18863);
or U21695 (N_21695,N_19294,N_19690);
xor U21696 (N_21696,N_18318,N_18913);
and U21697 (N_21697,N_18461,N_19188);
nor U21698 (N_21698,N_19332,N_18869);
nor U21699 (N_21699,N_18652,N_19024);
nand U21700 (N_21700,N_19600,N_18787);
nor U21701 (N_21701,N_19392,N_19902);
xnor U21702 (N_21702,N_19841,N_18872);
nand U21703 (N_21703,N_18702,N_19451);
and U21704 (N_21704,N_18651,N_19544);
nand U21705 (N_21705,N_18708,N_19451);
or U21706 (N_21706,N_19679,N_19451);
nor U21707 (N_21707,N_18869,N_18274);
nand U21708 (N_21708,N_18484,N_19835);
nor U21709 (N_21709,N_19001,N_19671);
nand U21710 (N_21710,N_19899,N_19894);
and U21711 (N_21711,N_18257,N_18948);
or U21712 (N_21712,N_18595,N_19000);
xor U21713 (N_21713,N_18331,N_18096);
nor U21714 (N_21714,N_19412,N_18411);
nor U21715 (N_21715,N_18421,N_18825);
or U21716 (N_21716,N_19203,N_18523);
and U21717 (N_21717,N_18295,N_18180);
or U21718 (N_21718,N_18313,N_19900);
and U21719 (N_21719,N_18870,N_19324);
or U21720 (N_21720,N_19591,N_19052);
nand U21721 (N_21721,N_18734,N_18772);
nand U21722 (N_21722,N_18161,N_18890);
or U21723 (N_21723,N_19901,N_19178);
xnor U21724 (N_21724,N_18707,N_18284);
and U21725 (N_21725,N_18058,N_19754);
or U21726 (N_21726,N_19422,N_19995);
or U21727 (N_21727,N_19410,N_18872);
nand U21728 (N_21728,N_18293,N_18252);
or U21729 (N_21729,N_19261,N_18147);
nand U21730 (N_21730,N_18502,N_19737);
xor U21731 (N_21731,N_19961,N_18256);
nor U21732 (N_21732,N_18963,N_19852);
nor U21733 (N_21733,N_18993,N_18132);
nor U21734 (N_21734,N_19062,N_19807);
nor U21735 (N_21735,N_19171,N_19012);
nor U21736 (N_21736,N_19190,N_19832);
nand U21737 (N_21737,N_19907,N_18356);
nor U21738 (N_21738,N_18926,N_19684);
and U21739 (N_21739,N_18322,N_19179);
and U21740 (N_21740,N_19703,N_19571);
nand U21741 (N_21741,N_18477,N_19685);
and U21742 (N_21742,N_18721,N_19061);
and U21743 (N_21743,N_19018,N_19891);
nand U21744 (N_21744,N_18716,N_19488);
nand U21745 (N_21745,N_19232,N_19091);
xnor U21746 (N_21746,N_19372,N_18049);
or U21747 (N_21747,N_18905,N_19393);
nand U21748 (N_21748,N_19428,N_18074);
nor U21749 (N_21749,N_18521,N_18328);
and U21750 (N_21750,N_18382,N_19595);
or U21751 (N_21751,N_18576,N_18164);
nor U21752 (N_21752,N_19174,N_19651);
nand U21753 (N_21753,N_19620,N_19567);
nor U21754 (N_21754,N_18086,N_18709);
xnor U21755 (N_21755,N_18560,N_19618);
nand U21756 (N_21756,N_18224,N_18340);
nor U21757 (N_21757,N_19332,N_19457);
nand U21758 (N_21758,N_19492,N_19010);
nand U21759 (N_21759,N_19052,N_19835);
nor U21760 (N_21760,N_19448,N_18420);
and U21761 (N_21761,N_18766,N_18353);
or U21762 (N_21762,N_18691,N_18705);
or U21763 (N_21763,N_18495,N_19632);
or U21764 (N_21764,N_18858,N_19547);
xor U21765 (N_21765,N_18551,N_19675);
xnor U21766 (N_21766,N_18701,N_18202);
or U21767 (N_21767,N_18199,N_19062);
nor U21768 (N_21768,N_19613,N_19810);
nor U21769 (N_21769,N_19554,N_18390);
nor U21770 (N_21770,N_18211,N_18810);
and U21771 (N_21771,N_18182,N_19441);
nor U21772 (N_21772,N_19873,N_19502);
and U21773 (N_21773,N_19511,N_19290);
nand U21774 (N_21774,N_18717,N_18285);
xor U21775 (N_21775,N_19871,N_19146);
nand U21776 (N_21776,N_18204,N_19988);
and U21777 (N_21777,N_18080,N_19277);
and U21778 (N_21778,N_19338,N_18232);
nor U21779 (N_21779,N_18056,N_19420);
or U21780 (N_21780,N_18730,N_18948);
nand U21781 (N_21781,N_19560,N_19767);
nor U21782 (N_21782,N_19990,N_19244);
nand U21783 (N_21783,N_18956,N_19675);
or U21784 (N_21784,N_18918,N_18184);
nor U21785 (N_21785,N_18563,N_19808);
xnor U21786 (N_21786,N_19217,N_18154);
or U21787 (N_21787,N_19874,N_19115);
xor U21788 (N_21788,N_18333,N_19787);
nand U21789 (N_21789,N_19846,N_19115);
nand U21790 (N_21790,N_18131,N_18431);
or U21791 (N_21791,N_18258,N_19359);
nor U21792 (N_21792,N_18469,N_18944);
or U21793 (N_21793,N_18248,N_18950);
and U21794 (N_21794,N_18408,N_18765);
and U21795 (N_21795,N_18644,N_19724);
nand U21796 (N_21796,N_19452,N_19295);
xnor U21797 (N_21797,N_18593,N_19015);
or U21798 (N_21798,N_18690,N_19522);
nor U21799 (N_21799,N_19250,N_18772);
or U21800 (N_21800,N_18170,N_19122);
xnor U21801 (N_21801,N_19711,N_19029);
nor U21802 (N_21802,N_19536,N_18336);
nand U21803 (N_21803,N_18190,N_18731);
nand U21804 (N_21804,N_19193,N_19008);
and U21805 (N_21805,N_18490,N_19491);
nand U21806 (N_21806,N_18358,N_18826);
and U21807 (N_21807,N_19547,N_18324);
nand U21808 (N_21808,N_19263,N_18610);
nor U21809 (N_21809,N_18272,N_18984);
xor U21810 (N_21810,N_18235,N_19994);
xnor U21811 (N_21811,N_18526,N_18248);
xor U21812 (N_21812,N_18499,N_19817);
nand U21813 (N_21813,N_19533,N_18181);
and U21814 (N_21814,N_19976,N_19492);
nor U21815 (N_21815,N_18099,N_19237);
and U21816 (N_21816,N_18532,N_19054);
xnor U21817 (N_21817,N_19709,N_18862);
and U21818 (N_21818,N_18688,N_18335);
and U21819 (N_21819,N_19426,N_19238);
and U21820 (N_21820,N_18655,N_18460);
nand U21821 (N_21821,N_19591,N_19225);
xnor U21822 (N_21822,N_19166,N_18000);
nand U21823 (N_21823,N_19018,N_19584);
nand U21824 (N_21824,N_18552,N_18896);
nand U21825 (N_21825,N_19772,N_18730);
nor U21826 (N_21826,N_18924,N_18470);
xor U21827 (N_21827,N_18001,N_19761);
nor U21828 (N_21828,N_19411,N_19953);
or U21829 (N_21829,N_18126,N_18868);
nand U21830 (N_21830,N_19249,N_18210);
or U21831 (N_21831,N_19552,N_19078);
and U21832 (N_21832,N_18439,N_19642);
xor U21833 (N_21833,N_18485,N_19223);
and U21834 (N_21834,N_19693,N_19406);
nor U21835 (N_21835,N_19435,N_19992);
or U21836 (N_21836,N_19553,N_19419);
nand U21837 (N_21837,N_19547,N_18139);
xnor U21838 (N_21838,N_18694,N_18669);
xnor U21839 (N_21839,N_19857,N_19187);
or U21840 (N_21840,N_18856,N_18811);
nor U21841 (N_21841,N_19808,N_19360);
nor U21842 (N_21842,N_19109,N_18598);
or U21843 (N_21843,N_18350,N_19277);
nand U21844 (N_21844,N_19502,N_19322);
nor U21845 (N_21845,N_19558,N_18311);
or U21846 (N_21846,N_18969,N_18290);
and U21847 (N_21847,N_18556,N_18002);
and U21848 (N_21848,N_18973,N_18926);
nand U21849 (N_21849,N_19741,N_19582);
xor U21850 (N_21850,N_19243,N_19832);
xnor U21851 (N_21851,N_18478,N_19710);
xor U21852 (N_21852,N_19715,N_19638);
xor U21853 (N_21853,N_19268,N_19482);
xor U21854 (N_21854,N_19656,N_19123);
xor U21855 (N_21855,N_18378,N_19102);
and U21856 (N_21856,N_18501,N_19744);
xnor U21857 (N_21857,N_19688,N_18052);
nor U21858 (N_21858,N_18105,N_19569);
nor U21859 (N_21859,N_18705,N_18207);
or U21860 (N_21860,N_19539,N_18759);
nor U21861 (N_21861,N_18734,N_19056);
or U21862 (N_21862,N_18155,N_18544);
and U21863 (N_21863,N_19909,N_18701);
or U21864 (N_21864,N_18930,N_18181);
xnor U21865 (N_21865,N_18309,N_18547);
nand U21866 (N_21866,N_18765,N_18763);
and U21867 (N_21867,N_18939,N_19080);
nand U21868 (N_21868,N_19520,N_19685);
xor U21869 (N_21869,N_19090,N_19249);
and U21870 (N_21870,N_19469,N_19781);
xnor U21871 (N_21871,N_18834,N_18581);
or U21872 (N_21872,N_19494,N_18971);
nor U21873 (N_21873,N_18111,N_18585);
nand U21874 (N_21874,N_19324,N_18868);
nor U21875 (N_21875,N_19752,N_19072);
nor U21876 (N_21876,N_18579,N_18045);
and U21877 (N_21877,N_18619,N_18310);
nand U21878 (N_21878,N_18573,N_19064);
and U21879 (N_21879,N_18324,N_18691);
nor U21880 (N_21880,N_18858,N_18632);
or U21881 (N_21881,N_18285,N_18272);
xor U21882 (N_21882,N_19083,N_18999);
nand U21883 (N_21883,N_19224,N_19973);
nor U21884 (N_21884,N_18352,N_19271);
or U21885 (N_21885,N_18181,N_18731);
and U21886 (N_21886,N_19465,N_18101);
and U21887 (N_21887,N_18457,N_19008);
nand U21888 (N_21888,N_19348,N_19290);
xnor U21889 (N_21889,N_18061,N_19265);
and U21890 (N_21890,N_19872,N_19189);
nand U21891 (N_21891,N_19882,N_18081);
or U21892 (N_21892,N_18615,N_19259);
xnor U21893 (N_21893,N_19076,N_18316);
nand U21894 (N_21894,N_18883,N_19239);
nor U21895 (N_21895,N_18747,N_18370);
nor U21896 (N_21896,N_19794,N_18796);
or U21897 (N_21897,N_18680,N_18280);
and U21898 (N_21898,N_18993,N_19169);
nor U21899 (N_21899,N_19274,N_19144);
and U21900 (N_21900,N_18695,N_18875);
or U21901 (N_21901,N_18210,N_18729);
nand U21902 (N_21902,N_18951,N_18357);
xnor U21903 (N_21903,N_18347,N_19320);
and U21904 (N_21904,N_19331,N_19367);
or U21905 (N_21905,N_19649,N_19399);
or U21906 (N_21906,N_19472,N_18496);
or U21907 (N_21907,N_18203,N_19042);
nand U21908 (N_21908,N_18071,N_19459);
nand U21909 (N_21909,N_18807,N_18838);
or U21910 (N_21910,N_18785,N_18166);
or U21911 (N_21911,N_18245,N_18102);
and U21912 (N_21912,N_18564,N_19368);
nor U21913 (N_21913,N_18112,N_18592);
and U21914 (N_21914,N_18025,N_19708);
nor U21915 (N_21915,N_19600,N_18394);
xnor U21916 (N_21916,N_19823,N_18903);
xor U21917 (N_21917,N_19102,N_18563);
nor U21918 (N_21918,N_19207,N_19151);
or U21919 (N_21919,N_19228,N_19435);
or U21920 (N_21920,N_18012,N_19732);
xnor U21921 (N_21921,N_18547,N_18448);
nand U21922 (N_21922,N_18947,N_19493);
nand U21923 (N_21923,N_19397,N_19172);
nand U21924 (N_21924,N_19411,N_19568);
nor U21925 (N_21925,N_19333,N_19087);
and U21926 (N_21926,N_18007,N_18567);
or U21927 (N_21927,N_18375,N_19587);
and U21928 (N_21928,N_19412,N_18485);
or U21929 (N_21929,N_19646,N_19010);
or U21930 (N_21930,N_18173,N_19701);
nor U21931 (N_21931,N_18243,N_18456);
nor U21932 (N_21932,N_19000,N_18381);
nor U21933 (N_21933,N_19336,N_19793);
or U21934 (N_21934,N_18965,N_18831);
and U21935 (N_21935,N_18800,N_18286);
nor U21936 (N_21936,N_19075,N_19249);
and U21937 (N_21937,N_19191,N_18479);
or U21938 (N_21938,N_18542,N_19035);
nand U21939 (N_21939,N_18735,N_19337);
nand U21940 (N_21940,N_19323,N_18296);
xor U21941 (N_21941,N_18061,N_19103);
xor U21942 (N_21942,N_18821,N_19741);
or U21943 (N_21943,N_19193,N_19699);
or U21944 (N_21944,N_18200,N_19668);
nand U21945 (N_21945,N_18454,N_19084);
xnor U21946 (N_21946,N_19700,N_18889);
or U21947 (N_21947,N_18502,N_19406);
nand U21948 (N_21948,N_18256,N_18604);
xnor U21949 (N_21949,N_18624,N_18110);
and U21950 (N_21950,N_18581,N_19710);
nor U21951 (N_21951,N_19618,N_18546);
xor U21952 (N_21952,N_18896,N_18946);
nor U21953 (N_21953,N_19223,N_19568);
and U21954 (N_21954,N_18490,N_19131);
or U21955 (N_21955,N_19392,N_18723);
nor U21956 (N_21956,N_18760,N_19364);
nor U21957 (N_21957,N_18304,N_19775);
nand U21958 (N_21958,N_18982,N_18523);
and U21959 (N_21959,N_18600,N_18608);
nor U21960 (N_21960,N_19695,N_19794);
nor U21961 (N_21961,N_18486,N_19081);
nand U21962 (N_21962,N_19246,N_18481);
or U21963 (N_21963,N_19014,N_19831);
xor U21964 (N_21964,N_18538,N_19418);
nor U21965 (N_21965,N_18254,N_19414);
nor U21966 (N_21966,N_19125,N_18728);
nor U21967 (N_21967,N_19009,N_18627);
or U21968 (N_21968,N_19809,N_19243);
xnor U21969 (N_21969,N_19443,N_18812);
and U21970 (N_21970,N_19217,N_18511);
nand U21971 (N_21971,N_19871,N_19669);
and U21972 (N_21972,N_19441,N_19082);
and U21973 (N_21973,N_18066,N_19989);
xor U21974 (N_21974,N_18894,N_19050);
nand U21975 (N_21975,N_19408,N_18031);
and U21976 (N_21976,N_19248,N_18769);
xnor U21977 (N_21977,N_18745,N_18039);
nor U21978 (N_21978,N_18618,N_18118);
and U21979 (N_21979,N_19987,N_19175);
nor U21980 (N_21980,N_19551,N_19038);
nand U21981 (N_21981,N_19933,N_19765);
nand U21982 (N_21982,N_19057,N_18304);
nand U21983 (N_21983,N_18520,N_19865);
xnor U21984 (N_21984,N_19308,N_18656);
or U21985 (N_21985,N_19818,N_19540);
nand U21986 (N_21986,N_19601,N_18370);
or U21987 (N_21987,N_19903,N_18479);
xnor U21988 (N_21988,N_18564,N_18425);
nor U21989 (N_21989,N_18132,N_19730);
or U21990 (N_21990,N_19287,N_19536);
and U21991 (N_21991,N_18571,N_18108);
xor U21992 (N_21992,N_19177,N_18165);
nor U21993 (N_21993,N_18554,N_18734);
nor U21994 (N_21994,N_18817,N_19588);
nor U21995 (N_21995,N_18980,N_19944);
nor U21996 (N_21996,N_18949,N_18257);
or U21997 (N_21997,N_18891,N_19424);
nor U21998 (N_21998,N_19957,N_19000);
and U21999 (N_21999,N_19541,N_18310);
nand U22000 (N_22000,N_21320,N_20394);
xor U22001 (N_22001,N_20665,N_20721);
or U22002 (N_22002,N_21685,N_20158);
nor U22003 (N_22003,N_20635,N_21105);
nor U22004 (N_22004,N_20609,N_20051);
or U22005 (N_22005,N_20432,N_21138);
and U22006 (N_22006,N_21281,N_21327);
or U22007 (N_22007,N_21280,N_20666);
nor U22008 (N_22008,N_20826,N_21383);
or U22009 (N_22009,N_20496,N_21227);
xor U22010 (N_22010,N_20195,N_21788);
nor U22011 (N_22011,N_20361,N_20799);
and U22012 (N_22012,N_20524,N_21220);
nand U22013 (N_22013,N_20773,N_20723);
xor U22014 (N_22014,N_20904,N_20812);
or U22015 (N_22015,N_21405,N_21576);
or U22016 (N_22016,N_20208,N_20276);
xnor U22017 (N_22017,N_20518,N_21474);
nor U22018 (N_22018,N_21987,N_20235);
nand U22019 (N_22019,N_21619,N_20820);
nor U22020 (N_22020,N_21560,N_20214);
and U22021 (N_22021,N_21497,N_20460);
xor U22022 (N_22022,N_21449,N_21346);
and U22023 (N_22023,N_21007,N_21000);
nor U22024 (N_22024,N_20996,N_20210);
or U22025 (N_22025,N_21230,N_20819);
xor U22026 (N_22026,N_21574,N_21924);
and U22027 (N_22027,N_21568,N_21855);
nand U22028 (N_22028,N_20964,N_21659);
nor U22029 (N_22029,N_21056,N_20308);
xor U22030 (N_22030,N_20075,N_21693);
or U22031 (N_22031,N_21861,N_20171);
nand U22032 (N_22032,N_21225,N_21233);
and U22033 (N_22033,N_21178,N_21340);
or U22034 (N_22034,N_21317,N_21650);
nor U22035 (N_22035,N_20226,N_21022);
xnor U22036 (N_22036,N_20835,N_21889);
xnor U22037 (N_22037,N_21587,N_21835);
nand U22038 (N_22038,N_20517,N_20753);
xnor U22039 (N_22039,N_20371,N_20786);
or U22040 (N_22040,N_20601,N_20804);
nand U22041 (N_22041,N_20341,N_21399);
nor U22042 (N_22042,N_20315,N_20652);
xnor U22043 (N_22043,N_20872,N_21442);
xnor U22044 (N_22044,N_21043,N_21503);
or U22045 (N_22045,N_21635,N_21342);
nor U22046 (N_22046,N_20752,N_21780);
and U22047 (N_22047,N_20718,N_20040);
xnor U22048 (N_22048,N_20623,N_20707);
xnor U22049 (N_22049,N_21535,N_20093);
nand U22050 (N_22050,N_20468,N_21100);
nor U22051 (N_22051,N_20574,N_21696);
and U22052 (N_22052,N_20270,N_20594);
nor U22053 (N_22053,N_20113,N_20547);
nand U22054 (N_22054,N_21931,N_21324);
or U22055 (N_22055,N_20245,N_21819);
xnor U22056 (N_22056,N_20381,N_20749);
nor U22057 (N_22057,N_20364,N_21948);
nand U22058 (N_22058,N_21637,N_21341);
or U22059 (N_22059,N_21168,N_20670);
or U22060 (N_22060,N_20626,N_20146);
xor U22061 (N_22061,N_20318,N_20661);
nand U22062 (N_22062,N_21212,N_20175);
nand U22063 (N_22063,N_20473,N_21257);
or U22064 (N_22064,N_21763,N_21395);
nor U22065 (N_22065,N_21925,N_20192);
nand U22066 (N_22066,N_21791,N_21407);
and U22067 (N_22067,N_21379,N_20454);
or U22068 (N_22068,N_21125,N_21837);
and U22069 (N_22069,N_20128,N_21963);
xnor U22070 (N_22070,N_21279,N_20023);
and U22071 (N_22071,N_21093,N_20005);
nor U22072 (N_22072,N_21103,N_20809);
nor U22073 (N_22073,N_20549,N_21027);
and U22074 (N_22074,N_20847,N_20922);
xor U22075 (N_22075,N_20448,N_21877);
nand U22076 (N_22076,N_21058,N_21081);
or U22077 (N_22077,N_20472,N_21588);
nand U22078 (N_22078,N_21648,N_21555);
xor U22079 (N_22079,N_20515,N_20330);
nor U22080 (N_22080,N_20566,N_21457);
and U22081 (N_22081,N_21228,N_21612);
and U22082 (N_22082,N_20926,N_20742);
xor U22083 (N_22083,N_21947,N_20941);
or U22084 (N_22084,N_21487,N_20933);
nand U22085 (N_22085,N_21695,N_21974);
xnor U22086 (N_22086,N_21831,N_21377);
nand U22087 (N_22087,N_21223,N_20047);
xor U22088 (N_22088,N_20359,N_21123);
and U22089 (N_22089,N_21332,N_20483);
xnor U22090 (N_22090,N_21301,N_20502);
nand U22091 (N_22091,N_21694,N_20862);
or U22092 (N_22092,N_21090,N_21372);
and U22093 (N_22093,N_20689,N_20015);
and U22094 (N_22094,N_20252,N_20519);
xnor U22095 (N_22095,N_20006,N_21794);
nand U22096 (N_22096,N_20918,N_20767);
nand U22097 (N_22097,N_20072,N_20376);
or U22098 (N_22098,N_20199,N_21864);
and U22099 (N_22099,N_20363,N_20266);
nand U22100 (N_22100,N_20755,N_21107);
and U22101 (N_22101,N_21716,N_21847);
and U22102 (N_22102,N_21381,N_20362);
nand U22103 (N_22103,N_21884,N_20928);
nor U22104 (N_22104,N_20054,N_20368);
and U22105 (N_22105,N_20938,N_21024);
and U22106 (N_22106,N_20043,N_21764);
nor U22107 (N_22107,N_21633,N_21744);
and U22108 (N_22108,N_21751,N_21786);
or U22109 (N_22109,N_21288,N_21293);
or U22110 (N_22110,N_20233,N_20818);
or U22111 (N_22111,N_20378,N_20148);
nor U22112 (N_22112,N_21718,N_21331);
nor U22113 (N_22113,N_21733,N_20232);
or U22114 (N_22114,N_20593,N_21537);
nand U22115 (N_22115,N_21185,N_21431);
or U22116 (N_22116,N_20372,N_21059);
or U22117 (N_22117,N_20281,N_21870);
nor U22118 (N_22118,N_21462,N_20781);
nand U22119 (N_22119,N_20296,N_21472);
or U22120 (N_22120,N_21805,N_20476);
xnor U22121 (N_22121,N_21708,N_20857);
nand U22122 (N_22122,N_21893,N_21964);
nor U22123 (N_22123,N_20414,N_20324);
nor U22124 (N_22124,N_20863,N_21008);
or U22125 (N_22125,N_20523,N_20614);
or U22126 (N_22126,N_20895,N_21769);
xnor U22127 (N_22127,N_20892,N_21486);
or U22128 (N_22128,N_21857,N_20706);
nor U22129 (N_22129,N_21760,N_21229);
and U22130 (N_22130,N_21358,N_21632);
or U22131 (N_22131,N_21347,N_21691);
xnor U22132 (N_22132,N_21810,N_20919);
nor U22133 (N_22133,N_21822,N_20693);
and U22134 (N_22134,N_20469,N_21993);
and U22135 (N_22135,N_20690,N_21130);
xnor U22136 (N_22136,N_21417,N_21552);
nor U22137 (N_22137,N_21839,N_21338);
and U22138 (N_22138,N_21018,N_20008);
or U22139 (N_22139,N_21912,N_21160);
nand U22140 (N_22140,N_20995,N_21918);
nand U22141 (N_22141,N_21600,N_20638);
or U22142 (N_22142,N_21894,N_21036);
nor U22143 (N_22143,N_21690,N_20772);
nor U22144 (N_22144,N_21732,N_21207);
nand U22145 (N_22145,N_20354,N_20189);
nor U22146 (N_22146,N_21531,N_21702);
and U22147 (N_22147,N_20708,N_20084);
nand U22148 (N_22148,N_21561,N_20916);
or U22149 (N_22149,N_20828,N_20866);
and U22150 (N_22150,N_21250,N_20878);
xnor U22151 (N_22151,N_20391,N_21887);
nand U22152 (N_22152,N_20177,N_20821);
nor U22153 (N_22153,N_20264,N_20736);
nand U22154 (N_22154,N_20420,N_20912);
xor U22155 (N_22155,N_20410,N_21583);
nor U22156 (N_22156,N_21916,N_21113);
and U22157 (N_22157,N_20568,N_21546);
nand U22158 (N_22158,N_21146,N_21570);
nor U22159 (N_22159,N_21674,N_21730);
nor U22160 (N_22160,N_21642,N_20145);
nand U22161 (N_22161,N_20747,N_20683);
nor U22162 (N_22162,N_20503,N_21011);
xor U22163 (N_22163,N_20358,N_20935);
xnor U22164 (N_22164,N_21832,N_21353);
and U22165 (N_22165,N_21269,N_20873);
or U22166 (N_22166,N_21796,N_21415);
nor U22167 (N_22167,N_20104,N_20312);
xor U22168 (N_22168,N_21958,N_20408);
or U22169 (N_22169,N_21823,N_21616);
nor U22170 (N_22170,N_21500,N_21048);
or U22171 (N_22171,N_20726,N_20830);
or U22172 (N_22172,N_21156,N_20013);
and U22173 (N_22173,N_20123,N_20196);
or U22174 (N_22174,N_21186,N_20621);
nor U22175 (N_22175,N_21840,N_20546);
xor U22176 (N_22176,N_21917,N_20012);
nor U22177 (N_22177,N_21014,N_20832);
nor U22178 (N_22178,N_20932,N_21858);
and U22179 (N_22179,N_20622,N_20393);
nand U22180 (N_22180,N_20882,N_21667);
nand U22181 (N_22181,N_20639,N_21554);
nor U22182 (N_22182,N_21152,N_21050);
xor U22183 (N_22183,N_21883,N_20495);
nor U22184 (N_22184,N_20314,N_21759);
and U22185 (N_22185,N_21770,N_21339);
or U22186 (N_22186,N_21793,N_21950);
or U22187 (N_22187,N_20944,N_20975);
nor U22188 (N_22188,N_21150,N_21905);
or U22189 (N_22189,N_21019,N_20852);
or U22190 (N_22190,N_20081,N_21191);
nand U22191 (N_22191,N_20778,N_21844);
or U22192 (N_22192,N_20466,N_20978);
nand U22193 (N_22193,N_20624,N_20530);
and U22194 (N_22194,N_20554,N_20541);
and U22195 (N_22195,N_20230,N_21393);
nand U22196 (N_22196,N_21362,N_21995);
xor U22197 (N_22197,N_21001,N_20389);
nand U22198 (N_22198,N_20610,N_21333);
or U22199 (N_22199,N_20717,N_21704);
or U22200 (N_22200,N_21971,N_21595);
xnor U22201 (N_22201,N_21656,N_21422);
or U22202 (N_22202,N_21491,N_20605);
and U22203 (N_22203,N_21128,N_21478);
nand U22204 (N_22204,N_20950,N_21663);
or U22205 (N_22205,N_21767,N_21578);
nand U22206 (N_22206,N_20691,N_20164);
xnor U22207 (N_22207,N_21041,N_21871);
or U22208 (N_22208,N_20563,N_20630);
and U22209 (N_22209,N_20029,N_20985);
and U22210 (N_22210,N_20141,N_20680);
nand U22211 (N_22211,N_20067,N_20289);
or U22212 (N_22212,N_21657,N_20887);
nor U22213 (N_22213,N_21376,N_20401);
and U22214 (N_22214,N_21412,N_20461);
nor U22215 (N_22215,N_21532,N_21572);
xnor U22216 (N_22216,N_20065,N_20556);
and U22217 (N_22217,N_21575,N_21458);
and U22218 (N_22218,N_21867,N_21030);
nor U22219 (N_22219,N_21804,N_20046);
xor U22220 (N_22220,N_20896,N_21444);
nand U22221 (N_22221,N_21611,N_20795);
or U22222 (N_22222,N_21569,N_21783);
nand U22223 (N_22223,N_20135,N_21741);
and U22224 (N_22224,N_21664,N_20567);
xnor U22225 (N_22225,N_21904,N_20322);
nand U22226 (N_22226,N_20783,N_21975);
nand U22227 (N_22227,N_21067,N_20026);
and U22228 (N_22228,N_20237,N_20740);
xnor U22229 (N_22229,N_21945,N_21826);
nand U22230 (N_22230,N_21304,N_20144);
nand U22231 (N_22231,N_21258,N_20422);
nand U22232 (N_22232,N_20036,N_21271);
nand U22233 (N_22233,N_21099,N_21721);
and U22234 (N_22234,N_21929,N_21647);
nand U22235 (N_22235,N_20894,N_21519);
or U22236 (N_22236,N_21521,N_21594);
nor U22237 (N_22237,N_21420,N_21003);
xor U22238 (N_22238,N_21498,N_21802);
xnor U22239 (N_22239,N_21911,N_20033);
or U22240 (N_22240,N_20038,N_21495);
nand U22241 (N_22241,N_20824,N_20434);
and U22242 (N_22242,N_21735,N_20679);
nor U22243 (N_22243,N_21455,N_21256);
nor U22244 (N_22244,N_21900,N_20790);
nor U22245 (N_22245,N_21179,N_20256);
xnor U22246 (N_22246,N_21678,N_21651);
nand U22247 (N_22247,N_20967,N_20599);
xnor U22248 (N_22248,N_20529,N_21591);
xor U22249 (N_22249,N_20577,N_21124);
nand U22250 (N_22250,N_21202,N_20475);
nand U22251 (N_22251,N_20711,N_20902);
and U22252 (N_22252,N_20842,N_21109);
xnor U22253 (N_22253,N_20240,N_21137);
and U22254 (N_22254,N_20991,N_20768);
xor U22255 (N_22255,N_21990,N_20152);
nor U22256 (N_22256,N_20987,N_21965);
and U22257 (N_22257,N_20265,N_21216);
or U22258 (N_22258,N_21969,N_21013);
nand U22259 (N_22259,N_21966,N_20485);
xor U22260 (N_22260,N_21687,N_20076);
or U22261 (N_22261,N_20989,N_20303);
nor U22262 (N_22262,N_21699,N_20027);
xor U22263 (N_22263,N_20032,N_20206);
xnor U22264 (N_22264,N_20913,N_20347);
nor U22265 (N_22265,N_20976,N_20096);
nor U22266 (N_22266,N_20672,N_20353);
and U22267 (N_22267,N_21860,N_21892);
and U22268 (N_22268,N_21490,N_21384);
nand U22269 (N_22269,N_20655,N_20544);
nand U22270 (N_22270,N_21471,N_21367);
nand U22271 (N_22271,N_20606,N_21937);
nor U22272 (N_22272,N_21941,N_21940);
nor U22273 (N_22273,N_21952,N_21558);
xor U22274 (N_22274,N_21209,N_21047);
or U22275 (N_22275,N_21590,N_20548);
nor U22276 (N_22276,N_20750,N_21511);
nand U22277 (N_22277,N_21245,N_20891);
nor U22278 (N_22278,N_21134,N_20701);
nor U22279 (N_22279,N_20911,N_21060);
xnor U22280 (N_22280,N_21875,N_20739);
and U22281 (N_22281,N_20823,N_21800);
or U22282 (N_22282,N_21213,N_21441);
nor U22283 (N_22283,N_20539,N_20219);
or U22284 (N_22284,N_20227,N_20540);
and U22285 (N_22285,N_21743,N_21972);
and U22286 (N_22286,N_20520,N_20600);
nor U22287 (N_22287,N_21747,N_20304);
nor U22288 (N_22288,N_21307,N_21928);
nor U22289 (N_22289,N_21758,N_21724);
and U22290 (N_22290,N_21448,N_20471);
and U22291 (N_22291,N_20977,N_20339);
and U22292 (N_22292,N_21456,N_21427);
xnor U22293 (N_22293,N_20129,N_20581);
xnor U22294 (N_22294,N_20584,N_21419);
and U22295 (N_22295,N_21533,N_20699);
xnor U22296 (N_22296,N_20961,N_21029);
xnor U22297 (N_22297,N_21640,N_21046);
or U22298 (N_22298,N_21818,N_20906);
and U22299 (N_22299,N_21715,N_21666);
xor U22300 (N_22300,N_21335,N_20771);
xor U22301 (N_22301,N_20774,N_20404);
or U22302 (N_22302,N_21599,N_21182);
nor U22303 (N_22303,N_20730,N_21418);
or U22304 (N_22304,N_21408,N_21841);
and U22305 (N_22305,N_21776,N_21660);
nand U22306 (N_22306,N_20814,N_21649);
or U22307 (N_22307,N_21254,N_20508);
xnor U22308 (N_22308,N_20255,N_21766);
nor U22309 (N_22309,N_21746,N_21210);
nand U22310 (N_22310,N_21604,N_20667);
nand U22311 (N_22311,N_21211,N_21066);
nor U22312 (N_22312,N_21914,N_21714);
xor U22313 (N_22313,N_21038,N_21275);
nand U22314 (N_22314,N_20557,N_20417);
and U22315 (N_22315,N_21015,N_20613);
nand U22316 (N_22316,N_20244,N_21825);
and U22317 (N_22317,N_20692,N_20806);
and U22318 (N_22318,N_21689,N_20236);
xnor U22319 (N_22319,N_20899,N_20439);
nor U22320 (N_22320,N_20827,N_20491);
xor U22321 (N_22321,N_21294,N_20653);
nor U22322 (N_22322,N_21998,N_20149);
xor U22323 (N_22323,N_21366,N_20431);
or U22324 (N_22324,N_20694,N_20182);
nand U22325 (N_22325,N_21201,N_21062);
xor U22326 (N_22326,N_21119,N_20014);
xor U22327 (N_22327,N_21540,N_21073);
nor U22328 (N_22328,N_21175,N_20555);
nand U22329 (N_22329,N_21483,N_20238);
or U22330 (N_22330,N_21135,N_20305);
and U22331 (N_22331,N_21195,N_20607);
nand U22332 (N_22332,N_20212,N_20561);
nor U22333 (N_22333,N_21527,N_20142);
and U22334 (N_22334,N_21446,N_20194);
nor U22335 (N_22335,N_21573,N_20139);
nand U22336 (N_22336,N_20467,N_20049);
nor U22337 (N_22337,N_21778,N_20766);
nand U22338 (N_22338,N_20796,N_20597);
nand U22339 (N_22339,N_21915,N_21820);
or U22340 (N_22340,N_20333,N_20440);
nor U22341 (N_22341,N_20720,N_20168);
nor U22342 (N_22342,N_20004,N_21801);
nand U22343 (N_22343,N_21181,N_20462);
nor U22344 (N_22344,N_20449,N_21224);
nor U22345 (N_22345,N_21082,N_21053);
and U22346 (N_22346,N_20170,N_21520);
nand U22347 (N_22347,N_21357,N_21609);
nand U22348 (N_22348,N_20041,N_21170);
and U22349 (N_22349,N_20565,N_21592);
xor U22350 (N_22350,N_21543,N_20514);
and U22351 (N_22351,N_20316,N_20161);
or U22352 (N_22352,N_20271,N_21432);
xor U22353 (N_22353,N_20868,N_20156);
or U22354 (N_22354,N_20810,N_20360);
nor U22355 (N_22355,N_20246,N_20438);
and U22356 (N_22356,N_20620,N_20703);
and U22357 (N_22357,N_20151,N_21754);
xor U22358 (N_22358,N_21827,N_20929);
or U22359 (N_22359,N_20335,N_20627);
and U22360 (N_22360,N_21094,N_21290);
or U22361 (N_22361,N_21547,N_20147);
xnor U22362 (N_22362,N_20193,N_21436);
nand U22363 (N_22363,N_21349,N_21232);
or U22364 (N_22364,N_21888,N_20656);
or U22365 (N_22365,N_21865,N_21516);
xnor U22366 (N_22366,N_20841,N_20336);
nor U22367 (N_22367,N_20780,N_21692);
nand U22368 (N_22368,N_21913,N_20838);
nand U22369 (N_22369,N_21378,N_21434);
or U22370 (N_22370,N_20114,N_21643);
nor U22371 (N_22371,N_20382,N_21740);
nor U22372 (N_22372,N_21961,N_21775);
nand U22373 (N_22373,N_20844,N_21171);
nand U22374 (N_22374,N_21979,N_21200);
and U22375 (N_22375,N_20998,N_21622);
nor U22376 (N_22376,N_21809,N_21453);
xnor U22377 (N_22377,N_20984,N_20295);
nor U22378 (N_22378,N_21266,N_20674);
and U22379 (N_22379,N_21899,N_21355);
nor U22380 (N_22380,N_20455,N_20272);
and U22381 (N_22381,N_21042,N_20850);
and U22382 (N_22382,N_21488,N_20300);
or U22383 (N_22383,N_21375,N_20110);
and U22384 (N_22384,N_20262,N_20052);
xor U22385 (N_22385,N_21194,N_20968);
and U22386 (N_22386,N_20095,N_20367);
xnor U22387 (N_22387,N_21943,N_20644);
nand U22388 (N_22388,N_21016,N_21454);
xor U22389 (N_22389,N_20534,N_21523);
and U22390 (N_22390,N_20450,N_21144);
and U22391 (N_22391,N_20947,N_20066);
nand U22392 (N_22392,N_21070,N_21553);
xnor U22393 (N_22393,N_21298,N_20634);
xor U22394 (N_22394,N_20558,N_21157);
nand U22395 (N_22395,N_21133,N_21240);
or U22396 (N_22396,N_20278,N_20187);
nor U22397 (N_22397,N_21978,N_20017);
xor U22398 (N_22398,N_20259,N_21946);
nor U22399 (N_22399,N_21538,N_20423);
and U22400 (N_22400,N_21414,N_20385);
and U22401 (N_22401,N_21634,N_21725);
nor U22402 (N_22402,N_20331,N_20490);
and U22403 (N_22403,N_21319,N_21798);
xor U22404 (N_22404,N_21145,N_21843);
xnor U22405 (N_22405,N_21882,N_21967);
and U22406 (N_22406,N_21314,N_20538);
and U22407 (N_22407,N_21944,N_20390);
and U22408 (N_22408,N_21010,N_20973);
and U22409 (N_22409,N_20031,N_20787);
xnor U22410 (N_22410,N_20019,N_20681);
and U22411 (N_22411,N_21938,N_20048);
or U22412 (N_22412,N_20320,N_20204);
or U22413 (N_22413,N_21154,N_21238);
nand U22414 (N_22414,N_21466,N_20260);
xnor U22415 (N_22415,N_20258,N_20411);
xnor U22416 (N_22416,N_21777,N_20784);
nand U22417 (N_22417,N_21068,N_20443);
nand U22418 (N_22418,N_20542,N_21489);
nor U22419 (N_22419,N_20834,N_21410);
or U22420 (N_22420,N_20294,N_20884);
and U22421 (N_22421,N_21957,N_21813);
and U22422 (N_22422,N_21421,N_21243);
and U22423 (N_22423,N_20971,N_21734);
nand U22424 (N_22424,N_21605,N_21092);
or U22425 (N_22425,N_21337,N_21748);
nor U22426 (N_22426,N_21954,N_20001);
xor U22427 (N_22427,N_21126,N_20988);
nor U22428 (N_22428,N_20646,N_20016);
nand U22429 (N_22429,N_21608,N_21476);
nor U22430 (N_22430,N_20945,N_21343);
nand U22431 (N_22431,N_21284,N_20885);
or U22432 (N_22432,N_20174,N_20618);
xor U22433 (N_22433,N_21557,N_20734);
nand U22434 (N_22434,N_20297,N_20531);
nor U22435 (N_22435,N_20344,N_20698);
xor U22436 (N_22436,N_20086,N_20228);
or U22437 (N_22437,N_21452,N_20659);
and U22438 (N_22438,N_20994,N_21768);
or U22439 (N_22439,N_20464,N_20397);
xnor U22440 (N_22440,N_21830,N_20917);
nand U22441 (N_22441,N_20586,N_20535);
or U22442 (N_22442,N_21143,N_21982);
xor U22443 (N_22443,N_20222,N_21617);
or U22444 (N_22444,N_21226,N_20116);
xor U22445 (N_22445,N_20167,N_20218);
or U22446 (N_22446,N_21728,N_21544);
xnor U22447 (N_22447,N_20074,N_21773);
or U22448 (N_22448,N_21564,N_20137);
and U22449 (N_22449,N_20356,N_20273);
nand U22450 (N_22450,N_21930,N_21772);
nor U22451 (N_22451,N_20611,N_20124);
nand U22452 (N_22452,N_21045,N_21328);
xnor U22453 (N_22453,N_21989,N_21189);
nand U22454 (N_22454,N_21757,N_20716);
and U22455 (N_22455,N_20418,N_20536);
or U22456 (N_22456,N_21854,N_20859);
xnor U22457 (N_22457,N_20855,N_21348);
and U22458 (N_22458,N_21549,N_20671);
nor U22459 (N_22459,N_21313,N_21579);
and U22460 (N_22460,N_20788,N_20327);
nor U22461 (N_22461,N_20106,N_21102);
or U22462 (N_22462,N_20754,N_21596);
nor U22463 (N_22463,N_21641,N_20836);
nand U22464 (N_22464,N_20954,N_21876);
nand U22465 (N_22465,N_21044,N_20101);
or U22466 (N_22466,N_20188,N_21976);
and U22467 (N_22467,N_21765,N_20657);
or U22468 (N_22468,N_21438,N_21009);
xnor U22469 (N_22469,N_21680,N_21681);
or U22470 (N_22470,N_21536,N_20745);
nor U22471 (N_22471,N_21795,N_20115);
nand U22472 (N_22472,N_20309,N_20969);
and U22473 (N_22473,N_21869,N_21196);
nand U22474 (N_22474,N_21086,N_20992);
or U22475 (N_22475,N_20791,N_21006);
nor U22476 (N_22476,N_21668,N_21518);
xnor U22477 (N_22477,N_20386,N_20059);
and U22478 (N_22478,N_21004,N_20365);
or U22479 (N_22479,N_20224,N_20760);
and U22480 (N_22480,N_21614,N_21122);
nor U22481 (N_22481,N_20424,N_20340);
nand U22482 (N_22482,N_20883,N_21514);
nand U22483 (N_22483,N_20881,N_20283);
nand U22484 (N_22484,N_21400,N_20522);
or U22485 (N_22485,N_20057,N_21252);
xnor U22486 (N_22486,N_21853,N_20588);
nand U22487 (N_22487,N_20136,N_20459);
or U22488 (N_22488,N_21712,N_20727);
and U22489 (N_22489,N_20590,N_21994);
nor U22490 (N_22490,N_20735,N_20504);
nor U22491 (N_22491,N_21909,N_20728);
or U22492 (N_22492,N_21606,N_21428);
or U22493 (N_22493,N_21953,N_21310);
or U22494 (N_22494,N_20993,N_21291);
and U22495 (N_22495,N_20936,N_21507);
and U22496 (N_22496,N_21545,N_20184);
nor U22497 (N_22497,N_20748,N_20299);
xnor U22498 (N_22498,N_21088,N_20267);
and U22499 (N_22499,N_20179,N_20183);
or U22500 (N_22500,N_20349,N_21688);
or U22501 (N_22501,N_20526,N_21286);
nor U22502 (N_22502,N_20831,N_21439);
and U22503 (N_22503,N_21385,N_21517);
and U22504 (N_22504,N_21559,N_20025);
or U22505 (N_22505,N_21264,N_21296);
or U22506 (N_22506,N_21705,N_21745);
nand U22507 (N_22507,N_21311,N_20088);
xor U22508 (N_22508,N_21390,N_21239);
nor U22509 (N_22509,N_20662,N_21509);
and U22510 (N_22510,N_21282,N_21214);
nand U22511 (N_22511,N_20409,N_21180);
nor U22512 (N_22512,N_20369,N_21625);
or U22513 (N_22513,N_20165,N_20890);
or U22514 (N_22514,N_20169,N_20619);
and U22515 (N_22515,N_21977,N_20126);
or U22516 (N_22516,N_20458,N_21155);
or U22517 (N_22517,N_21352,N_20970);
or U22518 (N_22518,N_20375,N_21999);
and U22519 (N_22519,N_21219,N_20091);
xnor U22520 (N_22520,N_20325,N_20400);
nand U22521 (N_22521,N_21292,N_21603);
xor U22522 (N_22522,N_20525,N_20190);
nor U22523 (N_22523,N_21880,N_21719);
xnor U22524 (N_22524,N_20090,N_21834);
xor U22525 (N_22525,N_21040,N_21817);
xnor U22526 (N_22526,N_21300,N_20654);
or U22527 (N_22527,N_21074,N_21988);
or U22528 (N_22528,N_20078,N_20893);
or U22529 (N_22529,N_21720,N_20392);
xor U22530 (N_22530,N_20507,N_21477);
and U22531 (N_22531,N_20301,N_21247);
or U22532 (N_22532,N_20903,N_20092);
or U22533 (N_22533,N_20553,N_21262);
xor U22534 (N_22534,N_20663,N_21949);
or U22535 (N_22535,N_20311,N_21049);
nand U22536 (N_22536,N_21984,N_20261);
or U22537 (N_22537,N_20447,N_20122);
and U22538 (N_22538,N_20550,N_20677);
xor U22539 (N_22539,N_20248,N_21515);
or U22540 (N_22540,N_20034,N_20501);
and U22541 (N_22541,N_21797,N_21147);
or U22542 (N_22542,N_20552,N_20348);
xor U22543 (N_22543,N_21429,N_20647);
nor U22544 (N_22544,N_20055,N_21661);
nor U22545 (N_22545,N_21459,N_20217);
xnor U22546 (N_22546,N_21198,N_20509);
nor U22547 (N_22547,N_21031,N_21848);
or U22548 (N_22548,N_20649,N_20481);
and U22549 (N_22549,N_20869,N_20279);
nor U22550 (N_22550,N_21968,N_20582);
and U22551 (N_22551,N_20761,N_21936);
or U22552 (N_22552,N_21508,N_21234);
xnor U22553 (N_22553,N_21682,N_21645);
and U22554 (N_22554,N_21629,N_21499);
xnor U22555 (N_22555,N_21076,N_21723);
nand U22556 (N_22556,N_20942,N_21140);
or U22557 (N_22557,N_21686,N_21469);
and U22558 (N_22558,N_21071,N_21850);
nand U22559 (N_22559,N_20130,N_20943);
xnor U22560 (N_22560,N_21184,N_20022);
or U22561 (N_22561,N_21033,N_20275);
or U22562 (N_22562,N_21387,N_21026);
xnor U22563 (N_22563,N_20250,N_20898);
or U22564 (N_22564,N_21162,N_21447);
or U22565 (N_22565,N_21753,N_21164);
nand U22566 (N_22566,N_20160,N_20910);
nand U22567 (N_22567,N_21302,N_21644);
nand U22568 (N_22568,N_21920,N_21997);
nor U22569 (N_22569,N_20071,N_21411);
nor U22570 (N_22570,N_21665,N_20100);
nor U22571 (N_22571,N_20478,N_20695);
or U22572 (N_22572,N_20660,N_20704);
or U22573 (N_22573,N_21110,N_20428);
nand U22574 (N_22574,N_21610,N_21960);
nand U22575 (N_22575,N_20516,N_21445);
xnor U22576 (N_22576,N_20762,N_20955);
or U22577 (N_22577,N_20480,N_20658);
xnor U22578 (N_22578,N_21752,N_21806);
nor U22579 (N_22579,N_21287,N_20722);
nand U22580 (N_22580,N_21316,N_21061);
or U22581 (N_22581,N_20426,N_21087);
nand U22582 (N_22582,N_20562,N_20811);
xnor U22583 (N_22583,N_20837,N_20758);
and U22584 (N_22584,N_21951,N_20415);
and U22585 (N_22585,N_20668,N_20243);
or U22586 (N_22586,N_20181,N_21707);
or U22587 (N_22587,N_21364,N_21846);
nand U22588 (N_22588,N_21556,N_21512);
nor U22589 (N_22589,N_21896,N_20650);
nor U22590 (N_22590,N_20532,N_20323);
xnor U22591 (N_22591,N_21812,N_20909);
nand U22592 (N_22592,N_21199,N_20198);
and U22593 (N_22593,N_20494,N_20633);
and U22594 (N_22594,N_21106,N_21217);
and U22595 (N_22595,N_20402,N_21601);
or U22596 (N_22596,N_20384,N_21350);
nand U22597 (N_22597,N_21117,N_20268);
or U22598 (N_22598,N_20277,N_21833);
xor U22599 (N_22599,N_20839,N_21700);
or U22600 (N_22600,N_21903,N_21244);
xor U22601 (N_22601,N_21485,N_21623);
and U22602 (N_22602,N_20203,N_20604);
or U22603 (N_22603,N_21295,N_21885);
or U22604 (N_22604,N_20682,N_21193);
xor U22605 (N_22605,N_20191,N_21465);
xor U22606 (N_22606,N_20082,N_21494);
nor U22607 (N_22607,N_21467,N_20905);
xnor U22608 (N_22608,N_21906,N_20856);
and U22609 (N_22609,N_20900,N_20713);
nor U22610 (N_22610,N_21192,N_20302);
or U22611 (N_22611,N_21939,N_21526);
xor U22612 (N_22612,N_20789,N_21108);
nand U22613 (N_22613,N_21072,N_21424);
and U22614 (N_22614,N_20953,N_21116);
or U22615 (N_22615,N_21277,N_20162);
nand U22616 (N_22616,N_20109,N_20710);
nand U22617 (N_22617,N_21701,N_21034);
or U22618 (N_22618,N_21115,N_21473);
or U22619 (N_22619,N_20957,N_20241);
xor U22620 (N_22620,N_21197,N_21078);
xor U22621 (N_22621,N_20732,N_20628);
xnor U22622 (N_22622,N_20875,N_21165);
and U22623 (N_22623,N_20050,N_20979);
nand U22624 (N_22624,N_20797,N_20453);
xor U22625 (N_22625,N_20225,N_21190);
nor U22626 (N_22626,N_21440,N_21373);
and U22627 (N_22627,N_20216,N_21173);
or U22628 (N_22628,N_21910,N_20445);
and U22629 (N_22629,N_20676,N_21323);
xor U22630 (N_22630,N_21139,N_21856);
xor U22631 (N_22631,N_21163,N_20962);
or U22632 (N_22632,N_21272,N_20685);
or U22633 (N_22633,N_20042,N_20021);
or U22634 (N_22634,N_20274,N_20247);
nor U22635 (N_22635,N_21799,N_20770);
xnor U22636 (N_22636,N_20785,N_21836);
and U22637 (N_22637,N_20121,N_21529);
xor U22638 (N_22638,N_20632,N_21739);
and U22639 (N_22639,N_20079,N_20925);
nor U22640 (N_22640,N_20383,N_20921);
nor U22641 (N_22641,N_21095,N_20457);
nor U22642 (N_22642,N_20551,N_20888);
nor U22643 (N_22643,N_20500,N_20688);
nor U22644 (N_22644,N_21069,N_21065);
or U22645 (N_22645,N_21112,N_20571);
and U22646 (N_22646,N_20479,N_20960);
nor U22647 (N_22647,N_21621,N_21204);
nand U22648 (N_22648,N_20153,N_21808);
nor U22649 (N_22649,N_20492,N_20782);
and U22650 (N_22650,N_21435,N_21513);
or U22651 (N_22651,N_20513,N_20028);
or U22652 (N_22652,N_21111,N_20880);
and U22653 (N_22653,N_20963,N_21627);
nor U22654 (N_22654,N_21562,N_20959);
xor U22655 (N_22655,N_20744,N_20986);
xor U22656 (N_22656,N_20010,N_20437);
or U22657 (N_22657,N_21237,N_21492);
xor U22658 (N_22658,N_21406,N_20374);
nor U22659 (N_22659,N_21278,N_20239);
and U22660 (N_22660,N_21828,N_20997);
and U22661 (N_22661,N_20280,N_20731);
xor U22662 (N_22662,N_20543,N_21382);
xnor U22663 (N_22663,N_21787,N_20351);
or U22664 (N_22664,N_20446,N_21654);
xnor U22665 (N_22665,N_20207,N_21585);
and U22666 (N_22666,N_20854,N_20290);
nand U22667 (N_22667,N_20039,N_21460);
nor U22668 (N_22668,N_21091,N_20527);
or U22669 (N_22669,N_20366,N_21359);
nor U22670 (N_22670,N_20105,N_20412);
xnor U22671 (N_22671,N_20512,N_20282);
xnor U22672 (N_22672,N_21638,N_20908);
nand U22673 (N_22673,N_20433,N_20343);
and U22674 (N_22674,N_21423,N_20242);
and U22675 (N_22675,N_21396,N_20877);
xnor U22676 (N_22676,N_20251,N_21677);
or U22677 (N_22677,N_21371,N_20560);
nand U22678 (N_22678,N_20405,N_20846);
xor U22679 (N_22679,N_20940,N_20775);
nor U22680 (N_22680,N_21221,N_20779);
nand U22681 (N_22681,N_20629,N_20948);
and U22682 (N_22682,N_20615,N_21602);
nand U22683 (N_22683,N_21131,N_21345);
nand U22684 (N_22684,N_20002,N_20286);
or U22685 (N_22685,N_21413,N_20651);
or U22686 (N_22686,N_20705,N_20980);
nand U22687 (N_22687,N_20070,N_21669);
xor U22688 (N_22688,N_20497,N_20403);
and U22689 (N_22689,N_21120,N_20608);
nor U22690 (N_22690,N_20801,N_20822);
nor U22691 (N_22691,N_20421,N_21852);
nor U22692 (N_22692,N_20035,N_20003);
nand U22693 (N_22693,N_21075,N_20511);
nor U22694 (N_22694,N_21908,N_20897);
or U22695 (N_22695,N_20060,N_20591);
nor U22696 (N_22696,N_21039,N_20570);
or U22697 (N_22697,N_20451,N_20045);
and U22698 (N_22698,N_21580,N_20637);
nand U22699 (N_22699,N_21032,N_21620);
nor U22700 (N_22700,N_20061,N_21589);
xor U22701 (N_22701,N_21386,N_20937);
and U22702 (N_22702,N_20825,N_21550);
or U22703 (N_22703,N_20173,N_21862);
nor U22704 (N_22704,N_20851,N_21481);
or U22705 (N_22705,N_21927,N_21208);
and U22706 (N_22706,N_20202,N_20537);
nand U22707 (N_22707,N_20853,N_20569);
nor U22708 (N_22708,N_20664,N_21932);
or U22709 (N_22709,N_21859,N_21807);
xor U22710 (N_22710,N_20724,N_21803);
nand U22711 (N_22711,N_21992,N_21370);
nor U22712 (N_22712,N_20140,N_20387);
nand U22713 (N_22713,N_20220,N_21475);
xor U22714 (N_22714,N_20696,N_20186);
xor U22715 (N_22715,N_20373,N_20083);
nand U22716 (N_22716,N_21374,N_21451);
and U22717 (N_22717,N_20598,N_21104);
nand U22718 (N_22718,N_20861,N_20352);
or U22719 (N_22719,N_20858,N_20956);
and U22720 (N_22720,N_21996,N_20648);
or U22721 (N_22721,N_20602,N_20924);
and U22722 (N_22722,N_20585,N_20510);
and U22723 (N_22723,N_21354,N_20737);
and U22724 (N_22724,N_20102,N_20573);
nor U22725 (N_22725,N_21789,N_20062);
or U22726 (N_22726,N_21866,N_20564);
and U22727 (N_22727,N_21890,N_21676);
nand U22728 (N_22728,N_20429,N_20719);
or U22729 (N_22729,N_20641,N_21679);
nor U22730 (N_22730,N_20575,N_21231);
nor U22731 (N_22731,N_21251,N_21729);
nor U22732 (N_22732,N_21970,N_20915);
nor U22733 (N_22733,N_21089,N_20310);
nand U22734 (N_22734,N_20489,N_20388);
and U22735 (N_22735,N_21898,N_21615);
or U22736 (N_22736,N_21242,N_20505);
or U22737 (N_22737,N_21020,N_20865);
and U22738 (N_22738,N_20958,N_21774);
xnor U22739 (N_22739,N_21085,N_21636);
nand U22740 (N_22740,N_21571,N_21149);
and U22741 (N_22741,N_21991,N_21551);
nand U22742 (N_22742,N_20684,N_21055);
and U22743 (N_22743,N_21934,N_20616);
nor U22744 (N_22744,N_21114,N_20642);
nor U22745 (N_22745,N_21394,N_21083);
xor U22746 (N_22746,N_20329,N_20803);
xnor U22747 (N_22747,N_21096,N_21923);
nor U22748 (N_22748,N_20625,N_20342);
nand U22749 (N_22749,N_21814,N_20293);
or U22750 (N_22750,N_21329,N_21057);
and U22751 (N_22751,N_21962,N_21790);
or U22752 (N_22752,N_20346,N_21935);
and U22753 (N_22753,N_20328,N_21738);
nor U22754 (N_22754,N_21653,N_21305);
nand U22755 (N_22755,N_20094,N_20355);
xnor U22756 (N_22756,N_20370,N_20185);
or U22757 (N_22757,N_21534,N_21215);
nor U22758 (N_22758,N_21222,N_21283);
and U22759 (N_22759,N_21129,N_21598);
nor U22760 (N_22760,N_21261,N_20406);
nor U22761 (N_22761,N_20506,N_20794);
nor U22762 (N_22762,N_21762,N_20776);
nor U22763 (N_22763,N_21779,N_20759);
or U22764 (N_22764,N_21816,N_21933);
xor U22765 (N_22765,N_20715,N_21166);
nor U22766 (N_22766,N_20377,N_21755);
or U22767 (N_22767,N_20617,N_20132);
nand U22768 (N_22768,N_21541,N_21586);
or U22769 (N_22769,N_21321,N_21675);
and U22770 (N_22770,N_20576,N_21461);
xnor U22771 (N_22771,N_20743,N_21336);
nand U22772 (N_22772,N_20673,N_20399);
and U22773 (N_22773,N_21717,N_21631);
xnor U22774 (N_22774,N_20817,N_20345);
xnor U22775 (N_22775,N_20298,N_20583);
nor U22776 (N_22776,N_20288,N_20436);
nand U22777 (N_22777,N_21959,N_20874);
nand U22778 (N_22778,N_20020,N_20125);
xor U22779 (N_22779,N_20843,N_21713);
or U22780 (N_22780,N_21901,N_20150);
and U22781 (N_22781,N_20640,N_20474);
xnor U22782 (N_22782,N_20254,N_21276);
xnor U22783 (N_22783,N_20867,N_21253);
nor U22784 (N_22784,N_20211,N_21522);
nor U22785 (N_22785,N_21736,N_21981);
xnor U22786 (N_22786,N_21821,N_21158);
and U22787 (N_22787,N_21330,N_21480);
nand U22788 (N_22788,N_20741,N_20612);
xor U22789 (N_22789,N_21167,N_21711);
nor U22790 (N_22790,N_21811,N_20545);
and U22791 (N_22791,N_21703,N_21922);
xor U22792 (N_22792,N_20223,N_20163);
nor U22793 (N_22793,N_20595,N_21363);
nor U22794 (N_22794,N_20456,N_21673);
nand U22795 (N_22795,N_21401,N_20037);
nand U22796 (N_22796,N_21709,N_21530);
or U22797 (N_22797,N_20209,N_21392);
or U22798 (N_22798,N_21504,N_21127);
or U22799 (N_22799,N_21142,N_21955);
nand U22800 (N_22800,N_20155,N_21493);
and U22801 (N_22801,N_20587,N_20119);
xnor U22802 (N_22802,N_20482,N_21051);
xor U22803 (N_22803,N_21662,N_20486);
nand U22804 (N_22804,N_21404,N_20493);
xnor U22805 (N_22805,N_21886,N_20159);
xor U22806 (N_22806,N_20064,N_21369);
xnor U22807 (N_22807,N_20172,N_21121);
and U22808 (N_22808,N_20138,N_20166);
nor U22809 (N_22809,N_20477,N_20965);
and U22810 (N_22810,N_20178,N_21593);
nor U22811 (N_22811,N_20808,N_21626);
nand U22812 (N_22812,N_21907,N_20757);
nor U22813 (N_22813,N_20133,N_20334);
nor U22814 (N_22814,N_20572,N_21658);
xnor U22815 (N_22815,N_20714,N_21726);
nand U22816 (N_22816,N_20927,N_21274);
nand U22817 (N_22817,N_20269,N_21079);
nor U22818 (N_22818,N_20763,N_21698);
or U22819 (N_22819,N_21652,N_20396);
nand U22820 (N_22820,N_20499,N_20487);
nand U22821 (N_22821,N_20077,N_21344);
or U22822 (N_22822,N_20407,N_20357);
and U22823 (N_22823,N_20678,N_21582);
nor U22824 (N_22824,N_20580,N_21670);
nor U22825 (N_22825,N_20379,N_20914);
and U22826 (N_22826,N_21710,N_20669);
or U22827 (N_22827,N_20069,N_20675);
nor U22828 (N_22828,N_21613,N_21365);
or U22829 (N_22829,N_20983,N_20056);
or U22830 (N_22830,N_21397,N_20845);
and U22831 (N_22831,N_20068,N_20700);
nand U22832 (N_22832,N_20291,N_21437);
and U22833 (N_22833,N_20920,N_21388);
xnor U22834 (N_22834,N_21784,N_20805);
nor U22835 (N_22835,N_21985,N_21851);
or U22836 (N_22836,N_21872,N_21023);
or U22837 (N_22837,N_21309,N_20939);
nand U22838 (N_22838,N_21052,N_20465);
xnor U22839 (N_22839,N_21464,N_20860);
and U22840 (N_22840,N_20319,N_20603);
and U22841 (N_22841,N_20578,N_21012);
xnor U22842 (N_22842,N_21398,N_20712);
xor U22843 (N_22843,N_20974,N_20498);
and U22844 (N_22844,N_20769,N_21080);
and U22845 (N_22845,N_20024,N_21980);
nand U22846 (N_22846,N_21325,N_21655);
nand U22847 (N_22847,N_20127,N_21322);
nand U22848 (N_22848,N_21502,N_20533);
or U22849 (N_22849,N_20321,N_21731);
xnor U22850 (N_22850,N_21169,N_21942);
and U22851 (N_22851,N_21506,N_21548);
nand U22852 (N_22852,N_21005,N_21897);
nor U22853 (N_22853,N_21403,N_21356);
or U22854 (N_22854,N_20946,N_20829);
nand U22855 (N_22855,N_20802,N_21183);
or U22856 (N_22856,N_21581,N_20111);
nor U22857 (N_22857,N_20073,N_20085);
nor U22858 (N_22858,N_21539,N_20229);
and U22859 (N_22859,N_21402,N_20907);
nor U22860 (N_22860,N_20215,N_21101);
and U22861 (N_22861,N_21021,N_20249);
nand U22862 (N_22862,N_21235,N_21315);
and U22863 (N_22863,N_21919,N_20559);
and U22864 (N_22864,N_20234,N_20018);
xor U22865 (N_22865,N_20528,N_21684);
and U22866 (N_22866,N_21824,N_21425);
nor U22867 (N_22867,N_20686,N_20645);
or U22868 (N_22868,N_20746,N_21308);
xor U22869 (N_22869,N_20435,N_21566);
nor U22870 (N_22870,N_20725,N_21630);
or U22871 (N_22871,N_20687,N_20864);
or U22872 (N_22872,N_20463,N_21505);
and U22873 (N_22873,N_21035,N_20488);
nor U22874 (N_22874,N_21037,N_20848);
xnor U22875 (N_22875,N_20521,N_21618);
and U22876 (N_22876,N_20833,N_21368);
and U22877 (N_22877,N_21203,N_20636);
nor U22878 (N_22878,N_20108,N_21098);
xnor U22879 (N_22879,N_20470,N_20756);
xnor U22880 (N_22880,N_20871,N_21672);
nand U22881 (N_22881,N_21153,N_20697);
nor U22882 (N_22882,N_20589,N_20120);
and U22883 (N_22883,N_21002,N_20231);
or U22884 (N_22884,N_21303,N_20205);
nand U22885 (N_22885,N_21236,N_20131);
or U22886 (N_22886,N_21727,N_20702);
and U22887 (N_22887,N_21484,N_21028);
and U22888 (N_22888,N_21289,N_21761);
or U22889 (N_22889,N_20143,N_21218);
nand U22890 (N_22890,N_20923,N_21077);
and U22891 (N_22891,N_21389,N_20416);
and U22892 (N_22892,N_20815,N_21815);
or U22893 (N_22893,N_20596,N_21756);
nand U22894 (N_22894,N_20338,N_21624);
and U22895 (N_22895,N_20949,N_21956);
nor U22896 (N_22896,N_21525,N_20427);
nor U22897 (N_22897,N_21161,N_21785);
and U22898 (N_22898,N_21017,N_20176);
or U22899 (N_22899,N_21433,N_21174);
nor U22900 (N_22900,N_21187,N_21084);
and U22901 (N_22901,N_21177,N_20800);
nor U22902 (N_22902,N_21132,N_21683);
xor U22903 (N_22903,N_20098,N_20337);
or U22904 (N_22904,N_21351,N_20000);
and U22905 (N_22905,N_20097,N_21118);
nor U22906 (N_22906,N_21706,N_20452);
and U22907 (N_22907,N_21297,N_21750);
or U22908 (N_22908,N_21416,N_20009);
and U22909 (N_22909,N_21479,N_20263);
nor U22910 (N_22910,N_20807,N_20764);
nor U22911 (N_22911,N_21510,N_21470);
or U22912 (N_22912,N_20087,N_20063);
or U22913 (N_22913,N_21926,N_20307);
nor U22914 (N_22914,N_21737,N_21849);
nor U22915 (N_22915,N_21463,N_21567);
nor U22916 (N_22916,N_20419,N_21496);
nor U22917 (N_22917,N_21097,N_21792);
nand U22918 (N_22918,N_21565,N_21265);
nor U22919 (N_22919,N_20777,N_21781);
nor U22920 (N_22920,N_20080,N_20253);
xor U22921 (N_22921,N_21273,N_20030);
nor U22922 (N_22922,N_21450,N_21136);
and U22923 (N_22923,N_21360,N_20999);
and U22924 (N_22924,N_21845,N_20765);
xor U22925 (N_22925,N_21380,N_21468);
nand U22926 (N_22926,N_21528,N_21025);
nand U22927 (N_22927,N_21879,N_21409);
or U22928 (N_22928,N_20292,N_21260);
or U22929 (N_22929,N_20430,N_20982);
nand U22930 (N_22930,N_20889,N_21361);
xor U22931 (N_22931,N_21771,N_20579);
xnor U22932 (N_22932,N_20813,N_21263);
nand U22933 (N_22933,N_21148,N_20380);
xor U22934 (N_22934,N_21782,N_20007);
and U22935 (N_22935,N_21749,N_21255);
nor U22936 (N_22936,N_21246,N_20840);
and U22937 (N_22937,N_21628,N_21986);
and U22938 (N_22938,N_21607,N_20306);
xor U22939 (N_22939,N_20332,N_21891);
and U22940 (N_22940,N_21318,N_20053);
or U22941 (N_22941,N_20413,N_20134);
nor U22942 (N_22942,N_21326,N_20107);
and U22943 (N_22943,N_21524,N_20738);
or U22944 (N_22944,N_20816,N_21838);
and U22945 (N_22945,N_21973,N_20631);
nand U22946 (N_22946,N_21868,N_20197);
nand U22947 (N_22947,N_21443,N_21205);
and U22948 (N_22948,N_21542,N_20441);
xor U22949 (N_22949,N_21267,N_20444);
nor U22950 (N_22950,N_21188,N_20952);
nand U22951 (N_22951,N_21176,N_21259);
nor U22952 (N_22952,N_20934,N_20213);
and U22953 (N_22953,N_20966,N_21697);
nand U22954 (N_22954,N_20886,N_21597);
xor U22955 (N_22955,N_20876,N_21983);
and U22956 (N_22956,N_21312,N_20484);
xnor U22957 (N_22957,N_21921,N_20044);
nand U22958 (N_22958,N_20930,N_20099);
xnor U22959 (N_22959,N_20951,N_20751);
nor U22960 (N_22960,N_20733,N_21248);
or U22961 (N_22961,N_21895,N_20200);
nor U22962 (N_22962,N_20317,N_20112);
nor U22963 (N_22963,N_21391,N_20285);
xnor U22964 (N_22964,N_21829,N_21584);
nand U22965 (N_22965,N_21334,N_20792);
nor U22966 (N_22966,N_20326,N_21671);
and U22967 (N_22967,N_20709,N_20643);
and U22968 (N_22968,N_21054,N_20879);
and U22969 (N_22969,N_20011,N_20395);
nand U22970 (N_22970,N_21241,N_21863);
nor U22971 (N_22971,N_21646,N_20117);
and U22972 (N_22972,N_21873,N_20157);
or U22973 (N_22973,N_20849,N_20981);
xnor U22974 (N_22974,N_20284,N_21206);
nor U22975 (N_22975,N_21172,N_20180);
nand U22976 (N_22976,N_20154,N_20103);
and U22977 (N_22977,N_21881,N_21639);
xnor U22978 (N_22978,N_20901,N_20089);
xnor U22979 (N_22979,N_21063,N_21878);
nor U22980 (N_22980,N_20058,N_20972);
nand U22981 (N_22981,N_21722,N_21285);
nand U22982 (N_22982,N_21742,N_21064);
nor U22983 (N_22983,N_20313,N_20350);
and U22984 (N_22984,N_20990,N_21299);
nand U22985 (N_22985,N_20287,N_20870);
nor U22986 (N_22986,N_21151,N_21141);
nand U22987 (N_22987,N_21577,N_21306);
xor U22988 (N_22988,N_20931,N_20425);
or U22989 (N_22989,N_21159,N_21902);
and U22990 (N_22990,N_21842,N_21874);
and U22991 (N_22991,N_20793,N_20257);
or U22992 (N_22992,N_21426,N_21270);
nor U22993 (N_22993,N_20442,N_21430);
nand U22994 (N_22994,N_21249,N_21501);
nor U22995 (N_22995,N_20729,N_20118);
nand U22996 (N_22996,N_20592,N_20221);
nor U22997 (N_22997,N_21563,N_21482);
nand U22998 (N_22998,N_20201,N_20398);
nand U22999 (N_22999,N_20798,N_21268);
nand U23000 (N_23000,N_21051,N_20514);
xnor U23001 (N_23001,N_21508,N_21780);
nor U23002 (N_23002,N_20078,N_21473);
nand U23003 (N_23003,N_21830,N_20700);
nand U23004 (N_23004,N_21890,N_21356);
and U23005 (N_23005,N_20063,N_20234);
nor U23006 (N_23006,N_21818,N_20974);
and U23007 (N_23007,N_21342,N_20043);
nand U23008 (N_23008,N_20614,N_21075);
nand U23009 (N_23009,N_21949,N_20296);
nand U23010 (N_23010,N_20543,N_20440);
xnor U23011 (N_23011,N_21379,N_20071);
xnor U23012 (N_23012,N_21052,N_20149);
nor U23013 (N_23013,N_20856,N_20943);
nor U23014 (N_23014,N_20597,N_21146);
xor U23015 (N_23015,N_20576,N_21161);
and U23016 (N_23016,N_21164,N_20244);
nor U23017 (N_23017,N_20172,N_20817);
or U23018 (N_23018,N_20170,N_20475);
xnor U23019 (N_23019,N_20556,N_20841);
nor U23020 (N_23020,N_21762,N_21809);
nor U23021 (N_23021,N_20922,N_20129);
and U23022 (N_23022,N_20051,N_21077);
nand U23023 (N_23023,N_20719,N_21519);
nor U23024 (N_23024,N_20186,N_20514);
and U23025 (N_23025,N_21302,N_20296);
and U23026 (N_23026,N_21723,N_21471);
or U23027 (N_23027,N_21944,N_21105);
nand U23028 (N_23028,N_21337,N_20537);
and U23029 (N_23029,N_20123,N_21074);
or U23030 (N_23030,N_21770,N_20845);
nand U23031 (N_23031,N_21368,N_20045);
xnor U23032 (N_23032,N_20496,N_21894);
or U23033 (N_23033,N_21546,N_21028);
nand U23034 (N_23034,N_20593,N_21477);
nor U23035 (N_23035,N_20199,N_21814);
or U23036 (N_23036,N_21077,N_21128);
or U23037 (N_23037,N_21995,N_21731);
nand U23038 (N_23038,N_21449,N_21608);
xnor U23039 (N_23039,N_21286,N_21501);
and U23040 (N_23040,N_20866,N_21738);
nand U23041 (N_23041,N_20177,N_20339);
xor U23042 (N_23042,N_21459,N_20358);
and U23043 (N_23043,N_21142,N_21929);
and U23044 (N_23044,N_21561,N_20110);
nand U23045 (N_23045,N_20930,N_20220);
or U23046 (N_23046,N_21443,N_20719);
or U23047 (N_23047,N_21424,N_21874);
xor U23048 (N_23048,N_20640,N_20692);
and U23049 (N_23049,N_20005,N_20281);
xor U23050 (N_23050,N_20232,N_21115);
nor U23051 (N_23051,N_21146,N_20383);
xor U23052 (N_23052,N_20525,N_20498);
nand U23053 (N_23053,N_20425,N_20249);
nand U23054 (N_23054,N_20393,N_20795);
and U23055 (N_23055,N_21369,N_20663);
xnor U23056 (N_23056,N_20952,N_20579);
or U23057 (N_23057,N_21567,N_21489);
or U23058 (N_23058,N_20153,N_20982);
nor U23059 (N_23059,N_20269,N_21296);
and U23060 (N_23060,N_20333,N_21961);
and U23061 (N_23061,N_21479,N_20949);
nand U23062 (N_23062,N_21763,N_20029);
nor U23063 (N_23063,N_20399,N_20634);
xor U23064 (N_23064,N_20505,N_20608);
xor U23065 (N_23065,N_21420,N_21660);
or U23066 (N_23066,N_21204,N_21759);
nor U23067 (N_23067,N_21303,N_20171);
xnor U23068 (N_23068,N_20133,N_20247);
nor U23069 (N_23069,N_21216,N_20860);
xor U23070 (N_23070,N_21525,N_21129);
nor U23071 (N_23071,N_21302,N_21513);
and U23072 (N_23072,N_21487,N_20008);
and U23073 (N_23073,N_21990,N_21734);
nand U23074 (N_23074,N_20310,N_21289);
nor U23075 (N_23075,N_20075,N_21875);
and U23076 (N_23076,N_20290,N_21824);
nor U23077 (N_23077,N_20811,N_20337);
or U23078 (N_23078,N_21692,N_20326);
nand U23079 (N_23079,N_21493,N_21389);
and U23080 (N_23080,N_20732,N_21865);
xor U23081 (N_23081,N_21023,N_20097);
and U23082 (N_23082,N_21360,N_20961);
and U23083 (N_23083,N_21307,N_20189);
nand U23084 (N_23084,N_20317,N_20532);
or U23085 (N_23085,N_20517,N_21522);
nor U23086 (N_23086,N_21168,N_20686);
or U23087 (N_23087,N_20222,N_21370);
nand U23088 (N_23088,N_21250,N_20296);
xor U23089 (N_23089,N_20553,N_21880);
or U23090 (N_23090,N_20628,N_20437);
and U23091 (N_23091,N_21991,N_20235);
and U23092 (N_23092,N_20378,N_21848);
nor U23093 (N_23093,N_21294,N_21204);
nand U23094 (N_23094,N_20903,N_21113);
or U23095 (N_23095,N_21059,N_21230);
nor U23096 (N_23096,N_21659,N_21309);
nor U23097 (N_23097,N_21034,N_20872);
nand U23098 (N_23098,N_20214,N_20781);
nand U23099 (N_23099,N_21958,N_21533);
or U23100 (N_23100,N_21886,N_20936);
xnor U23101 (N_23101,N_20258,N_20186);
xor U23102 (N_23102,N_20100,N_20073);
nor U23103 (N_23103,N_20162,N_21456);
nand U23104 (N_23104,N_21213,N_21399);
nand U23105 (N_23105,N_21016,N_21430);
xnor U23106 (N_23106,N_20982,N_21142);
nor U23107 (N_23107,N_20911,N_21703);
or U23108 (N_23108,N_21018,N_20066);
or U23109 (N_23109,N_20629,N_21289);
or U23110 (N_23110,N_20051,N_20599);
and U23111 (N_23111,N_20286,N_21600);
and U23112 (N_23112,N_20652,N_21876);
and U23113 (N_23113,N_20378,N_21605);
nand U23114 (N_23114,N_20941,N_20206);
nor U23115 (N_23115,N_20319,N_20461);
and U23116 (N_23116,N_20874,N_20260);
nor U23117 (N_23117,N_21504,N_20037);
xor U23118 (N_23118,N_21656,N_21405);
nand U23119 (N_23119,N_21486,N_21043);
or U23120 (N_23120,N_20768,N_20306);
nor U23121 (N_23121,N_21412,N_21987);
nand U23122 (N_23122,N_21566,N_20114);
xnor U23123 (N_23123,N_20361,N_20029);
xnor U23124 (N_23124,N_20416,N_20938);
xnor U23125 (N_23125,N_20933,N_20535);
nor U23126 (N_23126,N_20650,N_21507);
or U23127 (N_23127,N_20078,N_20453);
nor U23128 (N_23128,N_20777,N_21334);
and U23129 (N_23129,N_21271,N_21343);
xor U23130 (N_23130,N_20642,N_20844);
nand U23131 (N_23131,N_21028,N_21527);
nand U23132 (N_23132,N_21312,N_20342);
xor U23133 (N_23133,N_20163,N_21796);
or U23134 (N_23134,N_20809,N_20193);
nor U23135 (N_23135,N_20030,N_20815);
xnor U23136 (N_23136,N_20788,N_21357);
xor U23137 (N_23137,N_21762,N_21322);
or U23138 (N_23138,N_21645,N_21004);
nor U23139 (N_23139,N_20838,N_20799);
or U23140 (N_23140,N_21021,N_21245);
nand U23141 (N_23141,N_20584,N_20562);
or U23142 (N_23142,N_20867,N_21947);
nor U23143 (N_23143,N_20193,N_20418);
xor U23144 (N_23144,N_21904,N_20534);
nor U23145 (N_23145,N_20887,N_20395);
xor U23146 (N_23146,N_20655,N_21696);
nor U23147 (N_23147,N_21786,N_20228);
nor U23148 (N_23148,N_20495,N_21490);
xor U23149 (N_23149,N_21948,N_20091);
nand U23150 (N_23150,N_21655,N_21083);
xnor U23151 (N_23151,N_20669,N_20679);
nand U23152 (N_23152,N_20885,N_20517);
xnor U23153 (N_23153,N_21671,N_20937);
nand U23154 (N_23154,N_20958,N_21332);
or U23155 (N_23155,N_21323,N_21516);
nor U23156 (N_23156,N_21830,N_20880);
nand U23157 (N_23157,N_20916,N_20677);
or U23158 (N_23158,N_21706,N_20878);
xor U23159 (N_23159,N_21564,N_21143);
nor U23160 (N_23160,N_20160,N_20859);
nand U23161 (N_23161,N_20953,N_21622);
nand U23162 (N_23162,N_21571,N_21295);
nand U23163 (N_23163,N_20925,N_21834);
nand U23164 (N_23164,N_21104,N_20478);
nor U23165 (N_23165,N_20890,N_21673);
and U23166 (N_23166,N_20385,N_20965);
or U23167 (N_23167,N_21509,N_20943);
nand U23168 (N_23168,N_20888,N_21466);
or U23169 (N_23169,N_21491,N_21665);
nand U23170 (N_23170,N_21051,N_21942);
nand U23171 (N_23171,N_21022,N_21194);
xor U23172 (N_23172,N_21892,N_20494);
and U23173 (N_23173,N_21588,N_21749);
nor U23174 (N_23174,N_21643,N_21848);
and U23175 (N_23175,N_20093,N_21729);
nor U23176 (N_23176,N_21378,N_20597);
or U23177 (N_23177,N_21646,N_21933);
xnor U23178 (N_23178,N_20277,N_21622);
or U23179 (N_23179,N_20771,N_20442);
nor U23180 (N_23180,N_21942,N_21040);
and U23181 (N_23181,N_21528,N_20433);
or U23182 (N_23182,N_21909,N_20193);
xnor U23183 (N_23183,N_20047,N_21880);
and U23184 (N_23184,N_20408,N_21344);
and U23185 (N_23185,N_20227,N_21349);
nand U23186 (N_23186,N_20675,N_21963);
nand U23187 (N_23187,N_21040,N_21421);
or U23188 (N_23188,N_20981,N_21135);
xor U23189 (N_23189,N_21898,N_21344);
nor U23190 (N_23190,N_21636,N_20156);
nor U23191 (N_23191,N_21627,N_21020);
and U23192 (N_23192,N_21156,N_21899);
xnor U23193 (N_23193,N_20466,N_20947);
or U23194 (N_23194,N_21613,N_20846);
or U23195 (N_23195,N_21153,N_20336);
or U23196 (N_23196,N_21767,N_20175);
nor U23197 (N_23197,N_20738,N_20837);
nand U23198 (N_23198,N_20361,N_21630);
nor U23199 (N_23199,N_21780,N_21016);
or U23200 (N_23200,N_20698,N_21427);
nor U23201 (N_23201,N_21099,N_20209);
nor U23202 (N_23202,N_21627,N_20290);
and U23203 (N_23203,N_20517,N_21063);
nor U23204 (N_23204,N_20381,N_20268);
nor U23205 (N_23205,N_21953,N_21160);
nor U23206 (N_23206,N_21786,N_21316);
or U23207 (N_23207,N_21278,N_20177);
nor U23208 (N_23208,N_20421,N_20561);
nor U23209 (N_23209,N_21452,N_20627);
nand U23210 (N_23210,N_20700,N_21464);
nor U23211 (N_23211,N_21832,N_20645);
nand U23212 (N_23212,N_20283,N_20915);
nand U23213 (N_23213,N_20593,N_20338);
or U23214 (N_23214,N_21773,N_20455);
or U23215 (N_23215,N_21173,N_21177);
xnor U23216 (N_23216,N_20971,N_20742);
xor U23217 (N_23217,N_21365,N_21944);
xor U23218 (N_23218,N_21986,N_20911);
and U23219 (N_23219,N_20588,N_21027);
or U23220 (N_23220,N_21562,N_21697);
and U23221 (N_23221,N_21581,N_20598);
or U23222 (N_23222,N_20938,N_21183);
nand U23223 (N_23223,N_20370,N_21289);
or U23224 (N_23224,N_20572,N_21433);
xnor U23225 (N_23225,N_21202,N_20911);
xor U23226 (N_23226,N_20085,N_21938);
and U23227 (N_23227,N_21201,N_21992);
xor U23228 (N_23228,N_21457,N_21697);
nor U23229 (N_23229,N_20765,N_20556);
or U23230 (N_23230,N_21469,N_20981);
nand U23231 (N_23231,N_20769,N_20842);
or U23232 (N_23232,N_20306,N_20424);
nand U23233 (N_23233,N_20302,N_20119);
and U23234 (N_23234,N_21753,N_20089);
or U23235 (N_23235,N_21880,N_21585);
and U23236 (N_23236,N_21060,N_20346);
nor U23237 (N_23237,N_21696,N_20804);
and U23238 (N_23238,N_20785,N_21653);
nand U23239 (N_23239,N_20135,N_21984);
nand U23240 (N_23240,N_21074,N_21066);
nand U23241 (N_23241,N_20090,N_21007);
nor U23242 (N_23242,N_21576,N_20409);
or U23243 (N_23243,N_21569,N_20642);
and U23244 (N_23244,N_20529,N_21125);
xor U23245 (N_23245,N_20504,N_21386);
nor U23246 (N_23246,N_21171,N_21559);
xnor U23247 (N_23247,N_20515,N_20092);
or U23248 (N_23248,N_21896,N_20334);
or U23249 (N_23249,N_20563,N_21744);
and U23250 (N_23250,N_21195,N_21622);
or U23251 (N_23251,N_20698,N_21051);
nor U23252 (N_23252,N_20559,N_21334);
nand U23253 (N_23253,N_21142,N_21323);
xor U23254 (N_23254,N_20070,N_21367);
nand U23255 (N_23255,N_20889,N_20287);
nor U23256 (N_23256,N_21615,N_20744);
nor U23257 (N_23257,N_20829,N_21309);
or U23258 (N_23258,N_20787,N_20361);
or U23259 (N_23259,N_20366,N_20893);
and U23260 (N_23260,N_21058,N_21770);
or U23261 (N_23261,N_20447,N_21413);
xnor U23262 (N_23262,N_20064,N_21889);
or U23263 (N_23263,N_20333,N_21638);
and U23264 (N_23264,N_21758,N_20656);
xnor U23265 (N_23265,N_21685,N_21152);
xor U23266 (N_23266,N_20721,N_20338);
and U23267 (N_23267,N_20060,N_21095);
nor U23268 (N_23268,N_21860,N_21952);
xnor U23269 (N_23269,N_20423,N_20584);
nand U23270 (N_23270,N_21043,N_21898);
nor U23271 (N_23271,N_20116,N_21096);
or U23272 (N_23272,N_21368,N_21930);
or U23273 (N_23273,N_20922,N_20348);
xor U23274 (N_23274,N_21672,N_21621);
or U23275 (N_23275,N_21578,N_20636);
and U23276 (N_23276,N_20644,N_20260);
nand U23277 (N_23277,N_20365,N_21830);
nand U23278 (N_23278,N_21123,N_20934);
or U23279 (N_23279,N_20214,N_21448);
xnor U23280 (N_23280,N_21219,N_20194);
xnor U23281 (N_23281,N_20024,N_21062);
and U23282 (N_23282,N_20607,N_20034);
nand U23283 (N_23283,N_21391,N_20277);
nor U23284 (N_23284,N_21149,N_21980);
xnor U23285 (N_23285,N_20146,N_20696);
nand U23286 (N_23286,N_21852,N_20573);
xnor U23287 (N_23287,N_20876,N_20206);
or U23288 (N_23288,N_21703,N_20914);
and U23289 (N_23289,N_21793,N_21290);
xnor U23290 (N_23290,N_21983,N_21454);
nor U23291 (N_23291,N_20324,N_20440);
and U23292 (N_23292,N_21301,N_20052);
xnor U23293 (N_23293,N_21121,N_20242);
and U23294 (N_23294,N_20480,N_20620);
or U23295 (N_23295,N_20031,N_20669);
nand U23296 (N_23296,N_20841,N_21077);
nand U23297 (N_23297,N_20183,N_21235);
xnor U23298 (N_23298,N_21394,N_20019);
and U23299 (N_23299,N_21229,N_21795);
nand U23300 (N_23300,N_20968,N_20957);
or U23301 (N_23301,N_20864,N_20649);
and U23302 (N_23302,N_21502,N_20505);
and U23303 (N_23303,N_21471,N_20101);
or U23304 (N_23304,N_20935,N_20100);
and U23305 (N_23305,N_20051,N_20001);
xnor U23306 (N_23306,N_21459,N_20529);
xor U23307 (N_23307,N_21668,N_21427);
nor U23308 (N_23308,N_20305,N_20931);
and U23309 (N_23309,N_20994,N_21046);
or U23310 (N_23310,N_20873,N_20143);
and U23311 (N_23311,N_21252,N_20514);
nand U23312 (N_23312,N_20623,N_20716);
nand U23313 (N_23313,N_21499,N_21220);
nand U23314 (N_23314,N_21371,N_21948);
nand U23315 (N_23315,N_21215,N_20857);
nor U23316 (N_23316,N_21410,N_21352);
or U23317 (N_23317,N_21208,N_20801);
nand U23318 (N_23318,N_20942,N_21397);
and U23319 (N_23319,N_20721,N_20166);
nor U23320 (N_23320,N_21034,N_21358);
nand U23321 (N_23321,N_20919,N_21186);
or U23322 (N_23322,N_20267,N_20509);
or U23323 (N_23323,N_21688,N_20570);
and U23324 (N_23324,N_21501,N_20614);
or U23325 (N_23325,N_20335,N_20791);
xnor U23326 (N_23326,N_20516,N_20837);
xnor U23327 (N_23327,N_20601,N_21437);
or U23328 (N_23328,N_20333,N_21282);
nand U23329 (N_23329,N_21936,N_21346);
and U23330 (N_23330,N_20824,N_20959);
xor U23331 (N_23331,N_20831,N_21845);
and U23332 (N_23332,N_20574,N_20349);
nand U23333 (N_23333,N_20195,N_21745);
or U23334 (N_23334,N_21317,N_21695);
or U23335 (N_23335,N_20617,N_20444);
nor U23336 (N_23336,N_20910,N_21642);
and U23337 (N_23337,N_20810,N_20743);
nor U23338 (N_23338,N_21040,N_21115);
nor U23339 (N_23339,N_20540,N_20871);
nand U23340 (N_23340,N_20696,N_21689);
nand U23341 (N_23341,N_21583,N_20264);
and U23342 (N_23342,N_20677,N_20915);
and U23343 (N_23343,N_20317,N_20624);
nor U23344 (N_23344,N_21197,N_21188);
nand U23345 (N_23345,N_21067,N_20243);
nand U23346 (N_23346,N_20247,N_20256);
xnor U23347 (N_23347,N_20897,N_20088);
xnor U23348 (N_23348,N_21249,N_21023);
nor U23349 (N_23349,N_21145,N_20512);
nand U23350 (N_23350,N_20842,N_20631);
and U23351 (N_23351,N_20467,N_20628);
xnor U23352 (N_23352,N_20729,N_21572);
nand U23353 (N_23353,N_20813,N_21768);
xor U23354 (N_23354,N_20852,N_21616);
or U23355 (N_23355,N_20106,N_21227);
and U23356 (N_23356,N_20818,N_21876);
nand U23357 (N_23357,N_20844,N_21890);
or U23358 (N_23358,N_20588,N_20350);
or U23359 (N_23359,N_20502,N_20752);
nor U23360 (N_23360,N_20776,N_21955);
or U23361 (N_23361,N_20495,N_21893);
or U23362 (N_23362,N_21491,N_21851);
xor U23363 (N_23363,N_21363,N_20449);
nor U23364 (N_23364,N_20521,N_21873);
or U23365 (N_23365,N_20315,N_20387);
or U23366 (N_23366,N_21383,N_21553);
nor U23367 (N_23367,N_21435,N_20141);
xor U23368 (N_23368,N_21867,N_20824);
or U23369 (N_23369,N_21472,N_20133);
nand U23370 (N_23370,N_21540,N_21090);
xor U23371 (N_23371,N_21411,N_21303);
xnor U23372 (N_23372,N_20852,N_20661);
or U23373 (N_23373,N_21745,N_20312);
and U23374 (N_23374,N_20692,N_20021);
nand U23375 (N_23375,N_20983,N_20453);
nor U23376 (N_23376,N_21046,N_20118);
and U23377 (N_23377,N_21422,N_21294);
and U23378 (N_23378,N_20773,N_21426);
xor U23379 (N_23379,N_21208,N_21809);
or U23380 (N_23380,N_21169,N_20504);
xnor U23381 (N_23381,N_20443,N_20537);
nand U23382 (N_23382,N_20026,N_21339);
nand U23383 (N_23383,N_21588,N_21097);
and U23384 (N_23384,N_21899,N_21929);
xor U23385 (N_23385,N_20938,N_20059);
or U23386 (N_23386,N_20201,N_20487);
or U23387 (N_23387,N_21275,N_20773);
nand U23388 (N_23388,N_21801,N_20406);
nor U23389 (N_23389,N_20445,N_20880);
or U23390 (N_23390,N_21963,N_21753);
xnor U23391 (N_23391,N_21333,N_21782);
nand U23392 (N_23392,N_20184,N_21472);
xor U23393 (N_23393,N_21930,N_21447);
or U23394 (N_23394,N_20984,N_20132);
nor U23395 (N_23395,N_20231,N_21960);
and U23396 (N_23396,N_21406,N_21368);
or U23397 (N_23397,N_21108,N_20067);
nor U23398 (N_23398,N_21456,N_20007);
nand U23399 (N_23399,N_20987,N_20991);
nor U23400 (N_23400,N_20860,N_21957);
nand U23401 (N_23401,N_20298,N_21976);
nand U23402 (N_23402,N_20445,N_20868);
nand U23403 (N_23403,N_20526,N_21693);
nor U23404 (N_23404,N_21271,N_20118);
nand U23405 (N_23405,N_20937,N_21004);
nand U23406 (N_23406,N_21787,N_20120);
and U23407 (N_23407,N_21380,N_20689);
nor U23408 (N_23408,N_20824,N_20396);
and U23409 (N_23409,N_21137,N_20061);
nor U23410 (N_23410,N_21364,N_21623);
and U23411 (N_23411,N_21814,N_21960);
xnor U23412 (N_23412,N_20823,N_20299);
nor U23413 (N_23413,N_20442,N_21386);
xnor U23414 (N_23414,N_21965,N_20494);
xor U23415 (N_23415,N_20018,N_21511);
or U23416 (N_23416,N_21279,N_20176);
and U23417 (N_23417,N_20807,N_20964);
nor U23418 (N_23418,N_20506,N_21181);
or U23419 (N_23419,N_20496,N_20896);
and U23420 (N_23420,N_21122,N_21660);
nor U23421 (N_23421,N_20763,N_20320);
nor U23422 (N_23422,N_21246,N_20988);
and U23423 (N_23423,N_20368,N_21697);
xor U23424 (N_23424,N_21094,N_21777);
or U23425 (N_23425,N_21152,N_20047);
nor U23426 (N_23426,N_21452,N_20513);
xor U23427 (N_23427,N_20322,N_21443);
nand U23428 (N_23428,N_21344,N_20067);
xor U23429 (N_23429,N_21639,N_20217);
nor U23430 (N_23430,N_20247,N_21268);
and U23431 (N_23431,N_21368,N_21931);
xor U23432 (N_23432,N_20789,N_21307);
xnor U23433 (N_23433,N_20192,N_20126);
nand U23434 (N_23434,N_21019,N_20786);
nor U23435 (N_23435,N_21904,N_20630);
nand U23436 (N_23436,N_21042,N_20509);
nor U23437 (N_23437,N_21061,N_20495);
nand U23438 (N_23438,N_20459,N_21085);
nor U23439 (N_23439,N_20300,N_21961);
nand U23440 (N_23440,N_21769,N_21347);
or U23441 (N_23441,N_21456,N_20597);
or U23442 (N_23442,N_21129,N_20527);
nor U23443 (N_23443,N_21293,N_21396);
nor U23444 (N_23444,N_20037,N_21208);
nor U23445 (N_23445,N_20053,N_21510);
xnor U23446 (N_23446,N_20667,N_20989);
xnor U23447 (N_23447,N_20897,N_21115);
or U23448 (N_23448,N_20603,N_20544);
xor U23449 (N_23449,N_21893,N_21077);
nor U23450 (N_23450,N_20481,N_20538);
xor U23451 (N_23451,N_21966,N_20199);
nand U23452 (N_23452,N_21592,N_21238);
nor U23453 (N_23453,N_20673,N_21958);
and U23454 (N_23454,N_21339,N_20124);
xor U23455 (N_23455,N_21752,N_21158);
xor U23456 (N_23456,N_20136,N_20493);
and U23457 (N_23457,N_20840,N_20581);
nor U23458 (N_23458,N_20422,N_20187);
or U23459 (N_23459,N_21101,N_21405);
nor U23460 (N_23460,N_21957,N_21395);
nand U23461 (N_23461,N_21573,N_21284);
xor U23462 (N_23462,N_21753,N_20573);
and U23463 (N_23463,N_20816,N_21670);
nor U23464 (N_23464,N_20842,N_21553);
or U23465 (N_23465,N_20182,N_20343);
xnor U23466 (N_23466,N_20202,N_21021);
nand U23467 (N_23467,N_21865,N_20445);
and U23468 (N_23468,N_21665,N_21099);
nor U23469 (N_23469,N_21637,N_21990);
nor U23470 (N_23470,N_21098,N_20505);
nand U23471 (N_23471,N_21621,N_21383);
nand U23472 (N_23472,N_20376,N_21810);
nor U23473 (N_23473,N_20291,N_20627);
or U23474 (N_23474,N_21815,N_21392);
or U23475 (N_23475,N_21381,N_21436);
and U23476 (N_23476,N_20679,N_20396);
nand U23477 (N_23477,N_20846,N_20736);
or U23478 (N_23478,N_20663,N_20015);
and U23479 (N_23479,N_20182,N_21753);
nor U23480 (N_23480,N_21168,N_20569);
xnor U23481 (N_23481,N_21335,N_21112);
and U23482 (N_23482,N_21446,N_20548);
or U23483 (N_23483,N_21627,N_21187);
or U23484 (N_23484,N_20587,N_21343);
nand U23485 (N_23485,N_20794,N_20159);
nand U23486 (N_23486,N_20722,N_20265);
and U23487 (N_23487,N_20782,N_21985);
nand U23488 (N_23488,N_21366,N_20830);
xnor U23489 (N_23489,N_21987,N_20582);
or U23490 (N_23490,N_21649,N_21281);
xor U23491 (N_23491,N_21232,N_20344);
or U23492 (N_23492,N_21134,N_21569);
and U23493 (N_23493,N_20185,N_21783);
nor U23494 (N_23494,N_21896,N_20635);
or U23495 (N_23495,N_21553,N_20352);
xor U23496 (N_23496,N_20444,N_20803);
and U23497 (N_23497,N_21089,N_20304);
nor U23498 (N_23498,N_21374,N_20588);
xor U23499 (N_23499,N_21902,N_21480);
nand U23500 (N_23500,N_20941,N_21693);
nand U23501 (N_23501,N_21418,N_20518);
and U23502 (N_23502,N_21962,N_20161);
xor U23503 (N_23503,N_21677,N_20461);
nor U23504 (N_23504,N_21950,N_21370);
nor U23505 (N_23505,N_20037,N_21545);
xor U23506 (N_23506,N_21395,N_20596);
or U23507 (N_23507,N_20902,N_20732);
xnor U23508 (N_23508,N_20271,N_21000);
or U23509 (N_23509,N_20254,N_21567);
or U23510 (N_23510,N_20304,N_20050);
xnor U23511 (N_23511,N_20085,N_20064);
nand U23512 (N_23512,N_21207,N_21907);
xor U23513 (N_23513,N_21287,N_20666);
xor U23514 (N_23514,N_20566,N_20246);
nor U23515 (N_23515,N_21157,N_21533);
and U23516 (N_23516,N_20062,N_21911);
or U23517 (N_23517,N_21845,N_20972);
xor U23518 (N_23518,N_20850,N_20542);
and U23519 (N_23519,N_20058,N_21926);
nor U23520 (N_23520,N_21255,N_20837);
nand U23521 (N_23521,N_21176,N_20047);
or U23522 (N_23522,N_20941,N_20859);
nand U23523 (N_23523,N_21900,N_20041);
nor U23524 (N_23524,N_20409,N_20739);
xor U23525 (N_23525,N_20374,N_21612);
xnor U23526 (N_23526,N_20162,N_21193);
or U23527 (N_23527,N_20422,N_20807);
or U23528 (N_23528,N_20923,N_21539);
or U23529 (N_23529,N_21095,N_20022);
nor U23530 (N_23530,N_21263,N_20300);
nand U23531 (N_23531,N_20431,N_21309);
nand U23532 (N_23532,N_21096,N_21972);
xnor U23533 (N_23533,N_21035,N_21643);
nor U23534 (N_23534,N_20121,N_21978);
and U23535 (N_23535,N_21335,N_21179);
and U23536 (N_23536,N_20348,N_21448);
or U23537 (N_23537,N_21239,N_20102);
nor U23538 (N_23538,N_20654,N_20497);
xor U23539 (N_23539,N_20994,N_20013);
nand U23540 (N_23540,N_20111,N_21597);
and U23541 (N_23541,N_21562,N_21972);
or U23542 (N_23542,N_21456,N_21754);
nor U23543 (N_23543,N_20476,N_20548);
xnor U23544 (N_23544,N_21082,N_21033);
xor U23545 (N_23545,N_20774,N_21065);
or U23546 (N_23546,N_21222,N_21795);
xor U23547 (N_23547,N_20898,N_21641);
and U23548 (N_23548,N_21781,N_20819);
or U23549 (N_23549,N_21297,N_21175);
xnor U23550 (N_23550,N_21573,N_21515);
nand U23551 (N_23551,N_20066,N_20466);
and U23552 (N_23552,N_21357,N_20178);
xor U23553 (N_23553,N_21405,N_21683);
and U23554 (N_23554,N_21647,N_20139);
xnor U23555 (N_23555,N_21137,N_20056);
and U23556 (N_23556,N_20603,N_21835);
and U23557 (N_23557,N_21656,N_20341);
nor U23558 (N_23558,N_20520,N_20837);
or U23559 (N_23559,N_21421,N_21966);
nand U23560 (N_23560,N_21647,N_20430);
or U23561 (N_23561,N_21895,N_21662);
nor U23562 (N_23562,N_20215,N_21561);
nand U23563 (N_23563,N_21825,N_20016);
and U23564 (N_23564,N_20211,N_20112);
and U23565 (N_23565,N_20039,N_20382);
or U23566 (N_23566,N_21461,N_21082);
and U23567 (N_23567,N_20530,N_20330);
and U23568 (N_23568,N_20822,N_20277);
xnor U23569 (N_23569,N_21370,N_21020);
nor U23570 (N_23570,N_21420,N_21942);
nand U23571 (N_23571,N_20753,N_21178);
xnor U23572 (N_23572,N_20342,N_21917);
xor U23573 (N_23573,N_21165,N_21803);
xnor U23574 (N_23574,N_21614,N_20299);
nand U23575 (N_23575,N_21032,N_21162);
xor U23576 (N_23576,N_20699,N_21028);
nor U23577 (N_23577,N_20838,N_21575);
or U23578 (N_23578,N_20524,N_21047);
nor U23579 (N_23579,N_20876,N_21742);
nand U23580 (N_23580,N_20278,N_20265);
nand U23581 (N_23581,N_21720,N_20650);
and U23582 (N_23582,N_21504,N_21432);
nand U23583 (N_23583,N_21391,N_20645);
xnor U23584 (N_23584,N_20418,N_21217);
nor U23585 (N_23585,N_21174,N_20219);
or U23586 (N_23586,N_21495,N_21402);
or U23587 (N_23587,N_20906,N_20084);
nand U23588 (N_23588,N_21705,N_21770);
nand U23589 (N_23589,N_20513,N_21937);
xor U23590 (N_23590,N_20512,N_21934);
xnor U23591 (N_23591,N_21994,N_21301);
and U23592 (N_23592,N_21565,N_21709);
xor U23593 (N_23593,N_20157,N_21715);
and U23594 (N_23594,N_21247,N_20526);
or U23595 (N_23595,N_21783,N_20427);
nand U23596 (N_23596,N_21334,N_21878);
nand U23597 (N_23597,N_21874,N_20416);
xnor U23598 (N_23598,N_20872,N_21426);
nor U23599 (N_23599,N_21058,N_20459);
nand U23600 (N_23600,N_20372,N_21609);
nor U23601 (N_23601,N_20363,N_21629);
and U23602 (N_23602,N_21464,N_20930);
xnor U23603 (N_23603,N_20544,N_20901);
xor U23604 (N_23604,N_21871,N_21615);
nand U23605 (N_23605,N_21843,N_20251);
nor U23606 (N_23606,N_20167,N_21020);
xnor U23607 (N_23607,N_20073,N_20237);
and U23608 (N_23608,N_21377,N_20616);
nand U23609 (N_23609,N_20088,N_21762);
or U23610 (N_23610,N_21732,N_21431);
or U23611 (N_23611,N_20955,N_20859);
nand U23612 (N_23612,N_21473,N_20272);
or U23613 (N_23613,N_20206,N_20658);
nand U23614 (N_23614,N_21134,N_20661);
nand U23615 (N_23615,N_20095,N_21494);
and U23616 (N_23616,N_20359,N_20480);
nor U23617 (N_23617,N_20335,N_21599);
xor U23618 (N_23618,N_21340,N_20336);
nor U23619 (N_23619,N_21466,N_21272);
nand U23620 (N_23620,N_20381,N_20159);
nor U23621 (N_23621,N_20012,N_20534);
nor U23622 (N_23622,N_20025,N_20809);
or U23623 (N_23623,N_21026,N_20925);
and U23624 (N_23624,N_20318,N_21031);
or U23625 (N_23625,N_21501,N_21019);
or U23626 (N_23626,N_21342,N_21409);
xor U23627 (N_23627,N_21838,N_21702);
and U23628 (N_23628,N_21396,N_21964);
or U23629 (N_23629,N_20133,N_20353);
nand U23630 (N_23630,N_21369,N_21173);
nand U23631 (N_23631,N_21023,N_21504);
and U23632 (N_23632,N_20745,N_21071);
nand U23633 (N_23633,N_21894,N_21031);
or U23634 (N_23634,N_21562,N_20205);
and U23635 (N_23635,N_21099,N_21862);
or U23636 (N_23636,N_20925,N_21483);
nand U23637 (N_23637,N_20486,N_21316);
nand U23638 (N_23638,N_20278,N_20023);
and U23639 (N_23639,N_21139,N_20610);
or U23640 (N_23640,N_20838,N_21441);
and U23641 (N_23641,N_20825,N_20367);
or U23642 (N_23642,N_20347,N_20717);
nor U23643 (N_23643,N_20302,N_21559);
nand U23644 (N_23644,N_21255,N_20246);
and U23645 (N_23645,N_20973,N_20610);
nand U23646 (N_23646,N_20009,N_20489);
nand U23647 (N_23647,N_20504,N_21613);
and U23648 (N_23648,N_21658,N_20668);
nor U23649 (N_23649,N_20666,N_20852);
xnor U23650 (N_23650,N_21962,N_20580);
xnor U23651 (N_23651,N_20300,N_21977);
nor U23652 (N_23652,N_21534,N_20073);
nor U23653 (N_23653,N_21969,N_20634);
nor U23654 (N_23654,N_20739,N_21207);
nand U23655 (N_23655,N_21073,N_20027);
and U23656 (N_23656,N_20809,N_20926);
or U23657 (N_23657,N_20892,N_21189);
or U23658 (N_23658,N_20436,N_20667);
and U23659 (N_23659,N_21018,N_21535);
or U23660 (N_23660,N_20034,N_21576);
and U23661 (N_23661,N_21758,N_21093);
nor U23662 (N_23662,N_21490,N_20058);
xor U23663 (N_23663,N_20426,N_21138);
nand U23664 (N_23664,N_20358,N_20038);
and U23665 (N_23665,N_20749,N_20478);
xor U23666 (N_23666,N_21069,N_21438);
xor U23667 (N_23667,N_21432,N_20520);
nand U23668 (N_23668,N_21873,N_20322);
xor U23669 (N_23669,N_21682,N_20826);
nor U23670 (N_23670,N_20320,N_21753);
nor U23671 (N_23671,N_20497,N_21449);
and U23672 (N_23672,N_20211,N_21010);
nor U23673 (N_23673,N_20988,N_20647);
nor U23674 (N_23674,N_20481,N_21595);
or U23675 (N_23675,N_21000,N_21140);
xnor U23676 (N_23676,N_21561,N_21270);
nor U23677 (N_23677,N_21439,N_21240);
nor U23678 (N_23678,N_20595,N_21366);
or U23679 (N_23679,N_20100,N_21278);
and U23680 (N_23680,N_20281,N_20683);
and U23681 (N_23681,N_21661,N_21721);
nand U23682 (N_23682,N_21497,N_20462);
nand U23683 (N_23683,N_20582,N_21333);
or U23684 (N_23684,N_21273,N_20127);
nor U23685 (N_23685,N_21344,N_20955);
xor U23686 (N_23686,N_20832,N_20232);
or U23687 (N_23687,N_21242,N_20466);
nor U23688 (N_23688,N_21121,N_20889);
nand U23689 (N_23689,N_21348,N_21828);
xnor U23690 (N_23690,N_21476,N_20018);
or U23691 (N_23691,N_21871,N_20421);
nor U23692 (N_23692,N_21188,N_21817);
and U23693 (N_23693,N_21380,N_20207);
xor U23694 (N_23694,N_20770,N_20353);
nand U23695 (N_23695,N_20272,N_20886);
nor U23696 (N_23696,N_21768,N_21898);
xnor U23697 (N_23697,N_21534,N_21935);
or U23698 (N_23698,N_21751,N_20684);
nor U23699 (N_23699,N_21975,N_20953);
xnor U23700 (N_23700,N_20692,N_20482);
nor U23701 (N_23701,N_20877,N_21134);
and U23702 (N_23702,N_21448,N_21443);
nand U23703 (N_23703,N_21430,N_21864);
xnor U23704 (N_23704,N_20930,N_20171);
and U23705 (N_23705,N_20025,N_21781);
and U23706 (N_23706,N_21068,N_21723);
or U23707 (N_23707,N_20789,N_21012);
or U23708 (N_23708,N_20348,N_20321);
xor U23709 (N_23709,N_20784,N_21622);
nor U23710 (N_23710,N_20354,N_20341);
nand U23711 (N_23711,N_20068,N_21196);
or U23712 (N_23712,N_20663,N_21541);
nand U23713 (N_23713,N_21208,N_21764);
xnor U23714 (N_23714,N_21631,N_21584);
and U23715 (N_23715,N_21642,N_21442);
or U23716 (N_23716,N_21385,N_20280);
and U23717 (N_23717,N_20072,N_21915);
nor U23718 (N_23718,N_21180,N_21999);
and U23719 (N_23719,N_21689,N_21774);
and U23720 (N_23720,N_21066,N_20184);
or U23721 (N_23721,N_20932,N_20617);
or U23722 (N_23722,N_21355,N_20550);
xor U23723 (N_23723,N_21303,N_21185);
xor U23724 (N_23724,N_20162,N_20927);
or U23725 (N_23725,N_21659,N_20660);
or U23726 (N_23726,N_20684,N_21620);
or U23727 (N_23727,N_21677,N_21271);
nor U23728 (N_23728,N_20581,N_21044);
or U23729 (N_23729,N_21648,N_20128);
and U23730 (N_23730,N_20285,N_20265);
or U23731 (N_23731,N_20633,N_20906);
nand U23732 (N_23732,N_20762,N_20026);
and U23733 (N_23733,N_20464,N_20869);
xnor U23734 (N_23734,N_20817,N_21872);
and U23735 (N_23735,N_20829,N_21610);
xnor U23736 (N_23736,N_21670,N_21593);
nand U23737 (N_23737,N_20540,N_21096);
nand U23738 (N_23738,N_20906,N_20811);
and U23739 (N_23739,N_21966,N_20693);
nand U23740 (N_23740,N_21535,N_20072);
nand U23741 (N_23741,N_20704,N_20736);
or U23742 (N_23742,N_20838,N_21319);
or U23743 (N_23743,N_21553,N_21287);
and U23744 (N_23744,N_20499,N_21080);
xor U23745 (N_23745,N_21642,N_21854);
and U23746 (N_23746,N_20503,N_21133);
and U23747 (N_23747,N_20371,N_21867);
nor U23748 (N_23748,N_21091,N_20145);
and U23749 (N_23749,N_20820,N_21734);
nor U23750 (N_23750,N_20688,N_20472);
or U23751 (N_23751,N_20563,N_20221);
nand U23752 (N_23752,N_20584,N_20944);
nand U23753 (N_23753,N_21634,N_20162);
and U23754 (N_23754,N_21122,N_20015);
nor U23755 (N_23755,N_21543,N_20457);
nand U23756 (N_23756,N_21791,N_20260);
and U23757 (N_23757,N_21282,N_21988);
or U23758 (N_23758,N_20099,N_20078);
nor U23759 (N_23759,N_21940,N_20622);
xor U23760 (N_23760,N_20366,N_21924);
and U23761 (N_23761,N_20374,N_21726);
or U23762 (N_23762,N_20839,N_21230);
and U23763 (N_23763,N_20828,N_21296);
nor U23764 (N_23764,N_20163,N_21115);
nor U23765 (N_23765,N_21508,N_20412);
or U23766 (N_23766,N_20896,N_21697);
nor U23767 (N_23767,N_20467,N_21660);
nor U23768 (N_23768,N_21014,N_21201);
nor U23769 (N_23769,N_21496,N_21844);
nand U23770 (N_23770,N_21876,N_21748);
or U23771 (N_23771,N_20858,N_21375);
nor U23772 (N_23772,N_20627,N_21023);
or U23773 (N_23773,N_21463,N_20562);
nand U23774 (N_23774,N_21740,N_20508);
nor U23775 (N_23775,N_20264,N_21042);
nand U23776 (N_23776,N_21242,N_21813);
nand U23777 (N_23777,N_20848,N_21155);
or U23778 (N_23778,N_21162,N_21770);
xor U23779 (N_23779,N_20142,N_21410);
or U23780 (N_23780,N_20498,N_21545);
and U23781 (N_23781,N_20030,N_21306);
and U23782 (N_23782,N_20770,N_21320);
xor U23783 (N_23783,N_20807,N_20543);
nand U23784 (N_23784,N_21020,N_21262);
or U23785 (N_23785,N_21780,N_21407);
and U23786 (N_23786,N_20812,N_20862);
nor U23787 (N_23787,N_20855,N_20218);
and U23788 (N_23788,N_21827,N_20231);
or U23789 (N_23789,N_20525,N_21400);
or U23790 (N_23790,N_20662,N_21286);
or U23791 (N_23791,N_21497,N_21048);
nor U23792 (N_23792,N_20588,N_20120);
or U23793 (N_23793,N_21594,N_21503);
and U23794 (N_23794,N_21992,N_20479);
or U23795 (N_23795,N_21338,N_21436);
nand U23796 (N_23796,N_21107,N_21572);
xnor U23797 (N_23797,N_21831,N_21549);
nor U23798 (N_23798,N_20497,N_21562);
xor U23799 (N_23799,N_21192,N_21208);
nand U23800 (N_23800,N_21277,N_20010);
nand U23801 (N_23801,N_20501,N_20282);
nor U23802 (N_23802,N_21301,N_20198);
nor U23803 (N_23803,N_20858,N_21449);
and U23804 (N_23804,N_21163,N_21575);
nand U23805 (N_23805,N_21626,N_20425);
nand U23806 (N_23806,N_21175,N_21292);
xor U23807 (N_23807,N_21599,N_21091);
nand U23808 (N_23808,N_21956,N_20074);
nand U23809 (N_23809,N_21748,N_21621);
and U23810 (N_23810,N_20586,N_21726);
and U23811 (N_23811,N_20819,N_21616);
and U23812 (N_23812,N_20360,N_21303);
nand U23813 (N_23813,N_21025,N_20068);
nor U23814 (N_23814,N_21999,N_20654);
and U23815 (N_23815,N_20173,N_20233);
xnor U23816 (N_23816,N_20966,N_21565);
nand U23817 (N_23817,N_21958,N_20759);
or U23818 (N_23818,N_20238,N_20327);
and U23819 (N_23819,N_20323,N_20229);
nor U23820 (N_23820,N_20101,N_21267);
and U23821 (N_23821,N_21056,N_20553);
and U23822 (N_23822,N_20519,N_21081);
xor U23823 (N_23823,N_21335,N_20494);
nand U23824 (N_23824,N_21289,N_21054);
or U23825 (N_23825,N_21461,N_20435);
and U23826 (N_23826,N_20490,N_20924);
xnor U23827 (N_23827,N_20748,N_21382);
or U23828 (N_23828,N_21729,N_21885);
or U23829 (N_23829,N_20153,N_21476);
or U23830 (N_23830,N_20672,N_20138);
or U23831 (N_23831,N_21914,N_21917);
and U23832 (N_23832,N_20119,N_21069);
xor U23833 (N_23833,N_20343,N_21803);
nand U23834 (N_23834,N_20950,N_21705);
xnor U23835 (N_23835,N_20897,N_21769);
or U23836 (N_23836,N_20409,N_21743);
or U23837 (N_23837,N_21601,N_21621);
xor U23838 (N_23838,N_21575,N_21038);
and U23839 (N_23839,N_21211,N_21420);
xor U23840 (N_23840,N_21075,N_21439);
or U23841 (N_23841,N_20756,N_20793);
and U23842 (N_23842,N_20724,N_21404);
and U23843 (N_23843,N_20872,N_20573);
xnor U23844 (N_23844,N_20010,N_20384);
nor U23845 (N_23845,N_21682,N_20909);
xor U23846 (N_23846,N_20832,N_20862);
or U23847 (N_23847,N_20565,N_20272);
nor U23848 (N_23848,N_21099,N_20398);
nor U23849 (N_23849,N_21213,N_20981);
nor U23850 (N_23850,N_20887,N_21992);
nor U23851 (N_23851,N_21536,N_21895);
nand U23852 (N_23852,N_21127,N_21856);
nand U23853 (N_23853,N_21234,N_20705);
nor U23854 (N_23854,N_21198,N_21295);
and U23855 (N_23855,N_20503,N_21376);
or U23856 (N_23856,N_21090,N_21462);
and U23857 (N_23857,N_20277,N_21837);
or U23858 (N_23858,N_20370,N_20454);
nand U23859 (N_23859,N_21004,N_21906);
nor U23860 (N_23860,N_20632,N_21611);
xor U23861 (N_23861,N_20996,N_21408);
nor U23862 (N_23862,N_20895,N_20465);
or U23863 (N_23863,N_21407,N_20138);
or U23864 (N_23864,N_21208,N_21872);
and U23865 (N_23865,N_20833,N_20338);
nand U23866 (N_23866,N_20831,N_20647);
xor U23867 (N_23867,N_20972,N_21451);
and U23868 (N_23868,N_20846,N_21599);
and U23869 (N_23869,N_20135,N_20076);
nor U23870 (N_23870,N_21065,N_20114);
xnor U23871 (N_23871,N_21094,N_20246);
nand U23872 (N_23872,N_20217,N_20774);
or U23873 (N_23873,N_21184,N_21163);
or U23874 (N_23874,N_20533,N_21262);
nand U23875 (N_23875,N_21036,N_20903);
and U23876 (N_23876,N_21627,N_21281);
or U23877 (N_23877,N_20125,N_21353);
nand U23878 (N_23878,N_20010,N_20930);
nand U23879 (N_23879,N_20726,N_21832);
nand U23880 (N_23880,N_20812,N_21934);
or U23881 (N_23881,N_21505,N_20156);
xor U23882 (N_23882,N_20718,N_20557);
nand U23883 (N_23883,N_21451,N_21467);
nor U23884 (N_23884,N_21357,N_21306);
nor U23885 (N_23885,N_21685,N_20085);
and U23886 (N_23886,N_21526,N_20395);
and U23887 (N_23887,N_20524,N_20009);
nor U23888 (N_23888,N_20230,N_21157);
nand U23889 (N_23889,N_20992,N_21261);
nor U23890 (N_23890,N_21506,N_20530);
nand U23891 (N_23891,N_21758,N_21889);
xor U23892 (N_23892,N_21832,N_20452);
nor U23893 (N_23893,N_20684,N_20562);
and U23894 (N_23894,N_21543,N_21580);
nor U23895 (N_23895,N_21390,N_20930);
nor U23896 (N_23896,N_21995,N_20345);
nand U23897 (N_23897,N_21431,N_20458);
nor U23898 (N_23898,N_21923,N_20340);
nand U23899 (N_23899,N_21893,N_20030);
nor U23900 (N_23900,N_20203,N_20267);
nor U23901 (N_23901,N_20163,N_21540);
nor U23902 (N_23902,N_20593,N_20358);
nand U23903 (N_23903,N_21941,N_21646);
nand U23904 (N_23904,N_21233,N_20282);
xor U23905 (N_23905,N_21191,N_20603);
nor U23906 (N_23906,N_21852,N_20981);
and U23907 (N_23907,N_20455,N_21357);
or U23908 (N_23908,N_21416,N_21922);
or U23909 (N_23909,N_20909,N_20464);
xnor U23910 (N_23910,N_20270,N_20465);
and U23911 (N_23911,N_20441,N_21731);
xnor U23912 (N_23912,N_20342,N_21923);
nor U23913 (N_23913,N_21531,N_20283);
xor U23914 (N_23914,N_21438,N_21292);
xor U23915 (N_23915,N_21006,N_21344);
and U23916 (N_23916,N_21882,N_21549);
xor U23917 (N_23917,N_20508,N_21313);
nand U23918 (N_23918,N_21130,N_20868);
and U23919 (N_23919,N_20984,N_21216);
xor U23920 (N_23920,N_20484,N_21325);
and U23921 (N_23921,N_20397,N_21826);
or U23922 (N_23922,N_20479,N_21391);
nor U23923 (N_23923,N_21289,N_20037);
nor U23924 (N_23924,N_21461,N_20275);
nand U23925 (N_23925,N_20305,N_21704);
nand U23926 (N_23926,N_20282,N_21648);
and U23927 (N_23927,N_20861,N_20688);
nor U23928 (N_23928,N_21445,N_20751);
and U23929 (N_23929,N_21786,N_21667);
and U23930 (N_23930,N_21244,N_21483);
or U23931 (N_23931,N_20745,N_21007);
xor U23932 (N_23932,N_21781,N_21443);
nand U23933 (N_23933,N_20943,N_21324);
nor U23934 (N_23934,N_21382,N_20751);
and U23935 (N_23935,N_20484,N_21618);
xnor U23936 (N_23936,N_21956,N_20502);
nand U23937 (N_23937,N_20987,N_21258);
nand U23938 (N_23938,N_21206,N_21747);
xnor U23939 (N_23939,N_21689,N_21388);
nor U23940 (N_23940,N_21684,N_20096);
and U23941 (N_23941,N_20923,N_20297);
nand U23942 (N_23942,N_20755,N_20455);
xor U23943 (N_23943,N_20399,N_21722);
xor U23944 (N_23944,N_21415,N_21232);
or U23945 (N_23945,N_20623,N_20036);
and U23946 (N_23946,N_20954,N_21085);
and U23947 (N_23947,N_20039,N_20650);
xor U23948 (N_23948,N_20005,N_21751);
or U23949 (N_23949,N_20595,N_20664);
nand U23950 (N_23950,N_21188,N_20200);
nor U23951 (N_23951,N_21567,N_21540);
nor U23952 (N_23952,N_20534,N_21397);
xnor U23953 (N_23953,N_20674,N_21242);
and U23954 (N_23954,N_20402,N_20661);
nand U23955 (N_23955,N_20522,N_21785);
nor U23956 (N_23956,N_21146,N_21577);
or U23957 (N_23957,N_20570,N_21555);
xnor U23958 (N_23958,N_20390,N_21120);
nor U23959 (N_23959,N_21816,N_21295);
xor U23960 (N_23960,N_20088,N_21606);
and U23961 (N_23961,N_21473,N_20793);
xor U23962 (N_23962,N_21795,N_20686);
nand U23963 (N_23963,N_20817,N_21561);
and U23964 (N_23964,N_20618,N_21064);
and U23965 (N_23965,N_20757,N_20780);
nor U23966 (N_23966,N_20551,N_20809);
or U23967 (N_23967,N_21266,N_20170);
nand U23968 (N_23968,N_20852,N_20296);
xnor U23969 (N_23969,N_21717,N_20604);
xnor U23970 (N_23970,N_20811,N_21887);
and U23971 (N_23971,N_21441,N_21359);
nor U23972 (N_23972,N_20839,N_20836);
and U23973 (N_23973,N_21422,N_21870);
nor U23974 (N_23974,N_21019,N_21853);
and U23975 (N_23975,N_20903,N_21802);
xnor U23976 (N_23976,N_20674,N_20711);
or U23977 (N_23977,N_20956,N_20460);
nor U23978 (N_23978,N_20229,N_20755);
nand U23979 (N_23979,N_21832,N_21514);
and U23980 (N_23980,N_21874,N_20941);
nor U23981 (N_23981,N_21538,N_21243);
or U23982 (N_23982,N_21290,N_20696);
or U23983 (N_23983,N_20914,N_21070);
and U23984 (N_23984,N_21890,N_21848);
and U23985 (N_23985,N_20984,N_20739);
and U23986 (N_23986,N_21137,N_20874);
or U23987 (N_23987,N_21634,N_20014);
nor U23988 (N_23988,N_20700,N_21237);
nor U23989 (N_23989,N_20183,N_21631);
nand U23990 (N_23990,N_20716,N_20293);
nand U23991 (N_23991,N_21202,N_21244);
nor U23992 (N_23992,N_21917,N_20556);
xor U23993 (N_23993,N_20599,N_20459);
nor U23994 (N_23994,N_20378,N_21679);
nand U23995 (N_23995,N_21069,N_21678);
or U23996 (N_23996,N_21374,N_20664);
xnor U23997 (N_23997,N_20330,N_20827);
xor U23998 (N_23998,N_21570,N_20015);
nand U23999 (N_23999,N_20447,N_20438);
or U24000 (N_24000,N_23139,N_22557);
xor U24001 (N_24001,N_22114,N_23159);
nor U24002 (N_24002,N_22126,N_23121);
or U24003 (N_24003,N_22132,N_22334);
or U24004 (N_24004,N_23356,N_23216);
nand U24005 (N_24005,N_22220,N_22675);
nand U24006 (N_24006,N_22714,N_23850);
or U24007 (N_24007,N_22339,N_23550);
or U24008 (N_24008,N_23636,N_23720);
or U24009 (N_24009,N_23743,N_22036);
nor U24010 (N_24010,N_22607,N_23515);
nand U24011 (N_24011,N_23621,N_22191);
or U24012 (N_24012,N_23337,N_22628);
nand U24013 (N_24013,N_23832,N_23995);
nand U24014 (N_24014,N_23481,N_22273);
or U24015 (N_24015,N_23145,N_22935);
nand U24016 (N_24016,N_22410,N_23570);
or U24017 (N_24017,N_23360,N_22679);
and U24018 (N_24018,N_23651,N_23721);
or U24019 (N_24019,N_23306,N_23906);
nor U24020 (N_24020,N_22186,N_22544);
and U24021 (N_24021,N_22795,N_23050);
nor U24022 (N_24022,N_23445,N_23891);
nor U24023 (N_24023,N_23351,N_22589);
or U24024 (N_24024,N_22020,N_23184);
or U24025 (N_24025,N_22119,N_22377);
nand U24026 (N_24026,N_22025,N_23553);
xnor U24027 (N_24027,N_22817,N_23887);
nor U24028 (N_24028,N_22034,N_23375);
or U24029 (N_24029,N_22963,N_22363);
or U24030 (N_24030,N_23182,N_23158);
xnor U24031 (N_24031,N_22670,N_22088);
xnor U24032 (N_24032,N_22396,N_23512);
or U24033 (N_24033,N_22098,N_23770);
nor U24034 (N_24034,N_22669,N_22303);
and U24035 (N_24035,N_22414,N_23626);
nor U24036 (N_24036,N_23775,N_23568);
nand U24037 (N_24037,N_22183,N_22967);
nand U24038 (N_24038,N_23628,N_23263);
and U24039 (N_24039,N_22107,N_22285);
and U24040 (N_24040,N_22089,N_22786);
nor U24041 (N_24041,N_22282,N_22121);
nor U24042 (N_24042,N_22755,N_22968);
xnor U24043 (N_24043,N_23298,N_23187);
xnor U24044 (N_24044,N_23110,N_22863);
and U24045 (N_24045,N_23135,N_23190);
xor U24046 (N_24046,N_22641,N_22490);
nor U24047 (N_24047,N_22867,N_22317);
nand U24048 (N_24048,N_22274,N_22065);
nand U24049 (N_24049,N_22644,N_22151);
xnor U24050 (N_24050,N_22123,N_22656);
nor U24051 (N_24051,N_23044,N_22927);
xor U24052 (N_24052,N_23999,N_22615);
or U24053 (N_24053,N_23986,N_22995);
xnor U24054 (N_24054,N_23754,N_22591);
or U24055 (N_24055,N_23542,N_23885);
or U24056 (N_24056,N_23672,N_23259);
nand U24057 (N_24057,N_22320,N_22115);
and U24058 (N_24058,N_22150,N_22781);
nor U24059 (N_24059,N_22987,N_23883);
or U24060 (N_24060,N_23300,N_23059);
and U24061 (N_24061,N_23088,N_23027);
xor U24062 (N_24062,N_22224,N_23632);
xnor U24063 (N_24063,N_22402,N_22267);
nand U24064 (N_24064,N_23820,N_22925);
xor U24065 (N_24065,N_22019,N_23400);
nor U24066 (N_24066,N_23700,N_23489);
or U24067 (N_24067,N_23012,N_23544);
and U24068 (N_24068,N_22582,N_22000);
nor U24069 (N_24069,N_23030,N_22524);
nor U24070 (N_24070,N_22188,N_23691);
nand U24071 (N_24071,N_23797,N_23505);
or U24072 (N_24072,N_22821,N_23105);
xor U24073 (N_24073,N_23666,N_23742);
nand U24074 (N_24074,N_22558,N_23554);
xnor U24075 (N_24075,N_22498,N_22972);
and U24076 (N_24076,N_23177,N_22555);
nor U24077 (N_24077,N_22462,N_22838);
nand U24078 (N_24078,N_23443,N_22620);
nand U24079 (N_24079,N_23884,N_22773);
nor U24080 (N_24080,N_22829,N_22276);
or U24081 (N_24081,N_22057,N_22044);
and U24082 (N_24082,N_23384,N_22213);
nor U24083 (N_24083,N_22027,N_22288);
xnor U24084 (N_24084,N_22697,N_22311);
nor U24085 (N_24085,N_22031,N_22808);
nand U24086 (N_24086,N_23085,N_22793);
or U24087 (N_24087,N_23451,N_23004);
nand U24088 (N_24088,N_22281,N_23486);
xnor U24089 (N_24089,N_22194,N_23291);
nand U24090 (N_24090,N_22789,N_22278);
nor U24091 (N_24091,N_22102,N_23602);
nand U24092 (N_24092,N_23450,N_23961);
nand U24093 (N_24093,N_23620,N_23146);
or U24094 (N_24094,N_23881,N_23423);
and U24095 (N_24095,N_22095,N_22624);
and U24096 (N_24096,N_22051,N_23677);
or U24097 (N_24097,N_22949,N_23985);
xor U24098 (N_24098,N_23051,N_22295);
and U24099 (N_24099,N_23296,N_22309);
nor U24100 (N_24100,N_22692,N_23468);
and U24101 (N_24101,N_22042,N_22638);
nor U24102 (N_24102,N_23664,N_22212);
xnor U24103 (N_24103,N_22852,N_22242);
and U24104 (N_24104,N_23010,N_22552);
and U24105 (N_24105,N_23487,N_23814);
nor U24106 (N_24106,N_22381,N_22672);
nand U24107 (N_24107,N_22956,N_23740);
nor U24108 (N_24108,N_23975,N_23239);
or U24109 (N_24109,N_22064,N_23449);
nand U24110 (N_24110,N_22622,N_23096);
nor U24111 (N_24111,N_23840,N_23327);
nor U24112 (N_24112,N_23455,N_23822);
xnor U24113 (N_24113,N_22520,N_22342);
or U24114 (N_24114,N_22217,N_23900);
or U24115 (N_24115,N_23024,N_23454);
nor U24116 (N_24116,N_23957,N_23996);
xnor U24117 (N_24117,N_23582,N_23649);
xnor U24118 (N_24118,N_23000,N_23644);
nand U24119 (N_24119,N_22709,N_23907);
nor U24120 (N_24120,N_22120,N_23112);
or U24121 (N_24121,N_22237,N_23001);
nand U24122 (N_24122,N_23175,N_23904);
nand U24123 (N_24123,N_23988,N_23396);
xnor U24124 (N_24124,N_23790,N_23252);
or U24125 (N_24125,N_23330,N_23625);
or U24126 (N_24126,N_22354,N_23739);
and U24127 (N_24127,N_23359,N_23751);
nand U24128 (N_24128,N_22360,N_22685);
nor U24129 (N_24129,N_23962,N_23583);
or U24130 (N_24130,N_22657,N_23727);
nand U24131 (N_24131,N_22355,N_22594);
and U24132 (N_24132,N_23765,N_23747);
nor U24133 (N_24133,N_23695,N_22207);
nor U24134 (N_24134,N_23997,N_23369);
nand U24135 (N_24135,N_23439,N_23040);
nor U24136 (N_24136,N_22730,N_22632);
and U24137 (N_24137,N_22144,N_22668);
and U24138 (N_24138,N_23914,N_22616);
and U24139 (N_24139,N_22386,N_23331);
or U24140 (N_24140,N_22945,N_23075);
nand U24141 (N_24141,N_22055,N_23971);
nor U24142 (N_24142,N_22171,N_22388);
or U24143 (N_24143,N_23277,N_23854);
and U24144 (N_24144,N_22599,N_23825);
and U24145 (N_24145,N_22747,N_22340);
or U24146 (N_24146,N_22086,N_22008);
or U24147 (N_24147,N_22943,N_23471);
and U24148 (N_24148,N_23039,N_23188);
nor U24149 (N_24149,N_23019,N_22646);
nor U24150 (N_24150,N_23744,N_23060);
and U24151 (N_24151,N_23234,N_22313);
or U24152 (N_24152,N_22412,N_22152);
nor U24153 (N_24153,N_22459,N_23206);
or U24154 (N_24154,N_23398,N_23572);
nor U24155 (N_24155,N_22874,N_22181);
nand U24156 (N_24156,N_23577,N_23799);
xnor U24157 (N_24157,N_23448,N_22455);
and U24158 (N_24158,N_22839,N_22897);
or U24159 (N_24159,N_22523,N_23596);
nor U24160 (N_24160,N_23976,N_22227);
nor U24161 (N_24161,N_23475,N_22235);
xor U24162 (N_24162,N_23134,N_22940);
xnor U24163 (N_24163,N_22353,N_23103);
xor U24164 (N_24164,N_22296,N_22919);
xnor U24165 (N_24165,N_23686,N_23750);
nand U24166 (N_24166,N_23061,N_23438);
and U24167 (N_24167,N_22606,N_23054);
nand U24168 (N_24168,N_23590,N_23437);
and U24169 (N_24169,N_23560,N_22247);
xnor U24170 (N_24170,N_22976,N_22545);
or U24171 (N_24171,N_23511,N_22483);
nor U24172 (N_24172,N_23519,N_22394);
nand U24173 (N_24173,N_23767,N_23580);
nand U24174 (N_24174,N_22372,N_23682);
nand U24175 (N_24175,N_23735,N_22085);
and U24176 (N_24176,N_22243,N_23089);
and U24177 (N_24177,N_23414,N_23167);
xnor U24178 (N_24178,N_23482,N_23757);
and U24179 (N_24179,N_22040,N_22813);
xor U24180 (N_24180,N_23851,N_22752);
or U24181 (N_24181,N_22994,N_22571);
nand U24182 (N_24182,N_23272,N_22587);
or U24183 (N_24183,N_23616,N_22305);
nor U24184 (N_24184,N_23989,N_22634);
nand U24185 (N_24185,N_22422,N_23074);
and U24186 (N_24186,N_22988,N_23547);
xor U24187 (N_24187,N_23063,N_22712);
and U24188 (N_24188,N_23782,N_22721);
xor U24189 (N_24189,N_23631,N_22068);
or U24190 (N_24190,N_23275,N_23802);
xor U24191 (N_24191,N_23240,N_23416);
or U24192 (N_24192,N_22535,N_23132);
or U24193 (N_24193,N_22741,N_23441);
or U24194 (N_24194,N_23753,N_23761);
and U24195 (N_24195,N_23670,N_23502);
and U24196 (N_24196,N_23836,N_23779);
xor U24197 (N_24197,N_23383,N_23588);
and U24198 (N_24198,N_22516,N_22190);
or U24199 (N_24199,N_22087,N_23053);
nor U24200 (N_24200,N_23232,N_22700);
xnor U24201 (N_24201,N_22573,N_22018);
xnor U24202 (N_24202,N_22833,N_22491);
xor U24203 (N_24203,N_22200,N_23212);
xnor U24204 (N_24204,N_22233,N_22210);
nor U24205 (N_24205,N_22836,N_22985);
nand U24206 (N_24206,N_22508,N_22928);
and U24207 (N_24207,N_22333,N_23160);
xor U24208 (N_24208,N_22671,N_22447);
nand U24209 (N_24209,N_23784,N_23311);
nand U24210 (N_24210,N_22058,N_22173);
nand U24211 (N_24211,N_22827,N_22708);
and U24212 (N_24212,N_22244,N_23788);
or U24213 (N_24213,N_22739,N_23335);
xor U24214 (N_24214,N_22914,N_22862);
or U24215 (N_24215,N_22439,N_23425);
and U24216 (N_24216,N_22451,N_22532);
and U24217 (N_24217,N_23038,N_22865);
or U24218 (N_24218,N_22078,N_22264);
or U24219 (N_24219,N_22289,N_23114);
xor U24220 (N_24220,N_23133,N_22918);
or U24221 (N_24221,N_23610,N_22978);
nor U24222 (N_24222,N_23237,N_23390);
and U24223 (N_24223,N_23174,N_22780);
or U24224 (N_24224,N_22691,N_22134);
nor U24225 (N_24225,N_23849,N_23915);
or U24226 (N_24226,N_22346,N_23302);
nand U24227 (N_24227,N_22604,N_23342);
xnor U24228 (N_24228,N_22769,N_23090);
xor U24229 (N_24229,N_23338,N_22890);
and U24230 (N_24230,N_23729,N_22600);
and U24231 (N_24231,N_23171,N_23181);
and U24232 (N_24232,N_23941,N_23269);
or U24233 (N_24233,N_22218,N_23650);
nand U24234 (N_24234,N_22562,N_22481);
and U24235 (N_24235,N_22093,N_22383);
or U24236 (N_24236,N_23473,N_23172);
or U24237 (N_24237,N_22054,N_23320);
and U24238 (N_24238,N_23477,N_22478);
xnor U24239 (N_24239,N_22876,N_22291);
and U24240 (N_24240,N_23698,N_22182);
or U24241 (N_24241,N_22767,N_22053);
nand U24242 (N_24242,N_23209,N_23816);
and U24243 (N_24243,N_22735,N_22645);
nand U24244 (N_24244,N_22999,N_22837);
nand U24245 (N_24245,N_23407,N_22260);
or U24246 (N_24246,N_23210,N_23737);
or U24247 (N_24247,N_23215,N_22787);
nand U24248 (N_24248,N_22579,N_23122);
xnor U24249 (N_24249,N_22407,N_22762);
xnor U24250 (N_24250,N_23453,N_23857);
and U24251 (N_24251,N_22393,N_23864);
nand U24252 (N_24252,N_22184,N_23707);
xor U24253 (N_24253,N_23645,N_22122);
xor U24254 (N_24254,N_23049,N_22842);
xnor U24255 (N_24255,N_23768,N_22596);
and U24256 (N_24256,N_23657,N_23391);
or U24257 (N_24257,N_22778,N_23927);
nor U24258 (N_24258,N_22379,N_23618);
xnor U24259 (N_24259,N_22900,N_22467);
nor U24260 (N_24260,N_23260,N_22610);
nand U24261 (N_24261,N_23401,N_23348);
and U24262 (N_24262,N_22905,N_23523);
or U24263 (N_24263,N_23942,N_22921);
and U24264 (N_24264,N_22888,N_23633);
nor U24265 (N_24265,N_22546,N_22488);
and U24266 (N_24266,N_23289,N_23591);
and U24267 (N_24267,N_22626,N_22648);
nand U24268 (N_24268,N_23556,N_22933);
or U24269 (N_24269,N_22667,N_23752);
or U24270 (N_24270,N_23339,N_23783);
and U24271 (N_24271,N_23658,N_23460);
nor U24272 (N_24272,N_22209,N_23980);
and U24273 (N_24273,N_23009,N_22984);
or U24274 (N_24274,N_22323,N_23611);
or U24275 (N_24275,N_23222,N_23073);
nor U24276 (N_24276,N_23086,N_23329);
and U24277 (N_24277,N_22618,N_23336);
or U24278 (N_24278,N_22050,N_23969);
nand U24279 (N_24279,N_22856,N_23913);
nand U24280 (N_24280,N_23594,N_22981);
or U24281 (N_24281,N_22986,N_23678);
nand U24282 (N_24282,N_23756,N_22961);
or U24283 (N_24283,N_22904,N_23424);
xnor U24284 (N_24284,N_22306,N_22815);
or U24285 (N_24285,N_22497,N_23080);
or U24286 (N_24286,N_22344,N_22153);
nand U24287 (N_24287,N_22954,N_23166);
nor U24288 (N_24288,N_22814,N_23305);
nand U24289 (N_24289,N_22629,N_22090);
nor U24290 (N_24290,N_23253,N_22045);
or U24291 (N_24291,N_22436,N_23429);
or U24292 (N_24292,N_23943,N_23608);
and U24293 (N_24293,N_22633,N_23340);
and U24294 (N_24294,N_23373,N_22895);
or U24295 (N_24295,N_23071,N_22015);
and U24296 (N_24296,N_22105,N_22899);
and U24297 (N_24297,N_22109,N_23101);
xor U24298 (N_24298,N_23521,N_22418);
nor U24299 (N_24299,N_23223,N_22548);
nor U24300 (N_24300,N_22902,N_23692);
nand U24301 (N_24301,N_23273,N_22387);
nand U24302 (N_24302,N_22373,N_23680);
and U24303 (N_24303,N_22142,N_23876);
xnor U24304 (N_24304,N_22300,N_22732);
and U24305 (N_24305,N_23548,N_23806);
nand U24306 (N_24306,N_23108,N_23909);
nor U24307 (N_24307,N_23669,N_22328);
or U24308 (N_24308,N_22238,N_22137);
or U24309 (N_24309,N_22970,N_23056);
and U24310 (N_24310,N_22920,N_23270);
nor U24311 (N_24311,N_23488,N_23444);
or U24312 (N_24312,N_23880,N_22798);
or U24313 (N_24313,N_22229,N_23815);
or U24314 (N_24314,N_22463,N_22403);
nor U24315 (N_24315,N_22319,N_22287);
xor U24316 (N_24316,N_22683,N_22777);
nor U24317 (N_24317,N_23592,N_23821);
xor U24318 (N_24318,N_23042,N_23295);
xnor U24319 (N_24319,N_23893,N_22799);
nand U24320 (N_24320,N_23274,N_23852);
nand U24321 (N_24321,N_22775,N_23409);
xnor U24322 (N_24322,N_23358,N_22430);
or U24323 (N_24323,N_23624,N_22368);
and U24324 (N_24324,N_23354,N_22024);
xor U24325 (N_24325,N_22026,N_22887);
or U24326 (N_24326,N_22215,N_22621);
or U24327 (N_24327,N_23065,N_23813);
xnor U24328 (N_24328,N_22258,N_22894);
and U24329 (N_24329,N_22770,N_22757);
or U24330 (N_24330,N_22441,N_22494);
nor U24331 (N_24331,N_22469,N_22681);
nor U24332 (N_24332,N_22704,N_23955);
nand U24333 (N_24333,N_23224,N_22138);
xnor U24334 (N_24334,N_22653,N_22595);
nor U24335 (N_24335,N_23839,N_22046);
and U24336 (N_24336,N_23413,N_22160);
and U24337 (N_24337,N_23285,N_23665);
or U24338 (N_24338,N_22371,N_23655);
nor U24339 (N_24339,N_22140,N_22128);
nand U24340 (N_24340,N_22879,N_23983);
nand U24341 (N_24341,N_22245,N_22745);
xor U24342 (N_24342,N_23227,N_23531);
or U24343 (N_24343,N_22642,N_22841);
nor U24344 (N_24344,N_23702,N_23077);
and U24345 (N_24345,N_22030,N_23130);
and U24346 (N_24346,N_23901,N_23829);
nor U24347 (N_24347,N_23992,N_23192);
nor U24348 (N_24348,N_23169,N_22614);
and U24349 (N_24349,N_23036,N_23771);
xor U24350 (N_24350,N_23922,N_23524);
nor U24351 (N_24351,N_22710,N_23609);
nor U24352 (N_24352,N_23123,N_23179);
or U24353 (N_24353,N_23431,N_23456);
xor U24354 (N_24354,N_23968,N_22415);
nor U24355 (N_24355,N_22010,N_23510);
nand U24356 (N_24356,N_22947,N_23731);
nand U24357 (N_24357,N_22248,N_22885);
and U24358 (N_24358,N_23977,N_23026);
xnor U24359 (N_24359,N_22804,N_23235);
nand U24360 (N_24360,N_23613,N_22973);
or U24361 (N_24361,N_22146,N_23860);
nor U24362 (N_24362,N_22977,N_23370);
xor U24363 (N_24363,N_22964,N_23203);
or U24364 (N_24364,N_23705,N_23043);
nand U24365 (N_24365,N_22314,N_22543);
nor U24366 (N_24366,N_22910,N_23417);
nor U24367 (N_24367,N_23319,N_22529);
nor U24368 (N_24368,N_22574,N_23083);
and U24369 (N_24369,N_22148,N_22823);
or U24370 (N_24370,N_22851,N_23619);
nor U24371 (N_24371,N_22864,N_22004);
and U24372 (N_24372,N_23956,N_22484);
xnor U24373 (N_24373,N_23341,N_23662);
nand U24374 (N_24374,N_22435,N_23574);
nand U24375 (N_24375,N_23748,N_23102);
and U24376 (N_24376,N_23377,N_22909);
nand U24377 (N_24377,N_22991,N_22647);
nor U24378 (N_24378,N_22674,N_22474);
or U24379 (N_24379,N_22974,N_23925);
xor U24380 (N_24380,N_23463,N_23264);
xor U24381 (N_24381,N_23923,N_22052);
and U24382 (N_24382,N_23006,N_22992);
xor U24383 (N_24383,N_22500,N_23346);
and U24384 (N_24384,N_23379,N_23722);
nand U24385 (N_24385,N_23792,N_23536);
nand U24386 (N_24386,N_22577,N_23048);
or U24387 (N_24387,N_22660,N_22738);
or U24388 (N_24388,N_23343,N_22039);
nor U24389 (N_24389,N_22566,N_22601);
nand U24390 (N_24390,N_22416,N_23787);
nor U24391 (N_24391,N_23565,N_23776);
xnor U24392 (N_24392,N_23474,N_23738);
nand U24393 (N_24393,N_22161,N_23462);
or U24394 (N_24394,N_22445,N_23066);
and U24395 (N_24395,N_23562,N_22286);
or U24396 (N_24396,N_22680,N_22965);
xnor U24397 (N_24397,N_23890,N_22056);
xnor U24398 (N_24398,N_23525,N_23875);
xor U24399 (N_24399,N_23938,N_22017);
nor U24400 (N_24400,N_23954,N_22794);
nor U24401 (N_24401,N_22005,N_22944);
nor U24402 (N_24402,N_22756,N_23310);
nand U24403 (N_24403,N_23810,N_23516);
nor U24404 (N_24404,N_22203,N_23877);
xnor U24405 (N_24405,N_22409,N_23869);
and U24406 (N_24406,N_23945,N_23571);
or U24407 (N_24407,N_23663,N_23388);
and U24408 (N_24408,N_22982,N_22619);
and U24409 (N_24409,N_23903,N_22734);
nand U24410 (N_24410,N_23501,N_23419);
xor U24411 (N_24411,N_22460,N_22012);
xor U24412 (N_24412,N_22256,N_23733);
nand U24413 (N_24413,N_22617,N_23758);
xnor U24414 (N_24414,N_23076,N_23898);
nor U24415 (N_24415,N_22830,N_23585);
nand U24416 (N_24416,N_23189,N_23365);
xor U24417 (N_24417,N_22728,N_22292);
xnor U24418 (N_24418,N_22417,N_22891);
and U24419 (N_24419,N_22468,N_22406);
or U24420 (N_24420,N_22419,N_22263);
nand U24421 (N_24421,N_22784,N_23461);
nand U24422 (N_24422,N_22609,N_22037);
xnor U24423 (N_24423,N_22421,N_22092);
nand U24424 (N_24424,N_23848,N_23213);
or U24425 (N_24425,N_22958,N_22828);
and U24426 (N_24426,N_22438,N_22711);
nor U24427 (N_24427,N_22788,N_23315);
nand U24428 (N_24428,N_22850,N_22272);
xor U24429 (N_24429,N_23011,N_23833);
xor U24430 (N_24430,N_22509,N_22916);
and U24431 (N_24431,N_23458,N_23364);
or U24432 (N_24432,N_22826,N_23917);
or U24433 (N_24433,N_22774,N_22312);
or U24434 (N_24434,N_23068,N_23948);
nand U24435 (N_24435,N_22101,N_23126);
or U24436 (N_24436,N_22446,N_22597);
and U24437 (N_24437,N_23694,N_23667);
and U24438 (N_24438,N_23973,N_22689);
xnor U24439 (N_24439,N_23704,N_23967);
nor U24440 (N_24440,N_23124,N_22521);
nand U24441 (N_24441,N_23428,N_23452);
xnor U24442 (N_24442,N_22007,N_23207);
or U24443 (N_24443,N_23764,N_23991);
or U24444 (N_24444,N_22458,N_22185);
and U24445 (N_24445,N_22743,N_23037);
or U24446 (N_24446,N_22433,N_23817);
xnor U24447 (N_24447,N_22047,N_23022);
nor U24448 (N_24448,N_23870,N_22649);
and U24449 (N_24449,N_23144,N_22676);
and U24450 (N_24450,N_22650,N_23057);
nand U24451 (N_24451,N_23882,N_23229);
xnor U24452 (N_24452,N_22365,N_23293);
nand U24453 (N_24453,N_23023,N_22719);
nor U24454 (N_24454,N_22541,N_22753);
nand U24455 (N_24455,N_22698,N_22576);
or U24456 (N_24456,N_23500,N_23479);
nor U24457 (N_24457,N_22448,N_22096);
or U24458 (N_24458,N_23578,N_22136);
xor U24459 (N_24459,N_22080,N_23303);
xor U24460 (N_24460,N_23367,N_23828);
nand U24461 (N_24461,N_22389,N_23490);
and U24462 (N_24462,N_23033,N_23879);
nor U24463 (N_24463,N_22746,N_22907);
xor U24464 (N_24464,N_23537,N_22565);
nor U24465 (N_24465,N_23408,N_22104);
nand U24466 (N_24466,N_22337,N_22812);
xor U24467 (N_24467,N_22765,N_23557);
nor U24468 (N_24468,N_23469,N_22575);
xnor U24469 (N_24469,N_22528,N_22860);
xor U24470 (N_24470,N_22208,N_22375);
or U24471 (N_24471,N_22326,N_22911);
and U24472 (N_24472,N_22835,N_23862);
nand U24473 (N_24473,N_23154,N_23279);
xor U24474 (N_24474,N_22170,N_22875);
nand U24475 (N_24475,N_23219,N_23410);
nand U24476 (N_24476,N_22522,N_23601);
nand U24477 (N_24477,N_23604,N_22480);
nor U24478 (N_24478,N_23518,N_22923);
or U24479 (N_24479,N_22869,N_22525);
nand U24480 (N_24480,N_23195,N_23178);
and U24481 (N_24481,N_22790,N_22310);
xor U24482 (N_24482,N_22369,N_22062);
xor U24483 (N_24483,N_23345,N_23278);
xnor U24484 (N_24484,N_22748,N_23465);
xor U24485 (N_24485,N_23214,N_22112);
and U24486 (N_24486,N_22147,N_23393);
nand U24487 (N_24487,N_22651,N_22572);
and U24488 (N_24488,N_22392,N_23566);
nor U24489 (N_24489,N_22511,N_22948);
nand U24490 (N_24490,N_22726,N_22625);
or U24491 (N_24491,N_22444,N_23257);
and U24492 (N_24492,N_22032,N_22202);
xor U24493 (N_24493,N_23635,N_22125);
nor U24494 (N_24494,N_23246,N_23334);
xnor U24495 (N_24495,N_23120,N_22549);
or U24496 (N_24496,N_23161,N_23755);
nor U24497 (N_24497,N_23404,N_23286);
or U24498 (N_24498,N_22768,N_23918);
xor U24499 (N_24499,N_23642,N_23493);
nand U24500 (N_24500,N_23534,N_22507);
nand U24501 (N_24501,N_22338,N_23116);
nand U24502 (N_24502,N_22048,N_23007);
or U24503 (N_24503,N_22805,N_23946);
and U24504 (N_24504,N_22028,N_23094);
xor U24505 (N_24505,N_23830,N_22761);
and U24506 (N_24506,N_22825,N_22352);
nor U24507 (N_24507,N_22514,N_23844);
or U24508 (N_24508,N_23262,N_22846);
and U24509 (N_24509,N_22663,N_23380);
nand U24510 (N_24510,N_23386,N_23683);
xnor U24511 (N_24511,N_22779,N_22450);
or U24512 (N_24512,N_23713,N_22602);
and U24513 (N_24513,N_22021,N_23710);
nand U24514 (N_24514,N_22424,N_23540);
and U24515 (N_24515,N_22061,N_22586);
nor U24516 (N_24516,N_23606,N_23681);
xor U24517 (N_24517,N_22225,N_22560);
nor U24518 (N_24518,N_22423,N_23793);
or U24519 (N_24519,N_23517,N_23430);
or U24520 (N_24520,N_22512,N_22195);
nor U24521 (N_24521,N_23688,N_23297);
nor U24522 (N_24522,N_22942,N_23579);
nand U24523 (N_24523,N_22033,N_22637);
nor U24524 (N_24524,N_23064,N_23994);
nand U24525 (N_24525,N_22499,N_22703);
or U24526 (N_24526,N_22696,N_22640);
or U24527 (N_24527,N_23382,N_22744);
and U24528 (N_24528,N_23958,N_22420);
xnor U24529 (N_24529,N_22718,N_22737);
xor U24530 (N_24530,N_22325,N_22177);
nor U24531 (N_24531,N_22359,N_23576);
nand U24532 (N_24532,N_22496,N_22461);
and U24533 (N_24533,N_22693,N_22335);
or U24534 (N_24534,N_22236,N_22216);
or U24535 (N_24535,N_23387,N_22960);
or U24536 (N_24536,N_23878,N_23243);
nand U24537 (N_24537,N_22426,N_22307);
and U24538 (N_24538,N_22690,N_23935);
nand U24539 (N_24539,N_22391,N_22265);
xnor U24540 (N_24540,N_23711,N_22366);
and U24541 (N_24541,N_22706,N_22569);
and U24542 (N_24542,N_23800,N_23242);
or U24543 (N_24543,N_23622,N_23376);
or U24544 (N_24544,N_22515,N_22316);
or U24545 (N_24545,N_23115,N_22561);
xnor U24546 (N_24546,N_22831,N_22834);
xor U24547 (N_24547,N_22133,N_22156);
and U24548 (N_24548,N_22750,N_23982);
nand U24549 (N_24549,N_23818,N_22395);
nor U24550 (N_24550,N_22751,N_22580);
xor U24551 (N_24551,N_23687,N_23886);
and U24552 (N_24552,N_23589,N_23630);
or U24553 (N_24553,N_23165,N_22930);
nor U24554 (N_24554,N_23280,N_22197);
xnor U24555 (N_24555,N_23706,N_22298);
or U24556 (N_24556,N_22357,N_23406);
or U24557 (N_24557,N_23322,N_22946);
or U24558 (N_24558,N_22694,N_23838);
and U24559 (N_24559,N_23789,N_22882);
xnor U24560 (N_24560,N_23984,N_22878);
and U24561 (N_24561,N_22715,N_22477);
nand U24562 (N_24562,N_23427,N_23855);
nand U24563 (N_24563,N_22534,N_22157);
or U24564 (N_24564,N_23896,N_23378);
and U24565 (N_24565,N_22084,N_22428);
and U24566 (N_24566,N_22820,N_22075);
nand U24567 (N_24567,N_23638,N_23015);
and U24568 (N_24568,N_22702,N_23930);
nand U24569 (N_24569,N_22843,N_22329);
xnor U24570 (N_24570,N_22327,N_23905);
xor U24571 (N_24571,N_23936,N_23265);
and U24572 (N_24572,N_23432,N_22859);
xnor U24573 (N_24573,N_23457,N_23198);
nand U24574 (N_24574,N_23888,N_23173);
xor U24575 (N_24575,N_23522,N_22315);
and U24576 (N_24576,N_22536,N_23959);
or U24577 (N_24577,N_22749,N_22810);
nor U24578 (N_24578,N_22849,N_23598);
nand U24579 (N_24579,N_23953,N_22083);
nor U24580 (N_24580,N_23140,N_22180);
and U24581 (N_24581,N_22951,N_23564);
and U24582 (N_24582,N_23446,N_23484);
xor U24583 (N_24583,N_22519,N_22330);
and U24584 (N_24584,N_22608,N_23805);
xnor U24585 (N_24585,N_22431,N_23357);
nand U24586 (N_24586,N_22266,N_22966);
xnor U24587 (N_24587,N_22002,N_22427);
nor U24588 (N_24588,N_23865,N_23673);
nor U24589 (N_24589,N_23551,N_23241);
nand U24590 (N_24590,N_23530,N_23807);
nor U24591 (N_24591,N_22222,N_22013);
and U24592 (N_24592,N_22989,N_22517);
or U24593 (N_24593,N_22175,N_23156);
nand U24594 (N_24594,N_22639,N_23288);
xor U24595 (N_24595,N_23118,N_23020);
nand U24596 (N_24596,N_22023,N_23467);
nand U24597 (N_24597,N_23899,N_23003);
xor U24598 (N_24598,N_23464,N_22440);
nand U24599 (N_24599,N_23741,N_23433);
and U24600 (N_24600,N_22143,N_23304);
nand U24601 (N_24601,N_23614,N_22635);
and U24602 (N_24602,N_23503,N_22613);
and U24603 (N_24603,N_22695,N_22198);
nand U24604 (N_24604,N_23084,N_22998);
or U24605 (N_24605,N_23267,N_22955);
and U24606 (N_24606,N_22072,N_22772);
and U24607 (N_24607,N_23052,N_22035);
xnor U24608 (N_24608,N_23236,N_22802);
or U24609 (N_24609,N_23972,N_22168);
xnor U24610 (N_24610,N_23307,N_23283);
xnor U24611 (N_24611,N_22081,N_23251);
or U24612 (N_24612,N_22079,N_23660);
or U24613 (N_24613,N_22707,N_22908);
nor U24614 (N_24614,N_23593,N_23440);
nor U24615 (N_24615,N_23418,N_23889);
or U24616 (N_24616,N_22816,N_23823);
or U24617 (N_24617,N_23324,N_22506);
or U24618 (N_24618,N_22926,N_22495);
xor U24619 (N_24619,N_22271,N_23196);
and U24620 (N_24620,N_23087,N_22070);
nor U24621 (N_24621,N_23845,N_22259);
or U24622 (N_24622,N_22362,N_22666);
or U24623 (N_24623,N_22643,N_23526);
or U24624 (N_24624,N_23100,N_23328);
or U24625 (N_24625,N_22824,N_22892);
xor U24626 (N_24626,N_22819,N_23843);
nor U24627 (N_24627,N_23558,N_22673);
or U24628 (N_24628,N_23545,N_23586);
nor U24629 (N_24629,N_23069,N_23717);
and U24630 (N_24630,N_23491,N_22193);
and U24631 (N_24631,N_22350,N_22567);
nor U24632 (N_24632,N_23344,N_23931);
and U24633 (N_24633,N_22471,N_23021);
and U24634 (N_24634,N_23734,N_23506);
nor U24635 (N_24635,N_22871,N_23690);
nand U24636 (N_24636,N_22399,N_22556);
and U24637 (N_24637,N_22868,N_22370);
and U24638 (N_24638,N_22432,N_23719);
or U24639 (N_24639,N_23113,N_23648);
nand U24640 (N_24640,N_23697,N_23528);
nor U24641 (N_24641,N_23290,N_22530);
nor U24642 (N_24642,N_22108,N_22785);
or U24643 (N_24643,N_23034,N_23760);
nor U24644 (N_24644,N_23693,N_22442);
xor U24645 (N_24645,N_22145,N_22578);
nand U24646 (N_24646,N_22665,N_22590);
or U24647 (N_24647,N_23152,N_22797);
nand U24648 (N_24648,N_23361,N_22464);
or U24649 (N_24649,N_22701,N_23150);
xor U24650 (N_24650,N_23555,N_22939);
and U24651 (N_24651,N_22003,N_22922);
or U24652 (N_24652,N_23299,N_22174);
or U24653 (N_24653,N_22110,N_22934);
and U24654 (N_24654,N_22091,N_22302);
xnor U24655 (N_24655,N_22886,N_22593);
xor U24656 (N_24656,N_23549,N_23541);
nand U24657 (N_24657,N_23587,N_23403);
nand U24658 (N_24658,N_22166,N_22358);
or U24659 (N_24659,N_22912,N_22559);
and U24660 (N_24660,N_23653,N_22473);
nor U24661 (N_24661,N_22361,N_22343);
xnor U24662 (N_24662,N_22771,N_22038);
and U24663 (N_24663,N_23646,N_23372);
or U24664 (N_24664,N_22538,N_23919);
and U24665 (N_24665,N_23812,N_22503);
or U24666 (N_24666,N_23321,N_23960);
and U24667 (N_24667,N_23709,N_23868);
nor U24668 (N_24668,N_22290,N_23497);
nand U24669 (N_24669,N_23308,N_22189);
or U24670 (N_24670,N_22997,N_22452);
or U24671 (N_24671,N_22889,N_22723);
xnor U24672 (N_24672,N_23368,N_23546);
or U24673 (N_24673,N_22172,N_22382);
nor U24674 (N_24674,N_22592,N_22380);
or U24675 (N_24675,N_22022,N_23781);
nand U24676 (N_24676,N_22129,N_23412);
and U24677 (N_24677,N_23422,N_22106);
nor U24678 (N_24678,N_22141,N_23676);
and U24679 (N_24679,N_23895,N_23532);
and U24680 (N_24680,N_23476,N_22071);
nand U24681 (N_24681,N_23835,N_23402);
and U24682 (N_24682,N_22806,N_23035);
nand U24683 (N_24683,N_23912,N_23200);
and U24684 (N_24684,N_23397,N_22915);
and U24685 (N_24685,N_23186,N_23759);
xnor U24686 (N_24686,N_23249,N_22179);
nand U24687 (N_24687,N_22551,N_23002);
nor U24688 (N_24688,N_22434,N_23819);
and U24689 (N_24689,N_22223,N_22682);
or U24690 (N_24690,N_22766,N_23654);
nor U24691 (N_24691,N_23284,N_23392);
and U24692 (N_24692,N_23603,N_22113);
nand U24693 (N_24693,N_22280,N_22231);
and U24694 (N_24694,N_22117,N_23858);
xor U24695 (N_24695,N_22131,N_22526);
and U24696 (N_24696,N_22454,N_23689);
xnor U24697 (N_24697,N_23712,N_22466);
nor U24698 (N_24698,N_23092,N_23008);
nand U24699 (N_24699,N_22931,N_22049);
xor U24700 (N_24700,N_23831,N_23256);
or U24701 (N_24701,N_22733,N_22605);
nor U24702 (N_24702,N_22341,N_22896);
nor U24703 (N_24703,N_22652,N_23929);
nor U24704 (N_24704,N_22533,N_23032);
xor U24705 (N_24705,N_23911,N_22603);
xnor U24706 (N_24706,N_23193,N_22568);
nor U24707 (N_24707,N_22139,N_23151);
xor U24708 (N_24708,N_22832,N_22759);
or U24709 (N_24709,N_23138,N_23483);
nor U24710 (N_24710,N_23201,N_22776);
nand U24711 (N_24711,N_22853,N_22043);
nand U24712 (N_24712,N_22076,N_22727);
nand U24713 (N_24713,N_23993,N_22196);
nand U24714 (N_24714,N_23804,N_22717);
nand U24715 (N_24715,N_23933,N_23679);
nand U24716 (N_24716,N_22176,N_22932);
xnor U24717 (N_24717,N_23543,N_23902);
nand U24718 (N_24718,N_22493,N_23018);
and U24719 (N_24719,N_22901,N_23725);
xnor U24720 (N_24720,N_23226,N_23791);
xor U24721 (N_24721,N_22211,N_22159);
and U24722 (N_24722,N_23314,N_23990);
and U24723 (N_24723,N_22581,N_22763);
and U24724 (N_24724,N_23350,N_22623);
nand U24725 (N_24725,N_22262,N_22169);
xnor U24726 (N_24726,N_23162,N_22219);
nand U24727 (N_24727,N_23316,N_23106);
xnor U24728 (N_24728,N_22479,N_23939);
and U24729 (N_24729,N_23514,N_23950);
nor U24730 (N_24730,N_23640,N_22809);
nand U24731 (N_24731,N_23091,N_22199);
nor U24732 (N_24732,N_23723,N_23353);
nor U24733 (N_24733,N_22067,N_22400);
and U24734 (N_24734,N_23827,N_22230);
or U24735 (N_24735,N_23247,N_22687);
or U24736 (N_24736,N_23535,N_23029);
nor U24737 (N_24737,N_22742,N_23539);
or U24738 (N_24738,N_22489,N_23244);
nor U24739 (N_24739,N_23634,N_23567);
xnor U24740 (N_24740,N_23932,N_22760);
nor U24741 (N_24741,N_23231,N_23944);
xnor U24742 (N_24742,N_22598,N_23434);
nor U24743 (N_24743,N_23168,N_22542);
nand U24744 (N_24744,N_23301,N_23093);
or U24745 (N_24745,N_22800,N_23924);
nor U24746 (N_24746,N_22903,N_22214);
nand U24747 (N_24747,N_23573,N_23921);
or U24748 (N_24748,N_23874,N_22124);
and U24749 (N_24749,N_23312,N_22348);
nor U24750 (N_24750,N_22408,N_22127);
or U24751 (N_24751,N_22443,N_22066);
xnor U24752 (N_24752,N_22275,N_23426);
nand U24753 (N_24753,N_22699,N_22502);
and U24754 (N_24754,N_23785,N_22840);
nor U24755 (N_24755,N_22941,N_23317);
and U24756 (N_24756,N_23794,N_22165);
or U24757 (N_24757,N_23323,N_23326);
nand U24758 (N_24758,N_22118,N_23480);
nor U24759 (N_24759,N_23965,N_22531);
nand U24760 (N_24760,N_23472,N_22425);
xnor U24761 (N_24761,N_23318,N_23643);
or U24762 (N_24762,N_23217,N_23238);
and U24763 (N_24763,N_22178,N_23652);
xnor U24764 (N_24764,N_23394,N_22398);
nand U24765 (N_24765,N_23208,N_23520);
or U24766 (N_24766,N_22011,N_23157);
nor U24767 (N_24767,N_22111,N_23824);
and U24768 (N_24768,N_23674,N_22539);
and U24769 (N_24769,N_23866,N_22722);
and U24770 (N_24770,N_22397,N_22205);
xor U24771 (N_24771,N_23221,N_22584);
nand U24772 (N_24772,N_23595,N_22636);
nor U24773 (N_24773,N_23347,N_22251);
or U24774 (N_24774,N_23142,N_23732);
nand U24775 (N_24775,N_23363,N_23261);
nor U24776 (N_24776,N_22547,N_22082);
xor U24777 (N_24777,N_23671,N_22993);
and U24778 (N_24778,N_23947,N_22731);
or U24779 (N_24779,N_23325,N_22401);
nand U24780 (N_24780,N_23104,N_22226);
or U24781 (N_24781,N_23492,N_22664);
and U24782 (N_24782,N_23045,N_22950);
nor U24783 (N_24783,N_23668,N_23149);
nand U24784 (N_24784,N_22782,N_23803);
and U24785 (N_24785,N_23128,N_22374);
or U24786 (N_24786,N_22482,N_23979);
nand U24787 (N_24787,N_22201,N_23292);
nand U24788 (N_24788,N_23381,N_23067);
and U24789 (N_24789,N_22405,N_23963);
and U24790 (N_24790,N_22630,N_22801);
xor U24791 (N_24791,N_23395,N_22385);
and U24792 (N_24792,N_22001,N_23225);
nor U24793 (N_24793,N_23559,N_22906);
or U24794 (N_24794,N_23205,N_23867);
xnor U24795 (N_24795,N_22413,N_22881);
xnor U24796 (N_24796,N_23349,N_22204);
nor U24797 (N_24797,N_22376,N_23129);
nor U24798 (N_24798,N_22705,N_23276);
nor U24799 (N_24799,N_22487,N_23466);
and U24800 (N_24800,N_22009,N_22684);
xor U24801 (N_24801,N_22318,N_23708);
or U24802 (N_24802,N_22880,N_23684);
and U24803 (N_24803,N_22971,N_23107);
nor U24804 (N_24804,N_22807,N_22294);
nand U24805 (N_24805,N_22736,N_22324);
and U24806 (N_24806,N_22279,N_23204);
xnor U24807 (N_24807,N_23701,N_22364);
nand U24808 (N_24808,N_22073,N_23013);
and U24809 (N_24809,N_23255,N_23220);
nor U24810 (N_24810,N_22351,N_22990);
nor U24811 (N_24811,N_23581,N_22077);
xnor U24812 (N_24812,N_22270,N_23928);
and U24813 (N_24813,N_23746,N_22612);
and U24814 (N_24814,N_22253,N_22631);
and U24815 (N_24815,N_23730,N_22239);
and U24816 (N_24816,N_22570,N_22550);
nand U24817 (N_24817,N_23125,N_23856);
and U24818 (N_24818,N_23859,N_22135);
xnor U24819 (N_24819,N_23082,N_22857);
xnor U24820 (N_24820,N_22959,N_23436);
nor U24821 (N_24821,N_22537,N_23185);
xor U24822 (N_24822,N_23599,N_22261);
and U24823 (N_24823,N_23031,N_23079);
nor U24824 (N_24824,N_23194,N_22686);
nand U24825 (N_24825,N_22206,N_23998);
xor U24826 (N_24826,N_23442,N_22504);
nor U24827 (N_24827,N_23153,N_22983);
nand U24828 (N_24828,N_22783,N_22356);
and U24829 (N_24829,N_22979,N_22163);
nand U24830 (N_24830,N_23266,N_22898);
nand U24831 (N_24831,N_22116,N_22378);
xor U24832 (N_24832,N_23099,N_23268);
nand U24833 (N_24833,N_23773,N_22063);
nor U24834 (N_24834,N_23873,N_23248);
nor U24835 (N_24835,N_23795,N_23435);
nor U24836 (N_24836,N_22518,N_23504);
nor U24837 (N_24837,N_23191,N_22792);
or U24838 (N_24838,N_23798,N_23070);
xnor U24839 (N_24839,N_23281,N_22277);
and U24840 (N_24840,N_22936,N_23966);
xnor U24841 (N_24841,N_23951,N_22304);
nand U24842 (N_24842,N_23981,N_22938);
or U24843 (N_24843,N_23847,N_22268);
or U24844 (N_24844,N_22240,N_22758);
nor U24845 (N_24845,N_23250,N_23937);
or U24846 (N_24846,N_23017,N_23415);
nor U24847 (N_24847,N_23801,N_23459);
xor U24848 (N_24848,N_22250,N_22472);
or U24849 (N_24849,N_23846,N_22917);
and U24850 (N_24850,N_23411,N_23147);
nand U24851 (N_24851,N_22811,N_22969);
nand U24852 (N_24852,N_23841,N_22234);
or U24853 (N_24853,N_23872,N_23098);
xnor U24854 (N_24854,N_23637,N_23897);
xor U24855 (N_24855,N_22796,N_23842);
nor U24856 (N_24856,N_22861,N_23647);
nand U24857 (N_24857,N_22221,N_23014);
nand U24858 (N_24858,N_22347,N_22254);
nand U24859 (N_24859,N_23211,N_22957);
nand U24860 (N_24860,N_22014,N_23778);
nor U24861 (N_24861,N_22345,N_22349);
and U24862 (N_24862,N_22720,N_23180);
nor U24863 (N_24863,N_23777,N_23910);
and U24864 (N_24864,N_22041,N_23607);
nand U24865 (N_24865,N_22301,N_23940);
xor U24866 (N_24866,N_22847,N_22437);
nor U24867 (N_24867,N_23183,N_23916);
or U24868 (N_24868,N_22845,N_22485);
xor U24869 (N_24869,N_23254,N_22729);
and U24870 (N_24870,N_23605,N_23796);
or U24871 (N_24871,N_23699,N_22883);
or U24872 (N_24872,N_22390,N_22456);
nor U24873 (N_24873,N_23600,N_22232);
or U24874 (N_24874,N_22255,N_23109);
xnor U24875 (N_24875,N_22611,N_22540);
and U24876 (N_24876,N_22006,N_22367);
xor U24877 (N_24877,N_22870,N_22103);
nand U24878 (N_24878,N_22429,N_22158);
nor U24879 (N_24879,N_23362,N_22164);
xor U24880 (N_24880,N_22844,N_22449);
nor U24881 (N_24881,N_22384,N_22884);
or U24882 (N_24882,N_22069,N_22097);
nor U24883 (N_24883,N_22241,N_23233);
or U24884 (N_24884,N_23617,N_22016);
nand U24885 (N_24885,N_23726,N_23641);
nor U24886 (N_24886,N_22658,N_22913);
and U24887 (N_24887,N_23028,N_22975);
nand U24888 (N_24888,N_22249,N_23498);
nand U24889 (N_24889,N_23934,N_23786);
nor U24890 (N_24890,N_23584,N_23143);
and U24891 (N_24891,N_23202,N_23615);
xnor U24892 (N_24892,N_23228,N_22662);
nor U24893 (N_24893,N_23366,N_23563);
and U24894 (N_24894,N_22162,N_23352);
or U24895 (N_24895,N_22585,N_23371);
nand U24896 (N_24896,N_23309,N_23696);
nand U24897 (N_24897,N_23355,N_22553);
nand U24898 (N_24898,N_23447,N_22848);
xor U24899 (N_24899,N_22872,N_23127);
or U24900 (N_24900,N_22588,N_23970);
or U24901 (N_24901,N_23811,N_23724);
and U24902 (N_24902,N_23728,N_22060);
xnor U24903 (N_24903,N_22527,N_23627);
nand U24904 (N_24904,N_22293,N_22475);
xor U24905 (N_24905,N_22130,N_23148);
xor U24906 (N_24906,N_23508,N_22029);
xnor U24907 (N_24907,N_23495,N_22937);
and U24908 (N_24908,N_23041,N_23774);
or U24909 (N_24909,N_22299,N_22505);
xnor U24910 (N_24910,N_23964,N_22873);
xor U24911 (N_24911,N_23533,N_23058);
nand U24912 (N_24912,N_23141,N_23612);
nand U24913 (N_24913,N_22501,N_23569);
xor U24914 (N_24914,N_23716,N_23685);
nand U24915 (N_24915,N_22725,N_23176);
nand U24916 (N_24916,N_23808,N_23561);
xnor U24917 (N_24917,N_23809,N_23485);
xnor U24918 (N_24918,N_23949,N_22192);
nand U24919 (N_24919,N_23513,N_22678);
xnor U24920 (N_24920,N_23170,N_23478);
or U24921 (N_24921,N_23861,N_23509);
nand U24922 (N_24922,N_23470,N_23749);
or U24923 (N_24923,N_22492,N_23507);
xnor U24924 (N_24924,N_22929,N_22187);
nand U24925 (N_24925,N_23834,N_22167);
xnor U24926 (N_24926,N_22661,N_22677);
and U24927 (N_24927,N_22257,N_23766);
nor U24928 (N_24928,N_22996,N_22269);
nand U24929 (N_24929,N_22321,N_23062);
nor U24930 (N_24930,N_23136,N_23714);
nand U24931 (N_24931,N_22155,N_22059);
and U24932 (N_24932,N_23552,N_22094);
nand U24933 (N_24933,N_23597,N_23155);
xor U24934 (N_24934,N_23199,N_23780);
nand U24935 (N_24935,N_23736,N_22470);
nand U24936 (N_24936,N_22713,N_23072);
and U24937 (N_24937,N_22716,N_23046);
nor U24938 (N_24938,N_22854,N_22803);
and U24939 (N_24939,N_23769,N_22791);
xnor U24940 (N_24940,N_22564,N_22554);
nor U24941 (N_24941,N_23527,N_23389);
nor U24942 (N_24942,N_22411,N_22465);
or U24943 (N_24943,N_23421,N_22818);
and U24944 (N_24944,N_23218,N_23639);
nor U24945 (N_24945,N_23313,N_22924);
and U24946 (N_24946,N_23623,N_22252);
or U24947 (N_24947,N_23385,N_23926);
xnor U24948 (N_24948,N_23772,N_23016);
nor U24949 (N_24949,N_23763,N_23333);
nand U24950 (N_24950,N_22877,N_23081);
and U24951 (N_24951,N_23496,N_23494);
nand U24952 (N_24952,N_22246,N_23271);
and U24953 (N_24953,N_22563,N_23892);
or U24954 (N_24954,N_23853,N_22754);
or U24955 (N_24955,N_22404,N_22980);
xor U24956 (N_24956,N_22583,N_22740);
and U24957 (N_24957,N_23047,N_22331);
or U24958 (N_24958,N_23629,N_23718);
or U24959 (N_24959,N_22476,N_23230);
and U24960 (N_24960,N_23287,N_22154);
xnor U24961 (N_24961,N_23117,N_22952);
nor U24962 (N_24962,N_22953,N_23163);
or U24963 (N_24963,N_23837,N_23332);
xor U24964 (N_24964,N_23111,N_23164);
or U24965 (N_24965,N_23005,N_23762);
xnor U24966 (N_24966,N_23258,N_22486);
or U24967 (N_24967,N_22510,N_23405);
or U24968 (N_24968,N_22322,N_22297);
xor U24969 (N_24969,N_22724,N_23282);
nand U24970 (N_24970,N_22822,N_23197);
nor U24971 (N_24971,N_22659,N_23538);
xnor U24972 (N_24972,N_23420,N_23978);
nand U24973 (N_24973,N_23119,N_23078);
or U24974 (N_24974,N_22284,N_22655);
nand U24975 (N_24975,N_22962,N_22336);
and U24976 (N_24976,N_23575,N_23245);
and U24977 (N_24977,N_23703,N_23097);
xnor U24978 (N_24978,N_23826,N_23131);
xnor U24979 (N_24979,N_22893,N_23987);
and U24980 (N_24980,N_22099,N_23025);
nor U24981 (N_24981,N_22627,N_23661);
and U24982 (N_24982,N_23745,N_23137);
and U24983 (N_24983,N_23499,N_22283);
or U24984 (N_24984,N_22855,N_22688);
nor U24985 (N_24985,N_23055,N_22308);
or U24986 (N_24986,N_23294,N_22513);
and U24987 (N_24987,N_22457,N_22858);
nand U24988 (N_24988,N_23399,N_22764);
and U24989 (N_24989,N_22654,N_23374);
xnor U24990 (N_24990,N_22453,N_23908);
and U24991 (N_24991,N_23095,N_22228);
or U24992 (N_24992,N_23715,N_23974);
or U24993 (N_24993,N_23675,N_23952);
nor U24994 (N_24994,N_23920,N_23656);
and U24995 (N_24995,N_22866,N_23871);
nor U24996 (N_24996,N_23529,N_22332);
xnor U24997 (N_24997,N_22149,N_22074);
xnor U24998 (N_24998,N_22100,N_23894);
nand U24999 (N_24999,N_23659,N_23863);
nor U25000 (N_25000,N_22785,N_22271);
xnor U25001 (N_25001,N_23170,N_23847);
or U25002 (N_25002,N_22692,N_22569);
and U25003 (N_25003,N_22949,N_22429);
and U25004 (N_25004,N_22013,N_23731);
or U25005 (N_25005,N_22161,N_23651);
and U25006 (N_25006,N_22785,N_23456);
nand U25007 (N_25007,N_22074,N_23632);
and U25008 (N_25008,N_23344,N_23394);
nor U25009 (N_25009,N_23635,N_23934);
and U25010 (N_25010,N_23508,N_22055);
nor U25011 (N_25011,N_22812,N_22214);
xnor U25012 (N_25012,N_22677,N_22864);
nand U25013 (N_25013,N_22527,N_22975);
nor U25014 (N_25014,N_22049,N_23709);
nor U25015 (N_25015,N_23521,N_22641);
nor U25016 (N_25016,N_23609,N_23473);
nand U25017 (N_25017,N_22424,N_23655);
nor U25018 (N_25018,N_22191,N_23325);
or U25019 (N_25019,N_23680,N_22074);
or U25020 (N_25020,N_23858,N_22724);
and U25021 (N_25021,N_22104,N_23318);
nand U25022 (N_25022,N_23074,N_22324);
xnor U25023 (N_25023,N_23805,N_22105);
or U25024 (N_25024,N_22241,N_23213);
or U25025 (N_25025,N_23717,N_22399);
or U25026 (N_25026,N_23087,N_23950);
and U25027 (N_25027,N_22915,N_23388);
or U25028 (N_25028,N_22480,N_22042);
nand U25029 (N_25029,N_22856,N_22154);
nand U25030 (N_25030,N_22284,N_22197);
nand U25031 (N_25031,N_22053,N_22291);
nand U25032 (N_25032,N_22857,N_22346);
and U25033 (N_25033,N_22382,N_23944);
nand U25034 (N_25034,N_23944,N_23450);
or U25035 (N_25035,N_22965,N_22925);
nor U25036 (N_25036,N_22092,N_23107);
xnor U25037 (N_25037,N_23007,N_22881);
nor U25038 (N_25038,N_22507,N_23014);
nand U25039 (N_25039,N_23753,N_23675);
xnor U25040 (N_25040,N_23514,N_22805);
or U25041 (N_25041,N_23593,N_23918);
and U25042 (N_25042,N_22009,N_23727);
or U25043 (N_25043,N_22280,N_22176);
nand U25044 (N_25044,N_22775,N_22903);
nand U25045 (N_25045,N_22907,N_22327);
or U25046 (N_25046,N_23290,N_23149);
and U25047 (N_25047,N_23548,N_22737);
or U25048 (N_25048,N_23701,N_22823);
nand U25049 (N_25049,N_23791,N_23889);
and U25050 (N_25050,N_23661,N_23784);
xor U25051 (N_25051,N_23069,N_22470);
nor U25052 (N_25052,N_22369,N_22100);
or U25053 (N_25053,N_22588,N_22390);
nor U25054 (N_25054,N_22438,N_22706);
xnor U25055 (N_25055,N_23417,N_23642);
and U25056 (N_25056,N_23583,N_22163);
and U25057 (N_25057,N_23368,N_23427);
nor U25058 (N_25058,N_22628,N_23000);
nand U25059 (N_25059,N_23336,N_22435);
nand U25060 (N_25060,N_23292,N_23111);
nand U25061 (N_25061,N_23043,N_22526);
nor U25062 (N_25062,N_22317,N_23066);
xor U25063 (N_25063,N_22608,N_22916);
xnor U25064 (N_25064,N_22733,N_23689);
and U25065 (N_25065,N_23927,N_22013);
xor U25066 (N_25066,N_22604,N_22905);
or U25067 (N_25067,N_22455,N_23239);
nand U25068 (N_25068,N_23166,N_22091);
nor U25069 (N_25069,N_22545,N_23185);
nand U25070 (N_25070,N_22483,N_23362);
nor U25071 (N_25071,N_22918,N_23487);
nor U25072 (N_25072,N_23572,N_23683);
or U25073 (N_25073,N_23305,N_23912);
and U25074 (N_25074,N_22917,N_22116);
nand U25075 (N_25075,N_23845,N_22015);
or U25076 (N_25076,N_22667,N_23244);
nor U25077 (N_25077,N_23304,N_23726);
or U25078 (N_25078,N_23001,N_22336);
and U25079 (N_25079,N_23257,N_23038);
and U25080 (N_25080,N_23878,N_22745);
and U25081 (N_25081,N_23447,N_22093);
nor U25082 (N_25082,N_23289,N_23327);
nor U25083 (N_25083,N_23571,N_23924);
xnor U25084 (N_25084,N_22470,N_23173);
nor U25085 (N_25085,N_23189,N_23879);
or U25086 (N_25086,N_22714,N_23030);
xnor U25087 (N_25087,N_23778,N_23107);
nand U25088 (N_25088,N_23848,N_22626);
nor U25089 (N_25089,N_23460,N_22592);
and U25090 (N_25090,N_22221,N_22316);
nand U25091 (N_25091,N_23479,N_22208);
and U25092 (N_25092,N_23703,N_23387);
or U25093 (N_25093,N_22737,N_22910);
or U25094 (N_25094,N_22096,N_23844);
nand U25095 (N_25095,N_22617,N_22656);
nor U25096 (N_25096,N_23666,N_22223);
nor U25097 (N_25097,N_23303,N_23137);
or U25098 (N_25098,N_22898,N_22154);
nor U25099 (N_25099,N_23192,N_23151);
and U25100 (N_25100,N_22695,N_22072);
nand U25101 (N_25101,N_22130,N_22100);
xor U25102 (N_25102,N_23862,N_22021);
nor U25103 (N_25103,N_22979,N_23530);
xor U25104 (N_25104,N_23779,N_22995);
nand U25105 (N_25105,N_22286,N_22802);
nand U25106 (N_25106,N_22802,N_22190);
and U25107 (N_25107,N_22635,N_23861);
nand U25108 (N_25108,N_23610,N_22481);
or U25109 (N_25109,N_22611,N_23055);
or U25110 (N_25110,N_22769,N_23745);
xnor U25111 (N_25111,N_22252,N_22237);
or U25112 (N_25112,N_23521,N_22264);
xnor U25113 (N_25113,N_22994,N_22858);
and U25114 (N_25114,N_22173,N_22791);
nor U25115 (N_25115,N_22609,N_22010);
nor U25116 (N_25116,N_23808,N_23100);
xnor U25117 (N_25117,N_22252,N_22719);
xor U25118 (N_25118,N_22154,N_23011);
and U25119 (N_25119,N_22897,N_23668);
nor U25120 (N_25120,N_23841,N_23826);
or U25121 (N_25121,N_22421,N_22625);
nand U25122 (N_25122,N_22408,N_23548);
nand U25123 (N_25123,N_23707,N_22643);
or U25124 (N_25124,N_23692,N_22442);
and U25125 (N_25125,N_22836,N_23054);
nand U25126 (N_25126,N_22693,N_23407);
xnor U25127 (N_25127,N_22559,N_22592);
or U25128 (N_25128,N_22502,N_22822);
and U25129 (N_25129,N_22912,N_23565);
xnor U25130 (N_25130,N_23950,N_23612);
nand U25131 (N_25131,N_23902,N_22653);
nand U25132 (N_25132,N_23250,N_22518);
nor U25133 (N_25133,N_23366,N_23983);
and U25134 (N_25134,N_22159,N_22219);
or U25135 (N_25135,N_23479,N_23924);
or U25136 (N_25136,N_23476,N_22229);
and U25137 (N_25137,N_22068,N_23004);
nor U25138 (N_25138,N_22184,N_23373);
nor U25139 (N_25139,N_22668,N_22147);
nand U25140 (N_25140,N_22958,N_23071);
xor U25141 (N_25141,N_23970,N_23343);
nand U25142 (N_25142,N_23389,N_22366);
or U25143 (N_25143,N_23349,N_23231);
nand U25144 (N_25144,N_22586,N_22318);
and U25145 (N_25145,N_23530,N_22245);
and U25146 (N_25146,N_22673,N_22558);
or U25147 (N_25147,N_23762,N_22287);
nand U25148 (N_25148,N_23939,N_22754);
nor U25149 (N_25149,N_23443,N_22697);
xnor U25150 (N_25150,N_23851,N_23175);
nor U25151 (N_25151,N_22907,N_23361);
xnor U25152 (N_25152,N_23919,N_23316);
and U25153 (N_25153,N_23939,N_23199);
and U25154 (N_25154,N_22674,N_23984);
nand U25155 (N_25155,N_23740,N_22903);
and U25156 (N_25156,N_23059,N_22599);
xor U25157 (N_25157,N_22380,N_23145);
xor U25158 (N_25158,N_23509,N_23625);
nor U25159 (N_25159,N_23706,N_22409);
nor U25160 (N_25160,N_23065,N_22007);
or U25161 (N_25161,N_23520,N_22771);
nor U25162 (N_25162,N_23587,N_23827);
nand U25163 (N_25163,N_22725,N_22756);
and U25164 (N_25164,N_23622,N_23492);
xor U25165 (N_25165,N_23953,N_22237);
nand U25166 (N_25166,N_22777,N_22886);
and U25167 (N_25167,N_22778,N_22297);
nor U25168 (N_25168,N_23784,N_23602);
and U25169 (N_25169,N_22384,N_22057);
and U25170 (N_25170,N_23775,N_23141);
xnor U25171 (N_25171,N_23873,N_23787);
nor U25172 (N_25172,N_22417,N_22481);
nor U25173 (N_25173,N_23860,N_22079);
and U25174 (N_25174,N_22871,N_23426);
or U25175 (N_25175,N_22019,N_22174);
nor U25176 (N_25176,N_22838,N_23629);
nor U25177 (N_25177,N_22962,N_22900);
nor U25178 (N_25178,N_23184,N_22528);
nor U25179 (N_25179,N_22909,N_23646);
nand U25180 (N_25180,N_23475,N_22424);
xnor U25181 (N_25181,N_22105,N_23450);
and U25182 (N_25182,N_23557,N_22557);
xnor U25183 (N_25183,N_23684,N_22889);
or U25184 (N_25184,N_22007,N_23686);
or U25185 (N_25185,N_23530,N_22739);
or U25186 (N_25186,N_23974,N_22500);
nand U25187 (N_25187,N_22944,N_23997);
nor U25188 (N_25188,N_23514,N_22771);
or U25189 (N_25189,N_22010,N_23415);
and U25190 (N_25190,N_22869,N_22006);
nand U25191 (N_25191,N_22012,N_22066);
nand U25192 (N_25192,N_22489,N_22778);
nor U25193 (N_25193,N_22203,N_22922);
xor U25194 (N_25194,N_22740,N_23425);
or U25195 (N_25195,N_23495,N_23958);
xnor U25196 (N_25196,N_22376,N_22814);
and U25197 (N_25197,N_23179,N_23565);
xnor U25198 (N_25198,N_23966,N_22352);
and U25199 (N_25199,N_23627,N_23830);
xor U25200 (N_25200,N_23002,N_22287);
xnor U25201 (N_25201,N_23584,N_22601);
and U25202 (N_25202,N_22243,N_23104);
nor U25203 (N_25203,N_22595,N_23650);
xor U25204 (N_25204,N_22802,N_22472);
xor U25205 (N_25205,N_23407,N_23672);
xnor U25206 (N_25206,N_22221,N_22120);
nand U25207 (N_25207,N_23037,N_22763);
and U25208 (N_25208,N_23541,N_22560);
nor U25209 (N_25209,N_23728,N_22422);
xor U25210 (N_25210,N_22657,N_23159);
xnor U25211 (N_25211,N_22037,N_22682);
nand U25212 (N_25212,N_23614,N_22523);
nand U25213 (N_25213,N_22029,N_23063);
nand U25214 (N_25214,N_22798,N_22146);
and U25215 (N_25215,N_23593,N_23125);
nand U25216 (N_25216,N_23812,N_23249);
nand U25217 (N_25217,N_23842,N_23082);
and U25218 (N_25218,N_22944,N_23753);
nor U25219 (N_25219,N_23275,N_23625);
or U25220 (N_25220,N_23350,N_23879);
and U25221 (N_25221,N_23781,N_23901);
or U25222 (N_25222,N_22438,N_22354);
nor U25223 (N_25223,N_23206,N_23746);
nor U25224 (N_25224,N_23397,N_23915);
and U25225 (N_25225,N_22023,N_23045);
and U25226 (N_25226,N_22382,N_23025);
or U25227 (N_25227,N_22702,N_23762);
nand U25228 (N_25228,N_22563,N_23952);
nor U25229 (N_25229,N_23248,N_22244);
or U25230 (N_25230,N_22639,N_23850);
nand U25231 (N_25231,N_22178,N_22769);
xor U25232 (N_25232,N_23057,N_22249);
or U25233 (N_25233,N_23772,N_23761);
nor U25234 (N_25234,N_22632,N_23281);
and U25235 (N_25235,N_23254,N_22517);
nor U25236 (N_25236,N_23193,N_23508);
xnor U25237 (N_25237,N_23504,N_23797);
nand U25238 (N_25238,N_22117,N_23502);
nor U25239 (N_25239,N_23827,N_22302);
or U25240 (N_25240,N_22653,N_22709);
or U25241 (N_25241,N_23827,N_23220);
or U25242 (N_25242,N_23835,N_23227);
nand U25243 (N_25243,N_23587,N_22967);
or U25244 (N_25244,N_23879,N_23008);
nand U25245 (N_25245,N_23773,N_23426);
xnor U25246 (N_25246,N_22627,N_22536);
xor U25247 (N_25247,N_22763,N_22688);
nand U25248 (N_25248,N_23240,N_23682);
xnor U25249 (N_25249,N_22856,N_23622);
xnor U25250 (N_25250,N_22346,N_23159);
xnor U25251 (N_25251,N_22415,N_23995);
nor U25252 (N_25252,N_22737,N_22027);
nor U25253 (N_25253,N_22519,N_22308);
xor U25254 (N_25254,N_23726,N_23419);
or U25255 (N_25255,N_23503,N_23074);
nor U25256 (N_25256,N_22420,N_22086);
and U25257 (N_25257,N_23616,N_22983);
or U25258 (N_25258,N_22451,N_22156);
and U25259 (N_25259,N_22867,N_23330);
nor U25260 (N_25260,N_22132,N_23966);
and U25261 (N_25261,N_22637,N_22196);
nand U25262 (N_25262,N_23922,N_22511);
and U25263 (N_25263,N_23196,N_22006);
nor U25264 (N_25264,N_22141,N_23489);
xor U25265 (N_25265,N_22574,N_23502);
or U25266 (N_25266,N_23333,N_22879);
xnor U25267 (N_25267,N_23669,N_22279);
nand U25268 (N_25268,N_23569,N_23426);
nand U25269 (N_25269,N_23681,N_22001);
nor U25270 (N_25270,N_22576,N_22407);
nand U25271 (N_25271,N_22788,N_23832);
or U25272 (N_25272,N_23305,N_23639);
or U25273 (N_25273,N_23147,N_23862);
and U25274 (N_25274,N_23824,N_22958);
nor U25275 (N_25275,N_23827,N_23659);
nor U25276 (N_25276,N_22725,N_22808);
and U25277 (N_25277,N_23918,N_23166);
nor U25278 (N_25278,N_23888,N_22423);
nand U25279 (N_25279,N_23777,N_23218);
xnor U25280 (N_25280,N_22056,N_23058);
and U25281 (N_25281,N_23507,N_23225);
or U25282 (N_25282,N_23181,N_23316);
nor U25283 (N_25283,N_22582,N_22278);
nor U25284 (N_25284,N_23414,N_23738);
or U25285 (N_25285,N_23516,N_22905);
nor U25286 (N_25286,N_23718,N_23617);
nor U25287 (N_25287,N_22906,N_23805);
nor U25288 (N_25288,N_22714,N_23452);
nor U25289 (N_25289,N_23057,N_22885);
or U25290 (N_25290,N_23117,N_22780);
nand U25291 (N_25291,N_22090,N_22849);
nand U25292 (N_25292,N_22603,N_23908);
nand U25293 (N_25293,N_22381,N_23956);
nand U25294 (N_25294,N_23686,N_22167);
nor U25295 (N_25295,N_23553,N_22790);
and U25296 (N_25296,N_22834,N_22505);
or U25297 (N_25297,N_23367,N_23903);
nand U25298 (N_25298,N_22235,N_22823);
nor U25299 (N_25299,N_22339,N_23350);
or U25300 (N_25300,N_22228,N_23034);
nand U25301 (N_25301,N_23866,N_22371);
nand U25302 (N_25302,N_22597,N_23090);
nand U25303 (N_25303,N_22819,N_23209);
nor U25304 (N_25304,N_22834,N_22972);
nor U25305 (N_25305,N_22843,N_23598);
or U25306 (N_25306,N_22310,N_23943);
or U25307 (N_25307,N_23827,N_22192);
nor U25308 (N_25308,N_22428,N_23233);
or U25309 (N_25309,N_22401,N_23232);
nor U25310 (N_25310,N_22360,N_22902);
or U25311 (N_25311,N_22378,N_22162);
xor U25312 (N_25312,N_23498,N_22935);
nand U25313 (N_25313,N_23846,N_22707);
nor U25314 (N_25314,N_23878,N_22447);
and U25315 (N_25315,N_23850,N_22165);
xor U25316 (N_25316,N_22300,N_22394);
nand U25317 (N_25317,N_22353,N_22335);
and U25318 (N_25318,N_22188,N_22043);
nand U25319 (N_25319,N_23259,N_22880);
xor U25320 (N_25320,N_22954,N_22360);
xor U25321 (N_25321,N_23586,N_22188);
nand U25322 (N_25322,N_23275,N_23674);
xnor U25323 (N_25323,N_23713,N_22046);
and U25324 (N_25324,N_23486,N_23868);
and U25325 (N_25325,N_22685,N_22310);
and U25326 (N_25326,N_22473,N_23260);
nor U25327 (N_25327,N_23141,N_23516);
nand U25328 (N_25328,N_23234,N_22032);
nor U25329 (N_25329,N_23950,N_22830);
or U25330 (N_25330,N_22266,N_22954);
or U25331 (N_25331,N_23431,N_23427);
xnor U25332 (N_25332,N_23292,N_23723);
nand U25333 (N_25333,N_23611,N_22939);
nor U25334 (N_25334,N_23831,N_22742);
and U25335 (N_25335,N_22029,N_22365);
xor U25336 (N_25336,N_22443,N_23056);
xnor U25337 (N_25337,N_23702,N_22969);
or U25338 (N_25338,N_23265,N_22442);
xnor U25339 (N_25339,N_23858,N_22239);
or U25340 (N_25340,N_22921,N_23451);
xnor U25341 (N_25341,N_23746,N_22421);
nor U25342 (N_25342,N_23569,N_23032);
nand U25343 (N_25343,N_22884,N_22571);
and U25344 (N_25344,N_23877,N_23688);
xnor U25345 (N_25345,N_22530,N_23121);
or U25346 (N_25346,N_22481,N_23714);
or U25347 (N_25347,N_22159,N_23682);
or U25348 (N_25348,N_22796,N_22759);
and U25349 (N_25349,N_23544,N_22104);
xnor U25350 (N_25350,N_22380,N_23103);
nor U25351 (N_25351,N_22657,N_22493);
nand U25352 (N_25352,N_22482,N_23961);
nor U25353 (N_25353,N_22623,N_22952);
nor U25354 (N_25354,N_23998,N_22110);
nor U25355 (N_25355,N_22708,N_23814);
and U25356 (N_25356,N_22995,N_23252);
nor U25357 (N_25357,N_23649,N_22715);
nor U25358 (N_25358,N_22237,N_23260);
and U25359 (N_25359,N_23866,N_22009);
and U25360 (N_25360,N_22522,N_23900);
and U25361 (N_25361,N_23631,N_22192);
or U25362 (N_25362,N_22535,N_22391);
nand U25363 (N_25363,N_23456,N_23990);
nand U25364 (N_25364,N_23564,N_22728);
or U25365 (N_25365,N_23696,N_22607);
and U25366 (N_25366,N_23680,N_23332);
or U25367 (N_25367,N_22295,N_22940);
xnor U25368 (N_25368,N_23479,N_23635);
xor U25369 (N_25369,N_22560,N_22037);
xnor U25370 (N_25370,N_23238,N_23931);
nor U25371 (N_25371,N_22333,N_23362);
nand U25372 (N_25372,N_22189,N_23855);
xor U25373 (N_25373,N_23535,N_23820);
xor U25374 (N_25374,N_22345,N_22978);
or U25375 (N_25375,N_23604,N_22543);
or U25376 (N_25376,N_23502,N_22682);
and U25377 (N_25377,N_22440,N_22146);
nor U25378 (N_25378,N_22217,N_23738);
nand U25379 (N_25379,N_23145,N_23192);
or U25380 (N_25380,N_22116,N_22265);
or U25381 (N_25381,N_22069,N_22036);
nand U25382 (N_25382,N_23012,N_22040);
xnor U25383 (N_25383,N_23105,N_23042);
nand U25384 (N_25384,N_23342,N_22281);
or U25385 (N_25385,N_22103,N_22693);
nand U25386 (N_25386,N_22146,N_23152);
or U25387 (N_25387,N_22795,N_23400);
xor U25388 (N_25388,N_22020,N_23673);
nor U25389 (N_25389,N_22061,N_22118);
nand U25390 (N_25390,N_23901,N_23604);
nor U25391 (N_25391,N_23681,N_23218);
nor U25392 (N_25392,N_22321,N_23326);
or U25393 (N_25393,N_23478,N_23672);
nor U25394 (N_25394,N_23379,N_23196);
nor U25395 (N_25395,N_23556,N_23016);
and U25396 (N_25396,N_23665,N_22524);
nor U25397 (N_25397,N_23136,N_23810);
or U25398 (N_25398,N_22289,N_22238);
nor U25399 (N_25399,N_22594,N_23822);
nor U25400 (N_25400,N_22171,N_23289);
nand U25401 (N_25401,N_23030,N_22153);
and U25402 (N_25402,N_22378,N_22647);
or U25403 (N_25403,N_22786,N_22577);
xnor U25404 (N_25404,N_23154,N_23355);
and U25405 (N_25405,N_22944,N_22254);
nor U25406 (N_25406,N_23196,N_22069);
nand U25407 (N_25407,N_23076,N_23653);
nand U25408 (N_25408,N_23215,N_22870);
nand U25409 (N_25409,N_23114,N_23565);
nor U25410 (N_25410,N_22538,N_23098);
or U25411 (N_25411,N_23638,N_22835);
xnor U25412 (N_25412,N_23677,N_22782);
xnor U25413 (N_25413,N_23841,N_23330);
nand U25414 (N_25414,N_23840,N_23187);
nand U25415 (N_25415,N_23979,N_22352);
or U25416 (N_25416,N_22713,N_23688);
nand U25417 (N_25417,N_22498,N_23261);
nand U25418 (N_25418,N_22485,N_23672);
nand U25419 (N_25419,N_22925,N_23723);
and U25420 (N_25420,N_22911,N_22231);
or U25421 (N_25421,N_23165,N_22065);
xnor U25422 (N_25422,N_23566,N_22722);
or U25423 (N_25423,N_23549,N_22918);
or U25424 (N_25424,N_23339,N_22913);
or U25425 (N_25425,N_23330,N_23010);
or U25426 (N_25426,N_22504,N_22160);
xor U25427 (N_25427,N_22022,N_23014);
nor U25428 (N_25428,N_22226,N_23576);
and U25429 (N_25429,N_22467,N_22118);
and U25430 (N_25430,N_23239,N_23683);
and U25431 (N_25431,N_22353,N_22197);
nand U25432 (N_25432,N_22747,N_22168);
nor U25433 (N_25433,N_23646,N_23806);
nor U25434 (N_25434,N_22068,N_23113);
xor U25435 (N_25435,N_22811,N_22748);
or U25436 (N_25436,N_22454,N_22803);
or U25437 (N_25437,N_22622,N_23667);
nand U25438 (N_25438,N_23595,N_22777);
nand U25439 (N_25439,N_22191,N_22018);
nor U25440 (N_25440,N_22923,N_23933);
and U25441 (N_25441,N_23919,N_23941);
nand U25442 (N_25442,N_22196,N_22305);
or U25443 (N_25443,N_22694,N_23033);
xor U25444 (N_25444,N_22524,N_23562);
and U25445 (N_25445,N_23306,N_23603);
nand U25446 (N_25446,N_23981,N_23098);
nand U25447 (N_25447,N_22652,N_23751);
and U25448 (N_25448,N_23528,N_23600);
nor U25449 (N_25449,N_22990,N_22273);
or U25450 (N_25450,N_23565,N_22326);
nor U25451 (N_25451,N_23340,N_23040);
nand U25452 (N_25452,N_23364,N_22840);
xor U25453 (N_25453,N_23193,N_23454);
xnor U25454 (N_25454,N_23644,N_23441);
nor U25455 (N_25455,N_23088,N_22738);
xor U25456 (N_25456,N_23529,N_23604);
nor U25457 (N_25457,N_22231,N_22018);
xnor U25458 (N_25458,N_22435,N_22842);
and U25459 (N_25459,N_23205,N_22422);
xnor U25460 (N_25460,N_23028,N_22710);
or U25461 (N_25461,N_23490,N_23087);
or U25462 (N_25462,N_23110,N_23831);
xnor U25463 (N_25463,N_23154,N_23937);
and U25464 (N_25464,N_22916,N_22107);
or U25465 (N_25465,N_23460,N_23436);
and U25466 (N_25466,N_22611,N_22782);
xnor U25467 (N_25467,N_23301,N_23177);
or U25468 (N_25468,N_23420,N_23260);
nand U25469 (N_25469,N_22000,N_23500);
and U25470 (N_25470,N_22540,N_22349);
nor U25471 (N_25471,N_22912,N_23472);
and U25472 (N_25472,N_22728,N_22693);
or U25473 (N_25473,N_22189,N_23341);
and U25474 (N_25474,N_22211,N_22586);
xor U25475 (N_25475,N_22331,N_22226);
nor U25476 (N_25476,N_22361,N_23615);
nor U25477 (N_25477,N_23323,N_23832);
xor U25478 (N_25478,N_22075,N_23603);
xnor U25479 (N_25479,N_23140,N_22357);
or U25480 (N_25480,N_22805,N_23880);
nand U25481 (N_25481,N_23282,N_23148);
and U25482 (N_25482,N_23331,N_23576);
nand U25483 (N_25483,N_23146,N_23700);
or U25484 (N_25484,N_23037,N_23290);
and U25485 (N_25485,N_23071,N_22392);
xnor U25486 (N_25486,N_22121,N_23760);
nand U25487 (N_25487,N_22612,N_22153);
nand U25488 (N_25488,N_22856,N_23822);
xor U25489 (N_25489,N_22166,N_23029);
and U25490 (N_25490,N_23632,N_23725);
or U25491 (N_25491,N_23791,N_23377);
or U25492 (N_25492,N_23833,N_22434);
nand U25493 (N_25493,N_22966,N_23200);
or U25494 (N_25494,N_22385,N_22529);
or U25495 (N_25495,N_23707,N_23763);
and U25496 (N_25496,N_23596,N_23258);
xnor U25497 (N_25497,N_22205,N_22807);
nor U25498 (N_25498,N_22979,N_22880);
nand U25499 (N_25499,N_23698,N_22451);
and U25500 (N_25500,N_22880,N_22207);
xor U25501 (N_25501,N_23402,N_22366);
nor U25502 (N_25502,N_22666,N_22074);
and U25503 (N_25503,N_23679,N_23608);
nor U25504 (N_25504,N_22877,N_23099);
xnor U25505 (N_25505,N_23803,N_23717);
and U25506 (N_25506,N_22654,N_22271);
and U25507 (N_25507,N_22437,N_23044);
xor U25508 (N_25508,N_23480,N_23286);
xor U25509 (N_25509,N_23214,N_23537);
or U25510 (N_25510,N_23864,N_22048);
nand U25511 (N_25511,N_22116,N_22602);
or U25512 (N_25512,N_23829,N_22557);
xnor U25513 (N_25513,N_23374,N_23720);
and U25514 (N_25514,N_23402,N_22630);
or U25515 (N_25515,N_23204,N_22476);
nand U25516 (N_25516,N_23172,N_23390);
xor U25517 (N_25517,N_23471,N_22806);
and U25518 (N_25518,N_23042,N_23600);
nor U25519 (N_25519,N_23478,N_22440);
nand U25520 (N_25520,N_23344,N_22339);
or U25521 (N_25521,N_22174,N_23877);
and U25522 (N_25522,N_22389,N_22898);
nand U25523 (N_25523,N_23486,N_23467);
nor U25524 (N_25524,N_22070,N_22468);
and U25525 (N_25525,N_23536,N_22733);
or U25526 (N_25526,N_22363,N_23629);
xnor U25527 (N_25527,N_22675,N_22599);
xor U25528 (N_25528,N_22416,N_22736);
nor U25529 (N_25529,N_23334,N_22834);
xor U25530 (N_25530,N_22643,N_22220);
xnor U25531 (N_25531,N_22278,N_22392);
nand U25532 (N_25532,N_22302,N_23824);
and U25533 (N_25533,N_23002,N_22158);
xor U25534 (N_25534,N_23045,N_23235);
and U25535 (N_25535,N_23720,N_23541);
xor U25536 (N_25536,N_22004,N_22950);
nor U25537 (N_25537,N_23520,N_22080);
nand U25538 (N_25538,N_22191,N_22900);
nand U25539 (N_25539,N_22131,N_22483);
xor U25540 (N_25540,N_23211,N_22079);
xor U25541 (N_25541,N_23238,N_22581);
and U25542 (N_25542,N_22633,N_22175);
and U25543 (N_25543,N_22338,N_22624);
or U25544 (N_25544,N_22594,N_22656);
and U25545 (N_25545,N_23757,N_22315);
xnor U25546 (N_25546,N_22032,N_22662);
nand U25547 (N_25547,N_22832,N_22903);
nor U25548 (N_25548,N_22472,N_23183);
xor U25549 (N_25549,N_23094,N_23888);
xor U25550 (N_25550,N_22627,N_23999);
or U25551 (N_25551,N_23617,N_22581);
nand U25552 (N_25552,N_22271,N_23453);
nor U25553 (N_25553,N_22676,N_22228);
and U25554 (N_25554,N_22013,N_22407);
or U25555 (N_25555,N_22171,N_22986);
and U25556 (N_25556,N_22147,N_22456);
or U25557 (N_25557,N_22807,N_23688);
xnor U25558 (N_25558,N_23992,N_23875);
nor U25559 (N_25559,N_23904,N_23934);
nand U25560 (N_25560,N_22683,N_23409);
or U25561 (N_25561,N_22940,N_23676);
nand U25562 (N_25562,N_23806,N_22831);
or U25563 (N_25563,N_22055,N_23202);
or U25564 (N_25564,N_22607,N_23973);
and U25565 (N_25565,N_22095,N_22115);
or U25566 (N_25566,N_23890,N_22061);
or U25567 (N_25567,N_23645,N_22384);
nand U25568 (N_25568,N_22431,N_22700);
xor U25569 (N_25569,N_23651,N_23426);
nor U25570 (N_25570,N_22106,N_22675);
xnor U25571 (N_25571,N_22012,N_22191);
nand U25572 (N_25572,N_23300,N_22275);
nor U25573 (N_25573,N_23935,N_22914);
nand U25574 (N_25574,N_22349,N_23308);
and U25575 (N_25575,N_22218,N_23122);
nand U25576 (N_25576,N_23262,N_23821);
nor U25577 (N_25577,N_22895,N_23615);
xor U25578 (N_25578,N_22067,N_22549);
xnor U25579 (N_25579,N_23803,N_22020);
nor U25580 (N_25580,N_23138,N_22294);
nand U25581 (N_25581,N_22841,N_23283);
or U25582 (N_25582,N_23528,N_23674);
nor U25583 (N_25583,N_22106,N_23194);
nor U25584 (N_25584,N_23703,N_22912);
or U25585 (N_25585,N_23567,N_23345);
nor U25586 (N_25586,N_23650,N_22939);
nor U25587 (N_25587,N_23604,N_23403);
and U25588 (N_25588,N_22176,N_23324);
xor U25589 (N_25589,N_22350,N_23597);
and U25590 (N_25590,N_22211,N_22378);
and U25591 (N_25591,N_22821,N_22165);
or U25592 (N_25592,N_22825,N_22251);
nor U25593 (N_25593,N_22041,N_22599);
nor U25594 (N_25594,N_22147,N_23089);
and U25595 (N_25595,N_22327,N_22778);
nand U25596 (N_25596,N_22515,N_22570);
and U25597 (N_25597,N_22753,N_22009);
and U25598 (N_25598,N_23394,N_23251);
nand U25599 (N_25599,N_22202,N_23431);
or U25600 (N_25600,N_23275,N_23325);
nor U25601 (N_25601,N_23306,N_22222);
and U25602 (N_25602,N_23066,N_22672);
xnor U25603 (N_25603,N_23641,N_22456);
or U25604 (N_25604,N_22556,N_22644);
nor U25605 (N_25605,N_22640,N_22413);
and U25606 (N_25606,N_23593,N_22561);
nor U25607 (N_25607,N_23221,N_22179);
and U25608 (N_25608,N_23591,N_23981);
xor U25609 (N_25609,N_22790,N_22541);
and U25610 (N_25610,N_23685,N_23968);
xnor U25611 (N_25611,N_23685,N_22256);
xor U25612 (N_25612,N_22411,N_23211);
or U25613 (N_25613,N_22960,N_23489);
or U25614 (N_25614,N_22426,N_22956);
nor U25615 (N_25615,N_22422,N_23822);
nor U25616 (N_25616,N_23899,N_22271);
and U25617 (N_25617,N_22318,N_22111);
xor U25618 (N_25618,N_23983,N_22247);
or U25619 (N_25619,N_22582,N_22290);
and U25620 (N_25620,N_23938,N_23558);
nor U25621 (N_25621,N_23428,N_23445);
nand U25622 (N_25622,N_22290,N_22550);
or U25623 (N_25623,N_22257,N_23277);
nor U25624 (N_25624,N_23027,N_23790);
xnor U25625 (N_25625,N_23255,N_22587);
nand U25626 (N_25626,N_22526,N_23050);
nor U25627 (N_25627,N_22776,N_23793);
nand U25628 (N_25628,N_23233,N_22579);
and U25629 (N_25629,N_22523,N_22194);
or U25630 (N_25630,N_22564,N_23722);
or U25631 (N_25631,N_22199,N_22328);
nand U25632 (N_25632,N_23578,N_23004);
and U25633 (N_25633,N_23886,N_23564);
nand U25634 (N_25634,N_22146,N_22588);
xor U25635 (N_25635,N_22429,N_22616);
and U25636 (N_25636,N_23422,N_22627);
and U25637 (N_25637,N_23028,N_22452);
xnor U25638 (N_25638,N_23037,N_23963);
nand U25639 (N_25639,N_22699,N_22256);
xor U25640 (N_25640,N_22980,N_22490);
xor U25641 (N_25641,N_22574,N_23533);
nand U25642 (N_25642,N_23047,N_22770);
or U25643 (N_25643,N_22461,N_23116);
or U25644 (N_25644,N_22937,N_22808);
nand U25645 (N_25645,N_23858,N_23386);
xnor U25646 (N_25646,N_23605,N_23491);
nand U25647 (N_25647,N_23732,N_23262);
xor U25648 (N_25648,N_23335,N_23726);
or U25649 (N_25649,N_23903,N_23718);
and U25650 (N_25650,N_23464,N_23374);
and U25651 (N_25651,N_23713,N_23227);
xor U25652 (N_25652,N_22521,N_22764);
nor U25653 (N_25653,N_23602,N_23752);
nor U25654 (N_25654,N_22099,N_22102);
or U25655 (N_25655,N_22864,N_23057);
or U25656 (N_25656,N_23476,N_23746);
nand U25657 (N_25657,N_22998,N_22914);
nor U25658 (N_25658,N_22680,N_22990);
nand U25659 (N_25659,N_22090,N_22732);
and U25660 (N_25660,N_22810,N_23088);
or U25661 (N_25661,N_22840,N_22441);
and U25662 (N_25662,N_23085,N_22132);
and U25663 (N_25663,N_23625,N_22030);
and U25664 (N_25664,N_22851,N_22312);
xnor U25665 (N_25665,N_23359,N_22774);
nor U25666 (N_25666,N_22172,N_23120);
and U25667 (N_25667,N_22974,N_23028);
nor U25668 (N_25668,N_22763,N_22385);
or U25669 (N_25669,N_22842,N_23170);
xor U25670 (N_25670,N_22381,N_23121);
nand U25671 (N_25671,N_22163,N_23134);
and U25672 (N_25672,N_22692,N_22157);
nor U25673 (N_25673,N_23948,N_23769);
nand U25674 (N_25674,N_23410,N_23275);
xor U25675 (N_25675,N_22198,N_22147);
xnor U25676 (N_25676,N_23107,N_23338);
nor U25677 (N_25677,N_22619,N_23689);
nand U25678 (N_25678,N_22188,N_23962);
or U25679 (N_25679,N_22908,N_22543);
nor U25680 (N_25680,N_23523,N_22510);
or U25681 (N_25681,N_23957,N_22849);
nand U25682 (N_25682,N_22666,N_22276);
nand U25683 (N_25683,N_23998,N_22273);
and U25684 (N_25684,N_23710,N_22287);
or U25685 (N_25685,N_22373,N_22027);
xor U25686 (N_25686,N_23293,N_23913);
nand U25687 (N_25687,N_22205,N_23770);
or U25688 (N_25688,N_23714,N_23712);
and U25689 (N_25689,N_22249,N_22540);
xor U25690 (N_25690,N_22618,N_22800);
xor U25691 (N_25691,N_23955,N_23371);
or U25692 (N_25692,N_22350,N_23015);
nor U25693 (N_25693,N_22969,N_23491);
or U25694 (N_25694,N_22246,N_22615);
or U25695 (N_25695,N_23223,N_22804);
or U25696 (N_25696,N_22661,N_22508);
nor U25697 (N_25697,N_23594,N_23004);
nand U25698 (N_25698,N_22419,N_23116);
or U25699 (N_25699,N_23383,N_23925);
and U25700 (N_25700,N_22930,N_22840);
nand U25701 (N_25701,N_22795,N_22146);
xor U25702 (N_25702,N_23144,N_22448);
and U25703 (N_25703,N_23715,N_23489);
and U25704 (N_25704,N_22057,N_23462);
nor U25705 (N_25705,N_23952,N_23134);
and U25706 (N_25706,N_23569,N_22289);
nor U25707 (N_25707,N_23346,N_22448);
or U25708 (N_25708,N_23647,N_22157);
xor U25709 (N_25709,N_23548,N_23114);
xnor U25710 (N_25710,N_23714,N_23479);
nand U25711 (N_25711,N_23095,N_23624);
nor U25712 (N_25712,N_23257,N_22962);
nand U25713 (N_25713,N_23712,N_22507);
xor U25714 (N_25714,N_22432,N_23012);
nor U25715 (N_25715,N_23601,N_22716);
or U25716 (N_25716,N_23789,N_22427);
xnor U25717 (N_25717,N_22159,N_22068);
and U25718 (N_25718,N_23987,N_23007);
or U25719 (N_25719,N_23579,N_23413);
or U25720 (N_25720,N_22115,N_22502);
nand U25721 (N_25721,N_22680,N_23167);
nor U25722 (N_25722,N_22510,N_23146);
xnor U25723 (N_25723,N_22942,N_22445);
or U25724 (N_25724,N_23226,N_23056);
xnor U25725 (N_25725,N_23148,N_23974);
nor U25726 (N_25726,N_23331,N_23485);
xor U25727 (N_25727,N_23394,N_22673);
xor U25728 (N_25728,N_23521,N_22531);
xnor U25729 (N_25729,N_22128,N_23405);
nor U25730 (N_25730,N_22669,N_22178);
and U25731 (N_25731,N_22685,N_23023);
xnor U25732 (N_25732,N_22280,N_22981);
and U25733 (N_25733,N_23137,N_22727);
nand U25734 (N_25734,N_23034,N_23510);
xor U25735 (N_25735,N_23022,N_23229);
nand U25736 (N_25736,N_23137,N_22242);
and U25737 (N_25737,N_23726,N_23992);
and U25738 (N_25738,N_22802,N_22842);
xnor U25739 (N_25739,N_23187,N_23136);
nor U25740 (N_25740,N_23644,N_22911);
and U25741 (N_25741,N_22288,N_22250);
nor U25742 (N_25742,N_23495,N_23343);
xor U25743 (N_25743,N_22989,N_23474);
nor U25744 (N_25744,N_22171,N_23133);
or U25745 (N_25745,N_23342,N_22363);
or U25746 (N_25746,N_23709,N_22039);
xor U25747 (N_25747,N_23710,N_23609);
nand U25748 (N_25748,N_23838,N_23312);
nand U25749 (N_25749,N_23497,N_22080);
and U25750 (N_25750,N_23008,N_23029);
nand U25751 (N_25751,N_22102,N_23413);
and U25752 (N_25752,N_22861,N_22604);
and U25753 (N_25753,N_22566,N_22018);
xnor U25754 (N_25754,N_23980,N_23517);
or U25755 (N_25755,N_23643,N_23480);
nand U25756 (N_25756,N_23104,N_23335);
and U25757 (N_25757,N_22166,N_22550);
nand U25758 (N_25758,N_23543,N_23307);
xor U25759 (N_25759,N_23158,N_23359);
nand U25760 (N_25760,N_22534,N_23321);
nor U25761 (N_25761,N_23393,N_23401);
nand U25762 (N_25762,N_22165,N_23370);
nor U25763 (N_25763,N_22598,N_23428);
and U25764 (N_25764,N_22645,N_22699);
nand U25765 (N_25765,N_23329,N_22614);
and U25766 (N_25766,N_22743,N_23982);
or U25767 (N_25767,N_23301,N_23829);
xor U25768 (N_25768,N_23323,N_22379);
nor U25769 (N_25769,N_23834,N_22454);
and U25770 (N_25770,N_22264,N_23724);
and U25771 (N_25771,N_23626,N_23062);
and U25772 (N_25772,N_22049,N_23547);
nor U25773 (N_25773,N_22990,N_22247);
nor U25774 (N_25774,N_22682,N_23082);
and U25775 (N_25775,N_23958,N_23450);
xnor U25776 (N_25776,N_23210,N_23844);
nand U25777 (N_25777,N_23492,N_23734);
and U25778 (N_25778,N_23656,N_22698);
nor U25779 (N_25779,N_23739,N_22490);
or U25780 (N_25780,N_22907,N_23013);
nor U25781 (N_25781,N_22953,N_22637);
xnor U25782 (N_25782,N_22728,N_22205);
or U25783 (N_25783,N_22674,N_22238);
or U25784 (N_25784,N_22202,N_22460);
nand U25785 (N_25785,N_22448,N_23437);
and U25786 (N_25786,N_23700,N_22226);
and U25787 (N_25787,N_23583,N_22594);
or U25788 (N_25788,N_23071,N_23953);
or U25789 (N_25789,N_23709,N_22055);
xor U25790 (N_25790,N_23765,N_23744);
xor U25791 (N_25791,N_23888,N_23029);
and U25792 (N_25792,N_23840,N_22192);
and U25793 (N_25793,N_23925,N_22119);
nand U25794 (N_25794,N_22605,N_22949);
nand U25795 (N_25795,N_23469,N_23855);
nand U25796 (N_25796,N_23395,N_23113);
nor U25797 (N_25797,N_23430,N_22920);
and U25798 (N_25798,N_22986,N_22155);
nand U25799 (N_25799,N_22215,N_23921);
and U25800 (N_25800,N_22346,N_23917);
xor U25801 (N_25801,N_23317,N_22960);
and U25802 (N_25802,N_22483,N_22574);
nand U25803 (N_25803,N_23337,N_23272);
nand U25804 (N_25804,N_22072,N_23321);
nand U25805 (N_25805,N_22835,N_22136);
xor U25806 (N_25806,N_22725,N_23049);
nand U25807 (N_25807,N_22311,N_22434);
nand U25808 (N_25808,N_22872,N_22762);
nor U25809 (N_25809,N_23957,N_22878);
nand U25810 (N_25810,N_22555,N_23725);
or U25811 (N_25811,N_22933,N_23659);
xor U25812 (N_25812,N_22278,N_22334);
or U25813 (N_25813,N_23348,N_23616);
and U25814 (N_25814,N_22083,N_23240);
xor U25815 (N_25815,N_22567,N_23876);
nand U25816 (N_25816,N_23732,N_23376);
or U25817 (N_25817,N_23718,N_22846);
nand U25818 (N_25818,N_23895,N_22417);
xor U25819 (N_25819,N_23138,N_23453);
nor U25820 (N_25820,N_22333,N_22397);
nand U25821 (N_25821,N_22033,N_22615);
xnor U25822 (N_25822,N_22991,N_23021);
nor U25823 (N_25823,N_23622,N_23782);
nor U25824 (N_25824,N_22157,N_22999);
nor U25825 (N_25825,N_22483,N_23244);
nand U25826 (N_25826,N_22459,N_22927);
nor U25827 (N_25827,N_23516,N_22833);
nor U25828 (N_25828,N_22502,N_22825);
nor U25829 (N_25829,N_23030,N_22613);
and U25830 (N_25830,N_22444,N_22120);
nand U25831 (N_25831,N_23139,N_22373);
and U25832 (N_25832,N_23353,N_22499);
or U25833 (N_25833,N_23592,N_22377);
xnor U25834 (N_25834,N_23807,N_23251);
or U25835 (N_25835,N_23054,N_23487);
nand U25836 (N_25836,N_23036,N_23108);
and U25837 (N_25837,N_23848,N_23547);
or U25838 (N_25838,N_23276,N_23145);
or U25839 (N_25839,N_23575,N_22895);
and U25840 (N_25840,N_22729,N_23013);
or U25841 (N_25841,N_23839,N_23003);
xor U25842 (N_25842,N_22301,N_22206);
xnor U25843 (N_25843,N_23548,N_22430);
or U25844 (N_25844,N_23099,N_22996);
nor U25845 (N_25845,N_23164,N_22759);
nand U25846 (N_25846,N_23547,N_22536);
or U25847 (N_25847,N_23000,N_22724);
and U25848 (N_25848,N_23769,N_23397);
nor U25849 (N_25849,N_23164,N_22899);
and U25850 (N_25850,N_22864,N_22153);
or U25851 (N_25851,N_22437,N_22629);
and U25852 (N_25852,N_22878,N_22276);
or U25853 (N_25853,N_22442,N_23109);
and U25854 (N_25854,N_22887,N_23103);
xnor U25855 (N_25855,N_23956,N_22532);
xor U25856 (N_25856,N_23162,N_23835);
xnor U25857 (N_25857,N_22649,N_23066);
nor U25858 (N_25858,N_23073,N_23624);
nor U25859 (N_25859,N_23776,N_22702);
nand U25860 (N_25860,N_23857,N_23897);
or U25861 (N_25861,N_22029,N_22698);
nand U25862 (N_25862,N_22597,N_22020);
and U25863 (N_25863,N_23310,N_23551);
and U25864 (N_25864,N_22827,N_22685);
and U25865 (N_25865,N_23072,N_22209);
and U25866 (N_25866,N_23998,N_23823);
and U25867 (N_25867,N_23139,N_23956);
xnor U25868 (N_25868,N_23053,N_22205);
xnor U25869 (N_25869,N_23365,N_23470);
or U25870 (N_25870,N_23245,N_23041);
xnor U25871 (N_25871,N_22978,N_23251);
nor U25872 (N_25872,N_23518,N_23040);
or U25873 (N_25873,N_23468,N_23685);
nor U25874 (N_25874,N_22677,N_23582);
xnor U25875 (N_25875,N_22838,N_23948);
or U25876 (N_25876,N_22752,N_22647);
nor U25877 (N_25877,N_22762,N_22036);
or U25878 (N_25878,N_22779,N_23365);
and U25879 (N_25879,N_23527,N_23103);
and U25880 (N_25880,N_23774,N_22096);
nand U25881 (N_25881,N_23016,N_23234);
nor U25882 (N_25882,N_22485,N_22649);
and U25883 (N_25883,N_23600,N_22818);
or U25884 (N_25884,N_22685,N_23380);
and U25885 (N_25885,N_22813,N_22932);
nand U25886 (N_25886,N_22285,N_23296);
nor U25887 (N_25887,N_23025,N_23120);
nor U25888 (N_25888,N_23513,N_23546);
or U25889 (N_25889,N_22077,N_23636);
nor U25890 (N_25890,N_22502,N_23501);
xnor U25891 (N_25891,N_22364,N_22229);
nor U25892 (N_25892,N_23620,N_23340);
or U25893 (N_25893,N_23459,N_22489);
nand U25894 (N_25894,N_23557,N_23830);
and U25895 (N_25895,N_22082,N_22433);
or U25896 (N_25896,N_23771,N_23872);
nor U25897 (N_25897,N_23972,N_23705);
and U25898 (N_25898,N_22013,N_22992);
or U25899 (N_25899,N_23915,N_22520);
nand U25900 (N_25900,N_22590,N_22181);
xor U25901 (N_25901,N_22063,N_23416);
and U25902 (N_25902,N_22216,N_22347);
xor U25903 (N_25903,N_23335,N_22961);
and U25904 (N_25904,N_23165,N_22262);
or U25905 (N_25905,N_22335,N_22553);
xnor U25906 (N_25906,N_23315,N_22906);
and U25907 (N_25907,N_23655,N_23816);
or U25908 (N_25908,N_23165,N_23032);
nand U25909 (N_25909,N_22577,N_22092);
or U25910 (N_25910,N_23189,N_22137);
xnor U25911 (N_25911,N_23409,N_22073);
or U25912 (N_25912,N_23245,N_22030);
and U25913 (N_25913,N_22383,N_22191);
nand U25914 (N_25914,N_23061,N_22837);
nand U25915 (N_25915,N_23066,N_22012);
nor U25916 (N_25916,N_22255,N_23314);
nand U25917 (N_25917,N_22615,N_23538);
xnor U25918 (N_25918,N_23797,N_23735);
nor U25919 (N_25919,N_23513,N_22295);
xor U25920 (N_25920,N_23073,N_23713);
and U25921 (N_25921,N_23479,N_23662);
or U25922 (N_25922,N_22456,N_22722);
or U25923 (N_25923,N_23068,N_22695);
and U25924 (N_25924,N_22211,N_22591);
and U25925 (N_25925,N_22119,N_22791);
xor U25926 (N_25926,N_22708,N_23861);
xnor U25927 (N_25927,N_22024,N_23261);
or U25928 (N_25928,N_23624,N_23813);
and U25929 (N_25929,N_23329,N_22913);
nand U25930 (N_25930,N_23172,N_22785);
xnor U25931 (N_25931,N_23710,N_23062);
nor U25932 (N_25932,N_22846,N_22801);
and U25933 (N_25933,N_23417,N_22159);
and U25934 (N_25934,N_23372,N_22029);
xor U25935 (N_25935,N_23259,N_23360);
or U25936 (N_25936,N_22215,N_22360);
and U25937 (N_25937,N_23735,N_23196);
nor U25938 (N_25938,N_23400,N_23290);
and U25939 (N_25939,N_22357,N_23333);
xnor U25940 (N_25940,N_22653,N_23824);
and U25941 (N_25941,N_22366,N_23753);
and U25942 (N_25942,N_23663,N_22725);
nand U25943 (N_25943,N_23777,N_22963);
nor U25944 (N_25944,N_23199,N_23697);
nand U25945 (N_25945,N_23902,N_22974);
nand U25946 (N_25946,N_23763,N_23720);
or U25947 (N_25947,N_22069,N_22805);
xnor U25948 (N_25948,N_22672,N_22443);
nor U25949 (N_25949,N_23380,N_23867);
or U25950 (N_25950,N_22013,N_23333);
xnor U25951 (N_25951,N_22587,N_23909);
xor U25952 (N_25952,N_23865,N_23282);
xnor U25953 (N_25953,N_23816,N_23331);
nand U25954 (N_25954,N_23772,N_22844);
nand U25955 (N_25955,N_22437,N_23188);
and U25956 (N_25956,N_23189,N_22696);
xor U25957 (N_25957,N_23436,N_23708);
nand U25958 (N_25958,N_22701,N_22713);
and U25959 (N_25959,N_22459,N_22795);
or U25960 (N_25960,N_23678,N_22424);
nor U25961 (N_25961,N_22651,N_22368);
or U25962 (N_25962,N_22823,N_23482);
and U25963 (N_25963,N_23949,N_22716);
xor U25964 (N_25964,N_22920,N_22974);
nor U25965 (N_25965,N_23021,N_22571);
xor U25966 (N_25966,N_22550,N_23161);
and U25967 (N_25967,N_22443,N_23273);
xor U25968 (N_25968,N_22591,N_23622);
nand U25969 (N_25969,N_22573,N_23577);
and U25970 (N_25970,N_22917,N_23843);
nor U25971 (N_25971,N_23687,N_22283);
nand U25972 (N_25972,N_23393,N_22261);
nor U25973 (N_25973,N_23689,N_22789);
nor U25974 (N_25974,N_22889,N_22479);
and U25975 (N_25975,N_22149,N_22776);
and U25976 (N_25976,N_22058,N_23158);
xor U25977 (N_25977,N_23290,N_23801);
or U25978 (N_25978,N_22094,N_23341);
or U25979 (N_25979,N_23035,N_23130);
nand U25980 (N_25980,N_22584,N_23628);
nand U25981 (N_25981,N_23528,N_22047);
xor U25982 (N_25982,N_23576,N_23874);
xnor U25983 (N_25983,N_23096,N_22487);
xor U25984 (N_25984,N_23321,N_23636);
and U25985 (N_25985,N_22316,N_23379);
and U25986 (N_25986,N_22044,N_23818);
xor U25987 (N_25987,N_23012,N_22225);
xor U25988 (N_25988,N_22217,N_23355);
nor U25989 (N_25989,N_23210,N_22948);
nor U25990 (N_25990,N_23353,N_22917);
xor U25991 (N_25991,N_22927,N_22380);
nand U25992 (N_25992,N_23867,N_22084);
or U25993 (N_25993,N_22976,N_23239);
nor U25994 (N_25994,N_22818,N_22049);
xor U25995 (N_25995,N_22530,N_22732);
or U25996 (N_25996,N_22914,N_22717);
nand U25997 (N_25997,N_22426,N_23826);
and U25998 (N_25998,N_23049,N_23818);
and U25999 (N_25999,N_23167,N_23854);
nor U26000 (N_26000,N_24517,N_24258);
and U26001 (N_26001,N_24799,N_24073);
nand U26002 (N_26002,N_24233,N_25282);
nor U26003 (N_26003,N_25456,N_25170);
nor U26004 (N_26004,N_25213,N_25645);
nand U26005 (N_26005,N_24198,N_24087);
nor U26006 (N_26006,N_24278,N_24541);
xnor U26007 (N_26007,N_25537,N_25770);
and U26008 (N_26008,N_25006,N_24898);
nor U26009 (N_26009,N_24753,N_25246);
and U26010 (N_26010,N_25191,N_25382);
xor U26011 (N_26011,N_24165,N_24305);
nand U26012 (N_26012,N_24811,N_24132);
nand U26013 (N_26013,N_25872,N_25061);
or U26014 (N_26014,N_24442,N_24300);
or U26015 (N_26015,N_25990,N_25357);
or U26016 (N_26016,N_25577,N_24255);
xor U26017 (N_26017,N_25559,N_24622);
or U26018 (N_26018,N_25344,N_25153);
nand U26019 (N_26019,N_24341,N_25882);
xor U26020 (N_26020,N_25807,N_24130);
xnor U26021 (N_26021,N_24729,N_24352);
or U26022 (N_26022,N_25998,N_25301);
and U26023 (N_26023,N_25858,N_25830);
and U26024 (N_26024,N_25777,N_25734);
nor U26025 (N_26025,N_24791,N_24543);
and U26026 (N_26026,N_25556,N_25760);
or U26027 (N_26027,N_24146,N_24690);
nor U26028 (N_26028,N_25339,N_24206);
xor U26029 (N_26029,N_25322,N_25219);
xor U26030 (N_26030,N_25893,N_25319);
and U26031 (N_26031,N_24597,N_25944);
nand U26032 (N_26032,N_24518,N_24426);
or U26033 (N_26033,N_25979,N_25057);
nor U26034 (N_26034,N_25750,N_25673);
and U26035 (N_26035,N_24742,N_24997);
and U26036 (N_26036,N_25193,N_24557);
nand U26037 (N_26037,N_25054,N_24998);
and U26038 (N_26038,N_24814,N_24995);
nor U26039 (N_26039,N_25634,N_24480);
xor U26040 (N_26040,N_25294,N_24826);
or U26041 (N_26041,N_24065,N_24717);
or U26042 (N_26042,N_25343,N_25288);
and U26043 (N_26043,N_25171,N_25501);
or U26044 (N_26044,N_25936,N_24144);
and U26045 (N_26045,N_25692,N_25053);
xor U26046 (N_26046,N_25351,N_25355);
nand U26047 (N_26047,N_25894,N_25615);
xor U26048 (N_26048,N_24568,N_24931);
and U26049 (N_26049,N_25334,N_24909);
nand U26050 (N_26050,N_24281,N_25480);
nor U26051 (N_26051,N_24009,N_24266);
nand U26052 (N_26052,N_24496,N_25066);
xor U26053 (N_26053,N_25503,N_24743);
nand U26054 (N_26054,N_24611,N_24272);
and U26055 (N_26055,N_24421,N_24427);
or U26056 (N_26056,N_25557,N_25237);
nand U26057 (N_26057,N_25425,N_25426);
and U26058 (N_26058,N_25011,N_25534);
and U26059 (N_26059,N_25899,N_25100);
nand U26060 (N_26060,N_25746,N_25454);
or U26061 (N_26061,N_25012,N_24126);
nand U26062 (N_26062,N_24918,N_24225);
or U26063 (N_26063,N_25016,N_24306);
nor U26064 (N_26064,N_24121,N_24409);
and U26065 (N_26065,N_24714,N_25187);
nand U26066 (N_26066,N_25890,N_24755);
xor U26067 (N_26067,N_25423,N_25310);
nand U26068 (N_26068,N_24026,N_25867);
nor U26069 (N_26069,N_25010,N_24606);
nand U26070 (N_26070,N_25020,N_25044);
and U26071 (N_26071,N_24860,N_24882);
or U26072 (N_26072,N_25951,N_24808);
or U26073 (N_26073,N_25657,N_24946);
or U26074 (N_26074,N_24895,N_24941);
nor U26075 (N_26075,N_25045,N_24375);
xor U26076 (N_26076,N_25875,N_24044);
xor U26077 (N_26077,N_25140,N_24599);
and U26078 (N_26078,N_25749,N_24419);
or U26079 (N_26079,N_25983,N_24884);
xnor U26080 (N_26080,N_24361,N_24522);
and U26081 (N_26081,N_24360,N_25304);
xnor U26082 (N_26082,N_24962,N_24436);
nor U26083 (N_26083,N_24953,N_24711);
xor U26084 (N_26084,N_25421,N_24721);
nor U26085 (N_26085,N_24444,N_24822);
xnor U26086 (N_26086,N_24735,N_24745);
nor U26087 (N_26087,N_24561,N_25956);
xor U26088 (N_26088,N_25129,N_25758);
nor U26089 (N_26089,N_24046,N_25279);
and U26090 (N_26090,N_24581,N_24520);
and U26091 (N_26091,N_25218,N_25712);
nor U26092 (N_26092,N_24397,N_24900);
nor U26093 (N_26093,N_24944,N_25293);
xnor U26094 (N_26094,N_24798,N_24211);
xor U26095 (N_26095,N_24507,N_25119);
nand U26096 (N_26096,N_24182,N_25582);
nand U26097 (N_26097,N_24892,N_24927);
or U26098 (N_26098,N_25130,N_24293);
nand U26099 (N_26099,N_24567,N_25331);
or U26100 (N_26100,N_25654,N_25079);
xnor U26101 (N_26101,N_24777,N_24248);
or U26102 (N_26102,N_24772,N_24503);
and U26103 (N_26103,N_25623,N_25550);
or U26104 (N_26104,N_24949,N_24162);
nor U26105 (N_26105,N_25136,N_24118);
or U26106 (N_26106,N_25542,N_25833);
nor U26107 (N_26107,N_24940,N_25722);
nor U26108 (N_26108,N_25263,N_25624);
and U26109 (N_26109,N_24367,N_25483);
and U26110 (N_26110,N_25791,N_25773);
nor U26111 (N_26111,N_25707,N_25811);
nor U26112 (N_26112,N_24460,N_25589);
nand U26113 (N_26113,N_24045,N_24506);
or U26114 (N_26114,N_24191,N_24971);
xor U26115 (N_26115,N_25374,N_24230);
nand U26116 (N_26116,N_24369,N_24746);
nand U26117 (N_26117,N_24678,N_24539);
and U26118 (N_26118,N_24751,N_24353);
and U26119 (N_26119,N_25093,N_24364);
and U26120 (N_26120,N_25788,N_24488);
nor U26121 (N_26121,N_25470,N_25451);
nor U26122 (N_26122,N_25055,N_25766);
and U26123 (N_26123,N_24084,N_25461);
nand U26124 (N_26124,N_25243,N_24881);
nor U26125 (N_26125,N_24463,N_24373);
nor U26126 (N_26126,N_25853,N_24642);
and U26127 (N_26127,N_24587,N_25730);
nor U26128 (N_26128,N_25385,N_25447);
nor U26129 (N_26129,N_24528,N_24307);
nor U26130 (N_26130,N_25690,N_24580);
nor U26131 (N_26131,N_25650,N_24308);
and U26132 (N_26132,N_24846,N_25367);
nor U26133 (N_26133,N_24196,N_25158);
or U26134 (N_26134,N_24189,N_25271);
or U26135 (N_26135,N_24773,N_24842);
nand U26136 (N_26136,N_25023,N_25341);
xnor U26137 (N_26137,N_24806,N_25234);
xor U26138 (N_26138,N_24573,N_24035);
xor U26139 (N_26139,N_25786,N_24490);
and U26140 (N_26140,N_25030,N_24276);
nor U26141 (N_26141,N_25256,N_24183);
nor U26142 (N_26142,N_24322,N_24474);
and U26143 (N_26143,N_25849,N_24261);
xnor U26144 (N_26144,N_24218,N_24748);
nor U26145 (N_26145,N_24201,N_25092);
nand U26146 (N_26146,N_24874,N_25124);
and U26147 (N_26147,N_24256,N_25236);
nand U26148 (N_26148,N_24783,N_24075);
xnor U26149 (N_26149,N_25504,N_25659);
and U26150 (N_26150,N_24351,N_25142);
nor U26151 (N_26151,N_24801,N_24952);
or U26152 (N_26152,N_25688,N_24337);
nand U26153 (N_26153,N_24099,N_25097);
or U26154 (N_26154,N_24312,N_25772);
xnor U26155 (N_26155,N_24924,N_24184);
xnor U26156 (N_26156,N_25910,N_25937);
and U26157 (N_26157,N_24890,N_24238);
and U26158 (N_26158,N_24902,N_24487);
and U26159 (N_26159,N_25437,N_24453);
nand U26160 (N_26160,N_25802,N_25507);
or U26161 (N_26161,N_25047,N_24605);
xnor U26162 (N_26162,N_25695,N_25590);
nand U26163 (N_26163,N_25682,N_24468);
and U26164 (N_26164,N_24694,N_25723);
xnor U26165 (N_26165,N_24221,N_25354);
xor U26166 (N_26166,N_25675,N_25416);
xor U26167 (N_26167,N_24072,N_24023);
or U26168 (N_26168,N_24907,N_25596);
xor U26169 (N_26169,N_24164,N_24730);
or U26170 (N_26170,N_25139,N_24310);
and U26171 (N_26171,N_25822,N_25844);
nand U26172 (N_26172,N_24457,N_24534);
nand U26173 (N_26173,N_24876,N_25570);
xor U26174 (N_26174,N_24172,N_24289);
nor U26175 (N_26175,N_24240,N_25608);
and U26176 (N_26176,N_25535,N_24049);
nand U26177 (N_26177,N_25958,N_25434);
nand U26178 (N_26178,N_25088,N_25303);
xor U26179 (N_26179,N_24259,N_24631);
nand U26180 (N_26180,N_25151,N_25267);
or U26181 (N_26181,N_25729,N_25743);
and U26182 (N_26182,N_24537,N_24332);
and U26183 (N_26183,N_24471,N_25629);
and U26184 (N_26184,N_24736,N_25546);
and U26185 (N_26185,N_24664,N_24334);
or U26186 (N_26186,N_25498,N_24042);
xnor U26187 (N_26187,N_24370,N_24257);
and U26188 (N_26188,N_25185,N_25942);
nand U26189 (N_26189,N_24859,N_24790);
nor U26190 (N_26190,N_24731,N_25071);
nor U26191 (N_26191,N_25014,N_25389);
nand U26192 (N_26192,N_25027,N_24552);
xor U26193 (N_26193,N_24829,N_24869);
xnor U26194 (N_26194,N_25831,N_24142);
nor U26195 (N_26195,N_24173,N_24968);
and U26196 (N_26196,N_24283,N_24015);
nand U26197 (N_26197,N_25001,N_25476);
nand U26198 (N_26198,N_25689,N_24429);
or U26199 (N_26199,N_24269,N_25133);
or U26200 (N_26200,N_24657,N_24823);
nor U26201 (N_26201,N_24550,N_24708);
nand U26202 (N_26202,N_24591,N_24408);
xnor U26203 (N_26203,N_25453,N_25812);
nor U26204 (N_26204,N_25467,N_24595);
nand U26205 (N_26205,N_24616,N_25265);
or U26206 (N_26206,N_24394,N_24709);
nor U26207 (N_26207,N_25935,N_25806);
xnor U26208 (N_26208,N_25850,N_25363);
nor U26209 (N_26209,N_24200,N_25008);
or U26210 (N_26210,N_25863,N_24445);
or U26211 (N_26211,N_24809,N_25464);
nand U26212 (N_26212,N_24656,N_25189);
nand U26213 (N_26213,N_25360,N_24284);
nand U26214 (N_26214,N_25552,N_24400);
or U26215 (N_26215,N_24391,N_24066);
and U26216 (N_26216,N_24264,N_25004);
nand U26217 (N_26217,N_25593,N_24083);
or U26218 (N_26218,N_24835,N_25245);
and U26219 (N_26219,N_25261,N_24153);
xor U26220 (N_26220,N_24696,N_25522);
and U26221 (N_26221,N_24584,N_24039);
or U26222 (N_26222,N_24193,N_24626);
or U26223 (N_26223,N_25561,N_25819);
nor U26224 (N_26224,N_24020,N_24381);
and U26225 (N_26225,N_24855,N_25224);
and U26226 (N_26226,N_24638,N_24905);
nor U26227 (N_26227,N_24004,N_24672);
or U26228 (N_26228,N_24301,N_25832);
or U26229 (N_26229,N_24983,N_24151);
or U26230 (N_26230,N_25460,N_25961);
nor U26231 (N_26231,N_25443,N_24767);
nor U26232 (N_26232,N_24236,N_24190);
nor U26233 (N_26233,N_25636,N_25975);
nor U26234 (N_26234,N_24288,N_24123);
or U26235 (N_26235,N_24681,N_24270);
nor U26236 (N_26236,N_25953,N_24961);
nor U26237 (N_26237,N_25392,N_25720);
or U26238 (N_26238,N_25037,N_25250);
and U26239 (N_26239,N_24650,N_24462);
xor U26240 (N_26240,N_24761,N_25137);
and U26241 (N_26241,N_25487,N_25164);
and U26242 (N_26242,N_24987,N_24204);
xor U26243 (N_26243,N_25064,N_24390);
or U26244 (N_26244,N_24505,N_25817);
xnor U26245 (N_26245,N_24309,N_24077);
xor U26246 (N_26246,N_25672,N_25616);
nand U26247 (N_26247,N_24586,N_24800);
and U26248 (N_26248,N_24435,N_24486);
and U26249 (N_26249,N_25477,N_25586);
or U26250 (N_26250,N_25969,N_25548);
nor U26251 (N_26251,N_25335,N_24493);
nor U26252 (N_26252,N_25406,N_24824);
and U26253 (N_26253,N_24147,N_25328);
nor U26254 (N_26254,N_24841,N_25229);
xnor U26255 (N_26255,N_24074,N_25753);
or U26256 (N_26256,N_25524,N_24973);
xor U26257 (N_26257,N_24819,N_24199);
and U26258 (N_26258,N_24251,N_25254);
xor U26259 (N_26259,N_25326,N_24827);
and U26260 (N_26260,N_25926,N_24555);
and U26261 (N_26261,N_25275,N_24069);
nand U26262 (N_26262,N_24145,N_24679);
nand U26263 (N_26263,N_25489,N_24563);
and U26264 (N_26264,N_24935,N_24470);
nor U26265 (N_26265,N_24665,N_24768);
nor U26266 (N_26266,N_24250,N_24821);
or U26267 (N_26267,N_25838,N_24113);
or U26268 (N_26268,N_25502,N_24500);
xnor U26269 (N_26269,N_24302,N_24793);
or U26270 (N_26270,N_24440,N_24325);
xnor U26271 (N_26271,N_25717,N_24180);
or U26272 (N_26272,N_25143,N_24222);
or U26273 (N_26273,N_25852,N_24384);
nor U26274 (N_26274,N_24556,N_24095);
or U26275 (N_26275,N_24268,N_24691);
nand U26276 (N_26276,N_25747,N_25827);
xnor U26277 (N_26277,N_24643,N_24538);
or U26278 (N_26278,N_24852,N_24070);
nor U26279 (N_26279,N_24277,N_24870);
xor U26280 (N_26280,N_24707,N_25021);
nor U26281 (N_26281,N_25065,N_25134);
and U26282 (N_26282,N_24763,N_24569);
and U26283 (N_26283,N_25757,N_25317);
and U26284 (N_26284,N_24249,N_24728);
or U26285 (N_26285,N_25103,N_24774);
nand U26286 (N_26286,N_24553,N_25769);
nand U26287 (N_26287,N_24863,N_25078);
or U26288 (N_26288,N_24380,N_24904);
and U26289 (N_26289,N_24964,N_24451);
xnor U26290 (N_26290,N_25194,N_25718);
nor U26291 (N_26291,N_24896,N_24531);
and U26292 (N_26292,N_24911,N_25036);
nand U26293 (N_26293,N_24851,N_25086);
nand U26294 (N_26294,N_24788,N_24254);
nand U26295 (N_26295,N_25878,N_24727);
or U26296 (N_26296,N_25298,N_25728);
and U26297 (N_26297,N_25764,N_25399);
and U26298 (N_26298,N_24029,N_25022);
nand U26299 (N_26299,N_25835,N_24612);
nand U26300 (N_26300,N_25284,N_25127);
nand U26301 (N_26301,N_24661,N_24701);
and U26302 (N_26302,N_25876,N_24395);
and U26303 (N_26303,N_24738,N_25101);
or U26304 (N_26304,N_24733,N_25856);
nand U26305 (N_26305,N_24956,N_25619);
nand U26306 (N_26306,N_25272,N_24700);
xor U26307 (N_26307,N_24963,N_25923);
and U26308 (N_26308,N_25699,N_24689);
and U26309 (N_26309,N_24355,N_24933);
and U26310 (N_26310,N_25114,N_24232);
xnor U26311 (N_26311,N_25765,N_24234);
nand U26312 (N_26312,N_24106,N_24036);
nand U26313 (N_26313,N_25925,N_25631);
nand U26314 (N_26314,N_25493,N_25353);
nand U26315 (N_26315,N_25366,N_24131);
nor U26316 (N_26316,N_25735,N_24651);
xnor U26317 (N_26317,N_24051,N_25039);
xor U26318 (N_26318,N_25073,N_25420);
xnor U26319 (N_26319,N_25368,N_24125);
xnor U26320 (N_26320,N_25800,N_25528);
nor U26321 (N_26321,N_25580,N_24465);
nor U26322 (N_26322,N_25499,N_24385);
nand U26323 (N_26323,N_24014,N_24634);
or U26324 (N_26324,N_25273,N_25048);
xor U26325 (N_26325,N_25599,N_25824);
and U26326 (N_26326,N_24217,N_24785);
or U26327 (N_26327,N_24687,N_25560);
or U26328 (N_26328,N_24677,N_24923);
xnor U26329 (N_26329,N_25523,N_25803);
nand U26330 (N_26330,N_25783,N_25780);
or U26331 (N_26331,N_24022,N_24834);
or U26332 (N_26332,N_24529,N_24318);
nand U26333 (N_26333,N_24105,N_24313);
nor U26334 (N_26334,N_25940,N_25996);
nor U26335 (N_26335,N_24715,N_25080);
nand U26336 (N_26336,N_25763,N_25240);
and U26337 (N_26337,N_24406,N_24063);
or U26338 (N_26338,N_25538,N_24343);
nand U26339 (N_26339,N_24917,N_25211);
nor U26340 (N_26340,N_25517,N_24849);
or U26341 (N_26341,N_25052,N_25395);
xor U26342 (N_26342,N_24187,N_24446);
nand U26343 (N_26343,N_24787,N_24437);
or U26344 (N_26344,N_25733,N_24000);
nor U26345 (N_26345,N_25930,N_24702);
nand U26346 (N_26346,N_25452,N_25697);
nor U26347 (N_26347,N_25837,N_25215);
or U26348 (N_26348,N_24161,N_25286);
xnor U26349 (N_26349,N_25973,N_24166);
nand U26350 (N_26350,N_24698,N_25836);
nand U26351 (N_26351,N_24980,N_25247);
nor U26352 (N_26352,N_24363,N_24179);
nor U26353 (N_26353,N_25300,N_24867);
or U26354 (N_26354,N_25784,N_24646);
or U26355 (N_26355,N_24667,N_24958);
nor U26356 (N_26356,N_24438,N_25350);
nor U26357 (N_26357,N_24959,N_25627);
nand U26358 (N_26358,N_25144,N_25122);
or U26359 (N_26359,N_25290,N_24564);
nand U26360 (N_26360,N_24262,N_25315);
nor U26361 (N_26361,N_25933,N_25241);
nor U26362 (N_26362,N_25795,N_25521);
nand U26363 (N_26363,N_25174,N_24220);
and U26364 (N_26364,N_25081,N_25238);
nand U26365 (N_26365,N_24600,N_25960);
nor U26366 (N_26366,N_25040,N_24862);
and U26367 (N_26367,N_25518,N_24992);
nand U26368 (N_26368,N_25025,N_24158);
or U26369 (N_26369,N_25168,N_24002);
xor U26370 (N_26370,N_25232,N_24271);
or U26371 (N_26371,N_24176,N_25472);
xnor U26372 (N_26372,N_24540,N_25543);
or U26373 (N_26373,N_24868,N_24508);
and U26374 (N_26374,N_25292,N_25677);
nand U26375 (N_26375,N_25358,N_25128);
or U26376 (N_26376,N_25670,N_25056);
and U26377 (N_26377,N_25270,N_25741);
nor U26378 (N_26378,N_24452,N_25768);
and U26379 (N_26379,N_24719,N_24246);
xor U26380 (N_26380,N_24632,N_24459);
xnor U26381 (N_26381,N_25280,N_24280);
nand U26382 (N_26382,N_24292,N_24845);
or U26383 (N_26383,N_24875,N_25378);
and U26384 (N_26384,N_24954,N_25857);
and U26385 (N_26385,N_24660,N_24114);
and U26386 (N_26386,N_25660,N_25949);
nor U26387 (N_26387,N_24978,N_24025);
xor U26388 (N_26388,N_24475,N_24676);
xnor U26389 (N_26389,N_24879,N_24759);
or U26390 (N_26390,N_25051,N_24340);
xnor U26391 (N_26391,N_25253,N_24921);
nor U26392 (N_26392,N_25515,N_24416);
xnor U26393 (N_26393,N_24535,N_25554);
and U26394 (N_26394,N_25751,N_24775);
or U26395 (N_26395,N_25028,N_25438);
nand U26396 (N_26396,N_25600,N_25562);
xor U26397 (N_26397,N_24641,N_25323);
nand U26398 (N_26398,N_25816,N_25703);
or U26399 (N_26399,N_24710,N_24820);
nor U26400 (N_26400,N_25109,N_25711);
and U26401 (N_26401,N_24185,N_25694);
and U26402 (N_26402,N_24137,N_25906);
and U26403 (N_26403,N_24388,N_25919);
nand U26404 (N_26404,N_24135,N_25948);
nor U26405 (N_26405,N_25167,N_25687);
nor U26406 (N_26406,N_24295,N_24747);
nor U26407 (N_26407,N_24216,N_24315);
or U26408 (N_26408,N_24386,N_24304);
or U26409 (N_26409,N_25605,N_24048);
or U26410 (N_26410,N_25564,N_24327);
nor U26411 (N_26411,N_24865,N_25216);
nor U26412 (N_26412,N_25195,N_25620);
nor U26413 (N_26413,N_24119,N_25611);
nand U26414 (N_26414,N_25306,N_24703);
and U26415 (N_26415,N_24975,N_24514);
nand U26416 (N_26416,N_25644,N_25166);
xor U26417 (N_26417,N_24188,N_24996);
nor U26418 (N_26418,N_25277,N_24796);
nand U26419 (N_26419,N_25204,N_24950);
xnor U26420 (N_26420,N_24047,N_24558);
nor U26421 (N_26421,N_24516,N_25266);
and U26422 (N_26422,N_24494,N_24848);
xnor U26423 (N_26423,N_24285,N_25375);
and U26424 (N_26424,N_25150,N_25007);
xor U26425 (N_26425,N_25551,N_24919);
and U26426 (N_26426,N_25159,N_25312);
or U26427 (N_26427,N_25050,N_25967);
nand U26428 (N_26428,N_24619,N_25754);
and U26429 (N_26429,N_24024,N_24323);
xnor U26430 (N_26430,N_25814,N_25176);
nor U26431 (N_26431,N_25479,N_24878);
and U26432 (N_26432,N_24524,N_25356);
nand U26433 (N_26433,N_24644,N_24697);
xnor U26434 (N_26434,N_25952,N_25739);
and U26435 (N_26435,N_25278,N_24802);
and U26436 (N_26436,N_24912,N_24723);
nand U26437 (N_26437,N_24265,N_25519);
and U26438 (N_26438,N_25845,N_24120);
nor U26439 (N_26439,N_25681,N_25539);
and U26440 (N_26440,N_24521,N_25771);
or U26441 (N_26441,N_25448,N_24913);
and U26442 (N_26442,N_24925,N_24207);
and U26443 (N_26443,N_24392,N_24637);
nor U26444 (N_26444,N_25209,N_25716);
and U26445 (N_26445,N_24282,N_25839);
nor U26446 (N_26446,N_25896,N_25658);
nor U26447 (N_26447,N_25330,N_24447);
xor U26448 (N_26448,N_25465,N_24492);
nand U26449 (N_26449,N_25742,N_25778);
nor U26450 (N_26450,N_24129,N_24085);
or U26451 (N_26451,N_24916,N_24530);
and U26452 (N_26452,N_24476,N_25609);
and U26453 (N_26453,N_24333,N_24762);
xnor U26454 (N_26454,N_24673,N_25369);
nor U26455 (N_26455,N_25820,N_25513);
nand U26456 (N_26456,N_25070,N_25401);
and U26457 (N_26457,N_25640,N_24208);
or U26458 (N_26458,N_25662,N_24920);
nand U26459 (N_26459,N_25459,N_24377);
nor U26460 (N_26460,N_24559,N_24724);
nor U26461 (N_26461,N_25904,N_25032);
and U26462 (N_26462,N_25511,N_25865);
nand U26463 (N_26463,N_25096,N_25713);
and U26464 (N_26464,N_25442,N_24133);
or U26465 (N_26465,N_24136,N_25701);
nor U26466 (N_26466,N_25289,N_24016);
or U26467 (N_26467,N_25107,N_24549);
or U26468 (N_26468,N_24658,N_25927);
xnor U26469 (N_26469,N_24021,N_25413);
nor U26470 (N_26470,N_24630,N_25160);
nand U26471 (N_26471,N_25384,N_25393);
and U26472 (N_26472,N_24589,N_24290);
nor U26473 (N_26473,N_25509,N_24744);
and U26474 (N_26474,N_24003,N_24779);
nor U26475 (N_26475,N_24560,N_25019);
and U26476 (N_26476,N_24401,N_25678);
nor U26477 (N_26477,N_25762,N_24596);
xnor U26478 (N_26478,N_24897,N_25002);
xnor U26479 (N_26479,N_24140,N_24082);
xor U26480 (N_26480,N_25738,N_25468);
nand U26481 (N_26481,N_24888,N_24839);
or U26482 (N_26482,N_25362,N_25607);
nor U26483 (N_26483,N_24986,N_25540);
and U26484 (N_26484,N_25291,N_25598);
nand U26485 (N_26485,N_24393,N_25202);
nor U26486 (N_26486,N_25474,N_25005);
nand U26487 (N_26487,N_25484,N_25336);
xor U26488 (N_26488,N_24734,N_24491);
or U26489 (N_26489,N_25258,N_25233);
xor U26490 (N_26490,N_25939,N_24041);
and U26491 (N_26491,N_24803,N_25759);
xnor U26492 (N_26492,N_24756,N_25642);
nor U26493 (N_26493,N_24629,N_24455);
nor U26494 (N_26494,N_25297,N_24669);
xor U26495 (N_26495,N_24079,N_24057);
or U26496 (N_26496,N_24485,N_24339);
nor U26497 (N_26497,N_25201,N_24627);
and U26498 (N_26498,N_24575,N_24523);
or U26499 (N_26499,N_25536,N_24548);
xnor U26500 (N_26500,N_25921,N_24981);
xnor U26501 (N_26501,N_24346,N_25579);
and U26502 (N_26502,N_25976,N_24354);
and U26503 (N_26503,N_25862,N_25997);
xnor U26504 (N_26504,N_24321,N_25938);
nor U26505 (N_26505,N_25394,N_25525);
nor U26506 (N_26506,N_24011,N_24527);
nand U26507 (N_26507,N_24229,N_25646);
xor U26508 (N_26508,N_24947,N_25641);
and U26509 (N_26509,N_24458,N_24441);
or U26510 (N_26510,N_25628,N_25179);
nand U26511 (N_26511,N_25748,N_24850);
nand U26512 (N_26512,N_24297,N_24368);
and U26513 (N_26513,N_25775,N_24434);
xor U26514 (N_26514,N_25281,N_24252);
and U26515 (N_26515,N_25325,N_24607);
nand U26516 (N_26516,N_25945,N_24960);
nor U26517 (N_26517,N_25155,N_25494);
nor U26518 (N_26518,N_24449,N_24511);
nand U26519 (N_26519,N_25985,N_25505);
and U26520 (N_26520,N_24432,N_25573);
nand U26521 (N_26521,N_25592,N_25843);
or U26522 (N_26522,N_24407,N_25299);
nor U26523 (N_26523,N_25603,N_25138);
or U26524 (N_26524,N_25192,N_25486);
and U26525 (N_26525,N_25296,N_25316);
nand U26526 (N_26526,N_24286,N_24836);
or U26527 (N_26527,N_25033,N_24404);
nand U26528 (N_26528,N_24050,N_24861);
and U26529 (N_26529,N_24134,N_25475);
or U26530 (N_26530,N_25231,N_24097);
or U26531 (N_26531,N_25478,N_25018);
and U26532 (N_26532,N_25698,N_25987);
and U26533 (N_26533,N_24930,N_24609);
nor U26534 (N_26534,N_25941,N_24054);
xor U26535 (N_26535,N_24688,N_25991);
nor U26536 (N_26536,N_25541,N_25099);
nor U26537 (N_26537,N_25601,N_24148);
and U26538 (N_26538,N_24633,N_24413);
xor U26539 (N_26539,N_24562,N_25327);
nor U26540 (N_26540,N_25026,N_25587);
nand U26541 (N_26541,N_25809,N_24005);
nand U26542 (N_26542,N_25430,N_24122);
or U26543 (N_26543,N_25485,N_25062);
xor U26544 (N_26544,N_24326,N_25613);
xnor U26545 (N_26545,N_25929,N_25995);
nand U26546 (N_26546,N_24593,N_24273);
and U26547 (N_26547,N_24001,N_25132);
xnor U26548 (N_26548,N_24623,N_24214);
nor U26549 (N_26549,N_24805,N_24197);
or U26550 (N_26550,N_25950,N_25696);
nand U26551 (N_26551,N_25106,N_24317);
or U26552 (N_26552,N_24291,N_24565);
xnor U26553 (N_26553,N_24034,N_25886);
and U26554 (N_26554,N_24705,N_24830);
and U26555 (N_26555,N_25686,N_25283);
nand U26556 (N_26556,N_24171,N_25329);
xnor U26557 (N_26557,N_25861,N_25104);
or U26558 (N_26558,N_24857,N_25175);
nand U26559 (N_26559,N_25879,N_25003);
nand U26560 (N_26560,N_24342,N_25706);
and U26561 (N_26561,N_25668,N_24010);
xor U26562 (N_26562,N_25408,N_24583);
nand U26563 (N_26563,N_25617,N_24794);
and U26564 (N_26564,N_25226,N_24107);
nor U26565 (N_26565,N_24692,N_25994);
xor U26566 (N_26566,N_24915,N_25181);
and U26567 (N_26567,N_25649,N_25789);
or U26568 (N_26568,N_24052,N_25285);
and U26569 (N_26569,N_25090,N_25414);
and U26570 (N_26570,N_25197,N_25152);
or U26571 (N_26571,N_24818,N_25855);
nor U26572 (N_26572,N_24864,N_24328);
nand U26573 (N_26573,N_24668,N_24781);
nor U26574 (N_26574,N_25993,N_25038);
or U26575 (N_26575,N_24614,N_24484);
or U26576 (N_26576,N_25432,N_25555);
xor U26577 (N_26577,N_24032,N_25131);
and U26578 (N_26578,N_25891,N_24443);
and U26579 (N_26579,N_25665,N_25410);
xnor U26580 (N_26580,N_24792,N_25239);
nand U26581 (N_26581,N_25912,N_24038);
nand U26582 (N_26582,N_24467,N_24928);
nor U26583 (N_26583,N_24319,N_25915);
and U26584 (N_26584,N_25264,N_25041);
xor U26585 (N_26585,N_25077,N_25801);
nor U26586 (N_26586,N_25884,N_25563);
xor U26587 (N_26587,N_24056,N_25371);
and U26588 (N_26588,N_25901,N_24320);
and U26589 (N_26589,N_25402,N_25859);
nand U26590 (N_26590,N_24100,N_24716);
xnor U26591 (N_26591,N_24495,N_24152);
and U26592 (N_26592,N_25851,N_24725);
nor U26593 (N_26593,N_25165,N_24080);
and U26594 (N_26594,N_25571,N_25497);
and U26595 (N_26595,N_25146,N_24090);
xor U26596 (N_26596,N_24908,N_24833);
or U26597 (N_26597,N_25177,N_24985);
or U26598 (N_26598,N_25818,N_25977);
and U26599 (N_26599,N_24544,N_24582);
and U26600 (N_26600,N_25412,N_24778);
nor U26601 (N_26601,N_25125,N_24410);
and U26602 (N_26602,N_25429,N_24914);
nor U26603 (N_26603,N_24810,N_25223);
nor U26604 (N_26604,N_24982,N_25981);
and U26605 (N_26605,N_24376,N_25761);
nor U26606 (N_26606,N_25576,N_25508);
and U26607 (N_26607,N_25840,N_24431);
and U26608 (N_26608,N_24089,N_24415);
nor U26609 (N_26609,N_25999,N_24932);
nand U26610 (N_26610,N_25492,N_24566);
nor U26611 (N_26611,N_24713,N_24737);
xnor U26612 (N_26612,N_24350,N_24979);
nand U26613 (N_26613,N_25643,N_25813);
and U26614 (N_26614,N_25868,N_25404);
nand U26615 (N_26615,N_24356,N_25473);
nor U26616 (N_26616,N_25959,N_24590);
or U26617 (N_26617,N_24403,N_24167);
nand U26618 (N_26618,N_25897,N_24382);
nor U26619 (N_26619,N_25190,N_25972);
nor U26620 (N_26620,N_24138,N_25989);
and U26621 (N_26621,N_25147,N_25918);
nor U26622 (N_26622,N_24588,N_25349);
xor U26623 (N_26623,N_24067,N_24186);
or U26624 (N_26624,N_24922,N_24091);
nand U26625 (N_26625,N_25500,N_25710);
or U26626 (N_26626,N_25724,N_25269);
nand U26627 (N_26627,N_24017,N_25792);
or U26628 (N_26628,N_24275,N_24243);
xnor U26629 (N_26629,N_25829,N_25683);
and U26630 (N_26630,N_24012,N_25974);
nand U26631 (N_26631,N_24398,N_25680);
or U26632 (N_26632,N_25913,N_24178);
and U26633 (N_26633,N_24159,N_24966);
or U26634 (N_26634,N_25988,N_24533);
nor U26635 (N_26635,N_24081,N_25889);
xor U26636 (N_26636,N_25970,N_25200);
xnor U26637 (N_26637,N_24055,N_25373);
and U26638 (N_26638,N_25931,N_24610);
nor U26639 (N_26639,N_24906,N_24481);
nor U26640 (N_26640,N_25379,N_25512);
nand U26641 (N_26641,N_25495,N_25732);
nor U26642 (N_26642,N_24647,N_25095);
and U26643 (N_26643,N_25529,N_24260);
or U26644 (N_26644,N_24513,N_25808);
or U26645 (N_26645,N_25111,N_25595);
or U26646 (N_26646,N_24194,N_25340);
xor U26647 (N_26647,N_25567,N_24156);
and U26648 (N_26648,N_24402,N_24640);
and U26649 (N_26649,N_25075,N_25449);
nand U26650 (N_26650,N_25655,N_25920);
nor U26651 (N_26651,N_25965,N_25017);
and U26652 (N_26652,N_24366,N_24387);
nor U26653 (N_26653,N_25569,N_24239);
nand U26654 (N_26654,N_24347,N_24418);
nand U26655 (N_26655,N_24299,N_25400);
nor U26656 (N_26656,N_25156,N_24750);
nor U26657 (N_26657,N_25719,N_25902);
nand U26658 (N_26658,N_24477,N_24576);
nand U26659 (N_26659,N_24433,N_24483);
xor U26660 (N_26660,N_25042,N_25259);
nor U26661 (N_26661,N_25435,N_24345);
nor U26662 (N_26662,N_25034,N_24571);
and U26663 (N_26663,N_25205,N_24424);
and U26664 (N_26664,N_25203,N_25208);
or U26665 (N_26665,N_24938,N_24371);
or U26666 (N_26666,N_25964,N_25744);
nor U26667 (N_26667,N_25118,N_24224);
xor U26668 (N_26668,N_24329,N_25957);
and U26669 (N_26669,N_24989,N_25345);
nand U26670 (N_26670,N_24976,N_24215);
xor U26671 (N_26671,N_25116,N_25610);
or U26672 (N_26672,N_24464,N_25691);
nand U26673 (N_26673,N_25333,N_25574);
xor U26674 (N_26674,N_24999,N_25196);
nor U26675 (N_26675,N_25621,N_24872);
or U26676 (N_26676,N_24007,N_25934);
xnor U26677 (N_26677,N_25516,N_24498);
and U26678 (N_26678,N_24682,N_25346);
nand U26679 (N_26679,N_25207,N_25866);
or U26680 (N_26680,N_24936,N_25575);
nor U26681 (N_26681,N_25365,N_25321);
or U26682 (N_26682,N_24873,N_25947);
or U26683 (N_26683,N_24061,N_25161);
nand U26684 (N_26684,N_24499,N_24324);
and U26685 (N_26685,N_25230,N_25469);
xor U26686 (N_26686,N_24071,N_24684);
and U26687 (N_26687,N_24174,N_24279);
and U26688 (N_26688,N_24412,N_25268);
nand U26689 (N_26689,N_25907,N_25594);
xor U26690 (N_26690,N_24683,N_24815);
and U26691 (N_26691,N_24263,N_25332);
or U26692 (N_26692,N_24205,N_24102);
or U26693 (N_26693,N_25674,N_25083);
nor U26694 (N_26694,N_25110,N_24546);
or U26695 (N_26695,N_24227,N_24813);
nor U26696 (N_26696,N_25984,N_24532);
xor U26697 (N_26697,N_25794,N_24512);
and U26698 (N_26698,N_24096,N_25428);
nand U26699 (N_26699,N_25178,N_25248);
and U26700 (N_26700,N_25731,N_24117);
nor U26701 (N_26701,N_24237,N_25113);
and U26702 (N_26702,N_25186,N_25145);
nor U26703 (N_26703,N_25553,N_25679);
nor U26704 (N_26704,N_25639,N_24752);
nor U26705 (N_26705,N_24510,N_24109);
xnor U26706 (N_26706,N_24362,N_25917);
xnor U26707 (N_26707,N_24615,N_24770);
nand U26708 (N_26708,N_25024,N_25348);
and U26709 (N_26709,N_24901,N_24843);
or U26710 (N_26710,N_24974,N_24536);
xnor U26711 (N_26711,N_24115,N_25854);
nor U26712 (N_26712,N_25169,N_25225);
nand U26713 (N_26713,N_24502,N_25188);
xor U26714 (N_26714,N_25797,N_25094);
nor U26715 (N_26715,N_24749,N_25962);
or U26716 (N_26716,N_24396,N_24195);
nor U26717 (N_26717,N_24389,N_25235);
nor U26718 (N_26718,N_24635,N_24247);
nor U26719 (N_26719,N_25445,N_24602);
nor U26720 (N_26720,N_24984,N_25864);
xor U26721 (N_26721,N_24143,N_24726);
or U26722 (N_26722,N_25992,N_25978);
nand U26723 (N_26723,N_25826,N_25444);
or U26724 (N_26724,N_24450,N_24141);
and U26725 (N_26725,N_24478,N_24625);
nor U26726 (N_26726,N_25262,N_25387);
or U26727 (N_26727,N_24675,N_25102);
xnor U26728 (N_26728,N_24812,N_24192);
xor U26729 (N_26729,N_25584,N_24519);
xnor U26730 (N_26730,N_25249,N_25785);
xor U26731 (N_26731,N_25446,N_25834);
or U26732 (N_26732,N_24155,N_24298);
nor U26733 (N_26733,N_25431,N_25210);
nor U26734 (N_26734,N_24338,N_25671);
nand U26735 (N_26735,N_24653,N_25370);
nor U26736 (N_26736,N_24828,N_25422);
and U26737 (N_26737,N_25180,N_25121);
nand U26738 (N_26738,N_25046,N_24212);
and U26739 (N_26739,N_24655,N_25274);
and U26740 (N_26740,N_25514,N_25342);
or U26741 (N_26741,N_25585,N_25436);
nand U26742 (N_26742,N_24344,N_25488);
xnor U26743 (N_26743,N_24177,N_24303);
and U26744 (N_26744,N_24111,N_24294);
and U26745 (N_26745,N_25058,N_24101);
nor U26746 (N_26746,N_24613,N_24776);
and U26747 (N_26747,N_25533,N_25869);
and U26748 (N_26748,N_25663,N_25578);
nand U26749 (N_26749,N_25383,N_24030);
nand U26750 (N_26750,N_25909,N_24358);
nor U26751 (N_26751,N_25388,N_24754);
and U26752 (N_26752,N_25398,N_25305);
nor U26753 (N_26753,N_25588,N_25364);
nor U26754 (N_26754,N_25085,N_24988);
xor U26755 (N_26755,N_25928,N_25684);
and U26756 (N_26756,N_25082,N_25804);
nand U26757 (N_26757,N_25490,N_25295);
nor U26758 (N_26758,N_25661,N_24088);
or U26759 (N_26759,N_25900,N_24420);
nand U26760 (N_26760,N_24608,N_25221);
or U26761 (N_26761,N_25276,N_25871);
xor U26762 (N_26762,N_25946,N_25311);
xor U26763 (N_26763,N_24645,N_25781);
and U26764 (N_26764,N_24674,N_25466);
or U26765 (N_26765,N_24076,N_25860);
or U26766 (N_26766,N_25214,N_25898);
xnor U26767 (N_26767,N_25227,N_25481);
xnor U26768 (N_26768,N_24466,N_25409);
xor U26769 (N_26769,N_24649,N_25632);
xnor U26770 (N_26770,N_25779,N_25885);
xor U26771 (N_26771,N_25916,N_24685);
or U26772 (N_26772,N_24267,N_25526);
xor U26773 (N_26773,N_25287,N_24154);
nor U26774 (N_26774,N_24515,N_24757);
xnor U26775 (N_26775,N_24993,N_24695);
nor U26776 (N_26776,N_24570,N_25653);
xor U26777 (N_26777,N_24720,N_25652);
xnor U26778 (N_26778,N_25787,N_24739);
nand U26779 (N_26779,N_25685,N_25377);
or U26780 (N_26780,N_24501,N_25031);
nand U26781 (N_26781,N_25633,N_25704);
xor U26782 (N_26782,N_24128,N_25583);
nor U26783 (N_26783,N_24889,N_25648);
and U26784 (N_26784,N_25089,N_24168);
nor U26785 (N_26785,N_25841,N_24970);
and U26786 (N_26786,N_25163,N_25612);
or U26787 (N_26787,N_25637,N_25914);
nand U26788 (N_26788,N_24804,N_24740);
or U26789 (N_26789,N_25782,N_25530);
nand U26790 (N_26790,N_25098,N_25591);
xor U26791 (N_26791,N_25117,N_24336);
nor U26792 (N_26792,N_24027,N_24139);
nand U26793 (N_26793,N_25074,N_24127);
and U26794 (N_26794,N_25173,N_25572);
or U26795 (N_26795,N_24712,N_24817);
or U26796 (N_26796,N_24411,N_24456);
and U26797 (N_26797,N_25411,N_24854);
nor U26798 (N_26798,N_24718,N_25183);
and U26799 (N_26799,N_24086,N_24231);
or U26800 (N_26800,N_24621,N_24620);
and U26801 (N_26801,N_25361,N_25700);
and U26802 (N_26802,N_25545,N_24314);
nor U26803 (N_26803,N_25963,N_25549);
or U26804 (N_26804,N_25966,N_25892);
and U26805 (N_26805,N_24816,N_25372);
or U26806 (N_26806,N_25043,N_24359);
xnor U26807 (N_26807,N_24043,N_24853);
xnor U26808 (N_26808,N_24663,N_24893);
xor U26809 (N_26809,N_24955,N_24092);
nand U26810 (N_26810,N_24670,N_24648);
or U26811 (N_26811,N_24425,N_24068);
xor U26812 (N_26812,N_25112,N_25656);
and U26813 (N_26813,N_25120,N_24847);
nand U26814 (N_26814,N_24448,N_25220);
or U26815 (N_26815,N_25419,N_25821);
xnor U26816 (N_26816,N_24579,N_24977);
or U26817 (N_26817,N_25496,N_25149);
nor U26818 (N_26818,N_24430,N_24525);
xnor U26819 (N_26819,N_24693,N_25352);
xor U26820 (N_26820,N_24040,N_24316);
and U26821 (N_26821,N_24831,N_24926);
nor U26822 (N_26822,N_25457,N_24149);
nor U26823 (N_26823,N_24104,N_24542);
nand U26824 (N_26824,N_24245,N_24840);
nor U26825 (N_26825,N_24078,N_24019);
xor U26826 (N_26826,N_24365,N_24545);
xnor U26827 (N_26827,N_24399,N_24858);
and U26828 (N_26828,N_25796,N_25954);
nand U26829 (N_26829,N_25558,N_24160);
nor U26830 (N_26830,N_25602,N_24124);
nor U26831 (N_26831,N_25338,N_25924);
nor U26832 (N_26832,N_25076,N_24013);
nand U26833 (N_26833,N_24244,N_24348);
nand U26834 (N_26834,N_25666,N_24551);
or U26835 (N_26835,N_25302,N_24103);
nand U26836 (N_26836,N_25905,N_25427);
or U26837 (N_26837,N_25148,N_24423);
nor U26838 (N_26838,N_24226,N_25324);
xor U26839 (N_26839,N_24732,N_24760);
and U26840 (N_26840,N_24554,N_24866);
xnor U26841 (N_26841,N_25881,N_24379);
nand U26842 (N_26842,N_24887,N_25347);
and U26843 (N_26843,N_24150,N_25309);
or U26844 (N_26844,N_25482,N_25667);
xnor U26845 (N_26845,N_24585,N_25307);
or U26846 (N_26846,N_25029,N_24856);
xnor U26847 (N_26847,N_25708,N_25458);
or U26848 (N_26848,N_25774,N_25433);
nor U26849 (N_26849,N_24006,N_24624);
nor U26850 (N_26850,N_24844,N_24957);
nor U26851 (N_26851,N_24235,N_24473);
nor U26852 (N_26852,N_25199,N_24837);
xor U26853 (N_26853,N_25932,N_25887);
nand U26854 (N_26854,N_25638,N_25714);
nand U26855 (N_26855,N_25581,N_25390);
or U26856 (N_26856,N_24652,N_25842);
or U26857 (N_26857,N_25244,N_25318);
nand U26858 (N_26858,N_24671,N_24937);
nor U26859 (N_26859,N_25105,N_25123);
nand U26860 (N_26860,N_25874,N_24782);
nor U26861 (N_26861,N_24098,N_24780);
or U26862 (N_26862,N_24018,N_25943);
nor U26863 (N_26863,N_24945,N_25630);
or U26864 (N_26864,N_25527,N_25091);
and U26865 (N_26865,N_24578,N_25450);
xnor U26866 (N_26866,N_24378,N_24765);
and U26867 (N_26867,N_25848,N_24939);
or U26868 (N_26868,N_25060,N_24053);
nand U26869 (N_26869,N_25491,N_25669);
and U26870 (N_26870,N_24825,N_24482);
nor U26871 (N_26871,N_24241,N_25381);
nor U26872 (N_26872,N_25986,N_25847);
nor U26873 (N_26873,N_25126,N_25767);
or U26874 (N_26874,N_25568,N_25441);
nand U26875 (N_26875,N_25745,N_24934);
and U26876 (N_26876,N_24686,N_24058);
xor U26877 (N_26877,N_24209,N_25702);
nor U26878 (N_26878,N_24704,N_25980);
or U26879 (N_26879,N_24242,N_25776);
xnor U26880 (N_26880,N_25228,N_24414);
and U26881 (N_26881,N_24454,N_25424);
or U26882 (N_26882,N_25651,N_25115);
nand U26883 (N_26883,N_25597,N_24572);
xnor U26884 (N_26884,N_24405,N_24112);
nor U26885 (N_26885,N_25625,N_25725);
nor U26886 (N_26886,N_24428,N_25727);
or U26887 (N_26887,N_24374,N_24110);
and U26888 (N_26888,N_24064,N_24994);
xor U26889 (N_26889,N_25251,N_24349);
and U26890 (N_26890,N_24093,N_25798);
or U26891 (N_26891,N_24504,N_24639);
and U26892 (N_26892,N_25439,N_24601);
or U26893 (N_26893,N_24330,N_24033);
xnor U26894 (N_26894,N_24903,N_25793);
nor U26895 (N_26895,N_24991,N_24654);
xnor U26896 (N_26896,N_24877,N_25895);
and U26897 (N_26897,N_24786,N_24417);
or U26898 (N_26898,N_24169,N_25405);
nand U26899 (N_26899,N_25520,N_24951);
nand U26900 (N_26900,N_24181,N_25635);
nor U26901 (N_26901,N_25396,N_25626);
xnor U26902 (N_26902,N_24784,N_25510);
nor U26903 (N_26903,N_24990,N_25415);
xor U26904 (N_26904,N_25063,N_25067);
and U26905 (N_26905,N_25471,N_25506);
nor U26906 (N_26906,N_24598,N_24722);
nor U26907 (N_26907,N_25049,N_25184);
xor U26908 (N_26908,N_24967,N_25359);
nor U26909 (N_26909,N_25154,N_25531);
nor U26910 (N_26910,N_24618,N_24795);
xnor U26911 (N_26911,N_25715,N_24439);
xor U26912 (N_26912,N_24574,N_25873);
nand U26913 (N_26913,N_24910,N_24832);
and U26914 (N_26914,N_25709,N_24699);
and U26915 (N_26915,N_25386,N_24372);
or U26916 (N_26916,N_24942,N_24617);
xor U26917 (N_26917,N_24157,N_25810);
nand U26918 (N_26918,N_24253,N_24706);
nand U26919 (N_26919,N_24628,N_25308);
nand U26920 (N_26920,N_25035,N_25877);
nor U26921 (N_26921,N_25606,N_25068);
xnor U26922 (N_26922,N_25971,N_24287);
and U26923 (N_26923,N_24108,N_25693);
nor U26924 (N_26924,N_25622,N_24577);
or U26925 (N_26925,N_24741,N_24885);
or U26926 (N_26926,N_25825,N_24943);
xor U26927 (N_26927,N_25888,N_24497);
or U26928 (N_26928,N_25320,N_25141);
or U26929 (N_26929,N_24422,N_25440);
and U26930 (N_26930,N_24202,N_25072);
nor U26931 (N_26931,N_25883,N_24479);
and U26932 (N_26932,N_25618,N_25206);
nor U26933 (N_26933,N_24203,N_24213);
nor U26934 (N_26934,N_25911,N_25664);
nor U26935 (N_26935,N_25009,N_25737);
nand U26936 (N_26936,N_25182,N_24461);
nor U26937 (N_26937,N_25337,N_24031);
or U26938 (N_26938,N_24311,N_24838);
nor U26939 (N_26939,N_25756,N_24274);
nor U26940 (N_26940,N_25805,N_24871);
and U26941 (N_26941,N_25828,N_25380);
nand U26942 (N_26942,N_25604,N_24789);
or U26943 (N_26943,N_24636,N_25255);
and U26944 (N_26944,N_24170,N_24929);
or U26945 (N_26945,N_24680,N_24028);
and U26946 (N_26946,N_25736,N_24886);
nor U26947 (N_26947,N_24331,N_24894);
and U26948 (N_26948,N_25135,N_25968);
and U26949 (N_26949,N_24899,N_24094);
nand U26950 (N_26950,N_24766,N_24062);
nor U26951 (N_26951,N_24509,N_24666);
nand U26952 (N_26952,N_25403,N_25846);
and U26953 (N_26953,N_25908,N_24594);
nor U26954 (N_26954,N_25172,N_24163);
nor U26955 (N_26955,N_24880,N_24175);
and U26956 (N_26956,N_24592,N_25955);
nand U26957 (N_26957,N_24891,N_25647);
nor U26958 (N_26958,N_25417,N_25242);
and U26959 (N_26959,N_25260,N_25676);
or U26960 (N_26960,N_25922,N_25565);
nor U26961 (N_26961,N_24296,N_24472);
nor U26962 (N_26962,N_24758,N_25198);
nor U26963 (N_26963,N_25257,N_24037);
xnor U26964 (N_26964,N_25614,N_24662);
xnor U26965 (N_26965,N_25982,N_24383);
nor U26966 (N_26966,N_25544,N_25463);
nor U26967 (N_26967,N_25084,N_24604);
and U26968 (N_26968,N_25815,N_25013);
nor U26969 (N_26969,N_25418,N_24969);
xor U26970 (N_26970,N_25755,N_25547);
nand U26971 (N_26971,N_24769,N_24797);
nand U26972 (N_26972,N_25462,N_25397);
or U26973 (N_26973,N_25212,N_24948);
nand U26974 (N_26974,N_25059,N_25314);
and U26975 (N_26975,N_25790,N_25740);
nand U26976 (N_26976,N_25752,N_25726);
nand U26977 (N_26977,N_25000,N_25566);
xor U26978 (N_26978,N_24116,N_25162);
nor U26979 (N_26979,N_24965,N_24972);
nand U26980 (N_26980,N_24526,N_24223);
nor U26981 (N_26981,N_24228,N_25407);
and U26982 (N_26982,N_25721,N_25823);
or U26983 (N_26983,N_25069,N_25799);
xor U26984 (N_26984,N_24603,N_24883);
nor U26985 (N_26985,N_25903,N_24335);
xnor U26986 (N_26986,N_25108,N_25222);
or U26987 (N_26987,N_24547,N_25217);
nand U26988 (N_26988,N_25705,N_24357);
nor U26989 (N_26989,N_25455,N_25087);
xnor U26990 (N_26990,N_25015,N_25391);
nor U26991 (N_26991,N_24764,N_24807);
and U26992 (N_26992,N_25376,N_24219);
xor U26993 (N_26993,N_25880,N_24469);
xor U26994 (N_26994,N_24659,N_25252);
nor U26995 (N_26995,N_25870,N_24210);
and U26996 (N_26996,N_24059,N_24008);
nor U26997 (N_26997,N_24060,N_25532);
nor U26998 (N_26998,N_24771,N_25157);
nor U26999 (N_26999,N_24489,N_25313);
nor U27000 (N_27000,N_25263,N_25609);
and U27001 (N_27001,N_24316,N_24872);
and U27002 (N_27002,N_25527,N_25053);
or U27003 (N_27003,N_24893,N_24343);
nor U27004 (N_27004,N_25688,N_24751);
xnor U27005 (N_27005,N_25282,N_24296);
and U27006 (N_27006,N_24195,N_25890);
and U27007 (N_27007,N_24218,N_24920);
nand U27008 (N_27008,N_25057,N_25564);
nor U27009 (N_27009,N_25386,N_25754);
nand U27010 (N_27010,N_25280,N_25309);
nand U27011 (N_27011,N_24773,N_24715);
nor U27012 (N_27012,N_25485,N_24844);
and U27013 (N_27013,N_24315,N_24325);
nor U27014 (N_27014,N_25526,N_24639);
xor U27015 (N_27015,N_25962,N_25463);
nand U27016 (N_27016,N_25426,N_24515);
or U27017 (N_27017,N_24488,N_24472);
or U27018 (N_27018,N_24257,N_25766);
nand U27019 (N_27019,N_24722,N_25523);
and U27020 (N_27020,N_24380,N_24001);
and U27021 (N_27021,N_24092,N_24204);
and U27022 (N_27022,N_24942,N_25111);
or U27023 (N_27023,N_25135,N_25269);
xnor U27024 (N_27024,N_24431,N_24764);
or U27025 (N_27025,N_25440,N_25817);
nor U27026 (N_27026,N_25921,N_25934);
nor U27027 (N_27027,N_25446,N_25467);
nor U27028 (N_27028,N_24033,N_25034);
or U27029 (N_27029,N_25483,N_24574);
nand U27030 (N_27030,N_25560,N_24148);
nand U27031 (N_27031,N_24247,N_25196);
nand U27032 (N_27032,N_25601,N_25291);
or U27033 (N_27033,N_24016,N_25826);
nor U27034 (N_27034,N_25294,N_25654);
or U27035 (N_27035,N_24192,N_24502);
and U27036 (N_27036,N_25696,N_25104);
nor U27037 (N_27037,N_24731,N_25285);
xnor U27038 (N_27038,N_24471,N_24562);
xor U27039 (N_27039,N_24938,N_24247);
and U27040 (N_27040,N_25989,N_25862);
or U27041 (N_27041,N_25873,N_25810);
nand U27042 (N_27042,N_25508,N_25625);
nor U27043 (N_27043,N_24271,N_25169);
nor U27044 (N_27044,N_24960,N_24986);
xor U27045 (N_27045,N_25251,N_25681);
xor U27046 (N_27046,N_24938,N_25663);
xor U27047 (N_27047,N_25125,N_24301);
or U27048 (N_27048,N_24960,N_25175);
and U27049 (N_27049,N_24633,N_24675);
or U27050 (N_27050,N_24984,N_24594);
or U27051 (N_27051,N_25162,N_24234);
nand U27052 (N_27052,N_24960,N_24756);
nand U27053 (N_27053,N_25065,N_25697);
and U27054 (N_27054,N_24897,N_24131);
nor U27055 (N_27055,N_25437,N_25650);
and U27056 (N_27056,N_25859,N_25384);
nor U27057 (N_27057,N_24168,N_24966);
and U27058 (N_27058,N_25770,N_25667);
or U27059 (N_27059,N_25691,N_25307);
xor U27060 (N_27060,N_25236,N_25357);
nand U27061 (N_27061,N_25827,N_25042);
nor U27062 (N_27062,N_24698,N_24746);
nor U27063 (N_27063,N_24162,N_24581);
nand U27064 (N_27064,N_24046,N_25276);
nand U27065 (N_27065,N_25184,N_25995);
xor U27066 (N_27066,N_24414,N_24222);
nand U27067 (N_27067,N_25974,N_24081);
xnor U27068 (N_27068,N_24132,N_25787);
xor U27069 (N_27069,N_24807,N_24061);
xor U27070 (N_27070,N_24761,N_25891);
nand U27071 (N_27071,N_25490,N_25067);
nand U27072 (N_27072,N_25892,N_24819);
nand U27073 (N_27073,N_25660,N_24600);
nor U27074 (N_27074,N_24410,N_24905);
xor U27075 (N_27075,N_25107,N_24008);
nand U27076 (N_27076,N_25717,N_25926);
nand U27077 (N_27077,N_24832,N_24096);
nor U27078 (N_27078,N_25433,N_24651);
nand U27079 (N_27079,N_25266,N_25397);
nor U27080 (N_27080,N_24321,N_25176);
nand U27081 (N_27081,N_24364,N_24204);
nand U27082 (N_27082,N_24712,N_24809);
and U27083 (N_27083,N_24844,N_24048);
and U27084 (N_27084,N_24830,N_25984);
nand U27085 (N_27085,N_25687,N_24274);
and U27086 (N_27086,N_24150,N_25523);
or U27087 (N_27087,N_24199,N_25850);
or U27088 (N_27088,N_25894,N_24258);
nand U27089 (N_27089,N_25212,N_25002);
xnor U27090 (N_27090,N_25209,N_25326);
or U27091 (N_27091,N_25161,N_25802);
or U27092 (N_27092,N_24971,N_25661);
xor U27093 (N_27093,N_24204,N_24842);
nand U27094 (N_27094,N_25699,N_25921);
nand U27095 (N_27095,N_25320,N_24869);
and U27096 (N_27096,N_25989,N_24752);
nor U27097 (N_27097,N_24405,N_24300);
and U27098 (N_27098,N_24663,N_25465);
or U27099 (N_27099,N_25347,N_25987);
nand U27100 (N_27100,N_25221,N_25139);
and U27101 (N_27101,N_24358,N_25037);
xnor U27102 (N_27102,N_24372,N_24271);
and U27103 (N_27103,N_24390,N_24064);
nor U27104 (N_27104,N_24954,N_25078);
or U27105 (N_27105,N_25686,N_25015);
or U27106 (N_27106,N_24587,N_25133);
nor U27107 (N_27107,N_25346,N_25177);
nand U27108 (N_27108,N_25813,N_25155);
nor U27109 (N_27109,N_25699,N_24374);
or U27110 (N_27110,N_25281,N_25399);
nand U27111 (N_27111,N_24524,N_25747);
xor U27112 (N_27112,N_25140,N_24232);
and U27113 (N_27113,N_25403,N_24528);
xnor U27114 (N_27114,N_24062,N_25894);
or U27115 (N_27115,N_24040,N_25971);
or U27116 (N_27116,N_24298,N_25149);
nor U27117 (N_27117,N_25767,N_25174);
nor U27118 (N_27118,N_24863,N_25220);
and U27119 (N_27119,N_24554,N_24669);
nand U27120 (N_27120,N_24979,N_25986);
xnor U27121 (N_27121,N_24162,N_25880);
xor U27122 (N_27122,N_25892,N_24668);
and U27123 (N_27123,N_24317,N_24010);
nand U27124 (N_27124,N_25012,N_24188);
xnor U27125 (N_27125,N_25340,N_24591);
xnor U27126 (N_27126,N_25365,N_25950);
xor U27127 (N_27127,N_25333,N_24282);
nor U27128 (N_27128,N_25446,N_25073);
nand U27129 (N_27129,N_25207,N_25996);
nand U27130 (N_27130,N_24416,N_24996);
nor U27131 (N_27131,N_24451,N_25118);
or U27132 (N_27132,N_24704,N_24905);
and U27133 (N_27133,N_25888,N_25356);
and U27134 (N_27134,N_25266,N_24421);
xor U27135 (N_27135,N_24640,N_25121);
and U27136 (N_27136,N_24707,N_25724);
xnor U27137 (N_27137,N_24674,N_24113);
xor U27138 (N_27138,N_24636,N_25312);
nor U27139 (N_27139,N_25106,N_24221);
and U27140 (N_27140,N_24324,N_25767);
xnor U27141 (N_27141,N_24835,N_24909);
and U27142 (N_27142,N_24905,N_24542);
xor U27143 (N_27143,N_25350,N_24458);
nor U27144 (N_27144,N_25133,N_24974);
or U27145 (N_27145,N_24399,N_24795);
and U27146 (N_27146,N_25756,N_24250);
and U27147 (N_27147,N_25813,N_24133);
nor U27148 (N_27148,N_25554,N_24862);
or U27149 (N_27149,N_25629,N_25357);
and U27150 (N_27150,N_25934,N_25617);
xnor U27151 (N_27151,N_25447,N_25150);
nand U27152 (N_27152,N_25081,N_24061);
xor U27153 (N_27153,N_25385,N_25664);
nor U27154 (N_27154,N_25811,N_25853);
and U27155 (N_27155,N_25247,N_24450);
or U27156 (N_27156,N_25562,N_25781);
nand U27157 (N_27157,N_25423,N_24824);
nand U27158 (N_27158,N_24209,N_24189);
and U27159 (N_27159,N_24112,N_24821);
or U27160 (N_27160,N_24044,N_25286);
and U27161 (N_27161,N_25989,N_24579);
nor U27162 (N_27162,N_25295,N_24513);
or U27163 (N_27163,N_25042,N_25976);
nor U27164 (N_27164,N_25520,N_25910);
xnor U27165 (N_27165,N_25830,N_25413);
and U27166 (N_27166,N_25551,N_24325);
nand U27167 (N_27167,N_24838,N_25006);
xnor U27168 (N_27168,N_25663,N_25527);
or U27169 (N_27169,N_24995,N_25381);
nand U27170 (N_27170,N_25341,N_25673);
xor U27171 (N_27171,N_25612,N_24438);
nor U27172 (N_27172,N_24183,N_25490);
nand U27173 (N_27173,N_25470,N_24678);
and U27174 (N_27174,N_24380,N_24127);
and U27175 (N_27175,N_24362,N_25247);
nor U27176 (N_27176,N_25437,N_25276);
or U27177 (N_27177,N_24768,N_24288);
nor U27178 (N_27178,N_24965,N_24996);
and U27179 (N_27179,N_24273,N_25451);
nand U27180 (N_27180,N_25298,N_24515);
and U27181 (N_27181,N_24484,N_24483);
nor U27182 (N_27182,N_24062,N_25211);
nand U27183 (N_27183,N_25307,N_24038);
xor U27184 (N_27184,N_25489,N_24934);
xor U27185 (N_27185,N_25477,N_25825);
nand U27186 (N_27186,N_25261,N_25595);
or U27187 (N_27187,N_24487,N_24725);
and U27188 (N_27188,N_24885,N_24788);
and U27189 (N_27189,N_24443,N_25765);
or U27190 (N_27190,N_24670,N_25718);
and U27191 (N_27191,N_24274,N_25435);
and U27192 (N_27192,N_24296,N_24464);
and U27193 (N_27193,N_25834,N_25830);
nor U27194 (N_27194,N_24742,N_24666);
xnor U27195 (N_27195,N_25777,N_24094);
or U27196 (N_27196,N_24927,N_24188);
nand U27197 (N_27197,N_25565,N_25645);
and U27198 (N_27198,N_25063,N_25538);
or U27199 (N_27199,N_24405,N_24502);
xnor U27200 (N_27200,N_24893,N_25098);
nor U27201 (N_27201,N_25695,N_25562);
and U27202 (N_27202,N_25717,N_25519);
nor U27203 (N_27203,N_24133,N_24599);
or U27204 (N_27204,N_25084,N_24389);
nor U27205 (N_27205,N_25799,N_24314);
nor U27206 (N_27206,N_24516,N_24233);
xor U27207 (N_27207,N_24976,N_25175);
nor U27208 (N_27208,N_25706,N_24441);
nor U27209 (N_27209,N_25898,N_25962);
nor U27210 (N_27210,N_25215,N_24714);
or U27211 (N_27211,N_25437,N_25294);
nand U27212 (N_27212,N_25947,N_25575);
nor U27213 (N_27213,N_24831,N_24730);
nand U27214 (N_27214,N_25938,N_24860);
or U27215 (N_27215,N_25937,N_25626);
xnor U27216 (N_27216,N_25156,N_24016);
nor U27217 (N_27217,N_24601,N_25793);
xnor U27218 (N_27218,N_24397,N_24585);
nand U27219 (N_27219,N_25535,N_25686);
nand U27220 (N_27220,N_25556,N_24157);
xor U27221 (N_27221,N_25418,N_25421);
xor U27222 (N_27222,N_24261,N_25865);
and U27223 (N_27223,N_24695,N_25330);
or U27224 (N_27224,N_25586,N_24120);
nand U27225 (N_27225,N_24681,N_24051);
nand U27226 (N_27226,N_25929,N_25421);
xnor U27227 (N_27227,N_25021,N_24545);
xor U27228 (N_27228,N_24871,N_24760);
nor U27229 (N_27229,N_25025,N_24424);
nand U27230 (N_27230,N_24793,N_24357);
xor U27231 (N_27231,N_24249,N_24004);
or U27232 (N_27232,N_25308,N_24477);
xnor U27233 (N_27233,N_24845,N_24781);
nor U27234 (N_27234,N_24277,N_25467);
nand U27235 (N_27235,N_25448,N_25765);
xor U27236 (N_27236,N_24458,N_24120);
nand U27237 (N_27237,N_25342,N_24355);
nand U27238 (N_27238,N_25513,N_24285);
or U27239 (N_27239,N_24497,N_24099);
nand U27240 (N_27240,N_25727,N_24540);
and U27241 (N_27241,N_24987,N_25541);
nor U27242 (N_27242,N_25491,N_24217);
or U27243 (N_27243,N_25202,N_25127);
and U27244 (N_27244,N_24957,N_24208);
and U27245 (N_27245,N_24567,N_24013);
and U27246 (N_27246,N_24215,N_25484);
and U27247 (N_27247,N_25699,N_25655);
xnor U27248 (N_27248,N_24572,N_25595);
nor U27249 (N_27249,N_24029,N_24528);
and U27250 (N_27250,N_25484,N_24022);
and U27251 (N_27251,N_25787,N_24618);
xor U27252 (N_27252,N_25259,N_25927);
nor U27253 (N_27253,N_24380,N_25996);
or U27254 (N_27254,N_25678,N_24813);
nor U27255 (N_27255,N_24749,N_25944);
xnor U27256 (N_27256,N_25332,N_25529);
nand U27257 (N_27257,N_24700,N_25290);
nor U27258 (N_27258,N_25079,N_25735);
and U27259 (N_27259,N_24167,N_25131);
or U27260 (N_27260,N_24226,N_24489);
xnor U27261 (N_27261,N_25748,N_24746);
nand U27262 (N_27262,N_25740,N_25863);
or U27263 (N_27263,N_25618,N_24513);
xor U27264 (N_27264,N_25081,N_25432);
or U27265 (N_27265,N_25232,N_24488);
and U27266 (N_27266,N_25899,N_25353);
xor U27267 (N_27267,N_25125,N_25932);
or U27268 (N_27268,N_24545,N_24287);
xor U27269 (N_27269,N_25906,N_25834);
xor U27270 (N_27270,N_25203,N_25222);
nor U27271 (N_27271,N_24746,N_25255);
and U27272 (N_27272,N_25056,N_25412);
nor U27273 (N_27273,N_25705,N_24650);
and U27274 (N_27274,N_24496,N_25246);
or U27275 (N_27275,N_24782,N_24143);
nand U27276 (N_27276,N_25301,N_24788);
nor U27277 (N_27277,N_25899,N_25039);
nor U27278 (N_27278,N_24216,N_25322);
nand U27279 (N_27279,N_25151,N_25862);
nor U27280 (N_27280,N_24110,N_24526);
nand U27281 (N_27281,N_24120,N_24538);
or U27282 (N_27282,N_25339,N_24378);
and U27283 (N_27283,N_25915,N_24874);
nand U27284 (N_27284,N_24604,N_24829);
nand U27285 (N_27285,N_25735,N_25890);
nor U27286 (N_27286,N_25007,N_25094);
nor U27287 (N_27287,N_24149,N_24214);
nand U27288 (N_27288,N_25372,N_25841);
xor U27289 (N_27289,N_25401,N_24614);
or U27290 (N_27290,N_25602,N_24611);
nand U27291 (N_27291,N_24567,N_25009);
nor U27292 (N_27292,N_25300,N_25474);
xor U27293 (N_27293,N_25562,N_24702);
or U27294 (N_27294,N_25248,N_24898);
or U27295 (N_27295,N_24701,N_24568);
nand U27296 (N_27296,N_24100,N_25788);
nor U27297 (N_27297,N_25992,N_25187);
or U27298 (N_27298,N_25869,N_25365);
nand U27299 (N_27299,N_24982,N_25748);
nor U27300 (N_27300,N_25160,N_25999);
xnor U27301 (N_27301,N_24728,N_25279);
and U27302 (N_27302,N_25259,N_25180);
xnor U27303 (N_27303,N_24363,N_24732);
nand U27304 (N_27304,N_24714,N_24101);
nor U27305 (N_27305,N_24313,N_25472);
nand U27306 (N_27306,N_25028,N_24642);
nand U27307 (N_27307,N_24266,N_24944);
nand U27308 (N_27308,N_25142,N_25800);
xnor U27309 (N_27309,N_25193,N_25216);
nand U27310 (N_27310,N_24964,N_25095);
or U27311 (N_27311,N_24969,N_24987);
and U27312 (N_27312,N_24711,N_24517);
nand U27313 (N_27313,N_24670,N_25945);
nor U27314 (N_27314,N_24452,N_24165);
nand U27315 (N_27315,N_24227,N_25859);
nand U27316 (N_27316,N_24406,N_25194);
nand U27317 (N_27317,N_25692,N_25231);
xor U27318 (N_27318,N_24382,N_25040);
nor U27319 (N_27319,N_24460,N_25105);
nor U27320 (N_27320,N_24497,N_24081);
and U27321 (N_27321,N_24493,N_24580);
xnor U27322 (N_27322,N_24139,N_25150);
and U27323 (N_27323,N_25554,N_25556);
nor U27324 (N_27324,N_24641,N_24539);
nor U27325 (N_27325,N_25523,N_24625);
nand U27326 (N_27326,N_24916,N_24134);
nor U27327 (N_27327,N_24537,N_25152);
xor U27328 (N_27328,N_25376,N_25065);
nor U27329 (N_27329,N_25499,N_24709);
xor U27330 (N_27330,N_25244,N_25171);
nor U27331 (N_27331,N_25910,N_24217);
nor U27332 (N_27332,N_24554,N_24306);
nand U27333 (N_27333,N_24495,N_25995);
nor U27334 (N_27334,N_24719,N_25794);
xnor U27335 (N_27335,N_24235,N_25936);
xor U27336 (N_27336,N_24475,N_24661);
and U27337 (N_27337,N_25920,N_25460);
and U27338 (N_27338,N_24386,N_24584);
nand U27339 (N_27339,N_25221,N_24870);
nor U27340 (N_27340,N_24370,N_25374);
xnor U27341 (N_27341,N_24206,N_25278);
nor U27342 (N_27342,N_24965,N_25519);
xor U27343 (N_27343,N_25899,N_25106);
xor U27344 (N_27344,N_25818,N_25694);
nand U27345 (N_27345,N_24047,N_25685);
nor U27346 (N_27346,N_25973,N_25325);
nor U27347 (N_27347,N_25556,N_24559);
xor U27348 (N_27348,N_24574,N_25917);
or U27349 (N_27349,N_25569,N_25942);
or U27350 (N_27350,N_24521,N_25065);
or U27351 (N_27351,N_24369,N_24555);
nand U27352 (N_27352,N_25488,N_25089);
or U27353 (N_27353,N_25250,N_25913);
and U27354 (N_27354,N_24128,N_24563);
nand U27355 (N_27355,N_24111,N_25749);
nand U27356 (N_27356,N_24554,N_24793);
nand U27357 (N_27357,N_25991,N_25140);
and U27358 (N_27358,N_25681,N_25509);
and U27359 (N_27359,N_25502,N_24524);
and U27360 (N_27360,N_24220,N_24508);
and U27361 (N_27361,N_25711,N_24438);
nand U27362 (N_27362,N_24377,N_24929);
nand U27363 (N_27363,N_25558,N_24487);
or U27364 (N_27364,N_25080,N_25605);
xor U27365 (N_27365,N_25554,N_25229);
and U27366 (N_27366,N_25616,N_24625);
and U27367 (N_27367,N_25237,N_24015);
nand U27368 (N_27368,N_25491,N_24605);
nand U27369 (N_27369,N_25612,N_24790);
nand U27370 (N_27370,N_24822,N_25400);
or U27371 (N_27371,N_24479,N_24226);
and U27372 (N_27372,N_24776,N_25939);
and U27373 (N_27373,N_24965,N_25061);
nor U27374 (N_27374,N_25372,N_24978);
nand U27375 (N_27375,N_24799,N_24131);
nor U27376 (N_27376,N_25525,N_25713);
xnor U27377 (N_27377,N_24313,N_24608);
or U27378 (N_27378,N_25506,N_24797);
nor U27379 (N_27379,N_24637,N_24138);
xor U27380 (N_27380,N_24405,N_24808);
nand U27381 (N_27381,N_25430,N_24921);
xor U27382 (N_27382,N_25411,N_24154);
nor U27383 (N_27383,N_24802,N_25828);
or U27384 (N_27384,N_24702,N_25586);
or U27385 (N_27385,N_25458,N_25322);
or U27386 (N_27386,N_25054,N_25285);
xnor U27387 (N_27387,N_25288,N_24935);
nand U27388 (N_27388,N_24954,N_25478);
nor U27389 (N_27389,N_24639,N_24256);
and U27390 (N_27390,N_25413,N_24406);
and U27391 (N_27391,N_24311,N_25700);
nor U27392 (N_27392,N_25299,N_24084);
nor U27393 (N_27393,N_24526,N_24613);
nand U27394 (N_27394,N_24031,N_25439);
xnor U27395 (N_27395,N_24111,N_24242);
and U27396 (N_27396,N_24896,N_25038);
or U27397 (N_27397,N_24610,N_24886);
nor U27398 (N_27398,N_24315,N_25359);
or U27399 (N_27399,N_25908,N_25690);
nand U27400 (N_27400,N_25758,N_25388);
nand U27401 (N_27401,N_24749,N_25354);
and U27402 (N_27402,N_25159,N_24572);
xor U27403 (N_27403,N_24596,N_24993);
nor U27404 (N_27404,N_25589,N_24984);
xor U27405 (N_27405,N_24721,N_25082);
or U27406 (N_27406,N_25436,N_24073);
and U27407 (N_27407,N_24214,N_25465);
or U27408 (N_27408,N_24838,N_24758);
or U27409 (N_27409,N_24068,N_25755);
or U27410 (N_27410,N_25556,N_24079);
and U27411 (N_27411,N_25512,N_25906);
and U27412 (N_27412,N_25934,N_24370);
nor U27413 (N_27413,N_24150,N_25890);
or U27414 (N_27414,N_25390,N_25079);
nor U27415 (N_27415,N_24926,N_24604);
and U27416 (N_27416,N_25009,N_25330);
xnor U27417 (N_27417,N_25608,N_25306);
and U27418 (N_27418,N_25646,N_25559);
xnor U27419 (N_27419,N_24027,N_25993);
and U27420 (N_27420,N_24721,N_25368);
or U27421 (N_27421,N_24920,N_25452);
nand U27422 (N_27422,N_25219,N_25018);
nand U27423 (N_27423,N_25737,N_24784);
and U27424 (N_27424,N_24318,N_24212);
nand U27425 (N_27425,N_25145,N_24977);
nand U27426 (N_27426,N_24699,N_25639);
nor U27427 (N_27427,N_24426,N_25248);
nand U27428 (N_27428,N_24843,N_24870);
or U27429 (N_27429,N_24006,N_24260);
and U27430 (N_27430,N_25903,N_25801);
or U27431 (N_27431,N_25743,N_24990);
nand U27432 (N_27432,N_24676,N_24695);
nand U27433 (N_27433,N_24726,N_25953);
or U27434 (N_27434,N_24461,N_25238);
nand U27435 (N_27435,N_25277,N_24671);
xnor U27436 (N_27436,N_24555,N_25217);
and U27437 (N_27437,N_24073,N_24739);
nor U27438 (N_27438,N_24757,N_24468);
or U27439 (N_27439,N_24690,N_24351);
or U27440 (N_27440,N_25772,N_25006);
and U27441 (N_27441,N_25756,N_24349);
nor U27442 (N_27442,N_25904,N_25839);
and U27443 (N_27443,N_25821,N_24918);
nor U27444 (N_27444,N_25285,N_24821);
xor U27445 (N_27445,N_25641,N_25347);
nor U27446 (N_27446,N_25195,N_24354);
and U27447 (N_27447,N_25714,N_25487);
or U27448 (N_27448,N_24588,N_24275);
nor U27449 (N_27449,N_24664,N_24677);
and U27450 (N_27450,N_25247,N_25763);
or U27451 (N_27451,N_24909,N_25889);
and U27452 (N_27452,N_24537,N_25344);
nand U27453 (N_27453,N_24790,N_25098);
and U27454 (N_27454,N_25360,N_25878);
nor U27455 (N_27455,N_25289,N_24001);
or U27456 (N_27456,N_24397,N_25414);
and U27457 (N_27457,N_24306,N_24010);
nor U27458 (N_27458,N_24421,N_25128);
nand U27459 (N_27459,N_25157,N_25254);
xor U27460 (N_27460,N_24600,N_24825);
and U27461 (N_27461,N_25257,N_25032);
and U27462 (N_27462,N_25803,N_25301);
nand U27463 (N_27463,N_25332,N_24331);
nand U27464 (N_27464,N_24172,N_25050);
and U27465 (N_27465,N_25414,N_24096);
nor U27466 (N_27466,N_24720,N_25381);
nor U27467 (N_27467,N_24182,N_24880);
and U27468 (N_27468,N_25188,N_25183);
and U27469 (N_27469,N_25509,N_25311);
nand U27470 (N_27470,N_24719,N_25662);
and U27471 (N_27471,N_24703,N_25998);
nand U27472 (N_27472,N_24762,N_25270);
nand U27473 (N_27473,N_25841,N_24729);
xor U27474 (N_27474,N_25530,N_24935);
nand U27475 (N_27475,N_24675,N_24520);
or U27476 (N_27476,N_25844,N_25799);
nor U27477 (N_27477,N_24834,N_24632);
nand U27478 (N_27478,N_24232,N_25357);
xnor U27479 (N_27479,N_25605,N_24376);
xnor U27480 (N_27480,N_24463,N_24310);
nor U27481 (N_27481,N_24022,N_24465);
and U27482 (N_27482,N_25910,N_24025);
xnor U27483 (N_27483,N_24389,N_25597);
or U27484 (N_27484,N_25476,N_25576);
nand U27485 (N_27485,N_25245,N_24625);
or U27486 (N_27486,N_25320,N_25560);
xor U27487 (N_27487,N_25317,N_25535);
nand U27488 (N_27488,N_24928,N_24743);
nand U27489 (N_27489,N_24503,N_25224);
and U27490 (N_27490,N_25357,N_24222);
xnor U27491 (N_27491,N_24713,N_24545);
and U27492 (N_27492,N_24627,N_24675);
nand U27493 (N_27493,N_24645,N_24517);
or U27494 (N_27494,N_24014,N_25087);
nand U27495 (N_27495,N_25530,N_25039);
and U27496 (N_27496,N_25346,N_25407);
nor U27497 (N_27497,N_25963,N_24094);
nor U27498 (N_27498,N_25495,N_25514);
nor U27499 (N_27499,N_24468,N_25136);
and U27500 (N_27500,N_24415,N_25642);
or U27501 (N_27501,N_25506,N_25612);
and U27502 (N_27502,N_25559,N_25421);
and U27503 (N_27503,N_25185,N_24978);
or U27504 (N_27504,N_25056,N_25837);
and U27505 (N_27505,N_25993,N_25760);
or U27506 (N_27506,N_24700,N_25627);
and U27507 (N_27507,N_24317,N_25196);
and U27508 (N_27508,N_25449,N_24234);
nand U27509 (N_27509,N_24700,N_25168);
nor U27510 (N_27510,N_24605,N_24559);
and U27511 (N_27511,N_25940,N_25028);
and U27512 (N_27512,N_25049,N_24396);
and U27513 (N_27513,N_25141,N_25959);
or U27514 (N_27514,N_25398,N_25757);
nor U27515 (N_27515,N_25665,N_25688);
xor U27516 (N_27516,N_24204,N_25386);
xnor U27517 (N_27517,N_24396,N_24022);
or U27518 (N_27518,N_25280,N_24626);
xnor U27519 (N_27519,N_24551,N_25672);
xor U27520 (N_27520,N_24170,N_25510);
nor U27521 (N_27521,N_24716,N_25781);
and U27522 (N_27522,N_24822,N_25911);
nor U27523 (N_27523,N_24971,N_24044);
or U27524 (N_27524,N_24681,N_24363);
and U27525 (N_27525,N_24988,N_24280);
nor U27526 (N_27526,N_25252,N_25699);
xnor U27527 (N_27527,N_25224,N_24657);
nand U27528 (N_27528,N_24863,N_24140);
or U27529 (N_27529,N_24562,N_24619);
or U27530 (N_27530,N_24901,N_24402);
nor U27531 (N_27531,N_24431,N_24325);
nand U27532 (N_27532,N_24736,N_25028);
nand U27533 (N_27533,N_25573,N_25057);
nor U27534 (N_27534,N_24322,N_25738);
or U27535 (N_27535,N_24236,N_25813);
nor U27536 (N_27536,N_24283,N_24687);
nor U27537 (N_27537,N_24844,N_24869);
and U27538 (N_27538,N_25508,N_24429);
and U27539 (N_27539,N_24408,N_24929);
xor U27540 (N_27540,N_24859,N_24082);
and U27541 (N_27541,N_25665,N_24946);
nor U27542 (N_27542,N_25881,N_24566);
nand U27543 (N_27543,N_25944,N_24216);
xor U27544 (N_27544,N_25461,N_25749);
and U27545 (N_27545,N_24833,N_25720);
xor U27546 (N_27546,N_25518,N_25595);
and U27547 (N_27547,N_24428,N_25462);
nor U27548 (N_27548,N_25719,N_25355);
nand U27549 (N_27549,N_25232,N_24999);
nand U27550 (N_27550,N_25923,N_24063);
nand U27551 (N_27551,N_24482,N_24678);
nand U27552 (N_27552,N_24059,N_25446);
or U27553 (N_27553,N_25672,N_24947);
or U27554 (N_27554,N_24211,N_25315);
nand U27555 (N_27555,N_25621,N_25719);
xnor U27556 (N_27556,N_24001,N_24319);
nand U27557 (N_27557,N_24020,N_25883);
xor U27558 (N_27558,N_25119,N_25149);
and U27559 (N_27559,N_25151,N_24720);
xnor U27560 (N_27560,N_24433,N_24564);
and U27561 (N_27561,N_24379,N_25627);
nand U27562 (N_27562,N_25029,N_24296);
and U27563 (N_27563,N_25060,N_24295);
and U27564 (N_27564,N_24799,N_24984);
nand U27565 (N_27565,N_25372,N_25950);
xnor U27566 (N_27566,N_25893,N_25859);
and U27567 (N_27567,N_24474,N_24330);
or U27568 (N_27568,N_25485,N_25672);
xnor U27569 (N_27569,N_25588,N_24320);
and U27570 (N_27570,N_25883,N_25286);
nand U27571 (N_27571,N_24628,N_24334);
and U27572 (N_27572,N_25332,N_24343);
nand U27573 (N_27573,N_24786,N_24040);
nor U27574 (N_27574,N_25132,N_24126);
nand U27575 (N_27575,N_25270,N_25030);
and U27576 (N_27576,N_24811,N_25794);
nor U27577 (N_27577,N_24219,N_25047);
nand U27578 (N_27578,N_25165,N_24957);
nand U27579 (N_27579,N_25322,N_25273);
and U27580 (N_27580,N_24951,N_25108);
nor U27581 (N_27581,N_25853,N_24526);
nor U27582 (N_27582,N_25897,N_25351);
and U27583 (N_27583,N_24663,N_25304);
xnor U27584 (N_27584,N_24597,N_24721);
nand U27585 (N_27585,N_25884,N_25469);
or U27586 (N_27586,N_24190,N_25538);
nand U27587 (N_27587,N_25395,N_24237);
nand U27588 (N_27588,N_25363,N_25476);
or U27589 (N_27589,N_24806,N_25979);
and U27590 (N_27590,N_24512,N_24978);
xnor U27591 (N_27591,N_24996,N_25064);
nand U27592 (N_27592,N_25123,N_25401);
or U27593 (N_27593,N_24151,N_24744);
nand U27594 (N_27594,N_24676,N_24894);
nand U27595 (N_27595,N_24085,N_24835);
nor U27596 (N_27596,N_24076,N_25033);
nand U27597 (N_27597,N_24102,N_24231);
nand U27598 (N_27598,N_24841,N_24450);
or U27599 (N_27599,N_24640,N_25259);
or U27600 (N_27600,N_24238,N_24926);
or U27601 (N_27601,N_25619,N_25840);
or U27602 (N_27602,N_25905,N_24957);
nor U27603 (N_27603,N_24488,N_25056);
and U27604 (N_27604,N_25346,N_25539);
or U27605 (N_27605,N_24416,N_25901);
nor U27606 (N_27606,N_25162,N_24121);
xor U27607 (N_27607,N_24812,N_25426);
xnor U27608 (N_27608,N_25530,N_24971);
or U27609 (N_27609,N_24299,N_25977);
or U27610 (N_27610,N_24932,N_24139);
and U27611 (N_27611,N_24085,N_25131);
and U27612 (N_27612,N_25769,N_25639);
or U27613 (N_27613,N_24794,N_24842);
or U27614 (N_27614,N_24006,N_24050);
xor U27615 (N_27615,N_24904,N_25287);
or U27616 (N_27616,N_24121,N_25553);
nor U27617 (N_27617,N_24837,N_25665);
or U27618 (N_27618,N_25583,N_24462);
and U27619 (N_27619,N_24678,N_25760);
nand U27620 (N_27620,N_24025,N_24770);
xnor U27621 (N_27621,N_24597,N_24325);
nor U27622 (N_27622,N_24198,N_25905);
or U27623 (N_27623,N_25751,N_24021);
or U27624 (N_27624,N_24226,N_25228);
or U27625 (N_27625,N_25376,N_24961);
nand U27626 (N_27626,N_25062,N_25901);
and U27627 (N_27627,N_25265,N_24691);
nor U27628 (N_27628,N_24060,N_25924);
nand U27629 (N_27629,N_25643,N_24810);
xnor U27630 (N_27630,N_24168,N_24560);
xor U27631 (N_27631,N_24621,N_25793);
and U27632 (N_27632,N_25519,N_24763);
xor U27633 (N_27633,N_25746,N_25413);
xor U27634 (N_27634,N_25494,N_25787);
nor U27635 (N_27635,N_24946,N_25882);
nor U27636 (N_27636,N_25251,N_25353);
nand U27637 (N_27637,N_25383,N_25134);
xnor U27638 (N_27638,N_24337,N_24544);
xor U27639 (N_27639,N_25614,N_25300);
xor U27640 (N_27640,N_25092,N_25230);
and U27641 (N_27641,N_25227,N_25779);
and U27642 (N_27642,N_25981,N_24765);
nand U27643 (N_27643,N_25883,N_24768);
xor U27644 (N_27644,N_25549,N_24240);
or U27645 (N_27645,N_24213,N_24304);
nand U27646 (N_27646,N_24173,N_25008);
xor U27647 (N_27647,N_25012,N_25733);
or U27648 (N_27648,N_24903,N_24524);
nand U27649 (N_27649,N_25303,N_24275);
and U27650 (N_27650,N_25303,N_25947);
or U27651 (N_27651,N_24195,N_25184);
or U27652 (N_27652,N_25150,N_25122);
xnor U27653 (N_27653,N_24308,N_25537);
xnor U27654 (N_27654,N_25708,N_24092);
nor U27655 (N_27655,N_24047,N_25345);
nor U27656 (N_27656,N_24096,N_24638);
and U27657 (N_27657,N_24057,N_25314);
xor U27658 (N_27658,N_24579,N_25333);
nor U27659 (N_27659,N_24477,N_25783);
nor U27660 (N_27660,N_25672,N_24781);
nand U27661 (N_27661,N_24369,N_24289);
xor U27662 (N_27662,N_25199,N_24704);
or U27663 (N_27663,N_24325,N_24125);
or U27664 (N_27664,N_25349,N_24150);
xor U27665 (N_27665,N_24729,N_25090);
or U27666 (N_27666,N_24822,N_24797);
xor U27667 (N_27667,N_24395,N_24899);
or U27668 (N_27668,N_24193,N_24401);
nor U27669 (N_27669,N_24573,N_25263);
or U27670 (N_27670,N_24394,N_24998);
and U27671 (N_27671,N_24648,N_24156);
nor U27672 (N_27672,N_25517,N_24872);
and U27673 (N_27673,N_24010,N_25017);
nor U27674 (N_27674,N_25749,N_24601);
or U27675 (N_27675,N_24870,N_25819);
nand U27676 (N_27676,N_24564,N_25638);
nand U27677 (N_27677,N_24883,N_24625);
and U27678 (N_27678,N_24928,N_24391);
nor U27679 (N_27679,N_24549,N_25406);
nor U27680 (N_27680,N_25335,N_25080);
or U27681 (N_27681,N_25031,N_24971);
xor U27682 (N_27682,N_24103,N_25448);
nand U27683 (N_27683,N_25240,N_25405);
or U27684 (N_27684,N_24404,N_24289);
and U27685 (N_27685,N_24177,N_24509);
or U27686 (N_27686,N_25520,N_24202);
or U27687 (N_27687,N_25021,N_24815);
nand U27688 (N_27688,N_24512,N_25000);
nand U27689 (N_27689,N_25922,N_25673);
xnor U27690 (N_27690,N_25344,N_24825);
xor U27691 (N_27691,N_24963,N_25850);
or U27692 (N_27692,N_25698,N_25598);
or U27693 (N_27693,N_25740,N_24616);
nor U27694 (N_27694,N_24808,N_25606);
nand U27695 (N_27695,N_24077,N_25329);
nand U27696 (N_27696,N_25558,N_24886);
or U27697 (N_27697,N_25566,N_25922);
or U27698 (N_27698,N_24653,N_25178);
xor U27699 (N_27699,N_24798,N_24661);
nand U27700 (N_27700,N_25094,N_25737);
nand U27701 (N_27701,N_24734,N_25572);
nand U27702 (N_27702,N_24136,N_24427);
or U27703 (N_27703,N_25292,N_25894);
and U27704 (N_27704,N_24068,N_24921);
xnor U27705 (N_27705,N_25004,N_24891);
nand U27706 (N_27706,N_25609,N_24849);
and U27707 (N_27707,N_25292,N_25874);
and U27708 (N_27708,N_25685,N_25362);
or U27709 (N_27709,N_24326,N_24165);
nand U27710 (N_27710,N_25211,N_24624);
nor U27711 (N_27711,N_25100,N_24129);
nor U27712 (N_27712,N_24002,N_25297);
and U27713 (N_27713,N_25164,N_24598);
xor U27714 (N_27714,N_24577,N_25211);
or U27715 (N_27715,N_25660,N_24847);
or U27716 (N_27716,N_24546,N_25828);
nand U27717 (N_27717,N_24519,N_24927);
or U27718 (N_27718,N_24235,N_24569);
xnor U27719 (N_27719,N_25998,N_25209);
nand U27720 (N_27720,N_25963,N_25364);
nor U27721 (N_27721,N_25698,N_24694);
nand U27722 (N_27722,N_25497,N_25834);
xor U27723 (N_27723,N_24899,N_25873);
xnor U27724 (N_27724,N_24030,N_25317);
xor U27725 (N_27725,N_25757,N_25925);
or U27726 (N_27726,N_25826,N_25326);
and U27727 (N_27727,N_25888,N_24994);
nor U27728 (N_27728,N_24473,N_24168);
or U27729 (N_27729,N_24145,N_25788);
or U27730 (N_27730,N_24985,N_24010);
nor U27731 (N_27731,N_25561,N_25311);
nor U27732 (N_27732,N_24674,N_25424);
xor U27733 (N_27733,N_25649,N_25241);
xnor U27734 (N_27734,N_25017,N_24565);
nor U27735 (N_27735,N_24430,N_24723);
or U27736 (N_27736,N_24989,N_25705);
or U27737 (N_27737,N_24320,N_24873);
nand U27738 (N_27738,N_24024,N_25188);
or U27739 (N_27739,N_25727,N_24078);
nor U27740 (N_27740,N_25770,N_25338);
xor U27741 (N_27741,N_24654,N_24024);
xnor U27742 (N_27742,N_25990,N_25937);
nor U27743 (N_27743,N_24837,N_25895);
nor U27744 (N_27744,N_25921,N_24426);
and U27745 (N_27745,N_24172,N_24266);
nand U27746 (N_27746,N_25139,N_25424);
or U27747 (N_27747,N_24407,N_24538);
nor U27748 (N_27748,N_24590,N_25048);
nor U27749 (N_27749,N_24243,N_25537);
nor U27750 (N_27750,N_24904,N_24792);
or U27751 (N_27751,N_24776,N_25962);
and U27752 (N_27752,N_24765,N_25233);
xor U27753 (N_27753,N_25442,N_24380);
xor U27754 (N_27754,N_25182,N_24936);
or U27755 (N_27755,N_25411,N_24337);
and U27756 (N_27756,N_24044,N_25874);
and U27757 (N_27757,N_24520,N_24456);
nand U27758 (N_27758,N_25784,N_24576);
xnor U27759 (N_27759,N_24287,N_24269);
nand U27760 (N_27760,N_25105,N_25669);
or U27761 (N_27761,N_24117,N_25757);
nand U27762 (N_27762,N_25657,N_24624);
nor U27763 (N_27763,N_24486,N_24559);
nor U27764 (N_27764,N_24923,N_25170);
or U27765 (N_27765,N_24880,N_25981);
nand U27766 (N_27766,N_25042,N_25704);
or U27767 (N_27767,N_24925,N_24134);
and U27768 (N_27768,N_24908,N_24263);
or U27769 (N_27769,N_25359,N_25285);
nor U27770 (N_27770,N_25801,N_24999);
nor U27771 (N_27771,N_25648,N_25016);
nor U27772 (N_27772,N_24922,N_24949);
nor U27773 (N_27773,N_24797,N_24647);
or U27774 (N_27774,N_25396,N_25929);
nor U27775 (N_27775,N_25435,N_25575);
nand U27776 (N_27776,N_25857,N_24078);
and U27777 (N_27777,N_24233,N_25814);
and U27778 (N_27778,N_25482,N_24546);
or U27779 (N_27779,N_24328,N_25907);
or U27780 (N_27780,N_25203,N_24331);
and U27781 (N_27781,N_24516,N_24029);
xor U27782 (N_27782,N_25484,N_25572);
or U27783 (N_27783,N_24776,N_25863);
and U27784 (N_27784,N_25666,N_25632);
nand U27785 (N_27785,N_24172,N_24681);
nor U27786 (N_27786,N_24811,N_24012);
and U27787 (N_27787,N_24919,N_25867);
xnor U27788 (N_27788,N_24605,N_25629);
nor U27789 (N_27789,N_25822,N_25462);
and U27790 (N_27790,N_25079,N_24206);
xor U27791 (N_27791,N_25986,N_24431);
nor U27792 (N_27792,N_24104,N_24193);
nand U27793 (N_27793,N_24015,N_25537);
nand U27794 (N_27794,N_25980,N_25285);
xnor U27795 (N_27795,N_24384,N_24978);
or U27796 (N_27796,N_25128,N_25175);
or U27797 (N_27797,N_24019,N_25390);
or U27798 (N_27798,N_25689,N_24612);
or U27799 (N_27799,N_25838,N_25045);
nand U27800 (N_27800,N_25626,N_24541);
or U27801 (N_27801,N_24938,N_25191);
xnor U27802 (N_27802,N_24725,N_25166);
or U27803 (N_27803,N_24628,N_25175);
nor U27804 (N_27804,N_24057,N_25002);
and U27805 (N_27805,N_25481,N_25090);
or U27806 (N_27806,N_25827,N_24120);
nand U27807 (N_27807,N_25910,N_24062);
xnor U27808 (N_27808,N_24334,N_24632);
nand U27809 (N_27809,N_24446,N_24048);
or U27810 (N_27810,N_24119,N_24021);
or U27811 (N_27811,N_25366,N_25762);
xnor U27812 (N_27812,N_24660,N_24018);
or U27813 (N_27813,N_25564,N_24139);
xnor U27814 (N_27814,N_25860,N_25909);
or U27815 (N_27815,N_24626,N_25880);
xnor U27816 (N_27816,N_25311,N_24308);
xor U27817 (N_27817,N_24711,N_24941);
nand U27818 (N_27818,N_24448,N_24661);
or U27819 (N_27819,N_25011,N_24960);
and U27820 (N_27820,N_24916,N_24389);
xnor U27821 (N_27821,N_24803,N_24287);
nand U27822 (N_27822,N_24951,N_24986);
and U27823 (N_27823,N_25089,N_24037);
nor U27824 (N_27824,N_24809,N_25330);
nand U27825 (N_27825,N_25728,N_24944);
or U27826 (N_27826,N_25807,N_24807);
nor U27827 (N_27827,N_24246,N_24495);
or U27828 (N_27828,N_24779,N_25163);
or U27829 (N_27829,N_24185,N_24246);
nor U27830 (N_27830,N_25505,N_24040);
or U27831 (N_27831,N_24733,N_24867);
nor U27832 (N_27832,N_24915,N_25238);
and U27833 (N_27833,N_25448,N_25862);
and U27834 (N_27834,N_24612,N_24375);
and U27835 (N_27835,N_25247,N_25728);
nand U27836 (N_27836,N_24916,N_25647);
and U27837 (N_27837,N_24301,N_25706);
or U27838 (N_27838,N_25386,N_25378);
nor U27839 (N_27839,N_24915,N_25337);
xor U27840 (N_27840,N_25731,N_24685);
nand U27841 (N_27841,N_25942,N_25201);
nand U27842 (N_27842,N_24861,N_25733);
nor U27843 (N_27843,N_25236,N_24509);
and U27844 (N_27844,N_25659,N_24560);
xor U27845 (N_27845,N_24273,N_24171);
and U27846 (N_27846,N_25939,N_25507);
nand U27847 (N_27847,N_25480,N_25267);
xnor U27848 (N_27848,N_25371,N_25597);
xnor U27849 (N_27849,N_24920,N_24806);
xnor U27850 (N_27850,N_24462,N_24465);
nand U27851 (N_27851,N_24951,N_25281);
nand U27852 (N_27852,N_25961,N_24609);
or U27853 (N_27853,N_25752,N_24693);
or U27854 (N_27854,N_24158,N_24620);
nand U27855 (N_27855,N_24175,N_25431);
and U27856 (N_27856,N_25307,N_25224);
nand U27857 (N_27857,N_24621,N_25432);
nor U27858 (N_27858,N_25923,N_25998);
nand U27859 (N_27859,N_25734,N_24117);
nand U27860 (N_27860,N_25736,N_24503);
xnor U27861 (N_27861,N_24798,N_25046);
nand U27862 (N_27862,N_24453,N_24618);
nand U27863 (N_27863,N_25646,N_24302);
or U27864 (N_27864,N_25531,N_25624);
and U27865 (N_27865,N_24502,N_24198);
xor U27866 (N_27866,N_24816,N_24441);
nand U27867 (N_27867,N_24060,N_25570);
nand U27868 (N_27868,N_24056,N_25049);
and U27869 (N_27869,N_25592,N_24496);
nor U27870 (N_27870,N_25140,N_24528);
nor U27871 (N_27871,N_24422,N_24593);
nand U27872 (N_27872,N_24102,N_25731);
or U27873 (N_27873,N_25220,N_25860);
nor U27874 (N_27874,N_25046,N_24600);
nand U27875 (N_27875,N_25748,N_25472);
nor U27876 (N_27876,N_25187,N_25748);
nor U27877 (N_27877,N_24311,N_24778);
nor U27878 (N_27878,N_24784,N_24418);
nor U27879 (N_27879,N_25253,N_24713);
and U27880 (N_27880,N_24533,N_25136);
or U27881 (N_27881,N_24449,N_25312);
nor U27882 (N_27882,N_25271,N_25463);
nand U27883 (N_27883,N_25577,N_25541);
nand U27884 (N_27884,N_24318,N_25153);
and U27885 (N_27885,N_24572,N_25577);
or U27886 (N_27886,N_25087,N_24412);
nor U27887 (N_27887,N_25753,N_24550);
and U27888 (N_27888,N_25263,N_24350);
nor U27889 (N_27889,N_25711,N_25952);
or U27890 (N_27890,N_25986,N_25449);
and U27891 (N_27891,N_25795,N_24269);
xnor U27892 (N_27892,N_25243,N_24099);
nor U27893 (N_27893,N_25788,N_25533);
nor U27894 (N_27894,N_24420,N_25549);
nand U27895 (N_27895,N_25024,N_25231);
and U27896 (N_27896,N_24406,N_25840);
xor U27897 (N_27897,N_25358,N_24545);
xnor U27898 (N_27898,N_25884,N_24172);
nor U27899 (N_27899,N_24315,N_24487);
and U27900 (N_27900,N_25006,N_25621);
and U27901 (N_27901,N_24931,N_24037);
and U27902 (N_27902,N_24338,N_24778);
nor U27903 (N_27903,N_25477,N_24615);
and U27904 (N_27904,N_24767,N_25886);
and U27905 (N_27905,N_24102,N_25357);
xnor U27906 (N_27906,N_24782,N_25921);
xnor U27907 (N_27907,N_24145,N_25725);
or U27908 (N_27908,N_24653,N_24191);
or U27909 (N_27909,N_25803,N_25136);
xor U27910 (N_27910,N_24025,N_25182);
nand U27911 (N_27911,N_24236,N_25494);
xor U27912 (N_27912,N_25628,N_24175);
and U27913 (N_27913,N_24370,N_24164);
nor U27914 (N_27914,N_25197,N_24856);
or U27915 (N_27915,N_24352,N_25626);
or U27916 (N_27916,N_24755,N_24183);
and U27917 (N_27917,N_25015,N_25547);
or U27918 (N_27918,N_24821,N_24676);
and U27919 (N_27919,N_25446,N_25083);
nor U27920 (N_27920,N_25937,N_24565);
and U27921 (N_27921,N_25586,N_25195);
xor U27922 (N_27922,N_25776,N_25959);
and U27923 (N_27923,N_24222,N_25442);
or U27924 (N_27924,N_25321,N_25935);
nor U27925 (N_27925,N_25609,N_25735);
xnor U27926 (N_27926,N_25991,N_25656);
nor U27927 (N_27927,N_25825,N_25108);
or U27928 (N_27928,N_25051,N_25611);
nand U27929 (N_27929,N_25182,N_25031);
nand U27930 (N_27930,N_25194,N_25873);
xnor U27931 (N_27931,N_25513,N_25543);
xor U27932 (N_27932,N_25851,N_25985);
nand U27933 (N_27933,N_25937,N_25623);
nor U27934 (N_27934,N_24432,N_25523);
nand U27935 (N_27935,N_24420,N_24193);
or U27936 (N_27936,N_24660,N_25800);
or U27937 (N_27937,N_25647,N_24647);
and U27938 (N_27938,N_24423,N_24477);
nor U27939 (N_27939,N_24542,N_25482);
and U27940 (N_27940,N_24354,N_24334);
nand U27941 (N_27941,N_24669,N_24412);
or U27942 (N_27942,N_25409,N_25003);
nor U27943 (N_27943,N_24916,N_24800);
and U27944 (N_27944,N_24451,N_24945);
and U27945 (N_27945,N_25431,N_25307);
nor U27946 (N_27946,N_24049,N_24109);
nor U27947 (N_27947,N_24379,N_24671);
and U27948 (N_27948,N_25119,N_24022);
nand U27949 (N_27949,N_24716,N_25119);
or U27950 (N_27950,N_25105,N_24070);
nand U27951 (N_27951,N_24732,N_24154);
or U27952 (N_27952,N_25627,N_25398);
nand U27953 (N_27953,N_25816,N_24351);
nand U27954 (N_27954,N_24384,N_25741);
nand U27955 (N_27955,N_25783,N_25674);
or U27956 (N_27956,N_24051,N_25907);
xnor U27957 (N_27957,N_25231,N_24630);
nand U27958 (N_27958,N_25453,N_24437);
or U27959 (N_27959,N_24304,N_24170);
xor U27960 (N_27960,N_24407,N_25380);
nand U27961 (N_27961,N_24965,N_24908);
or U27962 (N_27962,N_25017,N_24337);
nand U27963 (N_27963,N_25145,N_25471);
nand U27964 (N_27964,N_24410,N_24565);
nor U27965 (N_27965,N_24343,N_24080);
or U27966 (N_27966,N_25384,N_24582);
and U27967 (N_27967,N_25297,N_25941);
and U27968 (N_27968,N_24639,N_25449);
nand U27969 (N_27969,N_25640,N_24089);
nand U27970 (N_27970,N_25426,N_25809);
and U27971 (N_27971,N_25013,N_25777);
xor U27972 (N_27972,N_24942,N_24487);
and U27973 (N_27973,N_24566,N_24388);
nor U27974 (N_27974,N_24545,N_25103);
nand U27975 (N_27975,N_25049,N_24103);
nand U27976 (N_27976,N_24193,N_25138);
xnor U27977 (N_27977,N_25056,N_25540);
or U27978 (N_27978,N_25630,N_25075);
nand U27979 (N_27979,N_24373,N_25934);
nor U27980 (N_27980,N_24710,N_24964);
and U27981 (N_27981,N_25806,N_25500);
or U27982 (N_27982,N_25782,N_25302);
or U27983 (N_27983,N_24201,N_24295);
and U27984 (N_27984,N_24795,N_24533);
and U27985 (N_27985,N_24563,N_24636);
or U27986 (N_27986,N_25831,N_25702);
nor U27987 (N_27987,N_24270,N_24192);
nor U27988 (N_27988,N_24700,N_24417);
nand U27989 (N_27989,N_24970,N_24360);
nor U27990 (N_27990,N_24068,N_25241);
or U27991 (N_27991,N_25440,N_25931);
nor U27992 (N_27992,N_25872,N_24123);
or U27993 (N_27993,N_25777,N_24107);
nand U27994 (N_27994,N_24218,N_25638);
and U27995 (N_27995,N_24025,N_24370);
nor U27996 (N_27996,N_25607,N_24087);
or U27997 (N_27997,N_24097,N_25643);
or U27998 (N_27998,N_24943,N_25963);
and U27999 (N_27999,N_25371,N_25289);
or U28000 (N_28000,N_26427,N_27605);
and U28001 (N_28001,N_26115,N_26622);
nand U28002 (N_28002,N_27186,N_27264);
nand U28003 (N_28003,N_26910,N_27749);
and U28004 (N_28004,N_27888,N_27787);
xor U28005 (N_28005,N_26957,N_27346);
and U28006 (N_28006,N_27543,N_27604);
nor U28007 (N_28007,N_27832,N_27699);
nor U28008 (N_28008,N_27139,N_26896);
xnor U28009 (N_28009,N_27815,N_26359);
and U28010 (N_28010,N_26300,N_27780);
nor U28011 (N_28011,N_26110,N_27172);
or U28012 (N_28012,N_26459,N_26731);
and U28013 (N_28013,N_26921,N_26837);
nand U28014 (N_28014,N_27753,N_27056);
nand U28015 (N_28015,N_26696,N_26217);
nand U28016 (N_28016,N_26749,N_27824);
nand U28017 (N_28017,N_27042,N_26079);
xnor U28018 (N_28018,N_26399,N_27043);
nand U28019 (N_28019,N_26833,N_27035);
or U28020 (N_28020,N_27334,N_27214);
xor U28021 (N_28021,N_26712,N_27872);
xor U28022 (N_28022,N_27222,N_26263);
or U28023 (N_28023,N_27251,N_27350);
nand U28024 (N_28024,N_27083,N_27565);
or U28025 (N_28025,N_27695,N_26353);
and U28026 (N_28026,N_26024,N_27986);
nand U28027 (N_28027,N_27521,N_27138);
nand U28028 (N_28028,N_26806,N_27449);
or U28029 (N_28029,N_27135,N_26893);
or U28030 (N_28030,N_27635,N_27512);
xor U28031 (N_28031,N_26343,N_27049);
and U28032 (N_28032,N_26069,N_26061);
xnor U28033 (N_28033,N_26598,N_27996);
nand U28034 (N_28034,N_27812,N_27528);
or U28035 (N_28035,N_27853,N_26911);
nor U28036 (N_28036,N_27638,N_26460);
and U28037 (N_28037,N_27538,N_26119);
or U28038 (N_28038,N_26129,N_27731);
xnor U28039 (N_28039,N_26416,N_27532);
xnor U28040 (N_28040,N_27050,N_27178);
nor U28041 (N_28041,N_27622,N_27240);
nand U28042 (N_28042,N_26941,N_26033);
nor U28043 (N_28043,N_26383,N_26456);
nand U28044 (N_28044,N_26778,N_27151);
nand U28045 (N_28045,N_27848,N_26093);
xor U28046 (N_28046,N_26496,N_26701);
or U28047 (N_28047,N_27886,N_27958);
xor U28048 (N_28048,N_27558,N_26603);
nand U28049 (N_28049,N_27307,N_27961);
nor U28050 (N_28050,N_26414,N_26591);
nand U28051 (N_28051,N_27205,N_27001);
nor U28052 (N_28052,N_27271,N_26873);
or U28053 (N_28053,N_26410,N_27202);
nor U28054 (N_28054,N_26729,N_26154);
and U28055 (N_28055,N_27182,N_26145);
nor U28056 (N_28056,N_26012,N_27450);
or U28057 (N_28057,N_26007,N_26286);
xnor U28058 (N_28058,N_26502,N_27073);
nand U28059 (N_28059,N_26651,N_27705);
and U28060 (N_28060,N_26567,N_26793);
nand U28061 (N_28061,N_26026,N_26962);
xnor U28062 (N_28062,N_26504,N_26705);
and U28063 (N_28063,N_27674,N_27746);
or U28064 (N_28064,N_26083,N_26657);
nand U28065 (N_28065,N_26091,N_27548);
and U28066 (N_28066,N_27319,N_26215);
nand U28067 (N_28067,N_26625,N_26718);
xor U28068 (N_28068,N_26411,N_27806);
xnor U28069 (N_28069,N_27870,N_27219);
or U28070 (N_28070,N_27022,N_27943);
nand U28071 (N_28071,N_27335,N_26108);
nor U28072 (N_28072,N_27134,N_27712);
xnor U28073 (N_28073,N_26754,N_26355);
and U28074 (N_28074,N_26758,N_27226);
nand U28075 (N_28075,N_27892,N_26248);
or U28076 (N_28076,N_26206,N_26076);
nand U28077 (N_28077,N_26085,N_27567);
nor U28078 (N_28078,N_26009,N_27589);
or U28079 (N_28079,N_26429,N_27951);
nand U28080 (N_28080,N_26196,N_27783);
nand U28081 (N_28081,N_27875,N_26054);
and U28082 (N_28082,N_26270,N_26236);
xnor U28083 (N_28083,N_26350,N_27137);
and U28084 (N_28084,N_26051,N_27663);
xor U28085 (N_28085,N_26136,N_27498);
and U28086 (N_28086,N_26272,N_27127);
and U28087 (N_28087,N_27725,N_27442);
nand U28088 (N_28088,N_27502,N_26711);
nor U28089 (N_28089,N_26821,N_27300);
and U28090 (N_28090,N_27244,N_26347);
and U28091 (N_28091,N_27189,N_26305);
nor U28092 (N_28092,N_27864,N_27614);
nand U28093 (N_28093,N_27509,N_27545);
xnor U28094 (N_28094,N_27715,N_26363);
nor U28095 (N_28095,N_26938,N_26838);
nor U28096 (N_28096,N_27929,N_26229);
xor U28097 (N_28097,N_26843,N_27945);
nand U28098 (N_28098,N_27418,N_26530);
nor U28099 (N_28099,N_27184,N_26317);
nand U28100 (N_28100,N_27341,N_26401);
nor U28101 (N_28101,N_26213,N_26223);
nor U28102 (N_28102,N_26249,N_27778);
and U28103 (N_28103,N_26855,N_26038);
and U28104 (N_28104,N_27713,N_27293);
nor U28105 (N_28105,N_26779,N_26785);
nand U28106 (N_28106,N_26207,N_26869);
nand U28107 (N_28107,N_27084,N_27131);
or U28108 (N_28108,N_27523,N_27484);
nor U28109 (N_28109,N_26074,N_26548);
and U28110 (N_28110,N_26037,N_26543);
xor U28111 (N_28111,N_27637,N_27036);
xor U28112 (N_28112,N_26694,N_27069);
and U28113 (N_28113,N_27594,N_27597);
nand U28114 (N_28114,N_26084,N_27174);
xor U28115 (N_28115,N_26589,N_27499);
nand U28116 (N_28116,N_27088,N_26916);
and U28117 (N_28117,N_27469,N_26588);
or U28118 (N_28118,N_27505,N_27006);
or U28119 (N_28119,N_26848,N_27018);
and U28120 (N_28120,N_26203,N_26010);
xor U28121 (N_28121,N_27800,N_27950);
nand U28122 (N_28122,N_26972,N_27694);
nand U28123 (N_28123,N_26936,N_27587);
nor U28124 (N_28124,N_27515,N_27145);
xor U28125 (N_28125,N_27889,N_27366);
nand U28126 (N_28126,N_26608,N_26040);
nor U28127 (N_28127,N_27629,N_27337);
xor U28128 (N_28128,N_26540,N_27033);
xnor U28129 (N_28129,N_26652,N_27369);
nand U28130 (N_28130,N_27031,N_26420);
xor U28131 (N_28131,N_26716,N_26755);
nor U28132 (N_28132,N_27267,N_26982);
and U28133 (N_28133,N_27061,N_27952);
xor U28134 (N_28134,N_26812,N_27039);
and U28135 (N_28135,N_27308,N_27243);
nand U28136 (N_28136,N_27852,N_26225);
nor U28137 (N_28137,N_26759,N_27011);
or U28138 (N_28138,N_26509,N_26137);
xnor U28139 (N_28139,N_27782,N_26049);
or U28140 (N_28140,N_26524,N_27680);
and U28141 (N_28141,N_26555,N_27093);
nor U28142 (N_28142,N_26887,N_27406);
or U28143 (N_28143,N_26200,N_27917);
or U28144 (N_28144,N_26708,N_26440);
nand U28145 (N_28145,N_26523,N_27736);
xor U28146 (N_28146,N_27737,N_27647);
xor U28147 (N_28147,N_26841,N_27352);
nand U28148 (N_28148,N_26082,N_26426);
nand U28149 (N_28149,N_27707,N_26304);
nor U28150 (N_28150,N_26547,N_27317);
and U28151 (N_28151,N_26807,N_26571);
and U28152 (N_28152,N_26597,N_27455);
xnor U28153 (N_28153,N_26665,N_26528);
nor U28154 (N_28154,N_27690,N_26782);
or U28155 (N_28155,N_27378,N_27381);
nand U28156 (N_28156,N_26538,N_27479);
nor U28157 (N_28157,N_27960,N_27197);
and U28158 (N_28158,N_26212,N_27171);
nand U28159 (N_28159,N_27314,N_27285);
xor U28160 (N_28160,N_26867,N_26802);
and U28161 (N_28161,N_27403,N_26556);
nand U28162 (N_28162,N_26211,N_27415);
nor U28163 (N_28163,N_26576,N_26089);
nand U28164 (N_28164,N_27908,N_26422);
or U28165 (N_28165,N_27072,N_27053);
nand U28166 (N_28166,N_27891,N_26158);
and U28167 (N_28167,N_26457,N_26011);
nor U28168 (N_28168,N_27054,N_26878);
and U28169 (N_28169,N_27631,N_27173);
nor U28170 (N_28170,N_27992,N_26258);
or U28171 (N_28171,N_27191,N_27600);
and U28172 (N_28172,N_26336,N_27164);
nand U28173 (N_28173,N_27693,N_26232);
nor U28174 (N_28174,N_27772,N_26561);
xor U28175 (N_28175,N_26617,N_27873);
and U28176 (N_28176,N_26455,N_27212);
nor U28177 (N_28177,N_26857,N_26851);
or U28178 (N_28178,N_27167,N_26393);
nand U28179 (N_28179,N_27497,N_27210);
xor U28180 (N_28180,N_26070,N_26021);
xnor U28181 (N_28181,N_27867,N_26606);
xor U28182 (N_28182,N_27291,N_26565);
xor U28183 (N_28183,N_27785,N_26402);
xnor U28184 (N_28184,N_27717,N_27642);
nor U28185 (N_28185,N_26053,N_26376);
nand U28186 (N_28186,N_26488,N_27862);
xnor U28187 (N_28187,N_27326,N_26473);
xnor U28188 (N_28188,N_27117,N_26319);
or U28189 (N_28189,N_26058,N_27048);
and U28190 (N_28190,N_26439,N_26193);
and U28191 (N_28191,N_26719,N_27492);
nand U28192 (N_28192,N_26739,N_27621);
nor U28193 (N_28193,N_26819,N_27411);
nor U28194 (N_28194,N_27767,N_26649);
xnor U28195 (N_28195,N_26486,N_27985);
xor U28196 (N_28196,N_27551,N_27322);
and U28197 (N_28197,N_26105,N_27994);
nand U28198 (N_28198,N_26480,N_27227);
nand U28199 (N_28199,N_27382,N_27420);
nand U28200 (N_28200,N_26859,N_27000);
nand U28201 (N_28201,N_26165,N_26358);
or U28202 (N_28202,N_27128,N_26333);
xor U28203 (N_28203,N_26640,N_26464);
or U28204 (N_28204,N_27355,N_27997);
xnor U28205 (N_28205,N_26844,N_26906);
or U28206 (N_28206,N_27801,N_26398);
xnor U28207 (N_28207,N_27234,N_26506);
xor U28208 (N_28208,N_26991,N_26299);
and U28209 (N_28209,N_26308,N_27585);
and U28210 (N_28210,N_26999,N_27866);
and U28211 (N_28211,N_26149,N_26043);
xor U28212 (N_28212,N_27909,N_27799);
or U28213 (N_28213,N_27067,N_26963);
or U28214 (N_28214,N_26901,N_26527);
nand U28215 (N_28215,N_26346,N_26512);
nand U28216 (N_28216,N_27125,N_27401);
and U28217 (N_28217,N_27550,N_27536);
nand U28218 (N_28218,N_27625,N_26418);
and U28219 (N_28219,N_27351,N_27910);
xor U28220 (N_28220,N_26500,N_27295);
nor U28221 (N_28221,N_26392,N_27620);
and U28222 (N_28222,N_26413,N_27461);
nor U28223 (N_28223,N_27196,N_26564);
and U28224 (N_28224,N_26094,N_26927);
nor U28225 (N_28225,N_26503,N_27796);
nor U28226 (N_28226,N_26192,N_27071);
and U28227 (N_28227,N_26202,N_26590);
or U28228 (N_28228,N_26792,N_27878);
or U28229 (N_28229,N_26604,N_27199);
xor U28230 (N_28230,N_26114,N_26293);
xor U28231 (N_28231,N_26948,N_26167);
and U28232 (N_28232,N_27412,N_27974);
and U28233 (N_28233,N_27379,N_26048);
nand U28234 (N_28234,N_27915,N_26148);
or U28235 (N_28235,N_26784,N_27896);
and U28236 (N_28236,N_26199,N_26288);
nand U28237 (N_28237,N_27108,N_26276);
nor U28238 (N_28238,N_26829,N_27390);
nand U28239 (N_28239,N_27204,N_27901);
nor U28240 (N_28240,N_27428,N_27590);
xnor U28241 (N_28241,N_27673,N_26747);
or U28242 (N_28242,N_27941,N_27903);
or U28243 (N_28243,N_27805,N_26198);
and U28244 (N_28244,N_27835,N_27274);
nand U28245 (N_28245,N_27270,N_26130);
or U28246 (N_28246,N_27656,N_27784);
and U28247 (N_28247,N_26680,N_27037);
and U28248 (N_28248,N_26297,N_26431);
nor U28249 (N_28249,N_27847,N_27678);
nand U28250 (N_28250,N_27028,N_27283);
or U28251 (N_28251,N_26075,N_27714);
and U28252 (N_28252,N_27467,N_26031);
and U28253 (N_28253,N_27679,N_27107);
xnor U28254 (N_28254,N_26474,N_26475);
nand U28255 (N_28255,N_26681,N_27819);
or U28256 (N_28256,N_26441,N_27702);
or U28257 (N_28257,N_27046,N_26435);
or U28258 (N_28258,N_26001,N_26790);
xnor U28259 (N_28259,N_26124,N_26808);
or U28260 (N_28260,N_26521,N_27761);
or U28261 (N_28261,N_26809,N_26235);
xnor U28262 (N_28262,N_27675,N_26645);
xnor U28263 (N_28263,N_26799,N_26780);
nor U28264 (N_28264,N_26955,N_26909);
xnor U28265 (N_28265,N_27115,N_26746);
or U28266 (N_28266,N_26531,N_26634);
nand U28267 (N_28267,N_27452,N_26394);
and U28268 (N_28268,N_26720,N_26926);
or U28269 (N_28269,N_27318,N_27561);
or U28270 (N_28270,N_26321,N_26077);
and U28271 (N_28271,N_27948,N_26269);
or U28272 (N_28272,N_27124,N_27681);
nor U28273 (N_28273,N_27798,N_27779);
nand U28274 (N_28274,N_26585,N_27123);
nor U28275 (N_28275,N_26357,N_27101);
and U28276 (N_28276,N_27474,N_26607);
and U28277 (N_28277,N_26632,N_27065);
nand U28278 (N_28278,N_27553,N_26481);
nor U28279 (N_28279,N_27354,N_27010);
nor U28280 (N_28280,N_26047,N_26677);
or U28281 (N_28281,N_27609,N_26143);
nand U28282 (N_28282,N_26157,N_27582);
nand U28283 (N_28283,N_26615,N_26939);
nand U28284 (N_28284,N_26772,N_26244);
or U28285 (N_28285,N_27836,N_26041);
nand U28286 (N_28286,N_27668,N_27162);
nand U28287 (N_28287,N_27791,N_26086);
or U28288 (N_28288,N_26757,N_27289);
and U28289 (N_28289,N_27788,N_27008);
and U28290 (N_28290,N_27444,N_27333);
nand U28291 (N_28291,N_27777,N_27920);
or U28292 (N_28292,N_26783,N_27813);
xnor U28293 (N_28293,N_26662,N_26195);
nand U28294 (N_28294,N_27094,N_27634);
nor U28295 (N_28295,N_26302,N_27932);
nor U28296 (N_28296,N_26903,N_26879);
xnor U28297 (N_28297,N_27651,N_26852);
or U28298 (N_28298,N_27988,N_26678);
and U28299 (N_28299,N_26522,N_26839);
and U28300 (N_28300,N_27064,N_27868);
xor U28301 (N_28301,N_26118,N_26593);
and U28302 (N_28302,N_26518,N_27472);
nand U28303 (N_28303,N_27670,N_26894);
or U28304 (N_28304,N_26624,N_27719);
or U28305 (N_28305,N_27682,N_27644);
or U28306 (N_28306,N_27934,N_26014);
nor U28307 (N_28307,N_26032,N_26151);
or U28308 (N_28308,N_26847,N_26368);
xnor U28309 (N_28309,N_27183,N_27716);
nand U28310 (N_28310,N_26865,N_27760);
nor U28311 (N_28311,N_26928,N_27016);
or U28312 (N_28312,N_27924,N_26324);
nand U28313 (N_28313,N_27809,N_27827);
nor U28314 (N_28314,N_27816,N_27030);
or U28315 (N_28315,N_26993,N_26765);
xnor U28316 (N_28316,N_26447,N_27987);
and U28317 (N_28317,N_26572,N_26382);
xor U28318 (N_28318,N_26536,N_27066);
xor U28319 (N_28319,N_26514,N_27388);
and U28320 (N_28320,N_27328,N_27744);
or U28321 (N_28321,N_26117,N_27342);
nor U28322 (N_28322,N_26810,N_27361);
or U28323 (N_28323,N_26419,N_26127);
xor U28324 (N_28324,N_27757,N_26344);
nor U28325 (N_28325,N_27007,N_26801);
xnor U28326 (N_28326,N_27236,N_26629);
xnor U28327 (N_28327,N_26626,N_27722);
nand U28328 (N_28328,N_27921,N_26914);
xor U28329 (N_28329,N_27849,N_27993);
or U28330 (N_28330,N_27102,N_26261);
xor U28331 (N_28331,N_26423,N_27911);
nor U28332 (N_28332,N_27844,N_27928);
xnor U28333 (N_28333,N_26998,N_27216);
and U28334 (N_28334,N_26967,N_27269);
nand U28335 (N_28335,N_27147,N_26295);
and U28336 (N_28336,N_26631,N_27607);
nand U28337 (N_28337,N_26836,N_27506);
nor U28338 (N_28338,N_26553,N_26562);
nor U28339 (N_28339,N_26688,N_27610);
nor U28340 (N_28340,N_26997,N_26691);
nor U28341 (N_28341,N_27306,N_26717);
and U28342 (N_28342,N_26144,N_26000);
and U28343 (N_28343,N_26811,N_27633);
nand U28344 (N_28344,N_26633,N_26330);
and U28345 (N_28345,N_27579,N_26959);
and U28346 (N_28346,N_27899,N_26654);
or U28347 (N_28347,N_27315,N_26919);
or U28348 (N_28348,N_26237,N_26449);
xnor U28349 (N_28349,N_27114,N_27581);
or U28350 (N_28350,N_26209,N_26513);
nand U28351 (N_28351,N_27936,N_27837);
nor U28352 (N_28352,N_27407,N_27735);
nor U28353 (N_28353,N_26899,N_27554);
nor U28354 (N_28354,N_27990,N_27684);
xnor U28355 (N_28355,N_26977,N_26882);
nand U28356 (N_28356,N_27465,N_26155);
or U28357 (N_28357,N_26684,N_26974);
and U28358 (N_28358,N_27488,N_26947);
xnor U28359 (N_28359,N_27953,N_26294);
xnor U28360 (N_28360,N_27459,N_26123);
xor U28361 (N_28361,N_27817,N_26275);
nand U28362 (N_28362,N_27508,N_27931);
xnor U28363 (N_28363,N_27973,N_26365);
nor U28364 (N_28364,N_27296,N_26113);
xnor U28365 (N_28365,N_26341,N_27246);
and U28366 (N_28366,N_26690,N_27275);
or U28367 (N_28367,N_26306,N_27981);
nor U28368 (N_28368,N_27962,N_26259);
xnor U28369 (N_28369,N_26682,N_26406);
nand U28370 (N_28370,N_27155,N_27615);
nand U28371 (N_28371,N_27068,N_26661);
and U28372 (N_28372,N_27454,N_27721);
and U28373 (N_28373,N_27978,N_27966);
nor U28374 (N_28374,N_27024,N_27169);
nand U28375 (N_28375,N_26642,N_26803);
or U28376 (N_28376,N_26039,N_27012);
or U28377 (N_28377,N_26566,N_27860);
or U28378 (N_28378,N_26723,N_27462);
nand U28379 (N_28379,N_26159,N_26845);
xor U28380 (N_28380,N_26254,N_27880);
xnor U28381 (N_28381,N_26609,N_27198);
or U28382 (N_28382,N_26619,N_26415);
nor U28383 (N_28383,N_27149,N_27116);
nor U28384 (N_28384,N_26954,N_27230);
and U28385 (N_28385,N_26314,N_26380);
nand U28386 (N_28386,N_26722,N_27009);
nor U28387 (N_28387,N_26296,N_27709);
nor U28388 (N_28388,N_27027,N_26933);
xnor U28389 (N_28389,N_26243,N_26262);
nor U28390 (N_28390,N_27483,N_27859);
nor U28391 (N_28391,N_27956,N_27095);
or U28392 (N_28392,N_27165,N_27766);
or U28393 (N_28393,N_27294,N_27413);
nand U28394 (N_28394,N_27794,N_26111);
or U28395 (N_28395,N_27762,N_27666);
or U28396 (N_28396,N_26292,N_26046);
and U28397 (N_28397,N_27259,N_26017);
and U28398 (N_28398,N_26886,N_27999);
xnor U28399 (N_28399,N_26517,N_27365);
or U28400 (N_28400,N_27419,N_26824);
or U28401 (N_28401,N_26025,N_26250);
or U28402 (N_28402,N_27299,N_26692);
xor U28403 (N_28403,N_26951,N_26109);
xor U28404 (N_28404,N_27998,N_27841);
and U28405 (N_28405,N_27305,N_27871);
nor U28406 (N_28406,N_26797,N_27424);
xor U28407 (N_28407,N_26417,N_27003);
or U28408 (N_28408,N_26771,N_26970);
and U28409 (N_28409,N_26871,N_26638);
nand U28410 (N_28410,N_26493,N_26374);
and U28411 (N_28411,N_26139,N_27534);
or U28412 (N_28412,N_27261,N_26854);
or U28413 (N_28413,N_27839,N_26988);
and U28414 (N_28414,N_26580,N_27552);
or U28415 (N_28415,N_27091,N_27949);
nor U28416 (N_28416,N_27795,N_26929);
nor U28417 (N_28417,N_27331,N_26958);
and U28418 (N_28418,N_26950,N_26183);
xnor U28419 (N_28419,N_26776,N_27747);
or U28420 (N_28420,N_26853,N_26730);
nand U28421 (N_28421,N_26541,N_26284);
and U28422 (N_28422,N_26194,N_27383);
or U28423 (N_28423,N_26877,N_27112);
nor U28424 (N_28424,N_26472,N_27229);
and U28425 (N_28425,N_27152,N_27211);
xor U28426 (N_28426,N_27510,N_26816);
nand U28427 (N_28427,N_26850,N_26052);
xor U28428 (N_28428,N_26240,N_27478);
xor U28429 (N_28429,N_27658,N_26822);
nor U28430 (N_28430,N_27393,N_26753);
xor U28431 (N_28431,N_27595,N_26366);
nor U28432 (N_28432,N_27970,N_26761);
nand U28433 (N_28433,N_26471,N_27738);
nand U28434 (N_28434,N_26030,N_26674);
and U28435 (N_28435,N_27623,N_27098);
nand U28436 (N_28436,N_27241,N_27537);
xnor U28437 (N_28437,N_27804,N_26981);
nand U28438 (N_28438,N_26191,N_26693);
and U28439 (N_28439,N_27220,N_27349);
and U28440 (N_28440,N_26301,N_26980);
xnor U28441 (N_28441,N_27159,N_27533);
nor U28442 (N_28442,N_26002,N_27818);
and U28443 (N_28443,N_27976,N_26242);
nand U28444 (N_28444,N_26059,N_26055);
xor U28445 (N_28445,N_26623,N_26160);
nor U28446 (N_28446,N_27154,N_27530);
nor U28447 (N_28447,N_27400,N_26814);
nor U28448 (N_28448,N_26364,N_26599);
nor U28449 (N_28449,N_27168,N_26029);
nor U28450 (N_28450,N_27877,N_27925);
nor U28451 (N_28451,N_26379,N_26768);
nor U28452 (N_28452,N_26329,N_26713);
or U28453 (N_28453,N_27755,N_26228);
or U28454 (N_28454,N_26740,N_27132);
xnor U28455 (N_28455,N_26057,N_27754);
and U28456 (N_28456,N_26327,N_26744);
or U28457 (N_28457,N_26282,N_27792);
nand U28458 (N_28458,N_26444,N_26096);
xor U28459 (N_28459,N_27570,N_27672);
or U28460 (N_28460,N_26386,N_27881);
and U28461 (N_28461,N_27448,N_26405);
xor U28462 (N_28462,N_27312,N_26430);
or U28463 (N_28463,N_27763,N_26796);
xnor U28464 (N_28464,N_27034,N_26320);
xor U28465 (N_28465,N_27580,N_26550);
nand U28466 (N_28466,N_27516,N_26019);
or U28467 (N_28467,N_26056,N_27213);
xnor U28468 (N_28468,N_27504,N_26611);
nor U28469 (N_28469,N_26161,N_26989);
nor U28470 (N_28470,N_27677,N_26125);
or U28471 (N_28471,N_27667,N_27330);
xnor U28472 (N_28472,N_26188,N_26979);
nor U28473 (N_28473,N_27628,N_26614);
nand U28474 (N_28474,N_26062,N_27060);
and U28475 (N_28475,N_27057,N_26602);
nor U28476 (N_28476,N_27922,N_26973);
nand U28477 (N_28477,N_26798,N_27741);
xor U28478 (N_28478,N_26763,N_27503);
xor U28479 (N_28479,N_27734,N_26104);
and U28480 (N_28480,N_26834,N_27616);
and U28481 (N_28481,N_27555,N_27939);
and U28482 (N_28482,N_27279,N_26184);
nand U28483 (N_28483,N_27689,N_27704);
and U28484 (N_28484,N_26815,N_26335);
nand U28485 (N_28485,N_27436,N_26081);
xor U28486 (N_28486,N_27136,N_26505);
xor U28487 (N_28487,N_27527,N_26732);
and U28488 (N_28488,N_26338,N_27397);
or U28489 (N_28489,N_26892,N_27287);
nand U28490 (N_28490,N_27402,N_27372);
nor U28491 (N_28491,N_27657,N_26434);
xnor U28492 (N_28492,N_26735,N_27608);
or U28493 (N_28493,N_26594,N_27514);
and U28494 (N_28494,N_26687,N_26066);
and U28495 (N_28495,N_27923,N_26526);
or U28496 (N_28496,N_26362,N_26099);
and U28497 (N_28497,N_26704,N_27256);
and U28498 (N_28498,N_27569,N_26361);
nand U28499 (N_28499,N_26210,N_26312);
xnor U28500 (N_28500,N_27058,N_26257);
nor U28501 (N_28501,N_26601,N_27468);
nor U28502 (N_28502,N_27414,N_27158);
nor U28503 (N_28503,N_27395,N_26498);
nor U28504 (N_28504,N_26990,N_27119);
nor U28505 (N_28505,N_27458,N_26656);
xor U28506 (N_28506,N_27641,N_27086);
or U28507 (N_28507,N_27052,N_27559);
xnor U28508 (N_28508,N_27089,N_26964);
xor U28509 (N_28509,N_26519,N_26064);
or U28510 (N_28510,N_27075,N_27433);
nand U28511 (N_28511,N_27258,N_27113);
xnor U28512 (N_28512,N_27730,N_26388);
and U28513 (N_28513,N_27564,N_27861);
nand U28514 (N_28514,N_27963,N_27727);
and U28515 (N_28515,N_26018,N_27654);
nor U28516 (N_28516,N_27964,N_27586);
or U28517 (N_28517,N_26310,N_27096);
and U28518 (N_28518,N_27099,N_26710);
nand U28519 (N_28519,N_26045,N_26817);
xnor U28520 (N_28520,N_26858,N_27141);
xor U28521 (N_28521,N_27904,N_27014);
or U28522 (N_28522,N_27288,N_26952);
and U28523 (N_28523,N_26781,N_27652);
or U28524 (N_28524,N_26373,N_26116);
nor U28525 (N_28525,N_27386,N_26573);
xnor U28526 (N_28526,N_27557,N_26908);
nand U28527 (N_28527,N_26214,N_27325);
nand U28528 (N_28528,N_26315,N_26570);
and U28529 (N_28529,N_26133,N_27930);
nor U28530 (N_28530,N_26126,N_26630);
nor U28531 (N_28531,N_26549,N_26351);
nand U28532 (N_28532,N_26985,N_26557);
nor U28533 (N_28533,N_27599,N_27272);
nand U28534 (N_28534,N_26849,N_26818);
and U28535 (N_28535,N_27769,N_26734);
nand U28536 (N_28536,N_27013,N_27445);
nand U28537 (N_28537,N_26996,N_26699);
xor U28538 (N_28538,N_26028,N_27215);
xor U28539 (N_28539,N_27897,N_26006);
nor U28540 (N_28540,N_26073,N_27982);
xnor U28541 (N_28541,N_26381,N_26050);
xnor U28542 (N_28542,N_27257,N_27732);
xor U28543 (N_28543,N_26702,N_27517);
and U28544 (N_28544,N_26279,N_27281);
nand U28545 (N_28545,N_27501,N_26227);
xnor U28546 (N_28546,N_27842,N_26285);
and U28547 (N_28547,N_26864,N_26995);
or U28548 (N_28548,N_26403,N_26542);
nand U28549 (N_28549,N_27063,N_27421);
nand U28550 (N_28550,N_26251,N_27476);
and U28551 (N_28551,N_26241,N_27983);
or U28552 (N_28552,N_27661,N_27121);
nand U28553 (N_28553,N_27260,N_26016);
and U28554 (N_28554,N_27487,N_26560);
nand U28555 (N_28555,N_27320,N_27830);
and U28556 (N_28556,N_27646,N_27002);
and U28557 (N_28557,N_27457,N_27150);
and U28558 (N_28558,N_26535,N_26264);
nor U28559 (N_28559,N_26485,N_26342);
and U28560 (N_28560,N_26683,N_26463);
or U28561 (N_28561,N_26356,N_27618);
xnor U28562 (N_28562,N_26961,N_26769);
nor U28563 (N_28563,N_27752,N_26583);
nor U28564 (N_28564,N_27937,N_27869);
nand U28565 (N_28565,N_26641,N_27218);
nor U28566 (N_28566,N_26433,N_27696);
and U28567 (N_28567,N_26384,N_26466);
nand U28568 (N_28568,N_27017,N_26216);
or U28569 (N_28569,N_26289,N_26408);
nand U28570 (N_28570,N_26231,N_27879);
nand U28571 (N_28571,N_26975,N_26171);
nand U28572 (N_28572,N_26291,N_26078);
nor U28573 (N_28573,N_27188,N_26670);
and U28574 (N_28574,N_27902,N_27571);
nand U28575 (N_28575,N_27362,N_27789);
or U28576 (N_28576,N_26960,N_27245);
nand U28577 (N_28577,N_27040,N_27770);
nand U28578 (N_28578,N_27810,N_27518);
xor U28579 (N_28579,N_26067,N_27263);
and U28580 (N_28580,N_26616,N_26372);
or U28581 (N_28581,N_26756,N_27055);
or U28582 (N_28582,N_27021,N_27426);
and U28583 (N_28583,N_26260,N_26986);
and U28584 (N_28584,N_26551,N_27373);
or U28585 (N_28585,N_27463,N_26660);
and U28586 (N_28586,N_26283,N_26581);
and U28587 (N_28587,N_26146,N_26946);
nor U28588 (N_28588,N_27774,N_26239);
nor U28589 (N_28589,N_27991,N_27627);
xor U28590 (N_28590,N_26828,N_27926);
and U28591 (N_28591,N_27650,N_27032);
or U28592 (N_28592,N_27460,N_26182);
or U28593 (N_28593,N_27268,N_27759);
or U28594 (N_28594,N_26390,N_27965);
nor U28595 (N_28595,N_27495,N_27611);
nand U28596 (N_28596,N_26863,N_27209);
nor U28597 (N_28597,N_26918,N_27519);
xnor U28598 (N_28598,N_26186,N_26620);
nand U28599 (N_28599,N_26103,N_27249);
or U28600 (N_28600,N_27708,N_26875);
xor U28601 (N_28601,N_26895,N_26582);
or U28602 (N_28602,N_26337,N_27201);
nor U28603 (N_28603,N_27751,N_26915);
and U28604 (N_28604,N_27980,N_27821);
nor U28605 (N_28605,N_26092,N_27729);
and U28606 (N_28606,N_26700,N_26234);
nand U28607 (N_28607,N_26492,N_27404);
xnor U28608 (N_28608,N_26432,N_27025);
nand U28609 (N_28609,N_26138,N_27535);
xor U28610 (N_28610,N_27905,N_26613);
and U28611 (N_28611,N_26469,N_27863);
and U28612 (N_28612,N_26253,N_27384);
or U28613 (N_28613,N_26377,N_27765);
or U28614 (N_28614,N_27814,N_27613);
nor U28615 (N_28615,N_26862,N_26458);
or U28616 (N_28616,N_26489,N_27041);
nand U28617 (N_28617,N_26268,N_27698);
nor U28618 (N_28618,N_26022,N_26904);
nand U28619 (N_28619,N_26994,N_27938);
nand U28620 (N_28620,N_26208,N_26791);
and U28621 (N_28621,N_26400,N_26728);
nor U28622 (N_28622,N_26467,N_27883);
or U28623 (N_28623,N_26360,N_27126);
xnor U28624 (N_28624,N_26750,N_26511);
xor U28625 (N_28625,N_27343,N_27464);
and U28626 (N_28626,N_27522,N_27250);
nor U28627 (N_28627,N_27718,N_26664);
or U28628 (N_28628,N_26409,N_27206);
xor U28629 (N_28629,N_27302,N_26741);
xor U28630 (N_28630,N_26760,N_26644);
and U28631 (N_28631,N_27371,N_26175);
xor U28632 (N_28632,N_27854,N_26924);
nor U28633 (N_28633,N_27122,N_26726);
and U28634 (N_28634,N_27513,N_26889);
and U28635 (N_28635,N_27688,N_27090);
nand U28636 (N_28636,N_27957,N_27750);
or U28637 (N_28637,N_26352,N_27919);
nand U28638 (N_28638,N_27252,N_26397);
and U28639 (N_28639,N_27446,N_27078);
nand U28640 (N_28640,N_26671,N_27425);
and U28641 (N_28641,N_26605,N_27360);
and U28642 (N_28642,N_27336,N_26445);
or U28643 (N_28643,N_26490,N_27405);
or U28644 (N_28644,N_26520,N_26676);
nor U28645 (N_28645,N_26584,N_27995);
and U28646 (N_28646,N_27524,N_26831);
xnor U28647 (N_28647,N_26221,N_27038);
nor U28648 (N_28648,N_27313,N_27153);
nand U28649 (N_28649,N_26313,N_27195);
nor U28650 (N_28650,N_27636,N_26787);
nor U28651 (N_28651,N_26088,N_26245);
nand U28652 (N_28652,N_26443,N_26872);
nand U28653 (N_28653,N_27768,N_26265);
xnor U28654 (N_28654,N_27645,N_26884);
and U28655 (N_28655,N_27142,N_26134);
xor U28656 (N_28656,N_26883,N_27092);
and U28657 (N_28657,N_27443,N_26179);
nor U28658 (N_28658,N_26482,N_26349);
xor U28659 (N_28659,N_27106,N_27884);
and U28660 (N_28660,N_26153,N_27496);
or U28661 (N_28661,N_27947,N_26003);
and U28662 (N_28662,N_27439,N_26529);
or U28663 (N_28663,N_27619,N_26281);
or U28664 (N_28664,N_27062,N_26569);
nand U28665 (N_28665,N_27895,N_27146);
nor U28666 (N_28666,N_26880,N_27435);
nand U28667 (N_28667,N_27309,N_26840);
xnor U28668 (N_28668,N_27385,N_26453);
and U28669 (N_28669,N_27664,N_27632);
and U28670 (N_28670,N_27077,N_26890);
or U28671 (N_28671,N_26846,N_27408);
and U28672 (N_28672,N_27793,N_26966);
and U28673 (N_28673,N_26412,N_26881);
and U28674 (N_28674,N_26823,N_26942);
nand U28675 (N_28675,N_26579,N_26098);
nand U28676 (N_28676,N_27825,N_27045);
or U28677 (N_28677,N_27491,N_27160);
xnor U28678 (N_28678,N_26256,N_27876);
and U28679 (N_28679,N_26900,N_27266);
or U28680 (N_28680,N_27612,N_26233);
or U28681 (N_28681,N_26491,N_26326);
nand U28682 (N_28682,N_26287,N_26112);
nor U28683 (N_28683,N_27562,N_26922);
nor U28684 (N_28684,N_26647,N_26902);
or U28685 (N_28685,N_26794,N_26586);
nand U28686 (N_28686,N_26805,N_27262);
or U28687 (N_28687,N_27797,N_26131);
xnor U28688 (N_28688,N_26015,N_27207);
or U28689 (N_28689,N_27906,N_26226);
or U28690 (N_28690,N_26005,N_27583);
nor U28691 (N_28691,N_26835,N_27838);
xnor U28692 (N_28692,N_27946,N_27624);
or U28693 (N_28693,N_26748,N_27723);
xor U28694 (N_28694,N_26655,N_26323);
xor U28695 (N_28695,N_26544,N_26943);
nor U28696 (N_28696,N_27163,N_27639);
nand U28697 (N_28697,N_27907,N_26907);
xor U28698 (N_28698,N_27560,N_27029);
nand U28699 (N_28699,N_27120,N_27858);
xor U28700 (N_28700,N_27265,N_26451);
nand U28701 (N_28701,N_26766,N_27015);
xor U28702 (N_28702,N_27023,N_27786);
nor U28703 (N_28703,N_27475,N_27855);
xnor U28704 (N_28704,N_26438,N_27047);
and U28705 (N_28705,N_27130,N_27348);
xor U28706 (N_28706,N_27748,N_27471);
nor U28707 (N_28707,N_26479,N_26197);
or U28708 (N_28708,N_26176,N_26087);
or U28709 (N_28709,N_26820,N_27726);
and U28710 (N_28710,N_26106,N_27955);
xnor U28711 (N_28711,N_27745,N_26659);
or U28712 (N_28712,N_27375,N_26178);
or U28713 (N_28713,N_26648,N_26931);
and U28714 (N_28714,N_26508,N_26721);
or U28715 (N_28715,N_27916,N_26023);
nand U28716 (N_28716,N_27566,N_27803);
nor U28717 (N_28717,N_27380,N_27104);
xnor U28718 (N_28718,N_27248,N_26992);
nor U28719 (N_28719,N_27026,N_27473);
nand U28720 (N_28720,N_27894,N_26554);
nor U28721 (N_28721,N_26826,N_26874);
and U28722 (N_28722,N_26367,N_26751);
or U28723 (N_28723,N_26706,N_27577);
and U28724 (N_28724,N_27284,N_26174);
or U28725 (N_28725,N_26940,N_26180);
xnor U28726 (N_28726,N_27572,N_27526);
nor U28727 (N_28727,N_26220,N_27208);
nor U28728 (N_28728,N_27347,N_27187);
nor U28729 (N_28729,N_26737,N_27097);
and U28730 (N_28730,N_27235,N_27546);
nand U28731 (N_28731,N_27979,N_27081);
nor U28732 (N_28732,N_26478,N_26063);
and U28733 (N_28733,N_27601,N_27655);
or U28734 (N_28734,N_26068,N_27598);
and U28735 (N_28735,N_26484,N_27710);
xor U28736 (N_28736,N_26147,N_27840);
or U28737 (N_28737,N_26122,N_26450);
nand U28738 (N_28738,N_26666,N_26968);
and U28739 (N_28739,N_27363,N_27823);
xor U28740 (N_28740,N_27588,N_27323);
xnor U28741 (N_28741,N_26596,N_26389);
nor U28742 (N_28742,N_26189,N_26866);
or U28743 (N_28743,N_26825,N_26574);
or U28744 (N_28744,N_27203,N_26698);
or U28745 (N_28745,N_26177,N_26953);
nand U28746 (N_28746,N_26230,N_26685);
and U28747 (N_28747,N_26354,N_27826);
or U28748 (N_28748,N_27019,N_27254);
or U28749 (N_28749,N_26653,N_26150);
or U28750 (N_28750,N_27606,N_26546);
nand U28751 (N_28751,N_26795,N_26483);
nand U28752 (N_28752,N_26743,N_27456);
and U28753 (N_28753,N_27972,N_27339);
xor U28754 (N_28754,N_26448,N_27059);
xnor U28755 (N_28755,N_27179,N_27232);
and U28756 (N_28756,N_27470,N_27367);
nor U28757 (N_28757,N_26575,N_27539);
nand U28758 (N_28758,N_26868,N_26303);
nor U28759 (N_28759,N_26913,N_26156);
or U28760 (N_28760,N_27846,N_26494);
nand U28761 (N_28761,N_26454,N_26345);
xnor U28762 (N_28762,N_26925,N_27324);
and U28763 (N_28763,N_26169,N_26738);
nand U28764 (N_28764,N_27085,N_27802);
xor U28765 (N_28765,N_27417,N_27685);
xnor U28766 (N_28766,N_27118,N_26238);
or U28767 (N_28767,N_27466,N_27176);
and U28768 (N_28768,N_26978,N_27531);
and U28769 (N_28769,N_27239,N_26773);
xor U28770 (N_28770,N_26725,N_26468);
and U28771 (N_28771,N_27529,N_26425);
and U28772 (N_28772,N_26424,N_27180);
nor U28773 (N_28773,N_26568,N_26695);
nand U28774 (N_28774,N_27161,N_27434);
or U28775 (N_28775,N_27332,N_27603);
or U28776 (N_28776,N_26724,N_27630);
and U28777 (N_28777,N_26905,N_27808);
nand U28778 (N_28778,N_26764,N_27316);
or U28779 (N_28779,N_27364,N_26714);
xnor U28780 (N_28780,N_26813,N_26923);
or U28781 (N_28781,N_26762,N_26334);
nor U28782 (N_28782,N_26421,N_27771);
xnor U28783 (N_28783,N_27422,N_27671);
and U28784 (N_28784,N_26166,N_27898);
nand U28785 (N_28785,N_27781,N_27843);
and U28786 (N_28786,N_27857,N_27935);
and U28787 (N_28787,N_27193,N_26152);
or U28788 (N_28788,N_27874,N_26532);
nor U28789 (N_28789,N_27648,N_27686);
nand U28790 (N_28790,N_26937,N_27649);
or U28791 (N_28791,N_27345,N_27353);
and U28792 (N_28792,N_26537,N_26311);
nor U28793 (N_28793,N_26578,N_27192);
nor U28794 (N_28794,N_27447,N_27311);
nor U28795 (N_28795,N_26181,N_27773);
nor U28796 (N_28796,N_27074,N_27396);
nand U28797 (N_28797,N_27944,N_26870);
nor U28798 (N_28798,N_26767,N_26804);
nand U28799 (N_28799,N_27556,N_26563);
or U28800 (N_28800,N_27157,N_27914);
xnor U28801 (N_28801,N_27640,N_26462);
or U28802 (N_28802,N_26318,N_26643);
xnor U28803 (N_28803,N_26736,N_26752);
nand U28804 (N_28804,N_27833,N_27278);
nand U28805 (N_28805,N_27887,N_26600);
xor U28806 (N_28806,N_26102,N_27756);
or U28807 (N_28807,N_27829,N_27392);
or U28808 (N_28808,N_26222,N_26072);
or U28809 (N_28809,N_27676,N_27724);
and U28810 (N_28810,N_26612,N_27807);
nor U28811 (N_28811,N_26786,N_26404);
nand U28812 (N_28812,N_27253,N_26162);
or U28813 (N_28813,N_26252,N_27574);
or U28814 (N_28814,N_26686,N_27584);
nor U28815 (N_28815,N_26487,N_26949);
xor U28816 (N_28816,N_26788,N_27103);
xor U28817 (N_28817,N_27968,N_26499);
nand U28818 (N_28818,N_26396,N_27225);
nor U28819 (N_28819,N_26733,N_27327);
or U28820 (N_28820,N_26034,N_26246);
and U28821 (N_28821,N_26170,N_27665);
xnor U28822 (N_28822,N_27578,N_26065);
nor U28823 (N_28823,N_26219,N_26375);
xor U28824 (N_28824,N_27374,N_27743);
or U28825 (N_28825,N_26271,N_26476);
and U28826 (N_28826,N_26930,N_26510);
and U28827 (N_28827,N_26672,N_27912);
or U28828 (N_28828,N_27653,N_27486);
and U28829 (N_28829,N_26789,N_26027);
or U28830 (N_28830,N_26774,N_27692);
and U28831 (N_28831,N_26534,N_26442);
nand U28832 (N_28832,N_27540,N_26008);
xnor U28833 (N_28833,N_27525,N_27733);
xor U28834 (N_28834,N_26121,N_27592);
and U28835 (N_28835,N_27591,N_27004);
nand U28836 (N_28836,N_27398,N_27148);
and U28837 (N_28837,N_27662,N_27304);
nand U28838 (N_28838,N_27477,N_26770);
xor U28839 (N_28839,N_27228,N_26668);
xnor U28840 (N_28840,N_27959,N_26976);
xnor U28841 (N_28841,N_26095,N_26168);
nand U28842 (N_28842,N_26101,N_27282);
xnor U28843 (N_28843,N_26587,N_27194);
and U28844 (N_28844,N_27890,N_27185);
xor U28845 (N_28845,N_27511,N_27359);
xnor U28846 (N_28846,N_27811,N_27277);
or U28847 (N_28847,N_27933,N_27489);
nor U28848 (N_28848,N_27882,N_27500);
nand U28849 (N_28849,N_26627,N_26842);
xnor U28850 (N_28850,N_27711,N_26507);
xor U28851 (N_28851,N_27493,N_27701);
nand U28852 (N_28852,N_27865,N_26371);
or U28853 (N_28853,N_26035,N_26465);
and U28854 (N_28854,N_26044,N_26004);
nor U28855 (N_28855,N_27387,N_27140);
xor U28856 (N_28856,N_27728,N_27358);
and U28857 (N_28857,N_26920,N_27740);
and U28858 (N_28858,N_26669,N_27775);
or U28859 (N_28859,N_26628,N_27166);
nor U28860 (N_28860,N_26984,N_27969);
or U28861 (N_28861,N_27399,N_26309);
nand U28862 (N_28862,N_26461,N_27758);
or U28863 (N_28863,N_27217,N_27143);
or U28864 (N_28864,N_27427,N_26577);
or U28865 (N_28865,N_26187,N_26912);
or U28866 (N_28866,N_27181,N_27394);
and U28867 (N_28867,N_27593,N_26945);
nor U28868 (N_28868,N_26255,N_26370);
or U28869 (N_28869,N_27423,N_26267);
nor U28870 (N_28870,N_27340,N_27441);
or U28871 (N_28871,N_27100,N_26832);
nand U28872 (N_28872,N_26539,N_27834);
nor U28873 (N_28873,N_26663,N_27298);
and U28874 (N_28874,N_27764,N_26658);
nor U28875 (N_28875,N_27547,N_27076);
and U28876 (N_28876,N_26860,N_27301);
nor U28877 (N_28877,N_27776,N_27051);
and U28878 (N_28878,N_27133,N_27596);
nand U28879 (N_28879,N_26830,N_26709);
nand U28880 (N_28880,N_27356,N_26090);
or U28881 (N_28881,N_27237,N_26452);
or U28882 (N_28882,N_26885,N_26339);
nor U28883 (N_28883,N_27409,N_27954);
or U28884 (N_28884,N_27290,N_26172);
nor U28885 (N_28885,N_26277,N_27856);
xor U28886 (N_28886,N_27542,N_26204);
or U28887 (N_28887,N_27416,N_26525);
nor U28888 (N_28888,N_27617,N_27984);
xnor U28889 (N_28889,N_26274,N_26775);
or U28890 (N_28890,N_26173,N_26280);
nor U28891 (N_28891,N_26891,N_27845);
xor U28892 (N_28892,N_27739,N_26201);
nor U28893 (N_28893,N_26100,N_27070);
nand U28894 (N_28894,N_26218,N_27568);
nor U28895 (N_28895,N_27190,N_27828);
nand U28896 (N_28896,N_26436,N_26331);
and U28897 (N_28897,N_27541,N_26639);
or U28898 (N_28898,N_27697,N_27438);
or U28899 (N_28899,N_26861,N_27310);
nor U28900 (N_28900,N_27223,N_27129);
nor U28901 (N_28901,N_27967,N_26340);
or U28902 (N_28902,N_26618,N_27942);
nand U28903 (N_28903,N_26673,N_26956);
and U28904 (N_28904,N_27110,N_27549);
and U28905 (N_28905,N_27233,N_26636);
and U28906 (N_28906,N_26559,N_27900);
xor U28907 (N_28907,N_26190,N_26742);
nor U28908 (N_28908,N_27706,N_26164);
nand U28909 (N_28909,N_26080,N_27485);
nor U28910 (N_28910,N_27273,N_27280);
nor U28911 (N_28911,N_26501,N_27918);
xor U28912 (N_28912,N_27989,N_26934);
and U28913 (N_28913,N_27927,N_26935);
and U28914 (N_28914,N_27544,N_27276);
and U28915 (N_28915,N_26932,N_26132);
xnor U28916 (N_28916,N_27602,N_27660);
nand U28917 (N_28917,N_26497,N_26369);
and U28918 (N_28918,N_27520,N_26107);
nor U28919 (N_28919,N_26777,N_26983);
xnor U28920 (N_28920,N_27044,N_27079);
nand U28921 (N_28921,N_27850,N_26407);
xor U28922 (N_28922,N_26042,N_26060);
xnor U28923 (N_28923,N_27144,N_26727);
and U28924 (N_28924,N_26827,N_27494);
and U28925 (N_28925,N_26290,N_27971);
or U28926 (N_28926,N_27913,N_27720);
or U28927 (N_28927,N_26322,N_27080);
or U28928 (N_28928,N_26266,N_27490);
xnor U28929 (N_28929,N_26637,N_27691);
xor U28930 (N_28930,N_26944,N_27432);
or U28931 (N_28931,N_26348,N_27231);
or U28932 (N_28932,N_26689,N_26552);
nand U28933 (N_28933,N_26969,N_27344);
or U28934 (N_28934,N_27087,N_26545);
nand U28935 (N_28935,N_26097,N_27224);
xor U28936 (N_28936,N_27082,N_27703);
or U28937 (N_28937,N_27431,N_26897);
and U28938 (N_28938,N_27790,N_27109);
xor U28939 (N_28939,N_26071,N_26595);
and U28940 (N_28940,N_26675,N_26715);
nor U28941 (N_28941,N_26163,N_26385);
and U28942 (N_28942,N_27286,N_27338);
and U28943 (N_28943,N_27481,N_26437);
nand U28944 (N_28944,N_26703,N_27329);
and U28945 (N_28945,N_27177,N_26646);
nor U28946 (N_28946,N_27321,N_27200);
xor U28947 (N_28947,N_27683,N_26387);
nand U28948 (N_28948,N_27156,N_27822);
or U28949 (N_28949,N_26395,N_26898);
nand U28950 (N_28950,N_26667,N_27507);
and U28951 (N_28951,N_27669,N_26495);
and U28952 (N_28952,N_27626,N_27451);
xnor U28953 (N_28953,N_26470,N_27247);
or U28954 (N_28954,N_27221,N_27453);
nand U28955 (N_28955,N_26013,N_26856);
nand U28956 (N_28956,N_26142,N_26477);
nor U28957 (N_28957,N_27111,N_26428);
and U28958 (N_28958,N_26745,N_26378);
or U28959 (N_28959,N_27563,N_27368);
xnor U28960 (N_28960,N_26917,N_26558);
xnor U28961 (N_28961,N_26516,N_27687);
and U28962 (N_28962,N_27238,N_27005);
nor U28963 (N_28963,N_26621,N_27255);
nand U28964 (N_28964,N_26876,N_27357);
nand U28965 (N_28965,N_26592,N_26610);
xnor U28966 (N_28966,N_26800,N_27659);
nand U28967 (N_28967,N_26247,N_27977);
nor U28968 (N_28968,N_26020,N_26391);
and U28969 (N_28969,N_26140,N_26120);
or U28970 (N_28970,N_26278,N_27643);
nand U28971 (N_28971,N_27429,N_27573);
nor U28972 (N_28972,N_26185,N_26635);
nor U28973 (N_28973,N_26316,N_27242);
nor U28974 (N_28974,N_27020,N_26971);
nor U28975 (N_28975,N_26332,N_26141);
and U28976 (N_28976,N_27391,N_26273);
or U28977 (N_28977,N_27893,N_27105);
and U28978 (N_28978,N_27820,N_27975);
nand U28979 (N_28979,N_27170,N_27831);
nor U28980 (N_28980,N_26298,N_27377);
nor U28981 (N_28981,N_27885,N_26135);
xnor U28982 (N_28982,N_26036,N_27437);
or U28983 (N_28983,N_27575,N_26325);
xor U28984 (N_28984,N_26987,N_27742);
nor U28985 (N_28985,N_26205,N_27482);
nand U28986 (N_28986,N_26679,N_26328);
nor U28987 (N_28987,N_27480,N_27851);
or U28988 (N_28988,N_27303,N_27376);
and U28989 (N_28989,N_26307,N_26533);
nor U28990 (N_28990,N_26515,N_27430);
nand U28991 (N_28991,N_26650,N_27370);
xnor U28992 (N_28992,N_26446,N_26888);
xor U28993 (N_28993,N_27940,N_27297);
and U28994 (N_28994,N_27175,N_27410);
and U28995 (N_28995,N_27576,N_27389);
and U28996 (N_28996,N_26224,N_26965);
and U28997 (N_28997,N_27292,N_26707);
or U28998 (N_28998,N_26128,N_27700);
nor U28999 (N_28999,N_26697,N_27440);
and U29000 (N_29000,N_26422,N_26702);
nand U29001 (N_29001,N_26124,N_26325);
and U29002 (N_29002,N_27486,N_26626);
xnor U29003 (N_29003,N_26078,N_27331);
and U29004 (N_29004,N_27804,N_27537);
and U29005 (N_29005,N_26213,N_27435);
and U29006 (N_29006,N_26891,N_27292);
nand U29007 (N_29007,N_27879,N_26619);
or U29008 (N_29008,N_26750,N_27772);
xor U29009 (N_29009,N_26409,N_26254);
nand U29010 (N_29010,N_26774,N_27127);
nor U29011 (N_29011,N_26615,N_26224);
xor U29012 (N_29012,N_27021,N_27816);
xnor U29013 (N_29013,N_26856,N_27556);
nand U29014 (N_29014,N_27165,N_26822);
xor U29015 (N_29015,N_27773,N_26886);
nor U29016 (N_29016,N_26401,N_27279);
and U29017 (N_29017,N_26740,N_26760);
nor U29018 (N_29018,N_27641,N_26840);
nand U29019 (N_29019,N_26481,N_27687);
nand U29020 (N_29020,N_26275,N_26181);
or U29021 (N_29021,N_26243,N_26779);
nor U29022 (N_29022,N_27935,N_26220);
xnor U29023 (N_29023,N_27058,N_26486);
nor U29024 (N_29024,N_26222,N_26518);
xnor U29025 (N_29025,N_27793,N_27205);
nand U29026 (N_29026,N_27259,N_27106);
nand U29027 (N_29027,N_26231,N_26132);
or U29028 (N_29028,N_26536,N_26100);
and U29029 (N_29029,N_26637,N_27212);
nand U29030 (N_29030,N_27633,N_26104);
nand U29031 (N_29031,N_27091,N_26625);
xnor U29032 (N_29032,N_27888,N_27519);
nand U29033 (N_29033,N_27320,N_27373);
xnor U29034 (N_29034,N_26675,N_27440);
xor U29035 (N_29035,N_27245,N_26773);
xor U29036 (N_29036,N_26825,N_26555);
xnor U29037 (N_29037,N_26320,N_27460);
xnor U29038 (N_29038,N_26191,N_27959);
and U29039 (N_29039,N_27519,N_26300);
or U29040 (N_29040,N_27432,N_26053);
nand U29041 (N_29041,N_26471,N_27671);
and U29042 (N_29042,N_27726,N_27457);
nor U29043 (N_29043,N_26399,N_26695);
or U29044 (N_29044,N_26513,N_26056);
xnor U29045 (N_29045,N_27394,N_27361);
nand U29046 (N_29046,N_26946,N_26291);
or U29047 (N_29047,N_26410,N_26057);
and U29048 (N_29048,N_26490,N_27663);
nor U29049 (N_29049,N_26948,N_27909);
xor U29050 (N_29050,N_26241,N_26886);
xnor U29051 (N_29051,N_26982,N_27946);
xor U29052 (N_29052,N_27832,N_26065);
or U29053 (N_29053,N_27303,N_27891);
xnor U29054 (N_29054,N_27398,N_27900);
xor U29055 (N_29055,N_27027,N_27772);
xor U29056 (N_29056,N_27146,N_26018);
nand U29057 (N_29057,N_26543,N_27022);
xnor U29058 (N_29058,N_27557,N_27703);
and U29059 (N_29059,N_26505,N_26848);
nor U29060 (N_29060,N_26171,N_27109);
nor U29061 (N_29061,N_26210,N_27375);
xnor U29062 (N_29062,N_27079,N_27252);
nand U29063 (N_29063,N_26942,N_27860);
or U29064 (N_29064,N_26317,N_27182);
and U29065 (N_29065,N_27885,N_26069);
or U29066 (N_29066,N_27991,N_26629);
xnor U29067 (N_29067,N_26609,N_26821);
xnor U29068 (N_29068,N_27205,N_27425);
nor U29069 (N_29069,N_26697,N_27850);
nand U29070 (N_29070,N_27483,N_26689);
nand U29071 (N_29071,N_27639,N_27361);
nor U29072 (N_29072,N_26708,N_26125);
and U29073 (N_29073,N_26563,N_26000);
nand U29074 (N_29074,N_26642,N_26774);
nand U29075 (N_29075,N_27099,N_27097);
nor U29076 (N_29076,N_27416,N_27793);
or U29077 (N_29077,N_26442,N_27362);
and U29078 (N_29078,N_27569,N_27752);
or U29079 (N_29079,N_26451,N_27690);
and U29080 (N_29080,N_27790,N_27980);
xnor U29081 (N_29081,N_27169,N_26404);
xor U29082 (N_29082,N_27652,N_26554);
nor U29083 (N_29083,N_27839,N_27739);
nor U29084 (N_29084,N_27471,N_26809);
or U29085 (N_29085,N_27942,N_27776);
or U29086 (N_29086,N_26010,N_27044);
or U29087 (N_29087,N_27060,N_26233);
and U29088 (N_29088,N_26387,N_26802);
or U29089 (N_29089,N_27654,N_26787);
xnor U29090 (N_29090,N_26313,N_26272);
xor U29091 (N_29091,N_26214,N_27422);
xor U29092 (N_29092,N_27874,N_26228);
nand U29093 (N_29093,N_26558,N_26062);
or U29094 (N_29094,N_26225,N_26928);
nor U29095 (N_29095,N_27041,N_26635);
nand U29096 (N_29096,N_27470,N_27951);
xor U29097 (N_29097,N_26990,N_26670);
and U29098 (N_29098,N_27141,N_27891);
nor U29099 (N_29099,N_26351,N_26138);
and U29100 (N_29100,N_27946,N_26437);
and U29101 (N_29101,N_27185,N_27311);
and U29102 (N_29102,N_27289,N_26552);
nand U29103 (N_29103,N_27744,N_26760);
or U29104 (N_29104,N_27866,N_26327);
nand U29105 (N_29105,N_26053,N_27829);
or U29106 (N_29106,N_26637,N_26575);
and U29107 (N_29107,N_26540,N_27049);
nor U29108 (N_29108,N_27652,N_26647);
nand U29109 (N_29109,N_26772,N_26784);
nor U29110 (N_29110,N_27815,N_26499);
xnor U29111 (N_29111,N_27161,N_27491);
nand U29112 (N_29112,N_26526,N_26330);
and U29113 (N_29113,N_26304,N_27609);
nor U29114 (N_29114,N_26475,N_27255);
nor U29115 (N_29115,N_27759,N_26821);
nand U29116 (N_29116,N_27457,N_26842);
xor U29117 (N_29117,N_26603,N_26873);
and U29118 (N_29118,N_26846,N_26230);
nor U29119 (N_29119,N_26724,N_26554);
and U29120 (N_29120,N_26618,N_26191);
and U29121 (N_29121,N_26286,N_26514);
nor U29122 (N_29122,N_26815,N_27627);
xnor U29123 (N_29123,N_27695,N_26492);
nor U29124 (N_29124,N_27378,N_27547);
xor U29125 (N_29125,N_27646,N_26872);
nor U29126 (N_29126,N_27426,N_26758);
xor U29127 (N_29127,N_26840,N_27723);
xor U29128 (N_29128,N_26776,N_27348);
nor U29129 (N_29129,N_26843,N_26683);
nand U29130 (N_29130,N_27532,N_26575);
and U29131 (N_29131,N_26047,N_26306);
nand U29132 (N_29132,N_27943,N_27528);
and U29133 (N_29133,N_27984,N_26037);
xor U29134 (N_29134,N_27937,N_26774);
or U29135 (N_29135,N_26680,N_26758);
or U29136 (N_29136,N_26696,N_26614);
nor U29137 (N_29137,N_26112,N_26607);
and U29138 (N_29138,N_26243,N_27943);
nand U29139 (N_29139,N_27072,N_26719);
nand U29140 (N_29140,N_27260,N_26780);
nand U29141 (N_29141,N_27607,N_27631);
and U29142 (N_29142,N_26174,N_27772);
nor U29143 (N_29143,N_27692,N_26007);
or U29144 (N_29144,N_27946,N_26786);
xor U29145 (N_29145,N_27780,N_27565);
or U29146 (N_29146,N_27837,N_27220);
nand U29147 (N_29147,N_26727,N_27707);
or U29148 (N_29148,N_27711,N_27340);
nand U29149 (N_29149,N_26588,N_26677);
and U29150 (N_29150,N_27051,N_27731);
and U29151 (N_29151,N_26897,N_26509);
and U29152 (N_29152,N_27526,N_26389);
nor U29153 (N_29153,N_26526,N_26403);
and U29154 (N_29154,N_27352,N_26330);
or U29155 (N_29155,N_27310,N_27743);
nand U29156 (N_29156,N_26853,N_26941);
and U29157 (N_29157,N_26718,N_27589);
or U29158 (N_29158,N_27481,N_26447);
nor U29159 (N_29159,N_27196,N_27788);
nand U29160 (N_29160,N_27560,N_27319);
xnor U29161 (N_29161,N_26703,N_26860);
and U29162 (N_29162,N_26807,N_27264);
xnor U29163 (N_29163,N_27536,N_26614);
xnor U29164 (N_29164,N_26989,N_26311);
nor U29165 (N_29165,N_27611,N_27819);
or U29166 (N_29166,N_27678,N_26425);
nand U29167 (N_29167,N_27703,N_26061);
xnor U29168 (N_29168,N_27358,N_26575);
or U29169 (N_29169,N_27819,N_26713);
xor U29170 (N_29170,N_26888,N_26358);
or U29171 (N_29171,N_27754,N_26216);
or U29172 (N_29172,N_27640,N_27631);
nand U29173 (N_29173,N_26521,N_27196);
and U29174 (N_29174,N_27053,N_27737);
or U29175 (N_29175,N_27356,N_26080);
nor U29176 (N_29176,N_26133,N_26270);
nand U29177 (N_29177,N_27026,N_27215);
nor U29178 (N_29178,N_27927,N_27474);
xnor U29179 (N_29179,N_27590,N_26077);
or U29180 (N_29180,N_26467,N_27363);
and U29181 (N_29181,N_26385,N_27952);
or U29182 (N_29182,N_27134,N_26346);
nand U29183 (N_29183,N_27605,N_26319);
xor U29184 (N_29184,N_27853,N_26495);
nand U29185 (N_29185,N_26663,N_27547);
and U29186 (N_29186,N_26878,N_27560);
xor U29187 (N_29187,N_26847,N_27553);
or U29188 (N_29188,N_27879,N_27200);
or U29189 (N_29189,N_27138,N_27450);
and U29190 (N_29190,N_26897,N_27120);
and U29191 (N_29191,N_26395,N_26545);
or U29192 (N_29192,N_26437,N_26870);
xnor U29193 (N_29193,N_26930,N_27127);
xnor U29194 (N_29194,N_27231,N_27580);
xnor U29195 (N_29195,N_27299,N_27525);
nor U29196 (N_29196,N_27625,N_27448);
nor U29197 (N_29197,N_27898,N_27044);
xnor U29198 (N_29198,N_26070,N_27404);
or U29199 (N_29199,N_26764,N_26601);
or U29200 (N_29200,N_27899,N_26553);
nand U29201 (N_29201,N_27057,N_27018);
nand U29202 (N_29202,N_26855,N_27865);
xor U29203 (N_29203,N_26265,N_27727);
nand U29204 (N_29204,N_26151,N_27785);
and U29205 (N_29205,N_27000,N_26000);
nand U29206 (N_29206,N_26742,N_27295);
nand U29207 (N_29207,N_27740,N_26902);
and U29208 (N_29208,N_26860,N_27657);
nand U29209 (N_29209,N_27096,N_26568);
xnor U29210 (N_29210,N_27109,N_26653);
xor U29211 (N_29211,N_27199,N_26756);
or U29212 (N_29212,N_26739,N_26912);
nor U29213 (N_29213,N_26198,N_27411);
or U29214 (N_29214,N_27425,N_27347);
nand U29215 (N_29215,N_26773,N_27294);
and U29216 (N_29216,N_26772,N_26728);
nand U29217 (N_29217,N_27145,N_27787);
and U29218 (N_29218,N_26198,N_27109);
nor U29219 (N_29219,N_26794,N_27113);
or U29220 (N_29220,N_26280,N_27829);
and U29221 (N_29221,N_26711,N_27570);
nand U29222 (N_29222,N_27201,N_26604);
nor U29223 (N_29223,N_26659,N_26515);
and U29224 (N_29224,N_26029,N_27810);
and U29225 (N_29225,N_27537,N_26440);
and U29226 (N_29226,N_26660,N_26462);
or U29227 (N_29227,N_27070,N_27143);
and U29228 (N_29228,N_26232,N_26975);
nor U29229 (N_29229,N_27132,N_26422);
nor U29230 (N_29230,N_26045,N_26314);
and U29231 (N_29231,N_27877,N_27191);
nor U29232 (N_29232,N_27410,N_26342);
nand U29233 (N_29233,N_26955,N_27698);
or U29234 (N_29234,N_27554,N_26674);
or U29235 (N_29235,N_26795,N_26901);
and U29236 (N_29236,N_26147,N_26467);
nand U29237 (N_29237,N_27448,N_26679);
or U29238 (N_29238,N_27804,N_27665);
or U29239 (N_29239,N_26153,N_27922);
or U29240 (N_29240,N_26710,N_26421);
or U29241 (N_29241,N_27991,N_27787);
nand U29242 (N_29242,N_26022,N_27364);
nor U29243 (N_29243,N_27462,N_27563);
or U29244 (N_29244,N_26269,N_26588);
nor U29245 (N_29245,N_27269,N_26778);
or U29246 (N_29246,N_27985,N_26646);
nor U29247 (N_29247,N_26415,N_27228);
nor U29248 (N_29248,N_26068,N_26157);
or U29249 (N_29249,N_27848,N_26472);
and U29250 (N_29250,N_27117,N_27104);
nor U29251 (N_29251,N_27316,N_27843);
nor U29252 (N_29252,N_26046,N_26261);
xor U29253 (N_29253,N_26351,N_27209);
or U29254 (N_29254,N_26606,N_26366);
or U29255 (N_29255,N_27524,N_26726);
nand U29256 (N_29256,N_26731,N_26836);
and U29257 (N_29257,N_27961,N_26789);
xnor U29258 (N_29258,N_26469,N_26486);
nand U29259 (N_29259,N_26065,N_27283);
or U29260 (N_29260,N_27879,N_27247);
or U29261 (N_29261,N_26592,N_27198);
xor U29262 (N_29262,N_27128,N_26732);
xnor U29263 (N_29263,N_27533,N_27549);
nand U29264 (N_29264,N_27281,N_26510);
nor U29265 (N_29265,N_27802,N_26145);
nor U29266 (N_29266,N_27540,N_26244);
nand U29267 (N_29267,N_26021,N_26173);
or U29268 (N_29268,N_26288,N_26212);
nor U29269 (N_29269,N_27877,N_27406);
nand U29270 (N_29270,N_26582,N_26298);
nand U29271 (N_29271,N_26375,N_26848);
and U29272 (N_29272,N_26825,N_27011);
nand U29273 (N_29273,N_26029,N_26126);
nand U29274 (N_29274,N_26566,N_27304);
xnor U29275 (N_29275,N_26485,N_27502);
nor U29276 (N_29276,N_26638,N_26583);
xnor U29277 (N_29277,N_27803,N_27607);
xnor U29278 (N_29278,N_26129,N_27763);
and U29279 (N_29279,N_26206,N_27501);
or U29280 (N_29280,N_27043,N_27954);
or U29281 (N_29281,N_26816,N_26681);
or U29282 (N_29282,N_26520,N_26490);
and U29283 (N_29283,N_26100,N_26429);
nor U29284 (N_29284,N_27453,N_26694);
and U29285 (N_29285,N_26628,N_26726);
nor U29286 (N_29286,N_27383,N_27194);
nand U29287 (N_29287,N_26734,N_26044);
and U29288 (N_29288,N_27338,N_27724);
nand U29289 (N_29289,N_26201,N_27365);
xor U29290 (N_29290,N_26871,N_26601);
xnor U29291 (N_29291,N_27712,N_26498);
or U29292 (N_29292,N_27358,N_27710);
nand U29293 (N_29293,N_26775,N_27410);
xnor U29294 (N_29294,N_27064,N_27747);
nor U29295 (N_29295,N_26499,N_27177);
xor U29296 (N_29296,N_27701,N_27090);
and U29297 (N_29297,N_26250,N_27146);
xor U29298 (N_29298,N_27908,N_26177);
xor U29299 (N_29299,N_27836,N_26373);
or U29300 (N_29300,N_26451,N_27845);
nor U29301 (N_29301,N_27424,N_27481);
and U29302 (N_29302,N_27350,N_27701);
or U29303 (N_29303,N_26777,N_26598);
nor U29304 (N_29304,N_27646,N_27602);
nor U29305 (N_29305,N_27679,N_26775);
xor U29306 (N_29306,N_27143,N_26429);
or U29307 (N_29307,N_26726,N_26641);
xor U29308 (N_29308,N_26562,N_27587);
xor U29309 (N_29309,N_26212,N_26446);
nor U29310 (N_29310,N_27803,N_26990);
or U29311 (N_29311,N_26250,N_26612);
or U29312 (N_29312,N_26820,N_27916);
nor U29313 (N_29313,N_26271,N_26842);
and U29314 (N_29314,N_27521,N_26832);
and U29315 (N_29315,N_27122,N_27379);
nor U29316 (N_29316,N_26220,N_26981);
and U29317 (N_29317,N_27019,N_26934);
xnor U29318 (N_29318,N_27764,N_26919);
or U29319 (N_29319,N_27608,N_26572);
xnor U29320 (N_29320,N_26947,N_26144);
xor U29321 (N_29321,N_26967,N_26904);
or U29322 (N_29322,N_26585,N_27198);
nand U29323 (N_29323,N_27618,N_26052);
nand U29324 (N_29324,N_26018,N_27818);
xor U29325 (N_29325,N_27271,N_26523);
and U29326 (N_29326,N_26508,N_26789);
or U29327 (N_29327,N_26982,N_27408);
nor U29328 (N_29328,N_27870,N_26125);
or U29329 (N_29329,N_27224,N_26857);
and U29330 (N_29330,N_27643,N_26175);
and U29331 (N_29331,N_26119,N_27963);
xnor U29332 (N_29332,N_27788,N_27946);
xor U29333 (N_29333,N_27942,N_26326);
xnor U29334 (N_29334,N_26943,N_26471);
or U29335 (N_29335,N_26875,N_26640);
nor U29336 (N_29336,N_27993,N_26804);
xnor U29337 (N_29337,N_27896,N_27827);
xor U29338 (N_29338,N_27971,N_26629);
xnor U29339 (N_29339,N_27138,N_26081);
and U29340 (N_29340,N_26807,N_27378);
or U29341 (N_29341,N_27496,N_26680);
or U29342 (N_29342,N_26888,N_27405);
nor U29343 (N_29343,N_26939,N_27464);
xnor U29344 (N_29344,N_26538,N_27751);
nand U29345 (N_29345,N_27234,N_26173);
and U29346 (N_29346,N_27985,N_26558);
nor U29347 (N_29347,N_26196,N_27948);
and U29348 (N_29348,N_27360,N_26564);
or U29349 (N_29349,N_27173,N_27826);
nand U29350 (N_29350,N_27210,N_26492);
or U29351 (N_29351,N_27629,N_27143);
and U29352 (N_29352,N_27470,N_26849);
xor U29353 (N_29353,N_26103,N_27928);
nor U29354 (N_29354,N_26217,N_26644);
nor U29355 (N_29355,N_27450,N_27231);
nor U29356 (N_29356,N_27228,N_26358);
or U29357 (N_29357,N_27177,N_26572);
and U29358 (N_29358,N_27067,N_27982);
or U29359 (N_29359,N_27212,N_26766);
or U29360 (N_29360,N_27873,N_26034);
nand U29361 (N_29361,N_27881,N_27581);
nand U29362 (N_29362,N_27619,N_26383);
nor U29363 (N_29363,N_27313,N_26806);
and U29364 (N_29364,N_27246,N_27560);
or U29365 (N_29365,N_26985,N_27072);
xnor U29366 (N_29366,N_26351,N_27223);
xnor U29367 (N_29367,N_27026,N_27689);
xor U29368 (N_29368,N_26207,N_26968);
xnor U29369 (N_29369,N_26502,N_26029);
xnor U29370 (N_29370,N_26430,N_27551);
nor U29371 (N_29371,N_27381,N_27633);
xor U29372 (N_29372,N_26512,N_27901);
xor U29373 (N_29373,N_26090,N_26571);
nand U29374 (N_29374,N_27807,N_27711);
and U29375 (N_29375,N_27689,N_27924);
nor U29376 (N_29376,N_26552,N_26754);
nor U29377 (N_29377,N_27832,N_27597);
nand U29378 (N_29378,N_26735,N_27894);
nor U29379 (N_29379,N_27282,N_27508);
nor U29380 (N_29380,N_27760,N_26054);
or U29381 (N_29381,N_26992,N_26309);
nand U29382 (N_29382,N_27427,N_27551);
and U29383 (N_29383,N_27658,N_26597);
nand U29384 (N_29384,N_26255,N_27147);
nand U29385 (N_29385,N_26496,N_26500);
and U29386 (N_29386,N_26955,N_26344);
nand U29387 (N_29387,N_27075,N_27188);
nand U29388 (N_29388,N_26569,N_26891);
nand U29389 (N_29389,N_26948,N_27880);
xnor U29390 (N_29390,N_26044,N_27989);
nand U29391 (N_29391,N_26572,N_27525);
and U29392 (N_29392,N_26085,N_27869);
or U29393 (N_29393,N_27680,N_27329);
and U29394 (N_29394,N_26267,N_27558);
xor U29395 (N_29395,N_26699,N_26326);
and U29396 (N_29396,N_27378,N_26041);
or U29397 (N_29397,N_27891,N_27922);
and U29398 (N_29398,N_26762,N_26451);
nor U29399 (N_29399,N_26361,N_27294);
xor U29400 (N_29400,N_27385,N_27106);
nor U29401 (N_29401,N_26535,N_26532);
xor U29402 (N_29402,N_26610,N_27775);
nor U29403 (N_29403,N_27822,N_26675);
xor U29404 (N_29404,N_27736,N_27375);
nor U29405 (N_29405,N_26070,N_27364);
or U29406 (N_29406,N_26089,N_26555);
nand U29407 (N_29407,N_27149,N_27438);
or U29408 (N_29408,N_27043,N_26496);
and U29409 (N_29409,N_27310,N_26818);
nor U29410 (N_29410,N_26945,N_26566);
nand U29411 (N_29411,N_27314,N_27949);
nand U29412 (N_29412,N_27645,N_27945);
nand U29413 (N_29413,N_26876,N_26584);
or U29414 (N_29414,N_26610,N_26109);
nand U29415 (N_29415,N_27009,N_27646);
or U29416 (N_29416,N_26098,N_27971);
nor U29417 (N_29417,N_27489,N_26673);
xnor U29418 (N_29418,N_26800,N_27307);
and U29419 (N_29419,N_27442,N_26598);
xnor U29420 (N_29420,N_26060,N_27133);
and U29421 (N_29421,N_26847,N_27995);
or U29422 (N_29422,N_27396,N_26019);
nor U29423 (N_29423,N_26958,N_27486);
xor U29424 (N_29424,N_26847,N_26388);
nor U29425 (N_29425,N_27326,N_27230);
or U29426 (N_29426,N_26803,N_27220);
nand U29427 (N_29427,N_27247,N_27019);
or U29428 (N_29428,N_27640,N_27831);
nor U29429 (N_29429,N_26908,N_26413);
nand U29430 (N_29430,N_26023,N_26153);
or U29431 (N_29431,N_26775,N_26532);
nor U29432 (N_29432,N_26425,N_27299);
or U29433 (N_29433,N_26037,N_27637);
and U29434 (N_29434,N_26740,N_26192);
or U29435 (N_29435,N_26319,N_27308);
and U29436 (N_29436,N_27528,N_26242);
and U29437 (N_29437,N_27692,N_27114);
and U29438 (N_29438,N_27578,N_26149);
nand U29439 (N_29439,N_26203,N_27785);
xnor U29440 (N_29440,N_27451,N_27631);
and U29441 (N_29441,N_27287,N_26573);
nor U29442 (N_29442,N_27087,N_26498);
and U29443 (N_29443,N_26273,N_27666);
and U29444 (N_29444,N_27319,N_26548);
nor U29445 (N_29445,N_27833,N_26604);
nand U29446 (N_29446,N_27393,N_27166);
nor U29447 (N_29447,N_26649,N_27634);
nand U29448 (N_29448,N_27795,N_27967);
nor U29449 (N_29449,N_27534,N_27028);
nand U29450 (N_29450,N_27013,N_26363);
nor U29451 (N_29451,N_27807,N_26132);
or U29452 (N_29452,N_27677,N_27106);
xor U29453 (N_29453,N_26799,N_26922);
nand U29454 (N_29454,N_26546,N_27804);
nand U29455 (N_29455,N_26827,N_27973);
and U29456 (N_29456,N_26441,N_26715);
nand U29457 (N_29457,N_26887,N_27413);
xor U29458 (N_29458,N_26278,N_26639);
nand U29459 (N_29459,N_26368,N_26681);
and U29460 (N_29460,N_27921,N_26304);
nand U29461 (N_29461,N_26399,N_26405);
and U29462 (N_29462,N_26327,N_26929);
nor U29463 (N_29463,N_27111,N_26654);
xnor U29464 (N_29464,N_26543,N_27000);
nor U29465 (N_29465,N_26499,N_27870);
nand U29466 (N_29466,N_26323,N_26430);
nor U29467 (N_29467,N_27016,N_26706);
and U29468 (N_29468,N_26628,N_27174);
or U29469 (N_29469,N_27398,N_27844);
and U29470 (N_29470,N_27241,N_27658);
and U29471 (N_29471,N_26666,N_27214);
and U29472 (N_29472,N_27634,N_27574);
or U29473 (N_29473,N_27182,N_26931);
and U29474 (N_29474,N_27246,N_26810);
nor U29475 (N_29475,N_27002,N_27659);
nor U29476 (N_29476,N_26213,N_27284);
and U29477 (N_29477,N_26736,N_26601);
nand U29478 (N_29478,N_27431,N_27882);
nand U29479 (N_29479,N_27967,N_26324);
nand U29480 (N_29480,N_27198,N_26345);
nor U29481 (N_29481,N_27618,N_27504);
xor U29482 (N_29482,N_26869,N_26149);
nand U29483 (N_29483,N_26284,N_26729);
or U29484 (N_29484,N_26142,N_26894);
nand U29485 (N_29485,N_27289,N_27017);
nor U29486 (N_29486,N_27004,N_27762);
nor U29487 (N_29487,N_27253,N_26319);
xor U29488 (N_29488,N_26628,N_26985);
and U29489 (N_29489,N_27551,N_27544);
xor U29490 (N_29490,N_27544,N_26517);
nor U29491 (N_29491,N_27130,N_26541);
nand U29492 (N_29492,N_26109,N_27815);
xnor U29493 (N_29493,N_26927,N_27140);
or U29494 (N_29494,N_27730,N_27071);
xnor U29495 (N_29495,N_27470,N_26403);
nor U29496 (N_29496,N_27349,N_27541);
xor U29497 (N_29497,N_27055,N_27296);
nand U29498 (N_29498,N_27599,N_26424);
or U29499 (N_29499,N_26667,N_26937);
or U29500 (N_29500,N_26767,N_26792);
or U29501 (N_29501,N_27785,N_27348);
or U29502 (N_29502,N_27934,N_26623);
or U29503 (N_29503,N_27571,N_27798);
nand U29504 (N_29504,N_26261,N_26866);
or U29505 (N_29505,N_27943,N_26283);
xor U29506 (N_29506,N_26490,N_26657);
and U29507 (N_29507,N_26077,N_27973);
or U29508 (N_29508,N_26772,N_26961);
nor U29509 (N_29509,N_26362,N_27539);
nand U29510 (N_29510,N_27154,N_27273);
nor U29511 (N_29511,N_26184,N_26141);
and U29512 (N_29512,N_26315,N_26707);
xnor U29513 (N_29513,N_27986,N_26372);
or U29514 (N_29514,N_26792,N_27939);
nor U29515 (N_29515,N_27289,N_26964);
and U29516 (N_29516,N_27220,N_27887);
or U29517 (N_29517,N_27243,N_27533);
or U29518 (N_29518,N_26891,N_27023);
or U29519 (N_29519,N_27905,N_26336);
and U29520 (N_29520,N_27126,N_27979);
and U29521 (N_29521,N_27181,N_27164);
xnor U29522 (N_29522,N_27806,N_27603);
nor U29523 (N_29523,N_26224,N_27415);
nor U29524 (N_29524,N_27458,N_27732);
and U29525 (N_29525,N_26638,N_26207);
nand U29526 (N_29526,N_27312,N_26851);
nor U29527 (N_29527,N_26670,N_26215);
or U29528 (N_29528,N_27051,N_27822);
nand U29529 (N_29529,N_26491,N_27699);
xnor U29530 (N_29530,N_26240,N_26807);
xor U29531 (N_29531,N_27277,N_27112);
nor U29532 (N_29532,N_27808,N_26966);
and U29533 (N_29533,N_26753,N_26977);
or U29534 (N_29534,N_27465,N_26448);
nand U29535 (N_29535,N_27267,N_27640);
xnor U29536 (N_29536,N_27367,N_26185);
xnor U29537 (N_29537,N_26192,N_27501);
and U29538 (N_29538,N_26855,N_26077);
or U29539 (N_29539,N_26993,N_27973);
or U29540 (N_29540,N_27085,N_26949);
nor U29541 (N_29541,N_27681,N_27039);
xnor U29542 (N_29542,N_26919,N_27124);
or U29543 (N_29543,N_27946,N_27821);
nor U29544 (N_29544,N_26217,N_27835);
nand U29545 (N_29545,N_26365,N_27270);
or U29546 (N_29546,N_26409,N_27884);
and U29547 (N_29547,N_26251,N_26896);
nand U29548 (N_29548,N_26528,N_27230);
and U29549 (N_29549,N_26496,N_27928);
nand U29550 (N_29550,N_26535,N_26508);
and U29551 (N_29551,N_26098,N_27793);
and U29552 (N_29552,N_26989,N_26548);
nor U29553 (N_29553,N_26152,N_27663);
or U29554 (N_29554,N_26020,N_26852);
nor U29555 (N_29555,N_27978,N_26929);
nor U29556 (N_29556,N_27694,N_27275);
nor U29557 (N_29557,N_27857,N_27392);
or U29558 (N_29558,N_26276,N_26205);
and U29559 (N_29559,N_26920,N_26692);
nand U29560 (N_29560,N_26715,N_27269);
nor U29561 (N_29561,N_26118,N_27033);
or U29562 (N_29562,N_26969,N_27193);
nand U29563 (N_29563,N_26879,N_27306);
and U29564 (N_29564,N_26972,N_26767);
and U29565 (N_29565,N_27252,N_27617);
and U29566 (N_29566,N_27732,N_26921);
nand U29567 (N_29567,N_27610,N_27362);
and U29568 (N_29568,N_26975,N_26363);
xor U29569 (N_29569,N_26091,N_26082);
and U29570 (N_29570,N_26051,N_26098);
nand U29571 (N_29571,N_26930,N_26488);
or U29572 (N_29572,N_26492,N_27444);
or U29573 (N_29573,N_27026,N_26762);
nor U29574 (N_29574,N_27261,N_27297);
nand U29575 (N_29575,N_27641,N_26144);
or U29576 (N_29576,N_27844,N_26796);
or U29577 (N_29577,N_26122,N_26329);
nor U29578 (N_29578,N_27053,N_27997);
or U29579 (N_29579,N_26152,N_27628);
nor U29580 (N_29580,N_26955,N_26411);
and U29581 (N_29581,N_26029,N_26662);
or U29582 (N_29582,N_26032,N_26794);
nor U29583 (N_29583,N_26800,N_27058);
nor U29584 (N_29584,N_26797,N_27049);
or U29585 (N_29585,N_27047,N_26264);
xnor U29586 (N_29586,N_26527,N_26803);
or U29587 (N_29587,N_27753,N_27758);
xnor U29588 (N_29588,N_27629,N_27368);
xnor U29589 (N_29589,N_27869,N_26198);
and U29590 (N_29590,N_27502,N_27400);
or U29591 (N_29591,N_26872,N_27718);
and U29592 (N_29592,N_27444,N_27782);
or U29593 (N_29593,N_26896,N_26465);
xor U29594 (N_29594,N_26997,N_26167);
nor U29595 (N_29595,N_27546,N_26285);
xnor U29596 (N_29596,N_27968,N_27335);
or U29597 (N_29597,N_26127,N_27946);
and U29598 (N_29598,N_26306,N_26421);
nand U29599 (N_29599,N_26756,N_26387);
nor U29600 (N_29600,N_26989,N_26881);
and U29601 (N_29601,N_26764,N_26504);
and U29602 (N_29602,N_26266,N_27771);
nor U29603 (N_29603,N_26660,N_26876);
nor U29604 (N_29604,N_26889,N_27919);
xnor U29605 (N_29605,N_26047,N_27676);
nand U29606 (N_29606,N_27550,N_27992);
or U29607 (N_29607,N_26672,N_26217);
xor U29608 (N_29608,N_27174,N_27399);
and U29609 (N_29609,N_27921,N_27435);
nand U29610 (N_29610,N_27557,N_26251);
nand U29611 (N_29611,N_27897,N_27880);
or U29612 (N_29612,N_26437,N_27802);
nor U29613 (N_29613,N_26918,N_26979);
and U29614 (N_29614,N_26614,N_27698);
nand U29615 (N_29615,N_26346,N_26378);
and U29616 (N_29616,N_27877,N_27170);
and U29617 (N_29617,N_27389,N_26380);
nand U29618 (N_29618,N_26893,N_27286);
xnor U29619 (N_29619,N_26695,N_27419);
or U29620 (N_29620,N_26690,N_27708);
nand U29621 (N_29621,N_26611,N_27819);
xnor U29622 (N_29622,N_26331,N_27701);
nand U29623 (N_29623,N_26273,N_26250);
xnor U29624 (N_29624,N_27969,N_27526);
and U29625 (N_29625,N_27542,N_27641);
or U29626 (N_29626,N_27908,N_26178);
xor U29627 (N_29627,N_26481,N_27431);
and U29628 (N_29628,N_26055,N_27332);
nor U29629 (N_29629,N_27645,N_27734);
and U29630 (N_29630,N_26373,N_27352);
or U29631 (N_29631,N_26552,N_26472);
or U29632 (N_29632,N_26138,N_26793);
xor U29633 (N_29633,N_26945,N_26393);
or U29634 (N_29634,N_27107,N_26073);
xnor U29635 (N_29635,N_27536,N_27390);
and U29636 (N_29636,N_27781,N_27598);
xor U29637 (N_29637,N_27538,N_26161);
and U29638 (N_29638,N_27873,N_27345);
nand U29639 (N_29639,N_26597,N_26549);
or U29640 (N_29640,N_26352,N_26219);
nand U29641 (N_29641,N_27655,N_26509);
and U29642 (N_29642,N_26335,N_26204);
xnor U29643 (N_29643,N_26868,N_27435);
xnor U29644 (N_29644,N_27422,N_27979);
and U29645 (N_29645,N_26964,N_26243);
nor U29646 (N_29646,N_27327,N_26694);
xnor U29647 (N_29647,N_26500,N_26721);
xnor U29648 (N_29648,N_26675,N_26380);
and U29649 (N_29649,N_26649,N_26233);
nand U29650 (N_29650,N_27910,N_26565);
and U29651 (N_29651,N_26922,N_26380);
nand U29652 (N_29652,N_26011,N_27723);
nor U29653 (N_29653,N_26649,N_26330);
nand U29654 (N_29654,N_26670,N_26509);
nor U29655 (N_29655,N_26969,N_26254);
nand U29656 (N_29656,N_27232,N_27306);
nor U29657 (N_29657,N_26384,N_27378);
nand U29658 (N_29658,N_27638,N_27319);
xor U29659 (N_29659,N_26465,N_26440);
xor U29660 (N_29660,N_26524,N_26662);
nand U29661 (N_29661,N_27135,N_27140);
xnor U29662 (N_29662,N_27262,N_26910);
or U29663 (N_29663,N_26726,N_26213);
and U29664 (N_29664,N_27496,N_26193);
nand U29665 (N_29665,N_26151,N_27401);
and U29666 (N_29666,N_26038,N_27658);
nor U29667 (N_29667,N_26162,N_27634);
nor U29668 (N_29668,N_27172,N_26888);
and U29669 (N_29669,N_26061,N_26551);
or U29670 (N_29670,N_27251,N_26133);
nand U29671 (N_29671,N_26850,N_26952);
or U29672 (N_29672,N_26756,N_26517);
nor U29673 (N_29673,N_26434,N_26665);
nand U29674 (N_29674,N_26681,N_26785);
and U29675 (N_29675,N_26312,N_26715);
or U29676 (N_29676,N_26032,N_26817);
nand U29677 (N_29677,N_27813,N_26695);
or U29678 (N_29678,N_27920,N_26922);
and U29679 (N_29679,N_27091,N_26726);
nor U29680 (N_29680,N_27901,N_27169);
and U29681 (N_29681,N_26788,N_26682);
nand U29682 (N_29682,N_27271,N_26995);
nor U29683 (N_29683,N_26566,N_27654);
or U29684 (N_29684,N_27995,N_26549);
or U29685 (N_29685,N_26788,N_26562);
nor U29686 (N_29686,N_27829,N_27251);
or U29687 (N_29687,N_27692,N_27598);
and U29688 (N_29688,N_27443,N_26682);
and U29689 (N_29689,N_27191,N_27740);
nor U29690 (N_29690,N_26569,N_26147);
nand U29691 (N_29691,N_26767,N_27146);
nor U29692 (N_29692,N_27612,N_27422);
or U29693 (N_29693,N_27465,N_26298);
xnor U29694 (N_29694,N_27177,N_27667);
nor U29695 (N_29695,N_27958,N_26860);
nand U29696 (N_29696,N_26688,N_27785);
nor U29697 (N_29697,N_26264,N_27036);
and U29698 (N_29698,N_26335,N_26503);
nand U29699 (N_29699,N_26268,N_27432);
or U29700 (N_29700,N_26753,N_27843);
nand U29701 (N_29701,N_26624,N_27174);
nor U29702 (N_29702,N_26468,N_26922);
and U29703 (N_29703,N_27225,N_27814);
xnor U29704 (N_29704,N_26642,N_26775);
nor U29705 (N_29705,N_26295,N_27051);
and U29706 (N_29706,N_26197,N_27927);
xnor U29707 (N_29707,N_27310,N_26864);
nand U29708 (N_29708,N_27889,N_26131);
or U29709 (N_29709,N_26433,N_27112);
or U29710 (N_29710,N_27522,N_26862);
or U29711 (N_29711,N_26275,N_26920);
or U29712 (N_29712,N_26897,N_27328);
xnor U29713 (N_29713,N_26822,N_27898);
xnor U29714 (N_29714,N_27170,N_26201);
or U29715 (N_29715,N_26829,N_27710);
xor U29716 (N_29716,N_27398,N_27740);
nor U29717 (N_29717,N_26148,N_26892);
nand U29718 (N_29718,N_26964,N_27385);
xnor U29719 (N_29719,N_27519,N_26559);
nor U29720 (N_29720,N_27339,N_27852);
and U29721 (N_29721,N_26578,N_27376);
and U29722 (N_29722,N_27685,N_26788);
nand U29723 (N_29723,N_26981,N_27628);
and U29724 (N_29724,N_27044,N_27381);
and U29725 (N_29725,N_26580,N_26812);
and U29726 (N_29726,N_27856,N_26531);
xnor U29727 (N_29727,N_26245,N_27671);
or U29728 (N_29728,N_26642,N_27556);
and U29729 (N_29729,N_27896,N_26902);
or U29730 (N_29730,N_26499,N_27996);
xor U29731 (N_29731,N_27739,N_27211);
nor U29732 (N_29732,N_26581,N_27236);
and U29733 (N_29733,N_26737,N_27206);
and U29734 (N_29734,N_27193,N_27067);
nand U29735 (N_29735,N_26113,N_27829);
nand U29736 (N_29736,N_26208,N_26165);
or U29737 (N_29737,N_27139,N_27132);
xnor U29738 (N_29738,N_27486,N_27500);
xor U29739 (N_29739,N_26541,N_27503);
and U29740 (N_29740,N_27444,N_26429);
nand U29741 (N_29741,N_26098,N_27072);
nand U29742 (N_29742,N_27643,N_26184);
xnor U29743 (N_29743,N_27433,N_27787);
nor U29744 (N_29744,N_27737,N_27289);
nand U29745 (N_29745,N_26704,N_26774);
nor U29746 (N_29746,N_27140,N_26518);
nand U29747 (N_29747,N_26587,N_26183);
nor U29748 (N_29748,N_27387,N_27755);
or U29749 (N_29749,N_27093,N_27840);
or U29750 (N_29750,N_27852,N_27799);
and U29751 (N_29751,N_26195,N_26064);
and U29752 (N_29752,N_26973,N_27068);
and U29753 (N_29753,N_27097,N_27584);
nand U29754 (N_29754,N_27072,N_26342);
nand U29755 (N_29755,N_26128,N_26456);
nand U29756 (N_29756,N_27356,N_27275);
nor U29757 (N_29757,N_27489,N_27896);
or U29758 (N_29758,N_26630,N_26022);
or U29759 (N_29759,N_27286,N_27841);
or U29760 (N_29760,N_26613,N_27303);
and U29761 (N_29761,N_26754,N_27432);
and U29762 (N_29762,N_26171,N_27642);
or U29763 (N_29763,N_26914,N_27856);
nand U29764 (N_29764,N_26328,N_27749);
and U29765 (N_29765,N_27056,N_27881);
xor U29766 (N_29766,N_26258,N_26336);
nand U29767 (N_29767,N_26087,N_26466);
xor U29768 (N_29768,N_26767,N_27899);
nor U29769 (N_29769,N_26580,N_27560);
xnor U29770 (N_29770,N_27328,N_27243);
nor U29771 (N_29771,N_26412,N_27217);
xor U29772 (N_29772,N_27447,N_27631);
or U29773 (N_29773,N_26566,N_26977);
nor U29774 (N_29774,N_26920,N_26694);
and U29775 (N_29775,N_26555,N_26546);
or U29776 (N_29776,N_27942,N_26708);
nand U29777 (N_29777,N_27721,N_27154);
or U29778 (N_29778,N_27989,N_27858);
xnor U29779 (N_29779,N_26563,N_27649);
xor U29780 (N_29780,N_27367,N_26295);
xor U29781 (N_29781,N_26757,N_27020);
nor U29782 (N_29782,N_26048,N_27682);
nand U29783 (N_29783,N_26860,N_26457);
or U29784 (N_29784,N_26343,N_27320);
nor U29785 (N_29785,N_26577,N_26070);
or U29786 (N_29786,N_27979,N_27414);
and U29787 (N_29787,N_27883,N_26563);
and U29788 (N_29788,N_26408,N_27858);
or U29789 (N_29789,N_27721,N_26059);
nand U29790 (N_29790,N_27583,N_27761);
or U29791 (N_29791,N_26121,N_26814);
or U29792 (N_29792,N_26899,N_26614);
xnor U29793 (N_29793,N_27276,N_27617);
nor U29794 (N_29794,N_26079,N_26142);
nor U29795 (N_29795,N_27071,N_27424);
nor U29796 (N_29796,N_27000,N_27601);
xor U29797 (N_29797,N_26354,N_27301);
and U29798 (N_29798,N_27148,N_27756);
or U29799 (N_29799,N_27609,N_26309);
nand U29800 (N_29800,N_26836,N_26541);
nand U29801 (N_29801,N_27873,N_27359);
nand U29802 (N_29802,N_27258,N_26502);
and U29803 (N_29803,N_27560,N_26811);
nand U29804 (N_29804,N_26377,N_26800);
nand U29805 (N_29805,N_27752,N_27679);
and U29806 (N_29806,N_27523,N_26004);
and U29807 (N_29807,N_26071,N_27759);
and U29808 (N_29808,N_26717,N_26409);
nor U29809 (N_29809,N_26300,N_27981);
xor U29810 (N_29810,N_27706,N_26894);
or U29811 (N_29811,N_27534,N_26661);
and U29812 (N_29812,N_26014,N_27299);
nor U29813 (N_29813,N_27822,N_27732);
and U29814 (N_29814,N_26073,N_26603);
or U29815 (N_29815,N_27206,N_27296);
or U29816 (N_29816,N_27415,N_27319);
xnor U29817 (N_29817,N_26503,N_26914);
nand U29818 (N_29818,N_27916,N_26157);
or U29819 (N_29819,N_26363,N_26124);
nand U29820 (N_29820,N_26215,N_26783);
nor U29821 (N_29821,N_26475,N_27520);
nand U29822 (N_29822,N_26759,N_27304);
nor U29823 (N_29823,N_27566,N_27493);
xor U29824 (N_29824,N_26644,N_26194);
xor U29825 (N_29825,N_26113,N_26825);
and U29826 (N_29826,N_27089,N_26607);
xor U29827 (N_29827,N_26943,N_27076);
xnor U29828 (N_29828,N_26190,N_26163);
nand U29829 (N_29829,N_27167,N_26085);
nand U29830 (N_29830,N_26502,N_26243);
nand U29831 (N_29831,N_27329,N_26147);
and U29832 (N_29832,N_27315,N_27295);
nor U29833 (N_29833,N_27309,N_26943);
or U29834 (N_29834,N_26364,N_26000);
xor U29835 (N_29835,N_27810,N_26721);
and U29836 (N_29836,N_27629,N_27548);
nor U29837 (N_29837,N_27829,N_27288);
nand U29838 (N_29838,N_27911,N_27248);
nor U29839 (N_29839,N_26192,N_26279);
nand U29840 (N_29840,N_27683,N_27631);
and U29841 (N_29841,N_27015,N_26810);
or U29842 (N_29842,N_27998,N_26909);
nand U29843 (N_29843,N_27760,N_27838);
or U29844 (N_29844,N_27704,N_27561);
or U29845 (N_29845,N_27368,N_27155);
nor U29846 (N_29846,N_26468,N_26941);
nand U29847 (N_29847,N_26890,N_27675);
or U29848 (N_29848,N_27860,N_27720);
nand U29849 (N_29849,N_26786,N_26882);
nand U29850 (N_29850,N_26879,N_27776);
nor U29851 (N_29851,N_26005,N_27120);
or U29852 (N_29852,N_27608,N_27776);
xnor U29853 (N_29853,N_27481,N_27727);
and U29854 (N_29854,N_27699,N_26768);
nand U29855 (N_29855,N_26107,N_27829);
nand U29856 (N_29856,N_27866,N_26217);
nor U29857 (N_29857,N_27417,N_26827);
nor U29858 (N_29858,N_26508,N_27007);
and U29859 (N_29859,N_27737,N_27204);
xor U29860 (N_29860,N_27437,N_27732);
xnor U29861 (N_29861,N_27343,N_26797);
and U29862 (N_29862,N_27473,N_26794);
and U29863 (N_29863,N_26317,N_26085);
and U29864 (N_29864,N_26391,N_26826);
nand U29865 (N_29865,N_27394,N_27486);
and U29866 (N_29866,N_27894,N_27059);
nor U29867 (N_29867,N_26114,N_27624);
nor U29868 (N_29868,N_26325,N_26922);
xnor U29869 (N_29869,N_27610,N_26729);
nand U29870 (N_29870,N_26278,N_26842);
nor U29871 (N_29871,N_26999,N_27256);
nor U29872 (N_29872,N_26230,N_27327);
nand U29873 (N_29873,N_26418,N_27825);
and U29874 (N_29874,N_26092,N_27266);
or U29875 (N_29875,N_27582,N_27337);
nand U29876 (N_29876,N_26212,N_26441);
xnor U29877 (N_29877,N_26092,N_26223);
nor U29878 (N_29878,N_26660,N_27744);
xor U29879 (N_29879,N_27369,N_26185);
and U29880 (N_29880,N_26409,N_26609);
or U29881 (N_29881,N_26952,N_27525);
and U29882 (N_29882,N_26392,N_27089);
nor U29883 (N_29883,N_27152,N_27806);
or U29884 (N_29884,N_27470,N_27948);
and U29885 (N_29885,N_27076,N_27556);
or U29886 (N_29886,N_27399,N_26893);
nor U29887 (N_29887,N_27943,N_27630);
and U29888 (N_29888,N_27283,N_27915);
nand U29889 (N_29889,N_27556,N_27432);
or U29890 (N_29890,N_26737,N_27629);
and U29891 (N_29891,N_27528,N_26088);
nor U29892 (N_29892,N_26999,N_26963);
and U29893 (N_29893,N_27032,N_27348);
nor U29894 (N_29894,N_26512,N_27813);
nor U29895 (N_29895,N_26110,N_26315);
nor U29896 (N_29896,N_26223,N_27699);
nand U29897 (N_29897,N_26514,N_27707);
xor U29898 (N_29898,N_26967,N_26158);
nand U29899 (N_29899,N_27378,N_27961);
nor U29900 (N_29900,N_27276,N_26205);
xnor U29901 (N_29901,N_26364,N_27862);
nor U29902 (N_29902,N_26842,N_26267);
and U29903 (N_29903,N_26956,N_27729);
xnor U29904 (N_29904,N_27034,N_26383);
nor U29905 (N_29905,N_26433,N_27215);
or U29906 (N_29906,N_27484,N_26848);
or U29907 (N_29907,N_26384,N_26812);
or U29908 (N_29908,N_26018,N_26812);
nand U29909 (N_29909,N_27872,N_27509);
nor U29910 (N_29910,N_27717,N_26432);
and U29911 (N_29911,N_27666,N_27685);
or U29912 (N_29912,N_26438,N_26082);
nor U29913 (N_29913,N_26757,N_26141);
xnor U29914 (N_29914,N_26928,N_26367);
and U29915 (N_29915,N_27897,N_26897);
nor U29916 (N_29916,N_27712,N_26344);
nand U29917 (N_29917,N_26024,N_26494);
nor U29918 (N_29918,N_27866,N_26166);
or U29919 (N_29919,N_27687,N_27850);
xor U29920 (N_29920,N_26554,N_27401);
xor U29921 (N_29921,N_27138,N_26801);
nand U29922 (N_29922,N_27891,N_26373);
nand U29923 (N_29923,N_26430,N_26681);
xnor U29924 (N_29924,N_27322,N_27008);
or U29925 (N_29925,N_26101,N_26141);
xor U29926 (N_29926,N_26916,N_26500);
and U29927 (N_29927,N_26995,N_27298);
or U29928 (N_29928,N_27265,N_27586);
nor U29929 (N_29929,N_27474,N_27324);
nor U29930 (N_29930,N_27895,N_27624);
or U29931 (N_29931,N_26843,N_27200);
xor U29932 (N_29932,N_26185,N_27622);
nand U29933 (N_29933,N_27937,N_27365);
or U29934 (N_29934,N_27114,N_26915);
or U29935 (N_29935,N_26250,N_26572);
or U29936 (N_29936,N_26676,N_27319);
or U29937 (N_29937,N_27492,N_27341);
nand U29938 (N_29938,N_27747,N_27968);
xor U29939 (N_29939,N_27870,N_27350);
nor U29940 (N_29940,N_27768,N_27101);
or U29941 (N_29941,N_26211,N_27152);
or U29942 (N_29942,N_27540,N_26177);
or U29943 (N_29943,N_26624,N_26078);
xnor U29944 (N_29944,N_26155,N_26520);
xor U29945 (N_29945,N_26085,N_27558);
xor U29946 (N_29946,N_26751,N_27500);
or U29947 (N_29947,N_27914,N_27190);
nor U29948 (N_29948,N_26098,N_26668);
nor U29949 (N_29949,N_27759,N_26974);
nand U29950 (N_29950,N_27542,N_26465);
and U29951 (N_29951,N_26036,N_26099);
and U29952 (N_29952,N_27897,N_27797);
nor U29953 (N_29953,N_26806,N_27877);
xnor U29954 (N_29954,N_27481,N_27029);
xor U29955 (N_29955,N_27416,N_26818);
nand U29956 (N_29956,N_27872,N_26451);
nand U29957 (N_29957,N_27355,N_27858);
xnor U29958 (N_29958,N_27587,N_27282);
or U29959 (N_29959,N_26758,N_27549);
and U29960 (N_29960,N_26478,N_26696);
xor U29961 (N_29961,N_26334,N_27109);
and U29962 (N_29962,N_26403,N_26784);
xnor U29963 (N_29963,N_26450,N_27141);
or U29964 (N_29964,N_26976,N_27039);
nand U29965 (N_29965,N_27936,N_27682);
and U29966 (N_29966,N_26713,N_27102);
or U29967 (N_29967,N_27906,N_27538);
nand U29968 (N_29968,N_26501,N_26824);
xnor U29969 (N_29969,N_26390,N_26038);
nor U29970 (N_29970,N_26425,N_26639);
or U29971 (N_29971,N_26683,N_27639);
xor U29972 (N_29972,N_26198,N_27999);
or U29973 (N_29973,N_26933,N_27702);
nor U29974 (N_29974,N_26812,N_26770);
xor U29975 (N_29975,N_26032,N_26415);
and U29976 (N_29976,N_26622,N_26941);
nor U29977 (N_29977,N_27257,N_26090);
nor U29978 (N_29978,N_26088,N_27553);
xor U29979 (N_29979,N_26787,N_26962);
or U29980 (N_29980,N_26294,N_27315);
xor U29981 (N_29981,N_26654,N_27134);
xnor U29982 (N_29982,N_27990,N_26631);
xnor U29983 (N_29983,N_26705,N_26286);
nand U29984 (N_29984,N_26059,N_26517);
or U29985 (N_29985,N_27257,N_27757);
nand U29986 (N_29986,N_26346,N_27936);
or U29987 (N_29987,N_27551,N_26686);
nor U29988 (N_29988,N_26483,N_26642);
nand U29989 (N_29989,N_26186,N_27105);
nand U29990 (N_29990,N_27717,N_26273);
or U29991 (N_29991,N_27725,N_26347);
xnor U29992 (N_29992,N_26550,N_27438);
xor U29993 (N_29993,N_26344,N_27030);
and U29994 (N_29994,N_27560,N_26945);
or U29995 (N_29995,N_27161,N_26364);
and U29996 (N_29996,N_26688,N_26664);
nand U29997 (N_29997,N_26629,N_27725);
nand U29998 (N_29998,N_26456,N_27257);
nand U29999 (N_29999,N_26611,N_27115);
nand UO_0 (O_0,N_29606,N_28449);
or UO_1 (O_1,N_28564,N_28391);
or UO_2 (O_2,N_29431,N_29321);
nor UO_3 (O_3,N_28371,N_28526);
xnor UO_4 (O_4,N_29986,N_28657);
nor UO_5 (O_5,N_29622,N_28732);
or UO_6 (O_6,N_29067,N_28326);
xor UO_7 (O_7,N_28224,N_28436);
nand UO_8 (O_8,N_29104,N_28033);
xor UO_9 (O_9,N_29946,N_29728);
and UO_10 (O_10,N_28053,N_29615);
nor UO_11 (O_11,N_29926,N_28807);
and UO_12 (O_12,N_28468,N_28548);
and UO_13 (O_13,N_29921,N_28621);
xnor UO_14 (O_14,N_28571,N_29937);
or UO_15 (O_15,N_28139,N_29400);
nand UO_16 (O_16,N_28533,N_28856);
or UO_17 (O_17,N_29865,N_29248);
and UO_18 (O_18,N_28274,N_29740);
nand UO_19 (O_19,N_29528,N_28034);
nor UO_20 (O_20,N_29358,N_28589);
nor UO_21 (O_21,N_28045,N_29648);
nand UO_22 (O_22,N_28538,N_28675);
and UO_23 (O_23,N_29057,N_28926);
nand UO_24 (O_24,N_29930,N_29639);
or UO_25 (O_25,N_28568,N_29656);
nand UO_26 (O_26,N_28836,N_28430);
or UO_27 (O_27,N_29823,N_29134);
nor UO_28 (O_28,N_28499,N_29430);
nand UO_29 (O_29,N_28464,N_29729);
nand UO_30 (O_30,N_29895,N_29064);
or UO_31 (O_31,N_28269,N_29672);
and UO_32 (O_32,N_29611,N_28427);
nor UO_33 (O_33,N_28388,N_29311);
xnor UO_34 (O_34,N_29890,N_28220);
and UO_35 (O_35,N_28349,N_29291);
nand UO_36 (O_36,N_28007,N_28990);
and UO_37 (O_37,N_29440,N_29395);
and UO_38 (O_38,N_28744,N_29893);
or UO_39 (O_39,N_29530,N_28176);
and UO_40 (O_40,N_28591,N_29715);
or UO_41 (O_41,N_29276,N_29344);
and UO_42 (O_42,N_29000,N_28212);
nand UO_43 (O_43,N_28615,N_29689);
or UO_44 (O_44,N_28480,N_29174);
and UO_45 (O_45,N_28179,N_28511);
nand UO_46 (O_46,N_28469,N_28201);
nor UO_47 (O_47,N_28437,N_28477);
xor UO_48 (O_48,N_29241,N_28902);
or UO_49 (O_49,N_28022,N_28539);
nand UO_50 (O_50,N_29201,N_29073);
nand UO_51 (O_51,N_28780,N_28654);
or UO_52 (O_52,N_28300,N_29742);
nor UO_53 (O_53,N_29447,N_28324);
nor UO_54 (O_54,N_29901,N_28550);
and UO_55 (O_55,N_29145,N_28878);
nand UO_56 (O_56,N_29014,N_29853);
or UO_57 (O_57,N_28206,N_28377);
nor UO_58 (O_58,N_28114,N_29065);
or UO_59 (O_59,N_28310,N_29956);
nand UO_60 (O_60,N_28473,N_29820);
nand UO_61 (O_61,N_29676,N_28241);
or UO_62 (O_62,N_29283,N_28000);
xnor UO_63 (O_63,N_29750,N_29347);
nor UO_64 (O_64,N_28655,N_28186);
nand UO_65 (O_65,N_28113,N_29580);
or UO_66 (O_66,N_29852,N_29380);
and UO_67 (O_67,N_29122,N_29984);
and UO_68 (O_68,N_28989,N_28998);
or UO_69 (O_69,N_29476,N_29391);
and UO_70 (O_70,N_28059,N_29668);
and UO_71 (O_71,N_29263,N_28008);
and UO_72 (O_72,N_29691,N_28669);
or UO_73 (O_73,N_29747,N_29878);
xor UO_74 (O_74,N_28535,N_29875);
nor UO_75 (O_75,N_29135,N_29749);
xnor UO_76 (O_76,N_28638,N_28058);
xor UO_77 (O_77,N_28685,N_28789);
nor UO_78 (O_78,N_28135,N_29339);
nor UO_79 (O_79,N_28646,N_29288);
nand UO_80 (O_80,N_28697,N_29109);
or UO_81 (O_81,N_29814,N_29120);
nand UO_82 (O_82,N_28573,N_28094);
and UO_83 (O_83,N_29766,N_29950);
or UO_84 (O_84,N_29218,N_28360);
nand UO_85 (O_85,N_29496,N_28439);
nor UO_86 (O_86,N_29474,N_29598);
xnor UO_87 (O_87,N_29577,N_28065);
nand UO_88 (O_88,N_29088,N_28040);
and UO_89 (O_89,N_28971,N_28277);
nand UO_90 (O_90,N_29962,N_29807);
nand UO_91 (O_91,N_28566,N_28854);
or UO_92 (O_92,N_29690,N_29557);
and UO_93 (O_93,N_29624,N_28808);
and UO_94 (O_94,N_29170,N_29848);
nor UO_95 (O_95,N_28041,N_29399);
nand UO_96 (O_96,N_28181,N_29157);
and UO_97 (O_97,N_29374,N_29702);
or UO_98 (O_98,N_28106,N_29303);
nand UO_99 (O_99,N_29082,N_29049);
and UO_100 (O_100,N_28500,N_29739);
nor UO_101 (O_101,N_28378,N_28947);
nor UO_102 (O_102,N_28081,N_28766);
and UO_103 (O_103,N_28927,N_29277);
and UO_104 (O_104,N_29491,N_28747);
xnor UO_105 (O_105,N_28024,N_28017);
and UO_106 (O_106,N_29970,N_29599);
nand UO_107 (O_107,N_28945,N_29841);
nand UO_108 (O_108,N_28231,N_29163);
nor UO_109 (O_109,N_28835,N_28859);
nand UO_110 (O_110,N_29963,N_28910);
and UO_111 (O_111,N_28524,N_29034);
nand UO_112 (O_112,N_28426,N_29454);
nand UO_113 (O_113,N_28215,N_29781);
and UO_114 (O_114,N_29269,N_29971);
or UO_115 (O_115,N_29942,N_29197);
and UO_116 (O_116,N_28664,N_29481);
and UO_117 (O_117,N_28598,N_29623);
and UO_118 (O_118,N_29189,N_29097);
and UO_119 (O_119,N_28559,N_29118);
and UO_120 (O_120,N_28012,N_28896);
nor UO_121 (O_121,N_28769,N_29386);
or UO_122 (O_122,N_29762,N_28949);
nor UO_123 (O_123,N_28811,N_28422);
xor UO_124 (O_124,N_28346,N_28184);
nand UO_125 (O_125,N_29954,N_28607);
nand UO_126 (O_126,N_28092,N_29500);
and UO_127 (O_127,N_28954,N_28537);
nor UO_128 (O_128,N_29645,N_28493);
or UO_129 (O_129,N_28818,N_29007);
nor UO_130 (O_130,N_28628,N_28466);
nand UO_131 (O_131,N_28384,N_28881);
or UO_132 (O_132,N_29364,N_29011);
and UO_133 (O_133,N_28907,N_28913);
nor UO_134 (O_134,N_28751,N_28547);
nor UO_135 (O_135,N_29153,N_28996);
and UO_136 (O_136,N_29405,N_29768);
xor UO_137 (O_137,N_28093,N_29552);
nor UO_138 (O_138,N_29774,N_29313);
and UO_139 (O_139,N_28062,N_28032);
xor UO_140 (O_140,N_29327,N_28492);
nor UO_141 (O_141,N_29085,N_28305);
and UO_142 (O_142,N_29056,N_29151);
or UO_143 (O_143,N_28904,N_29732);
xnor UO_144 (O_144,N_29009,N_28508);
nor UO_145 (O_145,N_28060,N_29404);
or UO_146 (O_146,N_28358,N_28642);
nor UO_147 (O_147,N_29289,N_28767);
and UO_148 (O_148,N_28972,N_28948);
xor UO_149 (O_149,N_28395,N_29526);
or UO_150 (O_150,N_29351,N_28627);
or UO_151 (O_151,N_29023,N_28157);
and UO_152 (O_152,N_29935,N_28775);
and UO_153 (O_153,N_28631,N_28737);
xor UO_154 (O_154,N_29166,N_28400);
nor UO_155 (O_155,N_29519,N_28741);
and UO_156 (O_156,N_28174,N_29026);
nand UO_157 (O_157,N_28719,N_29199);
xnor UO_158 (O_158,N_29809,N_28680);
nand UO_159 (O_159,N_28584,N_28455);
xnor UO_160 (O_160,N_29748,N_28278);
or UO_161 (O_161,N_29037,N_28216);
nand UO_162 (O_162,N_28997,N_28484);
xnor UO_163 (O_163,N_29059,N_29468);
or UO_164 (O_164,N_28286,N_29936);
nor UO_165 (O_165,N_29429,N_28031);
and UO_166 (O_166,N_29804,N_28935);
and UO_167 (O_167,N_29206,N_28233);
and UO_168 (O_168,N_28411,N_28699);
or UO_169 (O_169,N_28474,N_28299);
nand UO_170 (O_170,N_29638,N_28551);
nor UO_171 (O_171,N_28844,N_29955);
and UO_172 (O_172,N_28612,N_28529);
and UO_173 (O_173,N_29121,N_28504);
nand UO_174 (O_174,N_29232,N_28321);
or UO_175 (O_175,N_29038,N_29805);
nor UO_176 (O_176,N_28188,N_28848);
or UO_177 (O_177,N_28763,N_29521);
xnor UO_178 (O_178,N_28160,N_28984);
or UO_179 (O_179,N_28110,N_29022);
nand UO_180 (O_180,N_28428,N_29205);
nand UO_181 (O_181,N_29460,N_28246);
nor UO_182 (O_182,N_29483,N_28438);
nand UO_183 (O_183,N_28703,N_29512);
and UO_184 (O_184,N_28334,N_28235);
nor UO_185 (O_185,N_28796,N_28170);
nor UO_186 (O_186,N_29791,N_28330);
and UO_187 (O_187,N_28689,N_29900);
xnor UO_188 (O_188,N_29495,N_28893);
nor UO_189 (O_189,N_29362,N_28145);
xnor UO_190 (O_190,N_29424,N_29258);
xor UO_191 (O_191,N_28639,N_28602);
nor UO_192 (O_192,N_29734,N_28676);
nor UO_193 (O_193,N_28868,N_29188);
nor UO_194 (O_194,N_29249,N_29060);
and UO_195 (O_195,N_28218,N_29782);
nand UO_196 (O_196,N_29063,N_28922);
and UO_197 (O_197,N_29903,N_29209);
or UO_198 (O_198,N_29741,N_28051);
xnor UO_199 (O_199,N_29572,N_29941);
or UO_200 (O_200,N_29973,N_29301);
xnor UO_201 (O_201,N_28790,N_28852);
and UO_202 (O_202,N_28653,N_29200);
nand UO_203 (O_203,N_29670,N_28830);
nor UO_204 (O_204,N_29533,N_28341);
and UO_205 (O_205,N_28142,N_28006);
nand UO_206 (O_206,N_29196,N_29977);
and UO_207 (O_207,N_28660,N_28776);
and UO_208 (O_208,N_28123,N_29198);
nor UO_209 (O_209,N_28528,N_29256);
nand UO_210 (O_210,N_29334,N_29952);
xor UO_211 (O_211,N_29260,N_29994);
nand UO_212 (O_212,N_28347,N_29757);
xor UO_213 (O_213,N_29219,N_29630);
and UO_214 (O_214,N_28647,N_29824);
or UO_215 (O_215,N_29033,N_29195);
and UO_216 (O_216,N_28519,N_28923);
nand UO_217 (O_217,N_28541,N_28617);
xor UO_218 (O_218,N_29383,N_28293);
nand UO_219 (O_219,N_29695,N_29688);
xor UO_220 (O_220,N_28555,N_28292);
or UO_221 (O_221,N_29136,N_28667);
nor UO_222 (O_222,N_29981,N_28987);
xor UO_223 (O_223,N_28873,N_29158);
and UO_224 (O_224,N_29634,N_29112);
nand UO_225 (O_225,N_28725,N_29305);
xor UO_226 (O_226,N_28226,N_29990);
xor UO_227 (O_227,N_29746,N_29337);
xor UO_228 (O_228,N_28588,N_29040);
or UO_229 (O_229,N_28272,N_28066);
nor UO_230 (O_230,N_28822,N_28963);
or UO_231 (O_231,N_28857,N_28781);
xor UO_232 (O_232,N_28316,N_29148);
and UO_233 (O_233,N_28478,N_29646);
xor UO_234 (O_234,N_28824,N_28076);
or UO_235 (O_235,N_28821,N_29051);
xnor UO_236 (O_236,N_28942,N_29819);
and UO_237 (O_237,N_29192,N_28462);
and UO_238 (O_238,N_29662,N_29967);
nand UO_239 (O_239,N_29714,N_29231);
xor UO_240 (O_240,N_28648,N_28219);
and UO_241 (O_241,N_29379,N_28633);
nand UO_242 (O_242,N_28013,N_29564);
nand UO_243 (O_243,N_29003,N_28788);
nor UO_244 (O_244,N_29470,N_28026);
xor UO_245 (O_245,N_28086,N_28952);
xor UO_246 (O_246,N_29094,N_28661);
xor UO_247 (O_247,N_29242,N_29816);
and UO_248 (O_248,N_28682,N_29434);
nand UO_249 (O_249,N_28596,N_29870);
xor UO_250 (O_250,N_28151,N_28687);
xor UO_251 (O_251,N_28536,N_29610);
or UO_252 (O_252,N_28728,N_28916);
or UO_253 (O_253,N_29589,N_29250);
and UO_254 (O_254,N_28128,N_29832);
nand UO_255 (O_255,N_28713,N_29338);
or UO_256 (O_256,N_28275,N_28629);
nand UO_257 (O_257,N_29043,N_29008);
xor UO_258 (O_258,N_29324,N_29444);
xor UO_259 (O_259,N_29290,N_28879);
nor UO_260 (O_260,N_28105,N_28851);
nor UO_261 (O_261,N_29851,N_29329);
or UO_262 (O_262,N_29923,N_29382);
nand UO_263 (O_263,N_29132,N_29180);
xor UO_264 (O_264,N_28837,N_29708);
nor UO_265 (O_265,N_29932,N_29677);
nor UO_266 (O_266,N_29068,N_29091);
or UO_267 (O_267,N_28425,N_28716);
nor UO_268 (O_268,N_29278,N_29938);
xnor UO_269 (O_269,N_29764,N_29592);
xnor UO_270 (O_270,N_28173,N_28815);
or UO_271 (O_271,N_29562,N_28940);
and UO_272 (O_272,N_29463,N_28791);
nor UO_273 (O_273,N_28785,N_29234);
nand UO_274 (O_274,N_28369,N_29751);
nor UO_275 (O_275,N_28562,N_28577);
nand UO_276 (O_276,N_28283,N_29681);
xnor UO_277 (O_277,N_28574,N_28820);
or UO_278 (O_278,N_29540,N_29997);
nor UO_279 (O_279,N_29369,N_28995);
or UO_280 (O_280,N_29588,N_28928);
xor UO_281 (O_281,N_29911,N_29125);
nand UO_282 (O_282,N_28930,N_28208);
xnor UO_283 (O_283,N_29467,N_29511);
nor UO_284 (O_284,N_29368,N_29951);
nand UO_285 (O_285,N_29828,N_28625);
nand UO_286 (O_286,N_29266,N_29363);
xnor UO_287 (O_287,N_29129,N_29693);
nor UO_288 (O_288,N_28762,N_28244);
nor UO_289 (O_289,N_29015,N_29980);
or UO_290 (O_290,N_29272,N_28932);
xor UO_291 (O_291,N_29687,N_28297);
or UO_292 (O_292,N_29924,N_29866);
nand UO_293 (O_293,N_28523,N_29462);
nor UO_294 (O_294,N_29004,N_28485);
xnor UO_295 (O_295,N_29079,N_28759);
or UO_296 (O_296,N_28714,N_29896);
nand UO_297 (O_297,N_28800,N_29569);
nor UO_298 (O_298,N_28064,N_29076);
or UO_299 (O_299,N_29907,N_29953);
or UO_300 (O_300,N_28944,N_29867);
nand UO_301 (O_301,N_28946,N_29240);
nor UO_302 (O_302,N_29397,N_28214);
and UO_303 (O_303,N_28693,N_29760);
and UO_304 (O_304,N_28447,N_28498);
or UO_305 (O_305,N_28858,N_29767);
nor UO_306 (O_306,N_29210,N_28250);
nand UO_307 (O_307,N_28002,N_29046);
nor UO_308 (O_308,N_28921,N_28140);
nor UO_309 (O_309,N_28554,N_29909);
nor UO_310 (O_310,N_28943,N_29756);
or UO_311 (O_311,N_28071,N_29185);
and UO_312 (O_312,N_29947,N_29143);
xor UO_313 (O_313,N_29419,N_29720);
nand UO_314 (O_314,N_29054,N_28668);
xor UO_315 (O_315,N_28705,N_28175);
nor UO_316 (O_316,N_28882,N_29675);
xor UO_317 (O_317,N_28262,N_28581);
and UO_318 (O_318,N_28520,N_29617);
xor UO_319 (O_319,N_29510,N_29207);
nor UO_320 (O_320,N_29261,N_28479);
nand UO_321 (O_321,N_29513,N_28711);
xnor UO_322 (O_322,N_28959,N_29355);
and UO_323 (O_323,N_28784,N_29407);
nor UO_324 (O_324,N_29944,N_28599);
nor UO_325 (O_325,N_29711,N_29888);
nor UO_326 (O_326,N_28870,N_28252);
nand UO_327 (O_327,N_29803,N_29723);
and UO_328 (O_328,N_28080,N_29317);
or UO_329 (O_329,N_28163,N_29408);
xnor UO_330 (O_330,N_28295,N_29836);
nor UO_331 (O_331,N_29830,N_29945);
and UO_332 (O_332,N_29593,N_29092);
or UO_333 (O_333,N_28325,N_29307);
and UO_334 (O_334,N_29531,N_29846);
nand UO_335 (O_335,N_29680,N_29426);
and UO_336 (O_336,N_28553,N_29964);
nand UO_337 (O_337,N_29699,N_28649);
nor UO_338 (O_338,N_28409,N_29632);
nand UO_339 (O_339,N_29785,N_29243);
xor UO_340 (O_340,N_29108,N_28414);
nand UO_341 (O_341,N_29354,N_28307);
xnor UO_342 (O_342,N_29486,N_29403);
nand UO_343 (O_343,N_28379,N_28386);
xnor UO_344 (O_344,N_29503,N_29547);
and UO_345 (O_345,N_29822,N_28417);
nor UO_346 (O_346,N_28842,N_28476);
nor UO_347 (O_347,N_28756,N_28465);
xor UO_348 (O_348,N_29908,N_29124);
and UO_349 (O_349,N_28637,N_28150);
and UO_350 (O_350,N_29518,N_28770);
and UO_351 (O_351,N_29647,N_28825);
nand UO_352 (O_352,N_29152,N_29144);
or UO_353 (O_353,N_29071,N_28435);
and UO_354 (O_354,N_29775,N_29988);
nor UO_355 (O_355,N_28098,N_29139);
nor UO_356 (O_356,N_29817,N_28534);
and UO_357 (O_357,N_29758,N_28578);
xnor UO_358 (O_358,N_29031,N_28232);
or UO_359 (O_359,N_29826,N_29922);
nand UO_360 (O_360,N_29799,N_28593);
nor UO_361 (O_361,N_29709,N_28147);
nor UO_362 (O_362,N_28407,N_29464);
nand UO_363 (O_363,N_29727,N_28875);
and UO_364 (O_364,N_29275,N_28701);
nand UO_365 (O_365,N_28387,N_29456);
xor UO_366 (O_366,N_28068,N_28456);
xor UO_367 (O_367,N_29626,N_28494);
and UO_368 (O_368,N_28351,N_29897);
or UO_369 (O_369,N_28679,N_29889);
nor UO_370 (O_370,N_29235,N_28956);
nor UO_371 (O_371,N_29215,N_28595);
or UO_372 (O_372,N_28681,N_28396);
xor UO_373 (O_373,N_28953,N_29707);
xor UO_374 (O_374,N_28333,N_28515);
and UO_375 (O_375,N_28453,N_29735);
xor UO_376 (O_376,N_28799,N_29187);
or UO_377 (O_377,N_29162,N_28302);
xor UO_378 (O_378,N_29508,N_28199);
nand UO_379 (O_379,N_29300,N_29792);
nand UO_380 (O_380,N_29423,N_29323);
xor UO_381 (O_381,N_29566,N_28168);
nand UO_382 (O_382,N_29297,N_28936);
or UO_383 (O_383,N_29621,N_28889);
nor UO_384 (O_384,N_29585,N_29045);
and UO_385 (O_385,N_29265,N_29542);
xor UO_386 (O_386,N_28727,N_28223);
and UO_387 (O_387,N_29103,N_28684);
nor UO_388 (O_388,N_29372,N_29330);
xor UO_389 (O_389,N_29216,N_28306);
and UO_390 (O_390,N_29571,N_28416);
and UO_391 (O_391,N_29879,N_29126);
or UO_392 (O_392,N_28171,N_29925);
or UO_393 (O_393,N_28490,N_29722);
nor UO_394 (O_394,N_29072,N_28507);
xor UO_395 (O_395,N_28193,N_29696);
or UO_396 (O_396,N_29427,N_28644);
nand UO_397 (O_397,N_28354,N_28084);
nand UO_398 (O_398,N_28020,N_28606);
and UO_399 (O_399,N_28245,N_29357);
xor UO_400 (O_400,N_29812,N_29295);
and UO_401 (O_401,N_28517,N_29062);
nor UO_402 (O_402,N_28258,N_28254);
xnor UO_403 (O_403,N_29815,N_29560);
nor UO_404 (O_404,N_29349,N_28078);
and UO_405 (O_405,N_29413,N_29302);
nand UO_406 (O_406,N_29414,N_28243);
xor UO_407 (O_407,N_28707,N_29539);
nand UO_408 (O_408,N_28724,N_28828);
or UO_409 (O_409,N_29578,N_28885);
nand UO_410 (O_410,N_29021,N_28502);
and UO_411 (O_411,N_28804,N_28817);
xnor UO_412 (O_412,N_29299,N_29002);
and UO_413 (O_413,N_28154,N_29957);
xor UO_414 (O_414,N_28200,N_28225);
nand UO_415 (O_415,N_28318,N_29416);
or UO_416 (O_416,N_29227,N_28023);
xor UO_417 (O_417,N_28605,N_28015);
or UO_418 (O_418,N_29983,N_29590);
nand UO_419 (O_419,N_28813,N_28671);
and UO_420 (O_420,N_28700,N_28202);
and UO_421 (O_421,N_28563,N_28366);
nand UO_422 (O_422,N_28715,N_28290);
nand UO_423 (O_423,N_29459,N_28385);
or UO_424 (O_424,N_28843,N_29591);
and UO_425 (O_425,N_28883,N_29716);
xor UO_426 (O_426,N_29532,N_29501);
nand UO_427 (O_427,N_28792,N_29381);
nand UO_428 (O_428,N_28383,N_28733);
nor UO_429 (O_429,N_28937,N_29522);
nand UO_430 (O_430,N_28393,N_29497);
and UO_431 (O_431,N_28723,N_28382);
or UO_432 (O_432,N_28609,N_28442);
nand UO_433 (O_433,N_28116,N_29343);
or UO_434 (O_434,N_29341,N_29432);
xnor UO_435 (O_435,N_29107,N_28567);
or UO_436 (O_436,N_29361,N_28911);
xnor UO_437 (O_437,N_28014,N_28459);
nand UO_438 (O_438,N_28344,N_28753);
nor UO_439 (O_439,N_28810,N_28903);
and UO_440 (O_440,N_29529,N_28164);
xnor UO_441 (O_441,N_28522,N_29485);
nand UO_442 (O_442,N_29320,N_29721);
nor UO_443 (O_443,N_29884,N_28191);
nor UO_444 (O_444,N_29346,N_28692);
or UO_445 (O_445,N_29933,N_28748);
and UO_446 (O_446,N_28056,N_29348);
or UO_447 (O_447,N_29902,N_28153);
xnor UO_448 (O_448,N_29296,N_28118);
and UO_449 (O_449,N_29974,N_29371);
and UO_450 (O_450,N_29600,N_28827);
and UO_451 (O_451,N_28390,N_29736);
xor UO_452 (O_452,N_29582,N_28339);
or UO_453 (O_453,N_28194,N_29252);
nand UO_454 (O_454,N_28136,N_29154);
nand UO_455 (O_455,N_29827,N_28213);
nand UO_456 (O_456,N_28992,N_28565);
xnor UO_457 (O_457,N_28048,N_28542);
nand UO_458 (O_458,N_28892,N_28042);
xnor UO_459 (O_459,N_29969,N_28203);
and UO_460 (O_460,N_29664,N_29777);
nand UO_461 (O_461,N_29657,N_29527);
nor UO_462 (O_462,N_29948,N_28454);
or UO_463 (O_463,N_29442,N_29202);
nand UO_464 (O_464,N_29058,N_28061);
nor UO_465 (O_465,N_29917,N_29563);
and UO_466 (O_466,N_29683,N_28802);
nor UO_467 (O_467,N_29373,N_29978);
and UO_468 (O_468,N_28909,N_28688);
nor UO_469 (O_469,N_29452,N_29850);
or UO_470 (O_470,N_28444,N_29077);
nor UO_471 (O_471,N_28982,N_28557);
and UO_472 (O_472,N_28124,N_28090);
xnor UO_473 (O_473,N_29975,N_29465);
xor UO_474 (O_474,N_29319,N_28240);
or UO_475 (O_475,N_29553,N_28141);
and UO_476 (O_476,N_28125,N_29927);
nand UO_477 (O_477,N_29667,N_28976);
nor UO_478 (O_478,N_29451,N_29370);
or UO_479 (O_479,N_29417,N_29854);
nor UO_480 (O_480,N_29783,N_29469);
nor UO_481 (O_481,N_28758,N_28079);
nand UO_482 (O_482,N_28722,N_28083);
nor UO_483 (O_483,N_29184,N_28227);
nor UO_484 (O_484,N_28905,N_29894);
nand UO_485 (O_485,N_28755,N_28658);
or UO_486 (O_486,N_28036,N_29435);
and UO_487 (O_487,N_29268,N_29800);
or UO_488 (O_488,N_28399,N_28545);
xnor UO_489 (O_489,N_28918,N_28690);
xor UO_490 (O_490,N_28210,N_28100);
nand UO_491 (O_491,N_29259,N_28611);
xnor UO_492 (O_492,N_28472,N_29883);
and UO_493 (O_493,N_28331,N_29710);
and UO_494 (O_494,N_29471,N_28891);
or UO_495 (O_495,N_28424,N_29237);
xnor UO_496 (O_496,N_29918,N_29509);
and UO_497 (O_497,N_29765,N_29738);
or UO_498 (O_498,N_28457,N_29934);
and UO_499 (O_499,N_28717,N_29725);
xnor UO_500 (O_500,N_29081,N_28343);
nor UO_501 (O_501,N_28887,N_29834);
and UO_502 (O_502,N_29649,N_28010);
and UO_503 (O_503,N_28709,N_29795);
nor UO_504 (O_504,N_28683,N_29813);
and UO_505 (O_505,N_28234,N_28204);
and UO_506 (O_506,N_28643,N_28993);
or UO_507 (O_507,N_29780,N_29095);
and UO_508 (O_508,N_28257,N_28276);
or UO_509 (O_509,N_29704,N_28569);
nor UO_510 (O_510,N_28248,N_28877);
nand UO_511 (O_511,N_28067,N_28259);
and UO_512 (O_512,N_29692,N_29254);
and UO_513 (O_513,N_28619,N_28251);
nand UO_514 (O_514,N_29776,N_28624);
nor UO_515 (O_515,N_29601,N_29353);
or UO_516 (O_516,N_28475,N_28432);
and UO_517 (O_517,N_28576,N_28798);
and UO_518 (O_518,N_29770,N_29743);
nand UO_519 (O_519,N_28876,N_28718);
or UO_520 (O_520,N_29833,N_29331);
xor UO_521 (O_521,N_28115,N_28806);
xnor UO_522 (O_522,N_29253,N_28489);
and UO_523 (O_523,N_28801,N_29101);
xor UO_524 (O_524,N_29796,N_29779);
nor UO_525 (O_525,N_28180,N_28994);
or UO_526 (O_526,N_28372,N_29069);
nand UO_527 (O_527,N_28890,N_29644);
nand UO_528 (O_528,N_28710,N_29494);
xor UO_529 (O_529,N_28988,N_29390);
nand UO_530 (O_530,N_28483,N_29113);
xor UO_531 (O_531,N_29332,N_29411);
nand UO_532 (O_532,N_28745,N_29912);
nand UO_533 (O_533,N_28419,N_29613);
and UO_534 (O_534,N_29763,N_29394);
nor UO_535 (O_535,N_28312,N_28603);
nor UO_536 (O_536,N_28686,N_29309);
nor UO_537 (O_537,N_28301,N_28739);
nand UO_538 (O_538,N_28217,N_29958);
or UO_539 (O_539,N_28746,N_29385);
or UO_540 (O_540,N_29441,N_28367);
or UO_541 (O_541,N_29790,N_28678);
or UO_542 (O_542,N_29160,N_29137);
and UO_543 (O_543,N_28267,N_28107);
and UO_544 (O_544,N_29906,N_29472);
and UO_545 (O_545,N_29998,N_29279);
nor UO_546 (O_546,N_28146,N_29274);
nand UO_547 (O_547,N_28497,N_28166);
and UO_548 (O_548,N_28884,N_29028);
and UO_549 (O_549,N_28281,N_28506);
or UO_550 (O_550,N_29401,N_29966);
nand UO_551 (O_551,N_28665,N_28055);
xor UO_552 (O_552,N_29769,N_28803);
xor UO_553 (O_553,N_29115,N_28518);
nor UO_554 (O_554,N_28359,N_29844);
or UO_555 (O_555,N_28284,N_29433);
nand UO_556 (O_556,N_28038,N_29480);
nor UO_557 (O_557,N_28011,N_28734);
xor UO_558 (O_558,N_29753,N_28412);
or UO_559 (O_559,N_29730,N_28434);
nand UO_560 (O_560,N_29376,N_28162);
or UO_561 (O_561,N_29182,N_28304);
xor UO_562 (O_562,N_29633,N_28237);
and UO_563 (O_563,N_28178,N_29869);
and UO_564 (O_564,N_28074,N_28287);
nor UO_565 (O_565,N_29831,N_28880);
nand UO_566 (O_566,N_28979,N_29236);
xor UO_567 (O_567,N_28361,N_28912);
nand UO_568 (O_568,N_28404,N_28247);
or UO_569 (O_569,N_29384,N_29410);
nor UO_570 (O_570,N_29114,N_29224);
nand UO_571 (O_571,N_29789,N_29524);
and UO_572 (O_572,N_28632,N_29794);
nand UO_573 (O_573,N_29556,N_29377);
nor UO_574 (O_574,N_29620,N_28487);
xnor UO_575 (O_575,N_29847,N_29179);
and UO_576 (O_576,N_29388,N_28941);
and UO_577 (O_577,N_29147,N_28630);
or UO_578 (O_578,N_29345,N_28298);
or UO_579 (O_579,N_28091,N_29705);
and UO_580 (O_580,N_29579,N_29514);
nand UO_581 (O_581,N_29005,N_29335);
nor UO_582 (O_582,N_28674,N_29245);
or UO_583 (O_583,N_28320,N_29106);
nor UO_584 (O_584,N_29546,N_28618);
or UO_585 (O_585,N_28509,N_29418);
nor UO_586 (O_586,N_28543,N_29016);
or UO_587 (O_587,N_29943,N_29857);
or UO_588 (O_588,N_28864,N_29636);
and UO_589 (O_589,N_28104,N_29992);
xnor UO_590 (O_590,N_28336,N_29138);
xor UO_591 (O_591,N_28192,N_29133);
nor UO_592 (O_592,N_29492,N_28221);
or UO_593 (O_593,N_29913,N_29164);
nor UO_594 (O_594,N_28964,N_29558);
nand UO_595 (O_595,N_29650,N_28838);
nand UO_596 (O_596,N_28018,N_29223);
nand UO_597 (O_597,N_29719,N_28491);
xor UO_598 (O_598,N_28917,N_29169);
or UO_599 (O_599,N_28402,N_28981);
nand UO_600 (O_600,N_29194,N_29183);
nand UO_601 (O_601,N_28021,N_29534);
nand UO_602 (O_602,N_29538,N_29786);
or UO_603 (O_603,N_29336,N_28120);
nand UO_604 (O_604,N_28743,N_28754);
or UO_605 (O_605,N_28616,N_29246);
nand UO_606 (O_606,N_29450,N_28672);
nor UO_607 (O_607,N_28960,N_28398);
or UO_608 (O_608,N_28532,N_28317);
nand UO_609 (O_609,N_28119,N_28708);
and UO_610 (O_610,N_28005,N_29191);
and UO_611 (O_611,N_29161,N_28924);
nor UO_612 (O_612,N_29352,N_28253);
nor UO_613 (O_613,N_29387,N_29842);
nor UO_614 (O_614,N_29919,N_29996);
and UO_615 (O_615,N_28773,N_28027);
or UO_616 (O_616,N_29284,N_28239);
nand UO_617 (O_617,N_29421,N_28908);
xnor UO_618 (O_618,N_29304,N_28037);
xnor UO_619 (O_619,N_28777,N_29286);
and UO_620 (O_620,N_29586,N_29396);
nor UO_621 (O_621,N_28112,N_29181);
xnor UO_622 (O_622,N_28441,N_29325);
nand UO_623 (O_623,N_29378,N_28148);
and UO_624 (O_624,N_29642,N_28311);
or UO_625 (O_625,N_28131,N_29220);
nand UO_626 (O_626,N_29149,N_28418);
nor UO_627 (O_627,N_28263,N_29316);
and UO_628 (O_628,N_29455,N_28967);
nand UO_629 (O_629,N_28991,N_28211);
nor UO_630 (O_630,N_28364,N_28742);
xor UO_631 (O_631,N_29641,N_28951);
or UO_632 (O_632,N_29959,N_29665);
nand UO_633 (O_633,N_29328,N_28558);
or UO_634 (O_634,N_29653,N_28831);
nand UO_635 (O_635,N_28793,N_28450);
nor UO_636 (O_636,N_29609,N_29604);
nor UO_637 (O_637,N_29096,N_29517);
or UO_638 (O_638,N_28894,N_29554);
nand UO_639 (O_639,N_29825,N_28900);
nor UO_640 (O_640,N_29211,N_29123);
nor UO_641 (O_641,N_29712,N_28888);
xor UO_642 (O_642,N_29165,N_28587);
or UO_643 (O_643,N_28289,N_29087);
xnor UO_644 (O_644,N_28774,N_29287);
or UO_645 (O_645,N_29493,N_28075);
nor UO_646 (O_646,N_28832,N_29655);
nor UO_647 (O_647,N_28329,N_28406);
xnor UO_648 (O_648,N_29318,N_28514);
and UO_649 (O_649,N_28860,N_28268);
or UO_650 (O_650,N_28190,N_29239);
and UO_651 (O_651,N_29457,N_29629);
nand UO_652 (O_652,N_28920,N_28730);
and UO_653 (O_653,N_28337,N_28172);
and UO_654 (O_654,N_28256,N_29840);
nand UO_655 (O_655,N_28582,N_29731);
and UO_656 (O_656,N_28155,N_28122);
nor UO_657 (O_657,N_28285,N_28975);
nand UO_658 (O_658,N_28829,N_28265);
nor UO_659 (O_659,N_29084,N_29899);
and UO_660 (O_660,N_28270,N_29159);
nor UO_661 (O_661,N_28552,N_29616);
or UO_662 (O_662,N_29628,N_29772);
nor UO_663 (O_663,N_29713,N_28482);
nor UO_664 (O_664,N_28610,N_29920);
nand UO_665 (O_665,N_29845,N_29939);
or UO_666 (O_666,N_29267,N_29027);
or UO_667 (O_667,N_28696,N_29543);
and UO_668 (O_668,N_28871,N_29855);
and UO_669 (O_669,N_28600,N_28117);
nor UO_670 (O_670,N_28452,N_29535);
and UO_671 (O_671,N_29523,N_29987);
nand UO_672 (O_672,N_28082,N_28063);
nand UO_673 (O_673,N_28282,N_29873);
xor UO_674 (O_674,N_28029,N_28613);
xnor UO_675 (O_675,N_28255,N_28512);
and UO_676 (O_676,N_28260,N_28488);
and UO_677 (O_677,N_28764,N_29843);
and UO_678 (O_678,N_28392,N_29861);
xnor UO_679 (O_679,N_28389,N_29359);
or UO_680 (O_680,N_29801,N_28348);
or UO_681 (O_681,N_29342,N_28356);
nor UO_682 (O_682,N_28645,N_29083);
nor UO_683 (O_683,N_28513,N_28271);
and UO_684 (O_684,N_28583,N_28721);
and UO_685 (O_685,N_29117,N_28463);
nand UO_686 (O_686,N_29298,N_28039);
and UO_687 (O_687,N_28322,N_28397);
or UO_688 (O_688,N_28101,N_29315);
nor UO_689 (O_689,N_28375,N_29488);
nand UO_690 (O_690,N_28525,N_29490);
nand UO_691 (O_691,N_28955,N_29217);
xnor UO_692 (O_692,N_29838,N_29443);
and UO_693 (O_693,N_28765,N_29544);
or UO_694 (O_694,N_29281,N_29565);
nand UO_695 (O_695,N_29515,N_28853);
nor UO_696 (O_696,N_29102,N_29050);
xnor UO_697 (O_697,N_28899,N_28156);
or UO_698 (O_698,N_28077,N_29561);
and UO_699 (O_699,N_28401,N_29602);
and UO_700 (O_700,N_29788,N_28816);
xnor UO_701 (O_701,N_28132,N_29186);
nand UO_702 (O_702,N_29333,N_29306);
nor UO_703 (O_703,N_29439,N_28279);
nand UO_704 (O_704,N_28839,N_29915);
and UO_705 (O_705,N_29643,N_29111);
nor UO_706 (O_706,N_28294,N_29458);
nor UO_707 (O_707,N_29409,N_28706);
nand UO_708 (O_708,N_28999,N_28760);
or UO_709 (O_709,N_29190,N_28812);
nand UO_710 (O_710,N_29487,N_29100);
nand UO_711 (O_711,N_28035,N_29036);
or UO_712 (O_712,N_29504,N_29863);
xor UO_713 (O_713,N_28109,N_29887);
and UO_714 (O_714,N_29233,N_29916);
xnor UO_715 (O_715,N_29759,N_29965);
or UO_716 (O_716,N_28846,N_29718);
and UO_717 (O_717,N_29314,N_29548);
nor UO_718 (O_718,N_28046,N_29929);
and UO_719 (O_719,N_29466,N_28652);
nand UO_720 (O_720,N_28694,N_28726);
nand UO_721 (O_721,N_28394,N_29603);
nand UO_722 (O_722,N_29025,N_28350);
or UO_723 (O_723,N_28866,N_28230);
nor UO_724 (O_724,N_28471,N_28865);
nand UO_725 (O_725,N_28752,N_28429);
nand UO_726 (O_726,N_29700,N_29128);
or UO_727 (O_727,N_28403,N_28266);
nor UO_728 (O_728,N_29568,N_29204);
or UO_729 (O_729,N_29262,N_29860);
nor UO_730 (O_730,N_29904,N_28458);
nand UO_731 (O_731,N_29238,N_28814);
xnor UO_732 (O_732,N_28794,N_28635);
xor UO_733 (O_733,N_28778,N_28604);
or UO_734 (O_734,N_29874,N_28530);
nor UO_735 (O_735,N_28749,N_28729);
nor UO_736 (O_736,N_28365,N_28362);
xor UO_737 (O_737,N_29818,N_28313);
or UO_738 (O_738,N_28057,N_29047);
xor UO_739 (O_739,N_28712,N_29859);
nand UO_740 (O_740,N_29674,N_28261);
nor UO_741 (O_741,N_29446,N_28704);
nand UO_742 (O_742,N_28047,N_28368);
xor UO_743 (O_743,N_29886,N_28826);
or UO_744 (O_744,N_29761,N_28691);
and UO_745 (O_745,N_28443,N_28833);
or UO_746 (O_746,N_29856,N_29545);
or UO_747 (O_747,N_29264,N_29651);
nor UO_748 (O_748,N_29663,N_29039);
or UO_749 (O_749,N_29478,N_28030);
nand UO_750 (O_750,N_28303,N_28666);
nor UO_751 (O_751,N_28608,N_28169);
nand UO_752 (O_752,N_28841,N_29745);
xnor UO_753 (O_753,N_28809,N_29872);
xnor UO_754 (O_754,N_29017,N_29596);
xnor UO_755 (O_755,N_28914,N_29473);
and UO_756 (O_756,N_29326,N_28054);
nor UO_757 (O_757,N_29099,N_29898);
nand UO_758 (O_758,N_29972,N_28962);
and UO_759 (O_759,N_29366,N_29208);
and UO_760 (O_760,N_28958,N_29482);
or UO_761 (O_761,N_28138,N_29484);
or UO_762 (O_762,N_28740,N_28620);
nand UO_763 (O_763,N_29502,N_29150);
xnor UO_764 (O_764,N_28572,N_28757);
nand UO_765 (O_765,N_29652,N_29398);
nor UO_766 (O_766,N_29030,N_29116);
nand UO_767 (O_767,N_28121,N_29551);
nand UO_768 (O_768,N_28886,N_28222);
xor UO_769 (O_769,N_29282,N_29612);
and UO_770 (O_770,N_29222,N_28805);
nor UO_771 (O_771,N_28420,N_28531);
nor UO_772 (O_772,N_29006,N_29787);
and UO_773 (O_773,N_29802,N_29032);
or UO_774 (O_774,N_28849,N_28556);
and UO_775 (O_775,N_28440,N_29090);
nand UO_776 (O_776,N_29976,N_28415);
xor UO_777 (O_777,N_29717,N_29280);
or UO_778 (O_778,N_29402,N_29445);
nand UO_779 (O_779,N_29993,N_28486);
or UO_780 (O_780,N_28236,N_28872);
nor UO_781 (O_781,N_28229,N_28750);
and UO_782 (O_782,N_29605,N_29669);
nor UO_783 (O_783,N_28673,N_29308);
or UO_784 (O_784,N_29477,N_29985);
and UO_785 (O_785,N_28503,N_28405);
nand UO_786 (O_786,N_29864,N_29881);
nor UO_787 (O_787,N_29167,N_28408);
nand UO_788 (O_788,N_28787,N_29858);
nor UO_789 (O_789,N_29995,N_28088);
nand UO_790 (O_790,N_28161,N_28087);
nor UO_791 (O_791,N_29285,N_29271);
xnor UO_792 (O_792,N_28095,N_28586);
nor UO_793 (O_793,N_29024,N_29449);
and UO_794 (O_794,N_29961,N_29559);
or UO_795 (O_795,N_29891,N_28874);
or UO_796 (O_796,N_28834,N_29367);
and UO_797 (O_797,N_29453,N_28677);
nor UO_798 (O_798,N_28126,N_28919);
nand UO_799 (O_799,N_28738,N_28597);
and UO_800 (O_800,N_29146,N_28044);
xnor UO_801 (O_801,N_29979,N_29479);
and UO_802 (O_802,N_29041,N_28205);
nor UO_803 (O_803,N_28373,N_28238);
and UO_804 (O_804,N_29678,N_28288);
or UO_805 (O_805,N_29698,N_29176);
and UO_806 (O_806,N_29255,N_28096);
and UO_807 (O_807,N_28980,N_29356);
and UO_808 (O_808,N_28898,N_29244);
and UO_809 (O_809,N_28965,N_28189);
and UO_810 (O_810,N_28698,N_28332);
and UO_811 (O_811,N_29679,N_28782);
and UO_812 (O_812,N_29541,N_29310);
and UO_813 (O_813,N_29110,N_29755);
or UO_814 (O_814,N_29877,N_29461);
xnor UO_815 (O_815,N_29744,N_28198);
or UO_816 (O_816,N_29882,N_28451);
nor UO_817 (O_817,N_29230,N_29597);
and UO_818 (O_818,N_29155,N_28363);
nand UO_819 (O_819,N_28481,N_28969);
xnor UO_820 (O_820,N_29661,N_29685);
and UO_821 (O_821,N_29797,N_28925);
xor UO_822 (O_822,N_29614,N_28934);
xor UO_823 (O_823,N_29928,N_29130);
nand UO_824 (O_824,N_28973,N_28280);
nand UO_825 (O_825,N_29013,N_29949);
or UO_826 (O_826,N_28069,N_28357);
xor UO_827 (O_827,N_28467,N_29098);
and UO_828 (O_828,N_29422,N_28663);
nand UO_829 (O_829,N_28867,N_28273);
or UO_830 (O_830,N_29570,N_29660);
nor UO_831 (O_831,N_28043,N_28376);
xnor UO_832 (O_832,N_28614,N_29835);
xnor UO_833 (O_833,N_28433,N_29020);
nor UO_834 (O_834,N_28662,N_29055);
nand UO_835 (O_835,N_29573,N_29849);
xnor UO_836 (O_836,N_28049,N_28544);
nor UO_837 (O_837,N_28165,N_28579);
nor UO_838 (O_838,N_29905,N_29119);
or UO_839 (O_839,N_29567,N_29131);
nor UO_840 (O_840,N_28143,N_28847);
and UO_841 (O_841,N_29203,N_28130);
nor UO_842 (O_842,N_29213,N_28901);
or UO_843 (O_843,N_29576,N_28413);
xor UO_844 (O_844,N_29048,N_28209);
or UO_845 (O_845,N_29627,N_29671);
and UO_846 (O_846,N_29555,N_29340);
or UO_847 (O_847,N_29537,N_29412);
xor UO_848 (O_848,N_28003,N_28445);
nand UO_849 (O_849,N_28659,N_28025);
nand UO_850 (O_850,N_28470,N_29142);
nor UO_851 (O_851,N_28575,N_29105);
nand UO_852 (O_852,N_28510,N_29686);
and UO_853 (O_853,N_29516,N_29778);
or UO_854 (O_854,N_29829,N_29910);
or UO_855 (O_855,N_28089,N_28772);
and UO_856 (O_856,N_28196,N_29640);
nor UO_857 (O_857,N_28862,N_29733);
or UO_858 (O_858,N_29584,N_29658);
xor UO_859 (O_859,N_29393,N_28977);
xnor UO_860 (O_860,N_28768,N_28797);
and UO_861 (O_861,N_29706,N_28845);
xor UO_862 (O_862,N_29075,N_29520);
nor UO_863 (O_863,N_29607,N_29193);
nand UO_864 (O_864,N_28516,N_29177);
and UO_865 (O_865,N_28521,N_28129);
nand UO_866 (O_866,N_28966,N_28421);
and UO_867 (O_867,N_29078,N_28149);
nand UO_868 (O_868,N_29837,N_28950);
nor UO_869 (O_869,N_29694,N_29312);
nor UO_870 (O_870,N_29550,N_29798);
or UO_871 (O_871,N_29581,N_29808);
nand UO_872 (O_872,N_28108,N_29489);
nand UO_873 (O_873,N_29940,N_29549);
nor UO_874 (O_874,N_29625,N_28072);
nand UO_875 (O_875,N_29810,N_28228);
xnor UO_876 (O_876,N_28915,N_29171);
nand UO_877 (O_877,N_29583,N_29701);
and UO_878 (O_878,N_29737,N_28895);
nor UO_879 (O_879,N_29536,N_29042);
or UO_880 (O_880,N_28137,N_28050);
xor UO_881 (O_881,N_28570,N_29322);
or UO_882 (O_882,N_29406,N_28001);
xnor UO_883 (O_883,N_28127,N_29871);
or UO_884 (O_884,N_29029,N_29425);
xnor UO_885 (O_885,N_29294,N_28735);
or UO_886 (O_886,N_28823,N_29415);
or UO_887 (O_887,N_29914,N_29931);
nor UO_888 (O_888,N_29752,N_29389);
or UO_889 (O_889,N_28446,N_28315);
xor UO_890 (O_890,N_29012,N_28352);
nor UO_891 (O_891,N_28009,N_28720);
and UO_892 (O_892,N_28505,N_29438);
or UO_893 (O_893,N_28779,N_29574);
and UO_894 (O_894,N_28460,N_29175);
xor UO_895 (O_895,N_28242,N_29436);
nor UO_896 (O_896,N_28296,N_28197);
xor UO_897 (O_897,N_29703,N_28327);
nand UO_898 (O_898,N_28978,N_29619);
nand UO_899 (O_899,N_28929,N_28783);
or UO_900 (O_900,N_29892,N_29499);
xnor UO_901 (O_901,N_29659,N_29635);
nand UO_902 (O_902,N_29999,N_29053);
nor UO_903 (O_903,N_29784,N_28736);
nor UO_904 (O_904,N_28308,N_28731);
or UO_905 (O_905,N_29806,N_29618);
xor UO_906 (O_906,N_29637,N_28182);
xnor UO_907 (O_907,N_28423,N_28319);
and UO_908 (O_908,N_28933,N_28342);
nor UO_909 (O_909,N_29035,N_28795);
or UO_910 (O_910,N_29862,N_29066);
nor UO_911 (O_911,N_29350,N_29684);
nand UO_912 (O_912,N_28640,N_29420);
and UO_913 (O_913,N_28938,N_29880);
and UO_914 (O_914,N_28897,N_28592);
or UO_915 (O_915,N_29089,N_28855);
nand UO_916 (O_916,N_28183,N_29960);
or UO_917 (O_917,N_28328,N_29811);
xnor UO_918 (O_918,N_29168,N_29010);
or UO_919 (O_919,N_29885,N_28028);
or UO_920 (O_920,N_29968,N_29044);
xnor UO_921 (O_921,N_29052,N_28623);
nor UO_922 (O_922,N_29595,N_28195);
or UO_923 (O_923,N_29251,N_29631);
or UO_924 (O_924,N_28207,N_29989);
or UO_925 (O_925,N_28019,N_29229);
and UO_926 (O_926,N_28670,N_28340);
xor UO_927 (O_927,N_29141,N_28355);
or UO_928 (O_928,N_28546,N_29991);
and UO_929 (O_929,N_28099,N_28187);
xnor UO_930 (O_930,N_29086,N_28819);
and UO_931 (O_931,N_29839,N_29127);
or UO_932 (O_932,N_28159,N_28496);
xnor UO_933 (O_933,N_28869,N_28102);
and UO_934 (O_934,N_29475,N_29773);
nand UO_935 (O_935,N_28986,N_28370);
nor UO_936 (O_936,N_29172,N_29001);
and UO_937 (O_937,N_28560,N_29225);
nor UO_938 (O_938,N_28850,N_28410);
and UO_939 (O_939,N_28626,N_29375);
and UO_940 (O_940,N_29654,N_28974);
nand UO_941 (O_941,N_29070,N_28786);
or UO_942 (O_942,N_29061,N_28185);
or UO_943 (O_943,N_28291,N_28004);
or UO_944 (O_944,N_28103,N_29156);
xor UO_945 (O_945,N_28431,N_28097);
and UO_946 (O_946,N_29587,N_29392);
and UO_947 (O_947,N_29793,N_28939);
and UO_948 (O_948,N_28249,N_29594);
nand UO_949 (O_949,N_29505,N_28702);
and UO_950 (O_950,N_28656,N_29754);
xnor UO_951 (O_951,N_29821,N_28374);
xnor UO_952 (O_952,N_28931,N_28501);
nor UO_953 (O_953,N_28771,N_29173);
nand UO_954 (O_954,N_28863,N_28840);
and UO_955 (O_955,N_28968,N_28549);
nor UO_956 (O_956,N_29724,N_28323);
or UO_957 (O_957,N_28016,N_28636);
or UO_958 (O_958,N_29293,N_28695);
xnor UO_959 (O_959,N_28983,N_29221);
nor UO_960 (O_960,N_28970,N_29018);
nand UO_961 (O_961,N_28861,N_28085);
and UO_962 (O_962,N_29140,N_29257);
nand UO_963 (O_963,N_28957,N_28314);
and UO_964 (O_964,N_28650,N_29666);
and UO_965 (O_965,N_28158,N_29428);
xnor UO_966 (O_966,N_28345,N_28264);
and UO_967 (O_967,N_29525,N_29982);
and UO_968 (O_968,N_28641,N_29868);
and UO_969 (O_969,N_29212,N_28073);
nor UO_970 (O_970,N_29019,N_28580);
or UO_971 (O_971,N_28052,N_28134);
nand UO_972 (O_972,N_28622,N_29448);
nand UO_973 (O_973,N_28380,N_29093);
or UO_974 (O_974,N_28585,N_29697);
or UO_975 (O_975,N_29876,N_28111);
or UO_976 (O_976,N_29506,N_29365);
xor UO_977 (O_977,N_28461,N_29437);
or UO_978 (O_978,N_29771,N_28634);
xnor UO_979 (O_979,N_29673,N_28961);
and UO_980 (O_980,N_29726,N_28590);
and UO_981 (O_981,N_29498,N_28761);
nand UO_982 (O_982,N_28167,N_28381);
nand UO_983 (O_983,N_28985,N_29360);
nor UO_984 (O_984,N_28651,N_28152);
or UO_985 (O_985,N_28540,N_29178);
and UO_986 (O_986,N_29270,N_28144);
or UO_987 (O_987,N_29074,N_28338);
nor UO_988 (O_988,N_28448,N_29682);
xnor UO_989 (O_989,N_28133,N_28527);
nand UO_990 (O_990,N_28906,N_28561);
nor UO_991 (O_991,N_28601,N_28594);
xor UO_992 (O_992,N_29608,N_29507);
xnor UO_993 (O_993,N_28353,N_29214);
or UO_994 (O_994,N_29226,N_29273);
nor UO_995 (O_995,N_28309,N_29080);
or UO_996 (O_996,N_28495,N_28070);
xor UO_997 (O_997,N_29247,N_28177);
and UO_998 (O_998,N_28335,N_29228);
nor UO_999 (O_999,N_29575,N_29292);
nor UO_1000 (O_1000,N_28039,N_28644);
or UO_1001 (O_1001,N_29131,N_28939);
nor UO_1002 (O_1002,N_29002,N_29241);
nor UO_1003 (O_1003,N_28894,N_29465);
or UO_1004 (O_1004,N_28256,N_29306);
or UO_1005 (O_1005,N_29820,N_28567);
nor UO_1006 (O_1006,N_28627,N_28987);
xor UO_1007 (O_1007,N_28838,N_29554);
and UO_1008 (O_1008,N_29477,N_29195);
nor UO_1009 (O_1009,N_29350,N_28566);
nor UO_1010 (O_1010,N_29409,N_29334);
xor UO_1011 (O_1011,N_29982,N_28207);
and UO_1012 (O_1012,N_28928,N_28770);
or UO_1013 (O_1013,N_29116,N_29654);
and UO_1014 (O_1014,N_29045,N_28652);
or UO_1015 (O_1015,N_28871,N_28985);
nand UO_1016 (O_1016,N_28225,N_29857);
nand UO_1017 (O_1017,N_28018,N_29263);
nor UO_1018 (O_1018,N_29226,N_29959);
nor UO_1019 (O_1019,N_29939,N_29359);
xor UO_1020 (O_1020,N_29813,N_28632);
nand UO_1021 (O_1021,N_28750,N_29925);
xor UO_1022 (O_1022,N_28726,N_28084);
or UO_1023 (O_1023,N_29773,N_28880);
nor UO_1024 (O_1024,N_28961,N_28591);
xor UO_1025 (O_1025,N_29963,N_28727);
nand UO_1026 (O_1026,N_29929,N_28550);
or UO_1027 (O_1027,N_28833,N_28516);
or UO_1028 (O_1028,N_28641,N_29734);
xnor UO_1029 (O_1029,N_29854,N_29747);
xor UO_1030 (O_1030,N_29229,N_29398);
and UO_1031 (O_1031,N_29088,N_29806);
nor UO_1032 (O_1032,N_29699,N_28045);
nand UO_1033 (O_1033,N_29484,N_28317);
nor UO_1034 (O_1034,N_28686,N_28289);
nand UO_1035 (O_1035,N_28927,N_28988);
nand UO_1036 (O_1036,N_29135,N_28307);
or UO_1037 (O_1037,N_29796,N_28830);
nor UO_1038 (O_1038,N_29384,N_28122);
nand UO_1039 (O_1039,N_29509,N_28337);
xor UO_1040 (O_1040,N_28642,N_29660);
nor UO_1041 (O_1041,N_29533,N_29181);
nor UO_1042 (O_1042,N_28692,N_29794);
and UO_1043 (O_1043,N_28999,N_28227);
nand UO_1044 (O_1044,N_29045,N_29654);
and UO_1045 (O_1045,N_29788,N_29845);
nor UO_1046 (O_1046,N_28931,N_29069);
nor UO_1047 (O_1047,N_28231,N_29659);
nor UO_1048 (O_1048,N_28331,N_29450);
or UO_1049 (O_1049,N_28612,N_28754);
and UO_1050 (O_1050,N_28710,N_29018);
nor UO_1051 (O_1051,N_28589,N_29634);
and UO_1052 (O_1052,N_29788,N_29002);
xor UO_1053 (O_1053,N_29306,N_29262);
and UO_1054 (O_1054,N_29598,N_29428);
nor UO_1055 (O_1055,N_29723,N_28650);
or UO_1056 (O_1056,N_29986,N_29018);
or UO_1057 (O_1057,N_28761,N_28115);
xor UO_1058 (O_1058,N_29826,N_29115);
or UO_1059 (O_1059,N_28827,N_28819);
or UO_1060 (O_1060,N_29485,N_29471);
xnor UO_1061 (O_1061,N_29048,N_29125);
or UO_1062 (O_1062,N_29565,N_28530);
nor UO_1063 (O_1063,N_29502,N_29314);
or UO_1064 (O_1064,N_28494,N_29537);
and UO_1065 (O_1065,N_28527,N_28121);
and UO_1066 (O_1066,N_28278,N_28628);
and UO_1067 (O_1067,N_28249,N_29229);
nand UO_1068 (O_1068,N_29454,N_29679);
or UO_1069 (O_1069,N_29872,N_28469);
nand UO_1070 (O_1070,N_29318,N_29576);
or UO_1071 (O_1071,N_28435,N_28957);
xnor UO_1072 (O_1072,N_28794,N_28735);
and UO_1073 (O_1073,N_28942,N_29426);
nand UO_1074 (O_1074,N_29367,N_29541);
or UO_1075 (O_1075,N_29927,N_29437);
or UO_1076 (O_1076,N_29965,N_28793);
xnor UO_1077 (O_1077,N_28691,N_28847);
nand UO_1078 (O_1078,N_28276,N_28603);
nor UO_1079 (O_1079,N_28034,N_29435);
xor UO_1080 (O_1080,N_28240,N_28833);
and UO_1081 (O_1081,N_29191,N_28210);
xor UO_1082 (O_1082,N_29942,N_28783);
nor UO_1083 (O_1083,N_28646,N_28849);
xor UO_1084 (O_1084,N_28713,N_29106);
nor UO_1085 (O_1085,N_29187,N_28047);
nor UO_1086 (O_1086,N_28682,N_28839);
and UO_1087 (O_1087,N_29847,N_29497);
nor UO_1088 (O_1088,N_28772,N_28188);
xnor UO_1089 (O_1089,N_28281,N_28454);
and UO_1090 (O_1090,N_28800,N_29881);
or UO_1091 (O_1091,N_28102,N_28175);
nor UO_1092 (O_1092,N_29278,N_28381);
and UO_1093 (O_1093,N_29924,N_29039);
xor UO_1094 (O_1094,N_28636,N_29998);
or UO_1095 (O_1095,N_29897,N_28339);
and UO_1096 (O_1096,N_29027,N_29077);
nor UO_1097 (O_1097,N_28477,N_29772);
nand UO_1098 (O_1098,N_28798,N_28671);
or UO_1099 (O_1099,N_28430,N_29867);
nor UO_1100 (O_1100,N_29935,N_29542);
xnor UO_1101 (O_1101,N_28667,N_28288);
and UO_1102 (O_1102,N_29547,N_29861);
and UO_1103 (O_1103,N_28247,N_29876);
and UO_1104 (O_1104,N_28776,N_28370);
xnor UO_1105 (O_1105,N_28274,N_28782);
xor UO_1106 (O_1106,N_28355,N_28666);
or UO_1107 (O_1107,N_28783,N_29154);
and UO_1108 (O_1108,N_29332,N_29560);
nor UO_1109 (O_1109,N_29222,N_28636);
nor UO_1110 (O_1110,N_29011,N_29438);
nand UO_1111 (O_1111,N_29013,N_28623);
nand UO_1112 (O_1112,N_28554,N_28076);
or UO_1113 (O_1113,N_28008,N_29372);
and UO_1114 (O_1114,N_28010,N_28998);
xor UO_1115 (O_1115,N_29174,N_28930);
and UO_1116 (O_1116,N_29721,N_29201);
nor UO_1117 (O_1117,N_28326,N_28642);
nor UO_1118 (O_1118,N_29831,N_28998);
xnor UO_1119 (O_1119,N_29094,N_28529);
and UO_1120 (O_1120,N_28020,N_29234);
and UO_1121 (O_1121,N_28370,N_28811);
xor UO_1122 (O_1122,N_28489,N_28668);
nand UO_1123 (O_1123,N_28648,N_28872);
nor UO_1124 (O_1124,N_28104,N_29896);
nor UO_1125 (O_1125,N_29590,N_29063);
nor UO_1126 (O_1126,N_28685,N_29353);
nor UO_1127 (O_1127,N_29321,N_28143);
and UO_1128 (O_1128,N_29783,N_29983);
xor UO_1129 (O_1129,N_28963,N_28062);
xor UO_1130 (O_1130,N_29879,N_28462);
xnor UO_1131 (O_1131,N_29245,N_29790);
nand UO_1132 (O_1132,N_28820,N_28645);
nor UO_1133 (O_1133,N_29460,N_29687);
nor UO_1134 (O_1134,N_28151,N_28716);
nand UO_1135 (O_1135,N_28511,N_29417);
nand UO_1136 (O_1136,N_28141,N_29546);
nand UO_1137 (O_1137,N_29222,N_28525);
and UO_1138 (O_1138,N_28880,N_28234);
xor UO_1139 (O_1139,N_29983,N_29816);
nor UO_1140 (O_1140,N_29954,N_28257);
nor UO_1141 (O_1141,N_28054,N_28856);
and UO_1142 (O_1142,N_28290,N_28337);
or UO_1143 (O_1143,N_29658,N_28078);
xnor UO_1144 (O_1144,N_29890,N_29455);
nor UO_1145 (O_1145,N_28736,N_29528);
nor UO_1146 (O_1146,N_29496,N_28747);
nor UO_1147 (O_1147,N_29988,N_29334);
and UO_1148 (O_1148,N_29315,N_28281);
xor UO_1149 (O_1149,N_29218,N_29355);
or UO_1150 (O_1150,N_29868,N_28351);
xnor UO_1151 (O_1151,N_28580,N_29023);
and UO_1152 (O_1152,N_29648,N_28757);
or UO_1153 (O_1153,N_29186,N_28958);
nor UO_1154 (O_1154,N_29730,N_28307);
nand UO_1155 (O_1155,N_28455,N_29233);
nand UO_1156 (O_1156,N_29332,N_29408);
and UO_1157 (O_1157,N_29080,N_28777);
and UO_1158 (O_1158,N_29331,N_29932);
nor UO_1159 (O_1159,N_29434,N_29025);
xnor UO_1160 (O_1160,N_28437,N_29036);
nor UO_1161 (O_1161,N_28422,N_29690);
xnor UO_1162 (O_1162,N_28540,N_28739);
or UO_1163 (O_1163,N_29985,N_29905);
xnor UO_1164 (O_1164,N_29240,N_29748);
or UO_1165 (O_1165,N_28143,N_28386);
and UO_1166 (O_1166,N_29467,N_28667);
nor UO_1167 (O_1167,N_29148,N_28583);
nand UO_1168 (O_1168,N_29778,N_28586);
nand UO_1169 (O_1169,N_29666,N_29670);
nor UO_1170 (O_1170,N_28837,N_28485);
and UO_1171 (O_1171,N_28487,N_29131);
nand UO_1172 (O_1172,N_29251,N_29660);
or UO_1173 (O_1173,N_28743,N_29919);
nor UO_1174 (O_1174,N_28161,N_28860);
nand UO_1175 (O_1175,N_28136,N_28531);
and UO_1176 (O_1176,N_29086,N_28910);
nand UO_1177 (O_1177,N_29993,N_28113);
and UO_1178 (O_1178,N_29560,N_28712);
nand UO_1179 (O_1179,N_29081,N_28590);
or UO_1180 (O_1180,N_28988,N_28642);
nor UO_1181 (O_1181,N_28020,N_29624);
nor UO_1182 (O_1182,N_29760,N_29531);
nor UO_1183 (O_1183,N_28012,N_29932);
or UO_1184 (O_1184,N_29491,N_28308);
nand UO_1185 (O_1185,N_28497,N_28685);
nor UO_1186 (O_1186,N_28218,N_28666);
nor UO_1187 (O_1187,N_29721,N_29975);
and UO_1188 (O_1188,N_28324,N_29126);
nor UO_1189 (O_1189,N_29954,N_29000);
and UO_1190 (O_1190,N_28435,N_29462);
or UO_1191 (O_1191,N_28669,N_29716);
nand UO_1192 (O_1192,N_29280,N_28831);
or UO_1193 (O_1193,N_29658,N_28937);
xor UO_1194 (O_1194,N_29687,N_28082);
nand UO_1195 (O_1195,N_28525,N_28907);
xnor UO_1196 (O_1196,N_28696,N_29782);
xor UO_1197 (O_1197,N_28816,N_29084);
xnor UO_1198 (O_1198,N_29990,N_29477);
or UO_1199 (O_1199,N_29293,N_29186);
or UO_1200 (O_1200,N_28174,N_28231);
nand UO_1201 (O_1201,N_28673,N_28727);
nand UO_1202 (O_1202,N_29383,N_28735);
and UO_1203 (O_1203,N_28974,N_28154);
or UO_1204 (O_1204,N_28824,N_29560);
nor UO_1205 (O_1205,N_29687,N_29004);
and UO_1206 (O_1206,N_29980,N_28899);
nand UO_1207 (O_1207,N_28296,N_29363);
or UO_1208 (O_1208,N_29464,N_29164);
and UO_1209 (O_1209,N_29991,N_28530);
or UO_1210 (O_1210,N_28027,N_29552);
nand UO_1211 (O_1211,N_29940,N_28009);
nand UO_1212 (O_1212,N_29505,N_28497);
nor UO_1213 (O_1213,N_28041,N_29670);
nor UO_1214 (O_1214,N_28267,N_29503);
and UO_1215 (O_1215,N_29942,N_28612);
nand UO_1216 (O_1216,N_28940,N_28388);
and UO_1217 (O_1217,N_29154,N_28817);
and UO_1218 (O_1218,N_29003,N_28127);
nor UO_1219 (O_1219,N_28599,N_29503);
xnor UO_1220 (O_1220,N_28193,N_28819);
nand UO_1221 (O_1221,N_29342,N_28919);
and UO_1222 (O_1222,N_28851,N_29701);
nand UO_1223 (O_1223,N_28230,N_29805);
nand UO_1224 (O_1224,N_29370,N_28181);
nand UO_1225 (O_1225,N_28644,N_28334);
nor UO_1226 (O_1226,N_28149,N_28048);
or UO_1227 (O_1227,N_29562,N_28170);
xor UO_1228 (O_1228,N_28047,N_28704);
and UO_1229 (O_1229,N_29095,N_29426);
nor UO_1230 (O_1230,N_28393,N_29527);
and UO_1231 (O_1231,N_29403,N_29140);
or UO_1232 (O_1232,N_29107,N_29298);
or UO_1233 (O_1233,N_28539,N_28504);
and UO_1234 (O_1234,N_29636,N_28646);
or UO_1235 (O_1235,N_28901,N_28400);
xnor UO_1236 (O_1236,N_28604,N_29135);
and UO_1237 (O_1237,N_29858,N_28869);
xor UO_1238 (O_1238,N_29487,N_28527);
nand UO_1239 (O_1239,N_29330,N_29568);
or UO_1240 (O_1240,N_28846,N_28287);
and UO_1241 (O_1241,N_29137,N_28402);
nand UO_1242 (O_1242,N_29528,N_29285);
or UO_1243 (O_1243,N_28110,N_29339);
xor UO_1244 (O_1244,N_29772,N_29156);
xnor UO_1245 (O_1245,N_29341,N_29380);
nor UO_1246 (O_1246,N_29034,N_29187);
and UO_1247 (O_1247,N_29387,N_29532);
and UO_1248 (O_1248,N_29532,N_28192);
nand UO_1249 (O_1249,N_29659,N_28848);
xnor UO_1250 (O_1250,N_28320,N_29195);
nor UO_1251 (O_1251,N_29077,N_28659);
and UO_1252 (O_1252,N_29098,N_28192);
and UO_1253 (O_1253,N_29853,N_28570);
nand UO_1254 (O_1254,N_29389,N_29577);
or UO_1255 (O_1255,N_28220,N_29863);
xor UO_1256 (O_1256,N_28167,N_28065);
and UO_1257 (O_1257,N_28812,N_28509);
and UO_1258 (O_1258,N_29495,N_28949);
nor UO_1259 (O_1259,N_29096,N_29330);
or UO_1260 (O_1260,N_28689,N_29579);
nand UO_1261 (O_1261,N_29029,N_29315);
nand UO_1262 (O_1262,N_28823,N_28401);
xnor UO_1263 (O_1263,N_28584,N_28525);
xnor UO_1264 (O_1264,N_29270,N_29447);
or UO_1265 (O_1265,N_29928,N_29140);
and UO_1266 (O_1266,N_29491,N_29486);
nand UO_1267 (O_1267,N_28253,N_28264);
or UO_1268 (O_1268,N_28932,N_28326);
nand UO_1269 (O_1269,N_29389,N_28373);
and UO_1270 (O_1270,N_29832,N_29794);
nor UO_1271 (O_1271,N_29522,N_29062);
or UO_1272 (O_1272,N_29269,N_29544);
nor UO_1273 (O_1273,N_29868,N_29304);
nand UO_1274 (O_1274,N_28239,N_28073);
xor UO_1275 (O_1275,N_29084,N_28306);
nand UO_1276 (O_1276,N_29416,N_28517);
nand UO_1277 (O_1277,N_29094,N_28130);
nand UO_1278 (O_1278,N_29239,N_28952);
nand UO_1279 (O_1279,N_29994,N_28200);
nand UO_1280 (O_1280,N_29227,N_29901);
and UO_1281 (O_1281,N_28021,N_28423);
xnor UO_1282 (O_1282,N_28909,N_28136);
nand UO_1283 (O_1283,N_28888,N_29948);
xor UO_1284 (O_1284,N_28581,N_29822);
or UO_1285 (O_1285,N_29282,N_29334);
or UO_1286 (O_1286,N_28521,N_29959);
xnor UO_1287 (O_1287,N_28407,N_29289);
and UO_1288 (O_1288,N_29749,N_28324);
nand UO_1289 (O_1289,N_29481,N_29717);
or UO_1290 (O_1290,N_29634,N_29744);
nor UO_1291 (O_1291,N_28063,N_29734);
xnor UO_1292 (O_1292,N_29126,N_29575);
and UO_1293 (O_1293,N_29078,N_28803);
nand UO_1294 (O_1294,N_28647,N_29858);
nor UO_1295 (O_1295,N_29281,N_29650);
nand UO_1296 (O_1296,N_28144,N_28636);
and UO_1297 (O_1297,N_28119,N_28033);
or UO_1298 (O_1298,N_28319,N_28427);
xnor UO_1299 (O_1299,N_29299,N_28290);
xor UO_1300 (O_1300,N_28205,N_28033);
or UO_1301 (O_1301,N_28107,N_28695);
nand UO_1302 (O_1302,N_29245,N_29957);
xnor UO_1303 (O_1303,N_28330,N_29628);
nand UO_1304 (O_1304,N_28262,N_29006);
or UO_1305 (O_1305,N_28278,N_29284);
and UO_1306 (O_1306,N_29269,N_29975);
or UO_1307 (O_1307,N_29988,N_28127);
nor UO_1308 (O_1308,N_29746,N_28725);
nor UO_1309 (O_1309,N_29881,N_28298);
nand UO_1310 (O_1310,N_28606,N_28038);
and UO_1311 (O_1311,N_29709,N_28344);
or UO_1312 (O_1312,N_28460,N_28848);
and UO_1313 (O_1313,N_28463,N_29839);
nand UO_1314 (O_1314,N_29964,N_28908);
and UO_1315 (O_1315,N_29897,N_29964);
nor UO_1316 (O_1316,N_28334,N_29489);
xnor UO_1317 (O_1317,N_29578,N_28032);
and UO_1318 (O_1318,N_29218,N_28310);
and UO_1319 (O_1319,N_29775,N_29223);
nor UO_1320 (O_1320,N_29869,N_29628);
nand UO_1321 (O_1321,N_28001,N_28405);
and UO_1322 (O_1322,N_28443,N_29747);
nand UO_1323 (O_1323,N_28930,N_29137);
and UO_1324 (O_1324,N_28627,N_28035);
xnor UO_1325 (O_1325,N_28869,N_28334);
xor UO_1326 (O_1326,N_28495,N_28999);
xor UO_1327 (O_1327,N_29861,N_29998);
or UO_1328 (O_1328,N_28620,N_29220);
xor UO_1329 (O_1329,N_29681,N_28060);
xor UO_1330 (O_1330,N_29763,N_28536);
xor UO_1331 (O_1331,N_28783,N_28800);
and UO_1332 (O_1332,N_29171,N_28720);
or UO_1333 (O_1333,N_29898,N_29025);
or UO_1334 (O_1334,N_29602,N_29239);
and UO_1335 (O_1335,N_29868,N_28343);
or UO_1336 (O_1336,N_29269,N_28932);
nand UO_1337 (O_1337,N_28161,N_28155);
and UO_1338 (O_1338,N_29577,N_28467);
or UO_1339 (O_1339,N_29026,N_29141);
xnor UO_1340 (O_1340,N_29747,N_28839);
nand UO_1341 (O_1341,N_29288,N_29062);
xnor UO_1342 (O_1342,N_29735,N_28483);
and UO_1343 (O_1343,N_29792,N_28232);
and UO_1344 (O_1344,N_29156,N_28509);
nor UO_1345 (O_1345,N_29581,N_29166);
nand UO_1346 (O_1346,N_28162,N_28120);
nand UO_1347 (O_1347,N_28669,N_29033);
nor UO_1348 (O_1348,N_29012,N_29671);
nand UO_1349 (O_1349,N_29362,N_28688);
nand UO_1350 (O_1350,N_29177,N_28954);
or UO_1351 (O_1351,N_28352,N_28038);
and UO_1352 (O_1352,N_28683,N_28229);
nand UO_1353 (O_1353,N_28594,N_28313);
nor UO_1354 (O_1354,N_28757,N_29317);
nor UO_1355 (O_1355,N_29017,N_28694);
xor UO_1356 (O_1356,N_29969,N_29897);
and UO_1357 (O_1357,N_29070,N_28501);
and UO_1358 (O_1358,N_28155,N_29268);
or UO_1359 (O_1359,N_28269,N_29831);
and UO_1360 (O_1360,N_28274,N_29267);
and UO_1361 (O_1361,N_28689,N_28335);
or UO_1362 (O_1362,N_29836,N_28094);
nor UO_1363 (O_1363,N_28251,N_28001);
nand UO_1364 (O_1364,N_29226,N_29011);
xnor UO_1365 (O_1365,N_28404,N_29354);
and UO_1366 (O_1366,N_29013,N_29427);
xor UO_1367 (O_1367,N_28885,N_29748);
and UO_1368 (O_1368,N_28091,N_29751);
nor UO_1369 (O_1369,N_28425,N_28215);
xnor UO_1370 (O_1370,N_28220,N_28508);
xor UO_1371 (O_1371,N_28240,N_28446);
or UO_1372 (O_1372,N_29673,N_28544);
and UO_1373 (O_1373,N_29671,N_29492);
and UO_1374 (O_1374,N_29874,N_29207);
and UO_1375 (O_1375,N_29072,N_28617);
nand UO_1376 (O_1376,N_29986,N_28266);
and UO_1377 (O_1377,N_28101,N_29672);
nor UO_1378 (O_1378,N_29698,N_28488);
nor UO_1379 (O_1379,N_28471,N_29978);
and UO_1380 (O_1380,N_28989,N_28519);
xor UO_1381 (O_1381,N_29424,N_28615);
xnor UO_1382 (O_1382,N_28172,N_29107);
nand UO_1383 (O_1383,N_28094,N_28226);
or UO_1384 (O_1384,N_29240,N_29534);
xnor UO_1385 (O_1385,N_28977,N_29425);
xor UO_1386 (O_1386,N_29043,N_28771);
and UO_1387 (O_1387,N_29624,N_29463);
xor UO_1388 (O_1388,N_29175,N_28298);
nand UO_1389 (O_1389,N_28560,N_29116);
and UO_1390 (O_1390,N_28169,N_28319);
nor UO_1391 (O_1391,N_28243,N_29481);
and UO_1392 (O_1392,N_29064,N_28747);
or UO_1393 (O_1393,N_28184,N_28788);
nand UO_1394 (O_1394,N_29671,N_28258);
or UO_1395 (O_1395,N_28765,N_28498);
or UO_1396 (O_1396,N_29046,N_28852);
and UO_1397 (O_1397,N_28606,N_29696);
nor UO_1398 (O_1398,N_29532,N_28475);
nand UO_1399 (O_1399,N_29166,N_28267);
nand UO_1400 (O_1400,N_29162,N_28069);
nor UO_1401 (O_1401,N_29018,N_28167);
and UO_1402 (O_1402,N_29194,N_28207);
or UO_1403 (O_1403,N_29533,N_29424);
xnor UO_1404 (O_1404,N_29127,N_29750);
nand UO_1405 (O_1405,N_28288,N_28012);
nand UO_1406 (O_1406,N_28731,N_29221);
xnor UO_1407 (O_1407,N_29232,N_29561);
nor UO_1408 (O_1408,N_29764,N_29196);
or UO_1409 (O_1409,N_29907,N_29746);
and UO_1410 (O_1410,N_28028,N_28881);
xor UO_1411 (O_1411,N_29525,N_29465);
nor UO_1412 (O_1412,N_28485,N_28441);
or UO_1413 (O_1413,N_28920,N_29187);
or UO_1414 (O_1414,N_28657,N_29882);
and UO_1415 (O_1415,N_29285,N_28919);
nand UO_1416 (O_1416,N_29823,N_28723);
nand UO_1417 (O_1417,N_28157,N_28899);
nand UO_1418 (O_1418,N_29708,N_28534);
nor UO_1419 (O_1419,N_29579,N_28824);
xnor UO_1420 (O_1420,N_29126,N_28599);
nor UO_1421 (O_1421,N_29462,N_29720);
xor UO_1422 (O_1422,N_29115,N_28269);
nor UO_1423 (O_1423,N_29037,N_28967);
or UO_1424 (O_1424,N_29547,N_29443);
and UO_1425 (O_1425,N_28137,N_28833);
or UO_1426 (O_1426,N_28362,N_29245);
and UO_1427 (O_1427,N_28599,N_29787);
nor UO_1428 (O_1428,N_28624,N_28245);
nor UO_1429 (O_1429,N_29755,N_28209);
or UO_1430 (O_1430,N_29421,N_29233);
xor UO_1431 (O_1431,N_28010,N_28505);
or UO_1432 (O_1432,N_28068,N_28950);
nor UO_1433 (O_1433,N_28681,N_29550);
xnor UO_1434 (O_1434,N_29540,N_28903);
nand UO_1435 (O_1435,N_28639,N_28458);
nor UO_1436 (O_1436,N_29075,N_29932);
nand UO_1437 (O_1437,N_29098,N_28994);
xnor UO_1438 (O_1438,N_29566,N_29164);
nand UO_1439 (O_1439,N_29895,N_29106);
xnor UO_1440 (O_1440,N_28349,N_28623);
and UO_1441 (O_1441,N_28126,N_28909);
nand UO_1442 (O_1442,N_29586,N_28409);
xor UO_1443 (O_1443,N_28064,N_29745);
nand UO_1444 (O_1444,N_29880,N_28372);
or UO_1445 (O_1445,N_28008,N_29338);
nor UO_1446 (O_1446,N_29976,N_28842);
and UO_1447 (O_1447,N_28908,N_29000);
nor UO_1448 (O_1448,N_29930,N_29205);
nand UO_1449 (O_1449,N_28336,N_29208);
and UO_1450 (O_1450,N_28511,N_29905);
xnor UO_1451 (O_1451,N_29028,N_28918);
nor UO_1452 (O_1452,N_29078,N_28771);
xnor UO_1453 (O_1453,N_29651,N_29160);
nor UO_1454 (O_1454,N_29969,N_29299);
nor UO_1455 (O_1455,N_28482,N_28710);
nor UO_1456 (O_1456,N_28724,N_29927);
or UO_1457 (O_1457,N_28559,N_29629);
or UO_1458 (O_1458,N_29098,N_29710);
nor UO_1459 (O_1459,N_28572,N_29460);
xor UO_1460 (O_1460,N_29635,N_29420);
and UO_1461 (O_1461,N_29701,N_29409);
nor UO_1462 (O_1462,N_28395,N_29172);
xor UO_1463 (O_1463,N_28248,N_28220);
and UO_1464 (O_1464,N_29264,N_28146);
and UO_1465 (O_1465,N_28939,N_28318);
or UO_1466 (O_1466,N_28461,N_28759);
nand UO_1467 (O_1467,N_29433,N_28296);
nand UO_1468 (O_1468,N_28913,N_29343);
xor UO_1469 (O_1469,N_29357,N_28101);
and UO_1470 (O_1470,N_28362,N_28646);
xnor UO_1471 (O_1471,N_29665,N_28915);
nor UO_1472 (O_1472,N_29436,N_29249);
and UO_1473 (O_1473,N_28820,N_28368);
xnor UO_1474 (O_1474,N_28215,N_29850);
and UO_1475 (O_1475,N_29332,N_28899);
or UO_1476 (O_1476,N_28764,N_29769);
and UO_1477 (O_1477,N_28729,N_28505);
xnor UO_1478 (O_1478,N_29105,N_28360);
xnor UO_1479 (O_1479,N_29196,N_29585);
nor UO_1480 (O_1480,N_29418,N_29683);
nor UO_1481 (O_1481,N_28940,N_29832);
and UO_1482 (O_1482,N_28711,N_28896);
xor UO_1483 (O_1483,N_29680,N_29965);
nand UO_1484 (O_1484,N_28630,N_29275);
or UO_1485 (O_1485,N_28198,N_29890);
and UO_1486 (O_1486,N_29054,N_28992);
xnor UO_1487 (O_1487,N_28308,N_29002);
nand UO_1488 (O_1488,N_28006,N_28859);
and UO_1489 (O_1489,N_29362,N_28391);
xnor UO_1490 (O_1490,N_28155,N_28079);
and UO_1491 (O_1491,N_29407,N_29854);
nor UO_1492 (O_1492,N_28672,N_29152);
or UO_1493 (O_1493,N_28390,N_29302);
xor UO_1494 (O_1494,N_29428,N_28462);
nor UO_1495 (O_1495,N_28972,N_29788);
nand UO_1496 (O_1496,N_28442,N_29895);
xor UO_1497 (O_1497,N_29376,N_28906);
nand UO_1498 (O_1498,N_28990,N_29428);
xor UO_1499 (O_1499,N_28680,N_28154);
or UO_1500 (O_1500,N_28172,N_28738);
nor UO_1501 (O_1501,N_29219,N_28971);
nand UO_1502 (O_1502,N_29879,N_28752);
or UO_1503 (O_1503,N_29945,N_28908);
and UO_1504 (O_1504,N_29641,N_29695);
nand UO_1505 (O_1505,N_29487,N_29999);
and UO_1506 (O_1506,N_28852,N_28542);
xnor UO_1507 (O_1507,N_28032,N_28270);
nor UO_1508 (O_1508,N_29002,N_28602);
xnor UO_1509 (O_1509,N_28533,N_28563);
and UO_1510 (O_1510,N_28702,N_29961);
or UO_1511 (O_1511,N_28824,N_28719);
nand UO_1512 (O_1512,N_29623,N_29812);
nor UO_1513 (O_1513,N_28366,N_29553);
xnor UO_1514 (O_1514,N_29149,N_29378);
or UO_1515 (O_1515,N_29527,N_29621);
nand UO_1516 (O_1516,N_28210,N_28551);
and UO_1517 (O_1517,N_29892,N_29130);
nor UO_1518 (O_1518,N_28548,N_29220);
or UO_1519 (O_1519,N_29810,N_28196);
xnor UO_1520 (O_1520,N_29993,N_29872);
xor UO_1521 (O_1521,N_29273,N_28839);
xnor UO_1522 (O_1522,N_29339,N_29850);
nor UO_1523 (O_1523,N_28987,N_29478);
nand UO_1524 (O_1524,N_29652,N_29012);
nor UO_1525 (O_1525,N_28934,N_28272);
or UO_1526 (O_1526,N_29083,N_29982);
or UO_1527 (O_1527,N_29956,N_29441);
nand UO_1528 (O_1528,N_28314,N_29393);
nand UO_1529 (O_1529,N_28579,N_28089);
or UO_1530 (O_1530,N_29202,N_28914);
nand UO_1531 (O_1531,N_28195,N_28130);
nor UO_1532 (O_1532,N_28784,N_29331);
nor UO_1533 (O_1533,N_28803,N_28188);
or UO_1534 (O_1534,N_29571,N_28568);
and UO_1535 (O_1535,N_28496,N_28233);
nor UO_1536 (O_1536,N_28540,N_28581);
nand UO_1537 (O_1537,N_29610,N_28182);
and UO_1538 (O_1538,N_29189,N_29061);
or UO_1539 (O_1539,N_28901,N_29525);
or UO_1540 (O_1540,N_29209,N_29571);
xor UO_1541 (O_1541,N_29467,N_29161);
and UO_1542 (O_1542,N_29147,N_29960);
xnor UO_1543 (O_1543,N_29439,N_29015);
nand UO_1544 (O_1544,N_28084,N_29840);
or UO_1545 (O_1545,N_28471,N_29086);
xor UO_1546 (O_1546,N_28371,N_28959);
xor UO_1547 (O_1547,N_29075,N_29698);
nor UO_1548 (O_1548,N_29124,N_28209);
or UO_1549 (O_1549,N_29768,N_29307);
xnor UO_1550 (O_1550,N_29763,N_28457);
nand UO_1551 (O_1551,N_28788,N_29749);
xor UO_1552 (O_1552,N_28722,N_28759);
nor UO_1553 (O_1553,N_28527,N_28874);
or UO_1554 (O_1554,N_28871,N_29074);
or UO_1555 (O_1555,N_29550,N_28965);
and UO_1556 (O_1556,N_28561,N_29263);
nor UO_1557 (O_1557,N_29039,N_28815);
xnor UO_1558 (O_1558,N_28778,N_28618);
nor UO_1559 (O_1559,N_29108,N_28348);
nand UO_1560 (O_1560,N_29676,N_29968);
xnor UO_1561 (O_1561,N_28900,N_29690);
nor UO_1562 (O_1562,N_28684,N_28844);
and UO_1563 (O_1563,N_29994,N_28038);
or UO_1564 (O_1564,N_29802,N_29398);
and UO_1565 (O_1565,N_28128,N_28520);
nor UO_1566 (O_1566,N_28171,N_28385);
nand UO_1567 (O_1567,N_28675,N_29032);
and UO_1568 (O_1568,N_28524,N_28793);
xor UO_1569 (O_1569,N_29943,N_29922);
and UO_1570 (O_1570,N_29763,N_29477);
nor UO_1571 (O_1571,N_28716,N_29960);
and UO_1572 (O_1572,N_28748,N_28490);
and UO_1573 (O_1573,N_28714,N_29066);
nand UO_1574 (O_1574,N_28198,N_28096);
xor UO_1575 (O_1575,N_29236,N_28406);
nor UO_1576 (O_1576,N_28846,N_28803);
or UO_1577 (O_1577,N_28536,N_28241);
or UO_1578 (O_1578,N_29690,N_28719);
xor UO_1579 (O_1579,N_28770,N_28258);
xor UO_1580 (O_1580,N_28585,N_29450);
nor UO_1581 (O_1581,N_29497,N_28743);
xnor UO_1582 (O_1582,N_28188,N_28249);
xnor UO_1583 (O_1583,N_28480,N_28399);
or UO_1584 (O_1584,N_29945,N_28827);
nor UO_1585 (O_1585,N_29763,N_28497);
or UO_1586 (O_1586,N_29303,N_28942);
xor UO_1587 (O_1587,N_28686,N_28065);
xor UO_1588 (O_1588,N_29506,N_28322);
or UO_1589 (O_1589,N_29114,N_29725);
nor UO_1590 (O_1590,N_29672,N_29150);
and UO_1591 (O_1591,N_28310,N_28306);
and UO_1592 (O_1592,N_29767,N_28608);
or UO_1593 (O_1593,N_28893,N_28392);
nor UO_1594 (O_1594,N_28342,N_29162);
nand UO_1595 (O_1595,N_28256,N_28509);
nor UO_1596 (O_1596,N_28800,N_28449);
xor UO_1597 (O_1597,N_28095,N_28294);
nand UO_1598 (O_1598,N_29420,N_28153);
or UO_1599 (O_1599,N_28657,N_28468);
xnor UO_1600 (O_1600,N_28529,N_29734);
xor UO_1601 (O_1601,N_28201,N_28964);
nand UO_1602 (O_1602,N_29015,N_29829);
and UO_1603 (O_1603,N_28188,N_28683);
xnor UO_1604 (O_1604,N_28063,N_28971);
xnor UO_1605 (O_1605,N_29870,N_28764);
xor UO_1606 (O_1606,N_28901,N_28860);
and UO_1607 (O_1607,N_29906,N_29851);
nor UO_1608 (O_1608,N_29047,N_29855);
nor UO_1609 (O_1609,N_29038,N_28007);
nand UO_1610 (O_1610,N_29361,N_29910);
xor UO_1611 (O_1611,N_29862,N_28967);
or UO_1612 (O_1612,N_28724,N_28493);
nor UO_1613 (O_1613,N_29565,N_29765);
xor UO_1614 (O_1614,N_28363,N_29862);
nor UO_1615 (O_1615,N_28256,N_28475);
and UO_1616 (O_1616,N_29062,N_29802);
or UO_1617 (O_1617,N_29650,N_28638);
xor UO_1618 (O_1618,N_29033,N_28461);
nor UO_1619 (O_1619,N_28277,N_28735);
or UO_1620 (O_1620,N_29933,N_29242);
nor UO_1621 (O_1621,N_29501,N_28255);
nand UO_1622 (O_1622,N_28479,N_28713);
or UO_1623 (O_1623,N_28128,N_28990);
or UO_1624 (O_1624,N_29714,N_29087);
xor UO_1625 (O_1625,N_29349,N_29051);
xnor UO_1626 (O_1626,N_28950,N_29066);
xnor UO_1627 (O_1627,N_29238,N_28672);
nor UO_1628 (O_1628,N_29753,N_29955);
nand UO_1629 (O_1629,N_28847,N_28429);
nor UO_1630 (O_1630,N_29349,N_28187);
nand UO_1631 (O_1631,N_29398,N_29271);
or UO_1632 (O_1632,N_29322,N_29786);
xnor UO_1633 (O_1633,N_29355,N_29562);
and UO_1634 (O_1634,N_29064,N_29167);
xnor UO_1635 (O_1635,N_28072,N_29500);
or UO_1636 (O_1636,N_28521,N_28016);
or UO_1637 (O_1637,N_28946,N_28987);
nand UO_1638 (O_1638,N_29368,N_29282);
and UO_1639 (O_1639,N_28016,N_28479);
and UO_1640 (O_1640,N_29411,N_28794);
nand UO_1641 (O_1641,N_28563,N_28230);
and UO_1642 (O_1642,N_28713,N_28520);
nor UO_1643 (O_1643,N_28703,N_29442);
and UO_1644 (O_1644,N_28042,N_29587);
xnor UO_1645 (O_1645,N_29547,N_29770);
and UO_1646 (O_1646,N_28490,N_29800);
nor UO_1647 (O_1647,N_29706,N_29037);
xor UO_1648 (O_1648,N_29666,N_28601);
nand UO_1649 (O_1649,N_29863,N_28933);
or UO_1650 (O_1650,N_28368,N_28980);
nand UO_1651 (O_1651,N_28248,N_29987);
nand UO_1652 (O_1652,N_29620,N_29206);
or UO_1653 (O_1653,N_29759,N_28378);
and UO_1654 (O_1654,N_28607,N_29706);
or UO_1655 (O_1655,N_28968,N_28280);
nor UO_1656 (O_1656,N_29745,N_29104);
nor UO_1657 (O_1657,N_29673,N_29485);
nor UO_1658 (O_1658,N_28511,N_28046);
or UO_1659 (O_1659,N_28508,N_29230);
and UO_1660 (O_1660,N_28849,N_28623);
nor UO_1661 (O_1661,N_28257,N_29792);
xnor UO_1662 (O_1662,N_28033,N_29270);
and UO_1663 (O_1663,N_29253,N_28611);
or UO_1664 (O_1664,N_28415,N_28079);
xor UO_1665 (O_1665,N_28899,N_28038);
and UO_1666 (O_1666,N_28171,N_29690);
or UO_1667 (O_1667,N_29863,N_28736);
nand UO_1668 (O_1668,N_29736,N_29912);
xnor UO_1669 (O_1669,N_28435,N_28466);
nand UO_1670 (O_1670,N_28206,N_28600);
xor UO_1671 (O_1671,N_29221,N_29745);
and UO_1672 (O_1672,N_28092,N_29010);
nand UO_1673 (O_1673,N_29125,N_29907);
xnor UO_1674 (O_1674,N_29631,N_29738);
xnor UO_1675 (O_1675,N_29366,N_28286);
nand UO_1676 (O_1676,N_28363,N_28354);
nand UO_1677 (O_1677,N_28644,N_28791);
and UO_1678 (O_1678,N_29017,N_28422);
nand UO_1679 (O_1679,N_29955,N_29340);
nor UO_1680 (O_1680,N_28872,N_29134);
nand UO_1681 (O_1681,N_29840,N_29770);
nand UO_1682 (O_1682,N_29110,N_28548);
nand UO_1683 (O_1683,N_29860,N_29215);
nor UO_1684 (O_1684,N_29186,N_28217);
and UO_1685 (O_1685,N_28543,N_29847);
nand UO_1686 (O_1686,N_28186,N_29320);
nand UO_1687 (O_1687,N_28834,N_28791);
xnor UO_1688 (O_1688,N_28565,N_29266);
or UO_1689 (O_1689,N_28619,N_29914);
xnor UO_1690 (O_1690,N_28001,N_28772);
and UO_1691 (O_1691,N_29678,N_28970);
nand UO_1692 (O_1692,N_29080,N_28618);
nand UO_1693 (O_1693,N_28854,N_28124);
nor UO_1694 (O_1694,N_28315,N_29516);
nor UO_1695 (O_1695,N_28657,N_28656);
and UO_1696 (O_1696,N_29402,N_28571);
and UO_1697 (O_1697,N_29147,N_28567);
and UO_1698 (O_1698,N_28782,N_29123);
or UO_1699 (O_1699,N_29491,N_29218);
or UO_1700 (O_1700,N_28253,N_29849);
and UO_1701 (O_1701,N_29355,N_28406);
and UO_1702 (O_1702,N_28216,N_28484);
and UO_1703 (O_1703,N_28001,N_29384);
or UO_1704 (O_1704,N_29981,N_29725);
and UO_1705 (O_1705,N_28615,N_28172);
nand UO_1706 (O_1706,N_28136,N_29399);
xnor UO_1707 (O_1707,N_28235,N_28046);
nor UO_1708 (O_1708,N_28343,N_28811);
or UO_1709 (O_1709,N_28909,N_29875);
nand UO_1710 (O_1710,N_28948,N_28229);
or UO_1711 (O_1711,N_29073,N_29978);
and UO_1712 (O_1712,N_29386,N_29041);
nand UO_1713 (O_1713,N_29867,N_29246);
or UO_1714 (O_1714,N_29067,N_29359);
nand UO_1715 (O_1715,N_29430,N_29550);
nand UO_1716 (O_1716,N_29017,N_28135);
or UO_1717 (O_1717,N_29253,N_29111);
nor UO_1718 (O_1718,N_29729,N_28793);
or UO_1719 (O_1719,N_29297,N_28139);
nor UO_1720 (O_1720,N_28527,N_28324);
nand UO_1721 (O_1721,N_28379,N_29117);
xnor UO_1722 (O_1722,N_28851,N_29569);
nand UO_1723 (O_1723,N_29808,N_29053);
or UO_1724 (O_1724,N_29404,N_28458);
xor UO_1725 (O_1725,N_29562,N_29658);
xnor UO_1726 (O_1726,N_29359,N_29757);
or UO_1727 (O_1727,N_28920,N_28966);
nor UO_1728 (O_1728,N_28759,N_29238);
or UO_1729 (O_1729,N_29174,N_29564);
nor UO_1730 (O_1730,N_29584,N_28065);
and UO_1731 (O_1731,N_28084,N_28390);
or UO_1732 (O_1732,N_28568,N_29956);
xnor UO_1733 (O_1733,N_29772,N_28960);
or UO_1734 (O_1734,N_29814,N_29204);
xnor UO_1735 (O_1735,N_29831,N_28504);
or UO_1736 (O_1736,N_29104,N_29476);
xor UO_1737 (O_1737,N_28983,N_28689);
xor UO_1738 (O_1738,N_29390,N_29943);
or UO_1739 (O_1739,N_28315,N_29621);
nor UO_1740 (O_1740,N_28570,N_29593);
xnor UO_1741 (O_1741,N_28892,N_28877);
nand UO_1742 (O_1742,N_28603,N_28006);
or UO_1743 (O_1743,N_29025,N_28290);
and UO_1744 (O_1744,N_29370,N_29762);
nor UO_1745 (O_1745,N_28256,N_29429);
and UO_1746 (O_1746,N_29465,N_28083);
and UO_1747 (O_1747,N_28851,N_29430);
nand UO_1748 (O_1748,N_28038,N_28361);
nand UO_1749 (O_1749,N_28535,N_28262);
or UO_1750 (O_1750,N_29914,N_28419);
and UO_1751 (O_1751,N_28578,N_28000);
or UO_1752 (O_1752,N_29671,N_29563);
or UO_1753 (O_1753,N_29013,N_28224);
and UO_1754 (O_1754,N_29935,N_29435);
and UO_1755 (O_1755,N_29620,N_29852);
and UO_1756 (O_1756,N_29558,N_28920);
or UO_1757 (O_1757,N_28331,N_29184);
or UO_1758 (O_1758,N_28615,N_28950);
nor UO_1759 (O_1759,N_29442,N_28254);
nor UO_1760 (O_1760,N_29560,N_28030);
and UO_1761 (O_1761,N_29244,N_28494);
and UO_1762 (O_1762,N_29860,N_29227);
xor UO_1763 (O_1763,N_28509,N_28156);
or UO_1764 (O_1764,N_29258,N_29345);
nand UO_1765 (O_1765,N_29470,N_29807);
and UO_1766 (O_1766,N_28959,N_28127);
nand UO_1767 (O_1767,N_29804,N_29416);
nor UO_1768 (O_1768,N_29772,N_28911);
nor UO_1769 (O_1769,N_28506,N_28270);
xor UO_1770 (O_1770,N_29030,N_29795);
xor UO_1771 (O_1771,N_28729,N_28167);
nand UO_1772 (O_1772,N_29044,N_29640);
or UO_1773 (O_1773,N_29791,N_28414);
nand UO_1774 (O_1774,N_28475,N_28353);
nand UO_1775 (O_1775,N_29328,N_28584);
xor UO_1776 (O_1776,N_29411,N_29268);
xnor UO_1777 (O_1777,N_28315,N_29351);
nand UO_1778 (O_1778,N_29282,N_28226);
xor UO_1779 (O_1779,N_29893,N_28652);
and UO_1780 (O_1780,N_29001,N_29242);
or UO_1781 (O_1781,N_28326,N_29666);
xnor UO_1782 (O_1782,N_28254,N_29651);
nor UO_1783 (O_1783,N_29991,N_29695);
xor UO_1784 (O_1784,N_29201,N_29328);
nand UO_1785 (O_1785,N_28400,N_29188);
or UO_1786 (O_1786,N_28931,N_29872);
and UO_1787 (O_1787,N_28232,N_28616);
nor UO_1788 (O_1788,N_29798,N_28621);
nor UO_1789 (O_1789,N_28841,N_28229);
nor UO_1790 (O_1790,N_28985,N_29052);
or UO_1791 (O_1791,N_29606,N_28000);
nand UO_1792 (O_1792,N_28885,N_28968);
and UO_1793 (O_1793,N_28083,N_29883);
and UO_1794 (O_1794,N_29756,N_28963);
or UO_1795 (O_1795,N_28841,N_29585);
or UO_1796 (O_1796,N_28273,N_28511);
nand UO_1797 (O_1797,N_28638,N_28408);
nand UO_1798 (O_1798,N_28136,N_29538);
xor UO_1799 (O_1799,N_28908,N_29895);
nand UO_1800 (O_1800,N_29436,N_28156);
nand UO_1801 (O_1801,N_28323,N_28769);
and UO_1802 (O_1802,N_29754,N_28345);
xor UO_1803 (O_1803,N_29153,N_29526);
nand UO_1804 (O_1804,N_28954,N_29904);
xor UO_1805 (O_1805,N_29707,N_29695);
and UO_1806 (O_1806,N_28184,N_29132);
nor UO_1807 (O_1807,N_28674,N_29167);
or UO_1808 (O_1808,N_29116,N_28913);
nand UO_1809 (O_1809,N_28051,N_28656);
nor UO_1810 (O_1810,N_28405,N_28905);
nand UO_1811 (O_1811,N_29120,N_29392);
nand UO_1812 (O_1812,N_28398,N_28579);
and UO_1813 (O_1813,N_29565,N_29201);
nand UO_1814 (O_1814,N_28399,N_28056);
or UO_1815 (O_1815,N_29255,N_29364);
or UO_1816 (O_1816,N_29522,N_29459);
nand UO_1817 (O_1817,N_29071,N_28598);
and UO_1818 (O_1818,N_29976,N_28443);
nand UO_1819 (O_1819,N_28290,N_29578);
xor UO_1820 (O_1820,N_29343,N_29730);
nor UO_1821 (O_1821,N_29058,N_29084);
and UO_1822 (O_1822,N_29381,N_28395);
and UO_1823 (O_1823,N_28136,N_28997);
nand UO_1824 (O_1824,N_28239,N_28719);
xnor UO_1825 (O_1825,N_28503,N_29114);
nand UO_1826 (O_1826,N_28095,N_29457);
nor UO_1827 (O_1827,N_29190,N_29278);
or UO_1828 (O_1828,N_29790,N_29177);
xor UO_1829 (O_1829,N_28786,N_28553);
or UO_1830 (O_1830,N_28166,N_29646);
or UO_1831 (O_1831,N_29151,N_29518);
or UO_1832 (O_1832,N_28999,N_28496);
nand UO_1833 (O_1833,N_28777,N_29173);
nor UO_1834 (O_1834,N_29223,N_29484);
xnor UO_1835 (O_1835,N_29918,N_28542);
or UO_1836 (O_1836,N_28721,N_29099);
or UO_1837 (O_1837,N_29472,N_29558);
xnor UO_1838 (O_1838,N_29295,N_28461);
nor UO_1839 (O_1839,N_29067,N_28026);
nor UO_1840 (O_1840,N_28348,N_29510);
nor UO_1841 (O_1841,N_28664,N_29465);
or UO_1842 (O_1842,N_29828,N_28894);
xnor UO_1843 (O_1843,N_29600,N_28390);
nand UO_1844 (O_1844,N_28249,N_28979);
nor UO_1845 (O_1845,N_29358,N_28742);
or UO_1846 (O_1846,N_28970,N_28157);
nand UO_1847 (O_1847,N_29026,N_29812);
or UO_1848 (O_1848,N_29680,N_28821);
nand UO_1849 (O_1849,N_29280,N_28056);
or UO_1850 (O_1850,N_28413,N_29240);
nor UO_1851 (O_1851,N_28408,N_29755);
and UO_1852 (O_1852,N_29349,N_28501);
xnor UO_1853 (O_1853,N_28977,N_28559);
nand UO_1854 (O_1854,N_29013,N_29326);
nand UO_1855 (O_1855,N_28379,N_28629);
xor UO_1856 (O_1856,N_29034,N_29676);
xor UO_1857 (O_1857,N_29578,N_28448);
or UO_1858 (O_1858,N_29448,N_28775);
nor UO_1859 (O_1859,N_29404,N_29236);
and UO_1860 (O_1860,N_28692,N_29863);
or UO_1861 (O_1861,N_28553,N_29719);
nand UO_1862 (O_1862,N_28456,N_28977);
xnor UO_1863 (O_1863,N_28476,N_28607);
nor UO_1864 (O_1864,N_28116,N_29680);
nand UO_1865 (O_1865,N_28796,N_28043);
xor UO_1866 (O_1866,N_29229,N_28099);
nor UO_1867 (O_1867,N_28095,N_28744);
xor UO_1868 (O_1868,N_29650,N_28876);
nor UO_1869 (O_1869,N_29982,N_28733);
nand UO_1870 (O_1870,N_28389,N_28937);
nor UO_1871 (O_1871,N_28425,N_28066);
nand UO_1872 (O_1872,N_28248,N_29096);
or UO_1873 (O_1873,N_29836,N_28541);
and UO_1874 (O_1874,N_28662,N_29746);
nand UO_1875 (O_1875,N_29960,N_28404);
or UO_1876 (O_1876,N_29795,N_28416);
nor UO_1877 (O_1877,N_29095,N_28705);
and UO_1878 (O_1878,N_28920,N_28105);
or UO_1879 (O_1879,N_28873,N_29525);
nor UO_1880 (O_1880,N_28047,N_28738);
nor UO_1881 (O_1881,N_28864,N_29453);
xnor UO_1882 (O_1882,N_28665,N_29457);
nor UO_1883 (O_1883,N_28432,N_29484);
xnor UO_1884 (O_1884,N_29693,N_29504);
nor UO_1885 (O_1885,N_28488,N_28589);
nor UO_1886 (O_1886,N_28240,N_29179);
nor UO_1887 (O_1887,N_28918,N_28989);
xor UO_1888 (O_1888,N_28593,N_29326);
nor UO_1889 (O_1889,N_29914,N_29315);
and UO_1890 (O_1890,N_28841,N_28652);
or UO_1891 (O_1891,N_28439,N_28126);
xor UO_1892 (O_1892,N_28660,N_29183);
nor UO_1893 (O_1893,N_28668,N_29996);
or UO_1894 (O_1894,N_29946,N_28240);
and UO_1895 (O_1895,N_28711,N_29948);
nand UO_1896 (O_1896,N_29883,N_28001);
nor UO_1897 (O_1897,N_29460,N_29813);
xor UO_1898 (O_1898,N_29239,N_28222);
nand UO_1899 (O_1899,N_29032,N_28327);
xnor UO_1900 (O_1900,N_28288,N_28807);
or UO_1901 (O_1901,N_29045,N_29759);
nand UO_1902 (O_1902,N_28480,N_28770);
nand UO_1903 (O_1903,N_29636,N_28604);
and UO_1904 (O_1904,N_28128,N_28033);
nor UO_1905 (O_1905,N_28988,N_29445);
and UO_1906 (O_1906,N_29519,N_28589);
xnor UO_1907 (O_1907,N_29140,N_28825);
xnor UO_1908 (O_1908,N_28357,N_28555);
nand UO_1909 (O_1909,N_29700,N_29395);
nor UO_1910 (O_1910,N_28223,N_29038);
nor UO_1911 (O_1911,N_28426,N_28910);
and UO_1912 (O_1912,N_28221,N_29480);
xnor UO_1913 (O_1913,N_29856,N_29155);
and UO_1914 (O_1914,N_28486,N_29076);
and UO_1915 (O_1915,N_29838,N_28804);
and UO_1916 (O_1916,N_28561,N_28032);
xor UO_1917 (O_1917,N_28718,N_28525);
nor UO_1918 (O_1918,N_29845,N_28941);
or UO_1919 (O_1919,N_29649,N_28231);
nor UO_1920 (O_1920,N_29914,N_29050);
or UO_1921 (O_1921,N_28652,N_28302);
nor UO_1922 (O_1922,N_28659,N_28288);
nand UO_1923 (O_1923,N_29088,N_29087);
xnor UO_1924 (O_1924,N_29813,N_28756);
nand UO_1925 (O_1925,N_28604,N_29384);
and UO_1926 (O_1926,N_28146,N_29047);
nand UO_1927 (O_1927,N_29320,N_28998);
xnor UO_1928 (O_1928,N_28567,N_28131);
or UO_1929 (O_1929,N_28629,N_29274);
nor UO_1930 (O_1930,N_28121,N_28673);
or UO_1931 (O_1931,N_28054,N_29317);
xnor UO_1932 (O_1932,N_29912,N_28141);
xnor UO_1933 (O_1933,N_28922,N_28820);
or UO_1934 (O_1934,N_29211,N_28440);
xnor UO_1935 (O_1935,N_29414,N_28087);
and UO_1936 (O_1936,N_28588,N_28370);
nand UO_1937 (O_1937,N_29418,N_28735);
xnor UO_1938 (O_1938,N_29886,N_28126);
nand UO_1939 (O_1939,N_29687,N_29186);
and UO_1940 (O_1940,N_28818,N_28201);
and UO_1941 (O_1941,N_28483,N_29436);
xor UO_1942 (O_1942,N_29934,N_28162);
and UO_1943 (O_1943,N_28513,N_29940);
nand UO_1944 (O_1944,N_29057,N_28899);
nand UO_1945 (O_1945,N_29914,N_29276);
and UO_1946 (O_1946,N_28595,N_28225);
and UO_1947 (O_1947,N_28387,N_28185);
nor UO_1948 (O_1948,N_28556,N_28347);
or UO_1949 (O_1949,N_29778,N_28527);
nor UO_1950 (O_1950,N_29482,N_29982);
xor UO_1951 (O_1951,N_29252,N_28667);
nor UO_1952 (O_1952,N_28443,N_28459);
or UO_1953 (O_1953,N_28268,N_28481);
or UO_1954 (O_1954,N_29486,N_29216);
nand UO_1955 (O_1955,N_28546,N_28391);
nand UO_1956 (O_1956,N_28580,N_28995);
and UO_1957 (O_1957,N_29627,N_28392);
or UO_1958 (O_1958,N_29369,N_28268);
nor UO_1959 (O_1959,N_29413,N_28351);
and UO_1960 (O_1960,N_28174,N_29437);
or UO_1961 (O_1961,N_28991,N_29388);
nor UO_1962 (O_1962,N_29310,N_29220);
and UO_1963 (O_1963,N_29018,N_28441);
nor UO_1964 (O_1964,N_29856,N_28332);
or UO_1965 (O_1965,N_29819,N_28239);
nor UO_1966 (O_1966,N_28870,N_29014);
nand UO_1967 (O_1967,N_29682,N_28868);
and UO_1968 (O_1968,N_28505,N_29276);
or UO_1969 (O_1969,N_28251,N_28965);
nor UO_1970 (O_1970,N_29874,N_29845);
nor UO_1971 (O_1971,N_29997,N_29566);
nor UO_1972 (O_1972,N_29152,N_29427);
and UO_1973 (O_1973,N_28943,N_29850);
nand UO_1974 (O_1974,N_29017,N_29563);
or UO_1975 (O_1975,N_29552,N_28234);
and UO_1976 (O_1976,N_28791,N_29859);
nand UO_1977 (O_1977,N_28469,N_29390);
xnor UO_1978 (O_1978,N_28168,N_29826);
nor UO_1979 (O_1979,N_29665,N_29591);
xnor UO_1980 (O_1980,N_28226,N_29571);
xnor UO_1981 (O_1981,N_29182,N_28029);
or UO_1982 (O_1982,N_28140,N_29668);
and UO_1983 (O_1983,N_28735,N_29940);
nor UO_1984 (O_1984,N_29886,N_28232);
xor UO_1985 (O_1985,N_29079,N_28924);
xnor UO_1986 (O_1986,N_28603,N_28254);
xor UO_1987 (O_1987,N_29827,N_29017);
or UO_1988 (O_1988,N_29791,N_28155);
nand UO_1989 (O_1989,N_29686,N_29399);
nor UO_1990 (O_1990,N_28027,N_29172);
or UO_1991 (O_1991,N_28272,N_29429);
nor UO_1992 (O_1992,N_28086,N_28860);
and UO_1993 (O_1993,N_29457,N_29985);
nor UO_1994 (O_1994,N_28010,N_29733);
xnor UO_1995 (O_1995,N_28452,N_29997);
xor UO_1996 (O_1996,N_28055,N_28940);
and UO_1997 (O_1997,N_29826,N_29641);
nand UO_1998 (O_1998,N_29956,N_28267);
nand UO_1999 (O_1999,N_29109,N_29818);
nor UO_2000 (O_2000,N_29725,N_29411);
nand UO_2001 (O_2001,N_29676,N_29545);
nand UO_2002 (O_2002,N_29351,N_28781);
nand UO_2003 (O_2003,N_29972,N_28057);
nor UO_2004 (O_2004,N_29678,N_28122);
xnor UO_2005 (O_2005,N_28953,N_29041);
and UO_2006 (O_2006,N_28760,N_28725);
nand UO_2007 (O_2007,N_29392,N_29653);
and UO_2008 (O_2008,N_29878,N_28225);
nor UO_2009 (O_2009,N_28974,N_28917);
or UO_2010 (O_2010,N_29426,N_29311);
or UO_2011 (O_2011,N_28126,N_29110);
nor UO_2012 (O_2012,N_29522,N_28558);
and UO_2013 (O_2013,N_29480,N_28917);
and UO_2014 (O_2014,N_29658,N_29871);
xnor UO_2015 (O_2015,N_28668,N_28404);
nor UO_2016 (O_2016,N_28749,N_28908);
and UO_2017 (O_2017,N_29247,N_28768);
xor UO_2018 (O_2018,N_29674,N_28100);
nand UO_2019 (O_2019,N_28303,N_28416);
and UO_2020 (O_2020,N_29313,N_28143);
and UO_2021 (O_2021,N_29531,N_28360);
nor UO_2022 (O_2022,N_29735,N_29221);
and UO_2023 (O_2023,N_28998,N_29789);
xor UO_2024 (O_2024,N_29262,N_28907);
nand UO_2025 (O_2025,N_29286,N_28176);
or UO_2026 (O_2026,N_28692,N_29714);
nand UO_2027 (O_2027,N_29291,N_29836);
and UO_2028 (O_2028,N_28337,N_28331);
nand UO_2029 (O_2029,N_29670,N_28383);
nor UO_2030 (O_2030,N_28017,N_28906);
and UO_2031 (O_2031,N_29812,N_28935);
xnor UO_2032 (O_2032,N_28133,N_28776);
nor UO_2033 (O_2033,N_29375,N_28041);
or UO_2034 (O_2034,N_29141,N_29631);
xnor UO_2035 (O_2035,N_29971,N_28045);
xor UO_2036 (O_2036,N_29065,N_29474);
nor UO_2037 (O_2037,N_29198,N_28946);
nor UO_2038 (O_2038,N_29966,N_29778);
or UO_2039 (O_2039,N_29999,N_29059);
nand UO_2040 (O_2040,N_28814,N_29950);
xnor UO_2041 (O_2041,N_28418,N_28013);
nor UO_2042 (O_2042,N_29276,N_28151);
and UO_2043 (O_2043,N_29723,N_29462);
and UO_2044 (O_2044,N_28704,N_29703);
xnor UO_2045 (O_2045,N_28034,N_28062);
and UO_2046 (O_2046,N_28330,N_29566);
or UO_2047 (O_2047,N_28280,N_28082);
nand UO_2048 (O_2048,N_28685,N_28284);
nand UO_2049 (O_2049,N_28612,N_29992);
or UO_2050 (O_2050,N_28387,N_29669);
or UO_2051 (O_2051,N_29819,N_28487);
nor UO_2052 (O_2052,N_29421,N_28878);
and UO_2053 (O_2053,N_28696,N_29210);
and UO_2054 (O_2054,N_29285,N_29733);
and UO_2055 (O_2055,N_29381,N_29215);
xor UO_2056 (O_2056,N_28085,N_29774);
and UO_2057 (O_2057,N_28831,N_28119);
nand UO_2058 (O_2058,N_29561,N_28773);
or UO_2059 (O_2059,N_28910,N_29168);
or UO_2060 (O_2060,N_29400,N_28838);
nand UO_2061 (O_2061,N_29355,N_29421);
or UO_2062 (O_2062,N_29844,N_29063);
or UO_2063 (O_2063,N_28197,N_29847);
and UO_2064 (O_2064,N_29768,N_28227);
or UO_2065 (O_2065,N_29408,N_29195);
nor UO_2066 (O_2066,N_29855,N_29419);
or UO_2067 (O_2067,N_28705,N_29532);
or UO_2068 (O_2068,N_28124,N_29621);
xnor UO_2069 (O_2069,N_29631,N_29707);
nor UO_2070 (O_2070,N_29582,N_28995);
and UO_2071 (O_2071,N_29022,N_28427);
and UO_2072 (O_2072,N_29426,N_29589);
and UO_2073 (O_2073,N_29716,N_28890);
nand UO_2074 (O_2074,N_28849,N_28766);
or UO_2075 (O_2075,N_29146,N_29987);
nand UO_2076 (O_2076,N_28454,N_28277);
xnor UO_2077 (O_2077,N_29484,N_28180);
or UO_2078 (O_2078,N_28811,N_29525);
nor UO_2079 (O_2079,N_28767,N_28738);
xnor UO_2080 (O_2080,N_29358,N_29101);
nor UO_2081 (O_2081,N_28085,N_28936);
nand UO_2082 (O_2082,N_28919,N_28520);
xnor UO_2083 (O_2083,N_29835,N_28986);
or UO_2084 (O_2084,N_29603,N_29610);
nor UO_2085 (O_2085,N_29148,N_28245);
nand UO_2086 (O_2086,N_28426,N_29190);
and UO_2087 (O_2087,N_29804,N_28279);
or UO_2088 (O_2088,N_29196,N_28108);
or UO_2089 (O_2089,N_29407,N_29426);
or UO_2090 (O_2090,N_28748,N_29774);
xnor UO_2091 (O_2091,N_28628,N_28327);
or UO_2092 (O_2092,N_29227,N_29595);
or UO_2093 (O_2093,N_29107,N_29269);
nand UO_2094 (O_2094,N_28208,N_28878);
nand UO_2095 (O_2095,N_28282,N_28200);
nor UO_2096 (O_2096,N_29118,N_29677);
and UO_2097 (O_2097,N_29203,N_28036);
nand UO_2098 (O_2098,N_28819,N_29538);
nand UO_2099 (O_2099,N_28387,N_29883);
or UO_2100 (O_2100,N_29608,N_28038);
xnor UO_2101 (O_2101,N_28574,N_29851);
nand UO_2102 (O_2102,N_28979,N_28359);
nor UO_2103 (O_2103,N_28172,N_29838);
nor UO_2104 (O_2104,N_28404,N_28734);
nor UO_2105 (O_2105,N_28299,N_29557);
nand UO_2106 (O_2106,N_29379,N_29498);
xor UO_2107 (O_2107,N_29805,N_28847);
or UO_2108 (O_2108,N_28625,N_28602);
nand UO_2109 (O_2109,N_29108,N_29133);
and UO_2110 (O_2110,N_28830,N_28417);
nor UO_2111 (O_2111,N_29040,N_28558);
or UO_2112 (O_2112,N_29117,N_28268);
nand UO_2113 (O_2113,N_29851,N_29856);
nor UO_2114 (O_2114,N_29790,N_29152);
xnor UO_2115 (O_2115,N_28824,N_28948);
xnor UO_2116 (O_2116,N_29695,N_28540);
or UO_2117 (O_2117,N_28917,N_29793);
and UO_2118 (O_2118,N_29144,N_29647);
nand UO_2119 (O_2119,N_28480,N_28963);
or UO_2120 (O_2120,N_29693,N_29842);
or UO_2121 (O_2121,N_28851,N_28743);
nand UO_2122 (O_2122,N_29273,N_28682);
xor UO_2123 (O_2123,N_29104,N_28194);
nor UO_2124 (O_2124,N_29799,N_28938);
xnor UO_2125 (O_2125,N_28969,N_28273);
and UO_2126 (O_2126,N_29700,N_29219);
nand UO_2127 (O_2127,N_29770,N_28861);
and UO_2128 (O_2128,N_28886,N_28555);
nand UO_2129 (O_2129,N_29802,N_29921);
nor UO_2130 (O_2130,N_29036,N_28385);
nand UO_2131 (O_2131,N_29083,N_28596);
nor UO_2132 (O_2132,N_29207,N_28084);
nand UO_2133 (O_2133,N_29869,N_29844);
or UO_2134 (O_2134,N_28572,N_28319);
nand UO_2135 (O_2135,N_29703,N_28365);
nor UO_2136 (O_2136,N_28333,N_28160);
nor UO_2137 (O_2137,N_29746,N_28193);
or UO_2138 (O_2138,N_29638,N_29338);
or UO_2139 (O_2139,N_29890,N_29545);
xnor UO_2140 (O_2140,N_29335,N_28988);
or UO_2141 (O_2141,N_28350,N_29416);
and UO_2142 (O_2142,N_28959,N_28326);
and UO_2143 (O_2143,N_28731,N_29400);
and UO_2144 (O_2144,N_28295,N_28000);
nor UO_2145 (O_2145,N_28533,N_29809);
and UO_2146 (O_2146,N_29146,N_28937);
xnor UO_2147 (O_2147,N_29282,N_29653);
nand UO_2148 (O_2148,N_29026,N_29279);
and UO_2149 (O_2149,N_28037,N_28499);
xor UO_2150 (O_2150,N_28321,N_29547);
nand UO_2151 (O_2151,N_29068,N_29492);
xor UO_2152 (O_2152,N_28266,N_29960);
nor UO_2153 (O_2153,N_28297,N_28671);
xnor UO_2154 (O_2154,N_28641,N_28229);
and UO_2155 (O_2155,N_28437,N_29874);
xor UO_2156 (O_2156,N_28282,N_29514);
or UO_2157 (O_2157,N_28608,N_28184);
nor UO_2158 (O_2158,N_29404,N_29635);
nor UO_2159 (O_2159,N_29444,N_29119);
nor UO_2160 (O_2160,N_28879,N_28875);
or UO_2161 (O_2161,N_28650,N_29715);
nand UO_2162 (O_2162,N_28853,N_29202);
or UO_2163 (O_2163,N_28780,N_28246);
and UO_2164 (O_2164,N_28250,N_28975);
xnor UO_2165 (O_2165,N_28977,N_28889);
nor UO_2166 (O_2166,N_28378,N_28978);
nor UO_2167 (O_2167,N_29802,N_28754);
and UO_2168 (O_2168,N_29827,N_28707);
nor UO_2169 (O_2169,N_28016,N_29346);
nor UO_2170 (O_2170,N_29719,N_29960);
nand UO_2171 (O_2171,N_29835,N_28069);
and UO_2172 (O_2172,N_29083,N_28531);
and UO_2173 (O_2173,N_29200,N_29699);
and UO_2174 (O_2174,N_29544,N_28482);
xnor UO_2175 (O_2175,N_28368,N_28173);
nor UO_2176 (O_2176,N_28926,N_29546);
nand UO_2177 (O_2177,N_29385,N_29013);
xnor UO_2178 (O_2178,N_29851,N_28661);
and UO_2179 (O_2179,N_29623,N_28576);
or UO_2180 (O_2180,N_29858,N_28568);
xnor UO_2181 (O_2181,N_28244,N_28739);
nand UO_2182 (O_2182,N_28509,N_29812);
or UO_2183 (O_2183,N_28739,N_28335);
xor UO_2184 (O_2184,N_28490,N_29169);
nand UO_2185 (O_2185,N_29732,N_29411);
and UO_2186 (O_2186,N_29269,N_29005);
nor UO_2187 (O_2187,N_29637,N_28288);
nand UO_2188 (O_2188,N_28061,N_29695);
and UO_2189 (O_2189,N_29188,N_28199);
and UO_2190 (O_2190,N_28266,N_29946);
or UO_2191 (O_2191,N_29306,N_28482);
nor UO_2192 (O_2192,N_29205,N_28708);
nand UO_2193 (O_2193,N_28641,N_28193);
nand UO_2194 (O_2194,N_28190,N_28666);
nand UO_2195 (O_2195,N_28111,N_29112);
xor UO_2196 (O_2196,N_29625,N_28148);
xor UO_2197 (O_2197,N_28409,N_28293);
nand UO_2198 (O_2198,N_29249,N_29906);
and UO_2199 (O_2199,N_28317,N_28954);
nand UO_2200 (O_2200,N_29877,N_29826);
xnor UO_2201 (O_2201,N_28339,N_29654);
nor UO_2202 (O_2202,N_29234,N_29500);
and UO_2203 (O_2203,N_28353,N_29431);
nand UO_2204 (O_2204,N_29345,N_29692);
nand UO_2205 (O_2205,N_29939,N_29316);
nor UO_2206 (O_2206,N_29353,N_29056);
or UO_2207 (O_2207,N_29561,N_29564);
and UO_2208 (O_2208,N_29553,N_29910);
xnor UO_2209 (O_2209,N_28617,N_28196);
or UO_2210 (O_2210,N_28962,N_29012);
or UO_2211 (O_2211,N_28055,N_28365);
or UO_2212 (O_2212,N_28582,N_29532);
or UO_2213 (O_2213,N_28958,N_29663);
xnor UO_2214 (O_2214,N_28313,N_28445);
nand UO_2215 (O_2215,N_28002,N_28488);
xnor UO_2216 (O_2216,N_28853,N_29939);
and UO_2217 (O_2217,N_29214,N_28161);
xor UO_2218 (O_2218,N_29131,N_28604);
nor UO_2219 (O_2219,N_28171,N_29627);
xor UO_2220 (O_2220,N_29976,N_29583);
xor UO_2221 (O_2221,N_28975,N_28003);
nor UO_2222 (O_2222,N_28014,N_29639);
nand UO_2223 (O_2223,N_29969,N_29731);
or UO_2224 (O_2224,N_28136,N_28629);
xor UO_2225 (O_2225,N_28857,N_28375);
xnor UO_2226 (O_2226,N_28770,N_29128);
xnor UO_2227 (O_2227,N_29760,N_29599);
or UO_2228 (O_2228,N_28668,N_28366);
or UO_2229 (O_2229,N_28473,N_28242);
and UO_2230 (O_2230,N_29711,N_29396);
xnor UO_2231 (O_2231,N_28729,N_29031);
or UO_2232 (O_2232,N_29240,N_28518);
and UO_2233 (O_2233,N_28739,N_29029);
nor UO_2234 (O_2234,N_29651,N_28781);
nand UO_2235 (O_2235,N_29087,N_28314);
or UO_2236 (O_2236,N_29517,N_29138);
and UO_2237 (O_2237,N_29302,N_28211);
or UO_2238 (O_2238,N_28960,N_29846);
nand UO_2239 (O_2239,N_28578,N_28328);
nand UO_2240 (O_2240,N_28547,N_28887);
xnor UO_2241 (O_2241,N_28219,N_29096);
or UO_2242 (O_2242,N_29403,N_29124);
and UO_2243 (O_2243,N_29546,N_29245);
or UO_2244 (O_2244,N_29420,N_29999);
xor UO_2245 (O_2245,N_28215,N_28907);
nand UO_2246 (O_2246,N_29980,N_28711);
nor UO_2247 (O_2247,N_28305,N_29049);
nor UO_2248 (O_2248,N_29199,N_28432);
and UO_2249 (O_2249,N_28911,N_28292);
and UO_2250 (O_2250,N_28924,N_28475);
nand UO_2251 (O_2251,N_28271,N_28175);
nor UO_2252 (O_2252,N_28395,N_29055);
and UO_2253 (O_2253,N_29348,N_28789);
or UO_2254 (O_2254,N_28408,N_29732);
or UO_2255 (O_2255,N_29148,N_28402);
xor UO_2256 (O_2256,N_29940,N_29571);
xor UO_2257 (O_2257,N_28844,N_29676);
nor UO_2258 (O_2258,N_28510,N_28306);
xnor UO_2259 (O_2259,N_28097,N_28919);
xor UO_2260 (O_2260,N_29204,N_29882);
nand UO_2261 (O_2261,N_28593,N_28568);
or UO_2262 (O_2262,N_28194,N_29765);
or UO_2263 (O_2263,N_28909,N_28109);
nand UO_2264 (O_2264,N_29881,N_28041);
nand UO_2265 (O_2265,N_28559,N_28240);
and UO_2266 (O_2266,N_28166,N_28231);
xnor UO_2267 (O_2267,N_29615,N_29596);
xnor UO_2268 (O_2268,N_29586,N_28659);
or UO_2269 (O_2269,N_28790,N_29849);
nor UO_2270 (O_2270,N_28761,N_29486);
nor UO_2271 (O_2271,N_28668,N_28802);
and UO_2272 (O_2272,N_28118,N_29800);
xor UO_2273 (O_2273,N_29270,N_29450);
or UO_2274 (O_2274,N_28933,N_28213);
and UO_2275 (O_2275,N_29763,N_28064);
nor UO_2276 (O_2276,N_28479,N_29258);
and UO_2277 (O_2277,N_29860,N_29902);
nor UO_2278 (O_2278,N_29918,N_29731);
nor UO_2279 (O_2279,N_28920,N_29911);
xnor UO_2280 (O_2280,N_29361,N_29481);
and UO_2281 (O_2281,N_28197,N_28475);
and UO_2282 (O_2282,N_29528,N_29330);
nor UO_2283 (O_2283,N_28163,N_28768);
or UO_2284 (O_2284,N_29216,N_29570);
xor UO_2285 (O_2285,N_29284,N_28287);
nor UO_2286 (O_2286,N_29542,N_28731);
nand UO_2287 (O_2287,N_29692,N_29107);
nor UO_2288 (O_2288,N_28801,N_28038);
xnor UO_2289 (O_2289,N_28403,N_29149);
nand UO_2290 (O_2290,N_29412,N_29067);
or UO_2291 (O_2291,N_28511,N_28908);
nor UO_2292 (O_2292,N_28770,N_28574);
xor UO_2293 (O_2293,N_29977,N_29072);
and UO_2294 (O_2294,N_29343,N_28786);
xnor UO_2295 (O_2295,N_28604,N_29050);
and UO_2296 (O_2296,N_29874,N_28715);
or UO_2297 (O_2297,N_28801,N_29931);
xnor UO_2298 (O_2298,N_28674,N_29440);
nor UO_2299 (O_2299,N_28431,N_28885);
nor UO_2300 (O_2300,N_29080,N_29386);
nor UO_2301 (O_2301,N_28534,N_29236);
nand UO_2302 (O_2302,N_29290,N_28414);
or UO_2303 (O_2303,N_28530,N_28240);
nor UO_2304 (O_2304,N_29469,N_28673);
nor UO_2305 (O_2305,N_28400,N_29300);
and UO_2306 (O_2306,N_29366,N_29977);
and UO_2307 (O_2307,N_29863,N_29067);
nor UO_2308 (O_2308,N_29434,N_29312);
nand UO_2309 (O_2309,N_28286,N_28776);
nor UO_2310 (O_2310,N_28409,N_28374);
nor UO_2311 (O_2311,N_28582,N_28535);
nand UO_2312 (O_2312,N_28366,N_28663);
or UO_2313 (O_2313,N_29006,N_29365);
nor UO_2314 (O_2314,N_28619,N_28947);
nor UO_2315 (O_2315,N_29457,N_29140);
nand UO_2316 (O_2316,N_29463,N_28729);
xor UO_2317 (O_2317,N_28732,N_29708);
or UO_2318 (O_2318,N_28373,N_28786);
nand UO_2319 (O_2319,N_29832,N_28736);
nor UO_2320 (O_2320,N_29224,N_29011);
nor UO_2321 (O_2321,N_29689,N_29854);
nor UO_2322 (O_2322,N_29413,N_28129);
or UO_2323 (O_2323,N_29954,N_29283);
or UO_2324 (O_2324,N_28266,N_28760);
nand UO_2325 (O_2325,N_28439,N_28188);
and UO_2326 (O_2326,N_29684,N_28983);
nand UO_2327 (O_2327,N_28823,N_29244);
xnor UO_2328 (O_2328,N_28867,N_28145);
nor UO_2329 (O_2329,N_28573,N_28319);
nand UO_2330 (O_2330,N_29389,N_28005);
or UO_2331 (O_2331,N_28613,N_28130);
nand UO_2332 (O_2332,N_29255,N_28816);
or UO_2333 (O_2333,N_29801,N_29682);
or UO_2334 (O_2334,N_28017,N_28030);
or UO_2335 (O_2335,N_29322,N_28826);
xor UO_2336 (O_2336,N_28374,N_29168);
xor UO_2337 (O_2337,N_28508,N_28489);
or UO_2338 (O_2338,N_29416,N_29900);
xor UO_2339 (O_2339,N_28398,N_29142);
or UO_2340 (O_2340,N_29520,N_29196);
nor UO_2341 (O_2341,N_29859,N_28486);
or UO_2342 (O_2342,N_28971,N_29567);
xnor UO_2343 (O_2343,N_29635,N_29419);
or UO_2344 (O_2344,N_29298,N_28716);
nor UO_2345 (O_2345,N_29481,N_28883);
nor UO_2346 (O_2346,N_28826,N_28652);
nand UO_2347 (O_2347,N_28613,N_29476);
xor UO_2348 (O_2348,N_29481,N_29896);
or UO_2349 (O_2349,N_28026,N_28930);
xnor UO_2350 (O_2350,N_28933,N_29585);
and UO_2351 (O_2351,N_28208,N_28974);
and UO_2352 (O_2352,N_29464,N_29597);
xnor UO_2353 (O_2353,N_28396,N_29436);
nor UO_2354 (O_2354,N_28987,N_29348);
nor UO_2355 (O_2355,N_29018,N_28957);
xnor UO_2356 (O_2356,N_28612,N_28138);
and UO_2357 (O_2357,N_29450,N_28877);
or UO_2358 (O_2358,N_28468,N_28979);
nand UO_2359 (O_2359,N_28717,N_28410);
or UO_2360 (O_2360,N_29473,N_28529);
xnor UO_2361 (O_2361,N_28000,N_28802);
xnor UO_2362 (O_2362,N_29425,N_28408);
or UO_2363 (O_2363,N_28283,N_28544);
and UO_2364 (O_2364,N_29950,N_28019);
nor UO_2365 (O_2365,N_28937,N_28490);
or UO_2366 (O_2366,N_29429,N_28998);
xor UO_2367 (O_2367,N_29347,N_28874);
nand UO_2368 (O_2368,N_29765,N_28026);
xor UO_2369 (O_2369,N_29208,N_29456);
nor UO_2370 (O_2370,N_28789,N_28159);
nor UO_2371 (O_2371,N_28388,N_28540);
nor UO_2372 (O_2372,N_28358,N_29011);
or UO_2373 (O_2373,N_28728,N_29741);
or UO_2374 (O_2374,N_28562,N_29154);
and UO_2375 (O_2375,N_29735,N_29986);
and UO_2376 (O_2376,N_28270,N_28078);
nor UO_2377 (O_2377,N_28246,N_28555);
or UO_2378 (O_2378,N_28563,N_28609);
xnor UO_2379 (O_2379,N_29332,N_28267);
and UO_2380 (O_2380,N_29890,N_29013);
xor UO_2381 (O_2381,N_28831,N_28082);
and UO_2382 (O_2382,N_29438,N_29641);
nand UO_2383 (O_2383,N_28056,N_29595);
and UO_2384 (O_2384,N_29168,N_29683);
nor UO_2385 (O_2385,N_29868,N_29965);
xnor UO_2386 (O_2386,N_28538,N_29592);
xor UO_2387 (O_2387,N_28295,N_29315);
or UO_2388 (O_2388,N_28890,N_29440);
and UO_2389 (O_2389,N_28005,N_28378);
nor UO_2390 (O_2390,N_28929,N_29345);
nand UO_2391 (O_2391,N_29610,N_29237);
xor UO_2392 (O_2392,N_28492,N_28092);
nand UO_2393 (O_2393,N_29513,N_28560);
xnor UO_2394 (O_2394,N_28574,N_28719);
and UO_2395 (O_2395,N_28645,N_28047);
nor UO_2396 (O_2396,N_29904,N_29854);
nand UO_2397 (O_2397,N_29931,N_29326);
nor UO_2398 (O_2398,N_28312,N_28044);
or UO_2399 (O_2399,N_28927,N_29739);
and UO_2400 (O_2400,N_29076,N_29595);
and UO_2401 (O_2401,N_29882,N_29632);
xor UO_2402 (O_2402,N_29427,N_29092);
xnor UO_2403 (O_2403,N_29224,N_28417);
nand UO_2404 (O_2404,N_29746,N_29398);
or UO_2405 (O_2405,N_28244,N_28143);
and UO_2406 (O_2406,N_29125,N_28844);
nor UO_2407 (O_2407,N_29241,N_29663);
nor UO_2408 (O_2408,N_29874,N_29380);
or UO_2409 (O_2409,N_28653,N_28434);
nor UO_2410 (O_2410,N_28653,N_29240);
or UO_2411 (O_2411,N_29171,N_28177);
and UO_2412 (O_2412,N_29182,N_29001);
or UO_2413 (O_2413,N_29330,N_28561);
nand UO_2414 (O_2414,N_29036,N_29195);
or UO_2415 (O_2415,N_28127,N_28202);
nor UO_2416 (O_2416,N_28433,N_28690);
and UO_2417 (O_2417,N_28401,N_29488);
nor UO_2418 (O_2418,N_28848,N_29816);
nand UO_2419 (O_2419,N_28023,N_29576);
nor UO_2420 (O_2420,N_29483,N_29115);
nor UO_2421 (O_2421,N_29845,N_29034);
xor UO_2422 (O_2422,N_29810,N_29987);
and UO_2423 (O_2423,N_28204,N_29927);
or UO_2424 (O_2424,N_29965,N_29097);
nor UO_2425 (O_2425,N_28301,N_29449);
and UO_2426 (O_2426,N_28360,N_29705);
nor UO_2427 (O_2427,N_28649,N_28768);
nand UO_2428 (O_2428,N_29568,N_29931);
nor UO_2429 (O_2429,N_28832,N_28834);
and UO_2430 (O_2430,N_28803,N_28959);
or UO_2431 (O_2431,N_28599,N_28028);
or UO_2432 (O_2432,N_28054,N_29587);
nand UO_2433 (O_2433,N_29062,N_29471);
nand UO_2434 (O_2434,N_28730,N_28560);
and UO_2435 (O_2435,N_29648,N_29195);
nor UO_2436 (O_2436,N_29818,N_28117);
and UO_2437 (O_2437,N_28104,N_29566);
nand UO_2438 (O_2438,N_29248,N_28513);
and UO_2439 (O_2439,N_28337,N_28470);
and UO_2440 (O_2440,N_29827,N_28113);
or UO_2441 (O_2441,N_29489,N_29616);
or UO_2442 (O_2442,N_28037,N_29301);
xnor UO_2443 (O_2443,N_28479,N_28747);
and UO_2444 (O_2444,N_28407,N_28411);
nor UO_2445 (O_2445,N_28369,N_29388);
and UO_2446 (O_2446,N_29102,N_29441);
or UO_2447 (O_2447,N_29196,N_28522);
and UO_2448 (O_2448,N_28535,N_29855);
or UO_2449 (O_2449,N_29350,N_28104);
nor UO_2450 (O_2450,N_29899,N_29058);
or UO_2451 (O_2451,N_29752,N_29176);
xnor UO_2452 (O_2452,N_28363,N_29024);
nor UO_2453 (O_2453,N_29485,N_29153);
and UO_2454 (O_2454,N_28581,N_28112);
and UO_2455 (O_2455,N_28937,N_29711);
xnor UO_2456 (O_2456,N_29648,N_29227);
or UO_2457 (O_2457,N_28892,N_29814);
and UO_2458 (O_2458,N_28919,N_29383);
and UO_2459 (O_2459,N_28676,N_28985);
nor UO_2460 (O_2460,N_28177,N_29913);
nand UO_2461 (O_2461,N_29547,N_28276);
nand UO_2462 (O_2462,N_29879,N_29862);
nor UO_2463 (O_2463,N_29460,N_28577);
and UO_2464 (O_2464,N_28142,N_28193);
and UO_2465 (O_2465,N_28085,N_29789);
nor UO_2466 (O_2466,N_28578,N_29662);
nand UO_2467 (O_2467,N_29034,N_29747);
or UO_2468 (O_2468,N_28320,N_28939);
xor UO_2469 (O_2469,N_28965,N_29541);
nand UO_2470 (O_2470,N_29087,N_29147);
xor UO_2471 (O_2471,N_28774,N_29239);
nand UO_2472 (O_2472,N_28534,N_28439);
and UO_2473 (O_2473,N_28741,N_29249);
and UO_2474 (O_2474,N_28206,N_29692);
and UO_2475 (O_2475,N_28887,N_29180);
nor UO_2476 (O_2476,N_28692,N_28770);
xor UO_2477 (O_2477,N_28312,N_28419);
or UO_2478 (O_2478,N_28417,N_28857);
nand UO_2479 (O_2479,N_28497,N_29416);
and UO_2480 (O_2480,N_28233,N_28017);
and UO_2481 (O_2481,N_28124,N_28596);
nand UO_2482 (O_2482,N_29412,N_28668);
nand UO_2483 (O_2483,N_28097,N_28339);
nor UO_2484 (O_2484,N_28311,N_29566);
nor UO_2485 (O_2485,N_28404,N_28407);
xnor UO_2486 (O_2486,N_29372,N_29108);
nand UO_2487 (O_2487,N_28854,N_29660);
and UO_2488 (O_2488,N_28925,N_28185);
nor UO_2489 (O_2489,N_28288,N_29774);
nor UO_2490 (O_2490,N_29854,N_28845);
xnor UO_2491 (O_2491,N_29334,N_28313);
or UO_2492 (O_2492,N_29988,N_28152);
nand UO_2493 (O_2493,N_28470,N_29488);
xnor UO_2494 (O_2494,N_29714,N_28334);
xnor UO_2495 (O_2495,N_29455,N_29814);
nand UO_2496 (O_2496,N_28088,N_28760);
nor UO_2497 (O_2497,N_28060,N_29816);
xnor UO_2498 (O_2498,N_28096,N_29746);
and UO_2499 (O_2499,N_28978,N_29939);
xor UO_2500 (O_2500,N_28111,N_28258);
xnor UO_2501 (O_2501,N_28768,N_28582);
or UO_2502 (O_2502,N_29750,N_29558);
nand UO_2503 (O_2503,N_29108,N_29546);
nor UO_2504 (O_2504,N_29853,N_29019);
nor UO_2505 (O_2505,N_28918,N_28953);
and UO_2506 (O_2506,N_29977,N_28797);
or UO_2507 (O_2507,N_28397,N_28665);
nor UO_2508 (O_2508,N_28967,N_28356);
or UO_2509 (O_2509,N_28727,N_28005);
nor UO_2510 (O_2510,N_28287,N_29431);
nand UO_2511 (O_2511,N_28248,N_29929);
and UO_2512 (O_2512,N_28970,N_28253);
or UO_2513 (O_2513,N_28466,N_29127);
xor UO_2514 (O_2514,N_28626,N_29819);
nand UO_2515 (O_2515,N_28339,N_28807);
xor UO_2516 (O_2516,N_28626,N_29501);
and UO_2517 (O_2517,N_29387,N_28163);
nor UO_2518 (O_2518,N_29437,N_28407);
or UO_2519 (O_2519,N_29779,N_28699);
nand UO_2520 (O_2520,N_28799,N_28184);
xnor UO_2521 (O_2521,N_28327,N_28966);
xnor UO_2522 (O_2522,N_29185,N_28806);
nor UO_2523 (O_2523,N_28549,N_29557);
and UO_2524 (O_2524,N_29533,N_28747);
or UO_2525 (O_2525,N_28562,N_28774);
xnor UO_2526 (O_2526,N_29073,N_29338);
nand UO_2527 (O_2527,N_29889,N_29614);
nor UO_2528 (O_2528,N_28305,N_28701);
nor UO_2529 (O_2529,N_28665,N_28277);
nor UO_2530 (O_2530,N_28809,N_29399);
nor UO_2531 (O_2531,N_29591,N_28184);
nand UO_2532 (O_2532,N_28601,N_29545);
and UO_2533 (O_2533,N_28496,N_28217);
or UO_2534 (O_2534,N_28690,N_29913);
or UO_2535 (O_2535,N_29299,N_29767);
nand UO_2536 (O_2536,N_28295,N_28968);
nand UO_2537 (O_2537,N_28730,N_29503);
or UO_2538 (O_2538,N_28077,N_29295);
xor UO_2539 (O_2539,N_28571,N_29276);
and UO_2540 (O_2540,N_28613,N_29267);
xnor UO_2541 (O_2541,N_28065,N_28428);
nor UO_2542 (O_2542,N_28567,N_28524);
nor UO_2543 (O_2543,N_28075,N_29509);
and UO_2544 (O_2544,N_29965,N_29465);
xnor UO_2545 (O_2545,N_29256,N_28352);
and UO_2546 (O_2546,N_28091,N_29097);
nand UO_2547 (O_2547,N_28066,N_29861);
nor UO_2548 (O_2548,N_28680,N_28487);
or UO_2549 (O_2549,N_28317,N_29185);
or UO_2550 (O_2550,N_28507,N_28667);
nor UO_2551 (O_2551,N_28922,N_28445);
xnor UO_2552 (O_2552,N_28799,N_28256);
nand UO_2553 (O_2553,N_29331,N_29447);
nor UO_2554 (O_2554,N_29335,N_29517);
nor UO_2555 (O_2555,N_28058,N_28103);
xor UO_2556 (O_2556,N_28571,N_28494);
or UO_2557 (O_2557,N_29027,N_28753);
xor UO_2558 (O_2558,N_28241,N_29162);
nor UO_2559 (O_2559,N_29568,N_28626);
xor UO_2560 (O_2560,N_28285,N_28071);
xnor UO_2561 (O_2561,N_29787,N_29842);
nor UO_2562 (O_2562,N_28588,N_29639);
xor UO_2563 (O_2563,N_28176,N_28622);
xor UO_2564 (O_2564,N_28642,N_28452);
xor UO_2565 (O_2565,N_28068,N_29738);
nor UO_2566 (O_2566,N_28320,N_28192);
or UO_2567 (O_2567,N_28409,N_28729);
xnor UO_2568 (O_2568,N_29578,N_29069);
nor UO_2569 (O_2569,N_29215,N_28928);
nor UO_2570 (O_2570,N_28335,N_29162);
nand UO_2571 (O_2571,N_29913,N_28323);
or UO_2572 (O_2572,N_28455,N_28057);
or UO_2573 (O_2573,N_28718,N_28166);
nand UO_2574 (O_2574,N_29374,N_28889);
nor UO_2575 (O_2575,N_29805,N_29110);
nand UO_2576 (O_2576,N_28923,N_28523);
and UO_2577 (O_2577,N_29683,N_28133);
nor UO_2578 (O_2578,N_28512,N_28242);
xnor UO_2579 (O_2579,N_28404,N_28077);
nand UO_2580 (O_2580,N_29271,N_28450);
xor UO_2581 (O_2581,N_29858,N_29063);
or UO_2582 (O_2582,N_28500,N_29578);
or UO_2583 (O_2583,N_29363,N_28966);
xor UO_2584 (O_2584,N_28560,N_29768);
nand UO_2585 (O_2585,N_29499,N_29358);
nor UO_2586 (O_2586,N_29672,N_28291);
nor UO_2587 (O_2587,N_28487,N_29424);
and UO_2588 (O_2588,N_29873,N_28014);
nand UO_2589 (O_2589,N_29788,N_29135);
nand UO_2590 (O_2590,N_29599,N_29189);
nor UO_2591 (O_2591,N_29119,N_29167);
xnor UO_2592 (O_2592,N_29362,N_28732);
and UO_2593 (O_2593,N_28021,N_29811);
xor UO_2594 (O_2594,N_29428,N_29387);
nor UO_2595 (O_2595,N_28285,N_28543);
nor UO_2596 (O_2596,N_29826,N_28550);
and UO_2597 (O_2597,N_28325,N_28122);
nand UO_2598 (O_2598,N_29029,N_28318);
nor UO_2599 (O_2599,N_28168,N_28878);
and UO_2600 (O_2600,N_29978,N_28651);
nand UO_2601 (O_2601,N_28762,N_28658);
and UO_2602 (O_2602,N_29112,N_28628);
nor UO_2603 (O_2603,N_29596,N_28040);
and UO_2604 (O_2604,N_29751,N_29616);
or UO_2605 (O_2605,N_28871,N_28354);
or UO_2606 (O_2606,N_29879,N_28715);
xor UO_2607 (O_2607,N_29062,N_28195);
and UO_2608 (O_2608,N_29186,N_29759);
or UO_2609 (O_2609,N_29779,N_29832);
or UO_2610 (O_2610,N_29388,N_29802);
xnor UO_2611 (O_2611,N_29607,N_28980);
or UO_2612 (O_2612,N_29546,N_28201);
nand UO_2613 (O_2613,N_29430,N_29161);
or UO_2614 (O_2614,N_29514,N_28502);
or UO_2615 (O_2615,N_28495,N_28965);
nor UO_2616 (O_2616,N_28298,N_28580);
nor UO_2617 (O_2617,N_28239,N_29832);
nand UO_2618 (O_2618,N_28046,N_28062);
and UO_2619 (O_2619,N_28378,N_29894);
or UO_2620 (O_2620,N_28903,N_28956);
xnor UO_2621 (O_2621,N_28838,N_28419);
xnor UO_2622 (O_2622,N_28417,N_28202);
nand UO_2623 (O_2623,N_29285,N_28572);
nand UO_2624 (O_2624,N_28542,N_29053);
nand UO_2625 (O_2625,N_28758,N_29674);
nor UO_2626 (O_2626,N_29196,N_29344);
nor UO_2627 (O_2627,N_28519,N_28029);
or UO_2628 (O_2628,N_29444,N_29554);
and UO_2629 (O_2629,N_29702,N_29385);
nand UO_2630 (O_2630,N_28469,N_29306);
or UO_2631 (O_2631,N_29798,N_29473);
nor UO_2632 (O_2632,N_28115,N_29565);
and UO_2633 (O_2633,N_28661,N_29774);
or UO_2634 (O_2634,N_28761,N_29344);
xnor UO_2635 (O_2635,N_28107,N_28879);
nor UO_2636 (O_2636,N_29598,N_28150);
xnor UO_2637 (O_2637,N_28321,N_29937);
and UO_2638 (O_2638,N_28372,N_28284);
or UO_2639 (O_2639,N_29924,N_29535);
and UO_2640 (O_2640,N_28086,N_28366);
xnor UO_2641 (O_2641,N_28952,N_28643);
nor UO_2642 (O_2642,N_29985,N_29867);
nand UO_2643 (O_2643,N_29290,N_29408);
nor UO_2644 (O_2644,N_29141,N_28409);
and UO_2645 (O_2645,N_29634,N_29004);
or UO_2646 (O_2646,N_28683,N_28881);
xor UO_2647 (O_2647,N_28266,N_29030);
and UO_2648 (O_2648,N_29483,N_29655);
or UO_2649 (O_2649,N_28316,N_29747);
or UO_2650 (O_2650,N_28842,N_29113);
and UO_2651 (O_2651,N_29202,N_29828);
and UO_2652 (O_2652,N_28490,N_29087);
nor UO_2653 (O_2653,N_29849,N_29810);
nor UO_2654 (O_2654,N_28141,N_29046);
nand UO_2655 (O_2655,N_28682,N_29569);
nor UO_2656 (O_2656,N_29257,N_28972);
or UO_2657 (O_2657,N_28184,N_28285);
nor UO_2658 (O_2658,N_29968,N_29811);
and UO_2659 (O_2659,N_28927,N_29264);
or UO_2660 (O_2660,N_29763,N_29448);
nand UO_2661 (O_2661,N_28793,N_28448);
or UO_2662 (O_2662,N_28648,N_29899);
xor UO_2663 (O_2663,N_29271,N_29143);
xor UO_2664 (O_2664,N_29763,N_29683);
xor UO_2665 (O_2665,N_28027,N_28452);
or UO_2666 (O_2666,N_28149,N_28109);
nand UO_2667 (O_2667,N_29489,N_28415);
or UO_2668 (O_2668,N_28865,N_28004);
nand UO_2669 (O_2669,N_28403,N_28539);
nand UO_2670 (O_2670,N_29874,N_29803);
nand UO_2671 (O_2671,N_28484,N_29356);
and UO_2672 (O_2672,N_28932,N_29433);
nand UO_2673 (O_2673,N_28401,N_28222);
or UO_2674 (O_2674,N_29896,N_29343);
or UO_2675 (O_2675,N_29672,N_29489);
or UO_2676 (O_2676,N_28328,N_29367);
or UO_2677 (O_2677,N_29183,N_29949);
and UO_2678 (O_2678,N_29131,N_28719);
nor UO_2679 (O_2679,N_29729,N_29008);
nor UO_2680 (O_2680,N_29407,N_28052);
and UO_2681 (O_2681,N_28711,N_28407);
nand UO_2682 (O_2682,N_29455,N_28646);
nand UO_2683 (O_2683,N_28923,N_28154);
and UO_2684 (O_2684,N_28086,N_28429);
nor UO_2685 (O_2685,N_28000,N_28352);
xnor UO_2686 (O_2686,N_29020,N_29492);
and UO_2687 (O_2687,N_29335,N_29248);
or UO_2688 (O_2688,N_29365,N_29052);
nand UO_2689 (O_2689,N_29666,N_29349);
nand UO_2690 (O_2690,N_28415,N_28392);
nand UO_2691 (O_2691,N_29407,N_28594);
nand UO_2692 (O_2692,N_29169,N_28155);
or UO_2693 (O_2693,N_29686,N_28716);
nand UO_2694 (O_2694,N_28786,N_29243);
and UO_2695 (O_2695,N_28396,N_28990);
nor UO_2696 (O_2696,N_29774,N_28764);
nand UO_2697 (O_2697,N_28211,N_28929);
or UO_2698 (O_2698,N_29607,N_29611);
nor UO_2699 (O_2699,N_28710,N_29117);
and UO_2700 (O_2700,N_28140,N_28780);
and UO_2701 (O_2701,N_28134,N_28676);
and UO_2702 (O_2702,N_28185,N_29913);
nor UO_2703 (O_2703,N_28419,N_28329);
nor UO_2704 (O_2704,N_28431,N_28698);
nand UO_2705 (O_2705,N_29918,N_29890);
nand UO_2706 (O_2706,N_28514,N_28695);
or UO_2707 (O_2707,N_28469,N_28162);
nand UO_2708 (O_2708,N_28009,N_28312);
or UO_2709 (O_2709,N_28900,N_29914);
and UO_2710 (O_2710,N_29035,N_28638);
nor UO_2711 (O_2711,N_28699,N_28225);
nand UO_2712 (O_2712,N_28088,N_28849);
and UO_2713 (O_2713,N_28295,N_28169);
nor UO_2714 (O_2714,N_29303,N_28384);
nor UO_2715 (O_2715,N_29783,N_28607);
or UO_2716 (O_2716,N_29006,N_29658);
nand UO_2717 (O_2717,N_29662,N_29174);
xor UO_2718 (O_2718,N_28726,N_29454);
nor UO_2719 (O_2719,N_29980,N_28626);
nand UO_2720 (O_2720,N_29832,N_28686);
and UO_2721 (O_2721,N_29029,N_28804);
xor UO_2722 (O_2722,N_29721,N_29748);
xnor UO_2723 (O_2723,N_28441,N_29592);
nor UO_2724 (O_2724,N_29127,N_28160);
xnor UO_2725 (O_2725,N_29598,N_29747);
and UO_2726 (O_2726,N_29862,N_29417);
and UO_2727 (O_2727,N_28260,N_29087);
nor UO_2728 (O_2728,N_28353,N_29023);
xnor UO_2729 (O_2729,N_29720,N_28254);
xnor UO_2730 (O_2730,N_29980,N_29385);
xor UO_2731 (O_2731,N_29888,N_28744);
nor UO_2732 (O_2732,N_28195,N_29213);
xor UO_2733 (O_2733,N_28967,N_28823);
xor UO_2734 (O_2734,N_28890,N_29489);
nand UO_2735 (O_2735,N_29038,N_28023);
and UO_2736 (O_2736,N_29279,N_28307);
and UO_2737 (O_2737,N_28496,N_29497);
and UO_2738 (O_2738,N_28870,N_29668);
xnor UO_2739 (O_2739,N_28579,N_29647);
nand UO_2740 (O_2740,N_29700,N_29748);
or UO_2741 (O_2741,N_28573,N_29299);
nand UO_2742 (O_2742,N_29109,N_29926);
and UO_2743 (O_2743,N_28025,N_29836);
nor UO_2744 (O_2744,N_29027,N_28532);
xor UO_2745 (O_2745,N_29679,N_28237);
nand UO_2746 (O_2746,N_28646,N_28970);
and UO_2747 (O_2747,N_28073,N_29087);
or UO_2748 (O_2748,N_29475,N_29736);
xnor UO_2749 (O_2749,N_29081,N_28663);
and UO_2750 (O_2750,N_29586,N_29228);
xor UO_2751 (O_2751,N_29223,N_28853);
xor UO_2752 (O_2752,N_29054,N_28323);
nand UO_2753 (O_2753,N_28467,N_29279);
nand UO_2754 (O_2754,N_29244,N_29756);
nand UO_2755 (O_2755,N_28365,N_28661);
or UO_2756 (O_2756,N_28295,N_28877);
nor UO_2757 (O_2757,N_29259,N_28650);
or UO_2758 (O_2758,N_28984,N_28445);
xnor UO_2759 (O_2759,N_29927,N_29232);
and UO_2760 (O_2760,N_29629,N_29126);
xor UO_2761 (O_2761,N_29769,N_29458);
xor UO_2762 (O_2762,N_29270,N_28725);
or UO_2763 (O_2763,N_28161,N_29063);
and UO_2764 (O_2764,N_29317,N_28978);
xor UO_2765 (O_2765,N_28955,N_28032);
and UO_2766 (O_2766,N_29992,N_29122);
or UO_2767 (O_2767,N_29902,N_29703);
or UO_2768 (O_2768,N_29386,N_28495);
or UO_2769 (O_2769,N_29349,N_28619);
nand UO_2770 (O_2770,N_29108,N_28224);
xor UO_2771 (O_2771,N_28031,N_29264);
nor UO_2772 (O_2772,N_29323,N_28811);
xor UO_2773 (O_2773,N_28234,N_28184);
or UO_2774 (O_2774,N_28897,N_28652);
xnor UO_2775 (O_2775,N_29598,N_28408);
and UO_2776 (O_2776,N_28876,N_28189);
nor UO_2777 (O_2777,N_29999,N_28787);
nand UO_2778 (O_2778,N_28645,N_28341);
nand UO_2779 (O_2779,N_28303,N_28242);
and UO_2780 (O_2780,N_28559,N_28736);
xor UO_2781 (O_2781,N_29028,N_29659);
nand UO_2782 (O_2782,N_29479,N_29724);
xor UO_2783 (O_2783,N_29223,N_29027);
xnor UO_2784 (O_2784,N_28376,N_28011);
nor UO_2785 (O_2785,N_29709,N_29710);
nand UO_2786 (O_2786,N_28515,N_29499);
and UO_2787 (O_2787,N_28301,N_29962);
or UO_2788 (O_2788,N_28558,N_29576);
nor UO_2789 (O_2789,N_29190,N_29807);
or UO_2790 (O_2790,N_29150,N_28297);
or UO_2791 (O_2791,N_28618,N_29636);
or UO_2792 (O_2792,N_28777,N_28792);
and UO_2793 (O_2793,N_28365,N_29727);
xnor UO_2794 (O_2794,N_28426,N_29116);
and UO_2795 (O_2795,N_29154,N_29598);
nand UO_2796 (O_2796,N_28642,N_29021);
xor UO_2797 (O_2797,N_28053,N_29738);
nor UO_2798 (O_2798,N_29981,N_28034);
nand UO_2799 (O_2799,N_28004,N_29507);
nand UO_2800 (O_2800,N_28975,N_28779);
or UO_2801 (O_2801,N_29952,N_29554);
or UO_2802 (O_2802,N_29294,N_28211);
nor UO_2803 (O_2803,N_29552,N_29587);
or UO_2804 (O_2804,N_29439,N_29402);
nor UO_2805 (O_2805,N_28689,N_29219);
and UO_2806 (O_2806,N_28803,N_29302);
xor UO_2807 (O_2807,N_28357,N_28867);
nand UO_2808 (O_2808,N_28710,N_29079);
nand UO_2809 (O_2809,N_28586,N_28587);
and UO_2810 (O_2810,N_28036,N_29376);
or UO_2811 (O_2811,N_29731,N_29204);
xor UO_2812 (O_2812,N_28175,N_28407);
nor UO_2813 (O_2813,N_29184,N_28741);
and UO_2814 (O_2814,N_28522,N_29630);
nor UO_2815 (O_2815,N_28315,N_28132);
and UO_2816 (O_2816,N_28577,N_28872);
nor UO_2817 (O_2817,N_28058,N_28616);
and UO_2818 (O_2818,N_28344,N_28868);
or UO_2819 (O_2819,N_29954,N_29705);
or UO_2820 (O_2820,N_28203,N_29093);
xnor UO_2821 (O_2821,N_29407,N_29165);
nand UO_2822 (O_2822,N_29401,N_29459);
and UO_2823 (O_2823,N_28609,N_28495);
nand UO_2824 (O_2824,N_29630,N_28643);
nor UO_2825 (O_2825,N_28815,N_28369);
and UO_2826 (O_2826,N_28958,N_28486);
and UO_2827 (O_2827,N_29914,N_29503);
nand UO_2828 (O_2828,N_29521,N_29364);
nand UO_2829 (O_2829,N_28718,N_28218);
nand UO_2830 (O_2830,N_29537,N_29634);
nand UO_2831 (O_2831,N_28747,N_29080);
xnor UO_2832 (O_2832,N_28140,N_28787);
nor UO_2833 (O_2833,N_28338,N_29354);
nor UO_2834 (O_2834,N_29197,N_28059);
or UO_2835 (O_2835,N_29324,N_29296);
nand UO_2836 (O_2836,N_29830,N_28972);
or UO_2837 (O_2837,N_29653,N_28564);
xnor UO_2838 (O_2838,N_28621,N_29368);
or UO_2839 (O_2839,N_28369,N_29528);
xor UO_2840 (O_2840,N_29533,N_29600);
or UO_2841 (O_2841,N_28138,N_29337);
and UO_2842 (O_2842,N_29741,N_28235);
or UO_2843 (O_2843,N_29483,N_28989);
xor UO_2844 (O_2844,N_28453,N_29551);
xnor UO_2845 (O_2845,N_28581,N_28910);
or UO_2846 (O_2846,N_29100,N_29002);
xnor UO_2847 (O_2847,N_29037,N_28375);
nand UO_2848 (O_2848,N_28655,N_29485);
and UO_2849 (O_2849,N_28806,N_29583);
nand UO_2850 (O_2850,N_28402,N_29874);
nor UO_2851 (O_2851,N_28213,N_28695);
nor UO_2852 (O_2852,N_28381,N_28000);
xor UO_2853 (O_2853,N_28161,N_29180);
and UO_2854 (O_2854,N_29074,N_28777);
xnor UO_2855 (O_2855,N_28606,N_28218);
nand UO_2856 (O_2856,N_29863,N_28057);
nor UO_2857 (O_2857,N_28164,N_28028);
xnor UO_2858 (O_2858,N_29385,N_29423);
or UO_2859 (O_2859,N_29312,N_29417);
xor UO_2860 (O_2860,N_29096,N_29057);
or UO_2861 (O_2861,N_29350,N_28720);
xnor UO_2862 (O_2862,N_28310,N_28139);
nand UO_2863 (O_2863,N_28969,N_29379);
and UO_2864 (O_2864,N_28171,N_28571);
nand UO_2865 (O_2865,N_28469,N_28670);
nor UO_2866 (O_2866,N_28857,N_28720);
and UO_2867 (O_2867,N_28266,N_28424);
nand UO_2868 (O_2868,N_28481,N_28636);
and UO_2869 (O_2869,N_28352,N_28575);
and UO_2870 (O_2870,N_28509,N_28879);
or UO_2871 (O_2871,N_29648,N_28403);
nand UO_2872 (O_2872,N_28878,N_28877);
or UO_2873 (O_2873,N_29190,N_28772);
or UO_2874 (O_2874,N_28324,N_28033);
and UO_2875 (O_2875,N_28748,N_28920);
and UO_2876 (O_2876,N_28573,N_28390);
xnor UO_2877 (O_2877,N_28997,N_29987);
and UO_2878 (O_2878,N_28593,N_29003);
and UO_2879 (O_2879,N_28826,N_29797);
nor UO_2880 (O_2880,N_28015,N_29153);
xor UO_2881 (O_2881,N_28557,N_29142);
nor UO_2882 (O_2882,N_28804,N_28482);
nor UO_2883 (O_2883,N_28353,N_28992);
xor UO_2884 (O_2884,N_29670,N_28265);
or UO_2885 (O_2885,N_29731,N_28818);
and UO_2886 (O_2886,N_29505,N_28758);
and UO_2887 (O_2887,N_29444,N_28207);
nand UO_2888 (O_2888,N_29995,N_28296);
nor UO_2889 (O_2889,N_29582,N_29549);
nor UO_2890 (O_2890,N_28250,N_28290);
or UO_2891 (O_2891,N_29989,N_28146);
or UO_2892 (O_2892,N_29194,N_28047);
nand UO_2893 (O_2893,N_29450,N_29187);
nor UO_2894 (O_2894,N_28422,N_29866);
and UO_2895 (O_2895,N_29061,N_29863);
and UO_2896 (O_2896,N_28003,N_28060);
and UO_2897 (O_2897,N_29293,N_29484);
nand UO_2898 (O_2898,N_29748,N_28126);
or UO_2899 (O_2899,N_28310,N_29374);
and UO_2900 (O_2900,N_29564,N_29032);
xor UO_2901 (O_2901,N_29152,N_28294);
nor UO_2902 (O_2902,N_28736,N_29980);
xor UO_2903 (O_2903,N_28656,N_29584);
nor UO_2904 (O_2904,N_29423,N_29392);
nor UO_2905 (O_2905,N_28003,N_28124);
xnor UO_2906 (O_2906,N_28202,N_28364);
nor UO_2907 (O_2907,N_29907,N_29659);
nand UO_2908 (O_2908,N_28213,N_28193);
nor UO_2909 (O_2909,N_28974,N_28860);
nand UO_2910 (O_2910,N_28321,N_29467);
or UO_2911 (O_2911,N_28762,N_29426);
or UO_2912 (O_2912,N_29245,N_29682);
nand UO_2913 (O_2913,N_28640,N_28781);
or UO_2914 (O_2914,N_28284,N_29085);
xnor UO_2915 (O_2915,N_29011,N_28265);
and UO_2916 (O_2916,N_28045,N_28452);
nor UO_2917 (O_2917,N_28735,N_28363);
nand UO_2918 (O_2918,N_29235,N_29803);
nand UO_2919 (O_2919,N_28521,N_28962);
xor UO_2920 (O_2920,N_29928,N_29391);
and UO_2921 (O_2921,N_29168,N_28222);
and UO_2922 (O_2922,N_29257,N_29745);
and UO_2923 (O_2923,N_28876,N_28923);
or UO_2924 (O_2924,N_29604,N_28648);
nand UO_2925 (O_2925,N_29342,N_29796);
nor UO_2926 (O_2926,N_28481,N_29691);
xor UO_2927 (O_2927,N_29358,N_28938);
nand UO_2928 (O_2928,N_28616,N_28073);
or UO_2929 (O_2929,N_28780,N_28276);
nor UO_2930 (O_2930,N_28896,N_28302);
or UO_2931 (O_2931,N_29755,N_28651);
xor UO_2932 (O_2932,N_29562,N_29564);
nor UO_2933 (O_2933,N_28325,N_29693);
nand UO_2934 (O_2934,N_28674,N_28205);
and UO_2935 (O_2935,N_29441,N_28295);
nor UO_2936 (O_2936,N_29262,N_29891);
and UO_2937 (O_2937,N_29415,N_28046);
xor UO_2938 (O_2938,N_28440,N_28613);
or UO_2939 (O_2939,N_28926,N_29117);
and UO_2940 (O_2940,N_28298,N_28977);
or UO_2941 (O_2941,N_28188,N_29909);
nor UO_2942 (O_2942,N_29142,N_28631);
or UO_2943 (O_2943,N_29932,N_28696);
nor UO_2944 (O_2944,N_29213,N_29423);
and UO_2945 (O_2945,N_29522,N_29367);
and UO_2946 (O_2946,N_28004,N_29431);
xor UO_2947 (O_2947,N_29131,N_29913);
or UO_2948 (O_2948,N_29501,N_29095);
or UO_2949 (O_2949,N_29045,N_29171);
nand UO_2950 (O_2950,N_29599,N_28436);
nor UO_2951 (O_2951,N_29049,N_28977);
nand UO_2952 (O_2952,N_29266,N_29737);
nand UO_2953 (O_2953,N_28115,N_28797);
or UO_2954 (O_2954,N_28505,N_28237);
or UO_2955 (O_2955,N_29042,N_29577);
and UO_2956 (O_2956,N_29883,N_28228);
nor UO_2957 (O_2957,N_29475,N_28245);
nor UO_2958 (O_2958,N_29113,N_29584);
or UO_2959 (O_2959,N_28131,N_28992);
xnor UO_2960 (O_2960,N_28971,N_28196);
nor UO_2961 (O_2961,N_29571,N_29692);
nor UO_2962 (O_2962,N_28662,N_29634);
or UO_2963 (O_2963,N_29230,N_28533);
and UO_2964 (O_2964,N_29097,N_29130);
nand UO_2965 (O_2965,N_28169,N_28047);
nor UO_2966 (O_2966,N_28092,N_29486);
and UO_2967 (O_2967,N_29484,N_28383);
nand UO_2968 (O_2968,N_29647,N_29716);
and UO_2969 (O_2969,N_28851,N_29590);
nor UO_2970 (O_2970,N_28181,N_28409);
nor UO_2971 (O_2971,N_29078,N_29842);
and UO_2972 (O_2972,N_29992,N_28081);
and UO_2973 (O_2973,N_29713,N_29351);
and UO_2974 (O_2974,N_28787,N_28458);
and UO_2975 (O_2975,N_28581,N_29603);
xnor UO_2976 (O_2976,N_29760,N_29824);
or UO_2977 (O_2977,N_28184,N_28284);
and UO_2978 (O_2978,N_28303,N_29458);
nand UO_2979 (O_2979,N_28363,N_28697);
and UO_2980 (O_2980,N_29250,N_29782);
or UO_2981 (O_2981,N_28998,N_29191);
nand UO_2982 (O_2982,N_29312,N_29140);
nand UO_2983 (O_2983,N_28238,N_28807);
nand UO_2984 (O_2984,N_29366,N_28419);
or UO_2985 (O_2985,N_28642,N_29462);
nor UO_2986 (O_2986,N_28702,N_29714);
xor UO_2987 (O_2987,N_28722,N_28703);
and UO_2988 (O_2988,N_29259,N_28035);
nor UO_2989 (O_2989,N_28953,N_28610);
and UO_2990 (O_2990,N_28568,N_29490);
and UO_2991 (O_2991,N_28184,N_29727);
nor UO_2992 (O_2992,N_29128,N_28054);
nor UO_2993 (O_2993,N_29478,N_29957);
nand UO_2994 (O_2994,N_29926,N_29638);
nor UO_2995 (O_2995,N_29039,N_28204);
nand UO_2996 (O_2996,N_29904,N_29949);
xnor UO_2997 (O_2997,N_28191,N_28754);
nor UO_2998 (O_2998,N_28169,N_28788);
nor UO_2999 (O_2999,N_29981,N_28388);
xnor UO_3000 (O_3000,N_28201,N_28018);
nand UO_3001 (O_3001,N_29260,N_28720);
nand UO_3002 (O_3002,N_29212,N_28334);
nor UO_3003 (O_3003,N_29435,N_29507);
and UO_3004 (O_3004,N_28532,N_29974);
and UO_3005 (O_3005,N_28834,N_28453);
nand UO_3006 (O_3006,N_28985,N_28074);
and UO_3007 (O_3007,N_28859,N_29765);
nor UO_3008 (O_3008,N_28101,N_28120);
nor UO_3009 (O_3009,N_29783,N_28186);
nand UO_3010 (O_3010,N_29377,N_28085);
or UO_3011 (O_3011,N_28262,N_29310);
nand UO_3012 (O_3012,N_28773,N_28721);
xnor UO_3013 (O_3013,N_28107,N_28854);
or UO_3014 (O_3014,N_28251,N_29243);
and UO_3015 (O_3015,N_29917,N_29456);
nand UO_3016 (O_3016,N_28193,N_28045);
nand UO_3017 (O_3017,N_29074,N_28465);
or UO_3018 (O_3018,N_28612,N_29278);
nor UO_3019 (O_3019,N_29380,N_28864);
or UO_3020 (O_3020,N_28010,N_29247);
nand UO_3021 (O_3021,N_28260,N_28449);
nand UO_3022 (O_3022,N_29828,N_28358);
or UO_3023 (O_3023,N_29685,N_29359);
nor UO_3024 (O_3024,N_28541,N_29040);
or UO_3025 (O_3025,N_29350,N_28798);
or UO_3026 (O_3026,N_28308,N_29086);
and UO_3027 (O_3027,N_29632,N_28588);
nand UO_3028 (O_3028,N_29078,N_28195);
nand UO_3029 (O_3029,N_28225,N_29286);
nor UO_3030 (O_3030,N_28994,N_28393);
or UO_3031 (O_3031,N_29353,N_29643);
xor UO_3032 (O_3032,N_29333,N_29371);
xnor UO_3033 (O_3033,N_28516,N_29961);
nor UO_3034 (O_3034,N_29270,N_28323);
nor UO_3035 (O_3035,N_28058,N_29085);
xnor UO_3036 (O_3036,N_28851,N_29094);
xnor UO_3037 (O_3037,N_29213,N_28439);
nand UO_3038 (O_3038,N_29292,N_28421);
or UO_3039 (O_3039,N_28924,N_28396);
and UO_3040 (O_3040,N_28968,N_28893);
xor UO_3041 (O_3041,N_28616,N_29744);
or UO_3042 (O_3042,N_29085,N_28405);
nor UO_3043 (O_3043,N_29256,N_28831);
nand UO_3044 (O_3044,N_29717,N_28583);
nand UO_3045 (O_3045,N_28944,N_28899);
nand UO_3046 (O_3046,N_29259,N_28286);
and UO_3047 (O_3047,N_29782,N_28737);
nor UO_3048 (O_3048,N_28729,N_28780);
xnor UO_3049 (O_3049,N_28550,N_28976);
and UO_3050 (O_3050,N_29685,N_28955);
nor UO_3051 (O_3051,N_28295,N_28503);
nor UO_3052 (O_3052,N_29475,N_28980);
or UO_3053 (O_3053,N_29606,N_28496);
xnor UO_3054 (O_3054,N_29092,N_28429);
nand UO_3055 (O_3055,N_29621,N_28953);
nand UO_3056 (O_3056,N_29607,N_28080);
or UO_3057 (O_3057,N_29667,N_28671);
or UO_3058 (O_3058,N_28065,N_28632);
nor UO_3059 (O_3059,N_28648,N_28154);
xnor UO_3060 (O_3060,N_28800,N_29516);
nand UO_3061 (O_3061,N_29203,N_29752);
and UO_3062 (O_3062,N_28077,N_29702);
xor UO_3063 (O_3063,N_29391,N_28921);
and UO_3064 (O_3064,N_28374,N_29939);
nand UO_3065 (O_3065,N_28095,N_29073);
nand UO_3066 (O_3066,N_29325,N_29281);
nor UO_3067 (O_3067,N_28463,N_29065);
nor UO_3068 (O_3068,N_28400,N_29645);
or UO_3069 (O_3069,N_29366,N_28659);
xnor UO_3070 (O_3070,N_28825,N_28943);
nor UO_3071 (O_3071,N_29616,N_29739);
or UO_3072 (O_3072,N_28927,N_28259);
and UO_3073 (O_3073,N_28024,N_28991);
nand UO_3074 (O_3074,N_28685,N_29675);
and UO_3075 (O_3075,N_28262,N_28014);
nor UO_3076 (O_3076,N_29469,N_28968);
nor UO_3077 (O_3077,N_28453,N_28539);
xor UO_3078 (O_3078,N_28113,N_29137);
nor UO_3079 (O_3079,N_28514,N_29725);
nor UO_3080 (O_3080,N_28159,N_29710);
or UO_3081 (O_3081,N_28148,N_29043);
xor UO_3082 (O_3082,N_28859,N_29377);
xnor UO_3083 (O_3083,N_29243,N_29590);
or UO_3084 (O_3084,N_29624,N_28637);
nor UO_3085 (O_3085,N_29581,N_29655);
nor UO_3086 (O_3086,N_28802,N_29232);
xor UO_3087 (O_3087,N_29025,N_28080);
nor UO_3088 (O_3088,N_29276,N_28983);
and UO_3089 (O_3089,N_28188,N_28569);
nand UO_3090 (O_3090,N_29510,N_29063);
xnor UO_3091 (O_3091,N_29143,N_28244);
and UO_3092 (O_3092,N_29366,N_29074);
or UO_3093 (O_3093,N_28051,N_28982);
nor UO_3094 (O_3094,N_29465,N_28158);
xor UO_3095 (O_3095,N_28698,N_28055);
nand UO_3096 (O_3096,N_28676,N_29116);
and UO_3097 (O_3097,N_29140,N_29342);
xnor UO_3098 (O_3098,N_29893,N_29228);
nor UO_3099 (O_3099,N_29473,N_28890);
nand UO_3100 (O_3100,N_29602,N_29770);
xnor UO_3101 (O_3101,N_28697,N_28595);
and UO_3102 (O_3102,N_28512,N_28061);
nor UO_3103 (O_3103,N_28114,N_28751);
xnor UO_3104 (O_3104,N_29546,N_29543);
nor UO_3105 (O_3105,N_28539,N_28802);
xor UO_3106 (O_3106,N_28420,N_29331);
or UO_3107 (O_3107,N_29740,N_29244);
xor UO_3108 (O_3108,N_28701,N_29253);
xnor UO_3109 (O_3109,N_28226,N_29422);
xor UO_3110 (O_3110,N_28544,N_29809);
nor UO_3111 (O_3111,N_28007,N_29692);
or UO_3112 (O_3112,N_29975,N_28994);
nand UO_3113 (O_3113,N_28566,N_28051);
xor UO_3114 (O_3114,N_29524,N_28231);
nor UO_3115 (O_3115,N_29825,N_28895);
nand UO_3116 (O_3116,N_28843,N_29265);
and UO_3117 (O_3117,N_28879,N_29394);
nand UO_3118 (O_3118,N_28417,N_28631);
nor UO_3119 (O_3119,N_29778,N_28228);
or UO_3120 (O_3120,N_28158,N_28830);
nor UO_3121 (O_3121,N_28513,N_28759);
xnor UO_3122 (O_3122,N_28462,N_28082);
nand UO_3123 (O_3123,N_29851,N_29777);
or UO_3124 (O_3124,N_28289,N_29278);
xor UO_3125 (O_3125,N_28837,N_28716);
nor UO_3126 (O_3126,N_28554,N_29086);
nand UO_3127 (O_3127,N_29900,N_29399);
nand UO_3128 (O_3128,N_28996,N_28689);
xor UO_3129 (O_3129,N_29224,N_29467);
or UO_3130 (O_3130,N_28261,N_28734);
and UO_3131 (O_3131,N_29579,N_28801);
or UO_3132 (O_3132,N_29472,N_28808);
nor UO_3133 (O_3133,N_29544,N_28708);
nor UO_3134 (O_3134,N_29790,N_28095);
or UO_3135 (O_3135,N_28263,N_28790);
nor UO_3136 (O_3136,N_29692,N_29456);
nor UO_3137 (O_3137,N_29503,N_28788);
nor UO_3138 (O_3138,N_29896,N_28978);
xor UO_3139 (O_3139,N_28922,N_29120);
nand UO_3140 (O_3140,N_28458,N_28597);
and UO_3141 (O_3141,N_28049,N_28842);
nand UO_3142 (O_3142,N_28979,N_29608);
or UO_3143 (O_3143,N_29746,N_28629);
nor UO_3144 (O_3144,N_28931,N_29311);
nand UO_3145 (O_3145,N_29032,N_29990);
nand UO_3146 (O_3146,N_29960,N_29236);
and UO_3147 (O_3147,N_29070,N_29848);
and UO_3148 (O_3148,N_29535,N_29637);
nand UO_3149 (O_3149,N_29966,N_28070);
xor UO_3150 (O_3150,N_28598,N_29805);
xor UO_3151 (O_3151,N_28174,N_28208);
xor UO_3152 (O_3152,N_29262,N_28566);
nor UO_3153 (O_3153,N_28585,N_29216);
nand UO_3154 (O_3154,N_28701,N_28753);
nand UO_3155 (O_3155,N_28407,N_28842);
or UO_3156 (O_3156,N_29604,N_29579);
or UO_3157 (O_3157,N_29350,N_29180);
and UO_3158 (O_3158,N_29165,N_28630);
and UO_3159 (O_3159,N_29360,N_29269);
and UO_3160 (O_3160,N_29693,N_28121);
or UO_3161 (O_3161,N_28065,N_29772);
nor UO_3162 (O_3162,N_29447,N_28244);
xnor UO_3163 (O_3163,N_28057,N_28132);
xnor UO_3164 (O_3164,N_28362,N_28426);
xnor UO_3165 (O_3165,N_28459,N_29394);
nor UO_3166 (O_3166,N_28120,N_28268);
xor UO_3167 (O_3167,N_29798,N_28219);
or UO_3168 (O_3168,N_28850,N_29458);
xor UO_3169 (O_3169,N_29383,N_28060);
xor UO_3170 (O_3170,N_29868,N_29416);
and UO_3171 (O_3171,N_28037,N_29650);
nor UO_3172 (O_3172,N_29379,N_29173);
or UO_3173 (O_3173,N_28188,N_29215);
and UO_3174 (O_3174,N_29781,N_28533);
nor UO_3175 (O_3175,N_28632,N_29526);
or UO_3176 (O_3176,N_28006,N_29043);
and UO_3177 (O_3177,N_29565,N_28974);
nand UO_3178 (O_3178,N_28182,N_29779);
nor UO_3179 (O_3179,N_29610,N_29474);
or UO_3180 (O_3180,N_29284,N_29836);
nand UO_3181 (O_3181,N_29095,N_29613);
nor UO_3182 (O_3182,N_29527,N_29736);
xnor UO_3183 (O_3183,N_28914,N_28192);
xor UO_3184 (O_3184,N_29845,N_29271);
xnor UO_3185 (O_3185,N_28552,N_29513);
nand UO_3186 (O_3186,N_28297,N_28682);
or UO_3187 (O_3187,N_28978,N_28705);
and UO_3188 (O_3188,N_29441,N_29620);
xor UO_3189 (O_3189,N_29854,N_28447);
nor UO_3190 (O_3190,N_29540,N_28285);
or UO_3191 (O_3191,N_28516,N_29199);
or UO_3192 (O_3192,N_29740,N_29346);
and UO_3193 (O_3193,N_29353,N_29463);
xnor UO_3194 (O_3194,N_28317,N_29268);
or UO_3195 (O_3195,N_28908,N_29966);
or UO_3196 (O_3196,N_28912,N_28772);
or UO_3197 (O_3197,N_29130,N_28834);
or UO_3198 (O_3198,N_29956,N_29807);
nand UO_3199 (O_3199,N_29257,N_28804);
and UO_3200 (O_3200,N_28444,N_29539);
and UO_3201 (O_3201,N_28236,N_28454);
nand UO_3202 (O_3202,N_28625,N_29489);
nor UO_3203 (O_3203,N_28979,N_29965);
xor UO_3204 (O_3204,N_29568,N_29812);
and UO_3205 (O_3205,N_28024,N_29126);
xnor UO_3206 (O_3206,N_29600,N_28627);
nand UO_3207 (O_3207,N_28535,N_29652);
nor UO_3208 (O_3208,N_28158,N_28680);
xnor UO_3209 (O_3209,N_29375,N_28144);
xor UO_3210 (O_3210,N_28218,N_29843);
or UO_3211 (O_3211,N_29957,N_28550);
and UO_3212 (O_3212,N_29093,N_29766);
nand UO_3213 (O_3213,N_29744,N_29867);
xor UO_3214 (O_3214,N_28658,N_29233);
xor UO_3215 (O_3215,N_28071,N_28429);
and UO_3216 (O_3216,N_28712,N_29749);
nand UO_3217 (O_3217,N_29675,N_29364);
xor UO_3218 (O_3218,N_29562,N_28005);
nor UO_3219 (O_3219,N_29059,N_28308);
nand UO_3220 (O_3220,N_29336,N_29380);
nand UO_3221 (O_3221,N_28296,N_28281);
or UO_3222 (O_3222,N_28025,N_29438);
and UO_3223 (O_3223,N_29227,N_28611);
or UO_3224 (O_3224,N_29616,N_28395);
xor UO_3225 (O_3225,N_28125,N_29508);
nor UO_3226 (O_3226,N_29033,N_29574);
nand UO_3227 (O_3227,N_28088,N_29270);
nand UO_3228 (O_3228,N_29033,N_28915);
and UO_3229 (O_3229,N_28830,N_28986);
nand UO_3230 (O_3230,N_28812,N_29709);
and UO_3231 (O_3231,N_28071,N_29998);
or UO_3232 (O_3232,N_29773,N_29245);
nor UO_3233 (O_3233,N_28322,N_28378);
and UO_3234 (O_3234,N_29138,N_29218);
xor UO_3235 (O_3235,N_28367,N_29967);
xnor UO_3236 (O_3236,N_28194,N_28331);
nand UO_3237 (O_3237,N_29159,N_29440);
nand UO_3238 (O_3238,N_29714,N_28455);
nand UO_3239 (O_3239,N_29579,N_29256);
and UO_3240 (O_3240,N_29927,N_28895);
and UO_3241 (O_3241,N_29755,N_28592);
xnor UO_3242 (O_3242,N_28349,N_29833);
xnor UO_3243 (O_3243,N_28598,N_28826);
nand UO_3244 (O_3244,N_29212,N_29250);
xor UO_3245 (O_3245,N_28805,N_29756);
and UO_3246 (O_3246,N_29785,N_28509);
xnor UO_3247 (O_3247,N_29428,N_29550);
xnor UO_3248 (O_3248,N_28911,N_29637);
and UO_3249 (O_3249,N_28659,N_28759);
and UO_3250 (O_3250,N_28982,N_29466);
nand UO_3251 (O_3251,N_29006,N_28095);
and UO_3252 (O_3252,N_28427,N_28693);
and UO_3253 (O_3253,N_29335,N_29647);
xor UO_3254 (O_3254,N_29309,N_28646);
or UO_3255 (O_3255,N_28342,N_28174);
nor UO_3256 (O_3256,N_28962,N_29475);
and UO_3257 (O_3257,N_28854,N_29650);
nor UO_3258 (O_3258,N_29897,N_28367);
or UO_3259 (O_3259,N_28584,N_29022);
and UO_3260 (O_3260,N_28772,N_28602);
xnor UO_3261 (O_3261,N_28448,N_29497);
nor UO_3262 (O_3262,N_28420,N_29389);
xor UO_3263 (O_3263,N_28260,N_28769);
nor UO_3264 (O_3264,N_28814,N_28713);
nand UO_3265 (O_3265,N_29154,N_28184);
nand UO_3266 (O_3266,N_29017,N_28831);
or UO_3267 (O_3267,N_29592,N_29830);
and UO_3268 (O_3268,N_28339,N_29627);
nor UO_3269 (O_3269,N_29127,N_28841);
xor UO_3270 (O_3270,N_28786,N_29555);
xnor UO_3271 (O_3271,N_29949,N_29119);
nand UO_3272 (O_3272,N_28310,N_29279);
xnor UO_3273 (O_3273,N_29965,N_29121);
xor UO_3274 (O_3274,N_28190,N_28359);
nor UO_3275 (O_3275,N_28643,N_28512);
or UO_3276 (O_3276,N_28481,N_28297);
or UO_3277 (O_3277,N_28865,N_28217);
or UO_3278 (O_3278,N_28239,N_28317);
or UO_3279 (O_3279,N_28222,N_28236);
xor UO_3280 (O_3280,N_29983,N_29574);
xor UO_3281 (O_3281,N_29589,N_28357);
xor UO_3282 (O_3282,N_28729,N_28119);
nor UO_3283 (O_3283,N_28649,N_29758);
or UO_3284 (O_3284,N_28467,N_28920);
xnor UO_3285 (O_3285,N_29582,N_29338);
nor UO_3286 (O_3286,N_29136,N_29651);
and UO_3287 (O_3287,N_28295,N_29179);
nor UO_3288 (O_3288,N_28103,N_28382);
nand UO_3289 (O_3289,N_29113,N_28449);
and UO_3290 (O_3290,N_29553,N_29191);
nor UO_3291 (O_3291,N_28786,N_29625);
and UO_3292 (O_3292,N_28947,N_28576);
nand UO_3293 (O_3293,N_29093,N_29898);
or UO_3294 (O_3294,N_29605,N_29715);
nand UO_3295 (O_3295,N_29972,N_29453);
nand UO_3296 (O_3296,N_28778,N_28170);
or UO_3297 (O_3297,N_29201,N_29736);
or UO_3298 (O_3298,N_29561,N_28919);
and UO_3299 (O_3299,N_29262,N_28745);
xnor UO_3300 (O_3300,N_29098,N_29025);
nand UO_3301 (O_3301,N_28901,N_28778);
nand UO_3302 (O_3302,N_29570,N_29489);
or UO_3303 (O_3303,N_29609,N_29719);
and UO_3304 (O_3304,N_28250,N_28416);
nand UO_3305 (O_3305,N_28317,N_29695);
nand UO_3306 (O_3306,N_28992,N_28380);
or UO_3307 (O_3307,N_28668,N_29037);
nand UO_3308 (O_3308,N_29028,N_28407);
nor UO_3309 (O_3309,N_29295,N_29748);
or UO_3310 (O_3310,N_29921,N_29342);
and UO_3311 (O_3311,N_29677,N_29307);
nand UO_3312 (O_3312,N_29323,N_28435);
or UO_3313 (O_3313,N_28047,N_29839);
xnor UO_3314 (O_3314,N_28772,N_28041);
xor UO_3315 (O_3315,N_29909,N_29123);
nand UO_3316 (O_3316,N_29678,N_29224);
nand UO_3317 (O_3317,N_28025,N_28810);
xnor UO_3318 (O_3318,N_29232,N_29070);
or UO_3319 (O_3319,N_29617,N_29295);
or UO_3320 (O_3320,N_29956,N_28877);
xor UO_3321 (O_3321,N_29680,N_29823);
xor UO_3322 (O_3322,N_29039,N_29197);
and UO_3323 (O_3323,N_28621,N_28098);
and UO_3324 (O_3324,N_28653,N_28845);
and UO_3325 (O_3325,N_28703,N_29644);
nor UO_3326 (O_3326,N_28746,N_29929);
and UO_3327 (O_3327,N_29754,N_29193);
nand UO_3328 (O_3328,N_29661,N_28527);
nand UO_3329 (O_3329,N_29722,N_28312);
nor UO_3330 (O_3330,N_29276,N_28617);
and UO_3331 (O_3331,N_29233,N_28992);
or UO_3332 (O_3332,N_29164,N_29470);
and UO_3333 (O_3333,N_29858,N_29008);
and UO_3334 (O_3334,N_28962,N_28353);
or UO_3335 (O_3335,N_28630,N_28395);
nor UO_3336 (O_3336,N_29340,N_29716);
xor UO_3337 (O_3337,N_29092,N_29210);
or UO_3338 (O_3338,N_28597,N_28627);
nand UO_3339 (O_3339,N_29357,N_28493);
or UO_3340 (O_3340,N_29809,N_29453);
nor UO_3341 (O_3341,N_28405,N_29209);
xnor UO_3342 (O_3342,N_28034,N_29389);
and UO_3343 (O_3343,N_29798,N_28984);
xor UO_3344 (O_3344,N_28670,N_29963);
nand UO_3345 (O_3345,N_29992,N_28423);
nor UO_3346 (O_3346,N_29469,N_29850);
nor UO_3347 (O_3347,N_29316,N_28165);
or UO_3348 (O_3348,N_28474,N_29994);
or UO_3349 (O_3349,N_28732,N_29639);
and UO_3350 (O_3350,N_29067,N_28724);
and UO_3351 (O_3351,N_29285,N_28479);
or UO_3352 (O_3352,N_29723,N_28368);
nand UO_3353 (O_3353,N_28672,N_29116);
or UO_3354 (O_3354,N_28743,N_28334);
or UO_3355 (O_3355,N_29822,N_29036);
or UO_3356 (O_3356,N_29723,N_29140);
nor UO_3357 (O_3357,N_29919,N_29453);
xor UO_3358 (O_3358,N_28009,N_29949);
xor UO_3359 (O_3359,N_29436,N_28221);
or UO_3360 (O_3360,N_29491,N_29197);
nor UO_3361 (O_3361,N_29089,N_28145);
xor UO_3362 (O_3362,N_28473,N_29789);
or UO_3363 (O_3363,N_28993,N_28882);
nor UO_3364 (O_3364,N_29177,N_29698);
nand UO_3365 (O_3365,N_28116,N_28886);
xor UO_3366 (O_3366,N_29310,N_29212);
nand UO_3367 (O_3367,N_28089,N_29679);
and UO_3368 (O_3368,N_29196,N_29211);
or UO_3369 (O_3369,N_29631,N_28980);
nand UO_3370 (O_3370,N_29743,N_29595);
nand UO_3371 (O_3371,N_28811,N_28798);
nand UO_3372 (O_3372,N_29037,N_29063);
nand UO_3373 (O_3373,N_28450,N_28202);
nor UO_3374 (O_3374,N_29542,N_29112);
and UO_3375 (O_3375,N_28224,N_28978);
nor UO_3376 (O_3376,N_29527,N_28401);
and UO_3377 (O_3377,N_28195,N_29328);
xnor UO_3378 (O_3378,N_29170,N_28818);
or UO_3379 (O_3379,N_28523,N_28830);
and UO_3380 (O_3380,N_29746,N_29792);
or UO_3381 (O_3381,N_28584,N_28266);
or UO_3382 (O_3382,N_29447,N_28180);
nor UO_3383 (O_3383,N_29992,N_28964);
nand UO_3384 (O_3384,N_29798,N_29219);
nand UO_3385 (O_3385,N_28613,N_29951);
nand UO_3386 (O_3386,N_28806,N_29698);
xnor UO_3387 (O_3387,N_28869,N_29942);
and UO_3388 (O_3388,N_29997,N_29332);
nand UO_3389 (O_3389,N_29003,N_29981);
nand UO_3390 (O_3390,N_28010,N_28383);
nand UO_3391 (O_3391,N_28795,N_28533);
xnor UO_3392 (O_3392,N_29078,N_29617);
and UO_3393 (O_3393,N_29778,N_29502);
nand UO_3394 (O_3394,N_28836,N_28081);
nor UO_3395 (O_3395,N_29533,N_29329);
or UO_3396 (O_3396,N_28596,N_29606);
nor UO_3397 (O_3397,N_28219,N_28772);
or UO_3398 (O_3398,N_28923,N_29941);
nor UO_3399 (O_3399,N_28864,N_28241);
nand UO_3400 (O_3400,N_29774,N_29570);
or UO_3401 (O_3401,N_28575,N_29321);
or UO_3402 (O_3402,N_28617,N_29184);
or UO_3403 (O_3403,N_29760,N_28619);
nand UO_3404 (O_3404,N_29592,N_28372);
nand UO_3405 (O_3405,N_28241,N_28517);
xor UO_3406 (O_3406,N_29538,N_29374);
and UO_3407 (O_3407,N_28780,N_28927);
nor UO_3408 (O_3408,N_28817,N_28695);
and UO_3409 (O_3409,N_29647,N_29024);
nand UO_3410 (O_3410,N_29989,N_29577);
nand UO_3411 (O_3411,N_29970,N_28735);
and UO_3412 (O_3412,N_29722,N_28210);
or UO_3413 (O_3413,N_29266,N_28362);
nand UO_3414 (O_3414,N_28897,N_29068);
or UO_3415 (O_3415,N_28215,N_28415);
and UO_3416 (O_3416,N_29261,N_28851);
or UO_3417 (O_3417,N_28214,N_29286);
nor UO_3418 (O_3418,N_29399,N_29973);
nand UO_3419 (O_3419,N_29722,N_28673);
or UO_3420 (O_3420,N_28231,N_29630);
xor UO_3421 (O_3421,N_28211,N_29889);
xnor UO_3422 (O_3422,N_28335,N_28971);
nor UO_3423 (O_3423,N_29596,N_29641);
and UO_3424 (O_3424,N_28209,N_29499);
and UO_3425 (O_3425,N_29632,N_28314);
nand UO_3426 (O_3426,N_28462,N_28384);
xnor UO_3427 (O_3427,N_28888,N_29933);
nand UO_3428 (O_3428,N_29897,N_29880);
nor UO_3429 (O_3429,N_28367,N_29984);
or UO_3430 (O_3430,N_29895,N_28462);
or UO_3431 (O_3431,N_28723,N_29936);
or UO_3432 (O_3432,N_29061,N_29005);
nand UO_3433 (O_3433,N_28811,N_28009);
nor UO_3434 (O_3434,N_28992,N_28562);
and UO_3435 (O_3435,N_29483,N_29293);
xnor UO_3436 (O_3436,N_28065,N_28459);
or UO_3437 (O_3437,N_29810,N_29244);
and UO_3438 (O_3438,N_29923,N_29818);
or UO_3439 (O_3439,N_29727,N_28564);
and UO_3440 (O_3440,N_28732,N_28069);
nor UO_3441 (O_3441,N_29350,N_28102);
nand UO_3442 (O_3442,N_29317,N_28711);
nor UO_3443 (O_3443,N_28285,N_29232);
xor UO_3444 (O_3444,N_28972,N_28138);
xnor UO_3445 (O_3445,N_28854,N_28383);
xor UO_3446 (O_3446,N_28699,N_29806);
or UO_3447 (O_3447,N_28241,N_28026);
xor UO_3448 (O_3448,N_28263,N_29422);
nand UO_3449 (O_3449,N_28693,N_28354);
xnor UO_3450 (O_3450,N_28394,N_28213);
xnor UO_3451 (O_3451,N_28547,N_28852);
and UO_3452 (O_3452,N_28389,N_28755);
xnor UO_3453 (O_3453,N_29448,N_29150);
xor UO_3454 (O_3454,N_29803,N_29593);
and UO_3455 (O_3455,N_28747,N_28129);
or UO_3456 (O_3456,N_28657,N_28549);
and UO_3457 (O_3457,N_28918,N_28928);
or UO_3458 (O_3458,N_29872,N_29921);
and UO_3459 (O_3459,N_28532,N_29101);
xor UO_3460 (O_3460,N_29474,N_28527);
or UO_3461 (O_3461,N_28771,N_29310);
and UO_3462 (O_3462,N_28140,N_28860);
nor UO_3463 (O_3463,N_29188,N_28363);
and UO_3464 (O_3464,N_29866,N_29804);
and UO_3465 (O_3465,N_28933,N_29739);
and UO_3466 (O_3466,N_29849,N_29934);
xor UO_3467 (O_3467,N_29733,N_29744);
nor UO_3468 (O_3468,N_28118,N_29342);
xnor UO_3469 (O_3469,N_28182,N_28528);
nor UO_3470 (O_3470,N_28205,N_28107);
and UO_3471 (O_3471,N_28972,N_28353);
nor UO_3472 (O_3472,N_29520,N_28258);
nor UO_3473 (O_3473,N_29200,N_28905);
or UO_3474 (O_3474,N_29412,N_28756);
xor UO_3475 (O_3475,N_29225,N_28262);
nor UO_3476 (O_3476,N_28103,N_28285);
and UO_3477 (O_3477,N_28143,N_29030);
nor UO_3478 (O_3478,N_29227,N_29064);
nor UO_3479 (O_3479,N_28337,N_29630);
and UO_3480 (O_3480,N_28522,N_28898);
or UO_3481 (O_3481,N_29422,N_28581);
xor UO_3482 (O_3482,N_28230,N_29106);
nor UO_3483 (O_3483,N_29251,N_29733);
nor UO_3484 (O_3484,N_29150,N_28153);
nand UO_3485 (O_3485,N_29337,N_29078);
nand UO_3486 (O_3486,N_28689,N_28135);
nand UO_3487 (O_3487,N_28397,N_29087);
or UO_3488 (O_3488,N_29985,N_28434);
xor UO_3489 (O_3489,N_28956,N_29906);
and UO_3490 (O_3490,N_29584,N_28204);
nor UO_3491 (O_3491,N_29185,N_28730);
and UO_3492 (O_3492,N_29206,N_29839);
xor UO_3493 (O_3493,N_29924,N_28106);
nand UO_3494 (O_3494,N_28769,N_28184);
or UO_3495 (O_3495,N_29414,N_28392);
and UO_3496 (O_3496,N_29059,N_29801);
xnor UO_3497 (O_3497,N_28172,N_29196);
nand UO_3498 (O_3498,N_28814,N_29986);
xnor UO_3499 (O_3499,N_28150,N_28765);
endmodule